module basic_1000_10000_1500_2_levels_5xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5003,N_5004,N_5005,N_5006,N_5007,N_5010,N_5012,N_5013,N_5015,N_5017,N_5018,N_5020,N_5022,N_5024,N_5028,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5037,N_5041,N_5042,N_5043,N_5044,N_5045,N_5047,N_5049,N_5050,N_5053,N_5055,N_5056,N_5058,N_5059,N_5060,N_5061,N_5064,N_5066,N_5067,N_5068,N_5069,N_5070,N_5074,N_5076,N_5077,N_5078,N_5079,N_5081,N_5082,N_5083,N_5084,N_5087,N_5088,N_5089,N_5090,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5106,N_5110,N_5112,N_5115,N_5116,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5126,N_5128,N_5130,N_5131,N_5132,N_5135,N_5137,N_5141,N_5143,N_5144,N_5146,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5156,N_5157,N_5158,N_5159,N_5163,N_5164,N_5167,N_5170,N_5171,N_5172,N_5175,N_5178,N_5179,N_5180,N_5182,N_5184,N_5185,N_5186,N_5188,N_5189,N_5191,N_5192,N_5193,N_5194,N_5197,N_5199,N_5200,N_5203,N_5205,N_5206,N_5207,N_5209,N_5210,N_5211,N_5214,N_5216,N_5219,N_5223,N_5226,N_5227,N_5228,N_5229,N_5232,N_5233,N_5234,N_5235,N_5236,N_5238,N_5239,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5252,N_5253,N_5254,N_5258,N_5260,N_5261,N_5263,N_5264,N_5265,N_5266,N_5267,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5278,N_5279,N_5280,N_5281,N_5283,N_5285,N_5286,N_5288,N_5289,N_5290,N_5292,N_5295,N_5297,N_5301,N_5302,N_5304,N_5305,N_5306,N_5307,N_5308,N_5310,N_5313,N_5314,N_5315,N_5316,N_5317,N_5320,N_5323,N_5325,N_5326,N_5327,N_5329,N_5330,N_5336,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5348,N_5349,N_5351,N_5352,N_5359,N_5361,N_5362,N_5364,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5386,N_5388,N_5389,N_5391,N_5392,N_5394,N_5395,N_5397,N_5398,N_5401,N_5403,N_5405,N_5408,N_5409,N_5410,N_5412,N_5413,N_5414,N_5417,N_5418,N_5419,N_5422,N_5423,N_5424,N_5425,N_5428,N_5430,N_5432,N_5434,N_5436,N_5437,N_5439,N_5441,N_5443,N_5445,N_5449,N_5451,N_5455,N_5456,N_5457,N_5458,N_5460,N_5463,N_5464,N_5466,N_5467,N_5468,N_5470,N_5471,N_5473,N_5474,N_5475,N_5477,N_5478,N_5479,N_5480,N_5481,N_5483,N_5485,N_5487,N_5490,N_5491,N_5492,N_5493,N_5496,N_5497,N_5499,N_5503,N_5505,N_5507,N_5508,N_5510,N_5511,N_5512,N_5516,N_5517,N_5520,N_5521,N_5523,N_5524,N_5526,N_5528,N_5530,N_5531,N_5534,N_5536,N_5537,N_5539,N_5541,N_5543,N_5544,N_5546,N_5547,N_5548,N_5551,N_5552,N_5553,N_5554,N_5555,N_5557,N_5559,N_5560,N_5561,N_5562,N_5563,N_5565,N_5566,N_5568,N_5570,N_5571,N_5572,N_5573,N_5574,N_5578,N_5580,N_5582,N_5583,N_5585,N_5588,N_5590,N_5593,N_5594,N_5595,N_5596,N_5597,N_5599,N_5601,N_5602,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5622,N_5623,N_5624,N_5626,N_5628,N_5629,N_5631,N_5632,N_5633,N_5634,N_5635,N_5637,N_5640,N_5641,N_5649,N_5650,N_5651,N_5652,N_5655,N_5657,N_5658,N_5659,N_5661,N_5662,N_5663,N_5664,N_5666,N_5667,N_5668,N_5673,N_5674,N_5675,N_5676,N_5677,N_5682,N_5684,N_5686,N_5689,N_5690,N_5691,N_5692,N_5693,N_5697,N_5698,N_5702,N_5704,N_5705,N_5706,N_5707,N_5710,N_5711,N_5712,N_5714,N_5717,N_5718,N_5721,N_5726,N_5728,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5739,N_5740,N_5742,N_5745,N_5746,N_5750,N_5751,N_5752,N_5754,N_5759,N_5762,N_5763,N_5764,N_5765,N_5767,N_5768,N_5769,N_5770,N_5772,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5787,N_5788,N_5790,N_5791,N_5792,N_5793,N_5795,N_5799,N_5801,N_5802,N_5803,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5817,N_5824,N_5825,N_5826,N_5830,N_5831,N_5832,N_5833,N_5836,N_5838,N_5839,N_5840,N_5841,N_5843,N_5845,N_5852,N_5854,N_5855,N_5856,N_5857,N_5863,N_5864,N_5867,N_5869,N_5870,N_5871,N_5872,N_5873,N_5875,N_5876,N_5877,N_5881,N_5882,N_5884,N_5887,N_5890,N_5892,N_5894,N_5896,N_5899,N_5900,N_5901,N_5904,N_5908,N_5909,N_5910,N_5911,N_5915,N_5917,N_5919,N_5920,N_5922,N_5923,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5934,N_5935,N_5936,N_5939,N_5940,N_5941,N_5944,N_5945,N_5948,N_5950,N_5952,N_5954,N_5955,N_5956,N_5959,N_5961,N_5962,N_5963,N_5964,N_5965,N_5969,N_5973,N_5975,N_5976,N_5978,N_5979,N_5981,N_5985,N_5986,N_5987,N_5988,N_5990,N_5991,N_5993,N_5994,N_5996,N_5998,N_5999,N_6000,N_6001,N_6005,N_6006,N_6008,N_6010,N_6011,N_6012,N_6013,N_6016,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6030,N_6035,N_6036,N_6040,N_6041,N_6043,N_6044,N_6045,N_6047,N_6049,N_6053,N_6055,N_6056,N_6058,N_6059,N_6060,N_6062,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6076,N_6077,N_6078,N_6080,N_6081,N_6082,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6094,N_6097,N_6100,N_6101,N_6103,N_6104,N_6105,N_6106,N_6109,N_6112,N_6113,N_6114,N_6115,N_6116,N_6119,N_6120,N_6123,N_6124,N_6126,N_6128,N_6130,N_6132,N_6133,N_6136,N_6138,N_6141,N_6144,N_6147,N_6148,N_6149,N_6150,N_6153,N_6154,N_6155,N_6156,N_6157,N_6159,N_6164,N_6165,N_6166,N_6167,N_6168,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6179,N_6181,N_6187,N_6188,N_6191,N_6193,N_6195,N_6197,N_6198,N_6200,N_6203,N_6204,N_6205,N_6207,N_6209,N_6210,N_6212,N_6214,N_6215,N_6216,N_6221,N_6224,N_6225,N_6228,N_6229,N_6230,N_6231,N_6232,N_6235,N_6236,N_6238,N_6239,N_6240,N_6245,N_6246,N_6248,N_6249,N_6251,N_6252,N_6253,N_6254,N_6255,N_6257,N_6261,N_6265,N_6267,N_6269,N_6275,N_6276,N_6279,N_6280,N_6281,N_6282,N_6284,N_6285,N_6286,N_6287,N_6289,N_6291,N_6293,N_6294,N_6295,N_6296,N_6297,N_6299,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6310,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6319,N_6320,N_6321,N_6322,N_6323,N_6325,N_6327,N_6328,N_6330,N_6332,N_6333,N_6335,N_6336,N_6338,N_6340,N_6341,N_6342,N_6343,N_6346,N_6347,N_6348,N_6349,N_6350,N_6352,N_6353,N_6354,N_6361,N_6362,N_6363,N_6365,N_6366,N_6367,N_6371,N_6372,N_6373,N_6375,N_6376,N_6378,N_6379,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6389,N_6392,N_6394,N_6395,N_6396,N_6397,N_6399,N_6401,N_6402,N_6403,N_6404,N_6406,N_6407,N_6408,N_6410,N_6412,N_6414,N_6416,N_6418,N_6419,N_6420,N_6422,N_6423,N_6426,N_6429,N_6430,N_6431,N_6433,N_6439,N_6442,N_6443,N_6446,N_6448,N_6451,N_6452,N_6456,N_6457,N_6459,N_6460,N_6463,N_6465,N_6466,N_6467,N_6469,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6493,N_6495,N_6497,N_6498,N_6500,N_6501,N_6503,N_6504,N_6507,N_6508,N_6509,N_6510,N_6512,N_6513,N_6514,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6527,N_6528,N_6530,N_6531,N_6532,N_6537,N_6538,N_6539,N_6540,N_6542,N_6543,N_6545,N_6547,N_6549,N_6550,N_6552,N_6553,N_6554,N_6557,N_6558,N_6559,N_6561,N_6562,N_6563,N_6565,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6580,N_6582,N_6583,N_6584,N_6586,N_6588,N_6589,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6601,N_6603,N_6605,N_6606,N_6607,N_6608,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6621,N_6623,N_6624,N_6625,N_6626,N_6629,N_6632,N_6635,N_6638,N_6639,N_6644,N_6645,N_6646,N_6648,N_6650,N_6651,N_6653,N_6654,N_6656,N_6658,N_6661,N_6662,N_6663,N_6665,N_6666,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6677,N_6681,N_6684,N_6685,N_6688,N_6689,N_6690,N_6692,N_6694,N_6695,N_6696,N_6698,N_6699,N_6700,N_6703,N_6704,N_6705,N_6706,N_6708,N_6710,N_6712,N_6715,N_6716,N_6718,N_6719,N_6720,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6737,N_6738,N_6739,N_6740,N_6741,N_6746,N_6747,N_6748,N_6751,N_6754,N_6756,N_6759,N_6760,N_6761,N_6762,N_6764,N_6765,N_6766,N_6767,N_6770,N_6771,N_6772,N_6778,N_6780,N_6782,N_6785,N_6787,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6800,N_6801,N_6802,N_6805,N_6806,N_6807,N_6808,N_6811,N_6812,N_6814,N_6816,N_6817,N_6818,N_6819,N_6821,N_6822,N_6827,N_6828,N_6831,N_6834,N_6835,N_6836,N_6837,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6854,N_6855,N_6856,N_6860,N_6863,N_6867,N_6868,N_6869,N_6870,N_6872,N_6875,N_6877,N_6878,N_6879,N_6883,N_6884,N_6885,N_6888,N_6889,N_6891,N_6893,N_6895,N_6896,N_6897,N_6898,N_6900,N_6903,N_6904,N_6907,N_6908,N_6909,N_6911,N_6914,N_6915,N_6918,N_6919,N_6920,N_6922,N_6925,N_6926,N_6927,N_6928,N_6930,N_6931,N_6933,N_6934,N_6936,N_6938,N_6939,N_6940,N_6941,N_6946,N_6947,N_6948,N_6950,N_6952,N_6953,N_6954,N_6955,N_6956,N_6959,N_6960,N_6964,N_6965,N_6966,N_6968,N_6969,N_6970,N_6976,N_6978,N_6979,N_6981,N_6983,N_6986,N_6987,N_6989,N_6991,N_6994,N_6995,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7006,N_7007,N_7009,N_7010,N_7012,N_7014,N_7015,N_7016,N_7017,N_7019,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7029,N_7030,N_7031,N_7032,N_7036,N_7038,N_7040,N_7041,N_7043,N_7044,N_7046,N_7048,N_7051,N_7055,N_7057,N_7058,N_7059,N_7061,N_7066,N_7067,N_7072,N_7073,N_7076,N_7079,N_7082,N_7083,N_7084,N_7086,N_7088,N_7089,N_7090,N_7091,N_7093,N_7097,N_7099,N_7100,N_7101,N_7102,N_7103,N_7105,N_7106,N_7107,N_7108,N_7109,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7121,N_7122,N_7126,N_7129,N_7130,N_7132,N_7135,N_7137,N_7138,N_7139,N_7140,N_7141,N_7144,N_7147,N_7148,N_7149,N_7150,N_7151,N_7153,N_7154,N_7156,N_7159,N_7160,N_7161,N_7165,N_7166,N_7169,N_7170,N_7174,N_7177,N_7178,N_7179,N_7180,N_7182,N_7184,N_7185,N_7186,N_7187,N_7190,N_7191,N_7194,N_7197,N_7201,N_7202,N_7204,N_7206,N_7207,N_7208,N_7210,N_7211,N_7212,N_7214,N_7216,N_7217,N_7218,N_7220,N_7221,N_7223,N_7225,N_7227,N_7228,N_7232,N_7233,N_7235,N_7237,N_7238,N_7239,N_7240,N_7242,N_7243,N_7248,N_7249,N_7250,N_7252,N_7253,N_7254,N_7255,N_7257,N_7258,N_7260,N_7261,N_7263,N_7265,N_7267,N_7271,N_7277,N_7278,N_7279,N_7280,N_7282,N_7283,N_7284,N_7286,N_7288,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7301,N_7302,N_7304,N_7306,N_7307,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7316,N_7317,N_7318,N_7319,N_7323,N_7324,N_7327,N_7329,N_7330,N_7331,N_7333,N_7334,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7348,N_7350,N_7352,N_7353,N_7359,N_7360,N_7362,N_7364,N_7365,N_7366,N_7367,N_7368,N_7373,N_7374,N_7375,N_7376,N_7379,N_7381,N_7383,N_7386,N_7395,N_7398,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7412,N_7414,N_7415,N_7416,N_7418,N_7419,N_7428,N_7431,N_7432,N_7433,N_7434,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7448,N_7449,N_7452,N_7453,N_7454,N_7456,N_7457,N_7458,N_7463,N_7464,N_7467,N_7468,N_7473,N_7475,N_7476,N_7477,N_7482,N_7483,N_7484,N_7486,N_7488,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7498,N_7499,N_7501,N_7503,N_7504,N_7505,N_7506,N_7507,N_7509,N_7510,N_7511,N_7512,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7522,N_7524,N_7527,N_7528,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7538,N_7539,N_7540,N_7541,N_7542,N_7544,N_7546,N_7547,N_7548,N_7549,N_7551,N_7552,N_7553,N_7554,N_7556,N_7559,N_7560,N_7564,N_7565,N_7566,N_7568,N_7569,N_7572,N_7573,N_7574,N_7575,N_7577,N_7578,N_7580,N_7581,N_7583,N_7584,N_7585,N_7587,N_7588,N_7589,N_7590,N_7591,N_7593,N_7598,N_7599,N_7600,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7616,N_7619,N_7620,N_7623,N_7624,N_7626,N_7627,N_7630,N_7633,N_7636,N_7637,N_7640,N_7641,N_7643,N_7644,N_7647,N_7648,N_7649,N_7651,N_7652,N_7654,N_7656,N_7657,N_7660,N_7661,N_7662,N_7663,N_7666,N_7667,N_7668,N_7671,N_7673,N_7677,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7689,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7712,N_7713,N_7714,N_7716,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7728,N_7729,N_7731,N_7732,N_7736,N_7737,N_7738,N_7739,N_7740,N_7742,N_7745,N_7749,N_7751,N_7752,N_7753,N_7754,N_7755,N_7757,N_7758,N_7759,N_7760,N_7763,N_7764,N_7767,N_7769,N_7771,N_7774,N_7775,N_7776,N_7781,N_7782,N_7783,N_7785,N_7786,N_7787,N_7788,N_7790,N_7794,N_7796,N_7799,N_7802,N_7803,N_7806,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7816,N_7820,N_7821,N_7822,N_7823,N_7825,N_7826,N_7828,N_7829,N_7830,N_7832,N_7838,N_7841,N_7842,N_7843,N_7845,N_7846,N_7848,N_7850,N_7851,N_7854,N_7856,N_7857,N_7859,N_7861,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7876,N_7878,N_7879,N_7880,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7901,N_7902,N_7904,N_7907,N_7908,N_7910,N_7911,N_7912,N_7913,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7924,N_7925,N_7927,N_7929,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7939,N_7940,N_7944,N_7945,N_7947,N_7950,N_7951,N_7952,N_7954,N_7955,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7968,N_7969,N_7970,N_7972,N_7974,N_7977,N_7980,N_7981,N_7983,N_7986,N_7987,N_7989,N_7991,N_7992,N_7993,N_7994,N_7997,N_8000,N_8001,N_8002,N_8004,N_8006,N_8009,N_8010,N_8012,N_8013,N_8016,N_8017,N_8019,N_8020,N_8021,N_8022,N_8027,N_8029,N_8031,N_8037,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8056,N_8059,N_8064,N_8066,N_8067,N_8068,N_8070,N_8071,N_8072,N_8074,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8087,N_8088,N_8090,N_8093,N_8096,N_8097,N_8098,N_8099,N_8101,N_8104,N_8105,N_8106,N_8107,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8117,N_8119,N_8120,N_8121,N_8122,N_8126,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8135,N_8136,N_8137,N_8139,N_8143,N_8146,N_8147,N_8148,N_8152,N_8153,N_8154,N_8156,N_8158,N_8159,N_8161,N_8163,N_8165,N_8166,N_8168,N_8172,N_8173,N_8176,N_8178,N_8181,N_8182,N_8183,N_8184,N_8185,N_8187,N_8190,N_8192,N_8193,N_8195,N_8197,N_8198,N_8200,N_8203,N_8204,N_8206,N_8210,N_8212,N_8213,N_8214,N_8215,N_8217,N_8218,N_8219,N_8221,N_8223,N_8226,N_8228,N_8229,N_8231,N_8232,N_8235,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8254,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8265,N_8269,N_8271,N_8272,N_8274,N_8275,N_8276,N_8279,N_8281,N_8285,N_8286,N_8287,N_8288,N_8290,N_8292,N_8297,N_8299,N_8300,N_8301,N_8302,N_8303,N_8305,N_8306,N_8307,N_8312,N_8313,N_8316,N_8320,N_8321,N_8322,N_8323,N_8324,N_8326,N_8327,N_8328,N_8329,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8341,N_8343,N_8345,N_8347,N_8351,N_8353,N_8354,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8364,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8389,N_8390,N_8392,N_8393,N_8394,N_8395,N_8397,N_8399,N_8401,N_8402,N_8403,N_8405,N_8407,N_8408,N_8411,N_8413,N_8414,N_8415,N_8417,N_8418,N_8420,N_8423,N_8426,N_8428,N_8429,N_8430,N_8435,N_8438,N_8439,N_8442,N_8444,N_8445,N_8446,N_8448,N_8449,N_8451,N_8452,N_8453,N_8457,N_8458,N_8459,N_8460,N_8463,N_8464,N_8466,N_8467,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8478,N_8482,N_8488,N_8489,N_8490,N_8492,N_8493,N_8495,N_8496,N_8499,N_8500,N_8501,N_8502,N_8503,N_8508,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8520,N_8522,N_8523,N_8524,N_8525,N_8527,N_8533,N_8534,N_8535,N_8536,N_8538,N_8539,N_8540,N_8541,N_8544,N_8545,N_8546,N_8548,N_8552,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8563,N_8565,N_8566,N_8567,N_8569,N_8570,N_8571,N_8572,N_8575,N_8578,N_8581,N_8582,N_8584,N_8585,N_8588,N_8589,N_8591,N_8592,N_8593,N_8594,N_8595,N_8597,N_8598,N_8599,N_8600,N_8601,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8613,N_8615,N_8617,N_8618,N_8619,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8637,N_8638,N_8641,N_8642,N_8645,N_8646,N_8647,N_8649,N_8650,N_8652,N_8653,N_8654,N_8659,N_8660,N_8662,N_8663,N_8665,N_8667,N_8669,N_8670,N_8672,N_8673,N_8674,N_8675,N_8677,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8688,N_8689,N_8691,N_8693,N_8694,N_8695,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8705,N_8706,N_8707,N_8709,N_8710,N_8712,N_8716,N_8719,N_8721,N_8723,N_8725,N_8727,N_8728,N_8729,N_8730,N_8732,N_8733,N_8734,N_8735,N_8737,N_8738,N_8739,N_8743,N_8744,N_8745,N_8747,N_8748,N_8750,N_8751,N_8752,N_8753,N_8754,N_8758,N_8759,N_8761,N_8762,N_8763,N_8764,N_8765,N_8767,N_8768,N_8770,N_8772,N_8778,N_8779,N_8781,N_8782,N_8784,N_8785,N_8786,N_8789,N_8790,N_8791,N_8792,N_8793,N_8795,N_8796,N_8801,N_8803,N_8805,N_8806,N_8808,N_8810,N_8811,N_8812,N_8814,N_8815,N_8816,N_8817,N_8819,N_8820,N_8822,N_8823,N_8824,N_8826,N_8827,N_8828,N_8829,N_8831,N_8833,N_8834,N_8835,N_8836,N_8839,N_8840,N_8841,N_8842,N_8844,N_8845,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8855,N_8857,N_8859,N_8861,N_8862,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8872,N_8874,N_8875,N_8878,N_8879,N_8880,N_8882,N_8883,N_8885,N_8886,N_8887,N_8888,N_8891,N_8892,N_8893,N_8897,N_8898,N_8899,N_8900,N_8901,N_8904,N_8911,N_8914,N_8915,N_8917,N_8918,N_8919,N_8921,N_8922,N_8923,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8939,N_8941,N_8942,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8953,N_8954,N_8958,N_8960,N_8962,N_8963,N_8964,N_8966,N_8967,N_8970,N_8971,N_8972,N_8975,N_8977,N_8979,N_8980,N_8982,N_8984,N_8986,N_8987,N_8990,N_8991,N_8993,N_8994,N_8996,N_8998,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9020,N_9022,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9036,N_9039,N_9041,N_9042,N_9046,N_9047,N_9048,N_9049,N_9050,N_9052,N_9054,N_9055,N_9057,N_9058,N_9061,N_9062,N_9065,N_9066,N_9068,N_9069,N_9070,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9081,N_9082,N_9084,N_9087,N_9088,N_9096,N_9097,N_9098,N_9101,N_9102,N_9105,N_9107,N_9108,N_9109,N_9110,N_9112,N_9114,N_9116,N_9117,N_9118,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9131,N_9133,N_9136,N_9137,N_9138,N_9140,N_9141,N_9142,N_9144,N_9149,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9160,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9173,N_9174,N_9176,N_9177,N_9179,N_9181,N_9182,N_9183,N_9185,N_9190,N_9191,N_9192,N_9194,N_9196,N_9199,N_9200,N_9201,N_9202,N_9203,N_9205,N_9207,N_9208,N_9209,N_9210,N_9212,N_9213,N_9214,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9225,N_9226,N_9230,N_9231,N_9232,N_9233,N_9234,N_9236,N_9237,N_9238,N_9241,N_9242,N_9243,N_9244,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9253,N_9256,N_9257,N_9260,N_9264,N_9266,N_9267,N_9268,N_9271,N_9273,N_9274,N_9276,N_9277,N_9278,N_9279,N_9280,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9309,N_9311,N_9312,N_9313,N_9315,N_9321,N_9322,N_9324,N_9327,N_9328,N_9329,N_9330,N_9332,N_9333,N_9334,N_9338,N_9339,N_9340,N_9341,N_9342,N_9344,N_9345,N_9346,N_9347,N_9349,N_9353,N_9354,N_9355,N_9356,N_9359,N_9361,N_9365,N_9366,N_9368,N_9369,N_9370,N_9371,N_9373,N_9375,N_9376,N_9377,N_9379,N_9380,N_9382,N_9383,N_9386,N_9387,N_9388,N_9389,N_9394,N_9395,N_9398,N_9400,N_9402,N_9403,N_9405,N_9406,N_9407,N_9408,N_9409,N_9411,N_9414,N_9415,N_9417,N_9418,N_9420,N_9422,N_9423,N_9424,N_9425,N_9431,N_9432,N_9435,N_9437,N_9440,N_9443,N_9444,N_9445,N_9447,N_9448,N_9449,N_9452,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9464,N_9465,N_9466,N_9470,N_9471,N_9476,N_9477,N_9479,N_9480,N_9483,N_9484,N_9487,N_9489,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9502,N_9503,N_9504,N_9505,N_9506,N_9508,N_9509,N_9510,N_9511,N_9512,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9525,N_9528,N_9529,N_9530,N_9531,N_9533,N_9535,N_9537,N_9538,N_9539,N_9541,N_9543,N_9544,N_9547,N_9549,N_9550,N_9551,N_9552,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9561,N_9562,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9572,N_9576,N_9579,N_9581,N_9582,N_9584,N_9585,N_9586,N_9588,N_9593,N_9594,N_9595,N_9596,N_9597,N_9599,N_9600,N_9601,N_9602,N_9604,N_9605,N_9607,N_9608,N_9609,N_9612,N_9616,N_9617,N_9618,N_9619,N_9624,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9637,N_9638,N_9645,N_9646,N_9648,N_9650,N_9651,N_9654,N_9655,N_9656,N_9658,N_9660,N_9663,N_9668,N_9669,N_9672,N_9673,N_9674,N_9675,N_9677,N_9680,N_9681,N_9682,N_9684,N_9685,N_9686,N_9687,N_9688,N_9690,N_9692,N_9695,N_9699,N_9700,N_9701,N_9705,N_9706,N_9707,N_9708,N_9711,N_9712,N_9714,N_9715,N_9719,N_9723,N_9726,N_9727,N_9728,N_9729,N_9732,N_9733,N_9734,N_9735,N_9738,N_9740,N_9744,N_9745,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9756,N_9759,N_9760,N_9761,N_9765,N_9769,N_9770,N_9772,N_9774,N_9775,N_9776,N_9777,N_9779,N_9782,N_9783,N_9787,N_9788,N_9789,N_9790,N_9793,N_9794,N_9796,N_9797,N_9799,N_9805,N_9807,N_9809,N_9812,N_9813,N_9814,N_9815,N_9818,N_9819,N_9821,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9830,N_9832,N_9833,N_9835,N_9836,N_9838,N_9842,N_9843,N_9846,N_9847,N_9849,N_9852,N_9853,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9874,N_9875,N_9877,N_9879,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9890,N_9891,N_9892,N_9893,N_9896,N_9899,N_9900,N_9901,N_9902,N_9904,N_9906,N_9907,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9917,N_9920,N_9921,N_9925,N_9927,N_9928,N_9932,N_9935,N_9936,N_9937,N_9942,N_9943,N_9946,N_9947,N_9950,N_9951,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9961,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9972,N_9978,N_9979,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9999;
and U0 (N_0,In_412,In_671);
nand U1 (N_1,In_599,In_13);
xor U2 (N_2,In_369,In_908);
nor U3 (N_3,In_613,In_745);
nor U4 (N_4,In_674,In_27);
and U5 (N_5,In_500,In_359);
and U6 (N_6,In_151,In_646);
nor U7 (N_7,In_969,In_382);
nor U8 (N_8,In_538,In_300);
or U9 (N_9,In_329,In_708);
nor U10 (N_10,In_25,In_129);
xnor U11 (N_11,In_233,In_666);
or U12 (N_12,In_951,In_784);
and U13 (N_13,In_462,In_918);
xnor U14 (N_14,In_79,In_58);
nand U15 (N_15,In_688,In_477);
or U16 (N_16,In_935,In_832);
or U17 (N_17,In_324,In_450);
and U18 (N_18,In_746,In_710);
nand U19 (N_19,In_361,In_545);
xnor U20 (N_20,In_384,In_120);
xnor U21 (N_21,In_160,In_882);
or U22 (N_22,In_636,In_608);
nor U23 (N_23,In_568,In_611);
nand U24 (N_24,In_252,In_258);
and U25 (N_25,In_958,In_749);
nand U26 (N_26,In_442,In_215);
xor U27 (N_27,In_291,In_730);
nor U28 (N_28,In_108,In_839);
or U29 (N_29,In_93,In_288);
nand U30 (N_30,In_266,In_53);
xor U31 (N_31,In_530,In_645);
and U32 (N_32,In_718,In_897);
xnor U33 (N_33,In_584,In_470);
nand U34 (N_34,In_85,In_473);
nand U35 (N_35,In_837,In_242);
nor U36 (N_36,In_536,In_325);
nand U37 (N_37,In_446,In_320);
or U38 (N_38,In_961,In_142);
nand U39 (N_39,In_657,In_10);
and U40 (N_40,In_949,In_181);
or U41 (N_41,In_474,In_321);
nor U42 (N_42,In_720,In_368);
nor U43 (N_43,In_133,In_979);
xor U44 (N_44,In_743,In_587);
or U45 (N_45,In_654,In_457);
and U46 (N_46,In_63,In_676);
nor U47 (N_47,In_183,In_427);
nand U48 (N_48,In_344,In_930);
and U49 (N_49,In_943,In_413);
or U50 (N_50,In_261,In_356);
nor U51 (N_51,In_993,In_658);
nor U52 (N_52,In_747,In_48);
or U53 (N_53,In_39,In_857);
nand U54 (N_54,In_307,In_762);
and U55 (N_55,In_892,In_317);
nand U56 (N_56,In_206,In_402);
and U57 (N_57,In_728,In_460);
and U58 (N_58,In_420,In_647);
nor U59 (N_59,In_377,In_773);
nand U60 (N_60,In_804,In_813);
and U61 (N_61,In_737,In_879);
and U62 (N_62,In_526,In_744);
nand U63 (N_63,In_95,In_973);
nand U64 (N_64,In_861,In_4);
or U65 (N_65,In_899,In_630);
nand U66 (N_66,In_455,In_148);
nor U67 (N_67,In_945,In_727);
nor U68 (N_68,In_328,In_189);
nor U69 (N_69,In_337,In_692);
or U70 (N_70,In_884,In_724);
nor U71 (N_71,In_370,In_209);
nand U72 (N_72,In_953,In_162);
or U73 (N_73,In_509,In_916);
nand U74 (N_74,In_229,In_130);
and U75 (N_75,In_56,In_546);
and U76 (N_76,In_612,In_807);
nor U77 (N_77,In_865,In_137);
nor U78 (N_78,In_253,In_498);
nor U79 (N_79,In_572,In_482);
and U80 (N_80,In_83,In_964);
and U81 (N_81,In_158,In_302);
nand U82 (N_82,In_939,In_34);
and U83 (N_83,In_553,In_684);
nor U84 (N_84,In_641,In_136);
xor U85 (N_85,In_214,In_277);
nor U86 (N_86,In_962,In_991);
nor U87 (N_87,In_924,In_234);
nand U88 (N_88,In_6,In_703);
and U89 (N_89,In_904,In_776);
nand U90 (N_90,In_533,In_101);
and U91 (N_91,In_7,In_115);
xnor U92 (N_92,In_535,In_902);
xor U93 (N_93,In_15,In_583);
or U94 (N_94,In_581,In_281);
or U95 (N_95,In_673,In_187);
and U96 (N_96,In_208,In_319);
nand U97 (N_97,In_419,In_168);
nor U98 (N_98,In_268,In_850);
and U99 (N_99,In_686,In_704);
and U100 (N_100,In_653,In_367);
and U101 (N_101,In_540,In_487);
nor U102 (N_102,In_390,In_920);
nor U103 (N_103,In_371,In_393);
nand U104 (N_104,In_542,In_826);
or U105 (N_105,In_348,In_515);
nor U106 (N_106,In_503,In_18);
nand U107 (N_107,In_984,In_520);
nor U108 (N_108,In_228,In_912);
and U109 (N_109,In_527,In_875);
and U110 (N_110,In_995,In_311);
nand U111 (N_111,In_171,In_981);
or U112 (N_112,In_250,In_810);
and U113 (N_113,In_997,In_65);
xnor U114 (N_114,In_247,In_489);
nand U115 (N_115,In_105,In_788);
or U116 (N_116,In_852,In_550);
or U117 (N_117,In_580,In_680);
nor U118 (N_118,In_989,In_764);
nand U119 (N_119,In_855,In_28);
nand U120 (N_120,In_428,In_407);
or U121 (N_121,In_761,In_597);
nand U122 (N_122,In_833,In_92);
nand U123 (N_123,In_511,In_824);
or U124 (N_124,In_483,In_605);
or U125 (N_125,In_663,In_971);
nor U126 (N_126,In_591,In_600);
nand U127 (N_127,In_598,In_615);
and U128 (N_128,In_575,In_135);
xnor U129 (N_129,In_80,In_327);
xnor U130 (N_130,In_774,In_47);
or U131 (N_131,In_225,In_458);
and U132 (N_132,In_99,In_456);
or U133 (N_133,In_29,In_604);
and U134 (N_134,In_614,In_903);
nand U135 (N_135,In_888,In_845);
nand U136 (N_136,In_705,In_346);
and U137 (N_137,In_38,In_116);
nor U138 (N_138,In_891,In_765);
and U139 (N_139,In_400,In_878);
nor U140 (N_140,In_563,In_691);
and U141 (N_141,In_73,In_808);
and U142 (N_142,In_484,In_687);
and U143 (N_143,In_508,In_119);
nor U144 (N_144,In_131,In_632);
xnor U145 (N_145,In_987,In_436);
or U146 (N_146,In_738,In_312);
nor U147 (N_147,In_310,In_132);
nor U148 (N_148,In_635,In_957);
nand U149 (N_149,In_947,In_640);
and U150 (N_150,In_213,In_403);
or U151 (N_151,In_146,In_629);
and U152 (N_152,In_618,In_244);
xor U153 (N_153,In_585,In_357);
or U154 (N_154,In_841,In_224);
nor U155 (N_155,In_510,In_349);
xnor U156 (N_156,In_634,In_795);
or U157 (N_157,In_925,In_860);
nor U158 (N_158,In_143,In_755);
or U159 (N_159,In_998,In_862);
xnor U160 (N_160,In_933,In_111);
and U161 (N_161,In_670,In_256);
nor U162 (N_162,In_192,In_603);
nor U163 (N_163,In_24,In_323);
or U164 (N_164,In_164,In_851);
xor U165 (N_165,In_278,In_496);
xnor U166 (N_166,In_104,In_528);
and U167 (N_167,In_651,In_820);
nand U168 (N_168,In_78,In_923);
or U169 (N_169,In_975,In_492);
and U170 (N_170,In_926,In_963);
nor U171 (N_171,In_98,In_523);
or U172 (N_172,In_96,In_609);
xnor U173 (N_173,In_351,In_524);
nor U174 (N_174,In_990,In_153);
or U175 (N_175,In_955,In_309);
nor U176 (N_176,In_594,In_731);
and U177 (N_177,In_552,In_89);
nand U178 (N_178,In_842,In_70);
nor U179 (N_179,In_699,In_395);
nor U180 (N_180,In_453,In_757);
or U181 (N_181,In_828,In_922);
nor U182 (N_182,In_952,In_376);
and U183 (N_183,In_184,In_260);
nor U184 (N_184,In_946,In_801);
nor U185 (N_185,In_700,In_942);
nor U186 (N_186,In_831,In_434);
nor U187 (N_187,In_55,In_114);
or U188 (N_188,In_775,In_199);
or U189 (N_189,In_194,In_766);
and U190 (N_190,In_937,In_426);
nand U191 (N_191,In_54,In_235);
or U192 (N_192,In_112,In_280);
nand U193 (N_193,In_976,In_358);
or U194 (N_194,In_227,In_960);
nor U195 (N_195,In_205,In_306);
or U196 (N_196,In_562,In_631);
nand U197 (N_197,In_154,In_799);
and U198 (N_198,In_974,In_313);
nor U199 (N_199,In_432,In_293);
nand U200 (N_200,In_0,In_607);
nand U201 (N_201,In_849,In_725);
and U202 (N_202,In_733,In_781);
nor U203 (N_203,In_64,In_415);
or U204 (N_204,In_966,In_404);
and U205 (N_205,In_431,In_558);
and U206 (N_206,In_777,In_433);
nor U207 (N_207,In_372,In_188);
or U208 (N_208,In_829,In_23);
xor U209 (N_209,In_988,In_672);
or U210 (N_210,In_863,In_398);
xor U211 (N_211,In_32,In_785);
and U212 (N_212,In_203,In_163);
nor U213 (N_213,In_621,In_463);
or U214 (N_214,In_620,In_2);
nand U215 (N_215,In_238,In_493);
nor U216 (N_216,In_571,In_914);
nor U217 (N_217,In_502,In_573);
xor U218 (N_218,In_771,In_790);
nor U219 (N_219,In_195,In_986);
nand U220 (N_220,In_475,In_996);
nor U221 (N_221,In_868,In_134);
nor U222 (N_222,In_396,In_147);
or U223 (N_223,In_342,In_161);
or U224 (N_224,In_123,In_514);
nor U225 (N_225,In_566,In_994);
nand U226 (N_226,In_299,In_251);
xnor U227 (N_227,In_289,In_409);
or U228 (N_228,In_797,In_140);
and U229 (N_229,In_938,In_648);
nor U230 (N_230,In_144,In_532);
and U231 (N_231,In_716,In_956);
xnor U232 (N_232,In_876,In_735);
nand U233 (N_233,In_275,In_665);
and U234 (N_234,In_72,In_249);
nand U235 (N_235,In_117,In_90);
nand U236 (N_236,In_816,In_362);
and U237 (N_237,In_50,In_669);
or U238 (N_238,In_221,In_14);
nand U239 (N_239,In_754,In_750);
nor U240 (N_240,In_282,In_240);
and U241 (N_241,In_847,In_274);
nand U242 (N_242,In_838,In_819);
and U243 (N_243,In_723,In_341);
and U244 (N_244,In_675,In_86);
or U245 (N_245,In_459,In_805);
or U246 (N_246,In_363,In_410);
or U247 (N_247,In_165,In_698);
nor U248 (N_248,In_959,In_223);
nand U249 (N_249,In_896,In_389);
or U250 (N_250,In_732,In_20);
and U251 (N_251,In_338,In_157);
nand U252 (N_252,In_992,In_439);
and U253 (N_253,In_3,In_272);
xor U254 (N_254,In_210,In_791);
and U255 (N_255,In_919,In_21);
nor U256 (N_256,In_308,In_36);
or U257 (N_257,In_318,In_736);
and U258 (N_258,In_68,In_506);
nor U259 (N_259,In_980,In_139);
nand U260 (N_260,In_292,In_169);
nand U261 (N_261,In_619,In_531);
nand U262 (N_262,In_331,In_574);
nor U263 (N_263,In_786,In_52);
nor U264 (N_264,In_555,In_950);
or U265 (N_265,In_217,In_355);
nor U266 (N_266,In_471,In_373);
nor U267 (N_267,In_602,In_548);
nor U268 (N_268,In_889,In_915);
nand U269 (N_269,In_353,In_35);
nand U270 (N_270,In_122,In_516);
nand U271 (N_271,In_917,In_37);
nand U272 (N_272,In_59,In_444);
or U273 (N_273,In_569,In_248);
nor U274 (N_274,In_501,In_19);
nor U275 (N_275,In_394,In_269);
or U276 (N_276,In_650,In_827);
nand U277 (N_277,In_794,In_414);
nor U278 (N_278,In_760,In_835);
xnor U279 (N_279,In_190,In_742);
xnor U280 (N_280,In_682,In_340);
nand U281 (N_281,In_769,In_701);
and U282 (N_282,In_696,In_706);
and U283 (N_283,In_834,In_468);
or U284 (N_284,In_263,In_330);
or U285 (N_285,In_616,In_793);
nor U286 (N_286,In_322,In_286);
and U287 (N_287,In_787,In_385);
and U288 (N_288,In_447,In_121);
and U289 (N_289,In_534,In_740);
or U290 (N_290,In_211,In_811);
xnor U291 (N_291,In_57,In_259);
nor U292 (N_292,In_170,In_76);
or U293 (N_293,In_182,In_517);
nand U294 (N_294,In_220,In_124);
nand U295 (N_295,In_488,In_505);
and U296 (N_296,In_301,In_62);
nand U297 (N_297,In_499,In_42);
xnor U298 (N_298,In_397,In_931);
and U299 (N_299,In_544,In_551);
or U300 (N_300,In_840,In_176);
nor U301 (N_301,In_316,In_295);
nand U302 (N_302,In_929,In_352);
nor U303 (N_303,In_401,In_767);
or U304 (N_304,In_106,In_172);
nor U305 (N_305,In_814,In_138);
or U306 (N_306,In_717,In_335);
xnor U307 (N_307,In_557,In_270);
and U308 (N_308,In_360,In_554);
nor U309 (N_309,In_429,In_521);
and U310 (N_310,In_622,In_898);
and U311 (N_311,In_901,In_626);
xor U312 (N_312,In_118,In_751);
and U313 (N_313,In_69,In_714);
nor U314 (N_314,In_386,In_287);
nand U315 (N_315,In_380,In_913);
or U316 (N_316,In_454,In_354);
or U317 (N_317,In_792,In_954);
nand U318 (N_318,In_748,In_617);
and U319 (N_319,In_91,In_207);
nor U320 (N_320,In_513,In_273);
nand U321 (N_321,In_388,In_601);
nor U322 (N_322,In_549,In_237);
nor U323 (N_323,In_623,In_809);
and U324 (N_324,In_416,In_589);
xor U325 (N_325,In_9,In_518);
and U326 (N_326,In_763,In_294);
and U327 (N_327,In_75,In_830);
and U328 (N_328,In_848,In_218);
nand U329 (N_329,In_770,In_649);
xor U330 (N_330,In_709,In_911);
and U331 (N_331,In_877,In_625);
nor U332 (N_332,In_103,In_702);
or U333 (N_333,In_438,In_84);
nor U334 (N_334,In_464,In_721);
nand U335 (N_335,In_201,In_297);
nand U336 (N_336,In_880,In_494);
nor U337 (N_337,In_392,In_639);
nor U338 (N_338,In_866,In_507);
and U339 (N_339,In_381,In_12);
nand U340 (N_340,In_226,In_678);
or U341 (N_341,In_480,In_944);
and U342 (N_342,In_465,In_697);
xor U343 (N_343,In_296,In_582);
nand U344 (N_344,In_894,In_719);
nor U345 (N_345,In_800,In_683);
and U346 (N_346,In_539,In_643);
and U347 (N_347,In_408,In_596);
nor U348 (N_348,In_859,In_752);
and U349 (N_349,In_941,In_936);
nor U350 (N_350,In_418,In_910);
nand U351 (N_351,In_729,In_110);
or U352 (N_352,In_186,In_753);
and U353 (N_353,In_257,In_780);
nor U354 (N_354,In_734,In_178);
or U355 (N_355,In_668,In_383);
and U356 (N_356,In_978,In_406);
nor U357 (N_357,In_885,In_156);
xnor U358 (N_358,In_577,In_255);
and U359 (N_359,In_212,In_231);
nand U360 (N_360,In_204,In_825);
or U361 (N_361,In_758,In_437);
or U362 (N_362,In_159,In_202);
nand U363 (N_363,In_570,In_759);
or U364 (N_364,In_512,In_595);
or U365 (N_365,In_485,In_232);
nor U366 (N_366,In_783,In_8);
xnor U367 (N_367,In_336,In_26);
nor U368 (N_368,In_768,In_593);
nor U369 (N_369,In_1,In_177);
nand U370 (N_370,In_689,In_82);
and U371 (N_371,In_890,In_448);
xnor U372 (N_372,In_461,In_332);
and U373 (N_373,In_284,In_711);
xnor U374 (N_374,In_145,In_693);
nor U375 (N_375,In_590,In_491);
xnor U376 (N_376,In_909,In_440);
nand U377 (N_377,In_637,In_586);
or U378 (N_378,In_326,In_628);
xnor U379 (N_379,In_303,In_149);
nand U380 (N_380,In_490,In_347);
nor U381 (N_381,In_864,In_722);
xor U382 (N_382,In_940,In_71);
and U383 (N_383,In_578,In_999);
xor U384 (N_384,In_695,In_927);
and U385 (N_385,In_391,In_113);
nor U386 (N_386,In_315,In_968);
nand U387 (N_387,In_100,In_173);
and U388 (N_388,In_387,In_374);
nor U389 (N_389,In_267,In_60);
or U390 (N_390,In_102,In_561);
or U391 (N_391,In_466,In_817);
xnor U392 (N_392,In_662,In_472);
or U393 (N_393,In_967,In_196);
or U394 (N_394,In_934,In_5);
or U395 (N_395,In_469,In_174);
nand U396 (N_396,In_803,In_236);
xnor U397 (N_397,In_30,In_81);
and U398 (N_398,In_948,In_495);
or U399 (N_399,In_262,In_185);
nand U400 (N_400,In_906,In_40);
nand U401 (N_401,In_379,In_559);
xnor U402 (N_402,In_547,In_141);
or U403 (N_403,In_304,In_67);
nand U404 (N_404,In_856,In_900);
nand U405 (N_405,In_624,In_519);
xor U406 (N_406,In_127,In_125);
nand U407 (N_407,In_200,In_74);
nor U408 (N_408,In_965,In_667);
and U409 (N_409,In_739,In_150);
nor U410 (N_410,In_271,In_756);
xnor U411 (N_411,In_452,In_871);
nor U412 (N_412,In_565,In_254);
and U413 (N_413,In_33,In_345);
nor U414 (N_414,In_167,In_798);
and U415 (N_415,In_333,In_246);
or U416 (N_416,In_109,In_713);
or U417 (N_417,In_893,In_681);
and U418 (N_418,In_476,In_378);
nor U419 (N_419,In_592,In_726);
xnor U420 (N_420,In_411,In_707);
nor U421 (N_421,In_486,In_525);
or U422 (N_422,In_970,In_422);
or U423 (N_423,In_664,In_537);
and U424 (N_424,In_887,In_715);
nand U425 (N_425,In_435,In_425);
xnor U426 (N_426,In_822,In_198);
nand U427 (N_427,In_179,In_661);
nor U428 (N_428,In_283,In_928);
nand U429 (N_429,In_430,In_655);
or U430 (N_430,In_556,In_504);
and U431 (N_431,In_886,In_107);
nor U432 (N_432,In_222,In_853);
and U433 (N_433,In_606,In_579);
nand U434 (N_434,In_874,In_982);
or U435 (N_435,In_197,In_366);
or U436 (N_436,In_741,In_241);
nor U437 (N_437,In_467,In_239);
and U438 (N_438,In_51,In_644);
nand U439 (N_439,In_443,In_642);
nor U440 (N_440,In_972,In_97);
and U441 (N_441,In_193,In_61);
and U442 (N_442,In_659,In_867);
nand U443 (N_443,In_836,In_638);
or U444 (N_444,In_873,In_872);
xnor U445 (N_445,In_243,In_812);
xnor U446 (N_446,In_41,In_94);
nor U447 (N_447,In_276,In_543);
nor U448 (N_448,In_782,In_314);
or U449 (N_449,In_610,In_245);
or U450 (N_450,In_175,In_806);
nand U451 (N_451,In_424,In_49);
or U452 (N_452,In_350,In_298);
and U453 (N_453,In_126,In_405);
and U454 (N_454,In_985,In_633);
nand U455 (N_455,In_365,In_869);
nor U456 (N_456,In_155,In_815);
nand U457 (N_457,In_17,In_44);
or U458 (N_458,In_46,In_88);
or U459 (N_459,In_677,In_823);
nand U460 (N_460,In_576,In_230);
nor U461 (N_461,In_264,In_334);
nand U462 (N_462,In_451,In_779);
nand U463 (N_463,In_905,In_265);
nand U464 (N_464,In_529,In_481);
or U465 (N_465,In_449,In_627);
xnor U466 (N_466,In_364,In_983);
and U467 (N_467,In_564,In_560);
or U468 (N_468,In_31,In_152);
and U469 (N_469,In_895,In_685);
nand U470 (N_470,In_285,In_441);
or U471 (N_471,In_789,In_399);
nand U472 (N_472,In_907,In_128);
nor U473 (N_473,In_166,In_567);
or U474 (N_474,In_802,In_87);
or U475 (N_475,In_445,In_712);
nand U476 (N_476,In_883,In_305);
nor U477 (N_477,In_421,In_821);
nor U478 (N_478,In_679,In_843);
xnor U479 (N_479,In_343,In_881);
nor U480 (N_480,In_497,In_772);
and U481 (N_481,In_844,In_858);
and U482 (N_482,In_279,In_778);
nand U483 (N_483,In_588,In_478);
nor U484 (N_484,In_180,In_11);
and U485 (N_485,In_694,In_219);
or U486 (N_486,In_77,In_656);
and U487 (N_487,In_652,In_290);
or U488 (N_488,In_854,In_522);
and U489 (N_489,In_932,In_22);
and U490 (N_490,In_16,In_541);
xor U491 (N_491,In_423,In_796);
nand U492 (N_492,In_660,In_191);
and U493 (N_493,In_818,In_870);
nor U494 (N_494,In_690,In_846);
and U495 (N_495,In_216,In_45);
xnor U496 (N_496,In_43,In_66);
nand U497 (N_497,In_921,In_977);
or U498 (N_498,In_375,In_417);
nand U499 (N_499,In_479,In_339);
or U500 (N_500,In_800,In_908);
nand U501 (N_501,In_789,In_147);
and U502 (N_502,In_44,In_752);
and U503 (N_503,In_709,In_986);
xor U504 (N_504,In_204,In_484);
and U505 (N_505,In_535,In_230);
nand U506 (N_506,In_794,In_501);
or U507 (N_507,In_530,In_156);
nand U508 (N_508,In_3,In_110);
nor U509 (N_509,In_157,In_479);
xnor U510 (N_510,In_110,In_672);
or U511 (N_511,In_123,In_140);
nor U512 (N_512,In_366,In_404);
nand U513 (N_513,In_523,In_609);
and U514 (N_514,In_123,In_825);
xor U515 (N_515,In_617,In_163);
and U516 (N_516,In_134,In_929);
nor U517 (N_517,In_536,In_356);
xnor U518 (N_518,In_414,In_145);
and U519 (N_519,In_482,In_379);
or U520 (N_520,In_159,In_528);
or U521 (N_521,In_123,In_689);
and U522 (N_522,In_393,In_199);
and U523 (N_523,In_56,In_801);
and U524 (N_524,In_267,In_87);
and U525 (N_525,In_396,In_953);
nand U526 (N_526,In_300,In_253);
or U527 (N_527,In_606,In_781);
or U528 (N_528,In_403,In_609);
nor U529 (N_529,In_40,In_797);
or U530 (N_530,In_956,In_656);
nand U531 (N_531,In_199,In_683);
and U532 (N_532,In_596,In_510);
nand U533 (N_533,In_619,In_990);
and U534 (N_534,In_328,In_393);
or U535 (N_535,In_336,In_743);
nand U536 (N_536,In_394,In_602);
or U537 (N_537,In_777,In_732);
nand U538 (N_538,In_179,In_451);
xor U539 (N_539,In_287,In_319);
and U540 (N_540,In_893,In_657);
nor U541 (N_541,In_888,In_233);
nor U542 (N_542,In_772,In_369);
nand U543 (N_543,In_374,In_252);
nor U544 (N_544,In_22,In_280);
xor U545 (N_545,In_778,In_510);
nor U546 (N_546,In_985,In_796);
nor U547 (N_547,In_641,In_719);
nor U548 (N_548,In_469,In_244);
or U549 (N_549,In_479,In_947);
nand U550 (N_550,In_664,In_352);
xnor U551 (N_551,In_316,In_413);
nor U552 (N_552,In_174,In_110);
nand U553 (N_553,In_901,In_107);
nor U554 (N_554,In_648,In_278);
nor U555 (N_555,In_48,In_362);
or U556 (N_556,In_900,In_24);
and U557 (N_557,In_142,In_258);
nand U558 (N_558,In_930,In_738);
nand U559 (N_559,In_670,In_702);
and U560 (N_560,In_452,In_653);
xor U561 (N_561,In_407,In_384);
nand U562 (N_562,In_447,In_340);
xor U563 (N_563,In_480,In_223);
nand U564 (N_564,In_541,In_608);
and U565 (N_565,In_946,In_357);
or U566 (N_566,In_14,In_169);
xnor U567 (N_567,In_522,In_757);
or U568 (N_568,In_786,In_946);
nand U569 (N_569,In_665,In_425);
or U570 (N_570,In_175,In_408);
and U571 (N_571,In_822,In_97);
nor U572 (N_572,In_493,In_242);
or U573 (N_573,In_97,In_71);
nor U574 (N_574,In_209,In_825);
or U575 (N_575,In_552,In_257);
and U576 (N_576,In_746,In_887);
nand U577 (N_577,In_305,In_376);
and U578 (N_578,In_394,In_174);
and U579 (N_579,In_87,In_507);
and U580 (N_580,In_900,In_1);
nor U581 (N_581,In_191,In_930);
and U582 (N_582,In_979,In_578);
nor U583 (N_583,In_446,In_231);
nor U584 (N_584,In_274,In_635);
and U585 (N_585,In_329,In_77);
nand U586 (N_586,In_535,In_990);
nor U587 (N_587,In_247,In_318);
and U588 (N_588,In_945,In_328);
nand U589 (N_589,In_242,In_451);
xnor U590 (N_590,In_831,In_84);
xnor U591 (N_591,In_993,In_121);
nor U592 (N_592,In_264,In_505);
nor U593 (N_593,In_486,In_890);
nor U594 (N_594,In_676,In_265);
and U595 (N_595,In_37,In_516);
xnor U596 (N_596,In_81,In_454);
nor U597 (N_597,In_318,In_825);
and U598 (N_598,In_163,In_648);
nand U599 (N_599,In_886,In_808);
and U600 (N_600,In_487,In_990);
or U601 (N_601,In_414,In_136);
nor U602 (N_602,In_148,In_511);
or U603 (N_603,In_487,In_773);
nor U604 (N_604,In_502,In_147);
and U605 (N_605,In_285,In_79);
and U606 (N_606,In_890,In_813);
nand U607 (N_607,In_608,In_295);
or U608 (N_608,In_114,In_648);
and U609 (N_609,In_924,In_976);
and U610 (N_610,In_177,In_475);
nand U611 (N_611,In_909,In_51);
or U612 (N_612,In_134,In_309);
or U613 (N_613,In_245,In_377);
nand U614 (N_614,In_64,In_739);
and U615 (N_615,In_539,In_996);
or U616 (N_616,In_25,In_311);
nor U617 (N_617,In_154,In_807);
nand U618 (N_618,In_207,In_203);
nor U619 (N_619,In_265,In_392);
xnor U620 (N_620,In_155,In_779);
nand U621 (N_621,In_799,In_280);
and U622 (N_622,In_18,In_936);
or U623 (N_623,In_132,In_205);
nand U624 (N_624,In_767,In_140);
xnor U625 (N_625,In_710,In_704);
xnor U626 (N_626,In_495,In_402);
nor U627 (N_627,In_931,In_929);
or U628 (N_628,In_809,In_609);
or U629 (N_629,In_616,In_922);
xor U630 (N_630,In_903,In_549);
nand U631 (N_631,In_897,In_825);
xnor U632 (N_632,In_702,In_112);
or U633 (N_633,In_787,In_138);
or U634 (N_634,In_872,In_269);
and U635 (N_635,In_332,In_875);
nand U636 (N_636,In_270,In_176);
or U637 (N_637,In_720,In_646);
or U638 (N_638,In_217,In_442);
nor U639 (N_639,In_42,In_305);
nand U640 (N_640,In_13,In_32);
nand U641 (N_641,In_611,In_290);
or U642 (N_642,In_874,In_978);
and U643 (N_643,In_954,In_164);
nand U644 (N_644,In_32,In_882);
nor U645 (N_645,In_663,In_656);
and U646 (N_646,In_121,In_428);
nand U647 (N_647,In_712,In_377);
nand U648 (N_648,In_187,In_276);
or U649 (N_649,In_959,In_837);
xor U650 (N_650,In_117,In_86);
nor U651 (N_651,In_758,In_44);
and U652 (N_652,In_886,In_546);
nand U653 (N_653,In_751,In_640);
xnor U654 (N_654,In_499,In_413);
and U655 (N_655,In_117,In_600);
and U656 (N_656,In_722,In_875);
or U657 (N_657,In_13,In_585);
and U658 (N_658,In_252,In_471);
or U659 (N_659,In_322,In_952);
or U660 (N_660,In_25,In_696);
nor U661 (N_661,In_683,In_500);
or U662 (N_662,In_542,In_443);
nor U663 (N_663,In_824,In_822);
nor U664 (N_664,In_830,In_380);
nand U665 (N_665,In_467,In_930);
nand U666 (N_666,In_216,In_275);
xor U667 (N_667,In_537,In_201);
nand U668 (N_668,In_757,In_8);
and U669 (N_669,In_291,In_701);
xnor U670 (N_670,In_524,In_293);
and U671 (N_671,In_141,In_154);
xnor U672 (N_672,In_486,In_261);
nor U673 (N_673,In_511,In_909);
nor U674 (N_674,In_644,In_630);
nor U675 (N_675,In_307,In_452);
nand U676 (N_676,In_954,In_296);
nor U677 (N_677,In_102,In_341);
and U678 (N_678,In_551,In_935);
nor U679 (N_679,In_620,In_873);
and U680 (N_680,In_87,In_538);
or U681 (N_681,In_239,In_674);
or U682 (N_682,In_715,In_245);
xor U683 (N_683,In_888,In_322);
or U684 (N_684,In_804,In_707);
or U685 (N_685,In_526,In_722);
xnor U686 (N_686,In_949,In_927);
nand U687 (N_687,In_196,In_707);
and U688 (N_688,In_511,In_535);
nor U689 (N_689,In_536,In_97);
nand U690 (N_690,In_332,In_505);
or U691 (N_691,In_666,In_75);
nor U692 (N_692,In_20,In_187);
xor U693 (N_693,In_495,In_685);
and U694 (N_694,In_844,In_969);
and U695 (N_695,In_154,In_395);
nand U696 (N_696,In_706,In_648);
and U697 (N_697,In_643,In_746);
and U698 (N_698,In_950,In_910);
or U699 (N_699,In_282,In_293);
or U700 (N_700,In_890,In_438);
or U701 (N_701,In_681,In_776);
nand U702 (N_702,In_193,In_342);
or U703 (N_703,In_309,In_483);
or U704 (N_704,In_751,In_152);
nand U705 (N_705,In_84,In_750);
or U706 (N_706,In_80,In_893);
nand U707 (N_707,In_586,In_619);
and U708 (N_708,In_591,In_123);
or U709 (N_709,In_355,In_841);
nand U710 (N_710,In_601,In_572);
xor U711 (N_711,In_359,In_497);
and U712 (N_712,In_529,In_10);
nand U713 (N_713,In_233,In_172);
nor U714 (N_714,In_517,In_804);
and U715 (N_715,In_841,In_749);
and U716 (N_716,In_325,In_640);
and U717 (N_717,In_864,In_479);
and U718 (N_718,In_551,In_463);
nor U719 (N_719,In_235,In_498);
or U720 (N_720,In_403,In_411);
and U721 (N_721,In_895,In_911);
nand U722 (N_722,In_995,In_711);
or U723 (N_723,In_393,In_695);
nor U724 (N_724,In_231,In_174);
xnor U725 (N_725,In_44,In_326);
or U726 (N_726,In_804,In_120);
nand U727 (N_727,In_482,In_200);
and U728 (N_728,In_826,In_684);
nor U729 (N_729,In_993,In_219);
nor U730 (N_730,In_74,In_674);
and U731 (N_731,In_608,In_201);
nand U732 (N_732,In_413,In_353);
and U733 (N_733,In_334,In_157);
or U734 (N_734,In_752,In_750);
nor U735 (N_735,In_459,In_413);
and U736 (N_736,In_732,In_942);
nand U737 (N_737,In_546,In_448);
xor U738 (N_738,In_54,In_260);
or U739 (N_739,In_137,In_72);
or U740 (N_740,In_788,In_934);
or U741 (N_741,In_25,In_669);
or U742 (N_742,In_240,In_980);
nand U743 (N_743,In_23,In_409);
or U744 (N_744,In_12,In_715);
nand U745 (N_745,In_56,In_750);
nor U746 (N_746,In_573,In_172);
nor U747 (N_747,In_391,In_726);
nor U748 (N_748,In_278,In_502);
or U749 (N_749,In_694,In_432);
xor U750 (N_750,In_620,In_44);
nor U751 (N_751,In_857,In_348);
nor U752 (N_752,In_740,In_661);
or U753 (N_753,In_121,In_35);
and U754 (N_754,In_126,In_901);
or U755 (N_755,In_255,In_484);
nand U756 (N_756,In_28,In_240);
xnor U757 (N_757,In_977,In_326);
and U758 (N_758,In_121,In_996);
xnor U759 (N_759,In_351,In_197);
or U760 (N_760,In_846,In_224);
or U761 (N_761,In_292,In_550);
or U762 (N_762,In_282,In_635);
xor U763 (N_763,In_490,In_504);
xor U764 (N_764,In_21,In_544);
nand U765 (N_765,In_754,In_176);
xnor U766 (N_766,In_983,In_964);
or U767 (N_767,In_302,In_818);
xnor U768 (N_768,In_269,In_613);
nand U769 (N_769,In_357,In_781);
nand U770 (N_770,In_168,In_336);
or U771 (N_771,In_922,In_770);
nand U772 (N_772,In_951,In_651);
xnor U773 (N_773,In_43,In_257);
xor U774 (N_774,In_865,In_367);
nor U775 (N_775,In_700,In_996);
nand U776 (N_776,In_946,In_76);
and U777 (N_777,In_614,In_21);
and U778 (N_778,In_834,In_707);
and U779 (N_779,In_384,In_67);
nor U780 (N_780,In_139,In_919);
nand U781 (N_781,In_207,In_676);
and U782 (N_782,In_541,In_946);
xor U783 (N_783,In_413,In_771);
or U784 (N_784,In_836,In_358);
and U785 (N_785,In_675,In_880);
nand U786 (N_786,In_239,In_687);
or U787 (N_787,In_794,In_901);
and U788 (N_788,In_1,In_659);
nor U789 (N_789,In_189,In_78);
or U790 (N_790,In_827,In_298);
or U791 (N_791,In_311,In_569);
nor U792 (N_792,In_502,In_399);
and U793 (N_793,In_475,In_325);
or U794 (N_794,In_536,In_103);
nor U795 (N_795,In_875,In_292);
xor U796 (N_796,In_855,In_604);
nor U797 (N_797,In_478,In_978);
nor U798 (N_798,In_997,In_52);
and U799 (N_799,In_352,In_666);
and U800 (N_800,In_270,In_318);
and U801 (N_801,In_179,In_751);
nor U802 (N_802,In_417,In_391);
or U803 (N_803,In_324,In_17);
nor U804 (N_804,In_851,In_835);
nor U805 (N_805,In_531,In_980);
or U806 (N_806,In_499,In_545);
and U807 (N_807,In_323,In_917);
nor U808 (N_808,In_729,In_592);
nor U809 (N_809,In_519,In_350);
and U810 (N_810,In_961,In_548);
and U811 (N_811,In_575,In_666);
nor U812 (N_812,In_930,In_226);
and U813 (N_813,In_269,In_19);
xor U814 (N_814,In_430,In_412);
nor U815 (N_815,In_747,In_514);
or U816 (N_816,In_104,In_933);
or U817 (N_817,In_342,In_372);
nand U818 (N_818,In_888,In_287);
and U819 (N_819,In_575,In_848);
nand U820 (N_820,In_702,In_57);
nor U821 (N_821,In_52,In_334);
or U822 (N_822,In_180,In_537);
nor U823 (N_823,In_648,In_431);
xor U824 (N_824,In_697,In_740);
nand U825 (N_825,In_625,In_779);
or U826 (N_826,In_479,In_510);
or U827 (N_827,In_151,In_363);
nor U828 (N_828,In_556,In_764);
or U829 (N_829,In_60,In_153);
nor U830 (N_830,In_661,In_518);
or U831 (N_831,In_423,In_727);
nand U832 (N_832,In_131,In_590);
or U833 (N_833,In_640,In_800);
xor U834 (N_834,In_826,In_629);
nand U835 (N_835,In_251,In_25);
nor U836 (N_836,In_94,In_381);
nand U837 (N_837,In_181,In_394);
or U838 (N_838,In_16,In_923);
xor U839 (N_839,In_270,In_822);
or U840 (N_840,In_851,In_755);
or U841 (N_841,In_308,In_405);
or U842 (N_842,In_46,In_909);
or U843 (N_843,In_184,In_469);
nor U844 (N_844,In_340,In_432);
nand U845 (N_845,In_788,In_110);
nand U846 (N_846,In_736,In_812);
nor U847 (N_847,In_547,In_758);
nor U848 (N_848,In_835,In_267);
xnor U849 (N_849,In_827,In_692);
nand U850 (N_850,In_476,In_428);
and U851 (N_851,In_7,In_390);
and U852 (N_852,In_789,In_234);
nor U853 (N_853,In_536,In_580);
and U854 (N_854,In_702,In_987);
nor U855 (N_855,In_217,In_894);
or U856 (N_856,In_434,In_76);
or U857 (N_857,In_288,In_483);
and U858 (N_858,In_636,In_587);
or U859 (N_859,In_813,In_667);
or U860 (N_860,In_615,In_883);
nand U861 (N_861,In_990,In_851);
xor U862 (N_862,In_643,In_993);
nand U863 (N_863,In_92,In_206);
xor U864 (N_864,In_474,In_907);
nor U865 (N_865,In_818,In_656);
xnor U866 (N_866,In_66,In_552);
nand U867 (N_867,In_246,In_214);
and U868 (N_868,In_274,In_668);
xor U869 (N_869,In_569,In_553);
nand U870 (N_870,In_135,In_347);
or U871 (N_871,In_790,In_299);
nand U872 (N_872,In_223,In_553);
and U873 (N_873,In_797,In_240);
and U874 (N_874,In_600,In_950);
nand U875 (N_875,In_96,In_787);
nor U876 (N_876,In_341,In_711);
nand U877 (N_877,In_467,In_683);
nand U878 (N_878,In_186,In_537);
or U879 (N_879,In_667,In_513);
nand U880 (N_880,In_891,In_339);
xnor U881 (N_881,In_91,In_57);
or U882 (N_882,In_351,In_599);
and U883 (N_883,In_178,In_595);
or U884 (N_884,In_506,In_110);
nor U885 (N_885,In_892,In_20);
nand U886 (N_886,In_342,In_506);
nand U887 (N_887,In_647,In_451);
and U888 (N_888,In_722,In_1);
nor U889 (N_889,In_926,In_15);
or U890 (N_890,In_259,In_175);
and U891 (N_891,In_421,In_108);
nand U892 (N_892,In_731,In_831);
nor U893 (N_893,In_156,In_37);
nor U894 (N_894,In_729,In_654);
xor U895 (N_895,In_706,In_484);
or U896 (N_896,In_687,In_310);
nor U897 (N_897,In_493,In_290);
or U898 (N_898,In_784,In_400);
nor U899 (N_899,In_633,In_33);
or U900 (N_900,In_917,In_800);
nand U901 (N_901,In_187,In_682);
or U902 (N_902,In_504,In_354);
nand U903 (N_903,In_351,In_117);
or U904 (N_904,In_536,In_300);
nor U905 (N_905,In_29,In_583);
xnor U906 (N_906,In_854,In_19);
nor U907 (N_907,In_380,In_704);
and U908 (N_908,In_170,In_387);
nand U909 (N_909,In_776,In_653);
and U910 (N_910,In_809,In_484);
or U911 (N_911,In_724,In_389);
or U912 (N_912,In_162,In_498);
nand U913 (N_913,In_150,In_832);
nor U914 (N_914,In_106,In_396);
and U915 (N_915,In_258,In_418);
and U916 (N_916,In_39,In_307);
and U917 (N_917,In_706,In_192);
nor U918 (N_918,In_210,In_300);
and U919 (N_919,In_837,In_165);
nor U920 (N_920,In_54,In_166);
nor U921 (N_921,In_441,In_9);
nor U922 (N_922,In_199,In_954);
and U923 (N_923,In_21,In_185);
nor U924 (N_924,In_734,In_620);
and U925 (N_925,In_102,In_970);
or U926 (N_926,In_115,In_729);
or U927 (N_927,In_525,In_265);
nand U928 (N_928,In_178,In_742);
or U929 (N_929,In_994,In_606);
or U930 (N_930,In_48,In_949);
or U931 (N_931,In_829,In_589);
or U932 (N_932,In_878,In_710);
or U933 (N_933,In_500,In_19);
nand U934 (N_934,In_586,In_739);
or U935 (N_935,In_906,In_300);
or U936 (N_936,In_106,In_537);
nand U937 (N_937,In_494,In_392);
nor U938 (N_938,In_801,In_787);
nand U939 (N_939,In_591,In_8);
and U940 (N_940,In_453,In_404);
and U941 (N_941,In_554,In_621);
nand U942 (N_942,In_646,In_179);
nand U943 (N_943,In_722,In_391);
or U944 (N_944,In_771,In_615);
xnor U945 (N_945,In_27,In_919);
nor U946 (N_946,In_373,In_306);
or U947 (N_947,In_615,In_720);
xnor U948 (N_948,In_840,In_502);
or U949 (N_949,In_888,In_635);
and U950 (N_950,In_204,In_499);
nand U951 (N_951,In_642,In_983);
or U952 (N_952,In_864,In_987);
xnor U953 (N_953,In_516,In_795);
nand U954 (N_954,In_108,In_386);
nand U955 (N_955,In_490,In_532);
nor U956 (N_956,In_98,In_378);
or U957 (N_957,In_661,In_330);
xnor U958 (N_958,In_523,In_998);
nand U959 (N_959,In_571,In_318);
nor U960 (N_960,In_642,In_979);
nor U961 (N_961,In_981,In_128);
and U962 (N_962,In_898,In_306);
nand U963 (N_963,In_323,In_174);
and U964 (N_964,In_817,In_789);
and U965 (N_965,In_47,In_332);
nor U966 (N_966,In_653,In_216);
or U967 (N_967,In_185,In_106);
nand U968 (N_968,In_534,In_498);
or U969 (N_969,In_588,In_271);
nor U970 (N_970,In_656,In_826);
and U971 (N_971,In_964,In_143);
nor U972 (N_972,In_480,In_256);
or U973 (N_973,In_453,In_371);
nor U974 (N_974,In_601,In_779);
and U975 (N_975,In_428,In_715);
or U976 (N_976,In_373,In_564);
nor U977 (N_977,In_975,In_63);
and U978 (N_978,In_646,In_477);
and U979 (N_979,In_150,In_867);
and U980 (N_980,In_158,In_348);
nor U981 (N_981,In_116,In_545);
nor U982 (N_982,In_299,In_659);
and U983 (N_983,In_933,In_417);
xor U984 (N_984,In_624,In_648);
nor U985 (N_985,In_145,In_133);
nand U986 (N_986,In_972,In_808);
nand U987 (N_987,In_920,In_703);
nor U988 (N_988,In_83,In_122);
or U989 (N_989,In_816,In_109);
and U990 (N_990,In_223,In_794);
or U991 (N_991,In_862,In_48);
nor U992 (N_992,In_405,In_888);
nor U993 (N_993,In_356,In_318);
xnor U994 (N_994,In_501,In_397);
or U995 (N_995,In_875,In_478);
nor U996 (N_996,In_983,In_740);
and U997 (N_997,In_176,In_11);
nand U998 (N_998,In_916,In_520);
nand U999 (N_999,In_731,In_4);
nand U1000 (N_1000,In_96,In_904);
and U1001 (N_1001,In_782,In_538);
xnor U1002 (N_1002,In_122,In_107);
xor U1003 (N_1003,In_421,In_71);
nor U1004 (N_1004,In_838,In_879);
or U1005 (N_1005,In_150,In_247);
nor U1006 (N_1006,In_250,In_904);
and U1007 (N_1007,In_404,In_55);
nor U1008 (N_1008,In_747,In_236);
nor U1009 (N_1009,In_628,In_286);
or U1010 (N_1010,In_995,In_998);
xor U1011 (N_1011,In_247,In_557);
nor U1012 (N_1012,In_585,In_386);
nand U1013 (N_1013,In_573,In_367);
nor U1014 (N_1014,In_800,In_355);
or U1015 (N_1015,In_978,In_905);
nand U1016 (N_1016,In_117,In_731);
nand U1017 (N_1017,In_486,In_103);
and U1018 (N_1018,In_196,In_443);
and U1019 (N_1019,In_188,In_603);
and U1020 (N_1020,In_57,In_625);
xor U1021 (N_1021,In_931,In_196);
and U1022 (N_1022,In_814,In_755);
and U1023 (N_1023,In_152,In_330);
xor U1024 (N_1024,In_761,In_747);
and U1025 (N_1025,In_426,In_17);
nand U1026 (N_1026,In_904,In_232);
and U1027 (N_1027,In_292,In_996);
and U1028 (N_1028,In_337,In_481);
nand U1029 (N_1029,In_39,In_370);
nor U1030 (N_1030,In_898,In_539);
or U1031 (N_1031,In_354,In_569);
nor U1032 (N_1032,In_454,In_577);
and U1033 (N_1033,In_192,In_624);
nand U1034 (N_1034,In_555,In_776);
nor U1035 (N_1035,In_720,In_118);
or U1036 (N_1036,In_282,In_946);
xnor U1037 (N_1037,In_495,In_204);
or U1038 (N_1038,In_43,In_323);
and U1039 (N_1039,In_221,In_964);
nand U1040 (N_1040,In_982,In_956);
and U1041 (N_1041,In_117,In_154);
nor U1042 (N_1042,In_593,In_915);
nand U1043 (N_1043,In_341,In_715);
xnor U1044 (N_1044,In_475,In_777);
nor U1045 (N_1045,In_862,In_359);
or U1046 (N_1046,In_737,In_855);
xor U1047 (N_1047,In_180,In_597);
or U1048 (N_1048,In_912,In_550);
nor U1049 (N_1049,In_973,In_731);
nand U1050 (N_1050,In_765,In_917);
nand U1051 (N_1051,In_75,In_241);
xnor U1052 (N_1052,In_455,In_812);
or U1053 (N_1053,In_859,In_176);
nor U1054 (N_1054,In_376,In_896);
or U1055 (N_1055,In_9,In_820);
nand U1056 (N_1056,In_668,In_523);
nor U1057 (N_1057,In_756,In_392);
nand U1058 (N_1058,In_361,In_525);
nand U1059 (N_1059,In_832,In_881);
and U1060 (N_1060,In_411,In_228);
nor U1061 (N_1061,In_165,In_659);
and U1062 (N_1062,In_181,In_747);
nand U1063 (N_1063,In_912,In_748);
nand U1064 (N_1064,In_305,In_74);
and U1065 (N_1065,In_143,In_74);
nor U1066 (N_1066,In_732,In_46);
nand U1067 (N_1067,In_953,In_987);
and U1068 (N_1068,In_982,In_186);
xnor U1069 (N_1069,In_173,In_855);
xor U1070 (N_1070,In_301,In_586);
and U1071 (N_1071,In_0,In_241);
nor U1072 (N_1072,In_692,In_212);
nand U1073 (N_1073,In_273,In_343);
or U1074 (N_1074,In_737,In_958);
nor U1075 (N_1075,In_249,In_778);
or U1076 (N_1076,In_196,In_458);
nor U1077 (N_1077,In_354,In_804);
nand U1078 (N_1078,In_667,In_420);
nor U1079 (N_1079,In_451,In_253);
nand U1080 (N_1080,In_76,In_462);
nor U1081 (N_1081,In_667,In_562);
nor U1082 (N_1082,In_975,In_662);
nor U1083 (N_1083,In_32,In_955);
and U1084 (N_1084,In_827,In_792);
nand U1085 (N_1085,In_725,In_918);
nand U1086 (N_1086,In_395,In_690);
nor U1087 (N_1087,In_91,In_157);
nand U1088 (N_1088,In_917,In_901);
and U1089 (N_1089,In_264,In_634);
or U1090 (N_1090,In_181,In_777);
nand U1091 (N_1091,In_943,In_495);
and U1092 (N_1092,In_756,In_813);
and U1093 (N_1093,In_857,In_939);
or U1094 (N_1094,In_972,In_774);
or U1095 (N_1095,In_672,In_893);
xnor U1096 (N_1096,In_148,In_155);
and U1097 (N_1097,In_775,In_130);
nor U1098 (N_1098,In_602,In_165);
or U1099 (N_1099,In_367,In_989);
and U1100 (N_1100,In_665,In_122);
and U1101 (N_1101,In_29,In_57);
nand U1102 (N_1102,In_600,In_345);
xor U1103 (N_1103,In_718,In_406);
or U1104 (N_1104,In_261,In_306);
or U1105 (N_1105,In_313,In_587);
or U1106 (N_1106,In_269,In_441);
or U1107 (N_1107,In_180,In_30);
nand U1108 (N_1108,In_656,In_680);
nand U1109 (N_1109,In_560,In_207);
nand U1110 (N_1110,In_41,In_269);
and U1111 (N_1111,In_780,In_857);
nor U1112 (N_1112,In_555,In_460);
or U1113 (N_1113,In_211,In_339);
or U1114 (N_1114,In_291,In_496);
nand U1115 (N_1115,In_261,In_173);
nor U1116 (N_1116,In_260,In_114);
or U1117 (N_1117,In_189,In_408);
and U1118 (N_1118,In_217,In_592);
nor U1119 (N_1119,In_362,In_448);
xnor U1120 (N_1120,In_519,In_3);
and U1121 (N_1121,In_82,In_521);
nand U1122 (N_1122,In_933,In_142);
and U1123 (N_1123,In_825,In_684);
and U1124 (N_1124,In_626,In_880);
nor U1125 (N_1125,In_22,In_410);
nor U1126 (N_1126,In_926,In_824);
nor U1127 (N_1127,In_460,In_579);
nand U1128 (N_1128,In_576,In_141);
xor U1129 (N_1129,In_390,In_304);
or U1130 (N_1130,In_101,In_946);
nor U1131 (N_1131,In_112,In_562);
and U1132 (N_1132,In_834,In_356);
nor U1133 (N_1133,In_303,In_178);
nor U1134 (N_1134,In_786,In_950);
nand U1135 (N_1135,In_211,In_678);
nand U1136 (N_1136,In_223,In_363);
nand U1137 (N_1137,In_217,In_954);
xnor U1138 (N_1138,In_872,In_942);
or U1139 (N_1139,In_794,In_342);
xnor U1140 (N_1140,In_107,In_428);
nand U1141 (N_1141,In_314,In_606);
or U1142 (N_1142,In_160,In_239);
or U1143 (N_1143,In_923,In_346);
or U1144 (N_1144,In_555,In_529);
nor U1145 (N_1145,In_881,In_196);
nor U1146 (N_1146,In_114,In_854);
nor U1147 (N_1147,In_679,In_822);
or U1148 (N_1148,In_97,In_725);
or U1149 (N_1149,In_559,In_649);
nand U1150 (N_1150,In_445,In_620);
and U1151 (N_1151,In_140,In_269);
nor U1152 (N_1152,In_224,In_498);
nor U1153 (N_1153,In_902,In_302);
xnor U1154 (N_1154,In_335,In_91);
nand U1155 (N_1155,In_470,In_294);
and U1156 (N_1156,In_368,In_740);
nor U1157 (N_1157,In_988,In_334);
nand U1158 (N_1158,In_555,In_881);
or U1159 (N_1159,In_580,In_970);
nand U1160 (N_1160,In_145,In_566);
or U1161 (N_1161,In_116,In_867);
or U1162 (N_1162,In_275,In_395);
nor U1163 (N_1163,In_852,In_844);
nand U1164 (N_1164,In_220,In_461);
nand U1165 (N_1165,In_167,In_522);
and U1166 (N_1166,In_560,In_804);
or U1167 (N_1167,In_993,In_102);
nand U1168 (N_1168,In_692,In_614);
and U1169 (N_1169,In_350,In_208);
or U1170 (N_1170,In_236,In_162);
nor U1171 (N_1171,In_786,In_902);
or U1172 (N_1172,In_643,In_111);
nor U1173 (N_1173,In_774,In_345);
nor U1174 (N_1174,In_502,In_635);
nor U1175 (N_1175,In_13,In_342);
xor U1176 (N_1176,In_555,In_372);
and U1177 (N_1177,In_107,In_210);
nand U1178 (N_1178,In_187,In_862);
and U1179 (N_1179,In_834,In_730);
nor U1180 (N_1180,In_850,In_401);
nor U1181 (N_1181,In_785,In_169);
and U1182 (N_1182,In_6,In_81);
xor U1183 (N_1183,In_931,In_866);
nor U1184 (N_1184,In_274,In_922);
and U1185 (N_1185,In_486,In_54);
and U1186 (N_1186,In_429,In_275);
nand U1187 (N_1187,In_137,In_124);
nand U1188 (N_1188,In_992,In_457);
or U1189 (N_1189,In_322,In_292);
or U1190 (N_1190,In_947,In_600);
nor U1191 (N_1191,In_462,In_211);
nor U1192 (N_1192,In_343,In_729);
nor U1193 (N_1193,In_18,In_832);
nand U1194 (N_1194,In_10,In_923);
or U1195 (N_1195,In_535,In_836);
nand U1196 (N_1196,In_83,In_378);
nor U1197 (N_1197,In_313,In_566);
or U1198 (N_1198,In_311,In_142);
nor U1199 (N_1199,In_901,In_39);
nand U1200 (N_1200,In_753,In_5);
and U1201 (N_1201,In_731,In_668);
nor U1202 (N_1202,In_811,In_624);
nor U1203 (N_1203,In_993,In_206);
and U1204 (N_1204,In_694,In_372);
nor U1205 (N_1205,In_592,In_757);
nand U1206 (N_1206,In_261,In_132);
or U1207 (N_1207,In_651,In_508);
or U1208 (N_1208,In_476,In_441);
nor U1209 (N_1209,In_193,In_512);
and U1210 (N_1210,In_789,In_926);
or U1211 (N_1211,In_966,In_999);
or U1212 (N_1212,In_881,In_603);
and U1213 (N_1213,In_829,In_296);
and U1214 (N_1214,In_328,In_827);
or U1215 (N_1215,In_991,In_0);
and U1216 (N_1216,In_35,In_775);
and U1217 (N_1217,In_398,In_212);
and U1218 (N_1218,In_857,In_155);
and U1219 (N_1219,In_794,In_255);
nand U1220 (N_1220,In_8,In_57);
and U1221 (N_1221,In_766,In_755);
nand U1222 (N_1222,In_737,In_319);
nor U1223 (N_1223,In_330,In_6);
nor U1224 (N_1224,In_109,In_395);
nor U1225 (N_1225,In_806,In_274);
and U1226 (N_1226,In_822,In_247);
and U1227 (N_1227,In_845,In_263);
nor U1228 (N_1228,In_320,In_307);
nor U1229 (N_1229,In_92,In_86);
nand U1230 (N_1230,In_589,In_345);
nor U1231 (N_1231,In_481,In_599);
or U1232 (N_1232,In_960,In_93);
nand U1233 (N_1233,In_135,In_895);
xnor U1234 (N_1234,In_454,In_445);
or U1235 (N_1235,In_773,In_270);
nand U1236 (N_1236,In_358,In_500);
nor U1237 (N_1237,In_225,In_469);
nand U1238 (N_1238,In_514,In_904);
and U1239 (N_1239,In_36,In_839);
or U1240 (N_1240,In_941,In_710);
nand U1241 (N_1241,In_160,In_738);
nand U1242 (N_1242,In_604,In_764);
and U1243 (N_1243,In_252,In_933);
nor U1244 (N_1244,In_495,In_297);
nand U1245 (N_1245,In_947,In_394);
and U1246 (N_1246,In_331,In_380);
nand U1247 (N_1247,In_446,In_648);
or U1248 (N_1248,In_440,In_946);
and U1249 (N_1249,In_705,In_716);
and U1250 (N_1250,In_575,In_158);
and U1251 (N_1251,In_182,In_460);
and U1252 (N_1252,In_640,In_822);
and U1253 (N_1253,In_467,In_766);
and U1254 (N_1254,In_910,In_987);
and U1255 (N_1255,In_705,In_178);
nor U1256 (N_1256,In_460,In_230);
nand U1257 (N_1257,In_212,In_202);
xor U1258 (N_1258,In_521,In_479);
and U1259 (N_1259,In_814,In_383);
and U1260 (N_1260,In_988,In_442);
and U1261 (N_1261,In_812,In_203);
and U1262 (N_1262,In_536,In_129);
nand U1263 (N_1263,In_501,In_594);
nor U1264 (N_1264,In_219,In_503);
and U1265 (N_1265,In_149,In_490);
or U1266 (N_1266,In_805,In_886);
nand U1267 (N_1267,In_502,In_101);
and U1268 (N_1268,In_780,In_747);
nor U1269 (N_1269,In_265,In_824);
nand U1270 (N_1270,In_969,In_790);
and U1271 (N_1271,In_160,In_139);
nand U1272 (N_1272,In_823,In_630);
nor U1273 (N_1273,In_742,In_433);
or U1274 (N_1274,In_332,In_545);
or U1275 (N_1275,In_718,In_545);
nor U1276 (N_1276,In_344,In_84);
nand U1277 (N_1277,In_128,In_307);
and U1278 (N_1278,In_661,In_70);
nor U1279 (N_1279,In_861,In_966);
nor U1280 (N_1280,In_338,In_520);
nor U1281 (N_1281,In_906,In_665);
and U1282 (N_1282,In_459,In_174);
nand U1283 (N_1283,In_24,In_207);
nor U1284 (N_1284,In_950,In_981);
nor U1285 (N_1285,In_47,In_874);
nor U1286 (N_1286,In_627,In_597);
nor U1287 (N_1287,In_654,In_604);
or U1288 (N_1288,In_212,In_681);
and U1289 (N_1289,In_846,In_284);
nand U1290 (N_1290,In_254,In_385);
and U1291 (N_1291,In_226,In_325);
and U1292 (N_1292,In_349,In_138);
nand U1293 (N_1293,In_214,In_488);
or U1294 (N_1294,In_835,In_382);
nand U1295 (N_1295,In_638,In_683);
or U1296 (N_1296,In_113,In_667);
xnor U1297 (N_1297,In_877,In_917);
nor U1298 (N_1298,In_874,In_203);
or U1299 (N_1299,In_619,In_484);
nor U1300 (N_1300,In_345,In_99);
and U1301 (N_1301,In_631,In_549);
nor U1302 (N_1302,In_491,In_111);
and U1303 (N_1303,In_598,In_981);
nor U1304 (N_1304,In_199,In_964);
and U1305 (N_1305,In_924,In_180);
or U1306 (N_1306,In_534,In_909);
xnor U1307 (N_1307,In_386,In_96);
or U1308 (N_1308,In_71,In_346);
and U1309 (N_1309,In_441,In_578);
and U1310 (N_1310,In_232,In_684);
and U1311 (N_1311,In_301,In_662);
or U1312 (N_1312,In_279,In_110);
nand U1313 (N_1313,In_0,In_481);
or U1314 (N_1314,In_506,In_691);
or U1315 (N_1315,In_997,In_802);
and U1316 (N_1316,In_391,In_937);
nor U1317 (N_1317,In_41,In_449);
and U1318 (N_1318,In_962,In_260);
nor U1319 (N_1319,In_12,In_235);
nor U1320 (N_1320,In_330,In_236);
nor U1321 (N_1321,In_351,In_62);
nand U1322 (N_1322,In_659,In_580);
or U1323 (N_1323,In_882,In_163);
and U1324 (N_1324,In_82,In_42);
and U1325 (N_1325,In_167,In_615);
nand U1326 (N_1326,In_827,In_735);
nand U1327 (N_1327,In_296,In_78);
and U1328 (N_1328,In_355,In_73);
nand U1329 (N_1329,In_687,In_638);
nand U1330 (N_1330,In_140,In_599);
nand U1331 (N_1331,In_507,In_576);
or U1332 (N_1332,In_487,In_459);
nand U1333 (N_1333,In_751,In_57);
and U1334 (N_1334,In_374,In_467);
nor U1335 (N_1335,In_946,In_738);
and U1336 (N_1336,In_461,In_68);
and U1337 (N_1337,In_752,In_457);
or U1338 (N_1338,In_125,In_27);
nor U1339 (N_1339,In_88,In_651);
and U1340 (N_1340,In_736,In_329);
nor U1341 (N_1341,In_101,In_743);
or U1342 (N_1342,In_796,In_200);
and U1343 (N_1343,In_186,In_298);
and U1344 (N_1344,In_127,In_320);
and U1345 (N_1345,In_986,In_561);
nor U1346 (N_1346,In_454,In_487);
nand U1347 (N_1347,In_947,In_372);
or U1348 (N_1348,In_899,In_828);
and U1349 (N_1349,In_596,In_688);
nand U1350 (N_1350,In_380,In_930);
nand U1351 (N_1351,In_498,In_424);
xor U1352 (N_1352,In_523,In_237);
nor U1353 (N_1353,In_897,In_583);
or U1354 (N_1354,In_224,In_606);
nand U1355 (N_1355,In_272,In_512);
or U1356 (N_1356,In_656,In_590);
nor U1357 (N_1357,In_219,In_703);
and U1358 (N_1358,In_324,In_700);
or U1359 (N_1359,In_215,In_804);
nor U1360 (N_1360,In_511,In_902);
nand U1361 (N_1361,In_37,In_296);
nand U1362 (N_1362,In_215,In_632);
nand U1363 (N_1363,In_64,In_579);
nand U1364 (N_1364,In_522,In_998);
and U1365 (N_1365,In_570,In_752);
and U1366 (N_1366,In_239,In_945);
and U1367 (N_1367,In_56,In_392);
and U1368 (N_1368,In_985,In_70);
nor U1369 (N_1369,In_163,In_153);
or U1370 (N_1370,In_973,In_229);
and U1371 (N_1371,In_824,In_107);
nor U1372 (N_1372,In_107,In_587);
nor U1373 (N_1373,In_814,In_875);
or U1374 (N_1374,In_108,In_367);
nand U1375 (N_1375,In_921,In_392);
nand U1376 (N_1376,In_151,In_175);
or U1377 (N_1377,In_597,In_350);
and U1378 (N_1378,In_904,In_883);
or U1379 (N_1379,In_453,In_689);
xnor U1380 (N_1380,In_211,In_561);
nor U1381 (N_1381,In_511,In_204);
nand U1382 (N_1382,In_295,In_36);
or U1383 (N_1383,In_154,In_840);
nand U1384 (N_1384,In_585,In_446);
or U1385 (N_1385,In_478,In_919);
or U1386 (N_1386,In_912,In_233);
nor U1387 (N_1387,In_176,In_605);
nand U1388 (N_1388,In_606,In_791);
and U1389 (N_1389,In_164,In_614);
xor U1390 (N_1390,In_163,In_963);
nor U1391 (N_1391,In_154,In_342);
nor U1392 (N_1392,In_234,In_65);
or U1393 (N_1393,In_115,In_842);
and U1394 (N_1394,In_574,In_726);
nand U1395 (N_1395,In_560,In_679);
nand U1396 (N_1396,In_285,In_740);
or U1397 (N_1397,In_386,In_652);
nor U1398 (N_1398,In_783,In_89);
nand U1399 (N_1399,In_959,In_887);
and U1400 (N_1400,In_866,In_969);
nor U1401 (N_1401,In_723,In_797);
and U1402 (N_1402,In_18,In_677);
nor U1403 (N_1403,In_295,In_890);
nor U1404 (N_1404,In_496,In_211);
nor U1405 (N_1405,In_80,In_649);
xor U1406 (N_1406,In_466,In_668);
nor U1407 (N_1407,In_623,In_324);
xor U1408 (N_1408,In_142,In_234);
xnor U1409 (N_1409,In_454,In_690);
nand U1410 (N_1410,In_512,In_14);
or U1411 (N_1411,In_993,In_252);
xnor U1412 (N_1412,In_834,In_338);
or U1413 (N_1413,In_276,In_425);
xnor U1414 (N_1414,In_756,In_317);
nand U1415 (N_1415,In_56,In_172);
xor U1416 (N_1416,In_345,In_781);
nor U1417 (N_1417,In_818,In_999);
nor U1418 (N_1418,In_583,In_489);
nand U1419 (N_1419,In_860,In_174);
and U1420 (N_1420,In_67,In_293);
and U1421 (N_1421,In_690,In_520);
and U1422 (N_1422,In_679,In_94);
or U1423 (N_1423,In_909,In_773);
and U1424 (N_1424,In_486,In_608);
nand U1425 (N_1425,In_314,In_962);
or U1426 (N_1426,In_28,In_196);
xnor U1427 (N_1427,In_755,In_305);
nand U1428 (N_1428,In_425,In_155);
nand U1429 (N_1429,In_41,In_916);
nand U1430 (N_1430,In_59,In_232);
nor U1431 (N_1431,In_989,In_627);
nand U1432 (N_1432,In_517,In_778);
and U1433 (N_1433,In_180,In_497);
or U1434 (N_1434,In_672,In_413);
xor U1435 (N_1435,In_6,In_20);
nand U1436 (N_1436,In_948,In_674);
nand U1437 (N_1437,In_513,In_753);
nand U1438 (N_1438,In_211,In_194);
nand U1439 (N_1439,In_436,In_978);
and U1440 (N_1440,In_383,In_185);
or U1441 (N_1441,In_136,In_212);
and U1442 (N_1442,In_428,In_875);
or U1443 (N_1443,In_862,In_880);
or U1444 (N_1444,In_150,In_541);
nand U1445 (N_1445,In_663,In_865);
nor U1446 (N_1446,In_320,In_323);
nor U1447 (N_1447,In_126,In_19);
nand U1448 (N_1448,In_909,In_891);
and U1449 (N_1449,In_996,In_239);
nor U1450 (N_1450,In_170,In_943);
nand U1451 (N_1451,In_885,In_932);
nand U1452 (N_1452,In_855,In_409);
nor U1453 (N_1453,In_441,In_865);
nor U1454 (N_1454,In_85,In_937);
or U1455 (N_1455,In_360,In_928);
nor U1456 (N_1456,In_946,In_270);
or U1457 (N_1457,In_171,In_860);
and U1458 (N_1458,In_118,In_817);
nor U1459 (N_1459,In_4,In_49);
xor U1460 (N_1460,In_910,In_503);
xnor U1461 (N_1461,In_696,In_937);
nand U1462 (N_1462,In_457,In_883);
nand U1463 (N_1463,In_547,In_746);
and U1464 (N_1464,In_429,In_757);
or U1465 (N_1465,In_564,In_754);
and U1466 (N_1466,In_111,In_761);
nand U1467 (N_1467,In_88,In_18);
nor U1468 (N_1468,In_746,In_108);
nand U1469 (N_1469,In_827,In_978);
xor U1470 (N_1470,In_906,In_623);
nand U1471 (N_1471,In_446,In_738);
and U1472 (N_1472,In_258,In_150);
or U1473 (N_1473,In_179,In_734);
and U1474 (N_1474,In_105,In_261);
or U1475 (N_1475,In_996,In_344);
nand U1476 (N_1476,In_739,In_339);
nor U1477 (N_1477,In_459,In_662);
nand U1478 (N_1478,In_156,In_68);
nor U1479 (N_1479,In_299,In_745);
nand U1480 (N_1480,In_516,In_446);
nor U1481 (N_1481,In_710,In_392);
and U1482 (N_1482,In_302,In_150);
and U1483 (N_1483,In_547,In_608);
nor U1484 (N_1484,In_400,In_274);
or U1485 (N_1485,In_545,In_515);
or U1486 (N_1486,In_836,In_668);
or U1487 (N_1487,In_866,In_944);
nand U1488 (N_1488,In_528,In_369);
nand U1489 (N_1489,In_35,In_500);
or U1490 (N_1490,In_237,In_556);
xor U1491 (N_1491,In_236,In_844);
and U1492 (N_1492,In_251,In_814);
xnor U1493 (N_1493,In_489,In_974);
nand U1494 (N_1494,In_270,In_418);
or U1495 (N_1495,In_64,In_362);
or U1496 (N_1496,In_40,In_337);
nand U1497 (N_1497,In_715,In_638);
nand U1498 (N_1498,In_335,In_128);
or U1499 (N_1499,In_353,In_40);
or U1500 (N_1500,In_235,In_20);
and U1501 (N_1501,In_136,In_404);
and U1502 (N_1502,In_269,In_354);
nor U1503 (N_1503,In_635,In_578);
or U1504 (N_1504,In_325,In_178);
or U1505 (N_1505,In_504,In_909);
nand U1506 (N_1506,In_917,In_861);
nand U1507 (N_1507,In_641,In_82);
nand U1508 (N_1508,In_831,In_361);
nand U1509 (N_1509,In_37,In_97);
nand U1510 (N_1510,In_579,In_396);
nor U1511 (N_1511,In_242,In_127);
nor U1512 (N_1512,In_474,In_290);
and U1513 (N_1513,In_515,In_80);
or U1514 (N_1514,In_476,In_529);
nand U1515 (N_1515,In_217,In_105);
or U1516 (N_1516,In_143,In_862);
nand U1517 (N_1517,In_613,In_272);
or U1518 (N_1518,In_383,In_811);
and U1519 (N_1519,In_974,In_40);
and U1520 (N_1520,In_94,In_372);
or U1521 (N_1521,In_968,In_409);
nand U1522 (N_1522,In_756,In_11);
nor U1523 (N_1523,In_863,In_21);
xnor U1524 (N_1524,In_658,In_937);
nand U1525 (N_1525,In_277,In_661);
nand U1526 (N_1526,In_963,In_918);
or U1527 (N_1527,In_887,In_491);
nand U1528 (N_1528,In_698,In_734);
nand U1529 (N_1529,In_495,In_780);
or U1530 (N_1530,In_361,In_823);
nand U1531 (N_1531,In_355,In_53);
nand U1532 (N_1532,In_112,In_962);
and U1533 (N_1533,In_820,In_772);
nor U1534 (N_1534,In_932,In_309);
nor U1535 (N_1535,In_876,In_13);
or U1536 (N_1536,In_129,In_982);
nand U1537 (N_1537,In_886,In_888);
xor U1538 (N_1538,In_786,In_71);
nor U1539 (N_1539,In_217,In_953);
and U1540 (N_1540,In_562,In_786);
or U1541 (N_1541,In_4,In_650);
and U1542 (N_1542,In_472,In_624);
nand U1543 (N_1543,In_570,In_161);
or U1544 (N_1544,In_472,In_320);
or U1545 (N_1545,In_950,In_696);
nand U1546 (N_1546,In_488,In_593);
nand U1547 (N_1547,In_226,In_636);
and U1548 (N_1548,In_558,In_408);
nand U1549 (N_1549,In_346,In_332);
or U1550 (N_1550,In_45,In_964);
or U1551 (N_1551,In_496,In_746);
nand U1552 (N_1552,In_146,In_341);
or U1553 (N_1553,In_898,In_124);
or U1554 (N_1554,In_631,In_293);
or U1555 (N_1555,In_298,In_187);
xnor U1556 (N_1556,In_837,In_387);
and U1557 (N_1557,In_509,In_221);
and U1558 (N_1558,In_48,In_502);
xor U1559 (N_1559,In_775,In_675);
nand U1560 (N_1560,In_398,In_489);
nand U1561 (N_1561,In_377,In_840);
nand U1562 (N_1562,In_56,In_516);
and U1563 (N_1563,In_91,In_447);
and U1564 (N_1564,In_549,In_26);
and U1565 (N_1565,In_984,In_809);
and U1566 (N_1566,In_653,In_732);
nor U1567 (N_1567,In_47,In_922);
xor U1568 (N_1568,In_696,In_677);
and U1569 (N_1569,In_150,In_804);
nor U1570 (N_1570,In_537,In_31);
nor U1571 (N_1571,In_375,In_697);
nor U1572 (N_1572,In_190,In_609);
nor U1573 (N_1573,In_349,In_822);
nand U1574 (N_1574,In_78,In_309);
or U1575 (N_1575,In_722,In_59);
nand U1576 (N_1576,In_274,In_571);
xnor U1577 (N_1577,In_528,In_242);
or U1578 (N_1578,In_457,In_0);
nand U1579 (N_1579,In_970,In_934);
or U1580 (N_1580,In_261,In_836);
or U1581 (N_1581,In_713,In_402);
and U1582 (N_1582,In_615,In_211);
nand U1583 (N_1583,In_257,In_907);
or U1584 (N_1584,In_990,In_783);
nand U1585 (N_1585,In_702,In_747);
or U1586 (N_1586,In_761,In_976);
xnor U1587 (N_1587,In_99,In_249);
nand U1588 (N_1588,In_11,In_660);
nand U1589 (N_1589,In_889,In_395);
and U1590 (N_1590,In_86,In_10);
nor U1591 (N_1591,In_225,In_639);
and U1592 (N_1592,In_840,In_903);
nand U1593 (N_1593,In_684,In_396);
or U1594 (N_1594,In_708,In_736);
and U1595 (N_1595,In_526,In_962);
nor U1596 (N_1596,In_997,In_663);
and U1597 (N_1597,In_218,In_451);
xor U1598 (N_1598,In_167,In_459);
or U1599 (N_1599,In_363,In_192);
or U1600 (N_1600,In_402,In_765);
xnor U1601 (N_1601,In_577,In_628);
and U1602 (N_1602,In_516,In_964);
nand U1603 (N_1603,In_576,In_512);
or U1604 (N_1604,In_873,In_902);
xnor U1605 (N_1605,In_890,In_537);
nand U1606 (N_1606,In_986,In_341);
and U1607 (N_1607,In_537,In_237);
nor U1608 (N_1608,In_362,In_56);
nand U1609 (N_1609,In_937,In_268);
or U1610 (N_1610,In_866,In_926);
nor U1611 (N_1611,In_381,In_794);
or U1612 (N_1612,In_462,In_80);
nand U1613 (N_1613,In_678,In_306);
xor U1614 (N_1614,In_153,In_679);
nor U1615 (N_1615,In_36,In_371);
xnor U1616 (N_1616,In_78,In_217);
nor U1617 (N_1617,In_626,In_100);
nor U1618 (N_1618,In_239,In_565);
or U1619 (N_1619,In_494,In_336);
or U1620 (N_1620,In_920,In_805);
nor U1621 (N_1621,In_883,In_836);
nor U1622 (N_1622,In_512,In_961);
and U1623 (N_1623,In_993,In_163);
nand U1624 (N_1624,In_972,In_975);
nor U1625 (N_1625,In_646,In_306);
or U1626 (N_1626,In_750,In_692);
and U1627 (N_1627,In_453,In_175);
nand U1628 (N_1628,In_863,In_565);
nor U1629 (N_1629,In_466,In_244);
nand U1630 (N_1630,In_594,In_312);
nor U1631 (N_1631,In_256,In_681);
and U1632 (N_1632,In_157,In_315);
and U1633 (N_1633,In_20,In_73);
and U1634 (N_1634,In_245,In_597);
nand U1635 (N_1635,In_399,In_746);
xnor U1636 (N_1636,In_606,In_829);
and U1637 (N_1637,In_604,In_274);
and U1638 (N_1638,In_945,In_612);
nand U1639 (N_1639,In_817,In_150);
and U1640 (N_1640,In_938,In_243);
or U1641 (N_1641,In_724,In_79);
xnor U1642 (N_1642,In_573,In_535);
or U1643 (N_1643,In_864,In_303);
or U1644 (N_1644,In_596,In_752);
nand U1645 (N_1645,In_677,In_375);
or U1646 (N_1646,In_698,In_92);
nand U1647 (N_1647,In_963,In_989);
and U1648 (N_1648,In_213,In_786);
nand U1649 (N_1649,In_510,In_982);
xnor U1650 (N_1650,In_177,In_458);
nor U1651 (N_1651,In_385,In_921);
or U1652 (N_1652,In_202,In_405);
xor U1653 (N_1653,In_996,In_870);
and U1654 (N_1654,In_19,In_104);
or U1655 (N_1655,In_46,In_572);
nand U1656 (N_1656,In_451,In_694);
xor U1657 (N_1657,In_58,In_0);
nand U1658 (N_1658,In_426,In_911);
or U1659 (N_1659,In_121,In_645);
or U1660 (N_1660,In_413,In_585);
xnor U1661 (N_1661,In_221,In_957);
or U1662 (N_1662,In_766,In_659);
nand U1663 (N_1663,In_393,In_637);
and U1664 (N_1664,In_314,In_117);
or U1665 (N_1665,In_277,In_550);
nand U1666 (N_1666,In_583,In_631);
nand U1667 (N_1667,In_601,In_292);
and U1668 (N_1668,In_273,In_706);
or U1669 (N_1669,In_188,In_185);
and U1670 (N_1670,In_985,In_649);
nor U1671 (N_1671,In_337,In_82);
nor U1672 (N_1672,In_963,In_523);
nor U1673 (N_1673,In_928,In_943);
or U1674 (N_1674,In_734,In_326);
and U1675 (N_1675,In_470,In_290);
nor U1676 (N_1676,In_512,In_556);
nand U1677 (N_1677,In_105,In_52);
and U1678 (N_1678,In_786,In_843);
and U1679 (N_1679,In_856,In_682);
nand U1680 (N_1680,In_319,In_959);
nor U1681 (N_1681,In_582,In_56);
xnor U1682 (N_1682,In_12,In_693);
nand U1683 (N_1683,In_597,In_60);
nor U1684 (N_1684,In_602,In_588);
and U1685 (N_1685,In_281,In_650);
nand U1686 (N_1686,In_261,In_175);
nor U1687 (N_1687,In_198,In_210);
or U1688 (N_1688,In_633,In_881);
nand U1689 (N_1689,In_381,In_469);
or U1690 (N_1690,In_874,In_117);
nand U1691 (N_1691,In_764,In_473);
or U1692 (N_1692,In_0,In_743);
nor U1693 (N_1693,In_176,In_527);
and U1694 (N_1694,In_289,In_379);
or U1695 (N_1695,In_516,In_967);
nor U1696 (N_1696,In_785,In_199);
xnor U1697 (N_1697,In_581,In_647);
or U1698 (N_1698,In_544,In_56);
and U1699 (N_1699,In_450,In_837);
or U1700 (N_1700,In_196,In_149);
nor U1701 (N_1701,In_318,In_188);
and U1702 (N_1702,In_885,In_6);
or U1703 (N_1703,In_373,In_377);
nor U1704 (N_1704,In_12,In_787);
nand U1705 (N_1705,In_722,In_578);
nor U1706 (N_1706,In_491,In_974);
xor U1707 (N_1707,In_269,In_532);
or U1708 (N_1708,In_832,In_181);
or U1709 (N_1709,In_396,In_536);
or U1710 (N_1710,In_173,In_906);
or U1711 (N_1711,In_585,In_95);
xnor U1712 (N_1712,In_922,In_205);
nor U1713 (N_1713,In_143,In_615);
and U1714 (N_1714,In_717,In_166);
nand U1715 (N_1715,In_5,In_577);
nand U1716 (N_1716,In_385,In_308);
nand U1717 (N_1717,In_717,In_320);
and U1718 (N_1718,In_502,In_254);
nor U1719 (N_1719,In_394,In_884);
nor U1720 (N_1720,In_342,In_806);
nand U1721 (N_1721,In_112,In_348);
nor U1722 (N_1722,In_778,In_947);
and U1723 (N_1723,In_588,In_913);
or U1724 (N_1724,In_559,In_450);
or U1725 (N_1725,In_814,In_56);
nor U1726 (N_1726,In_483,In_699);
and U1727 (N_1727,In_795,In_425);
nand U1728 (N_1728,In_304,In_637);
nor U1729 (N_1729,In_65,In_516);
and U1730 (N_1730,In_848,In_4);
nand U1731 (N_1731,In_729,In_339);
nand U1732 (N_1732,In_388,In_509);
and U1733 (N_1733,In_434,In_29);
nand U1734 (N_1734,In_368,In_459);
nor U1735 (N_1735,In_877,In_943);
or U1736 (N_1736,In_174,In_586);
and U1737 (N_1737,In_823,In_895);
nand U1738 (N_1738,In_372,In_675);
nand U1739 (N_1739,In_285,In_243);
and U1740 (N_1740,In_259,In_445);
or U1741 (N_1741,In_468,In_447);
or U1742 (N_1742,In_921,In_660);
nor U1743 (N_1743,In_894,In_839);
nand U1744 (N_1744,In_865,In_353);
and U1745 (N_1745,In_330,In_238);
and U1746 (N_1746,In_181,In_877);
or U1747 (N_1747,In_752,In_348);
and U1748 (N_1748,In_446,In_828);
xnor U1749 (N_1749,In_192,In_73);
nor U1750 (N_1750,In_210,In_142);
or U1751 (N_1751,In_245,In_109);
and U1752 (N_1752,In_6,In_463);
nand U1753 (N_1753,In_590,In_51);
nor U1754 (N_1754,In_448,In_447);
nor U1755 (N_1755,In_405,In_465);
nand U1756 (N_1756,In_179,In_261);
nand U1757 (N_1757,In_938,In_198);
nor U1758 (N_1758,In_83,In_207);
and U1759 (N_1759,In_512,In_483);
and U1760 (N_1760,In_12,In_232);
nand U1761 (N_1761,In_936,In_547);
xor U1762 (N_1762,In_595,In_318);
nand U1763 (N_1763,In_834,In_592);
nand U1764 (N_1764,In_968,In_525);
or U1765 (N_1765,In_332,In_870);
and U1766 (N_1766,In_430,In_973);
and U1767 (N_1767,In_485,In_369);
xor U1768 (N_1768,In_787,In_859);
or U1769 (N_1769,In_461,In_307);
nand U1770 (N_1770,In_550,In_319);
and U1771 (N_1771,In_61,In_786);
xnor U1772 (N_1772,In_936,In_865);
nor U1773 (N_1773,In_426,In_14);
or U1774 (N_1774,In_86,In_64);
or U1775 (N_1775,In_117,In_758);
or U1776 (N_1776,In_241,In_400);
nand U1777 (N_1777,In_913,In_886);
or U1778 (N_1778,In_854,In_283);
nor U1779 (N_1779,In_236,In_766);
and U1780 (N_1780,In_692,In_10);
nand U1781 (N_1781,In_196,In_498);
and U1782 (N_1782,In_163,In_16);
and U1783 (N_1783,In_393,In_419);
and U1784 (N_1784,In_65,In_677);
xor U1785 (N_1785,In_928,In_754);
nor U1786 (N_1786,In_473,In_117);
nor U1787 (N_1787,In_891,In_847);
nor U1788 (N_1788,In_106,In_62);
or U1789 (N_1789,In_539,In_593);
or U1790 (N_1790,In_553,In_396);
or U1791 (N_1791,In_873,In_73);
or U1792 (N_1792,In_553,In_394);
and U1793 (N_1793,In_619,In_1);
nor U1794 (N_1794,In_589,In_522);
xor U1795 (N_1795,In_802,In_53);
xnor U1796 (N_1796,In_878,In_526);
nor U1797 (N_1797,In_778,In_64);
nor U1798 (N_1798,In_611,In_264);
nor U1799 (N_1799,In_884,In_923);
or U1800 (N_1800,In_783,In_502);
and U1801 (N_1801,In_14,In_20);
nand U1802 (N_1802,In_678,In_574);
xnor U1803 (N_1803,In_560,In_35);
and U1804 (N_1804,In_572,In_392);
and U1805 (N_1805,In_178,In_760);
nand U1806 (N_1806,In_622,In_955);
or U1807 (N_1807,In_781,In_685);
xor U1808 (N_1808,In_700,In_261);
nor U1809 (N_1809,In_638,In_603);
nand U1810 (N_1810,In_876,In_566);
nor U1811 (N_1811,In_50,In_236);
nand U1812 (N_1812,In_14,In_995);
nor U1813 (N_1813,In_585,In_915);
or U1814 (N_1814,In_947,In_601);
nand U1815 (N_1815,In_245,In_127);
nand U1816 (N_1816,In_316,In_39);
nor U1817 (N_1817,In_510,In_747);
nand U1818 (N_1818,In_709,In_713);
or U1819 (N_1819,In_184,In_249);
xor U1820 (N_1820,In_99,In_234);
nor U1821 (N_1821,In_647,In_492);
nand U1822 (N_1822,In_954,In_888);
nand U1823 (N_1823,In_816,In_912);
or U1824 (N_1824,In_569,In_257);
nand U1825 (N_1825,In_202,In_251);
or U1826 (N_1826,In_287,In_79);
nand U1827 (N_1827,In_719,In_328);
nand U1828 (N_1828,In_321,In_841);
and U1829 (N_1829,In_79,In_62);
nor U1830 (N_1830,In_367,In_867);
nand U1831 (N_1831,In_972,In_425);
nand U1832 (N_1832,In_118,In_591);
nor U1833 (N_1833,In_329,In_698);
nand U1834 (N_1834,In_486,In_599);
nor U1835 (N_1835,In_985,In_251);
and U1836 (N_1836,In_267,In_433);
or U1837 (N_1837,In_667,In_534);
and U1838 (N_1838,In_260,In_899);
or U1839 (N_1839,In_970,In_904);
or U1840 (N_1840,In_898,In_955);
and U1841 (N_1841,In_366,In_219);
and U1842 (N_1842,In_621,In_988);
nand U1843 (N_1843,In_345,In_514);
and U1844 (N_1844,In_102,In_391);
nor U1845 (N_1845,In_196,In_511);
nor U1846 (N_1846,In_418,In_336);
nand U1847 (N_1847,In_647,In_548);
and U1848 (N_1848,In_173,In_567);
and U1849 (N_1849,In_926,In_227);
or U1850 (N_1850,In_591,In_394);
or U1851 (N_1851,In_822,In_854);
or U1852 (N_1852,In_34,In_805);
nor U1853 (N_1853,In_696,In_27);
nor U1854 (N_1854,In_584,In_342);
or U1855 (N_1855,In_863,In_206);
xnor U1856 (N_1856,In_166,In_762);
xor U1857 (N_1857,In_249,In_151);
and U1858 (N_1858,In_85,In_943);
and U1859 (N_1859,In_977,In_558);
and U1860 (N_1860,In_341,In_717);
or U1861 (N_1861,In_166,In_393);
and U1862 (N_1862,In_979,In_77);
xor U1863 (N_1863,In_188,In_665);
nand U1864 (N_1864,In_743,In_133);
nand U1865 (N_1865,In_511,In_867);
or U1866 (N_1866,In_432,In_514);
nor U1867 (N_1867,In_752,In_928);
and U1868 (N_1868,In_224,In_220);
nand U1869 (N_1869,In_887,In_436);
nor U1870 (N_1870,In_39,In_459);
nor U1871 (N_1871,In_571,In_590);
nor U1872 (N_1872,In_775,In_402);
or U1873 (N_1873,In_808,In_28);
xnor U1874 (N_1874,In_852,In_154);
and U1875 (N_1875,In_397,In_251);
nand U1876 (N_1876,In_958,In_92);
and U1877 (N_1877,In_860,In_758);
and U1878 (N_1878,In_68,In_157);
nor U1879 (N_1879,In_490,In_474);
nand U1880 (N_1880,In_862,In_77);
or U1881 (N_1881,In_505,In_538);
or U1882 (N_1882,In_989,In_38);
and U1883 (N_1883,In_651,In_929);
and U1884 (N_1884,In_945,In_189);
or U1885 (N_1885,In_540,In_823);
nor U1886 (N_1886,In_795,In_64);
nand U1887 (N_1887,In_256,In_3);
nand U1888 (N_1888,In_351,In_173);
nor U1889 (N_1889,In_160,In_147);
or U1890 (N_1890,In_977,In_700);
or U1891 (N_1891,In_454,In_277);
and U1892 (N_1892,In_820,In_11);
nand U1893 (N_1893,In_795,In_615);
xor U1894 (N_1894,In_574,In_237);
or U1895 (N_1895,In_167,In_130);
nand U1896 (N_1896,In_231,In_440);
or U1897 (N_1897,In_298,In_241);
nor U1898 (N_1898,In_464,In_723);
and U1899 (N_1899,In_664,In_694);
and U1900 (N_1900,In_856,In_257);
nand U1901 (N_1901,In_187,In_361);
xnor U1902 (N_1902,In_514,In_421);
xnor U1903 (N_1903,In_441,In_826);
or U1904 (N_1904,In_79,In_121);
or U1905 (N_1905,In_564,In_319);
or U1906 (N_1906,In_865,In_808);
nor U1907 (N_1907,In_613,In_35);
xor U1908 (N_1908,In_380,In_553);
nor U1909 (N_1909,In_132,In_255);
nor U1910 (N_1910,In_294,In_519);
nand U1911 (N_1911,In_854,In_853);
nor U1912 (N_1912,In_612,In_931);
and U1913 (N_1913,In_914,In_608);
nor U1914 (N_1914,In_997,In_782);
nand U1915 (N_1915,In_90,In_654);
or U1916 (N_1916,In_732,In_633);
and U1917 (N_1917,In_581,In_689);
nor U1918 (N_1918,In_310,In_923);
nand U1919 (N_1919,In_971,In_41);
nand U1920 (N_1920,In_667,In_408);
and U1921 (N_1921,In_11,In_621);
nand U1922 (N_1922,In_989,In_424);
nor U1923 (N_1923,In_401,In_189);
or U1924 (N_1924,In_97,In_205);
and U1925 (N_1925,In_331,In_736);
nand U1926 (N_1926,In_130,In_119);
nand U1927 (N_1927,In_501,In_127);
nor U1928 (N_1928,In_542,In_390);
nand U1929 (N_1929,In_150,In_367);
or U1930 (N_1930,In_692,In_207);
nand U1931 (N_1931,In_698,In_125);
and U1932 (N_1932,In_2,In_797);
or U1933 (N_1933,In_76,In_192);
or U1934 (N_1934,In_599,In_256);
or U1935 (N_1935,In_918,In_854);
nor U1936 (N_1936,In_555,In_735);
or U1937 (N_1937,In_350,In_645);
nor U1938 (N_1938,In_331,In_608);
or U1939 (N_1939,In_378,In_21);
xnor U1940 (N_1940,In_874,In_642);
nor U1941 (N_1941,In_990,In_177);
nand U1942 (N_1942,In_947,In_644);
or U1943 (N_1943,In_341,In_120);
nand U1944 (N_1944,In_684,In_817);
nor U1945 (N_1945,In_703,In_433);
nor U1946 (N_1946,In_975,In_706);
and U1947 (N_1947,In_565,In_793);
nor U1948 (N_1948,In_448,In_8);
nor U1949 (N_1949,In_252,In_722);
and U1950 (N_1950,In_993,In_31);
xor U1951 (N_1951,In_847,In_65);
and U1952 (N_1952,In_422,In_89);
and U1953 (N_1953,In_784,In_340);
or U1954 (N_1954,In_32,In_784);
or U1955 (N_1955,In_571,In_954);
nor U1956 (N_1956,In_472,In_206);
xor U1957 (N_1957,In_437,In_90);
and U1958 (N_1958,In_571,In_435);
xnor U1959 (N_1959,In_178,In_118);
xnor U1960 (N_1960,In_669,In_993);
nand U1961 (N_1961,In_832,In_499);
or U1962 (N_1962,In_523,In_881);
nor U1963 (N_1963,In_232,In_915);
and U1964 (N_1964,In_139,In_459);
or U1965 (N_1965,In_564,In_639);
and U1966 (N_1966,In_726,In_70);
nor U1967 (N_1967,In_866,In_992);
and U1968 (N_1968,In_319,In_665);
nand U1969 (N_1969,In_146,In_203);
and U1970 (N_1970,In_892,In_363);
nand U1971 (N_1971,In_758,In_111);
nor U1972 (N_1972,In_472,In_800);
or U1973 (N_1973,In_119,In_938);
and U1974 (N_1974,In_458,In_369);
or U1975 (N_1975,In_707,In_334);
or U1976 (N_1976,In_590,In_770);
nand U1977 (N_1977,In_911,In_217);
nor U1978 (N_1978,In_446,In_891);
xor U1979 (N_1979,In_132,In_266);
nand U1980 (N_1980,In_471,In_906);
xnor U1981 (N_1981,In_513,In_101);
xor U1982 (N_1982,In_285,In_229);
nor U1983 (N_1983,In_613,In_459);
nor U1984 (N_1984,In_653,In_784);
nor U1985 (N_1985,In_685,In_604);
or U1986 (N_1986,In_127,In_652);
nor U1987 (N_1987,In_316,In_294);
nor U1988 (N_1988,In_311,In_914);
xor U1989 (N_1989,In_920,In_499);
and U1990 (N_1990,In_752,In_855);
nor U1991 (N_1991,In_119,In_296);
nor U1992 (N_1992,In_534,In_659);
xor U1993 (N_1993,In_887,In_947);
xor U1994 (N_1994,In_671,In_933);
nand U1995 (N_1995,In_598,In_816);
nand U1996 (N_1996,In_503,In_580);
nand U1997 (N_1997,In_151,In_21);
and U1998 (N_1998,In_277,In_95);
nand U1999 (N_1999,In_727,In_400);
nor U2000 (N_2000,In_331,In_723);
and U2001 (N_2001,In_949,In_115);
nand U2002 (N_2002,In_590,In_774);
nand U2003 (N_2003,In_779,In_138);
and U2004 (N_2004,In_763,In_492);
or U2005 (N_2005,In_118,In_717);
or U2006 (N_2006,In_416,In_786);
and U2007 (N_2007,In_557,In_547);
xor U2008 (N_2008,In_273,In_345);
nor U2009 (N_2009,In_51,In_553);
nand U2010 (N_2010,In_852,In_694);
xnor U2011 (N_2011,In_148,In_489);
nand U2012 (N_2012,In_627,In_523);
nand U2013 (N_2013,In_475,In_984);
nand U2014 (N_2014,In_809,In_554);
nor U2015 (N_2015,In_957,In_88);
and U2016 (N_2016,In_790,In_36);
and U2017 (N_2017,In_296,In_950);
nand U2018 (N_2018,In_276,In_279);
or U2019 (N_2019,In_571,In_285);
or U2020 (N_2020,In_700,In_816);
xnor U2021 (N_2021,In_785,In_758);
and U2022 (N_2022,In_998,In_340);
nor U2023 (N_2023,In_188,In_720);
nand U2024 (N_2024,In_185,In_114);
xnor U2025 (N_2025,In_914,In_842);
or U2026 (N_2026,In_726,In_852);
and U2027 (N_2027,In_617,In_627);
nand U2028 (N_2028,In_16,In_794);
nor U2029 (N_2029,In_648,In_813);
nand U2030 (N_2030,In_486,In_875);
or U2031 (N_2031,In_804,In_429);
or U2032 (N_2032,In_229,In_158);
or U2033 (N_2033,In_65,In_12);
nand U2034 (N_2034,In_187,In_27);
nor U2035 (N_2035,In_312,In_692);
nor U2036 (N_2036,In_255,In_241);
and U2037 (N_2037,In_196,In_577);
xnor U2038 (N_2038,In_655,In_57);
nand U2039 (N_2039,In_778,In_940);
or U2040 (N_2040,In_789,In_218);
xor U2041 (N_2041,In_228,In_226);
nor U2042 (N_2042,In_643,In_920);
nor U2043 (N_2043,In_387,In_533);
or U2044 (N_2044,In_514,In_921);
or U2045 (N_2045,In_606,In_480);
or U2046 (N_2046,In_850,In_353);
and U2047 (N_2047,In_253,In_573);
and U2048 (N_2048,In_288,In_513);
and U2049 (N_2049,In_21,In_27);
xor U2050 (N_2050,In_99,In_52);
and U2051 (N_2051,In_68,In_815);
nor U2052 (N_2052,In_250,In_327);
nor U2053 (N_2053,In_469,In_157);
nor U2054 (N_2054,In_545,In_961);
and U2055 (N_2055,In_840,In_751);
nor U2056 (N_2056,In_659,In_101);
and U2057 (N_2057,In_799,In_310);
nand U2058 (N_2058,In_56,In_394);
xnor U2059 (N_2059,In_440,In_22);
nor U2060 (N_2060,In_696,In_856);
nor U2061 (N_2061,In_37,In_209);
nor U2062 (N_2062,In_47,In_894);
or U2063 (N_2063,In_59,In_315);
and U2064 (N_2064,In_430,In_894);
nor U2065 (N_2065,In_440,In_758);
or U2066 (N_2066,In_498,In_520);
or U2067 (N_2067,In_79,In_539);
and U2068 (N_2068,In_804,In_7);
and U2069 (N_2069,In_809,In_397);
nand U2070 (N_2070,In_827,In_763);
nand U2071 (N_2071,In_695,In_691);
nor U2072 (N_2072,In_244,In_874);
nor U2073 (N_2073,In_559,In_235);
xnor U2074 (N_2074,In_96,In_402);
or U2075 (N_2075,In_693,In_532);
or U2076 (N_2076,In_476,In_392);
and U2077 (N_2077,In_105,In_980);
nand U2078 (N_2078,In_948,In_340);
and U2079 (N_2079,In_392,In_935);
nand U2080 (N_2080,In_111,In_120);
nor U2081 (N_2081,In_172,In_117);
nor U2082 (N_2082,In_653,In_889);
and U2083 (N_2083,In_220,In_7);
xnor U2084 (N_2084,In_744,In_25);
and U2085 (N_2085,In_611,In_182);
nor U2086 (N_2086,In_262,In_470);
xnor U2087 (N_2087,In_41,In_735);
or U2088 (N_2088,In_913,In_543);
and U2089 (N_2089,In_298,In_357);
nand U2090 (N_2090,In_181,In_836);
and U2091 (N_2091,In_235,In_433);
and U2092 (N_2092,In_119,In_860);
nor U2093 (N_2093,In_656,In_914);
nand U2094 (N_2094,In_226,In_230);
or U2095 (N_2095,In_126,In_178);
and U2096 (N_2096,In_583,In_718);
nand U2097 (N_2097,In_929,In_322);
and U2098 (N_2098,In_380,In_243);
nor U2099 (N_2099,In_465,In_858);
nand U2100 (N_2100,In_247,In_594);
xnor U2101 (N_2101,In_102,In_520);
or U2102 (N_2102,In_773,In_969);
nand U2103 (N_2103,In_77,In_818);
nand U2104 (N_2104,In_740,In_737);
or U2105 (N_2105,In_194,In_542);
and U2106 (N_2106,In_502,In_202);
nor U2107 (N_2107,In_90,In_465);
nor U2108 (N_2108,In_73,In_446);
and U2109 (N_2109,In_354,In_651);
or U2110 (N_2110,In_436,In_746);
xnor U2111 (N_2111,In_742,In_959);
and U2112 (N_2112,In_849,In_556);
nor U2113 (N_2113,In_265,In_952);
and U2114 (N_2114,In_358,In_535);
and U2115 (N_2115,In_414,In_154);
xor U2116 (N_2116,In_717,In_791);
or U2117 (N_2117,In_704,In_587);
or U2118 (N_2118,In_732,In_729);
nand U2119 (N_2119,In_217,In_352);
nand U2120 (N_2120,In_965,In_227);
xor U2121 (N_2121,In_99,In_778);
nand U2122 (N_2122,In_176,In_808);
nor U2123 (N_2123,In_742,In_708);
nand U2124 (N_2124,In_328,In_86);
or U2125 (N_2125,In_407,In_234);
or U2126 (N_2126,In_542,In_600);
nor U2127 (N_2127,In_329,In_716);
or U2128 (N_2128,In_631,In_777);
xnor U2129 (N_2129,In_307,In_532);
nand U2130 (N_2130,In_934,In_770);
nor U2131 (N_2131,In_959,In_936);
or U2132 (N_2132,In_336,In_607);
nand U2133 (N_2133,In_12,In_987);
and U2134 (N_2134,In_623,In_359);
and U2135 (N_2135,In_427,In_54);
or U2136 (N_2136,In_946,In_151);
or U2137 (N_2137,In_667,In_71);
nor U2138 (N_2138,In_100,In_822);
nand U2139 (N_2139,In_481,In_64);
or U2140 (N_2140,In_732,In_523);
nor U2141 (N_2141,In_719,In_584);
or U2142 (N_2142,In_829,In_44);
nor U2143 (N_2143,In_419,In_505);
and U2144 (N_2144,In_901,In_541);
xnor U2145 (N_2145,In_299,In_863);
and U2146 (N_2146,In_432,In_540);
or U2147 (N_2147,In_686,In_362);
and U2148 (N_2148,In_956,In_810);
nor U2149 (N_2149,In_633,In_420);
and U2150 (N_2150,In_140,In_276);
and U2151 (N_2151,In_947,In_287);
and U2152 (N_2152,In_960,In_564);
or U2153 (N_2153,In_640,In_403);
nor U2154 (N_2154,In_515,In_894);
and U2155 (N_2155,In_673,In_818);
nor U2156 (N_2156,In_837,In_30);
and U2157 (N_2157,In_695,In_587);
and U2158 (N_2158,In_583,In_113);
and U2159 (N_2159,In_15,In_166);
xor U2160 (N_2160,In_18,In_75);
nand U2161 (N_2161,In_476,In_801);
or U2162 (N_2162,In_51,In_579);
and U2163 (N_2163,In_897,In_160);
xnor U2164 (N_2164,In_371,In_715);
and U2165 (N_2165,In_678,In_589);
nor U2166 (N_2166,In_427,In_936);
nor U2167 (N_2167,In_918,In_527);
nor U2168 (N_2168,In_710,In_566);
and U2169 (N_2169,In_592,In_797);
nand U2170 (N_2170,In_948,In_802);
or U2171 (N_2171,In_339,In_506);
xor U2172 (N_2172,In_97,In_315);
nand U2173 (N_2173,In_152,In_559);
nand U2174 (N_2174,In_708,In_650);
nor U2175 (N_2175,In_303,In_915);
and U2176 (N_2176,In_573,In_333);
or U2177 (N_2177,In_782,In_726);
or U2178 (N_2178,In_653,In_817);
or U2179 (N_2179,In_510,In_835);
or U2180 (N_2180,In_270,In_288);
and U2181 (N_2181,In_710,In_736);
nor U2182 (N_2182,In_687,In_252);
and U2183 (N_2183,In_701,In_899);
xnor U2184 (N_2184,In_139,In_297);
xor U2185 (N_2185,In_258,In_861);
or U2186 (N_2186,In_787,In_858);
or U2187 (N_2187,In_373,In_873);
nor U2188 (N_2188,In_830,In_468);
or U2189 (N_2189,In_863,In_960);
nor U2190 (N_2190,In_612,In_183);
nand U2191 (N_2191,In_454,In_239);
and U2192 (N_2192,In_929,In_543);
and U2193 (N_2193,In_438,In_888);
or U2194 (N_2194,In_626,In_949);
and U2195 (N_2195,In_976,In_140);
nor U2196 (N_2196,In_288,In_683);
and U2197 (N_2197,In_861,In_333);
xnor U2198 (N_2198,In_199,In_828);
nand U2199 (N_2199,In_586,In_355);
nor U2200 (N_2200,In_29,In_839);
nor U2201 (N_2201,In_257,In_122);
nor U2202 (N_2202,In_530,In_513);
or U2203 (N_2203,In_461,In_79);
or U2204 (N_2204,In_788,In_899);
and U2205 (N_2205,In_270,In_179);
nor U2206 (N_2206,In_84,In_592);
or U2207 (N_2207,In_896,In_475);
nor U2208 (N_2208,In_274,In_285);
nor U2209 (N_2209,In_415,In_904);
xor U2210 (N_2210,In_966,In_762);
or U2211 (N_2211,In_994,In_9);
or U2212 (N_2212,In_231,In_928);
and U2213 (N_2213,In_993,In_271);
nand U2214 (N_2214,In_146,In_14);
xnor U2215 (N_2215,In_492,In_464);
nor U2216 (N_2216,In_974,In_95);
or U2217 (N_2217,In_833,In_982);
nand U2218 (N_2218,In_537,In_914);
and U2219 (N_2219,In_69,In_905);
nor U2220 (N_2220,In_310,In_674);
or U2221 (N_2221,In_143,In_586);
nand U2222 (N_2222,In_45,In_527);
nand U2223 (N_2223,In_217,In_730);
nand U2224 (N_2224,In_149,In_854);
xor U2225 (N_2225,In_648,In_542);
nand U2226 (N_2226,In_424,In_529);
or U2227 (N_2227,In_581,In_571);
or U2228 (N_2228,In_409,In_676);
or U2229 (N_2229,In_148,In_661);
and U2230 (N_2230,In_28,In_406);
nor U2231 (N_2231,In_197,In_265);
nand U2232 (N_2232,In_17,In_84);
nor U2233 (N_2233,In_467,In_995);
nor U2234 (N_2234,In_30,In_656);
and U2235 (N_2235,In_16,In_306);
nand U2236 (N_2236,In_231,In_180);
nor U2237 (N_2237,In_338,In_99);
nand U2238 (N_2238,In_148,In_998);
nor U2239 (N_2239,In_98,In_232);
or U2240 (N_2240,In_459,In_33);
nand U2241 (N_2241,In_654,In_855);
or U2242 (N_2242,In_682,In_122);
nand U2243 (N_2243,In_178,In_799);
and U2244 (N_2244,In_308,In_562);
and U2245 (N_2245,In_805,In_457);
and U2246 (N_2246,In_230,In_59);
nand U2247 (N_2247,In_926,In_691);
and U2248 (N_2248,In_749,In_121);
or U2249 (N_2249,In_667,In_878);
and U2250 (N_2250,In_737,In_998);
or U2251 (N_2251,In_749,In_889);
nand U2252 (N_2252,In_494,In_552);
xnor U2253 (N_2253,In_411,In_140);
or U2254 (N_2254,In_871,In_261);
and U2255 (N_2255,In_793,In_678);
or U2256 (N_2256,In_935,In_123);
or U2257 (N_2257,In_256,In_203);
nor U2258 (N_2258,In_421,In_107);
or U2259 (N_2259,In_362,In_441);
or U2260 (N_2260,In_317,In_178);
nand U2261 (N_2261,In_100,In_300);
or U2262 (N_2262,In_850,In_638);
nor U2263 (N_2263,In_131,In_871);
or U2264 (N_2264,In_952,In_541);
and U2265 (N_2265,In_309,In_975);
nor U2266 (N_2266,In_900,In_446);
or U2267 (N_2267,In_806,In_410);
nor U2268 (N_2268,In_806,In_54);
xnor U2269 (N_2269,In_303,In_502);
and U2270 (N_2270,In_904,In_203);
or U2271 (N_2271,In_334,In_547);
nand U2272 (N_2272,In_617,In_323);
and U2273 (N_2273,In_12,In_458);
nor U2274 (N_2274,In_513,In_709);
and U2275 (N_2275,In_133,In_563);
and U2276 (N_2276,In_982,In_933);
or U2277 (N_2277,In_908,In_971);
or U2278 (N_2278,In_74,In_418);
nand U2279 (N_2279,In_351,In_21);
or U2280 (N_2280,In_660,In_377);
and U2281 (N_2281,In_247,In_535);
nor U2282 (N_2282,In_587,In_839);
and U2283 (N_2283,In_926,In_178);
or U2284 (N_2284,In_157,In_155);
xnor U2285 (N_2285,In_130,In_76);
nand U2286 (N_2286,In_719,In_351);
nor U2287 (N_2287,In_590,In_39);
nor U2288 (N_2288,In_206,In_841);
or U2289 (N_2289,In_735,In_129);
nor U2290 (N_2290,In_461,In_986);
and U2291 (N_2291,In_827,In_712);
xnor U2292 (N_2292,In_875,In_894);
xnor U2293 (N_2293,In_709,In_169);
and U2294 (N_2294,In_263,In_387);
or U2295 (N_2295,In_623,In_901);
or U2296 (N_2296,In_71,In_991);
nor U2297 (N_2297,In_478,In_790);
nor U2298 (N_2298,In_720,In_628);
or U2299 (N_2299,In_201,In_995);
xnor U2300 (N_2300,In_368,In_422);
nand U2301 (N_2301,In_350,In_946);
or U2302 (N_2302,In_206,In_98);
nor U2303 (N_2303,In_746,In_181);
or U2304 (N_2304,In_179,In_156);
nand U2305 (N_2305,In_989,In_980);
nor U2306 (N_2306,In_469,In_219);
xnor U2307 (N_2307,In_468,In_475);
nand U2308 (N_2308,In_560,In_722);
nor U2309 (N_2309,In_955,In_71);
nor U2310 (N_2310,In_383,In_169);
and U2311 (N_2311,In_452,In_937);
nor U2312 (N_2312,In_836,In_760);
xnor U2313 (N_2313,In_234,In_854);
nor U2314 (N_2314,In_13,In_561);
and U2315 (N_2315,In_542,In_555);
nor U2316 (N_2316,In_23,In_818);
or U2317 (N_2317,In_350,In_222);
nor U2318 (N_2318,In_722,In_665);
and U2319 (N_2319,In_464,In_781);
nor U2320 (N_2320,In_970,In_733);
and U2321 (N_2321,In_433,In_681);
nor U2322 (N_2322,In_213,In_730);
nor U2323 (N_2323,In_399,In_99);
nand U2324 (N_2324,In_654,In_342);
nand U2325 (N_2325,In_27,In_342);
or U2326 (N_2326,In_692,In_463);
and U2327 (N_2327,In_866,In_431);
and U2328 (N_2328,In_731,In_356);
nand U2329 (N_2329,In_359,In_852);
and U2330 (N_2330,In_271,In_789);
nor U2331 (N_2331,In_358,In_961);
or U2332 (N_2332,In_131,In_432);
and U2333 (N_2333,In_498,In_597);
or U2334 (N_2334,In_231,In_492);
and U2335 (N_2335,In_68,In_127);
or U2336 (N_2336,In_102,In_997);
or U2337 (N_2337,In_22,In_248);
and U2338 (N_2338,In_796,In_169);
nand U2339 (N_2339,In_949,In_375);
nor U2340 (N_2340,In_995,In_935);
or U2341 (N_2341,In_226,In_425);
nor U2342 (N_2342,In_888,In_479);
or U2343 (N_2343,In_682,In_659);
xnor U2344 (N_2344,In_279,In_274);
nor U2345 (N_2345,In_126,In_214);
xnor U2346 (N_2346,In_240,In_730);
nor U2347 (N_2347,In_216,In_975);
or U2348 (N_2348,In_384,In_383);
nand U2349 (N_2349,In_290,In_904);
nand U2350 (N_2350,In_264,In_959);
nor U2351 (N_2351,In_81,In_520);
and U2352 (N_2352,In_808,In_23);
nor U2353 (N_2353,In_416,In_721);
nand U2354 (N_2354,In_555,In_958);
nand U2355 (N_2355,In_660,In_302);
nand U2356 (N_2356,In_94,In_722);
and U2357 (N_2357,In_479,In_36);
and U2358 (N_2358,In_839,In_568);
and U2359 (N_2359,In_937,In_815);
and U2360 (N_2360,In_141,In_557);
and U2361 (N_2361,In_288,In_320);
xnor U2362 (N_2362,In_940,In_867);
and U2363 (N_2363,In_995,In_96);
xor U2364 (N_2364,In_413,In_105);
nor U2365 (N_2365,In_384,In_982);
nor U2366 (N_2366,In_466,In_572);
or U2367 (N_2367,In_244,In_706);
xnor U2368 (N_2368,In_251,In_252);
nand U2369 (N_2369,In_995,In_967);
and U2370 (N_2370,In_449,In_496);
nand U2371 (N_2371,In_242,In_138);
nor U2372 (N_2372,In_77,In_236);
or U2373 (N_2373,In_601,In_68);
nand U2374 (N_2374,In_926,In_311);
or U2375 (N_2375,In_494,In_91);
and U2376 (N_2376,In_265,In_637);
and U2377 (N_2377,In_324,In_616);
and U2378 (N_2378,In_423,In_776);
xor U2379 (N_2379,In_687,In_547);
xnor U2380 (N_2380,In_677,In_585);
and U2381 (N_2381,In_853,In_751);
and U2382 (N_2382,In_934,In_73);
or U2383 (N_2383,In_368,In_388);
or U2384 (N_2384,In_623,In_592);
nand U2385 (N_2385,In_917,In_82);
xnor U2386 (N_2386,In_951,In_813);
nand U2387 (N_2387,In_118,In_752);
nand U2388 (N_2388,In_947,In_82);
or U2389 (N_2389,In_22,In_883);
nor U2390 (N_2390,In_702,In_863);
nor U2391 (N_2391,In_682,In_232);
nor U2392 (N_2392,In_643,In_130);
or U2393 (N_2393,In_63,In_505);
nand U2394 (N_2394,In_888,In_316);
nand U2395 (N_2395,In_902,In_379);
nor U2396 (N_2396,In_660,In_983);
and U2397 (N_2397,In_35,In_884);
nand U2398 (N_2398,In_649,In_307);
or U2399 (N_2399,In_331,In_363);
xnor U2400 (N_2400,In_884,In_347);
nand U2401 (N_2401,In_319,In_8);
nor U2402 (N_2402,In_767,In_685);
nor U2403 (N_2403,In_819,In_205);
nor U2404 (N_2404,In_8,In_900);
nor U2405 (N_2405,In_72,In_10);
nor U2406 (N_2406,In_727,In_812);
or U2407 (N_2407,In_48,In_803);
or U2408 (N_2408,In_174,In_536);
or U2409 (N_2409,In_404,In_21);
or U2410 (N_2410,In_725,In_236);
nor U2411 (N_2411,In_1,In_692);
nor U2412 (N_2412,In_566,In_468);
and U2413 (N_2413,In_951,In_836);
and U2414 (N_2414,In_176,In_324);
nor U2415 (N_2415,In_845,In_732);
xnor U2416 (N_2416,In_778,In_330);
nand U2417 (N_2417,In_208,In_569);
and U2418 (N_2418,In_839,In_326);
and U2419 (N_2419,In_853,In_710);
and U2420 (N_2420,In_918,In_340);
or U2421 (N_2421,In_267,In_143);
or U2422 (N_2422,In_806,In_799);
and U2423 (N_2423,In_144,In_456);
or U2424 (N_2424,In_552,In_973);
nor U2425 (N_2425,In_566,In_371);
or U2426 (N_2426,In_143,In_581);
and U2427 (N_2427,In_876,In_941);
or U2428 (N_2428,In_631,In_474);
and U2429 (N_2429,In_737,In_49);
xor U2430 (N_2430,In_467,In_241);
xor U2431 (N_2431,In_791,In_684);
nand U2432 (N_2432,In_200,In_238);
or U2433 (N_2433,In_896,In_493);
xnor U2434 (N_2434,In_353,In_14);
and U2435 (N_2435,In_726,In_394);
and U2436 (N_2436,In_43,In_881);
xor U2437 (N_2437,In_137,In_209);
or U2438 (N_2438,In_578,In_201);
nor U2439 (N_2439,In_784,In_211);
nor U2440 (N_2440,In_648,In_195);
nor U2441 (N_2441,In_37,In_533);
and U2442 (N_2442,In_410,In_263);
xor U2443 (N_2443,In_958,In_188);
nor U2444 (N_2444,In_935,In_926);
or U2445 (N_2445,In_513,In_326);
nor U2446 (N_2446,In_770,In_578);
or U2447 (N_2447,In_206,In_699);
or U2448 (N_2448,In_725,In_585);
nand U2449 (N_2449,In_393,In_241);
nor U2450 (N_2450,In_724,In_291);
or U2451 (N_2451,In_21,In_762);
or U2452 (N_2452,In_532,In_287);
or U2453 (N_2453,In_251,In_416);
or U2454 (N_2454,In_934,In_881);
nand U2455 (N_2455,In_120,In_988);
or U2456 (N_2456,In_182,In_623);
and U2457 (N_2457,In_182,In_664);
nor U2458 (N_2458,In_389,In_495);
or U2459 (N_2459,In_227,In_905);
nor U2460 (N_2460,In_574,In_169);
or U2461 (N_2461,In_420,In_336);
nor U2462 (N_2462,In_950,In_940);
nor U2463 (N_2463,In_278,In_375);
and U2464 (N_2464,In_28,In_509);
nor U2465 (N_2465,In_152,In_27);
or U2466 (N_2466,In_7,In_344);
and U2467 (N_2467,In_487,In_302);
xor U2468 (N_2468,In_83,In_626);
and U2469 (N_2469,In_510,In_417);
and U2470 (N_2470,In_921,In_980);
nor U2471 (N_2471,In_692,In_228);
nor U2472 (N_2472,In_195,In_137);
nand U2473 (N_2473,In_980,In_323);
nor U2474 (N_2474,In_541,In_752);
or U2475 (N_2475,In_501,In_686);
nand U2476 (N_2476,In_717,In_556);
or U2477 (N_2477,In_575,In_479);
and U2478 (N_2478,In_625,In_961);
nand U2479 (N_2479,In_379,In_479);
nand U2480 (N_2480,In_719,In_660);
nor U2481 (N_2481,In_950,In_665);
xnor U2482 (N_2482,In_590,In_908);
nand U2483 (N_2483,In_285,In_829);
nand U2484 (N_2484,In_346,In_817);
and U2485 (N_2485,In_257,In_558);
nor U2486 (N_2486,In_158,In_495);
nor U2487 (N_2487,In_497,In_93);
and U2488 (N_2488,In_358,In_380);
nor U2489 (N_2489,In_138,In_596);
nor U2490 (N_2490,In_313,In_291);
or U2491 (N_2491,In_151,In_209);
or U2492 (N_2492,In_159,In_71);
nand U2493 (N_2493,In_325,In_32);
xor U2494 (N_2494,In_61,In_319);
nand U2495 (N_2495,In_344,In_352);
nor U2496 (N_2496,In_394,In_756);
xor U2497 (N_2497,In_783,In_594);
and U2498 (N_2498,In_424,In_521);
nor U2499 (N_2499,In_324,In_737);
xor U2500 (N_2500,In_663,In_551);
and U2501 (N_2501,In_818,In_464);
nand U2502 (N_2502,In_686,In_451);
nand U2503 (N_2503,In_322,In_987);
and U2504 (N_2504,In_714,In_165);
nand U2505 (N_2505,In_684,In_649);
xor U2506 (N_2506,In_454,In_200);
nor U2507 (N_2507,In_138,In_472);
nor U2508 (N_2508,In_66,In_447);
and U2509 (N_2509,In_850,In_466);
or U2510 (N_2510,In_936,In_351);
or U2511 (N_2511,In_473,In_233);
nor U2512 (N_2512,In_514,In_593);
and U2513 (N_2513,In_46,In_813);
nand U2514 (N_2514,In_185,In_66);
or U2515 (N_2515,In_698,In_561);
nor U2516 (N_2516,In_633,In_45);
nand U2517 (N_2517,In_310,In_27);
or U2518 (N_2518,In_945,In_607);
and U2519 (N_2519,In_463,In_796);
and U2520 (N_2520,In_674,In_569);
nor U2521 (N_2521,In_137,In_975);
or U2522 (N_2522,In_737,In_636);
nor U2523 (N_2523,In_671,In_687);
nand U2524 (N_2524,In_757,In_41);
or U2525 (N_2525,In_735,In_347);
nor U2526 (N_2526,In_423,In_120);
and U2527 (N_2527,In_348,In_814);
nor U2528 (N_2528,In_268,In_81);
nor U2529 (N_2529,In_636,In_717);
nand U2530 (N_2530,In_550,In_736);
and U2531 (N_2531,In_242,In_298);
or U2532 (N_2532,In_714,In_362);
or U2533 (N_2533,In_857,In_172);
xnor U2534 (N_2534,In_546,In_959);
or U2535 (N_2535,In_457,In_575);
nor U2536 (N_2536,In_984,In_688);
nor U2537 (N_2537,In_645,In_493);
nand U2538 (N_2538,In_617,In_300);
and U2539 (N_2539,In_287,In_514);
nand U2540 (N_2540,In_673,In_327);
xnor U2541 (N_2541,In_613,In_819);
nand U2542 (N_2542,In_598,In_433);
nor U2543 (N_2543,In_304,In_814);
and U2544 (N_2544,In_461,In_947);
and U2545 (N_2545,In_658,In_248);
nand U2546 (N_2546,In_44,In_864);
or U2547 (N_2547,In_329,In_24);
and U2548 (N_2548,In_885,In_37);
or U2549 (N_2549,In_219,In_451);
nand U2550 (N_2550,In_161,In_552);
and U2551 (N_2551,In_577,In_436);
or U2552 (N_2552,In_941,In_505);
nand U2553 (N_2553,In_135,In_626);
nand U2554 (N_2554,In_297,In_991);
or U2555 (N_2555,In_715,In_465);
xor U2556 (N_2556,In_899,In_484);
xnor U2557 (N_2557,In_976,In_611);
nor U2558 (N_2558,In_327,In_868);
and U2559 (N_2559,In_244,In_16);
or U2560 (N_2560,In_2,In_755);
nand U2561 (N_2561,In_806,In_656);
nand U2562 (N_2562,In_419,In_552);
nor U2563 (N_2563,In_596,In_233);
or U2564 (N_2564,In_897,In_605);
nand U2565 (N_2565,In_415,In_813);
nor U2566 (N_2566,In_901,In_225);
nand U2567 (N_2567,In_833,In_804);
nor U2568 (N_2568,In_370,In_337);
nand U2569 (N_2569,In_296,In_294);
nor U2570 (N_2570,In_851,In_888);
nand U2571 (N_2571,In_784,In_830);
nand U2572 (N_2572,In_391,In_815);
or U2573 (N_2573,In_202,In_719);
or U2574 (N_2574,In_560,In_483);
or U2575 (N_2575,In_110,In_219);
or U2576 (N_2576,In_527,In_612);
or U2577 (N_2577,In_959,In_33);
and U2578 (N_2578,In_566,In_587);
nor U2579 (N_2579,In_107,In_408);
xor U2580 (N_2580,In_609,In_76);
and U2581 (N_2581,In_505,In_658);
nor U2582 (N_2582,In_977,In_196);
nor U2583 (N_2583,In_227,In_966);
and U2584 (N_2584,In_672,In_639);
xor U2585 (N_2585,In_98,In_544);
nor U2586 (N_2586,In_785,In_94);
xnor U2587 (N_2587,In_439,In_196);
or U2588 (N_2588,In_884,In_364);
or U2589 (N_2589,In_538,In_357);
nor U2590 (N_2590,In_821,In_10);
nand U2591 (N_2591,In_905,In_554);
and U2592 (N_2592,In_787,In_191);
or U2593 (N_2593,In_834,In_283);
nor U2594 (N_2594,In_302,In_431);
and U2595 (N_2595,In_111,In_901);
nand U2596 (N_2596,In_737,In_193);
xnor U2597 (N_2597,In_78,In_404);
nor U2598 (N_2598,In_185,In_668);
and U2599 (N_2599,In_458,In_463);
xor U2600 (N_2600,In_364,In_944);
nand U2601 (N_2601,In_279,In_633);
or U2602 (N_2602,In_207,In_531);
nand U2603 (N_2603,In_359,In_845);
nor U2604 (N_2604,In_201,In_753);
and U2605 (N_2605,In_276,In_956);
or U2606 (N_2606,In_632,In_750);
or U2607 (N_2607,In_383,In_583);
nand U2608 (N_2608,In_913,In_263);
nor U2609 (N_2609,In_349,In_929);
or U2610 (N_2610,In_255,In_490);
nand U2611 (N_2611,In_991,In_881);
nand U2612 (N_2612,In_803,In_309);
nand U2613 (N_2613,In_66,In_799);
nand U2614 (N_2614,In_913,In_602);
or U2615 (N_2615,In_430,In_1);
or U2616 (N_2616,In_752,In_284);
nor U2617 (N_2617,In_793,In_885);
nor U2618 (N_2618,In_137,In_44);
or U2619 (N_2619,In_262,In_316);
or U2620 (N_2620,In_854,In_201);
nor U2621 (N_2621,In_941,In_812);
or U2622 (N_2622,In_954,In_401);
nand U2623 (N_2623,In_613,In_237);
and U2624 (N_2624,In_788,In_267);
nor U2625 (N_2625,In_834,In_620);
or U2626 (N_2626,In_786,In_569);
nand U2627 (N_2627,In_86,In_685);
and U2628 (N_2628,In_376,In_751);
nand U2629 (N_2629,In_596,In_99);
nand U2630 (N_2630,In_445,In_772);
xor U2631 (N_2631,In_567,In_770);
nand U2632 (N_2632,In_184,In_661);
or U2633 (N_2633,In_638,In_327);
and U2634 (N_2634,In_986,In_938);
and U2635 (N_2635,In_942,In_639);
nor U2636 (N_2636,In_197,In_516);
or U2637 (N_2637,In_116,In_908);
xor U2638 (N_2638,In_873,In_134);
nand U2639 (N_2639,In_857,In_34);
and U2640 (N_2640,In_204,In_806);
nor U2641 (N_2641,In_407,In_12);
nand U2642 (N_2642,In_298,In_78);
nand U2643 (N_2643,In_352,In_155);
and U2644 (N_2644,In_77,In_318);
or U2645 (N_2645,In_779,In_340);
or U2646 (N_2646,In_880,In_106);
nand U2647 (N_2647,In_67,In_919);
nor U2648 (N_2648,In_258,In_749);
nand U2649 (N_2649,In_397,In_29);
or U2650 (N_2650,In_941,In_153);
or U2651 (N_2651,In_307,In_143);
nor U2652 (N_2652,In_389,In_725);
nor U2653 (N_2653,In_745,In_427);
nor U2654 (N_2654,In_783,In_474);
nand U2655 (N_2655,In_747,In_206);
nand U2656 (N_2656,In_252,In_835);
nand U2657 (N_2657,In_150,In_332);
nor U2658 (N_2658,In_405,In_72);
nand U2659 (N_2659,In_792,In_994);
nand U2660 (N_2660,In_192,In_635);
and U2661 (N_2661,In_301,In_395);
and U2662 (N_2662,In_128,In_340);
nand U2663 (N_2663,In_150,In_402);
nor U2664 (N_2664,In_333,In_613);
and U2665 (N_2665,In_733,In_293);
xnor U2666 (N_2666,In_129,In_523);
and U2667 (N_2667,In_662,In_794);
or U2668 (N_2668,In_657,In_179);
nand U2669 (N_2669,In_569,In_541);
and U2670 (N_2670,In_577,In_95);
nand U2671 (N_2671,In_119,In_259);
nor U2672 (N_2672,In_224,In_573);
and U2673 (N_2673,In_605,In_594);
nand U2674 (N_2674,In_236,In_572);
nor U2675 (N_2675,In_613,In_756);
nand U2676 (N_2676,In_58,In_339);
or U2677 (N_2677,In_793,In_938);
and U2678 (N_2678,In_839,In_494);
or U2679 (N_2679,In_164,In_237);
or U2680 (N_2680,In_810,In_335);
and U2681 (N_2681,In_693,In_834);
nand U2682 (N_2682,In_270,In_14);
nand U2683 (N_2683,In_761,In_666);
or U2684 (N_2684,In_382,In_21);
nor U2685 (N_2685,In_252,In_588);
and U2686 (N_2686,In_458,In_366);
xnor U2687 (N_2687,In_427,In_547);
and U2688 (N_2688,In_357,In_443);
nand U2689 (N_2689,In_538,In_692);
or U2690 (N_2690,In_771,In_404);
nand U2691 (N_2691,In_689,In_899);
and U2692 (N_2692,In_404,In_208);
nor U2693 (N_2693,In_391,In_414);
nor U2694 (N_2694,In_408,In_507);
nor U2695 (N_2695,In_951,In_796);
nor U2696 (N_2696,In_843,In_75);
nand U2697 (N_2697,In_587,In_387);
or U2698 (N_2698,In_293,In_93);
nor U2699 (N_2699,In_556,In_195);
and U2700 (N_2700,In_456,In_892);
or U2701 (N_2701,In_467,In_696);
or U2702 (N_2702,In_650,In_249);
nand U2703 (N_2703,In_862,In_592);
nand U2704 (N_2704,In_52,In_322);
xor U2705 (N_2705,In_922,In_58);
nor U2706 (N_2706,In_873,In_535);
and U2707 (N_2707,In_615,In_653);
and U2708 (N_2708,In_827,In_172);
nor U2709 (N_2709,In_872,In_654);
or U2710 (N_2710,In_387,In_829);
nor U2711 (N_2711,In_501,In_98);
nand U2712 (N_2712,In_495,In_364);
nand U2713 (N_2713,In_111,In_436);
and U2714 (N_2714,In_204,In_25);
nor U2715 (N_2715,In_806,In_844);
or U2716 (N_2716,In_12,In_47);
or U2717 (N_2717,In_31,In_158);
nand U2718 (N_2718,In_830,In_961);
nor U2719 (N_2719,In_47,In_932);
and U2720 (N_2720,In_195,In_233);
nand U2721 (N_2721,In_364,In_124);
and U2722 (N_2722,In_575,In_180);
nor U2723 (N_2723,In_672,In_567);
nor U2724 (N_2724,In_386,In_114);
or U2725 (N_2725,In_117,In_551);
nor U2726 (N_2726,In_524,In_552);
and U2727 (N_2727,In_928,In_671);
and U2728 (N_2728,In_935,In_655);
and U2729 (N_2729,In_570,In_121);
nand U2730 (N_2730,In_161,In_685);
or U2731 (N_2731,In_739,In_736);
nand U2732 (N_2732,In_404,In_499);
nor U2733 (N_2733,In_83,In_104);
or U2734 (N_2734,In_517,In_319);
nand U2735 (N_2735,In_439,In_314);
nor U2736 (N_2736,In_185,In_430);
nand U2737 (N_2737,In_225,In_242);
and U2738 (N_2738,In_276,In_406);
nor U2739 (N_2739,In_66,In_976);
nor U2740 (N_2740,In_40,In_384);
nand U2741 (N_2741,In_56,In_175);
or U2742 (N_2742,In_214,In_453);
and U2743 (N_2743,In_137,In_82);
or U2744 (N_2744,In_29,In_455);
nand U2745 (N_2745,In_1,In_668);
and U2746 (N_2746,In_926,In_200);
nand U2747 (N_2747,In_426,In_293);
or U2748 (N_2748,In_683,In_906);
nor U2749 (N_2749,In_242,In_259);
nor U2750 (N_2750,In_246,In_669);
or U2751 (N_2751,In_915,In_894);
and U2752 (N_2752,In_903,In_774);
xnor U2753 (N_2753,In_803,In_246);
nor U2754 (N_2754,In_231,In_167);
or U2755 (N_2755,In_538,In_864);
and U2756 (N_2756,In_60,In_318);
or U2757 (N_2757,In_346,In_875);
and U2758 (N_2758,In_291,In_521);
nor U2759 (N_2759,In_691,In_619);
nand U2760 (N_2760,In_501,In_408);
or U2761 (N_2761,In_105,In_944);
nand U2762 (N_2762,In_170,In_555);
and U2763 (N_2763,In_162,In_86);
or U2764 (N_2764,In_867,In_568);
or U2765 (N_2765,In_479,In_621);
nor U2766 (N_2766,In_395,In_423);
or U2767 (N_2767,In_43,In_65);
or U2768 (N_2768,In_85,In_234);
nand U2769 (N_2769,In_824,In_952);
xnor U2770 (N_2770,In_135,In_703);
or U2771 (N_2771,In_162,In_373);
nor U2772 (N_2772,In_79,In_810);
xor U2773 (N_2773,In_861,In_336);
nand U2774 (N_2774,In_477,In_5);
nand U2775 (N_2775,In_581,In_827);
or U2776 (N_2776,In_901,In_600);
nor U2777 (N_2777,In_279,In_350);
nor U2778 (N_2778,In_404,In_550);
or U2779 (N_2779,In_945,In_706);
nor U2780 (N_2780,In_512,In_720);
nand U2781 (N_2781,In_453,In_723);
nor U2782 (N_2782,In_419,In_79);
nand U2783 (N_2783,In_542,In_508);
nor U2784 (N_2784,In_278,In_538);
nand U2785 (N_2785,In_481,In_449);
nand U2786 (N_2786,In_324,In_210);
and U2787 (N_2787,In_386,In_236);
and U2788 (N_2788,In_852,In_707);
xor U2789 (N_2789,In_317,In_25);
or U2790 (N_2790,In_673,In_864);
nand U2791 (N_2791,In_434,In_50);
and U2792 (N_2792,In_103,In_409);
nor U2793 (N_2793,In_556,In_166);
and U2794 (N_2794,In_505,In_617);
xor U2795 (N_2795,In_704,In_506);
nor U2796 (N_2796,In_335,In_771);
nor U2797 (N_2797,In_156,In_623);
nand U2798 (N_2798,In_707,In_452);
and U2799 (N_2799,In_331,In_416);
nor U2800 (N_2800,In_731,In_92);
xnor U2801 (N_2801,In_614,In_562);
nor U2802 (N_2802,In_802,In_856);
nand U2803 (N_2803,In_30,In_523);
and U2804 (N_2804,In_894,In_659);
nor U2805 (N_2805,In_946,In_564);
or U2806 (N_2806,In_227,In_626);
nand U2807 (N_2807,In_562,In_445);
and U2808 (N_2808,In_662,In_655);
or U2809 (N_2809,In_816,In_141);
or U2810 (N_2810,In_865,In_927);
and U2811 (N_2811,In_220,In_810);
or U2812 (N_2812,In_99,In_674);
nand U2813 (N_2813,In_938,In_654);
or U2814 (N_2814,In_544,In_295);
and U2815 (N_2815,In_113,In_799);
xnor U2816 (N_2816,In_132,In_72);
nand U2817 (N_2817,In_446,In_601);
and U2818 (N_2818,In_714,In_787);
or U2819 (N_2819,In_799,In_595);
or U2820 (N_2820,In_47,In_90);
nand U2821 (N_2821,In_433,In_377);
or U2822 (N_2822,In_296,In_824);
or U2823 (N_2823,In_369,In_647);
nand U2824 (N_2824,In_964,In_23);
nand U2825 (N_2825,In_379,In_897);
nand U2826 (N_2826,In_157,In_673);
and U2827 (N_2827,In_378,In_171);
nor U2828 (N_2828,In_346,In_355);
and U2829 (N_2829,In_758,In_532);
and U2830 (N_2830,In_110,In_449);
nand U2831 (N_2831,In_348,In_657);
or U2832 (N_2832,In_773,In_422);
and U2833 (N_2833,In_537,In_968);
nor U2834 (N_2834,In_487,In_380);
or U2835 (N_2835,In_934,In_585);
or U2836 (N_2836,In_694,In_338);
and U2837 (N_2837,In_78,In_13);
or U2838 (N_2838,In_766,In_418);
and U2839 (N_2839,In_648,In_100);
and U2840 (N_2840,In_238,In_578);
or U2841 (N_2841,In_871,In_816);
nor U2842 (N_2842,In_361,In_706);
xor U2843 (N_2843,In_611,In_880);
and U2844 (N_2844,In_575,In_969);
xor U2845 (N_2845,In_605,In_600);
xnor U2846 (N_2846,In_261,In_628);
nand U2847 (N_2847,In_299,In_435);
or U2848 (N_2848,In_861,In_906);
nand U2849 (N_2849,In_203,In_771);
xnor U2850 (N_2850,In_833,In_546);
or U2851 (N_2851,In_525,In_501);
nand U2852 (N_2852,In_982,In_644);
nand U2853 (N_2853,In_752,In_413);
or U2854 (N_2854,In_640,In_938);
nand U2855 (N_2855,In_728,In_726);
or U2856 (N_2856,In_564,In_113);
and U2857 (N_2857,In_256,In_281);
nor U2858 (N_2858,In_193,In_257);
nand U2859 (N_2859,In_280,In_487);
or U2860 (N_2860,In_877,In_878);
nor U2861 (N_2861,In_726,In_472);
or U2862 (N_2862,In_610,In_476);
or U2863 (N_2863,In_785,In_423);
and U2864 (N_2864,In_688,In_504);
or U2865 (N_2865,In_346,In_52);
and U2866 (N_2866,In_846,In_590);
nor U2867 (N_2867,In_572,In_564);
nand U2868 (N_2868,In_936,In_740);
nand U2869 (N_2869,In_987,In_65);
xnor U2870 (N_2870,In_437,In_206);
nor U2871 (N_2871,In_720,In_78);
xnor U2872 (N_2872,In_45,In_123);
and U2873 (N_2873,In_581,In_525);
and U2874 (N_2874,In_936,In_411);
and U2875 (N_2875,In_397,In_378);
nand U2876 (N_2876,In_123,In_888);
xnor U2877 (N_2877,In_95,In_796);
nand U2878 (N_2878,In_122,In_102);
or U2879 (N_2879,In_718,In_218);
and U2880 (N_2880,In_287,In_627);
and U2881 (N_2881,In_337,In_357);
nand U2882 (N_2882,In_989,In_898);
xnor U2883 (N_2883,In_323,In_477);
xnor U2884 (N_2884,In_198,In_800);
nor U2885 (N_2885,In_458,In_361);
nand U2886 (N_2886,In_245,In_397);
nand U2887 (N_2887,In_279,In_30);
nand U2888 (N_2888,In_793,In_740);
or U2889 (N_2889,In_278,In_846);
nor U2890 (N_2890,In_648,In_776);
or U2891 (N_2891,In_20,In_562);
nor U2892 (N_2892,In_719,In_869);
nor U2893 (N_2893,In_353,In_570);
nor U2894 (N_2894,In_754,In_33);
nand U2895 (N_2895,In_860,In_44);
nand U2896 (N_2896,In_367,In_54);
and U2897 (N_2897,In_893,In_669);
and U2898 (N_2898,In_401,In_886);
or U2899 (N_2899,In_222,In_243);
nand U2900 (N_2900,In_359,In_67);
or U2901 (N_2901,In_485,In_59);
xor U2902 (N_2902,In_467,In_905);
or U2903 (N_2903,In_631,In_565);
and U2904 (N_2904,In_113,In_933);
nor U2905 (N_2905,In_527,In_73);
and U2906 (N_2906,In_186,In_669);
nor U2907 (N_2907,In_130,In_698);
nand U2908 (N_2908,In_138,In_131);
xor U2909 (N_2909,In_28,In_69);
nor U2910 (N_2910,In_190,In_659);
or U2911 (N_2911,In_70,In_507);
nor U2912 (N_2912,In_977,In_221);
nor U2913 (N_2913,In_281,In_950);
nand U2914 (N_2914,In_473,In_260);
or U2915 (N_2915,In_555,In_124);
or U2916 (N_2916,In_869,In_746);
or U2917 (N_2917,In_299,In_520);
nand U2918 (N_2918,In_995,In_959);
or U2919 (N_2919,In_598,In_300);
nor U2920 (N_2920,In_996,In_233);
nand U2921 (N_2921,In_298,In_480);
nand U2922 (N_2922,In_478,In_866);
nor U2923 (N_2923,In_826,In_710);
nand U2924 (N_2924,In_559,In_374);
or U2925 (N_2925,In_196,In_897);
and U2926 (N_2926,In_715,In_494);
nor U2927 (N_2927,In_848,In_455);
and U2928 (N_2928,In_844,In_224);
and U2929 (N_2929,In_920,In_263);
nand U2930 (N_2930,In_74,In_34);
or U2931 (N_2931,In_916,In_529);
nor U2932 (N_2932,In_903,In_822);
or U2933 (N_2933,In_974,In_169);
xor U2934 (N_2934,In_624,In_317);
nor U2935 (N_2935,In_142,In_526);
nor U2936 (N_2936,In_567,In_384);
nand U2937 (N_2937,In_295,In_945);
and U2938 (N_2938,In_249,In_371);
nand U2939 (N_2939,In_895,In_546);
nand U2940 (N_2940,In_425,In_486);
or U2941 (N_2941,In_535,In_684);
nand U2942 (N_2942,In_343,In_974);
and U2943 (N_2943,In_41,In_655);
and U2944 (N_2944,In_978,In_238);
or U2945 (N_2945,In_381,In_88);
and U2946 (N_2946,In_807,In_589);
nor U2947 (N_2947,In_743,In_855);
and U2948 (N_2948,In_918,In_710);
nand U2949 (N_2949,In_619,In_193);
or U2950 (N_2950,In_638,In_901);
nor U2951 (N_2951,In_280,In_137);
nand U2952 (N_2952,In_235,In_732);
or U2953 (N_2953,In_523,In_796);
and U2954 (N_2954,In_765,In_320);
or U2955 (N_2955,In_588,In_803);
nor U2956 (N_2956,In_97,In_112);
and U2957 (N_2957,In_472,In_154);
and U2958 (N_2958,In_615,In_614);
nor U2959 (N_2959,In_866,In_600);
nor U2960 (N_2960,In_185,In_616);
or U2961 (N_2961,In_836,In_920);
and U2962 (N_2962,In_796,In_604);
or U2963 (N_2963,In_810,In_741);
nor U2964 (N_2964,In_830,In_634);
xor U2965 (N_2965,In_736,In_758);
nor U2966 (N_2966,In_952,In_960);
nor U2967 (N_2967,In_770,In_643);
nor U2968 (N_2968,In_922,In_530);
and U2969 (N_2969,In_653,In_171);
nand U2970 (N_2970,In_734,In_739);
nor U2971 (N_2971,In_376,In_888);
and U2972 (N_2972,In_600,In_46);
or U2973 (N_2973,In_531,In_127);
or U2974 (N_2974,In_444,In_778);
and U2975 (N_2975,In_457,In_416);
nand U2976 (N_2976,In_200,In_183);
and U2977 (N_2977,In_390,In_788);
and U2978 (N_2978,In_270,In_686);
nor U2979 (N_2979,In_308,In_7);
xor U2980 (N_2980,In_113,In_669);
and U2981 (N_2981,In_81,In_170);
nand U2982 (N_2982,In_567,In_535);
xnor U2983 (N_2983,In_341,In_419);
nand U2984 (N_2984,In_166,In_780);
or U2985 (N_2985,In_618,In_563);
nand U2986 (N_2986,In_542,In_943);
nor U2987 (N_2987,In_853,In_257);
nor U2988 (N_2988,In_838,In_66);
nand U2989 (N_2989,In_589,In_572);
and U2990 (N_2990,In_993,In_451);
nor U2991 (N_2991,In_23,In_19);
and U2992 (N_2992,In_819,In_634);
and U2993 (N_2993,In_271,In_131);
and U2994 (N_2994,In_413,In_227);
nor U2995 (N_2995,In_41,In_740);
nor U2996 (N_2996,In_75,In_575);
and U2997 (N_2997,In_477,In_458);
xnor U2998 (N_2998,In_555,In_770);
xnor U2999 (N_2999,In_344,In_153);
and U3000 (N_3000,In_41,In_496);
nor U3001 (N_3001,In_802,In_233);
and U3002 (N_3002,In_964,In_857);
or U3003 (N_3003,In_632,In_853);
and U3004 (N_3004,In_726,In_54);
nor U3005 (N_3005,In_228,In_610);
xor U3006 (N_3006,In_345,In_199);
nand U3007 (N_3007,In_561,In_34);
nand U3008 (N_3008,In_708,In_126);
and U3009 (N_3009,In_333,In_14);
and U3010 (N_3010,In_843,In_856);
nor U3011 (N_3011,In_820,In_152);
and U3012 (N_3012,In_220,In_590);
or U3013 (N_3013,In_642,In_52);
or U3014 (N_3014,In_558,In_80);
or U3015 (N_3015,In_865,In_6);
nand U3016 (N_3016,In_52,In_813);
nor U3017 (N_3017,In_893,In_291);
nand U3018 (N_3018,In_930,In_958);
or U3019 (N_3019,In_153,In_32);
or U3020 (N_3020,In_170,In_499);
or U3021 (N_3021,In_683,In_405);
nor U3022 (N_3022,In_727,In_954);
nor U3023 (N_3023,In_360,In_410);
and U3024 (N_3024,In_526,In_780);
xnor U3025 (N_3025,In_587,In_0);
nor U3026 (N_3026,In_778,In_271);
or U3027 (N_3027,In_485,In_454);
and U3028 (N_3028,In_849,In_161);
nand U3029 (N_3029,In_968,In_826);
xnor U3030 (N_3030,In_187,In_224);
nor U3031 (N_3031,In_278,In_465);
and U3032 (N_3032,In_48,In_644);
nand U3033 (N_3033,In_109,In_257);
and U3034 (N_3034,In_895,In_999);
and U3035 (N_3035,In_877,In_867);
and U3036 (N_3036,In_900,In_308);
or U3037 (N_3037,In_113,In_786);
or U3038 (N_3038,In_923,In_472);
and U3039 (N_3039,In_509,In_443);
nand U3040 (N_3040,In_53,In_758);
and U3041 (N_3041,In_562,In_840);
and U3042 (N_3042,In_9,In_148);
or U3043 (N_3043,In_223,In_63);
and U3044 (N_3044,In_428,In_634);
nor U3045 (N_3045,In_666,In_64);
and U3046 (N_3046,In_156,In_347);
nand U3047 (N_3047,In_417,In_777);
nor U3048 (N_3048,In_159,In_160);
or U3049 (N_3049,In_685,In_106);
or U3050 (N_3050,In_453,In_53);
nor U3051 (N_3051,In_882,In_985);
nor U3052 (N_3052,In_656,In_293);
and U3053 (N_3053,In_647,In_267);
and U3054 (N_3054,In_659,In_658);
and U3055 (N_3055,In_104,In_92);
or U3056 (N_3056,In_19,In_20);
nand U3057 (N_3057,In_230,In_920);
nand U3058 (N_3058,In_299,In_677);
or U3059 (N_3059,In_892,In_118);
and U3060 (N_3060,In_569,In_770);
and U3061 (N_3061,In_541,In_44);
nor U3062 (N_3062,In_575,In_522);
and U3063 (N_3063,In_554,In_268);
nand U3064 (N_3064,In_802,In_885);
nand U3065 (N_3065,In_423,In_865);
nand U3066 (N_3066,In_134,In_953);
and U3067 (N_3067,In_621,In_656);
nand U3068 (N_3068,In_168,In_653);
nand U3069 (N_3069,In_454,In_222);
xnor U3070 (N_3070,In_285,In_417);
nor U3071 (N_3071,In_555,In_923);
or U3072 (N_3072,In_563,In_401);
or U3073 (N_3073,In_597,In_371);
xnor U3074 (N_3074,In_223,In_872);
and U3075 (N_3075,In_96,In_409);
nor U3076 (N_3076,In_480,In_29);
and U3077 (N_3077,In_893,In_903);
or U3078 (N_3078,In_970,In_513);
nor U3079 (N_3079,In_274,In_298);
and U3080 (N_3080,In_559,In_457);
nor U3081 (N_3081,In_474,In_48);
nand U3082 (N_3082,In_564,In_257);
nor U3083 (N_3083,In_495,In_271);
or U3084 (N_3084,In_801,In_981);
and U3085 (N_3085,In_585,In_456);
xor U3086 (N_3086,In_237,In_837);
or U3087 (N_3087,In_553,In_340);
and U3088 (N_3088,In_68,In_998);
xnor U3089 (N_3089,In_356,In_283);
nor U3090 (N_3090,In_985,In_461);
nand U3091 (N_3091,In_351,In_95);
or U3092 (N_3092,In_322,In_32);
or U3093 (N_3093,In_123,In_379);
and U3094 (N_3094,In_447,In_408);
and U3095 (N_3095,In_4,In_608);
xnor U3096 (N_3096,In_834,In_200);
nor U3097 (N_3097,In_795,In_843);
or U3098 (N_3098,In_838,In_684);
or U3099 (N_3099,In_795,In_30);
or U3100 (N_3100,In_584,In_997);
nand U3101 (N_3101,In_336,In_772);
or U3102 (N_3102,In_600,In_911);
nand U3103 (N_3103,In_634,In_799);
nand U3104 (N_3104,In_401,In_860);
xor U3105 (N_3105,In_53,In_105);
or U3106 (N_3106,In_819,In_898);
and U3107 (N_3107,In_432,In_858);
nand U3108 (N_3108,In_1,In_113);
nor U3109 (N_3109,In_292,In_217);
and U3110 (N_3110,In_932,In_700);
xor U3111 (N_3111,In_614,In_387);
nand U3112 (N_3112,In_947,In_368);
and U3113 (N_3113,In_488,In_530);
and U3114 (N_3114,In_915,In_626);
nand U3115 (N_3115,In_719,In_560);
and U3116 (N_3116,In_823,In_727);
and U3117 (N_3117,In_432,In_71);
and U3118 (N_3118,In_905,In_536);
xnor U3119 (N_3119,In_7,In_402);
and U3120 (N_3120,In_805,In_503);
and U3121 (N_3121,In_102,In_584);
nor U3122 (N_3122,In_99,In_148);
and U3123 (N_3123,In_686,In_167);
nor U3124 (N_3124,In_820,In_808);
and U3125 (N_3125,In_661,In_452);
or U3126 (N_3126,In_923,In_169);
nor U3127 (N_3127,In_688,In_64);
nand U3128 (N_3128,In_267,In_558);
nor U3129 (N_3129,In_761,In_68);
nor U3130 (N_3130,In_460,In_723);
nor U3131 (N_3131,In_599,In_947);
and U3132 (N_3132,In_42,In_629);
xor U3133 (N_3133,In_986,In_1);
nand U3134 (N_3134,In_804,In_513);
nor U3135 (N_3135,In_511,In_801);
nor U3136 (N_3136,In_433,In_740);
nand U3137 (N_3137,In_89,In_966);
or U3138 (N_3138,In_636,In_732);
xor U3139 (N_3139,In_700,In_494);
or U3140 (N_3140,In_525,In_470);
nand U3141 (N_3141,In_802,In_533);
nand U3142 (N_3142,In_25,In_576);
nor U3143 (N_3143,In_909,In_211);
xor U3144 (N_3144,In_271,In_664);
nor U3145 (N_3145,In_820,In_40);
nand U3146 (N_3146,In_187,In_695);
and U3147 (N_3147,In_561,In_873);
and U3148 (N_3148,In_479,In_436);
nor U3149 (N_3149,In_302,In_3);
or U3150 (N_3150,In_154,In_365);
or U3151 (N_3151,In_926,In_314);
nor U3152 (N_3152,In_117,In_612);
nor U3153 (N_3153,In_145,In_844);
or U3154 (N_3154,In_403,In_774);
nand U3155 (N_3155,In_915,In_172);
or U3156 (N_3156,In_176,In_500);
nor U3157 (N_3157,In_922,In_970);
or U3158 (N_3158,In_396,In_616);
nand U3159 (N_3159,In_180,In_688);
nand U3160 (N_3160,In_949,In_440);
and U3161 (N_3161,In_873,In_110);
and U3162 (N_3162,In_339,In_581);
nor U3163 (N_3163,In_551,In_789);
nor U3164 (N_3164,In_599,In_269);
xnor U3165 (N_3165,In_417,In_899);
nor U3166 (N_3166,In_475,In_547);
or U3167 (N_3167,In_467,In_982);
and U3168 (N_3168,In_633,In_72);
nand U3169 (N_3169,In_957,In_275);
nand U3170 (N_3170,In_703,In_376);
and U3171 (N_3171,In_36,In_757);
or U3172 (N_3172,In_336,In_175);
nand U3173 (N_3173,In_479,In_322);
and U3174 (N_3174,In_246,In_958);
or U3175 (N_3175,In_883,In_199);
and U3176 (N_3176,In_851,In_204);
or U3177 (N_3177,In_99,In_292);
xnor U3178 (N_3178,In_560,In_869);
and U3179 (N_3179,In_994,In_485);
nor U3180 (N_3180,In_269,In_84);
and U3181 (N_3181,In_370,In_628);
and U3182 (N_3182,In_664,In_818);
and U3183 (N_3183,In_683,In_212);
nor U3184 (N_3184,In_650,In_115);
or U3185 (N_3185,In_782,In_353);
nor U3186 (N_3186,In_839,In_184);
nor U3187 (N_3187,In_117,In_192);
nor U3188 (N_3188,In_701,In_391);
and U3189 (N_3189,In_545,In_188);
nor U3190 (N_3190,In_330,In_142);
xor U3191 (N_3191,In_37,In_823);
xor U3192 (N_3192,In_262,In_130);
and U3193 (N_3193,In_549,In_135);
nand U3194 (N_3194,In_143,In_629);
nand U3195 (N_3195,In_475,In_377);
xor U3196 (N_3196,In_998,In_94);
nor U3197 (N_3197,In_53,In_61);
xnor U3198 (N_3198,In_545,In_347);
and U3199 (N_3199,In_343,In_321);
nand U3200 (N_3200,In_480,In_323);
and U3201 (N_3201,In_812,In_569);
nor U3202 (N_3202,In_500,In_895);
and U3203 (N_3203,In_356,In_585);
or U3204 (N_3204,In_898,In_51);
nand U3205 (N_3205,In_542,In_467);
and U3206 (N_3206,In_350,In_339);
and U3207 (N_3207,In_300,In_524);
and U3208 (N_3208,In_221,In_244);
or U3209 (N_3209,In_381,In_155);
or U3210 (N_3210,In_644,In_252);
or U3211 (N_3211,In_311,In_416);
or U3212 (N_3212,In_51,In_311);
and U3213 (N_3213,In_231,In_31);
nor U3214 (N_3214,In_436,In_358);
or U3215 (N_3215,In_424,In_115);
and U3216 (N_3216,In_982,In_810);
nand U3217 (N_3217,In_663,In_220);
and U3218 (N_3218,In_305,In_679);
nand U3219 (N_3219,In_846,In_318);
nand U3220 (N_3220,In_664,In_978);
and U3221 (N_3221,In_899,In_441);
xnor U3222 (N_3222,In_645,In_875);
or U3223 (N_3223,In_426,In_601);
or U3224 (N_3224,In_445,In_996);
or U3225 (N_3225,In_73,In_658);
nor U3226 (N_3226,In_389,In_494);
or U3227 (N_3227,In_943,In_702);
nand U3228 (N_3228,In_410,In_988);
nor U3229 (N_3229,In_620,In_698);
nand U3230 (N_3230,In_86,In_23);
xnor U3231 (N_3231,In_486,In_455);
and U3232 (N_3232,In_514,In_585);
nand U3233 (N_3233,In_449,In_841);
nand U3234 (N_3234,In_996,In_647);
nand U3235 (N_3235,In_926,In_385);
and U3236 (N_3236,In_66,In_49);
nor U3237 (N_3237,In_884,In_667);
nand U3238 (N_3238,In_937,In_892);
or U3239 (N_3239,In_615,In_385);
xor U3240 (N_3240,In_840,In_795);
and U3241 (N_3241,In_636,In_555);
or U3242 (N_3242,In_171,In_248);
xnor U3243 (N_3243,In_725,In_663);
and U3244 (N_3244,In_337,In_592);
nand U3245 (N_3245,In_549,In_270);
or U3246 (N_3246,In_392,In_204);
nand U3247 (N_3247,In_934,In_911);
or U3248 (N_3248,In_669,In_782);
nor U3249 (N_3249,In_844,In_750);
nand U3250 (N_3250,In_232,In_127);
or U3251 (N_3251,In_41,In_327);
xor U3252 (N_3252,In_700,In_338);
nand U3253 (N_3253,In_931,In_175);
or U3254 (N_3254,In_620,In_933);
nor U3255 (N_3255,In_737,In_663);
and U3256 (N_3256,In_789,In_556);
and U3257 (N_3257,In_383,In_909);
and U3258 (N_3258,In_351,In_904);
or U3259 (N_3259,In_787,In_87);
nand U3260 (N_3260,In_121,In_497);
nand U3261 (N_3261,In_450,In_161);
and U3262 (N_3262,In_681,In_96);
or U3263 (N_3263,In_224,In_452);
nor U3264 (N_3264,In_591,In_294);
xnor U3265 (N_3265,In_271,In_511);
or U3266 (N_3266,In_715,In_253);
or U3267 (N_3267,In_44,In_547);
and U3268 (N_3268,In_536,In_864);
nand U3269 (N_3269,In_30,In_47);
nor U3270 (N_3270,In_826,In_433);
nand U3271 (N_3271,In_74,In_151);
nor U3272 (N_3272,In_736,In_852);
or U3273 (N_3273,In_867,In_861);
or U3274 (N_3274,In_302,In_234);
or U3275 (N_3275,In_956,In_185);
nand U3276 (N_3276,In_276,In_40);
nand U3277 (N_3277,In_697,In_880);
or U3278 (N_3278,In_408,In_12);
and U3279 (N_3279,In_328,In_346);
or U3280 (N_3280,In_939,In_340);
and U3281 (N_3281,In_604,In_293);
nor U3282 (N_3282,In_816,In_773);
nor U3283 (N_3283,In_681,In_758);
nor U3284 (N_3284,In_732,In_17);
or U3285 (N_3285,In_254,In_387);
or U3286 (N_3286,In_793,In_692);
nand U3287 (N_3287,In_581,In_507);
and U3288 (N_3288,In_818,In_983);
or U3289 (N_3289,In_275,In_48);
or U3290 (N_3290,In_695,In_217);
nor U3291 (N_3291,In_369,In_393);
and U3292 (N_3292,In_563,In_276);
nor U3293 (N_3293,In_736,In_294);
or U3294 (N_3294,In_383,In_643);
or U3295 (N_3295,In_871,In_32);
or U3296 (N_3296,In_263,In_976);
and U3297 (N_3297,In_724,In_823);
and U3298 (N_3298,In_771,In_289);
or U3299 (N_3299,In_180,In_558);
nand U3300 (N_3300,In_797,In_187);
nand U3301 (N_3301,In_158,In_841);
nor U3302 (N_3302,In_580,In_353);
nor U3303 (N_3303,In_422,In_405);
nand U3304 (N_3304,In_948,In_412);
nand U3305 (N_3305,In_356,In_825);
xor U3306 (N_3306,In_931,In_944);
and U3307 (N_3307,In_86,In_245);
or U3308 (N_3308,In_765,In_148);
or U3309 (N_3309,In_534,In_734);
xor U3310 (N_3310,In_39,In_455);
or U3311 (N_3311,In_613,In_252);
and U3312 (N_3312,In_621,In_222);
xor U3313 (N_3313,In_965,In_398);
or U3314 (N_3314,In_217,In_623);
xnor U3315 (N_3315,In_68,In_891);
nor U3316 (N_3316,In_110,In_460);
or U3317 (N_3317,In_199,In_830);
or U3318 (N_3318,In_670,In_605);
and U3319 (N_3319,In_403,In_16);
or U3320 (N_3320,In_511,In_157);
or U3321 (N_3321,In_434,In_333);
nor U3322 (N_3322,In_441,In_546);
and U3323 (N_3323,In_251,In_566);
and U3324 (N_3324,In_455,In_240);
nor U3325 (N_3325,In_670,In_389);
and U3326 (N_3326,In_92,In_455);
or U3327 (N_3327,In_994,In_462);
nand U3328 (N_3328,In_584,In_511);
nand U3329 (N_3329,In_731,In_270);
nor U3330 (N_3330,In_797,In_317);
and U3331 (N_3331,In_442,In_598);
xnor U3332 (N_3332,In_966,In_106);
and U3333 (N_3333,In_792,In_714);
xnor U3334 (N_3334,In_245,In_392);
nor U3335 (N_3335,In_642,In_803);
nand U3336 (N_3336,In_740,In_679);
xor U3337 (N_3337,In_741,In_884);
and U3338 (N_3338,In_164,In_234);
nor U3339 (N_3339,In_780,In_160);
and U3340 (N_3340,In_87,In_36);
xor U3341 (N_3341,In_515,In_170);
nor U3342 (N_3342,In_369,In_164);
nand U3343 (N_3343,In_715,In_205);
and U3344 (N_3344,In_980,In_424);
or U3345 (N_3345,In_975,In_639);
or U3346 (N_3346,In_242,In_895);
and U3347 (N_3347,In_123,In_86);
or U3348 (N_3348,In_900,In_462);
nor U3349 (N_3349,In_674,In_370);
and U3350 (N_3350,In_827,In_422);
nor U3351 (N_3351,In_301,In_892);
and U3352 (N_3352,In_924,In_649);
nand U3353 (N_3353,In_812,In_649);
and U3354 (N_3354,In_818,In_253);
or U3355 (N_3355,In_516,In_533);
and U3356 (N_3356,In_499,In_787);
xnor U3357 (N_3357,In_241,In_994);
or U3358 (N_3358,In_407,In_564);
or U3359 (N_3359,In_67,In_524);
nand U3360 (N_3360,In_848,In_898);
nand U3361 (N_3361,In_477,In_864);
and U3362 (N_3362,In_481,In_62);
and U3363 (N_3363,In_987,In_772);
nor U3364 (N_3364,In_360,In_702);
nor U3365 (N_3365,In_345,In_267);
xnor U3366 (N_3366,In_502,In_240);
or U3367 (N_3367,In_205,In_445);
nor U3368 (N_3368,In_282,In_638);
or U3369 (N_3369,In_317,In_41);
nor U3370 (N_3370,In_461,In_466);
nor U3371 (N_3371,In_119,In_977);
xnor U3372 (N_3372,In_949,In_370);
and U3373 (N_3373,In_284,In_475);
nand U3374 (N_3374,In_960,In_950);
nor U3375 (N_3375,In_574,In_558);
nand U3376 (N_3376,In_903,In_634);
and U3377 (N_3377,In_214,In_612);
xnor U3378 (N_3378,In_686,In_572);
or U3379 (N_3379,In_488,In_28);
and U3380 (N_3380,In_65,In_877);
or U3381 (N_3381,In_699,In_123);
and U3382 (N_3382,In_462,In_745);
nor U3383 (N_3383,In_831,In_186);
nor U3384 (N_3384,In_177,In_532);
or U3385 (N_3385,In_576,In_335);
or U3386 (N_3386,In_969,In_672);
xnor U3387 (N_3387,In_774,In_602);
or U3388 (N_3388,In_216,In_522);
nor U3389 (N_3389,In_367,In_115);
or U3390 (N_3390,In_556,In_748);
nand U3391 (N_3391,In_376,In_55);
and U3392 (N_3392,In_96,In_252);
xor U3393 (N_3393,In_518,In_574);
and U3394 (N_3394,In_306,In_245);
nor U3395 (N_3395,In_342,In_191);
xor U3396 (N_3396,In_329,In_431);
or U3397 (N_3397,In_533,In_738);
nor U3398 (N_3398,In_29,In_417);
and U3399 (N_3399,In_964,In_555);
nor U3400 (N_3400,In_844,In_267);
nand U3401 (N_3401,In_436,In_972);
or U3402 (N_3402,In_784,In_650);
or U3403 (N_3403,In_571,In_654);
and U3404 (N_3404,In_634,In_559);
xor U3405 (N_3405,In_782,In_823);
or U3406 (N_3406,In_581,In_197);
nor U3407 (N_3407,In_575,In_253);
or U3408 (N_3408,In_664,In_234);
and U3409 (N_3409,In_199,In_620);
xor U3410 (N_3410,In_676,In_822);
and U3411 (N_3411,In_767,In_725);
and U3412 (N_3412,In_61,In_889);
and U3413 (N_3413,In_508,In_97);
nor U3414 (N_3414,In_241,In_554);
nand U3415 (N_3415,In_370,In_440);
or U3416 (N_3416,In_638,In_214);
nand U3417 (N_3417,In_898,In_838);
and U3418 (N_3418,In_79,In_693);
or U3419 (N_3419,In_776,In_319);
or U3420 (N_3420,In_974,In_821);
and U3421 (N_3421,In_122,In_623);
or U3422 (N_3422,In_228,In_184);
or U3423 (N_3423,In_730,In_983);
nand U3424 (N_3424,In_440,In_918);
nand U3425 (N_3425,In_892,In_532);
or U3426 (N_3426,In_771,In_503);
or U3427 (N_3427,In_54,In_556);
xnor U3428 (N_3428,In_813,In_387);
xor U3429 (N_3429,In_276,In_289);
nor U3430 (N_3430,In_993,In_745);
nor U3431 (N_3431,In_367,In_120);
or U3432 (N_3432,In_778,In_954);
xor U3433 (N_3433,In_760,In_378);
nand U3434 (N_3434,In_131,In_562);
nand U3435 (N_3435,In_59,In_804);
nor U3436 (N_3436,In_93,In_251);
xor U3437 (N_3437,In_868,In_544);
and U3438 (N_3438,In_830,In_840);
nor U3439 (N_3439,In_941,In_91);
nor U3440 (N_3440,In_986,In_684);
and U3441 (N_3441,In_229,In_673);
nand U3442 (N_3442,In_804,In_909);
nand U3443 (N_3443,In_859,In_900);
nand U3444 (N_3444,In_14,In_653);
nor U3445 (N_3445,In_265,In_212);
or U3446 (N_3446,In_880,In_123);
or U3447 (N_3447,In_322,In_736);
or U3448 (N_3448,In_493,In_566);
and U3449 (N_3449,In_531,In_574);
and U3450 (N_3450,In_475,In_401);
nor U3451 (N_3451,In_705,In_880);
or U3452 (N_3452,In_352,In_343);
and U3453 (N_3453,In_513,In_857);
and U3454 (N_3454,In_897,In_208);
or U3455 (N_3455,In_105,In_358);
or U3456 (N_3456,In_220,In_192);
and U3457 (N_3457,In_315,In_681);
and U3458 (N_3458,In_258,In_826);
and U3459 (N_3459,In_104,In_642);
or U3460 (N_3460,In_746,In_616);
nand U3461 (N_3461,In_705,In_593);
nor U3462 (N_3462,In_900,In_428);
nand U3463 (N_3463,In_347,In_961);
or U3464 (N_3464,In_168,In_959);
and U3465 (N_3465,In_359,In_723);
or U3466 (N_3466,In_260,In_512);
nand U3467 (N_3467,In_479,In_200);
nand U3468 (N_3468,In_916,In_572);
or U3469 (N_3469,In_247,In_417);
nor U3470 (N_3470,In_787,In_808);
nor U3471 (N_3471,In_766,In_213);
or U3472 (N_3472,In_224,In_914);
or U3473 (N_3473,In_816,In_705);
or U3474 (N_3474,In_528,In_548);
or U3475 (N_3475,In_378,In_84);
or U3476 (N_3476,In_785,In_104);
and U3477 (N_3477,In_385,In_982);
and U3478 (N_3478,In_548,In_551);
or U3479 (N_3479,In_124,In_30);
nand U3480 (N_3480,In_731,In_49);
xor U3481 (N_3481,In_88,In_5);
or U3482 (N_3482,In_741,In_896);
or U3483 (N_3483,In_552,In_59);
and U3484 (N_3484,In_107,In_171);
nor U3485 (N_3485,In_95,In_396);
nor U3486 (N_3486,In_104,In_484);
nor U3487 (N_3487,In_832,In_774);
nor U3488 (N_3488,In_579,In_851);
and U3489 (N_3489,In_967,In_441);
and U3490 (N_3490,In_769,In_957);
nand U3491 (N_3491,In_743,In_484);
nor U3492 (N_3492,In_358,In_137);
nor U3493 (N_3493,In_634,In_328);
nor U3494 (N_3494,In_966,In_365);
nand U3495 (N_3495,In_397,In_922);
or U3496 (N_3496,In_313,In_22);
nand U3497 (N_3497,In_419,In_520);
or U3498 (N_3498,In_497,In_606);
and U3499 (N_3499,In_754,In_106);
or U3500 (N_3500,In_378,In_926);
nor U3501 (N_3501,In_597,In_582);
or U3502 (N_3502,In_778,In_659);
nor U3503 (N_3503,In_62,In_811);
and U3504 (N_3504,In_367,In_374);
nor U3505 (N_3505,In_148,In_222);
xor U3506 (N_3506,In_88,In_250);
xnor U3507 (N_3507,In_803,In_801);
and U3508 (N_3508,In_604,In_958);
nand U3509 (N_3509,In_189,In_428);
or U3510 (N_3510,In_133,In_42);
or U3511 (N_3511,In_826,In_996);
or U3512 (N_3512,In_293,In_123);
or U3513 (N_3513,In_332,In_142);
xor U3514 (N_3514,In_416,In_158);
nand U3515 (N_3515,In_102,In_295);
and U3516 (N_3516,In_127,In_841);
and U3517 (N_3517,In_717,In_585);
and U3518 (N_3518,In_535,In_450);
or U3519 (N_3519,In_679,In_876);
or U3520 (N_3520,In_870,In_499);
or U3521 (N_3521,In_169,In_63);
nor U3522 (N_3522,In_353,In_508);
or U3523 (N_3523,In_545,In_45);
and U3524 (N_3524,In_438,In_217);
nand U3525 (N_3525,In_284,In_921);
nand U3526 (N_3526,In_713,In_833);
nor U3527 (N_3527,In_639,In_977);
nand U3528 (N_3528,In_334,In_671);
and U3529 (N_3529,In_329,In_32);
or U3530 (N_3530,In_784,In_982);
nor U3531 (N_3531,In_610,In_132);
and U3532 (N_3532,In_130,In_165);
nand U3533 (N_3533,In_442,In_646);
xnor U3534 (N_3534,In_212,In_385);
xnor U3535 (N_3535,In_26,In_120);
nor U3536 (N_3536,In_381,In_666);
nand U3537 (N_3537,In_837,In_806);
nor U3538 (N_3538,In_55,In_207);
xor U3539 (N_3539,In_375,In_845);
or U3540 (N_3540,In_735,In_768);
nand U3541 (N_3541,In_284,In_368);
nand U3542 (N_3542,In_202,In_167);
and U3543 (N_3543,In_434,In_815);
nand U3544 (N_3544,In_40,In_601);
nand U3545 (N_3545,In_834,In_109);
or U3546 (N_3546,In_89,In_774);
and U3547 (N_3547,In_22,In_250);
or U3548 (N_3548,In_389,In_751);
nand U3549 (N_3549,In_117,In_596);
xor U3550 (N_3550,In_435,In_24);
and U3551 (N_3551,In_743,In_759);
and U3552 (N_3552,In_513,In_407);
nor U3553 (N_3553,In_331,In_325);
nor U3554 (N_3554,In_964,In_513);
xnor U3555 (N_3555,In_185,In_183);
and U3556 (N_3556,In_73,In_719);
nor U3557 (N_3557,In_32,In_245);
or U3558 (N_3558,In_213,In_949);
and U3559 (N_3559,In_110,In_902);
or U3560 (N_3560,In_45,In_190);
and U3561 (N_3561,In_93,In_82);
nand U3562 (N_3562,In_63,In_305);
nor U3563 (N_3563,In_990,In_278);
or U3564 (N_3564,In_52,In_445);
nor U3565 (N_3565,In_743,In_721);
xor U3566 (N_3566,In_823,In_624);
nand U3567 (N_3567,In_343,In_111);
xor U3568 (N_3568,In_996,In_639);
nor U3569 (N_3569,In_523,In_63);
nand U3570 (N_3570,In_542,In_7);
and U3571 (N_3571,In_870,In_220);
nand U3572 (N_3572,In_414,In_728);
or U3573 (N_3573,In_980,In_945);
and U3574 (N_3574,In_510,In_259);
or U3575 (N_3575,In_828,In_641);
and U3576 (N_3576,In_163,In_519);
nor U3577 (N_3577,In_910,In_765);
nand U3578 (N_3578,In_712,In_797);
or U3579 (N_3579,In_405,In_199);
nor U3580 (N_3580,In_542,In_772);
xnor U3581 (N_3581,In_147,In_903);
and U3582 (N_3582,In_270,In_362);
nor U3583 (N_3583,In_361,In_209);
nor U3584 (N_3584,In_221,In_566);
and U3585 (N_3585,In_24,In_941);
or U3586 (N_3586,In_200,In_120);
and U3587 (N_3587,In_293,In_485);
and U3588 (N_3588,In_315,In_391);
xor U3589 (N_3589,In_4,In_664);
nand U3590 (N_3590,In_865,In_741);
or U3591 (N_3591,In_251,In_47);
and U3592 (N_3592,In_957,In_476);
and U3593 (N_3593,In_194,In_99);
nand U3594 (N_3594,In_737,In_171);
nor U3595 (N_3595,In_939,In_245);
nand U3596 (N_3596,In_12,In_835);
or U3597 (N_3597,In_966,In_460);
and U3598 (N_3598,In_756,In_263);
nor U3599 (N_3599,In_362,In_306);
nand U3600 (N_3600,In_6,In_640);
and U3601 (N_3601,In_233,In_4);
and U3602 (N_3602,In_265,In_827);
nand U3603 (N_3603,In_451,In_325);
or U3604 (N_3604,In_139,In_474);
xnor U3605 (N_3605,In_384,In_790);
nor U3606 (N_3606,In_721,In_206);
or U3607 (N_3607,In_227,In_238);
and U3608 (N_3608,In_738,In_408);
and U3609 (N_3609,In_237,In_769);
nor U3610 (N_3610,In_986,In_910);
or U3611 (N_3611,In_244,In_959);
and U3612 (N_3612,In_832,In_608);
nor U3613 (N_3613,In_514,In_427);
nand U3614 (N_3614,In_253,In_990);
nand U3615 (N_3615,In_352,In_468);
nor U3616 (N_3616,In_736,In_781);
nand U3617 (N_3617,In_30,In_884);
nor U3618 (N_3618,In_40,In_304);
and U3619 (N_3619,In_413,In_273);
nand U3620 (N_3620,In_293,In_933);
nor U3621 (N_3621,In_528,In_642);
nor U3622 (N_3622,In_250,In_875);
and U3623 (N_3623,In_324,In_22);
or U3624 (N_3624,In_254,In_798);
or U3625 (N_3625,In_590,In_599);
nand U3626 (N_3626,In_885,In_433);
and U3627 (N_3627,In_897,In_688);
nor U3628 (N_3628,In_998,In_67);
nand U3629 (N_3629,In_48,In_222);
nor U3630 (N_3630,In_606,In_828);
or U3631 (N_3631,In_858,In_2);
xnor U3632 (N_3632,In_380,In_959);
and U3633 (N_3633,In_347,In_10);
and U3634 (N_3634,In_779,In_384);
or U3635 (N_3635,In_720,In_479);
or U3636 (N_3636,In_298,In_402);
nor U3637 (N_3637,In_277,In_139);
or U3638 (N_3638,In_725,In_52);
nand U3639 (N_3639,In_225,In_236);
nand U3640 (N_3640,In_549,In_76);
nor U3641 (N_3641,In_134,In_777);
and U3642 (N_3642,In_670,In_103);
nand U3643 (N_3643,In_544,In_359);
nand U3644 (N_3644,In_582,In_927);
nand U3645 (N_3645,In_541,In_881);
xor U3646 (N_3646,In_790,In_602);
xnor U3647 (N_3647,In_10,In_309);
and U3648 (N_3648,In_193,In_1);
and U3649 (N_3649,In_405,In_12);
or U3650 (N_3650,In_706,In_559);
and U3651 (N_3651,In_880,In_641);
nand U3652 (N_3652,In_600,In_344);
and U3653 (N_3653,In_770,In_308);
nor U3654 (N_3654,In_808,In_427);
and U3655 (N_3655,In_252,In_184);
and U3656 (N_3656,In_469,In_356);
nand U3657 (N_3657,In_704,In_303);
and U3658 (N_3658,In_743,In_648);
or U3659 (N_3659,In_272,In_106);
and U3660 (N_3660,In_237,In_26);
or U3661 (N_3661,In_907,In_150);
nor U3662 (N_3662,In_350,In_840);
nand U3663 (N_3663,In_119,In_135);
nand U3664 (N_3664,In_393,In_414);
nand U3665 (N_3665,In_564,In_270);
nand U3666 (N_3666,In_139,In_831);
or U3667 (N_3667,In_524,In_81);
and U3668 (N_3668,In_713,In_297);
nand U3669 (N_3669,In_362,In_128);
nor U3670 (N_3670,In_788,In_920);
or U3671 (N_3671,In_718,In_685);
nor U3672 (N_3672,In_104,In_366);
nand U3673 (N_3673,In_374,In_164);
or U3674 (N_3674,In_759,In_30);
xnor U3675 (N_3675,In_76,In_134);
nor U3676 (N_3676,In_429,In_960);
xnor U3677 (N_3677,In_537,In_63);
and U3678 (N_3678,In_173,In_858);
nor U3679 (N_3679,In_362,In_352);
nor U3680 (N_3680,In_263,In_45);
and U3681 (N_3681,In_825,In_529);
or U3682 (N_3682,In_422,In_460);
and U3683 (N_3683,In_295,In_597);
or U3684 (N_3684,In_705,In_449);
or U3685 (N_3685,In_111,In_435);
and U3686 (N_3686,In_606,In_988);
nand U3687 (N_3687,In_982,In_999);
xor U3688 (N_3688,In_338,In_189);
nand U3689 (N_3689,In_514,In_190);
nand U3690 (N_3690,In_966,In_670);
nor U3691 (N_3691,In_169,In_882);
or U3692 (N_3692,In_981,In_928);
nor U3693 (N_3693,In_200,In_715);
nand U3694 (N_3694,In_322,In_812);
xor U3695 (N_3695,In_211,In_872);
or U3696 (N_3696,In_419,In_628);
and U3697 (N_3697,In_241,In_771);
or U3698 (N_3698,In_814,In_990);
nor U3699 (N_3699,In_509,In_483);
nor U3700 (N_3700,In_287,In_674);
xor U3701 (N_3701,In_430,In_499);
or U3702 (N_3702,In_426,In_466);
and U3703 (N_3703,In_134,In_556);
nor U3704 (N_3704,In_565,In_979);
nor U3705 (N_3705,In_222,In_268);
nor U3706 (N_3706,In_89,In_343);
and U3707 (N_3707,In_279,In_907);
xnor U3708 (N_3708,In_614,In_920);
nor U3709 (N_3709,In_205,In_299);
and U3710 (N_3710,In_256,In_934);
and U3711 (N_3711,In_362,In_815);
xor U3712 (N_3712,In_226,In_238);
and U3713 (N_3713,In_695,In_494);
or U3714 (N_3714,In_331,In_291);
and U3715 (N_3715,In_313,In_867);
and U3716 (N_3716,In_335,In_330);
nor U3717 (N_3717,In_447,In_95);
or U3718 (N_3718,In_22,In_183);
or U3719 (N_3719,In_259,In_261);
or U3720 (N_3720,In_374,In_992);
and U3721 (N_3721,In_310,In_152);
and U3722 (N_3722,In_853,In_517);
nand U3723 (N_3723,In_750,In_687);
xor U3724 (N_3724,In_105,In_700);
nand U3725 (N_3725,In_184,In_474);
and U3726 (N_3726,In_983,In_371);
xnor U3727 (N_3727,In_156,In_167);
and U3728 (N_3728,In_668,In_333);
and U3729 (N_3729,In_107,In_768);
and U3730 (N_3730,In_630,In_339);
nor U3731 (N_3731,In_9,In_787);
and U3732 (N_3732,In_540,In_650);
or U3733 (N_3733,In_253,In_532);
nor U3734 (N_3734,In_258,In_437);
nand U3735 (N_3735,In_483,In_553);
and U3736 (N_3736,In_436,In_977);
nor U3737 (N_3737,In_102,In_955);
or U3738 (N_3738,In_820,In_775);
nand U3739 (N_3739,In_317,In_304);
or U3740 (N_3740,In_217,In_617);
nand U3741 (N_3741,In_772,In_774);
nor U3742 (N_3742,In_395,In_780);
xnor U3743 (N_3743,In_441,In_97);
or U3744 (N_3744,In_971,In_817);
and U3745 (N_3745,In_297,In_746);
or U3746 (N_3746,In_393,In_296);
nor U3747 (N_3747,In_935,In_510);
and U3748 (N_3748,In_974,In_451);
or U3749 (N_3749,In_817,In_680);
xor U3750 (N_3750,In_971,In_614);
nor U3751 (N_3751,In_673,In_16);
nor U3752 (N_3752,In_888,In_622);
nand U3753 (N_3753,In_954,In_621);
nand U3754 (N_3754,In_263,In_948);
and U3755 (N_3755,In_242,In_885);
and U3756 (N_3756,In_906,In_150);
nand U3757 (N_3757,In_724,In_330);
nor U3758 (N_3758,In_276,In_978);
or U3759 (N_3759,In_317,In_438);
nand U3760 (N_3760,In_417,In_667);
nand U3761 (N_3761,In_329,In_858);
nor U3762 (N_3762,In_325,In_179);
or U3763 (N_3763,In_37,In_682);
nor U3764 (N_3764,In_259,In_705);
nand U3765 (N_3765,In_237,In_471);
nand U3766 (N_3766,In_653,In_954);
and U3767 (N_3767,In_300,In_134);
or U3768 (N_3768,In_711,In_805);
or U3769 (N_3769,In_409,In_62);
nand U3770 (N_3770,In_773,In_809);
nand U3771 (N_3771,In_551,In_136);
nand U3772 (N_3772,In_925,In_258);
and U3773 (N_3773,In_985,In_599);
nor U3774 (N_3774,In_254,In_813);
xor U3775 (N_3775,In_444,In_967);
nand U3776 (N_3776,In_695,In_48);
nand U3777 (N_3777,In_967,In_52);
or U3778 (N_3778,In_261,In_148);
nand U3779 (N_3779,In_723,In_250);
nor U3780 (N_3780,In_441,In_455);
nand U3781 (N_3781,In_192,In_22);
xor U3782 (N_3782,In_930,In_846);
and U3783 (N_3783,In_622,In_265);
or U3784 (N_3784,In_936,In_521);
nand U3785 (N_3785,In_302,In_698);
nor U3786 (N_3786,In_746,In_919);
xnor U3787 (N_3787,In_836,In_1);
xor U3788 (N_3788,In_62,In_713);
nor U3789 (N_3789,In_194,In_544);
or U3790 (N_3790,In_855,In_705);
xor U3791 (N_3791,In_516,In_577);
or U3792 (N_3792,In_129,In_102);
nand U3793 (N_3793,In_542,In_685);
or U3794 (N_3794,In_623,In_665);
or U3795 (N_3795,In_19,In_862);
and U3796 (N_3796,In_742,In_388);
nor U3797 (N_3797,In_124,In_626);
and U3798 (N_3798,In_326,In_813);
nor U3799 (N_3799,In_53,In_505);
or U3800 (N_3800,In_198,In_763);
nand U3801 (N_3801,In_597,In_447);
or U3802 (N_3802,In_888,In_367);
nand U3803 (N_3803,In_755,In_951);
or U3804 (N_3804,In_440,In_134);
nand U3805 (N_3805,In_44,In_945);
nand U3806 (N_3806,In_470,In_149);
or U3807 (N_3807,In_799,In_644);
nand U3808 (N_3808,In_135,In_292);
nand U3809 (N_3809,In_487,In_383);
nand U3810 (N_3810,In_771,In_701);
and U3811 (N_3811,In_577,In_711);
nor U3812 (N_3812,In_390,In_156);
nor U3813 (N_3813,In_821,In_804);
or U3814 (N_3814,In_414,In_383);
xnor U3815 (N_3815,In_93,In_660);
or U3816 (N_3816,In_768,In_905);
or U3817 (N_3817,In_31,In_807);
and U3818 (N_3818,In_933,In_71);
and U3819 (N_3819,In_184,In_701);
or U3820 (N_3820,In_500,In_522);
or U3821 (N_3821,In_571,In_196);
or U3822 (N_3822,In_300,In_172);
nand U3823 (N_3823,In_764,In_913);
and U3824 (N_3824,In_450,In_58);
nand U3825 (N_3825,In_786,In_125);
and U3826 (N_3826,In_56,In_690);
nor U3827 (N_3827,In_574,In_5);
and U3828 (N_3828,In_272,In_567);
and U3829 (N_3829,In_750,In_379);
nor U3830 (N_3830,In_537,In_477);
or U3831 (N_3831,In_558,In_727);
nand U3832 (N_3832,In_347,In_874);
nand U3833 (N_3833,In_797,In_577);
xor U3834 (N_3834,In_976,In_265);
nor U3835 (N_3835,In_2,In_366);
or U3836 (N_3836,In_586,In_243);
or U3837 (N_3837,In_417,In_962);
and U3838 (N_3838,In_642,In_308);
and U3839 (N_3839,In_351,In_414);
and U3840 (N_3840,In_888,In_66);
nor U3841 (N_3841,In_810,In_666);
nand U3842 (N_3842,In_465,In_642);
nand U3843 (N_3843,In_19,In_106);
nand U3844 (N_3844,In_13,In_971);
or U3845 (N_3845,In_905,In_929);
or U3846 (N_3846,In_775,In_891);
nor U3847 (N_3847,In_75,In_534);
or U3848 (N_3848,In_440,In_409);
or U3849 (N_3849,In_992,In_48);
or U3850 (N_3850,In_410,In_894);
xnor U3851 (N_3851,In_85,In_908);
and U3852 (N_3852,In_313,In_773);
and U3853 (N_3853,In_69,In_759);
nor U3854 (N_3854,In_996,In_119);
nor U3855 (N_3855,In_101,In_160);
nor U3856 (N_3856,In_308,In_141);
nor U3857 (N_3857,In_54,In_52);
nand U3858 (N_3858,In_742,In_823);
or U3859 (N_3859,In_421,In_689);
nor U3860 (N_3860,In_260,In_62);
and U3861 (N_3861,In_906,In_620);
and U3862 (N_3862,In_970,In_974);
nor U3863 (N_3863,In_816,In_552);
or U3864 (N_3864,In_725,In_920);
and U3865 (N_3865,In_815,In_955);
nand U3866 (N_3866,In_115,In_439);
or U3867 (N_3867,In_692,In_679);
nand U3868 (N_3868,In_237,In_504);
nand U3869 (N_3869,In_147,In_308);
nor U3870 (N_3870,In_598,In_756);
or U3871 (N_3871,In_770,In_12);
and U3872 (N_3872,In_933,In_655);
nand U3873 (N_3873,In_331,In_381);
or U3874 (N_3874,In_762,In_764);
and U3875 (N_3875,In_283,In_188);
nor U3876 (N_3876,In_753,In_656);
or U3877 (N_3877,In_417,In_801);
and U3878 (N_3878,In_204,In_769);
nand U3879 (N_3879,In_374,In_98);
and U3880 (N_3880,In_730,In_921);
xnor U3881 (N_3881,In_199,In_442);
nor U3882 (N_3882,In_304,In_422);
and U3883 (N_3883,In_293,In_285);
nor U3884 (N_3884,In_861,In_142);
nor U3885 (N_3885,In_263,In_156);
nor U3886 (N_3886,In_40,In_715);
nor U3887 (N_3887,In_759,In_560);
or U3888 (N_3888,In_663,In_534);
and U3889 (N_3889,In_496,In_779);
nand U3890 (N_3890,In_478,In_767);
nand U3891 (N_3891,In_217,In_856);
nor U3892 (N_3892,In_735,In_783);
and U3893 (N_3893,In_447,In_853);
xnor U3894 (N_3894,In_903,In_385);
nor U3895 (N_3895,In_717,In_736);
and U3896 (N_3896,In_995,In_513);
and U3897 (N_3897,In_243,In_128);
or U3898 (N_3898,In_490,In_229);
and U3899 (N_3899,In_938,In_852);
or U3900 (N_3900,In_618,In_152);
or U3901 (N_3901,In_434,In_705);
nand U3902 (N_3902,In_466,In_785);
or U3903 (N_3903,In_384,In_294);
nand U3904 (N_3904,In_927,In_484);
and U3905 (N_3905,In_295,In_705);
xor U3906 (N_3906,In_820,In_869);
nor U3907 (N_3907,In_631,In_397);
nand U3908 (N_3908,In_927,In_432);
and U3909 (N_3909,In_154,In_500);
or U3910 (N_3910,In_512,In_419);
or U3911 (N_3911,In_934,In_885);
and U3912 (N_3912,In_834,In_778);
or U3913 (N_3913,In_232,In_124);
nand U3914 (N_3914,In_892,In_946);
nor U3915 (N_3915,In_200,In_634);
nand U3916 (N_3916,In_720,In_651);
nand U3917 (N_3917,In_806,In_758);
or U3918 (N_3918,In_316,In_357);
xor U3919 (N_3919,In_809,In_285);
xor U3920 (N_3920,In_319,In_948);
and U3921 (N_3921,In_842,In_412);
or U3922 (N_3922,In_200,In_908);
nor U3923 (N_3923,In_749,In_479);
or U3924 (N_3924,In_564,In_397);
nand U3925 (N_3925,In_961,In_397);
and U3926 (N_3926,In_26,In_245);
and U3927 (N_3927,In_721,In_732);
or U3928 (N_3928,In_485,In_260);
nor U3929 (N_3929,In_746,In_618);
nand U3930 (N_3930,In_447,In_847);
or U3931 (N_3931,In_231,In_340);
or U3932 (N_3932,In_874,In_27);
nand U3933 (N_3933,In_446,In_839);
xor U3934 (N_3934,In_686,In_867);
nand U3935 (N_3935,In_206,In_964);
xor U3936 (N_3936,In_54,In_183);
nand U3937 (N_3937,In_369,In_806);
or U3938 (N_3938,In_746,In_918);
or U3939 (N_3939,In_605,In_659);
nand U3940 (N_3940,In_71,In_246);
xor U3941 (N_3941,In_749,In_813);
and U3942 (N_3942,In_704,In_382);
nor U3943 (N_3943,In_621,In_52);
and U3944 (N_3944,In_541,In_978);
nand U3945 (N_3945,In_771,In_343);
nor U3946 (N_3946,In_162,In_562);
or U3947 (N_3947,In_847,In_570);
nor U3948 (N_3948,In_156,In_767);
xor U3949 (N_3949,In_922,In_396);
nor U3950 (N_3950,In_381,In_281);
and U3951 (N_3951,In_64,In_950);
nand U3952 (N_3952,In_327,In_832);
or U3953 (N_3953,In_897,In_886);
nand U3954 (N_3954,In_11,In_846);
and U3955 (N_3955,In_428,In_582);
or U3956 (N_3956,In_250,In_816);
and U3957 (N_3957,In_138,In_721);
nand U3958 (N_3958,In_752,In_497);
nand U3959 (N_3959,In_890,In_635);
and U3960 (N_3960,In_72,In_234);
nor U3961 (N_3961,In_782,In_142);
and U3962 (N_3962,In_473,In_974);
nor U3963 (N_3963,In_490,In_222);
nor U3964 (N_3964,In_836,In_671);
nor U3965 (N_3965,In_398,In_962);
and U3966 (N_3966,In_340,In_249);
and U3967 (N_3967,In_417,In_85);
and U3968 (N_3968,In_25,In_969);
and U3969 (N_3969,In_618,In_406);
nand U3970 (N_3970,In_439,In_316);
and U3971 (N_3971,In_813,In_446);
nand U3972 (N_3972,In_331,In_420);
and U3973 (N_3973,In_210,In_123);
and U3974 (N_3974,In_405,In_891);
or U3975 (N_3975,In_988,In_46);
xnor U3976 (N_3976,In_771,In_420);
and U3977 (N_3977,In_449,In_53);
and U3978 (N_3978,In_568,In_496);
nand U3979 (N_3979,In_872,In_160);
nand U3980 (N_3980,In_973,In_354);
nand U3981 (N_3981,In_809,In_92);
nand U3982 (N_3982,In_111,In_219);
or U3983 (N_3983,In_563,In_100);
or U3984 (N_3984,In_270,In_931);
and U3985 (N_3985,In_9,In_91);
and U3986 (N_3986,In_609,In_336);
nand U3987 (N_3987,In_83,In_318);
nand U3988 (N_3988,In_16,In_149);
xor U3989 (N_3989,In_555,In_358);
nand U3990 (N_3990,In_443,In_700);
nor U3991 (N_3991,In_292,In_583);
or U3992 (N_3992,In_590,In_987);
or U3993 (N_3993,In_336,In_240);
and U3994 (N_3994,In_910,In_532);
nor U3995 (N_3995,In_404,In_511);
or U3996 (N_3996,In_995,In_181);
xnor U3997 (N_3997,In_53,In_626);
or U3998 (N_3998,In_198,In_122);
and U3999 (N_3999,In_415,In_884);
nand U4000 (N_4000,In_84,In_15);
nor U4001 (N_4001,In_69,In_343);
or U4002 (N_4002,In_267,In_354);
and U4003 (N_4003,In_564,In_323);
and U4004 (N_4004,In_136,In_292);
nor U4005 (N_4005,In_739,In_741);
and U4006 (N_4006,In_597,In_419);
nand U4007 (N_4007,In_936,In_153);
or U4008 (N_4008,In_312,In_757);
or U4009 (N_4009,In_606,In_374);
or U4010 (N_4010,In_331,In_954);
nor U4011 (N_4011,In_329,In_548);
nand U4012 (N_4012,In_710,In_813);
nor U4013 (N_4013,In_952,In_141);
nor U4014 (N_4014,In_139,In_664);
or U4015 (N_4015,In_653,In_988);
and U4016 (N_4016,In_525,In_692);
nor U4017 (N_4017,In_165,In_146);
or U4018 (N_4018,In_20,In_906);
nor U4019 (N_4019,In_443,In_419);
and U4020 (N_4020,In_915,In_497);
nand U4021 (N_4021,In_172,In_883);
xnor U4022 (N_4022,In_745,In_254);
nor U4023 (N_4023,In_12,In_428);
nor U4024 (N_4024,In_140,In_232);
and U4025 (N_4025,In_213,In_333);
or U4026 (N_4026,In_374,In_233);
or U4027 (N_4027,In_39,In_372);
and U4028 (N_4028,In_222,In_168);
or U4029 (N_4029,In_136,In_716);
or U4030 (N_4030,In_833,In_544);
and U4031 (N_4031,In_325,In_439);
nand U4032 (N_4032,In_690,In_412);
or U4033 (N_4033,In_742,In_499);
and U4034 (N_4034,In_396,In_74);
nand U4035 (N_4035,In_464,In_707);
nand U4036 (N_4036,In_530,In_785);
and U4037 (N_4037,In_585,In_316);
nor U4038 (N_4038,In_241,In_937);
nand U4039 (N_4039,In_575,In_377);
and U4040 (N_4040,In_95,In_555);
and U4041 (N_4041,In_307,In_921);
nor U4042 (N_4042,In_230,In_263);
or U4043 (N_4043,In_472,In_433);
nor U4044 (N_4044,In_993,In_336);
and U4045 (N_4045,In_203,In_895);
nand U4046 (N_4046,In_395,In_872);
and U4047 (N_4047,In_26,In_514);
nor U4048 (N_4048,In_623,In_723);
nor U4049 (N_4049,In_258,In_399);
xor U4050 (N_4050,In_118,In_399);
or U4051 (N_4051,In_927,In_747);
nor U4052 (N_4052,In_694,In_428);
and U4053 (N_4053,In_482,In_587);
and U4054 (N_4054,In_57,In_36);
nand U4055 (N_4055,In_759,In_442);
xnor U4056 (N_4056,In_521,In_626);
nand U4057 (N_4057,In_495,In_283);
and U4058 (N_4058,In_138,In_359);
and U4059 (N_4059,In_418,In_622);
nor U4060 (N_4060,In_941,In_983);
nand U4061 (N_4061,In_745,In_389);
nand U4062 (N_4062,In_268,In_484);
xor U4063 (N_4063,In_180,In_335);
nor U4064 (N_4064,In_345,In_709);
and U4065 (N_4065,In_315,In_544);
nor U4066 (N_4066,In_221,In_260);
nor U4067 (N_4067,In_274,In_840);
nor U4068 (N_4068,In_758,In_311);
and U4069 (N_4069,In_31,In_604);
or U4070 (N_4070,In_69,In_348);
nand U4071 (N_4071,In_697,In_36);
or U4072 (N_4072,In_235,In_360);
xor U4073 (N_4073,In_752,In_233);
nand U4074 (N_4074,In_684,In_619);
nor U4075 (N_4075,In_635,In_23);
nor U4076 (N_4076,In_658,In_296);
and U4077 (N_4077,In_98,In_669);
and U4078 (N_4078,In_542,In_624);
and U4079 (N_4079,In_323,In_734);
or U4080 (N_4080,In_646,In_699);
and U4081 (N_4081,In_828,In_527);
and U4082 (N_4082,In_532,In_338);
nor U4083 (N_4083,In_865,In_364);
nand U4084 (N_4084,In_6,In_299);
and U4085 (N_4085,In_964,In_786);
nor U4086 (N_4086,In_879,In_944);
and U4087 (N_4087,In_78,In_44);
and U4088 (N_4088,In_443,In_679);
and U4089 (N_4089,In_219,In_237);
and U4090 (N_4090,In_525,In_602);
xnor U4091 (N_4091,In_797,In_368);
or U4092 (N_4092,In_131,In_307);
or U4093 (N_4093,In_300,In_88);
and U4094 (N_4094,In_324,In_172);
nor U4095 (N_4095,In_358,In_525);
nand U4096 (N_4096,In_1,In_852);
nand U4097 (N_4097,In_135,In_846);
xnor U4098 (N_4098,In_815,In_982);
and U4099 (N_4099,In_314,In_870);
or U4100 (N_4100,In_792,In_444);
xnor U4101 (N_4101,In_932,In_865);
or U4102 (N_4102,In_502,In_835);
nor U4103 (N_4103,In_898,In_425);
and U4104 (N_4104,In_322,In_452);
nor U4105 (N_4105,In_877,In_756);
nor U4106 (N_4106,In_918,In_457);
or U4107 (N_4107,In_276,In_103);
or U4108 (N_4108,In_720,In_517);
or U4109 (N_4109,In_132,In_394);
nand U4110 (N_4110,In_684,In_323);
nand U4111 (N_4111,In_397,In_301);
nor U4112 (N_4112,In_848,In_518);
nor U4113 (N_4113,In_210,In_399);
nor U4114 (N_4114,In_929,In_91);
or U4115 (N_4115,In_21,In_59);
or U4116 (N_4116,In_670,In_199);
xnor U4117 (N_4117,In_694,In_832);
xor U4118 (N_4118,In_682,In_735);
xnor U4119 (N_4119,In_782,In_114);
and U4120 (N_4120,In_908,In_892);
nor U4121 (N_4121,In_66,In_971);
or U4122 (N_4122,In_214,In_147);
nand U4123 (N_4123,In_715,In_435);
nand U4124 (N_4124,In_911,In_837);
xor U4125 (N_4125,In_277,In_427);
and U4126 (N_4126,In_917,In_725);
xnor U4127 (N_4127,In_788,In_677);
or U4128 (N_4128,In_578,In_989);
and U4129 (N_4129,In_467,In_455);
nor U4130 (N_4130,In_324,In_801);
or U4131 (N_4131,In_495,In_682);
xnor U4132 (N_4132,In_239,In_737);
or U4133 (N_4133,In_365,In_497);
nand U4134 (N_4134,In_664,In_873);
nand U4135 (N_4135,In_279,In_716);
or U4136 (N_4136,In_65,In_421);
and U4137 (N_4137,In_576,In_341);
and U4138 (N_4138,In_958,In_574);
or U4139 (N_4139,In_853,In_428);
or U4140 (N_4140,In_617,In_695);
or U4141 (N_4141,In_476,In_781);
or U4142 (N_4142,In_832,In_333);
and U4143 (N_4143,In_839,In_896);
nor U4144 (N_4144,In_273,In_691);
nor U4145 (N_4145,In_374,In_368);
nand U4146 (N_4146,In_427,In_864);
or U4147 (N_4147,In_169,In_509);
xnor U4148 (N_4148,In_64,In_110);
nand U4149 (N_4149,In_636,In_719);
nor U4150 (N_4150,In_461,In_297);
nand U4151 (N_4151,In_601,In_636);
or U4152 (N_4152,In_435,In_388);
and U4153 (N_4153,In_933,In_333);
and U4154 (N_4154,In_85,In_88);
or U4155 (N_4155,In_489,In_268);
xor U4156 (N_4156,In_744,In_388);
nand U4157 (N_4157,In_146,In_414);
nor U4158 (N_4158,In_583,In_507);
and U4159 (N_4159,In_276,In_938);
nor U4160 (N_4160,In_60,In_185);
nand U4161 (N_4161,In_573,In_642);
and U4162 (N_4162,In_949,In_498);
nand U4163 (N_4163,In_366,In_854);
or U4164 (N_4164,In_814,In_129);
nand U4165 (N_4165,In_414,In_853);
or U4166 (N_4166,In_526,In_937);
or U4167 (N_4167,In_749,In_392);
nor U4168 (N_4168,In_893,In_795);
and U4169 (N_4169,In_82,In_77);
and U4170 (N_4170,In_636,In_98);
nor U4171 (N_4171,In_365,In_737);
or U4172 (N_4172,In_57,In_159);
xor U4173 (N_4173,In_706,In_315);
nand U4174 (N_4174,In_141,In_929);
nand U4175 (N_4175,In_360,In_342);
nand U4176 (N_4176,In_13,In_502);
and U4177 (N_4177,In_249,In_737);
nor U4178 (N_4178,In_549,In_277);
and U4179 (N_4179,In_854,In_749);
nand U4180 (N_4180,In_391,In_340);
nand U4181 (N_4181,In_687,In_573);
nor U4182 (N_4182,In_575,In_132);
nand U4183 (N_4183,In_48,In_828);
or U4184 (N_4184,In_128,In_78);
and U4185 (N_4185,In_678,In_600);
or U4186 (N_4186,In_772,In_398);
nand U4187 (N_4187,In_183,In_539);
and U4188 (N_4188,In_747,In_474);
or U4189 (N_4189,In_417,In_683);
nor U4190 (N_4190,In_163,In_829);
and U4191 (N_4191,In_780,In_187);
or U4192 (N_4192,In_44,In_851);
nor U4193 (N_4193,In_496,In_208);
and U4194 (N_4194,In_818,In_585);
xor U4195 (N_4195,In_928,In_188);
or U4196 (N_4196,In_539,In_270);
or U4197 (N_4197,In_646,In_422);
nand U4198 (N_4198,In_738,In_205);
or U4199 (N_4199,In_342,In_99);
nor U4200 (N_4200,In_453,In_167);
and U4201 (N_4201,In_229,In_524);
nand U4202 (N_4202,In_225,In_263);
or U4203 (N_4203,In_819,In_990);
nand U4204 (N_4204,In_231,In_541);
nor U4205 (N_4205,In_46,In_796);
or U4206 (N_4206,In_217,In_638);
and U4207 (N_4207,In_188,In_752);
or U4208 (N_4208,In_434,In_575);
nand U4209 (N_4209,In_842,In_1);
xor U4210 (N_4210,In_996,In_492);
and U4211 (N_4211,In_203,In_446);
xor U4212 (N_4212,In_727,In_504);
nand U4213 (N_4213,In_146,In_584);
or U4214 (N_4214,In_238,In_338);
and U4215 (N_4215,In_807,In_765);
nor U4216 (N_4216,In_742,In_588);
or U4217 (N_4217,In_512,In_216);
and U4218 (N_4218,In_325,In_89);
or U4219 (N_4219,In_128,In_24);
and U4220 (N_4220,In_322,In_354);
and U4221 (N_4221,In_767,In_665);
nand U4222 (N_4222,In_133,In_276);
or U4223 (N_4223,In_954,In_980);
xnor U4224 (N_4224,In_257,In_198);
and U4225 (N_4225,In_901,In_235);
nand U4226 (N_4226,In_896,In_291);
nor U4227 (N_4227,In_276,In_660);
xor U4228 (N_4228,In_247,In_564);
nand U4229 (N_4229,In_569,In_21);
nor U4230 (N_4230,In_918,In_233);
nand U4231 (N_4231,In_216,In_50);
nand U4232 (N_4232,In_301,In_262);
or U4233 (N_4233,In_710,In_816);
and U4234 (N_4234,In_845,In_184);
nand U4235 (N_4235,In_101,In_566);
or U4236 (N_4236,In_231,In_247);
or U4237 (N_4237,In_302,In_100);
and U4238 (N_4238,In_930,In_424);
nand U4239 (N_4239,In_527,In_18);
and U4240 (N_4240,In_609,In_988);
nand U4241 (N_4241,In_266,In_566);
and U4242 (N_4242,In_550,In_961);
nand U4243 (N_4243,In_426,In_497);
and U4244 (N_4244,In_713,In_16);
and U4245 (N_4245,In_32,In_141);
or U4246 (N_4246,In_547,In_964);
or U4247 (N_4247,In_782,In_44);
and U4248 (N_4248,In_310,In_251);
and U4249 (N_4249,In_185,In_195);
nand U4250 (N_4250,In_919,In_782);
and U4251 (N_4251,In_280,In_634);
nor U4252 (N_4252,In_648,In_445);
nand U4253 (N_4253,In_865,In_218);
nor U4254 (N_4254,In_727,In_480);
nand U4255 (N_4255,In_81,In_853);
and U4256 (N_4256,In_720,In_403);
and U4257 (N_4257,In_309,In_239);
xor U4258 (N_4258,In_996,In_638);
xor U4259 (N_4259,In_570,In_509);
xor U4260 (N_4260,In_604,In_863);
or U4261 (N_4261,In_110,In_304);
nor U4262 (N_4262,In_568,In_691);
nand U4263 (N_4263,In_521,In_9);
nor U4264 (N_4264,In_494,In_70);
and U4265 (N_4265,In_966,In_556);
and U4266 (N_4266,In_849,In_642);
and U4267 (N_4267,In_568,In_6);
or U4268 (N_4268,In_404,In_281);
nand U4269 (N_4269,In_360,In_499);
nor U4270 (N_4270,In_826,In_904);
xor U4271 (N_4271,In_991,In_499);
or U4272 (N_4272,In_520,In_919);
nand U4273 (N_4273,In_41,In_723);
and U4274 (N_4274,In_566,In_808);
or U4275 (N_4275,In_117,In_300);
nand U4276 (N_4276,In_856,In_157);
nor U4277 (N_4277,In_441,In_678);
and U4278 (N_4278,In_83,In_297);
xnor U4279 (N_4279,In_256,In_825);
nand U4280 (N_4280,In_256,In_249);
nor U4281 (N_4281,In_4,In_183);
and U4282 (N_4282,In_811,In_128);
nor U4283 (N_4283,In_576,In_816);
nand U4284 (N_4284,In_807,In_826);
nand U4285 (N_4285,In_431,In_849);
nor U4286 (N_4286,In_337,In_702);
nand U4287 (N_4287,In_259,In_646);
or U4288 (N_4288,In_370,In_884);
nor U4289 (N_4289,In_347,In_378);
or U4290 (N_4290,In_794,In_145);
and U4291 (N_4291,In_994,In_127);
or U4292 (N_4292,In_217,In_754);
nor U4293 (N_4293,In_630,In_775);
or U4294 (N_4294,In_834,In_575);
and U4295 (N_4295,In_603,In_858);
nor U4296 (N_4296,In_911,In_337);
and U4297 (N_4297,In_170,In_641);
nor U4298 (N_4298,In_631,In_25);
nand U4299 (N_4299,In_574,In_104);
nand U4300 (N_4300,In_352,In_146);
nor U4301 (N_4301,In_689,In_481);
nand U4302 (N_4302,In_741,In_382);
xnor U4303 (N_4303,In_772,In_494);
xor U4304 (N_4304,In_570,In_514);
nand U4305 (N_4305,In_455,In_461);
nor U4306 (N_4306,In_204,In_852);
nor U4307 (N_4307,In_256,In_707);
nand U4308 (N_4308,In_571,In_264);
or U4309 (N_4309,In_901,In_949);
and U4310 (N_4310,In_850,In_424);
xor U4311 (N_4311,In_373,In_488);
nor U4312 (N_4312,In_48,In_340);
and U4313 (N_4313,In_774,In_207);
or U4314 (N_4314,In_987,In_450);
and U4315 (N_4315,In_900,In_5);
nor U4316 (N_4316,In_50,In_871);
nor U4317 (N_4317,In_665,In_460);
or U4318 (N_4318,In_869,In_74);
and U4319 (N_4319,In_760,In_387);
nand U4320 (N_4320,In_5,In_256);
or U4321 (N_4321,In_716,In_634);
or U4322 (N_4322,In_408,In_102);
and U4323 (N_4323,In_745,In_637);
nor U4324 (N_4324,In_474,In_965);
or U4325 (N_4325,In_499,In_726);
or U4326 (N_4326,In_985,In_66);
or U4327 (N_4327,In_336,In_735);
nand U4328 (N_4328,In_724,In_645);
or U4329 (N_4329,In_159,In_580);
or U4330 (N_4330,In_888,In_143);
nor U4331 (N_4331,In_608,In_629);
and U4332 (N_4332,In_965,In_219);
nand U4333 (N_4333,In_5,In_736);
and U4334 (N_4334,In_275,In_122);
nor U4335 (N_4335,In_921,In_219);
or U4336 (N_4336,In_214,In_915);
or U4337 (N_4337,In_893,In_426);
or U4338 (N_4338,In_490,In_333);
and U4339 (N_4339,In_859,In_307);
nor U4340 (N_4340,In_700,In_368);
and U4341 (N_4341,In_68,In_799);
nor U4342 (N_4342,In_36,In_726);
or U4343 (N_4343,In_615,In_676);
nand U4344 (N_4344,In_502,In_116);
nand U4345 (N_4345,In_636,In_630);
or U4346 (N_4346,In_310,In_314);
nand U4347 (N_4347,In_183,In_793);
nand U4348 (N_4348,In_460,In_59);
nand U4349 (N_4349,In_409,In_81);
and U4350 (N_4350,In_223,In_301);
xor U4351 (N_4351,In_744,In_265);
or U4352 (N_4352,In_485,In_382);
nor U4353 (N_4353,In_237,In_88);
or U4354 (N_4354,In_621,In_852);
or U4355 (N_4355,In_542,In_491);
nand U4356 (N_4356,In_221,In_243);
and U4357 (N_4357,In_910,In_942);
and U4358 (N_4358,In_151,In_349);
nor U4359 (N_4359,In_824,In_98);
or U4360 (N_4360,In_741,In_137);
nor U4361 (N_4361,In_933,In_902);
or U4362 (N_4362,In_982,In_780);
xnor U4363 (N_4363,In_597,In_130);
and U4364 (N_4364,In_680,In_810);
or U4365 (N_4365,In_897,In_592);
and U4366 (N_4366,In_524,In_843);
or U4367 (N_4367,In_616,In_465);
nor U4368 (N_4368,In_331,In_283);
or U4369 (N_4369,In_456,In_667);
nand U4370 (N_4370,In_467,In_593);
xnor U4371 (N_4371,In_688,In_75);
nor U4372 (N_4372,In_769,In_0);
or U4373 (N_4373,In_247,In_175);
and U4374 (N_4374,In_369,In_951);
nand U4375 (N_4375,In_346,In_772);
nor U4376 (N_4376,In_231,In_992);
and U4377 (N_4377,In_928,In_810);
or U4378 (N_4378,In_457,In_566);
or U4379 (N_4379,In_847,In_505);
nor U4380 (N_4380,In_360,In_496);
nand U4381 (N_4381,In_774,In_229);
nor U4382 (N_4382,In_618,In_554);
or U4383 (N_4383,In_260,In_679);
nor U4384 (N_4384,In_407,In_877);
nor U4385 (N_4385,In_915,In_922);
and U4386 (N_4386,In_8,In_675);
nor U4387 (N_4387,In_968,In_750);
or U4388 (N_4388,In_691,In_465);
nand U4389 (N_4389,In_679,In_907);
nand U4390 (N_4390,In_742,In_147);
nand U4391 (N_4391,In_312,In_728);
or U4392 (N_4392,In_667,In_755);
or U4393 (N_4393,In_229,In_877);
or U4394 (N_4394,In_741,In_809);
or U4395 (N_4395,In_437,In_301);
and U4396 (N_4396,In_488,In_646);
and U4397 (N_4397,In_261,In_298);
xor U4398 (N_4398,In_511,In_421);
or U4399 (N_4399,In_387,In_78);
nand U4400 (N_4400,In_591,In_562);
nand U4401 (N_4401,In_934,In_953);
or U4402 (N_4402,In_484,In_173);
or U4403 (N_4403,In_242,In_899);
or U4404 (N_4404,In_881,In_441);
or U4405 (N_4405,In_187,In_478);
xnor U4406 (N_4406,In_365,In_31);
or U4407 (N_4407,In_501,In_588);
and U4408 (N_4408,In_911,In_474);
nor U4409 (N_4409,In_96,In_282);
and U4410 (N_4410,In_374,In_26);
nand U4411 (N_4411,In_427,In_377);
or U4412 (N_4412,In_82,In_841);
nor U4413 (N_4413,In_195,In_270);
nor U4414 (N_4414,In_830,In_722);
or U4415 (N_4415,In_980,In_66);
and U4416 (N_4416,In_496,In_907);
or U4417 (N_4417,In_632,In_4);
and U4418 (N_4418,In_234,In_147);
xnor U4419 (N_4419,In_135,In_824);
xor U4420 (N_4420,In_60,In_188);
or U4421 (N_4421,In_562,In_804);
and U4422 (N_4422,In_518,In_82);
nand U4423 (N_4423,In_423,In_685);
nand U4424 (N_4424,In_718,In_392);
nand U4425 (N_4425,In_305,In_515);
xor U4426 (N_4426,In_304,In_859);
or U4427 (N_4427,In_17,In_109);
xor U4428 (N_4428,In_950,In_537);
nor U4429 (N_4429,In_506,In_923);
and U4430 (N_4430,In_723,In_23);
and U4431 (N_4431,In_723,In_24);
and U4432 (N_4432,In_357,In_997);
nor U4433 (N_4433,In_961,In_289);
and U4434 (N_4434,In_704,In_689);
nand U4435 (N_4435,In_310,In_618);
or U4436 (N_4436,In_839,In_442);
or U4437 (N_4437,In_584,In_521);
and U4438 (N_4438,In_637,In_830);
nand U4439 (N_4439,In_329,In_817);
and U4440 (N_4440,In_879,In_574);
or U4441 (N_4441,In_91,In_270);
nor U4442 (N_4442,In_645,In_367);
xnor U4443 (N_4443,In_566,In_641);
and U4444 (N_4444,In_416,In_460);
and U4445 (N_4445,In_532,In_723);
or U4446 (N_4446,In_850,In_630);
or U4447 (N_4447,In_106,In_831);
and U4448 (N_4448,In_96,In_754);
and U4449 (N_4449,In_892,In_933);
and U4450 (N_4450,In_0,In_305);
and U4451 (N_4451,In_962,In_288);
nor U4452 (N_4452,In_816,In_116);
xor U4453 (N_4453,In_141,In_810);
xnor U4454 (N_4454,In_727,In_719);
nor U4455 (N_4455,In_577,In_468);
xnor U4456 (N_4456,In_85,In_850);
and U4457 (N_4457,In_605,In_325);
nor U4458 (N_4458,In_731,In_517);
nand U4459 (N_4459,In_265,In_749);
and U4460 (N_4460,In_297,In_134);
and U4461 (N_4461,In_442,In_5);
xor U4462 (N_4462,In_231,In_349);
xor U4463 (N_4463,In_406,In_594);
nand U4464 (N_4464,In_812,In_7);
nor U4465 (N_4465,In_865,In_465);
xnor U4466 (N_4466,In_427,In_232);
and U4467 (N_4467,In_319,In_12);
or U4468 (N_4468,In_547,In_63);
nand U4469 (N_4469,In_9,In_758);
nor U4470 (N_4470,In_400,In_920);
or U4471 (N_4471,In_659,In_782);
nand U4472 (N_4472,In_999,In_642);
or U4473 (N_4473,In_76,In_210);
nand U4474 (N_4474,In_493,In_292);
and U4475 (N_4475,In_948,In_363);
and U4476 (N_4476,In_783,In_326);
or U4477 (N_4477,In_830,In_567);
xor U4478 (N_4478,In_841,In_525);
and U4479 (N_4479,In_534,In_177);
or U4480 (N_4480,In_334,In_784);
nor U4481 (N_4481,In_899,In_276);
nand U4482 (N_4482,In_524,In_168);
and U4483 (N_4483,In_780,In_609);
and U4484 (N_4484,In_530,In_988);
nor U4485 (N_4485,In_633,In_17);
and U4486 (N_4486,In_71,In_689);
nand U4487 (N_4487,In_553,In_124);
xnor U4488 (N_4488,In_105,In_803);
and U4489 (N_4489,In_917,In_294);
and U4490 (N_4490,In_602,In_382);
or U4491 (N_4491,In_431,In_318);
nand U4492 (N_4492,In_974,In_460);
and U4493 (N_4493,In_946,In_215);
or U4494 (N_4494,In_672,In_704);
nand U4495 (N_4495,In_406,In_4);
xor U4496 (N_4496,In_454,In_116);
nor U4497 (N_4497,In_292,In_919);
xor U4498 (N_4498,In_198,In_693);
and U4499 (N_4499,In_371,In_289);
or U4500 (N_4500,In_337,In_176);
nand U4501 (N_4501,In_296,In_848);
nor U4502 (N_4502,In_772,In_451);
or U4503 (N_4503,In_823,In_807);
nand U4504 (N_4504,In_676,In_350);
nand U4505 (N_4505,In_77,In_360);
nand U4506 (N_4506,In_781,In_445);
nand U4507 (N_4507,In_771,In_283);
nand U4508 (N_4508,In_749,In_550);
or U4509 (N_4509,In_310,In_664);
nand U4510 (N_4510,In_575,In_858);
and U4511 (N_4511,In_898,In_428);
nor U4512 (N_4512,In_889,In_575);
nor U4513 (N_4513,In_452,In_734);
xnor U4514 (N_4514,In_237,In_964);
or U4515 (N_4515,In_727,In_883);
xor U4516 (N_4516,In_723,In_63);
nand U4517 (N_4517,In_101,In_706);
nor U4518 (N_4518,In_454,In_312);
nor U4519 (N_4519,In_169,In_17);
and U4520 (N_4520,In_982,In_468);
nand U4521 (N_4521,In_402,In_447);
and U4522 (N_4522,In_4,In_93);
or U4523 (N_4523,In_69,In_74);
nor U4524 (N_4524,In_673,In_655);
nand U4525 (N_4525,In_238,In_549);
and U4526 (N_4526,In_35,In_945);
xnor U4527 (N_4527,In_844,In_649);
nor U4528 (N_4528,In_296,In_159);
or U4529 (N_4529,In_843,In_620);
and U4530 (N_4530,In_406,In_696);
and U4531 (N_4531,In_394,In_927);
and U4532 (N_4532,In_837,In_857);
or U4533 (N_4533,In_253,In_267);
nand U4534 (N_4534,In_536,In_790);
nand U4535 (N_4535,In_560,In_356);
and U4536 (N_4536,In_937,In_585);
or U4537 (N_4537,In_4,In_240);
nand U4538 (N_4538,In_381,In_777);
nor U4539 (N_4539,In_531,In_20);
nand U4540 (N_4540,In_244,In_651);
xor U4541 (N_4541,In_801,In_122);
or U4542 (N_4542,In_499,In_339);
and U4543 (N_4543,In_214,In_275);
nor U4544 (N_4544,In_492,In_306);
and U4545 (N_4545,In_261,In_600);
and U4546 (N_4546,In_120,In_710);
nand U4547 (N_4547,In_89,In_331);
nand U4548 (N_4548,In_468,In_144);
and U4549 (N_4549,In_686,In_154);
or U4550 (N_4550,In_483,In_268);
nor U4551 (N_4551,In_599,In_609);
or U4552 (N_4552,In_352,In_874);
nand U4553 (N_4553,In_524,In_987);
and U4554 (N_4554,In_261,In_451);
and U4555 (N_4555,In_373,In_201);
or U4556 (N_4556,In_955,In_843);
and U4557 (N_4557,In_713,In_244);
nor U4558 (N_4558,In_724,In_860);
nand U4559 (N_4559,In_10,In_965);
or U4560 (N_4560,In_986,In_321);
nor U4561 (N_4561,In_931,In_885);
and U4562 (N_4562,In_945,In_659);
and U4563 (N_4563,In_924,In_535);
nand U4564 (N_4564,In_795,In_758);
nand U4565 (N_4565,In_782,In_654);
and U4566 (N_4566,In_978,In_428);
and U4567 (N_4567,In_685,In_770);
and U4568 (N_4568,In_877,In_60);
nor U4569 (N_4569,In_600,In_314);
xnor U4570 (N_4570,In_248,In_446);
xor U4571 (N_4571,In_714,In_170);
or U4572 (N_4572,In_317,In_657);
and U4573 (N_4573,In_829,In_997);
or U4574 (N_4574,In_465,In_491);
and U4575 (N_4575,In_735,In_160);
or U4576 (N_4576,In_453,In_943);
xor U4577 (N_4577,In_453,In_308);
nor U4578 (N_4578,In_515,In_136);
nor U4579 (N_4579,In_926,In_942);
nand U4580 (N_4580,In_517,In_951);
nand U4581 (N_4581,In_737,In_525);
or U4582 (N_4582,In_405,In_373);
nand U4583 (N_4583,In_58,In_992);
and U4584 (N_4584,In_262,In_758);
or U4585 (N_4585,In_660,In_485);
and U4586 (N_4586,In_950,In_252);
xnor U4587 (N_4587,In_489,In_748);
and U4588 (N_4588,In_151,In_331);
and U4589 (N_4589,In_85,In_516);
xor U4590 (N_4590,In_955,In_478);
or U4591 (N_4591,In_599,In_150);
nand U4592 (N_4592,In_457,In_253);
or U4593 (N_4593,In_788,In_367);
or U4594 (N_4594,In_213,In_194);
or U4595 (N_4595,In_679,In_971);
nand U4596 (N_4596,In_631,In_410);
nor U4597 (N_4597,In_708,In_803);
and U4598 (N_4598,In_718,In_727);
and U4599 (N_4599,In_478,In_93);
xor U4600 (N_4600,In_190,In_364);
and U4601 (N_4601,In_207,In_575);
nor U4602 (N_4602,In_143,In_430);
or U4603 (N_4603,In_808,In_257);
or U4604 (N_4604,In_333,In_728);
or U4605 (N_4605,In_391,In_767);
nand U4606 (N_4606,In_172,In_404);
or U4607 (N_4607,In_855,In_915);
nor U4608 (N_4608,In_410,In_993);
nand U4609 (N_4609,In_356,In_934);
nand U4610 (N_4610,In_585,In_460);
or U4611 (N_4611,In_296,In_90);
nand U4612 (N_4612,In_253,In_733);
and U4613 (N_4613,In_453,In_183);
or U4614 (N_4614,In_425,In_473);
nand U4615 (N_4615,In_247,In_39);
nand U4616 (N_4616,In_559,In_471);
nand U4617 (N_4617,In_340,In_515);
nand U4618 (N_4618,In_351,In_575);
nor U4619 (N_4619,In_108,In_621);
nand U4620 (N_4620,In_285,In_538);
nor U4621 (N_4621,In_429,In_494);
or U4622 (N_4622,In_697,In_235);
nor U4623 (N_4623,In_419,In_24);
nor U4624 (N_4624,In_241,In_453);
nor U4625 (N_4625,In_372,In_482);
nor U4626 (N_4626,In_638,In_347);
or U4627 (N_4627,In_488,In_454);
or U4628 (N_4628,In_203,In_162);
and U4629 (N_4629,In_616,In_763);
and U4630 (N_4630,In_594,In_528);
and U4631 (N_4631,In_204,In_299);
nor U4632 (N_4632,In_624,In_714);
and U4633 (N_4633,In_671,In_372);
nand U4634 (N_4634,In_994,In_149);
or U4635 (N_4635,In_815,In_308);
nand U4636 (N_4636,In_953,In_6);
or U4637 (N_4637,In_577,In_532);
and U4638 (N_4638,In_946,In_646);
or U4639 (N_4639,In_320,In_516);
or U4640 (N_4640,In_229,In_391);
xor U4641 (N_4641,In_777,In_327);
or U4642 (N_4642,In_836,In_56);
or U4643 (N_4643,In_22,In_843);
or U4644 (N_4644,In_561,In_145);
or U4645 (N_4645,In_496,In_123);
or U4646 (N_4646,In_64,In_516);
xor U4647 (N_4647,In_402,In_222);
or U4648 (N_4648,In_229,In_346);
nor U4649 (N_4649,In_289,In_211);
or U4650 (N_4650,In_977,In_964);
nand U4651 (N_4651,In_52,In_858);
nor U4652 (N_4652,In_73,In_179);
nor U4653 (N_4653,In_351,In_919);
xor U4654 (N_4654,In_392,In_380);
nand U4655 (N_4655,In_655,In_312);
nand U4656 (N_4656,In_985,In_960);
nor U4657 (N_4657,In_671,In_890);
and U4658 (N_4658,In_269,In_668);
or U4659 (N_4659,In_395,In_736);
xnor U4660 (N_4660,In_324,In_808);
nand U4661 (N_4661,In_724,In_20);
nor U4662 (N_4662,In_104,In_893);
and U4663 (N_4663,In_707,In_392);
nand U4664 (N_4664,In_641,In_418);
or U4665 (N_4665,In_777,In_40);
and U4666 (N_4666,In_649,In_615);
or U4667 (N_4667,In_711,In_960);
nand U4668 (N_4668,In_434,In_761);
and U4669 (N_4669,In_773,In_542);
nor U4670 (N_4670,In_175,In_777);
nor U4671 (N_4671,In_69,In_456);
nand U4672 (N_4672,In_672,In_66);
nand U4673 (N_4673,In_885,In_336);
or U4674 (N_4674,In_466,In_926);
nor U4675 (N_4675,In_884,In_120);
xor U4676 (N_4676,In_731,In_473);
or U4677 (N_4677,In_18,In_159);
nor U4678 (N_4678,In_778,In_951);
and U4679 (N_4679,In_730,In_387);
nand U4680 (N_4680,In_642,In_121);
nor U4681 (N_4681,In_749,In_540);
xor U4682 (N_4682,In_199,In_314);
and U4683 (N_4683,In_49,In_414);
nor U4684 (N_4684,In_958,In_639);
xor U4685 (N_4685,In_147,In_778);
or U4686 (N_4686,In_269,In_285);
and U4687 (N_4687,In_855,In_293);
or U4688 (N_4688,In_215,In_463);
nand U4689 (N_4689,In_454,In_588);
and U4690 (N_4690,In_763,In_37);
and U4691 (N_4691,In_501,In_826);
nand U4692 (N_4692,In_365,In_548);
or U4693 (N_4693,In_520,In_773);
and U4694 (N_4694,In_143,In_113);
nand U4695 (N_4695,In_112,In_890);
nand U4696 (N_4696,In_825,In_656);
or U4697 (N_4697,In_217,In_240);
nand U4698 (N_4698,In_79,In_763);
nor U4699 (N_4699,In_680,In_474);
or U4700 (N_4700,In_525,In_497);
nand U4701 (N_4701,In_337,In_41);
or U4702 (N_4702,In_689,In_979);
or U4703 (N_4703,In_74,In_870);
nand U4704 (N_4704,In_828,In_894);
xor U4705 (N_4705,In_996,In_926);
or U4706 (N_4706,In_730,In_307);
or U4707 (N_4707,In_707,In_518);
nand U4708 (N_4708,In_994,In_382);
and U4709 (N_4709,In_820,In_447);
and U4710 (N_4710,In_134,In_919);
xor U4711 (N_4711,In_791,In_75);
xnor U4712 (N_4712,In_918,In_976);
xor U4713 (N_4713,In_759,In_984);
nor U4714 (N_4714,In_688,In_231);
or U4715 (N_4715,In_375,In_636);
nand U4716 (N_4716,In_478,In_414);
nor U4717 (N_4717,In_406,In_426);
nand U4718 (N_4718,In_488,In_804);
and U4719 (N_4719,In_182,In_689);
nand U4720 (N_4720,In_51,In_561);
or U4721 (N_4721,In_526,In_640);
and U4722 (N_4722,In_357,In_386);
and U4723 (N_4723,In_327,In_795);
xor U4724 (N_4724,In_478,In_775);
or U4725 (N_4725,In_354,In_837);
nor U4726 (N_4726,In_469,In_644);
nor U4727 (N_4727,In_8,In_366);
and U4728 (N_4728,In_142,In_747);
or U4729 (N_4729,In_788,In_502);
nor U4730 (N_4730,In_917,In_867);
nor U4731 (N_4731,In_650,In_709);
nand U4732 (N_4732,In_464,In_88);
nand U4733 (N_4733,In_758,In_214);
nand U4734 (N_4734,In_843,In_389);
nor U4735 (N_4735,In_378,In_996);
and U4736 (N_4736,In_453,In_22);
and U4737 (N_4737,In_996,In_584);
or U4738 (N_4738,In_513,In_32);
and U4739 (N_4739,In_617,In_212);
and U4740 (N_4740,In_133,In_712);
nor U4741 (N_4741,In_955,In_909);
nand U4742 (N_4742,In_477,In_656);
nand U4743 (N_4743,In_733,In_707);
and U4744 (N_4744,In_155,In_768);
or U4745 (N_4745,In_246,In_225);
nand U4746 (N_4746,In_358,In_462);
nor U4747 (N_4747,In_222,In_420);
nand U4748 (N_4748,In_142,In_508);
nor U4749 (N_4749,In_196,In_427);
nand U4750 (N_4750,In_498,In_344);
nor U4751 (N_4751,In_397,In_413);
and U4752 (N_4752,In_375,In_310);
or U4753 (N_4753,In_301,In_919);
nand U4754 (N_4754,In_41,In_537);
or U4755 (N_4755,In_388,In_471);
or U4756 (N_4756,In_114,In_844);
and U4757 (N_4757,In_578,In_125);
and U4758 (N_4758,In_910,In_784);
and U4759 (N_4759,In_651,In_167);
or U4760 (N_4760,In_779,In_568);
nor U4761 (N_4761,In_942,In_524);
nor U4762 (N_4762,In_602,In_284);
nand U4763 (N_4763,In_288,In_907);
or U4764 (N_4764,In_799,In_758);
xnor U4765 (N_4765,In_598,In_98);
or U4766 (N_4766,In_386,In_584);
nor U4767 (N_4767,In_844,In_980);
nand U4768 (N_4768,In_14,In_954);
nand U4769 (N_4769,In_232,In_428);
and U4770 (N_4770,In_803,In_723);
or U4771 (N_4771,In_5,In_851);
nand U4772 (N_4772,In_672,In_732);
and U4773 (N_4773,In_149,In_48);
and U4774 (N_4774,In_367,In_859);
or U4775 (N_4775,In_332,In_499);
and U4776 (N_4776,In_922,In_802);
nand U4777 (N_4777,In_831,In_892);
or U4778 (N_4778,In_450,In_702);
nand U4779 (N_4779,In_108,In_514);
or U4780 (N_4780,In_639,In_15);
and U4781 (N_4781,In_553,In_473);
nand U4782 (N_4782,In_314,In_427);
nand U4783 (N_4783,In_598,In_132);
and U4784 (N_4784,In_194,In_183);
nand U4785 (N_4785,In_749,In_682);
and U4786 (N_4786,In_78,In_160);
or U4787 (N_4787,In_0,In_595);
xor U4788 (N_4788,In_392,In_299);
nand U4789 (N_4789,In_290,In_691);
and U4790 (N_4790,In_66,In_104);
and U4791 (N_4791,In_583,In_135);
nand U4792 (N_4792,In_19,In_721);
and U4793 (N_4793,In_707,In_276);
and U4794 (N_4794,In_533,In_203);
and U4795 (N_4795,In_464,In_439);
or U4796 (N_4796,In_670,In_316);
and U4797 (N_4797,In_234,In_893);
nand U4798 (N_4798,In_573,In_945);
nor U4799 (N_4799,In_466,In_856);
nor U4800 (N_4800,In_680,In_152);
nand U4801 (N_4801,In_54,In_116);
xor U4802 (N_4802,In_296,In_774);
xor U4803 (N_4803,In_36,In_544);
nor U4804 (N_4804,In_203,In_959);
nor U4805 (N_4805,In_606,In_842);
nand U4806 (N_4806,In_624,In_602);
and U4807 (N_4807,In_325,In_836);
and U4808 (N_4808,In_790,In_416);
nor U4809 (N_4809,In_780,In_948);
xor U4810 (N_4810,In_181,In_39);
nor U4811 (N_4811,In_636,In_285);
xor U4812 (N_4812,In_922,In_276);
or U4813 (N_4813,In_714,In_609);
nand U4814 (N_4814,In_21,In_903);
nand U4815 (N_4815,In_490,In_909);
nor U4816 (N_4816,In_297,In_77);
nor U4817 (N_4817,In_125,In_132);
and U4818 (N_4818,In_184,In_863);
nor U4819 (N_4819,In_344,In_180);
nor U4820 (N_4820,In_913,In_24);
xnor U4821 (N_4821,In_369,In_893);
nand U4822 (N_4822,In_806,In_542);
nand U4823 (N_4823,In_920,In_403);
nor U4824 (N_4824,In_509,In_147);
nand U4825 (N_4825,In_862,In_196);
nand U4826 (N_4826,In_723,In_115);
nor U4827 (N_4827,In_396,In_578);
or U4828 (N_4828,In_816,In_486);
or U4829 (N_4829,In_513,In_808);
or U4830 (N_4830,In_825,In_15);
nor U4831 (N_4831,In_294,In_572);
and U4832 (N_4832,In_419,In_31);
nor U4833 (N_4833,In_430,In_636);
and U4834 (N_4834,In_320,In_161);
and U4835 (N_4835,In_852,In_836);
xor U4836 (N_4836,In_243,In_847);
and U4837 (N_4837,In_343,In_345);
or U4838 (N_4838,In_505,In_838);
and U4839 (N_4839,In_298,In_589);
nor U4840 (N_4840,In_623,In_859);
xor U4841 (N_4841,In_100,In_942);
or U4842 (N_4842,In_728,In_423);
and U4843 (N_4843,In_533,In_693);
and U4844 (N_4844,In_291,In_749);
nand U4845 (N_4845,In_960,In_618);
nor U4846 (N_4846,In_948,In_983);
nor U4847 (N_4847,In_113,In_724);
nor U4848 (N_4848,In_428,In_606);
nand U4849 (N_4849,In_623,In_768);
or U4850 (N_4850,In_548,In_828);
and U4851 (N_4851,In_666,In_287);
nand U4852 (N_4852,In_332,In_701);
nor U4853 (N_4853,In_290,In_852);
nor U4854 (N_4854,In_289,In_482);
or U4855 (N_4855,In_531,In_744);
nand U4856 (N_4856,In_832,In_379);
nand U4857 (N_4857,In_668,In_445);
and U4858 (N_4858,In_700,In_596);
and U4859 (N_4859,In_103,In_743);
xor U4860 (N_4860,In_985,In_635);
and U4861 (N_4861,In_49,In_447);
or U4862 (N_4862,In_499,In_746);
nand U4863 (N_4863,In_777,In_670);
nor U4864 (N_4864,In_624,In_621);
nand U4865 (N_4865,In_392,In_915);
nor U4866 (N_4866,In_384,In_549);
or U4867 (N_4867,In_276,In_659);
and U4868 (N_4868,In_142,In_547);
and U4869 (N_4869,In_304,In_217);
and U4870 (N_4870,In_630,In_12);
or U4871 (N_4871,In_53,In_522);
or U4872 (N_4872,In_672,In_662);
nand U4873 (N_4873,In_315,In_821);
nor U4874 (N_4874,In_173,In_853);
nand U4875 (N_4875,In_557,In_469);
nor U4876 (N_4876,In_859,In_337);
nand U4877 (N_4877,In_917,In_579);
xnor U4878 (N_4878,In_444,In_410);
and U4879 (N_4879,In_986,In_402);
and U4880 (N_4880,In_846,In_600);
xnor U4881 (N_4881,In_895,In_737);
xnor U4882 (N_4882,In_770,In_718);
nor U4883 (N_4883,In_151,In_922);
or U4884 (N_4884,In_732,In_496);
nor U4885 (N_4885,In_868,In_63);
or U4886 (N_4886,In_108,In_201);
nand U4887 (N_4887,In_105,In_911);
xnor U4888 (N_4888,In_241,In_229);
nand U4889 (N_4889,In_916,In_596);
and U4890 (N_4890,In_90,In_327);
nand U4891 (N_4891,In_963,In_999);
and U4892 (N_4892,In_601,In_887);
and U4893 (N_4893,In_161,In_690);
nand U4894 (N_4894,In_105,In_496);
nand U4895 (N_4895,In_247,In_78);
and U4896 (N_4896,In_237,In_200);
and U4897 (N_4897,In_905,In_455);
nor U4898 (N_4898,In_523,In_204);
xnor U4899 (N_4899,In_340,In_30);
xor U4900 (N_4900,In_230,In_929);
nor U4901 (N_4901,In_467,In_919);
or U4902 (N_4902,In_414,In_28);
and U4903 (N_4903,In_701,In_476);
nor U4904 (N_4904,In_481,In_305);
nand U4905 (N_4905,In_396,In_918);
nor U4906 (N_4906,In_517,In_196);
and U4907 (N_4907,In_558,In_398);
or U4908 (N_4908,In_260,In_92);
or U4909 (N_4909,In_433,In_761);
xnor U4910 (N_4910,In_113,In_70);
or U4911 (N_4911,In_898,In_17);
nor U4912 (N_4912,In_13,In_246);
or U4913 (N_4913,In_936,In_581);
or U4914 (N_4914,In_532,In_574);
nor U4915 (N_4915,In_290,In_54);
nand U4916 (N_4916,In_178,In_311);
and U4917 (N_4917,In_258,In_787);
or U4918 (N_4918,In_139,In_574);
or U4919 (N_4919,In_381,In_228);
or U4920 (N_4920,In_413,In_473);
nor U4921 (N_4921,In_705,In_65);
or U4922 (N_4922,In_411,In_903);
nand U4923 (N_4923,In_936,In_1);
nor U4924 (N_4924,In_741,In_714);
nand U4925 (N_4925,In_111,In_669);
and U4926 (N_4926,In_765,In_271);
nand U4927 (N_4927,In_467,In_402);
xnor U4928 (N_4928,In_175,In_312);
nand U4929 (N_4929,In_386,In_160);
and U4930 (N_4930,In_893,In_756);
and U4931 (N_4931,In_770,In_612);
xnor U4932 (N_4932,In_898,In_531);
nand U4933 (N_4933,In_256,In_478);
or U4934 (N_4934,In_474,In_371);
nor U4935 (N_4935,In_2,In_343);
nor U4936 (N_4936,In_930,In_759);
and U4937 (N_4937,In_243,In_302);
nor U4938 (N_4938,In_685,In_734);
or U4939 (N_4939,In_773,In_353);
and U4940 (N_4940,In_475,In_640);
nor U4941 (N_4941,In_87,In_169);
nand U4942 (N_4942,In_186,In_503);
nand U4943 (N_4943,In_129,In_230);
nor U4944 (N_4944,In_903,In_548);
nor U4945 (N_4945,In_581,In_72);
xnor U4946 (N_4946,In_246,In_410);
or U4947 (N_4947,In_927,In_455);
and U4948 (N_4948,In_850,In_894);
nor U4949 (N_4949,In_385,In_438);
nor U4950 (N_4950,In_188,In_916);
nor U4951 (N_4951,In_159,In_867);
nor U4952 (N_4952,In_298,In_44);
and U4953 (N_4953,In_781,In_174);
or U4954 (N_4954,In_643,In_446);
and U4955 (N_4955,In_116,In_259);
or U4956 (N_4956,In_662,In_302);
nand U4957 (N_4957,In_285,In_149);
nand U4958 (N_4958,In_133,In_885);
and U4959 (N_4959,In_914,In_530);
nand U4960 (N_4960,In_490,In_847);
and U4961 (N_4961,In_309,In_256);
nand U4962 (N_4962,In_502,In_76);
xor U4963 (N_4963,In_278,In_170);
xnor U4964 (N_4964,In_45,In_850);
or U4965 (N_4965,In_993,In_299);
nand U4966 (N_4966,In_591,In_989);
nand U4967 (N_4967,In_889,In_341);
or U4968 (N_4968,In_254,In_488);
or U4969 (N_4969,In_637,In_686);
xnor U4970 (N_4970,In_625,In_741);
or U4971 (N_4971,In_78,In_80);
or U4972 (N_4972,In_269,In_101);
nor U4973 (N_4973,In_693,In_349);
nand U4974 (N_4974,In_634,In_517);
nand U4975 (N_4975,In_23,In_970);
nor U4976 (N_4976,In_390,In_591);
nand U4977 (N_4977,In_45,In_513);
nor U4978 (N_4978,In_672,In_731);
nor U4979 (N_4979,In_75,In_851);
xor U4980 (N_4980,In_918,In_966);
and U4981 (N_4981,In_649,In_67);
nor U4982 (N_4982,In_517,In_32);
xor U4983 (N_4983,In_98,In_723);
nor U4984 (N_4984,In_471,In_586);
and U4985 (N_4985,In_619,In_163);
nand U4986 (N_4986,In_769,In_195);
nor U4987 (N_4987,In_603,In_936);
or U4988 (N_4988,In_949,In_804);
nor U4989 (N_4989,In_386,In_567);
nor U4990 (N_4990,In_472,In_613);
nor U4991 (N_4991,In_210,In_457);
or U4992 (N_4992,In_787,In_741);
nand U4993 (N_4993,In_995,In_926);
xnor U4994 (N_4994,In_566,In_44);
and U4995 (N_4995,In_176,In_698);
or U4996 (N_4996,In_384,In_887);
nand U4997 (N_4997,In_70,In_178);
and U4998 (N_4998,In_882,In_165);
and U4999 (N_4999,In_143,In_424);
nand U5000 (N_5000,N_4129,N_2261);
nand U5001 (N_5001,N_2298,N_4389);
or U5002 (N_5002,N_2970,N_2587);
nor U5003 (N_5003,N_3557,N_3691);
or U5004 (N_5004,N_2734,N_2711);
and U5005 (N_5005,N_452,N_2500);
nor U5006 (N_5006,N_1904,N_1446);
and U5007 (N_5007,N_4326,N_1896);
and U5008 (N_5008,N_3439,N_2764);
and U5009 (N_5009,N_4633,N_3820);
and U5010 (N_5010,N_2015,N_3734);
and U5011 (N_5011,N_3620,N_197);
nor U5012 (N_5012,N_4844,N_784);
nand U5013 (N_5013,N_208,N_3462);
nand U5014 (N_5014,N_1353,N_3002);
or U5015 (N_5015,N_2930,N_1911);
and U5016 (N_5016,N_569,N_2851);
and U5017 (N_5017,N_3019,N_566);
and U5018 (N_5018,N_1409,N_133);
and U5019 (N_5019,N_1354,N_533);
and U5020 (N_5020,N_4727,N_1421);
or U5021 (N_5021,N_3355,N_2749);
xor U5022 (N_5022,N_69,N_4851);
or U5023 (N_5023,N_2598,N_1618);
nand U5024 (N_5024,N_2957,N_2714);
nand U5025 (N_5025,N_4086,N_808);
and U5026 (N_5026,N_316,N_1096);
and U5027 (N_5027,N_4678,N_3366);
and U5028 (N_5028,N_1413,N_2388);
and U5029 (N_5029,N_962,N_413);
and U5030 (N_5030,N_4380,N_2637);
or U5031 (N_5031,N_188,N_1633);
nor U5032 (N_5032,N_371,N_4765);
nand U5033 (N_5033,N_3265,N_4336);
nor U5034 (N_5034,N_933,N_3096);
and U5035 (N_5035,N_2421,N_3376);
xnor U5036 (N_5036,N_4609,N_4206);
or U5037 (N_5037,N_1532,N_168);
and U5038 (N_5038,N_2748,N_4871);
nand U5039 (N_5039,N_4147,N_3473);
or U5040 (N_5040,N_1542,N_2408);
nand U5041 (N_5041,N_3252,N_2457);
nor U5042 (N_5042,N_1712,N_826);
xor U5043 (N_5043,N_3505,N_4724);
or U5044 (N_5044,N_966,N_1714);
and U5045 (N_5045,N_3759,N_3465);
xnor U5046 (N_5046,N_3698,N_2493);
nand U5047 (N_5047,N_4707,N_4733);
nor U5048 (N_5048,N_3735,N_1047);
and U5049 (N_5049,N_3203,N_3534);
nor U5050 (N_5050,N_1190,N_2081);
or U5051 (N_5051,N_2596,N_1098);
and U5052 (N_5052,N_4210,N_3486);
nor U5053 (N_5053,N_1253,N_779);
or U5054 (N_5054,N_3843,N_2439);
xor U5055 (N_5055,N_3222,N_4907);
nand U5056 (N_5056,N_714,N_899);
and U5057 (N_5057,N_3240,N_4556);
xor U5058 (N_5058,N_3730,N_2316);
and U5059 (N_5059,N_2757,N_1246);
xnor U5060 (N_5060,N_2726,N_1495);
nand U5061 (N_5061,N_1311,N_4679);
nand U5062 (N_5062,N_2713,N_11);
nand U5063 (N_5063,N_2869,N_2833);
nor U5064 (N_5064,N_2514,N_2969);
and U5065 (N_5065,N_1772,N_3255);
or U5066 (N_5066,N_4261,N_1033);
xor U5067 (N_5067,N_4714,N_2667);
and U5068 (N_5068,N_2007,N_4876);
xnor U5069 (N_5069,N_2831,N_2622);
nor U5070 (N_5070,N_2110,N_3765);
xor U5071 (N_5071,N_4391,N_1068);
nand U5072 (N_5072,N_1999,N_2903);
and U5073 (N_5073,N_3297,N_3409);
nor U5074 (N_5074,N_3681,N_4295);
nor U5075 (N_5075,N_3290,N_3024);
xor U5076 (N_5076,N_4070,N_4974);
nand U5077 (N_5077,N_3242,N_4761);
nand U5078 (N_5078,N_2498,N_4832);
nor U5079 (N_5079,N_4066,N_3530);
nor U5080 (N_5080,N_3960,N_2156);
and U5081 (N_5081,N_4032,N_4209);
nor U5082 (N_5082,N_2504,N_1721);
nand U5083 (N_5083,N_1523,N_2280);
and U5084 (N_5084,N_428,N_1458);
or U5085 (N_5085,N_1473,N_1244);
or U5086 (N_5086,N_4596,N_1436);
and U5087 (N_5087,N_4578,N_2818);
nand U5088 (N_5088,N_957,N_3151);
nand U5089 (N_5089,N_4589,N_1137);
or U5090 (N_5090,N_1742,N_4008);
xor U5091 (N_5091,N_821,N_4890);
nor U5092 (N_5092,N_406,N_3042);
nor U5093 (N_5093,N_3635,N_4619);
nor U5094 (N_5094,N_1329,N_3933);
and U5095 (N_5095,N_4370,N_3496);
or U5096 (N_5096,N_2387,N_1386);
nand U5097 (N_5097,N_1502,N_205);
and U5098 (N_5098,N_2306,N_4669);
nor U5099 (N_5099,N_1653,N_397);
and U5100 (N_5100,N_2299,N_2509);
nor U5101 (N_5101,N_4971,N_588);
and U5102 (N_5102,N_362,N_3440);
nor U5103 (N_5103,N_1320,N_283);
nand U5104 (N_5104,N_4927,N_2894);
and U5105 (N_5105,N_30,N_1583);
or U5106 (N_5106,N_4401,N_3443);
nor U5107 (N_5107,N_4170,N_4011);
nand U5108 (N_5108,N_1148,N_4176);
nand U5109 (N_5109,N_1312,N_4012);
nor U5110 (N_5110,N_2750,N_4910);
nor U5111 (N_5111,N_4361,N_128);
and U5112 (N_5112,N_4037,N_2131);
nor U5113 (N_5113,N_4813,N_4899);
xor U5114 (N_5114,N_1063,N_1955);
nand U5115 (N_5115,N_3041,N_4660);
or U5116 (N_5116,N_2349,N_3060);
nand U5117 (N_5117,N_121,N_2135);
nor U5118 (N_5118,N_1025,N_4508);
and U5119 (N_5119,N_3246,N_1467);
or U5120 (N_5120,N_1303,N_238);
and U5121 (N_5121,N_1321,N_805);
nor U5122 (N_5122,N_2792,N_2270);
or U5123 (N_5123,N_3111,N_1704);
nand U5124 (N_5124,N_4959,N_4985);
and U5125 (N_5125,N_256,N_2255);
or U5126 (N_5126,N_1044,N_1871);
nor U5127 (N_5127,N_3651,N_1609);
nor U5128 (N_5128,N_2758,N_1408);
or U5129 (N_5129,N_2644,N_2835);
nor U5130 (N_5130,N_4978,N_967);
nand U5131 (N_5131,N_1179,N_2410);
or U5132 (N_5132,N_4888,N_1638);
nand U5133 (N_5133,N_3118,N_4148);
nand U5134 (N_5134,N_676,N_1754);
nor U5135 (N_5135,N_4809,N_4515);
nor U5136 (N_5136,N_3160,N_3772);
nand U5137 (N_5137,N_169,N_1572);
and U5138 (N_5138,N_2429,N_3086);
nor U5139 (N_5139,N_2663,N_1974);
and U5140 (N_5140,N_4360,N_1533);
nor U5141 (N_5141,N_4334,N_435);
xor U5142 (N_5142,N_2973,N_2057);
or U5143 (N_5143,N_3179,N_645);
nor U5144 (N_5144,N_2183,N_3892);
xor U5145 (N_5145,N_1128,N_2745);
nand U5146 (N_5146,N_2570,N_2064);
or U5147 (N_5147,N_1689,N_2454);
and U5148 (N_5148,N_4926,N_836);
and U5149 (N_5149,N_509,N_4886);
or U5150 (N_5150,N_323,N_4302);
or U5151 (N_5151,N_360,N_4192);
xor U5152 (N_5152,N_799,N_191);
xnor U5153 (N_5153,N_4098,N_3555);
nor U5154 (N_5154,N_3670,N_4885);
nand U5155 (N_5155,N_4081,N_274);
nor U5156 (N_5156,N_2516,N_4415);
nor U5157 (N_5157,N_4721,N_2247);
nor U5158 (N_5158,N_3447,N_4085);
or U5159 (N_5159,N_4940,N_1953);
or U5160 (N_5160,N_3381,N_776);
xor U5161 (N_5161,N_2508,N_1921);
nor U5162 (N_5162,N_2628,N_2941);
and U5163 (N_5163,N_2134,N_932);
or U5164 (N_5164,N_1782,N_2654);
or U5165 (N_5165,N_4426,N_1182);
or U5166 (N_5166,N_4053,N_3070);
nor U5167 (N_5167,N_3622,N_1392);
xnor U5168 (N_5168,N_2609,N_3221);
and U5169 (N_5169,N_2657,N_522);
xnor U5170 (N_5170,N_1674,N_2790);
nand U5171 (N_5171,N_3148,N_3781);
xor U5172 (N_5172,N_3900,N_2452);
and U5173 (N_5173,N_241,N_2370);
or U5174 (N_5174,N_3858,N_1357);
nand U5175 (N_5175,N_2097,N_3954);
and U5176 (N_5176,N_4156,N_1920);
or U5177 (N_5177,N_1892,N_1693);
or U5178 (N_5178,N_4004,N_3527);
nand U5179 (N_5179,N_4713,N_3586);
or U5180 (N_5180,N_2167,N_3278);
nand U5181 (N_5181,N_3747,N_2677);
or U5182 (N_5182,N_4655,N_3309);
or U5183 (N_5183,N_1091,N_1763);
nand U5184 (N_5184,N_624,N_2271);
or U5185 (N_5185,N_4997,N_503);
nand U5186 (N_5186,N_4625,N_2579);
nor U5187 (N_5187,N_1541,N_2291);
nor U5188 (N_5188,N_4339,N_3834);
and U5189 (N_5189,N_3236,N_2550);
or U5190 (N_5190,N_4812,N_90);
or U5191 (N_5191,N_1133,N_4279);
nand U5192 (N_5192,N_3628,N_127);
or U5193 (N_5193,N_4347,N_2947);
nand U5194 (N_5194,N_3008,N_771);
nor U5195 (N_5195,N_4635,N_3660);
or U5196 (N_5196,N_2779,N_1587);
or U5197 (N_5197,N_1787,N_3626);
nand U5198 (N_5198,N_139,N_2811);
nand U5199 (N_5199,N_2767,N_1812);
and U5200 (N_5200,N_2158,N_4058);
and U5201 (N_5201,N_2463,N_1239);
and U5202 (N_5202,N_3048,N_3972);
nand U5203 (N_5203,N_4403,N_1451);
or U5204 (N_5204,N_2661,N_3342);
or U5205 (N_5205,N_4990,N_4087);
nor U5206 (N_5206,N_3122,N_1435);
and U5207 (N_5207,N_571,N_79);
nand U5208 (N_5208,N_2681,N_544);
or U5209 (N_5209,N_1626,N_3247);
xnor U5210 (N_5210,N_504,N_691);
nand U5211 (N_5211,N_147,N_4740);
and U5212 (N_5212,N_231,N_1582);
nor U5213 (N_5213,N_4205,N_303);
nor U5214 (N_5214,N_3183,N_1792);
nand U5215 (N_5215,N_2958,N_4981);
nand U5216 (N_5216,N_334,N_3187);
or U5217 (N_5217,N_3846,N_4349);
or U5218 (N_5218,N_1290,N_618);
nor U5219 (N_5219,N_3384,N_4617);
nor U5220 (N_5220,N_665,N_574);
nor U5221 (N_5221,N_1255,N_3499);
nand U5222 (N_5222,N_4172,N_3804);
xnor U5223 (N_5223,N_2000,N_2279);
nand U5224 (N_5224,N_4128,N_2806);
nand U5225 (N_5225,N_2394,N_2563);
nand U5226 (N_5226,N_959,N_1732);
nor U5227 (N_5227,N_759,N_3103);
or U5228 (N_5228,N_1794,N_134);
nor U5229 (N_5229,N_2177,N_4542);
xnor U5230 (N_5230,N_4989,N_209);
nand U5231 (N_5231,N_818,N_3708);
nor U5232 (N_5232,N_3885,N_4031);
nand U5233 (N_5233,N_4686,N_174);
or U5234 (N_5234,N_1725,N_2936);
and U5235 (N_5235,N_3271,N_3062);
and U5236 (N_5236,N_4584,N_4750);
and U5237 (N_5237,N_4550,N_602);
and U5238 (N_5238,N_1646,N_151);
nand U5239 (N_5239,N_547,N_4801);
or U5240 (N_5240,N_336,N_4788);
or U5241 (N_5241,N_3040,N_1416);
or U5242 (N_5242,N_2418,N_2397);
and U5243 (N_5243,N_4648,N_1186);
nor U5244 (N_5244,N_439,N_1457);
nor U5245 (N_5245,N_929,N_3225);
nor U5246 (N_5246,N_3344,N_3894);
or U5247 (N_5247,N_4875,N_3579);
nor U5248 (N_5248,N_4757,N_1838);
nor U5249 (N_5249,N_1370,N_3992);
nand U5250 (N_5250,N_3649,N_4963);
nor U5251 (N_5251,N_3185,N_1000);
nor U5252 (N_5252,N_2829,N_4395);
and U5253 (N_5253,N_2816,N_281);
and U5254 (N_5254,N_2744,N_3390);
and U5255 (N_5255,N_4725,N_2216);
and U5256 (N_5256,N_3867,N_4623);
and U5257 (N_5257,N_2868,N_2467);
or U5258 (N_5258,N_814,N_3851);
nand U5259 (N_5259,N_3710,N_2664);
and U5260 (N_5260,N_736,N_4882);
nand U5261 (N_5261,N_2254,N_964);
or U5262 (N_5262,N_717,N_2176);
or U5263 (N_5263,N_388,N_1858);
nor U5264 (N_5264,N_225,N_2486);
xor U5265 (N_5265,N_1954,N_849);
or U5266 (N_5266,N_202,N_4717);
nor U5267 (N_5267,N_2478,N_4807);
and U5268 (N_5268,N_4588,N_3146);
or U5269 (N_5269,N_3169,N_2031);
or U5270 (N_5270,N_847,N_1594);
and U5271 (N_5271,N_3561,N_800);
nand U5272 (N_5272,N_3379,N_2539);
nor U5273 (N_5273,N_1611,N_1374);
nand U5274 (N_5274,N_242,N_2268);
nand U5275 (N_5275,N_1996,N_1511);
or U5276 (N_5276,N_340,N_4568);
nor U5277 (N_5277,N_1129,N_1165);
or U5278 (N_5278,N_260,N_1340);
or U5279 (N_5279,N_1139,N_510);
and U5280 (N_5280,N_1883,N_1987);
nor U5281 (N_5281,N_2554,N_3418);
and U5282 (N_5282,N_2450,N_3969);
or U5283 (N_5283,N_3454,N_690);
nor U5284 (N_5284,N_3196,N_2971);
nor U5285 (N_5285,N_3890,N_1931);
nand U5286 (N_5286,N_3669,N_558);
nand U5287 (N_5287,N_3931,N_240);
nor U5288 (N_5288,N_1298,N_1943);
nor U5289 (N_5289,N_2342,N_253);
nor U5290 (N_5290,N_2094,N_2848);
and U5291 (N_5291,N_1877,N_3982);
nand U5292 (N_5292,N_184,N_1134);
nor U5293 (N_5293,N_1417,N_3206);
nand U5294 (N_5294,N_894,N_2643);
nor U5295 (N_5295,N_4728,N_2945);
nor U5296 (N_5296,N_661,N_1146);
or U5297 (N_5297,N_4581,N_954);
nand U5298 (N_5298,N_3030,N_2368);
xnor U5299 (N_5299,N_4699,N_555);
and U5300 (N_5300,N_2093,N_4739);
or U5301 (N_5301,N_2328,N_2647);
nand U5302 (N_5302,N_791,N_2083);
nor U5303 (N_5303,N_1088,N_1059);
or U5304 (N_5304,N_2464,N_3047);
and U5305 (N_5305,N_3839,N_1575);
and U5306 (N_5306,N_4576,N_3322);
or U5307 (N_5307,N_232,N_2519);
and U5308 (N_5308,N_1160,N_3777);
or U5309 (N_5309,N_4487,N_185);
nand U5310 (N_5310,N_3945,N_3549);
nor U5311 (N_5311,N_3364,N_3827);
xor U5312 (N_5312,N_2112,N_404);
and U5313 (N_5313,N_306,N_1141);
and U5314 (N_5314,N_3633,N_1548);
nand U5315 (N_5315,N_2518,N_255);
or U5316 (N_5316,N_3791,N_4276);
or U5317 (N_5317,N_2905,N_1703);
nand U5318 (N_5318,N_2558,N_696);
nand U5319 (N_5319,N_637,N_4898);
xor U5320 (N_5320,N_4554,N_3090);
xnor U5321 (N_5321,N_511,N_4454);
and U5322 (N_5322,N_1514,N_4586);
and U5323 (N_5323,N_1066,N_1324);
and U5324 (N_5324,N_1115,N_359);
and U5325 (N_5325,N_4796,N_3058);
nand U5326 (N_5326,N_693,N_2787);
xor U5327 (N_5327,N_4993,N_834);
nand U5328 (N_5328,N_2171,N_23);
nor U5329 (N_5329,N_173,N_2440);
nor U5330 (N_5330,N_3458,N_3617);
and U5331 (N_5331,N_1775,N_3091);
and U5332 (N_5332,N_1891,N_3902);
xnor U5333 (N_5333,N_32,N_628);
and U5334 (N_5334,N_4693,N_3871);
and U5335 (N_5335,N_3916,N_4074);
nor U5336 (N_5336,N_3880,N_441);
nand U5337 (N_5337,N_2589,N_4569);
and U5338 (N_5338,N_4273,N_486);
nand U5339 (N_5339,N_4411,N_4649);
nor U5340 (N_5340,N_3550,N_1017);
or U5341 (N_5341,N_138,N_2234);
nor U5342 (N_5342,N_2658,N_1328);
nor U5343 (N_5343,N_73,N_1684);
nor U5344 (N_5344,N_2300,N_1676);
xnor U5345 (N_5345,N_2357,N_4951);
nor U5346 (N_5346,N_4145,N_1530);
or U5347 (N_5347,N_968,N_1472);
nand U5348 (N_5348,N_3373,N_4445);
nand U5349 (N_5349,N_2003,N_29);
nor U5350 (N_5350,N_2593,N_363);
nand U5351 (N_5351,N_3536,N_3789);
and U5352 (N_5352,N_2861,N_2877);
and U5353 (N_5353,N_4518,N_3372);
and U5354 (N_5354,N_2582,N_4294);
and U5355 (N_5355,N_2733,N_2798);
and U5356 (N_5356,N_3877,N_341);
xnor U5357 (N_5357,N_684,N_4121);
nor U5358 (N_5358,N_3343,N_2099);
xor U5359 (N_5359,N_3560,N_4611);
nor U5360 (N_5360,N_577,N_2016);
or U5361 (N_5361,N_2325,N_1961);
nand U5362 (N_5362,N_670,N_2312);
and U5363 (N_5363,N_2295,N_2712);
and U5364 (N_5364,N_2233,N_2351);
and U5365 (N_5365,N_2781,N_4522);
and U5366 (N_5366,N_333,N_4622);
or U5367 (N_5367,N_3737,N_60);
or U5368 (N_5368,N_1391,N_3662);
nand U5369 (N_5369,N_1655,N_1325);
nand U5370 (N_5370,N_2220,N_1993);
nand U5371 (N_5371,N_77,N_1570);
or U5372 (N_5372,N_3718,N_732);
nand U5373 (N_5373,N_2529,N_462);
nor U5374 (N_5374,N_2438,N_3562);
nand U5375 (N_5375,N_4689,N_387);
and U5376 (N_5376,N_99,N_913);
nand U5377 (N_5377,N_2121,N_1737);
or U5378 (N_5378,N_87,N_585);
and U5379 (N_5379,N_2120,N_414);
nand U5380 (N_5380,N_4471,N_4041);
or U5381 (N_5381,N_1699,N_4565);
nand U5382 (N_5382,N_4097,N_55);
nor U5383 (N_5383,N_3816,N_685);
nand U5384 (N_5384,N_2213,N_2547);
nand U5385 (N_5385,N_3218,N_2690);
and U5386 (N_5386,N_4709,N_2446);
nor U5387 (N_5387,N_936,N_3085);
nor U5388 (N_5388,N_2343,N_224);
nand U5389 (N_5389,N_3580,N_523);
or U5390 (N_5390,N_3491,N_158);
and U5391 (N_5391,N_337,N_4025);
nand U5392 (N_5392,N_2926,N_3724);
or U5393 (N_5393,N_1827,N_1997);
nor U5394 (N_5394,N_123,N_287);
nand U5395 (N_5395,N_4266,N_2235);
or U5396 (N_5396,N_1661,N_2577);
nor U5397 (N_5397,N_2686,N_2383);
and U5398 (N_5398,N_4764,N_2460);
nor U5399 (N_5399,N_3251,N_461);
nand U5400 (N_5400,N_2047,N_2739);
xnor U5401 (N_5401,N_3201,N_2885);
and U5402 (N_5402,N_3404,N_4902);
nand U5403 (N_5403,N_1937,N_4972);
nand U5404 (N_5404,N_1230,N_2290);
or U5405 (N_5405,N_4218,N_2495);
nor U5406 (N_5406,N_3300,N_2165);
nand U5407 (N_5407,N_2178,N_425);
nor U5408 (N_5408,N_183,N_2765);
xnor U5409 (N_5409,N_464,N_1579);
nor U5410 (N_5410,N_453,N_2656);
nor U5411 (N_5411,N_1310,N_1121);
nand U5412 (N_5412,N_417,N_3956);
nand U5413 (N_5413,N_3298,N_4333);
and U5414 (N_5414,N_296,N_3646);
nor U5415 (N_5415,N_2374,N_4327);
nand U5416 (N_5416,N_2545,N_4745);
or U5417 (N_5417,N_731,N_4343);
and U5418 (N_5418,N_1500,N_247);
or U5419 (N_5419,N_2159,N_3901);
or U5420 (N_5420,N_4193,N_1166);
nor U5421 (N_5421,N_2573,N_236);
and U5422 (N_5422,N_4760,N_3985);
and U5423 (N_5423,N_2055,N_1142);
or U5424 (N_5424,N_4219,N_2685);
or U5425 (N_5425,N_3369,N_3627);
nor U5426 (N_5426,N_4904,N_1450);
nor U5427 (N_5427,N_3779,N_3406);
xor U5428 (N_5428,N_83,N_2544);
or U5429 (N_5429,N_620,N_4400);
and U5430 (N_5430,N_2068,N_113);
or U5431 (N_5431,N_3519,N_57);
or U5432 (N_5432,N_2489,N_4616);
nor U5433 (N_5433,N_436,N_3887);
nand U5434 (N_5434,N_3093,N_4366);
nor U5435 (N_5435,N_2339,N_746);
and U5436 (N_5436,N_1765,N_4191);
nor U5437 (N_5437,N_2272,N_497);
or U5438 (N_5438,N_2182,N_426);
nand U5439 (N_5439,N_2096,N_1962);
nor U5440 (N_5440,N_212,N_2889);
nand U5441 (N_5441,N_934,N_3405);
and U5442 (N_5442,N_4591,N_2140);
or U5443 (N_5443,N_4592,N_1149);
nand U5444 (N_5444,N_1107,N_1224);
nand U5445 (N_5445,N_2297,N_4230);
or U5446 (N_5446,N_2684,N_1199);
or U5447 (N_5447,N_2997,N_1104);
nor U5448 (N_5448,N_4523,N_4475);
nor U5449 (N_5449,N_2538,N_1164);
nand U5450 (N_5450,N_2257,N_2492);
nand U5451 (N_5451,N_1231,N_4831);
nor U5452 (N_5452,N_1727,N_1613);
nor U5453 (N_5453,N_563,N_3276);
or U5454 (N_5454,N_1358,N_4906);
xnor U5455 (N_5455,N_4,N_1735);
xor U5456 (N_5456,N_148,N_2933);
nand U5457 (N_5457,N_2528,N_3711);
or U5458 (N_5458,N_2990,N_4390);
nand U5459 (N_5459,N_1818,N_1816);
nand U5460 (N_5460,N_4132,N_1934);
nor U5461 (N_5461,N_1398,N_1745);
xnor U5462 (N_5462,N_1665,N_2569);
nand U5463 (N_5463,N_1475,N_2778);
xor U5464 (N_5464,N_367,N_3910);
nor U5465 (N_5465,N_1057,N_617);
nor U5466 (N_5466,N_4892,N_3073);
nand U5467 (N_5467,N_81,N_1881);
and U5468 (N_5468,N_3205,N_4119);
or U5469 (N_5469,N_4911,N_3207);
or U5470 (N_5470,N_905,N_2030);
or U5471 (N_5471,N_2180,N_3361);
and U5472 (N_5472,N_2754,N_4486);
or U5473 (N_5473,N_3483,N_1990);
nand U5474 (N_5474,N_2882,N_3989);
nor U5475 (N_5475,N_3680,N_2395);
or U5476 (N_5476,N_1127,N_537);
nand U5477 (N_5477,N_2303,N_1879);
nor U5478 (N_5478,N_2753,N_423);
nand U5479 (N_5479,N_2723,N_1487);
xnor U5480 (N_5480,N_1539,N_1811);
nor U5481 (N_5481,N_1062,N_2301);
and U5482 (N_5482,N_4930,N_4778);
or U5483 (N_5483,N_3150,N_1885);
nand U5484 (N_5484,N_502,N_3668);
and U5485 (N_5485,N_327,N_2888);
or U5486 (N_5486,N_2608,N_1276);
xnor U5487 (N_5487,N_1259,N_2902);
or U5488 (N_5488,N_4626,N_804);
nand U5489 (N_5489,N_1368,N_1733);
nor U5490 (N_5490,N_2771,N_1946);
nand U5491 (N_5491,N_1364,N_2128);
or U5492 (N_5492,N_1893,N_4536);
xnor U5493 (N_5493,N_4413,N_1173);
nand U5494 (N_5494,N_4941,N_3587);
nand U5495 (N_5495,N_1844,N_2362);
nand U5496 (N_5496,N_431,N_1052);
nor U5497 (N_5497,N_810,N_488);
and U5498 (N_5498,N_44,N_2824);
nor U5499 (N_5499,N_152,N_1029);
nor U5500 (N_5500,N_798,N_4300);
nor U5501 (N_5501,N_4934,N_4237);
nor U5502 (N_5502,N_1598,N_149);
or U5503 (N_5503,N_3007,N_3217);
nand U5504 (N_5504,N_4269,N_2063);
and U5505 (N_5505,N_548,N_3383);
nor U5506 (N_5506,N_3808,N_565);
nand U5507 (N_5507,N_4073,N_3881);
or U5508 (N_5508,N_3479,N_285);
nor U5509 (N_5509,N_2435,N_1257);
nand U5510 (N_5510,N_796,N_679);
nor U5511 (N_5511,N_3727,N_4723);
or U5512 (N_5512,N_377,N_3805);
nor U5513 (N_5513,N_4214,N_2427);
xor U5514 (N_5514,N_4593,N_1861);
nand U5515 (N_5515,N_4239,N_196);
nor U5516 (N_5516,N_3585,N_4002);
and U5517 (N_5517,N_2580,N_1867);
nor U5518 (N_5518,N_4688,N_3911);
nand U5519 (N_5519,N_1747,N_2944);
nand U5520 (N_5520,N_3657,N_2975);
nor U5521 (N_5521,N_383,N_3524);
xor U5522 (N_5522,N_4063,N_3244);
and U5523 (N_5523,N_1766,N_4045);
nand U5524 (N_5524,N_1988,N_2696);
xnor U5525 (N_5525,N_2005,N_2501);
and U5526 (N_5526,N_179,N_2611);
and U5527 (N_5527,N_4384,N_4551);
nand U5528 (N_5528,N_2223,N_2447);
xnor U5529 (N_5529,N_2974,N_663);
nor U5530 (N_5530,N_3666,N_1209);
nand U5531 (N_5531,N_2858,N_875);
xnor U5532 (N_5532,N_4248,N_2708);
xor U5533 (N_5533,N_2595,N_4396);
or U5534 (N_5534,N_1786,N_3744);
xor U5535 (N_5535,N_2769,N_1073);
nor U5536 (N_5536,N_4781,N_2285);
nand U5537 (N_5537,N_3023,N_4381);
nor U5538 (N_5538,N_2566,N_638);
nand U5539 (N_5539,N_346,N_3568);
and U5540 (N_5540,N_712,N_1256);
or U5541 (N_5541,N_4553,N_2921);
or U5542 (N_5542,N_3603,N_3640);
or U5543 (N_5543,N_35,N_39);
nand U5544 (N_5544,N_4077,N_1343);
and U5545 (N_5545,N_3799,N_1669);
or U5546 (N_5546,N_144,N_613);
and U5547 (N_5547,N_3866,N_3335);
nor U5548 (N_5548,N_3424,N_4600);
xnor U5549 (N_5549,N_3776,N_1820);
nor U5550 (N_5550,N_2113,N_1327);
nor U5551 (N_5551,N_3347,N_171);
nor U5552 (N_5552,N_1872,N_739);
xor U5553 (N_5553,N_405,N_4787);
nor U5554 (N_5554,N_890,N_3955);
and U5555 (N_5555,N_4697,N_1082);
or U5556 (N_5556,N_3135,N_2634);
or U5557 (N_5557,N_2127,N_268);
nor U5558 (N_5558,N_1319,N_2241);
nor U5559 (N_5559,N_4134,N_364);
nor U5560 (N_5560,N_3348,N_3778);
nor U5561 (N_5561,N_2282,N_3828);
nand U5562 (N_5562,N_3375,N_623);
and U5563 (N_5563,N_481,N_4557);
nand U5564 (N_5564,N_2018,N_3604);
nand U5565 (N_5565,N_1595,N_911);
or U5566 (N_5566,N_1243,N_182);
and U5567 (N_5567,N_1379,N_619);
nand U5568 (N_5568,N_3136,N_3790);
xnor U5569 (N_5569,N_3688,N_1252);
nor U5570 (N_5570,N_3864,N_4869);
xor U5571 (N_5571,N_916,N_672);
nor U5572 (N_5572,N_500,N_1700);
nor U5573 (N_5573,N_2335,N_116);
or U5574 (N_5574,N_2172,N_1852);
nor U5575 (N_5575,N_91,N_1422);
nand U5576 (N_5576,N_110,N_4007);
and U5577 (N_5577,N_2666,N_2604);
nor U5578 (N_5578,N_4474,N_4544);
nor U5579 (N_5579,N_2679,N_2791);
and U5580 (N_5580,N_1886,N_4356);
or U5581 (N_5581,N_4759,N_1660);
nand U5582 (N_5582,N_2904,N_908);
and U5583 (N_5583,N_2557,N_1929);
xnor U5584 (N_5584,N_4949,N_115);
nor U5585 (N_5585,N_4977,N_4425);
nor U5586 (N_5586,N_4224,N_3199);
nor U5587 (N_5587,N_4316,N_3842);
nor U5588 (N_5588,N_4657,N_4015);
or U5589 (N_5589,N_3618,N_3484);
xor U5590 (N_5590,N_3512,N_2386);
nand U5591 (N_5591,N_4317,N_178);
and U5592 (N_5592,N_3821,N_2054);
or U5593 (N_5593,N_2952,N_1282);
nor U5594 (N_5594,N_1219,N_3517);
and U5595 (N_5595,N_49,N_2225);
and U5596 (N_5596,N_109,N_4767);
or U5597 (N_5597,N_3337,N_4254);
nand U5598 (N_5598,N_3020,N_994);
and U5599 (N_5599,N_1679,N_678);
or U5600 (N_5600,N_4197,N_4151);
and U5601 (N_5601,N_2471,N_839);
and U5602 (N_5602,N_4116,N_124);
or U5603 (N_5603,N_189,N_4737);
or U5604 (N_5604,N_809,N_2364);
nor U5605 (N_5605,N_1543,N_4964);
or U5606 (N_5606,N_743,N_248);
nand U5607 (N_5607,N_4856,N_27);
xnor U5608 (N_5608,N_2117,N_4570);
or U5609 (N_5609,N_4992,N_3700);
or U5610 (N_5610,N_3043,N_54);
and U5611 (N_5611,N_4558,N_3077);
and U5612 (N_5612,N_4644,N_969);
nand U5613 (N_5613,N_517,N_264);
or U5614 (N_5614,N_4372,N_1781);
or U5615 (N_5615,N_1713,N_21);
xor U5616 (N_5616,N_494,N_2897);
nor U5617 (N_5617,N_1399,N_2963);
and U5618 (N_5618,N_396,N_2549);
or U5619 (N_5619,N_4124,N_4141);
or U5620 (N_5620,N_3464,N_4329);
nor U5621 (N_5621,N_4213,N_4443);
or U5622 (N_5622,N_3814,N_4287);
nor U5623 (N_5623,N_737,N_4873);
and U5624 (N_5624,N_4301,N_1720);
and U5625 (N_5625,N_2051,N_1360);
nand U5626 (N_5626,N_3953,N_992);
nand U5627 (N_5627,N_862,N_313);
nor U5628 (N_5628,N_2959,N_4674);
nor U5629 (N_5629,N_2309,N_4304);
nand U5630 (N_5630,N_2988,N_1237);
nor U5631 (N_5631,N_3665,N_1323);
or U5632 (N_5632,N_1631,N_2511);
and U5633 (N_5633,N_802,N_3125);
nor U5634 (N_5634,N_4804,N_1823);
and U5635 (N_5635,N_419,N_2455);
xnor U5636 (N_5636,N_560,N_941);
nand U5637 (N_5637,N_1034,N_2794);
nor U5638 (N_5638,N_2953,N_1998);
and U5639 (N_5639,N_1862,N_4185);
xnor U5640 (N_5640,N_1210,N_1842);
xnor U5641 (N_5641,N_842,N_1798);
nand U5642 (N_5642,N_2828,N_2919);
and U5643 (N_5643,N_667,N_2668);
nor U5644 (N_5644,N_828,N_1228);
nor U5645 (N_5645,N_904,N_651);
nand U5646 (N_5646,N_2040,N_1901);
nand U5647 (N_5647,N_3163,N_1534);
nand U5648 (N_5648,N_401,N_512);
nand U5649 (N_5649,N_3393,N_1978);
and U5650 (N_5650,N_3531,N_4847);
and U5651 (N_5651,N_3899,N_2553);
and U5652 (N_5652,N_1078,N_507);
nand U5653 (N_5653,N_2735,N_1280);
or U5654 (N_5654,N_4286,N_3606);
nand U5655 (N_5655,N_3940,N_3837);
nand U5656 (N_5656,N_531,N_3213);
nor U5657 (N_5657,N_2507,N_4182);
nand U5658 (N_5658,N_2635,N_4095);
nand U5659 (N_5659,N_4021,N_2943);
and U5660 (N_5660,N_3056,N_321);
or U5661 (N_5661,N_4816,N_2939);
xnor U5662 (N_5662,N_1690,N_4406);
or U5663 (N_5663,N_4912,N_1456);
and U5664 (N_5664,N_411,N_1116);
and U5665 (N_5665,N_4606,N_3248);
nand U5666 (N_5666,N_2431,N_4830);
or U5667 (N_5667,N_4549,N_444);
nand U5668 (N_5668,N_2678,N_3216);
nand U5669 (N_5669,N_2506,N_792);
nor U5670 (N_5670,N_553,N_1201);
nor U5671 (N_5671,N_3861,N_2729);
and U5672 (N_5672,N_3612,N_4427);
or U5673 (N_5673,N_1326,N_2669);
and U5674 (N_5674,N_3045,N_4923);
and U5675 (N_5675,N_4632,N_3003);
and U5676 (N_5676,N_4253,N_3468);
or U5677 (N_5677,N_4942,N_3083);
xnor U5678 (N_5678,N_106,N_343);
or U5679 (N_5679,N_1145,N_2526);
nand U5680 (N_5680,N_3682,N_1509);
and U5681 (N_5681,N_4325,N_956);
nand U5682 (N_5682,N_1630,N_2617);
or U5683 (N_5683,N_3489,N_1215);
and U5684 (N_5684,N_4202,N_1602);
nand U5685 (N_5685,N_2319,N_289);
nor U5686 (N_5686,N_2197,N_1577);
nor U5687 (N_5687,N_3239,N_1254);
nand U5688 (N_5688,N_4365,N_1415);
nand U5689 (N_5689,N_2718,N_2774);
nand U5690 (N_5690,N_4416,N_3291);
or U5691 (N_5691,N_1671,N_606);
and U5692 (N_5692,N_142,N_1632);
xnor U5693 (N_5693,N_2369,N_470);
or U5694 (N_5694,N_1444,N_3738);
nand U5695 (N_5695,N_1189,N_3306);
nor U5696 (N_5696,N_4038,N_1288);
nand U5697 (N_5697,N_15,N_926);
nor U5698 (N_5698,N_2262,N_3162);
and U5699 (N_5699,N_4083,N_3882);
xor U5700 (N_5700,N_1649,N_3504);
xnor U5701 (N_5701,N_2626,N_545);
nor U5702 (N_5702,N_3903,N_456);
or U5703 (N_5703,N_3141,N_1991);
nor U5704 (N_5704,N_330,N_4962);
nand U5705 (N_5705,N_10,N_1306);
or U5706 (N_5706,N_823,N_1169);
and U5707 (N_5707,N_3292,N_2462);
nor U5708 (N_5708,N_2991,N_1499);
and U5709 (N_5709,N_13,N_1658);
and U5710 (N_5710,N_4520,N_4958);
nand U5711 (N_5711,N_2680,N_1300);
and U5712 (N_5712,N_2048,N_603);
xor U5713 (N_5713,N_1708,N_673);
nor U5714 (N_5714,N_830,N_4006);
or U5715 (N_5715,N_119,N_2804);
nor U5716 (N_5716,N_4091,N_2106);
or U5717 (N_5717,N_4233,N_549);
and U5718 (N_5718,N_1839,N_3302);
nand U5719 (N_5719,N_4509,N_4775);
or U5720 (N_5720,N_1948,N_1637);
nand U5721 (N_5721,N_3134,N_3189);
nor U5722 (N_5722,N_786,N_4732);
or U5723 (N_5723,N_1048,N_2049);
nor U5724 (N_5724,N_4180,N_965);
nor U5725 (N_5725,N_2322,N_2533);
xnor U5726 (N_5726,N_4620,N_1984);
or U5727 (N_5727,N_659,N_1791);
and U5728 (N_5728,N_986,N_4136);
and U5729 (N_5729,N_498,N_4817);
or U5730 (N_5730,N_2348,N_4453);
nand U5731 (N_5731,N_2330,N_3986);
nand U5732 (N_5732,N_3569,N_137);
or U5733 (N_5733,N_3815,N_1447);
or U5734 (N_5734,N_263,N_3129);
nand U5735 (N_5735,N_3362,N_1829);
nand U5736 (N_5736,N_3672,N_3689);
or U5737 (N_5737,N_652,N_1847);
nand U5738 (N_5738,N_3600,N_3349);
or U5739 (N_5739,N_4258,N_42);
nor U5740 (N_5740,N_1375,N_243);
and U5741 (N_5741,N_3243,N_427);
nand U5742 (N_5742,N_1743,N_2210);
or U5743 (N_5743,N_3752,N_3119);
nand U5744 (N_5744,N_2087,N_1233);
and U5745 (N_5745,N_3448,N_1865);
xor U5746 (N_5746,N_790,N_3212);
xor U5747 (N_5747,N_1203,N_1100);
nand U5748 (N_5748,N_1869,N_3005);
xnor U5749 (N_5749,N_923,N_2091);
or U5750 (N_5750,N_951,N_2625);
and U5751 (N_5751,N_1527,N_1010);
or U5752 (N_5752,N_105,N_2327);
xnor U5753 (N_5753,N_1083,N_4332);
nand U5754 (N_5754,N_3421,N_4506);
or U5755 (N_5755,N_2924,N_1356);
nor U5756 (N_5756,N_1977,N_1557);
and U5757 (N_5757,N_118,N_4252);
or U5758 (N_5758,N_4459,N_616);
and U5759 (N_5759,N_3220,N_2211);
or U5760 (N_5760,N_4952,N_4822);
nand U5761 (N_5761,N_3382,N_4954);
or U5762 (N_5762,N_865,N_1264);
xnor U5763 (N_5763,N_2474,N_1449);
and U5764 (N_5764,N_3736,N_2993);
or U5765 (N_5765,N_1774,N_2927);
or U5766 (N_5766,N_3540,N_3054);
and U5767 (N_5767,N_3094,N_4359);
xnor U5768 (N_5768,N_1544,N_4975);
xnor U5769 (N_5769,N_366,N_2072);
or U5770 (N_5770,N_4292,N_2414);
and U5771 (N_5771,N_765,N_3771);
or U5772 (N_5772,N_3608,N_4010);
nor U5773 (N_5773,N_711,N_1505);
nand U5774 (N_5774,N_2356,N_25);
and U5775 (N_5775,N_4879,N_4236);
or U5776 (N_5776,N_279,N_3132);
nor U5777 (N_5777,N_4200,N_1749);
nand U5778 (N_5778,N_356,N_4792);
or U5779 (N_5779,N_2004,N_4624);
or U5780 (N_5780,N_982,N_4186);
nor U5781 (N_5781,N_1898,N_2917);
nand U5782 (N_5782,N_4392,N_1686);
nor U5783 (N_5783,N_460,N_2423);
or U5784 (N_5784,N_3551,N_2188);
xor U5785 (N_5785,N_2610,N_4852);
xor U5786 (N_5786,N_24,N_3611);
or U5787 (N_5787,N_1909,N_4548);
nor U5788 (N_5788,N_3266,N_3434);
and U5789 (N_5789,N_3676,N_2481);
xor U5790 (N_5790,N_2281,N_254);
or U5791 (N_5791,N_1302,N_609);
nand U5792 (N_5792,N_4341,N_3018);
and U5793 (N_5793,N_4695,N_246);
nor U5794 (N_5794,N_1973,N_4824);
or U5795 (N_5795,N_756,N_4970);
nand U5796 (N_5796,N_4489,N_1517);
nand U5797 (N_5797,N_4692,N_3365);
xor U5798 (N_5798,N_920,N_3695);
and U5799 (N_5799,N_727,N_1419);
nor U5800 (N_5800,N_787,N_437);
xor U5801 (N_5801,N_3511,N_2801);
xor U5802 (N_5802,N_1503,N_3234);
or U5803 (N_5803,N_817,N_2965);
xor U5804 (N_5804,N_2025,N_4507);
xor U5805 (N_5805,N_4956,N_4994);
xnor U5806 (N_5806,N_4889,N_2721);
and U5807 (N_5807,N_3396,N_4656);
or U5808 (N_5808,N_4458,N_3064);
nor U5809 (N_5809,N_1117,N_2441);
and U5810 (N_5810,N_3112,N_538);
nand U5811 (N_5811,N_2204,N_4634);
nand U5812 (N_5812,N_376,N_2855);
nand U5813 (N_5813,N_176,N_3705);
and U5814 (N_5814,N_1890,N_3598);
and U5815 (N_5815,N_3327,N_4440);
and U5816 (N_5816,N_2659,N_4867);
or U5817 (N_5817,N_922,N_1843);
nor U5818 (N_5818,N_170,N_1606);
and U5819 (N_5819,N_3948,N_1295);
and U5820 (N_5820,N_3478,N_681);
xnor U5821 (N_5821,N_2510,N_3760);
nor U5822 (N_5822,N_4690,N_4541);
or U5823 (N_5823,N_4666,N_4834);
and U5824 (N_5824,N_2513,N_2168);
or U5825 (N_5825,N_469,N_4052);
nor U5826 (N_5826,N_1113,N_4155);
xor U5827 (N_5827,N_2682,N_1793);
or U5828 (N_5828,N_4220,N_3010);
nor U5829 (N_5829,N_3970,N_2638);
or U5830 (N_5830,N_3313,N_4621);
nand U5831 (N_5831,N_4881,N_3709);
and U5832 (N_5832,N_4383,N_3050);
xnor U5833 (N_5833,N_4322,N_3445);
nand U5834 (N_5834,N_317,N_1521);
nor U5835 (N_5835,N_4683,N_8);
or U5836 (N_5836,N_4791,N_2813);
nor U5837 (N_5837,N_4763,N_3884);
nor U5838 (N_5838,N_1670,N_793);
nor U5839 (N_5839,N_2525,N_1941);
and U5840 (N_5840,N_3507,N_2649);
nor U5841 (N_5841,N_4495,N_1191);
nor U5842 (N_5842,N_433,N_514);
nor U5843 (N_5843,N_869,N_1266);
or U5844 (N_5844,N_3848,N_996);
or U5845 (N_5845,N_64,N_4969);
nor U5846 (N_5846,N_3172,N_1589);
nand U5847 (N_5847,N_4613,N_615);
nand U5848 (N_5848,N_3658,N_2629);
xor U5849 (N_5849,N_220,N_1673);
and U5850 (N_5850,N_3316,N_1597);
and U5851 (N_5851,N_2619,N_2174);
nor U5852 (N_5852,N_3938,N_3971);
and U5853 (N_5853,N_1814,N_4514);
or U5854 (N_5854,N_3182,N_2908);
nand U5855 (N_5855,N_1151,N_2038);
nand U5856 (N_5856,N_1640,N_4826);
or U5857 (N_5857,N_2161,N_4932);
nand U5858 (N_5858,N_2612,N_3637);
xor U5859 (N_5859,N_3862,N_280);
and U5860 (N_5860,N_4654,N_1959);
nor U5861 (N_5861,N_1227,N_4594);
xor U5862 (N_5862,N_3497,N_1950);
nand U5863 (N_5863,N_2531,N_3400);
nand U5864 (N_5864,N_68,N_4769);
nand U5865 (N_5865,N_2821,N_947);
and U5866 (N_5866,N_2599,N_4663);
or U5867 (N_5867,N_4933,N_554);
xnor U5868 (N_5868,N_3998,N_1039);
or U5869 (N_5869,N_3968,N_3663);
nor U5870 (N_5870,N_3476,N_4701);
or U5871 (N_5871,N_837,N_788);
nand U5872 (N_5872,N_3363,N_4005);
nand U5873 (N_5873,N_3333,N_4436);
nor U5874 (N_5874,N_3190,N_4163);
nor U5875 (N_5875,N_1,N_1672);
nor U5876 (N_5876,N_4516,N_4315);
or U5877 (N_5877,N_3939,N_1428);
and U5878 (N_5878,N_4909,N_1969);
nand U5879 (N_5879,N_4950,N_1418);
nand U5880 (N_5880,N_1845,N_1410);
or U5881 (N_5881,N_499,N_4101);
or U5882 (N_5882,N_2938,N_2430);
nand U5883 (N_5883,N_876,N_2037);
nand U5884 (N_5884,N_1889,N_4884);
xnor U5885 (N_5885,N_3756,N_3208);
and U5886 (N_5886,N_3079,N_3004);
nor U5887 (N_5887,N_1402,N_4208);
or U5888 (N_5888,N_4929,N_2400);
nand U5889 (N_5889,N_4492,N_262);
nand U5890 (N_5890,N_2676,N_1420);
nor U5891 (N_5891,N_2250,N_861);
nor U5892 (N_5892,N_1564,N_2137);
nor U5893 (N_5893,N_1371,N_605);
and U5894 (N_5894,N_1109,N_3338);
and U5895 (N_5895,N_2377,N_3029);
nand U5896 (N_5896,N_1783,N_1344);
xnor U5897 (N_5897,N_2665,N_2320);
nor U5898 (N_5898,N_2163,N_1338);
or U5899 (N_5899,N_136,N_1138);
nand U5900 (N_5900,N_1695,N_1235);
and U5901 (N_5901,N_764,N_1412);
or U5902 (N_5902,N_34,N_3692);
nand U5903 (N_5903,N_108,N_1007);
nor U5904 (N_5904,N_273,N_4953);
and U5905 (N_5905,N_4094,N_845);
or U5906 (N_5906,N_2624,N_781);
or U5907 (N_5907,N_4984,N_723);
or U5908 (N_5908,N_833,N_3233);
nor U5909 (N_5909,N_1522,N_4810);
or U5910 (N_5910,N_1476,N_2173);
nand U5911 (N_5911,N_3453,N_4441);
xor U5912 (N_5912,N_2491,N_738);
and U5913 (N_5913,N_4028,N_584);
and U5914 (N_5914,N_4498,N_974);
or U5915 (N_5915,N_2568,N_320);
and U5916 (N_5916,N_2731,N_2411);
xor U5917 (N_5917,N_3697,N_3329);
nor U5918 (N_5918,N_4351,N_4271);
or U5919 (N_5919,N_1454,N_1994);
or U5920 (N_5920,N_4080,N_477);
nor U5921 (N_5921,N_2562,N_2832);
or U5922 (N_5922,N_1489,N_1178);
or U5923 (N_5923,N_3287,N_2763);
nand U5924 (N_5924,N_2212,N_3235);
and U5925 (N_5925,N_1538,N_4448);
and U5926 (N_5926,N_2983,N_1008);
or U5927 (N_5927,N_3909,N_4338);
or U5928 (N_5928,N_2591,N_4639);
nand U5929 (N_5929,N_1756,N_701);
and U5930 (N_5930,N_3227,N_2273);
nor U5931 (N_5931,N_1285,N_3294);
nor U5932 (N_5932,N_3193,N_1697);
and U5933 (N_5933,N_2071,N_1232);
nand U5934 (N_5934,N_870,N_2565);
or U5935 (N_5935,N_3260,N_4571);
xor U5936 (N_5936,N_971,N_484);
nor U5937 (N_5937,N_4840,N_2189);
nor U5938 (N_5938,N_375,N_579);
nor U5939 (N_5939,N_2532,N_3643);
nand U5940 (N_5940,N_3456,N_3703);
xnor U5941 (N_5941,N_2253,N_1752);
or U5942 (N_5942,N_1394,N_305);
or U5943 (N_5943,N_3906,N_1565);
and U5944 (N_5944,N_1619,N_3889);
nor U5945 (N_5945,N_2909,N_520);
nor U5946 (N_5946,N_1198,N_50);
xnor U5947 (N_5947,N_1834,N_726);
nor U5948 (N_5948,N_740,N_4353);
nor U5949 (N_5949,N_1728,N_1830);
or U5950 (N_5950,N_3386,N_754);
xnor U5951 (N_5951,N_4580,N_1213);
nor U5952 (N_5952,N_2227,N_4746);
or U5953 (N_5953,N_2198,N_3121);
or U5954 (N_5954,N_120,N_2482);
or U5955 (N_5955,N_852,N_4054);
nor U5956 (N_5956,N_4046,N_1907);
nand U5957 (N_5957,N_352,N_4324);
nand U5958 (N_5958,N_267,N_1277);
nor U5959 (N_5959,N_3558,N_1395);
nand U5960 (N_5960,N_3027,N_36);
nand U5961 (N_5961,N_252,N_213);
nor U5962 (N_5962,N_1363,N_660);
and U5963 (N_5963,N_3690,N_1981);
and U5964 (N_5964,N_1967,N_2671);
nor U5965 (N_5965,N_3601,N_1739);
nor U5966 (N_5966,N_1854,N_1644);
xnor U5967 (N_5967,N_4718,N_1677);
nand U5968 (N_5968,N_1225,N_3516);
nand U5969 (N_5969,N_4374,N_3308);
and U5970 (N_5970,N_1060,N_4118);
and U5971 (N_5971,N_755,N_314);
nor U5972 (N_5972,N_769,N_200);
nand U5973 (N_5973,N_1154,N_2077);
and U5974 (N_5974,N_1377,N_999);
nor U5975 (N_5975,N_1106,N_1887);
nand U5976 (N_5976,N_3444,N_879);
and U5977 (N_5977,N_3143,N_557);
nor U5978 (N_5978,N_4583,N_112);
and U5979 (N_5979,N_4477,N_3990);
nor U5980 (N_5980,N_4234,N_1908);
nand U5981 (N_5981,N_580,N_550);
nand U5982 (N_5982,N_3293,N_2892);
and U5983 (N_5983,N_863,N_780);
or U5984 (N_5984,N_3052,N_4423);
nor U5985 (N_5985,N_4394,N_1382);
and U5986 (N_5986,N_1664,N_1580);
nand U5987 (N_5987,N_2152,N_4106);
nor U5988 (N_5988,N_1486,N_2742);
nor U5989 (N_5989,N_4035,N_2358);
or U5990 (N_5990,N_2727,N_186);
nor U5991 (N_5991,N_4187,N_155);
nand U5992 (N_5992,N_1119,N_3716);
and U5993 (N_5993,N_361,N_312);
nor U5994 (N_5994,N_1293,N_3720);
or U5995 (N_5995,N_1229,N_4829);
and U5996 (N_5996,N_2826,N_4671);
and U5997 (N_5997,N_4026,N_3397);
or U5998 (N_5998,N_4521,N_1335);
or U5999 (N_5999,N_4637,N_2913);
or U6000 (N_6000,N_1855,N_166);
and U6001 (N_6001,N_4704,N_1848);
nor U6002 (N_6002,N_4947,N_94);
and U6003 (N_6003,N_688,N_2308);
and U6004 (N_6004,N_4117,N_2219);
xor U6005 (N_6005,N_3693,N_919);
nand U6006 (N_6006,N_1938,N_392);
nor U6007 (N_6007,N_682,N_973);
nand U6008 (N_6008,N_2728,N_4398);
nor U6009 (N_6009,N_2246,N_1615);
nand U6010 (N_6010,N_3200,N_1018);
nor U6011 (N_6011,N_2741,N_721);
and U6012 (N_6012,N_2451,N_3947);
and U6013 (N_6013,N_1813,N_513);
xnor U6014 (N_6014,N_4587,N_310);
nand U6015 (N_6015,N_1217,N_2691);
nor U6016 (N_6016,N_2221,N_2490);
or U6017 (N_6017,N_2854,N_2752);
nor U6018 (N_6018,N_1031,N_3176);
nand U6019 (N_6019,N_2296,N_3623);
or U6020 (N_6020,N_1831,N_3279);
nor U6021 (N_6021,N_3800,N_3571);
xor U6022 (N_6022,N_1801,N_1510);
xnor U6023 (N_6023,N_1729,N_3168);
nand U6024 (N_6024,N_607,N_2694);
or U6025 (N_6025,N_438,N_896);
or U6026 (N_6026,N_379,N_1214);
nand U6027 (N_6027,N_446,N_4766);
nand U6028 (N_6028,N_4399,N_910);
or U6029 (N_6029,N_373,N_3987);
nor U6030 (N_6030,N_4485,N_249);
nor U6031 (N_6031,N_1140,N_2772);
or U6032 (N_6032,N_2413,N_483);
or U6033 (N_6033,N_1975,N_2834);
and U6034 (N_6034,N_4161,N_650);
nand U6035 (N_6035,N_2224,N_190);
nand U6036 (N_6036,N_4442,N_372);
nor U6037 (N_6037,N_4377,N_883);
nand U6038 (N_6038,N_3171,N_1222);
nand U6039 (N_6039,N_4125,N_2843);
nor U6040 (N_6040,N_2217,N_3452);
nor U6041 (N_6041,N_1952,N_4555);
nand U6042 (N_6042,N_1762,N_2820);
nor U6043 (N_6043,N_1053,N_859);
and U6044 (N_6044,N_4795,N_3742);
nand U6045 (N_6045,N_2065,N_2080);
nor U6046 (N_6046,N_1709,N_1913);
and U6047 (N_6047,N_2466,N_125);
nand U6048 (N_6048,N_3031,N_349);
nand U6049 (N_6049,N_692,N_1494);
nand U6050 (N_6050,N_2483,N_3874);
or U6051 (N_6051,N_1207,N_2145);
nand U6052 (N_6052,N_1016,N_1396);
nand U6053 (N_6053,N_4597,N_3069);
nand U6054 (N_6054,N_1656,N_3195);
nor U6055 (N_6055,N_28,N_3973);
and U6056 (N_6056,N_505,N_2840);
or U6057 (N_6057,N_2600,N_3262);
nand U6058 (N_6058,N_2010,N_2318);
nor U6059 (N_6059,N_1223,N_4604);
and U6060 (N_6060,N_4488,N_1868);
nand U6061 (N_6061,N_4573,N_2886);
nor U6062 (N_6062,N_3191,N_3976);
nand U6063 (N_6063,N_1005,N_2035);
nor U6064 (N_6064,N_3671,N_1185);
or U6065 (N_6065,N_2951,N_284);
and U6066 (N_6066,N_311,N_3891);
nand U6067 (N_6067,N_1218,N_2797);
nor U6068 (N_6068,N_2720,N_4736);
or U6069 (N_6069,N_1349,N_2108);
xor U6070 (N_6070,N_4530,N_335);
nor U6071 (N_6071,N_4256,N_1287);
nand U6072 (N_6072,N_1188,N_4496);
xor U6073 (N_6073,N_4913,N_4849);
or U6074 (N_6074,N_3878,N_3832);
nand U6075 (N_6075,N_3630,N_1824);
nor U6076 (N_6076,N_4310,N_2590);
nand U6077 (N_6077,N_2688,N_4681);
or U6078 (N_6078,N_3783,N_1378);
and U6079 (N_6079,N_4040,N_2695);
and U6080 (N_6080,N_1352,N_1464);
nand U6081 (N_6081,N_309,N_1089);
and U6082 (N_6082,N_1927,N_1723);
nand U6083 (N_6083,N_2961,N_877);
nor U6084 (N_6084,N_1297,N_4561);
nor U6085 (N_6085,N_1481,N_1439);
xnor U6086 (N_6086,N_4067,N_1400);
nand U6087 (N_6087,N_4154,N_1275);
xnor U6088 (N_6088,N_812,N_3721);
nor U6089 (N_6089,N_2085,N_2715);
or U6090 (N_6090,N_2540,N_4217);
nor U6091 (N_6091,N_1221,N_261);
and U6092 (N_6092,N_2887,N_4741);
and U6093 (N_6093,N_783,N_4285);
and U6094 (N_6094,N_1158,N_1162);
and U6095 (N_6095,N_1815,N_2352);
nand U6096 (N_6096,N_1348,N_1870);
nor U6097 (N_6097,N_2581,N_2190);
or U6098 (N_6098,N_991,N_3389);
nand U6099 (N_6099,N_1600,N_4060);
or U6100 (N_6100,N_4264,N_4762);
or U6101 (N_6101,N_2675,N_1860);
and U6102 (N_6102,N_3983,N_3999);
and U6103 (N_6103,N_3026,N_2315);
and U6104 (N_6104,N_984,N_4603);
nand U6105 (N_6105,N_3614,N_1850);
or U6106 (N_6106,N_2379,N_3679);
nor U6107 (N_6107,N_1496,N_292);
nand U6108 (N_6108,N_2815,N_1807);
and U6109 (N_6109,N_3438,N_3650);
or U6110 (N_6110,N_1520,N_3763);
nor U6111 (N_6111,N_596,N_4159);
nor U6112 (N_6112,N_3596,N_782);
nor U6113 (N_6113,N_2788,N_420);
and U6114 (N_6114,N_2104,N_101);
nor U6115 (N_6115,N_2879,N_157);
and U6116 (N_6116,N_909,N_4241);
or U6117 (N_6117,N_1571,N_970);
nor U6118 (N_6118,N_2893,N_351);
or U6119 (N_6119,N_4371,N_4935);
and U6120 (N_6120,N_4169,N_1507);
nor U6121 (N_6121,N_4042,N_562);
or U6122 (N_6122,N_2633,N_3425);
nand U6123 (N_6123,N_4988,N_3037);
nand U6124 (N_6124,N_1554,N_2770);
nor U6125 (N_6125,N_3634,N_3952);
nor U6126 (N_6126,N_2006,N_4874);
or U6127 (N_6127,N_1064,N_1805);
nor U6128 (N_6128,N_6,N_2155);
nand U6129 (N_6129,N_1857,N_4729);
or U6130 (N_6130,N_3797,N_4168);
nand U6131 (N_6131,N_4866,N_1332);
nand U6132 (N_6132,N_4284,N_2245);
and U6133 (N_6133,N_3115,N_1069);
xnor U6134 (N_6134,N_308,N_2433);
nand U6135 (N_6135,N_636,N_4404);
xnor U6136 (N_6136,N_230,N_3461);
nor U6137 (N_6137,N_4482,N_2724);
xnor U6138 (N_6138,N_687,N_2830);
xnor U6139 (N_6139,N_634,N_2523);
or U6140 (N_6140,N_1897,N_2426);
or U6141 (N_6141,N_1401,N_2073);
or U6142 (N_6142,N_4525,N_2136);
nor U6143 (N_6143,N_3441,N_1776);
xor U6144 (N_6144,N_600,N_4362);
nor U6145 (N_6145,N_2181,N_1167);
nand U6146 (N_6146,N_2857,N_3869);
nand U6147 (N_6147,N_1731,N_3155);
or U6148 (N_6148,N_1715,N_1849);
nor U6149 (N_6149,N_4651,N_3673);
and U6150 (N_6150,N_2672,N_2294);
nor U6151 (N_6151,N_4642,N_215);
nand U6152 (N_6152,N_3401,N_4647);
and U6153 (N_6153,N_1960,N_1049);
nor U6154 (N_6154,N_3564,N_4127);
xnor U6155 (N_6155,N_2034,N_3466);
nand U6156 (N_6156,N_72,N_2086);
nor U6157 (N_6157,N_203,N_4113);
nand U6158 (N_6158,N_4308,N_2910);
nor U6159 (N_6159,N_4702,N_4244);
nor U6160 (N_6160,N_4773,N_611);
nand U6161 (N_6161,N_1682,N_2615);
and U6162 (N_6162,N_1825,N_1004);
nor U6163 (N_6163,N_4793,N_3009);
nand U6164 (N_6164,N_4179,N_840);
nor U6165 (N_6165,N_150,N_3503);
or U6166 (N_6166,N_2631,N_2572);
and U6167 (N_6167,N_2898,N_429);
nand U6168 (N_6168,N_1427,N_1607);
nor U6169 (N_6169,N_3794,N_223);
nand U6170 (N_6170,N_4064,N_1289);
and U6171 (N_6171,N_3656,N_389);
nand U6172 (N_6172,N_3013,N_2192);
or U6173 (N_6173,N_1090,N_71);
nor U6174 (N_6174,N_131,N_3795);
xnor U6175 (N_6175,N_4105,N_632);
nor U6176 (N_6176,N_1092,N_4968);
nand U6177 (N_6177,N_3326,N_3272);
xnor U6178 (N_6178,N_2942,N_977);
or U6179 (N_6179,N_872,N_3514);
nor U6180 (N_6180,N_244,N_275);
nor U6181 (N_6181,N_3539,N_1143);
or U6182 (N_6182,N_4883,N_4652);
and U6183 (N_6183,N_4999,N_4178);
nand U6184 (N_6184,N_831,N_2337);
or U6185 (N_6185,N_4870,N_1125);
or U6186 (N_6186,N_3934,N_204);
nor U6187 (N_6187,N_4770,N_2169);
or U6188 (N_6188,N_3574,N_2436);
or U6189 (N_6189,N_1393,N_1634);
and U6190 (N_6190,N_3104,N_187);
nor U6191 (N_6191,N_2045,N_627);
nor U6192 (N_6192,N_2627,N_4533);
nand U6193 (N_6193,N_318,N_4062);
or U6194 (N_6194,N_4980,N_4451);
nand U6195 (N_6195,N_43,N_2122);
nand U6196 (N_6196,N_2867,N_3460);
nand U6197 (N_6197,N_568,N_2267);
xor U6198 (N_6198,N_4535,N_1687);
and U6199 (N_6199,N_1478,N_4661);
or U6200 (N_6200,N_1738,N_3368);
nand U6201 (N_6201,N_1468,N_4730);
and U6202 (N_6202,N_2119,N_3748);
nor U6203 (N_6203,N_4149,N_3683);
or U6204 (N_6204,N_4720,N_3639);
xor U6205 (N_6205,N_750,N_3879);
and U6206 (N_6206,N_878,N_1350);
xnor U6207 (N_6207,N_4240,N_4449);
nand U6208 (N_6208,N_4900,N_140);
or U6209 (N_6209,N_3378,N_2470);
or U6210 (N_6210,N_1680,N_4564);
and U6211 (N_6211,N_2996,N_2251);
or U6212 (N_6212,N_3357,N_276);
nor U6213 (N_6213,N_2895,N_530);
and U6214 (N_6214,N_3749,N_2084);
nor U6215 (N_6215,N_3959,N_591);
xnor U6216 (N_6216,N_2670,N_141);
nand U6217 (N_6217,N_198,N_3525);
xnor U6218 (N_6218,N_4493,N_3853);
nor U6219 (N_6219,N_815,N_824);
and U6220 (N_6220,N_1965,N_4018);
and U6221 (N_6221,N_589,N_226);
or U6222 (N_6222,N_194,N_914);
and U6223 (N_6223,N_3782,N_2132);
or U6224 (N_6224,N_2193,N_4131);
or U6225 (N_6225,N_1668,N_162);
or U6226 (N_6226,N_592,N_983);
or U6227 (N_6227,N_3184,N_3857);
nor U6228 (N_6228,N_3813,N_3746);
and U6229 (N_6229,N_4255,N_4457);
or U6230 (N_6230,N_3936,N_931);
or U6231 (N_6231,N_4476,N_3107);
nand U6232 (N_6232,N_307,N_3993);
and U6233 (N_6233,N_4450,N_93);
or U6234 (N_6234,N_3714,N_3537);
nand U6235 (N_6235,N_5,N_1730);
xnor U6236 (N_6236,N_944,N_3967);
or U6237 (N_6237,N_370,N_3459);
nor U6238 (N_6238,N_4700,N_745);
nor U6239 (N_6239,N_4976,N_3865);
nand U6240 (N_6240,N_2355,N_3833);
or U6241 (N_6241,N_1617,N_4221);
nand U6242 (N_6242,N_3592,N_4166);
and U6243 (N_6243,N_2036,N_357);
nor U6244 (N_6244,N_3164,N_3863);
nand U6245 (N_6245,N_622,N_1878);
nor U6246 (N_6246,N_1620,N_1461);
or U6247 (N_6247,N_2802,N_3607);
nand U6248 (N_6248,N_1261,N_2710);
or U6249 (N_6249,N_3253,N_3082);
xor U6250 (N_6250,N_1307,N_195);
xnor U6251 (N_6251,N_4352,N_4504);
nand U6252 (N_6252,N_1910,N_3038);
nand U6253 (N_6253,N_2881,N_4369);
and U6254 (N_6254,N_1009,N_1906);
xor U6255 (N_6255,N_2517,N_2240);
and U6256 (N_6256,N_3488,N_3725);
nand U6257 (N_6257,N_4605,N_2527);
nor U6258 (N_6258,N_4665,N_1482);
or U6259 (N_6259,N_1453,N_129);
and U6260 (N_6260,N_266,N_987);
and U6261 (N_6261,N_1315,N_4051);
or U6262 (N_6262,N_3250,N_3423);
nand U6263 (N_6263,N_3430,N_2616);
and U6264 (N_6264,N_4397,N_864);
nor U6265 (N_6265,N_2740,N_4194);
and U6266 (N_6266,N_3826,N_1012);
nor U6267 (N_6267,N_4854,N_4575);
nor U6268 (N_6268,N_1568,N_2883);
nor U6269 (N_6269,N_2719,N_1905);
nand U6270 (N_6270,N_4722,N_844);
nor U6271 (N_6271,N_1314,N_3625);
or U6272 (N_6272,N_671,N_4685);
or U6273 (N_6273,N_3768,N_2972);
nand U6274 (N_6274,N_3249,N_4808);
nand U6275 (N_6275,N_4893,N_4354);
and U6276 (N_6276,N_2884,N_2199);
nand U6277 (N_6277,N_4270,N_1014);
or U6278 (N_6278,N_4393,N_4422);
or U6279 (N_6279,N_2803,N_4152);
or U6280 (N_6280,N_741,N_694);
xnor U6281 (N_6281,N_37,N_4201);
or U6282 (N_6282,N_3624,N_4430);
nand U6283 (N_6283,N_716,N_1586);
nor U6284 (N_6284,N_3664,N_2044);
and U6285 (N_6285,N_2954,N_2124);
or U6286 (N_6286,N_286,N_2743);
nor U6287 (N_6287,N_1284,N_3067);
or U6288 (N_6288,N_2149,N_4668);
nand U6289 (N_6289,N_2476,N_1599);
nand U6290 (N_6290,N_97,N_2393);
and U6291 (N_6291,N_4502,N_1755);
or U6292 (N_6292,N_2391,N_1123);
and U6293 (N_6293,N_410,N_3433);
or U6294 (N_6294,N_635,N_2215);
nand U6295 (N_6295,N_4114,N_4109);
nand U6296 (N_6296,N_2416,N_2636);
nand U6297 (N_6297,N_1576,N_322);
nand U6298 (N_6298,N_4845,N_4298);
nor U6299 (N_6299,N_3859,N_4858);
or U6300 (N_6300,N_4023,N_532);
or U6301 (N_6301,N_3156,N_3263);
nand U6302 (N_6302,N_4278,N_4572);
or U6303 (N_6303,N_1269,N_4198);
or U6304 (N_6304,N_3699,N_3792);
nand U6305 (N_6305,N_2329,N_3101);
or U6306 (N_6306,N_4190,N_3194);
and U6307 (N_6307,N_1933,N_3341);
nor U6308 (N_6308,N_1072,N_2800);
nand U6309 (N_6309,N_3809,N_902);
nor U6310 (N_6310,N_2844,N_4014);
xor U6311 (N_6311,N_4524,N_3166);
or U6312 (N_6312,N_3305,N_1681);
and U6313 (N_6313,N_2584,N_4139);
or U6314 (N_6314,N_3463,N_3647);
or U6315 (N_6315,N_3145,N_4478);
and U6316 (N_6316,N_2502,N_2862);
nand U6317 (N_6317,N_598,N_3573);
or U6318 (N_6318,N_1647,N_4242);
or U6319 (N_6319,N_604,N_2150);
nand U6320 (N_6320,N_368,N_3523);
nor U6321 (N_6321,N_3065,N_493);
or U6322 (N_6322,N_440,N_1079);
or U6323 (N_6323,N_689,N_2810);
nor U6324 (N_6324,N_2157,N_1211);
nor U6325 (N_6325,N_92,N_2548);
xor U6326 (N_6326,N_1074,N_402);
and U6327 (N_6327,N_3204,N_4367);
nor U6328 (N_6328,N_4921,N_686);
or U6329 (N_6329,N_1388,N_2784);
and U6330 (N_6330,N_4908,N_221);
or U6331 (N_6331,N_4877,N_506);
or U6332 (N_6332,N_2485,N_1985);
and U6333 (N_6333,N_2141,N_2807);
or U6334 (N_6334,N_1524,N_3553);
nor U6335 (N_6335,N_4547,N_1716);
nor U6336 (N_6336,N_860,N_3351);
xnor U6337 (N_6337,N_4160,N_1171);
and U6338 (N_6338,N_3961,N_3949);
nor U6339 (N_6339,N_751,N_3589);
nor U6340 (N_6340,N_47,N_2618);
and U6341 (N_6341,N_214,N_2747);
nand U6342 (N_6342,N_608,N_4966);
nand U6343 (N_6343,N_612,N_630);
xnor U6344 (N_6344,N_1777,N_1986);
and U6345 (N_6345,N_2350,N_4337);
and U6346 (N_6346,N_3230,N_3493);
nor U6347 (N_6347,N_4331,N_3850);
nor U6348 (N_6348,N_1362,N_3282);
nand U6349 (N_6349,N_1685,N_455);
nand U6350 (N_6350,N_2164,N_4566);
and U6351 (N_6351,N_3494,N_1759);
xnor U6352 (N_6352,N_16,N_3480);
or U6353 (N_6353,N_3593,N_1809);
xnor U6354 (N_6354,N_1103,N_2012);
nor U6355 (N_6355,N_2911,N_866);
nor U6356 (N_6356,N_4138,N_4102);
and U6357 (N_6357,N_1945,N_4072);
and U6358 (N_6358,N_4090,N_4839);
or U6359 (N_6359,N_4274,N_1077);
nor U6360 (N_6360,N_868,N_1526);
xor U6361 (N_6361,N_2111,N_3995);
and U6362 (N_6362,N_4465,N_912);
or U6363 (N_6363,N_906,N_2574);
nand U6364 (N_6364,N_1958,N_1790);
nor U6365 (N_6365,N_2808,N_3149);
nor U6366 (N_6366,N_3563,N_2901);
and U6367 (N_6367,N_1054,N_4986);
xnor U6368 (N_6368,N_4348,N_3996);
nand U6369 (N_6369,N_237,N_4470);
xnor U6370 (N_6370,N_3412,N_2773);
and U6371 (N_6371,N_2453,N_1675);
and U6372 (N_6372,N_2333,N_3769);
or U6373 (N_6373,N_324,N_4111);
and U6374 (N_6374,N_1558,N_4357);
or U6375 (N_6375,N_3502,N_3988);
nor U6376 (N_6376,N_508,N_4943);
nor U6377 (N_6377,N_1513,N_1922);
nor U6378 (N_6378,N_4142,N_1884);
nor U6379 (N_6379,N_4735,N_4560);
and U6380 (N_6380,N_891,N_4410);
nor U6381 (N_6381,N_345,N_3917);
nor U6382 (N_6382,N_1202,N_4123);
or U6383 (N_6383,N_744,N_412);
nor U6384 (N_6384,N_3371,N_1152);
or U6385 (N_6385,N_2512,N_3161);
nor U6386 (N_6386,N_3588,N_259);
nor U6387 (N_6387,N_895,N_1346);
or U6388 (N_6388,N_4013,N_621);
and U6389 (N_6389,N_2642,N_4079);
nor U6390 (N_6390,N_2768,N_2814);
nor U6391 (N_6391,N_3167,N_421);
nor U6392 (N_6392,N_4924,N_4126);
nor U6393 (N_6393,N_2175,N_2796);
nand U6394 (N_6394,N_1135,N_2836);
or U6395 (N_6395,N_4385,N_3035);
nor U6396 (N_6396,N_2955,N_811);
or U6397 (N_6397,N_3751,N_3395);
nor U6398 (N_6398,N_582,N_2918);
nand U6399 (N_6399,N_3426,N_1070);
nand U6400 (N_6400,N_4694,N_1433);
and U6401 (N_6401,N_4939,N_725);
or U6402 (N_6402,N_3829,N_1094);
nor U6403 (N_6403,N_4313,N_1050);
nor U6404 (N_6404,N_952,N_2982);
nand U6405 (N_6405,N_1220,N_819);
nor U6406 (N_6406,N_3345,N_135);
nor U6407 (N_6407,N_742,N_680);
nor U6408 (N_6408,N_4267,N_978);
nor U6409 (N_6409,N_3924,N_2448);
or U6410 (N_6410,N_581,N_2940);
and U6411 (N_6411,N_2332,N_2288);
nand U6412 (N_6412,N_2313,N_86);
nand U6413 (N_6413,N_67,N_677);
nand U6414 (N_6414,N_4417,N_4903);
nor U6415 (N_6415,N_2420,N_1455);
nand U6416 (N_6416,N_3576,N_1942);
nand U6417 (N_6417,N_803,N_2166);
or U6418 (N_6418,N_4664,N_2074);
or U6419 (N_6419,N_96,N_1506);
nor U6420 (N_6420,N_2542,N_1924);
and U6421 (N_6421,N_1902,N_4246);
or U6422 (N_6422,N_2776,N_4318);
or U6423 (N_6423,N_1546,N_2521);
or U6424 (N_6424,N_2259,N_1963);
or U6425 (N_6425,N_4920,N_2730);
and U6426 (N_6426,N_4931,N_704);
nand U6427 (N_6427,N_2070,N_4065);
or U6428 (N_6428,N_1124,N_3684);
nor U6429 (N_6429,N_760,N_4305);
or U6430 (N_6430,N_4527,N_4165);
or U6431 (N_6431,N_586,N_1635);
and U6432 (N_6432,N_1424,N_1132);
xor U6433 (N_6433,N_2402,N_53);
and U6434 (N_6434,N_3508,N_2095);
nor U6435 (N_6435,N_3429,N_3046);
nor U6436 (N_6436,N_2494,N_1471);
xor U6437 (N_6437,N_2907,N_4894);
or U6438 (N_6438,N_575,N_3807);
xor U6439 (N_6439,N_3228,N_2585);
or U6440 (N_6440,N_950,N_3538);
or U6441 (N_6441,N_2286,N_4076);
xnor U6442 (N_6442,N_4122,N_3332);
nand U6443 (N_6443,N_78,N_4245);
and U6444 (N_6444,N_1206,N_885);
xor U6445 (N_6445,N_4670,N_2125);
nor U6446 (N_6446,N_3130,N_1194);
nor U6447 (N_6447,N_2899,N_272);
and U6448 (N_6448,N_2977,N_354);
nor U6449 (N_6449,N_2650,N_4460);
nand U6450 (N_6450,N_4868,N_3728);
xnor U6451 (N_6451,N_3615,N_729);
nor U6452 (N_6452,N_2950,N_2321);
nor U6453 (N_6453,N_1168,N_3219);
and U6454 (N_6454,N_3675,N_945);
nor U6455 (N_6455,N_656,N_26);
and U6456 (N_6456,N_4996,N_449);
nor U6457 (N_6457,N_2989,N_3277);
and U6458 (N_6458,N_1504,N_84);
nand U6459 (N_6459,N_889,N_1181);
and U6460 (N_6460,N_1717,N_2856);
or U6461 (N_6461,N_1081,N_390);
nand U6462 (N_6462,N_2347,N_536);
or U6463 (N_6463,N_31,N_4783);
or U6464 (N_6464,N_1085,N_1013);
or U6465 (N_6465,N_4501,N_2027);
nor U6466 (N_6466,N_3930,N_2203);
and U6467 (N_6467,N_4918,N_1939);
nor U6468 (N_6468,N_3022,N_3084);
nor U6469 (N_6469,N_2278,N_2674);
or U6470 (N_6470,N_816,N_3729);
nand U6471 (N_6471,N_1448,N_1804);
or U6472 (N_6472,N_1550,N_1157);
nor U6473 (N_6473,N_1683,N_2029);
nor U6474 (N_6474,N_2520,N_2645);
xor U6475 (N_6475,N_4311,N_1309);
nand U6476 (N_6476,N_4345,N_2992);
xnor U6477 (N_6477,N_3286,N_2129);
or U6478 (N_6478,N_2780,N_1584);
or U6479 (N_6479,N_2849,N_3870);
nor U6480 (N_6480,N_2354,N_3957);
and U6481 (N_6481,N_1035,N_4257);
or U6482 (N_6482,N_3740,N_1028);
and U6483 (N_6483,N_2283,N_758);
or U6484 (N_6484,N_1245,N_4402);
nor U6485 (N_6485,N_2311,N_4872);
or U6486 (N_6486,N_4282,N_2699);
and U6487 (N_6487,N_4590,N_713);
nor U6488 (N_6488,N_4529,N_4409);
and U6489 (N_6489,N_3852,N_2536);
nor U6490 (N_6490,N_2648,N_95);
and U6491 (N_6491,N_4444,N_1006);
nor U6492 (N_6492,N_3,N_3898);
or U6493 (N_6493,N_2020,N_4280);
and U6494 (N_6494,N_2412,N_391);
or U6495 (N_6495,N_1112,N_4658);
nand U6496 (N_6496,N_2872,N_3068);
nor U6497 (N_6497,N_217,N_172);
nor U6498 (N_6498,N_2505,N_855);
nand U6499 (N_6499,N_1916,N_662);
nand U6500 (N_6500,N_540,N_551);
xor U6501 (N_6501,N_4272,N_2360);
or U6502 (N_6502,N_2378,N_1061);
nor U6503 (N_6503,N_1097,N_699);
nor U6504 (N_6504,N_181,N_3106);
nand U6505 (N_6505,N_724,N_2766);
and U6506 (N_6506,N_4433,N_4229);
nor U6507 (N_6507,N_3745,N_1351);
or U6508 (N_6508,N_733,N_1573);
or U6509 (N_6509,N_4585,N_2948);
xor U6510 (N_6510,N_2307,N_3097);
nand U6511 (N_6511,N_297,N_4667);
and U6512 (N_6512,N_3977,N_3232);
nand U6513 (N_6513,N_1802,N_4027);
nand U6514 (N_6514,N_3773,N_4715);
nor U6515 (N_6515,N_156,N_893);
and U6516 (N_6516,N_1989,N_1566);
nor U6517 (N_6517,N_3014,N_854);
or U6518 (N_6518,N_48,N_3352);
xnor U6519 (N_6519,N_3385,N_2052);
or U6520 (N_6520,N_2275,N_4790);
xnor U6521 (N_6521,N_4293,N_1273);
or U6522 (N_6522,N_4789,N_4755);
or U6523 (N_6523,N_1102,N_2);
nor U6524 (N_6524,N_1895,N_1260);
and U6525 (N_6525,N_2863,N_4891);
xor U6526 (N_6526,N_3528,N_1212);
and U6527 (N_6527,N_3295,N_1819);
nand U6528 (N_6528,N_4850,N_2703);
or U6529 (N_6529,N_3450,N_4069);
nand U6530 (N_6530,N_3109,N_2998);
or U6531 (N_6531,N_3229,N_3039);
and U6532 (N_6532,N_3590,N_4439);
or U6533 (N_6533,N_3214,N_4756);
or U6534 (N_6534,N_1528,N_211);
nor U6535 (N_6535,N_4650,N_2597);
nor U6536 (N_6536,N_2979,N_1249);
and U6537 (N_6537,N_1236,N_4751);
nor U6538 (N_6538,N_4437,N_2487);
and U6539 (N_6539,N_2274,N_491);
xor U6540 (N_6540,N_1095,N_1785);
and U6541 (N_6541,N_3619,N_4199);
and U6542 (N_6542,N_981,N_4653);
nor U6543 (N_6543,N_4979,N_18);
nor U6544 (N_6544,N_3509,N_4368);
nor U6545 (N_6545,N_2444,N_1020);
and U6546 (N_6546,N_3522,N_2469);
nand U6547 (N_6547,N_2702,N_2056);
or U6548 (N_6548,N_3057,N_3399);
nand U6549 (N_6549,N_829,N_2133);
or U6550 (N_6550,N_2043,N_2284);
nor U6551 (N_6551,N_1108,N_1150);
xor U6552 (N_6552,N_567,N_2479);
or U6553 (N_6553,N_1751,N_4948);
or U6554 (N_6554,N_4283,N_2147);
nand U6555 (N_6555,N_646,N_3380);
or U6556 (N_6556,N_4627,N_3314);
nor U6557 (N_6557,N_1397,N_1779);
nor U6558 (N_6558,N_4946,N_4312);
and U6559 (N_6559,N_1111,N_2218);
or U6560 (N_6560,N_1590,N_3733);
and U6561 (N_6561,N_928,N_344);
xor U6562 (N_6562,N_3403,N_3687);
or U6563 (N_6563,N_1336,N_2248);
and U6564 (N_6564,N_2381,N_2380);
and U6565 (N_6565,N_4820,N_4631);
or U6566 (N_6566,N_4107,N_1894);
and U6567 (N_6567,N_3259,N_2555);
nor U6568 (N_6568,N_4708,N_1710);
nor U6569 (N_6569,N_4428,N_4029);
xor U6570 (N_6570,N_4146,N_2324);
nor U6571 (N_6571,N_1056,N_4296);
nor U6572 (N_6572,N_206,N_2107);
or U6573 (N_6573,N_2660,N_1001);
or U6574 (N_6574,N_385,N_4919);
and U6575 (N_6575,N_1330,N_3415);
or U6576 (N_6576,N_2515,N_3686);
nand U6577 (N_6577,N_2396,N_1650);
nand U6578 (N_6578,N_3707,N_3824);
nor U6579 (N_6579,N_3178,N_529);
nor U6580 (N_6580,N_474,N_2384);
xor U6581 (N_6581,N_3331,N_3677);
or U6582 (N_6582,N_3835,N_3793);
nor U6583 (N_6583,N_3997,N_3209);
and U6584 (N_6584,N_2846,N_3559);
and U6585 (N_6585,N_1058,N_111);
and U6586 (N_6586,N_4340,N_1624);
nand U6587 (N_6587,N_2162,N_4249);
nor U6588 (N_6588,N_3575,N_709);
nor U6589 (N_6589,N_1432,N_130);
or U6590 (N_6590,N_2146,N_1174);
and U6591 (N_6591,N_2756,N_2875);
nand U6592 (N_6592,N_2345,N_1856);
nand U6593 (N_6593,N_2401,N_1956);
xnor U6594 (N_6594,N_3138,N_3317);
nor U6595 (N_6595,N_1826,N_3554);
xor U6596 (N_6596,N_2499,N_4610);
or U6597 (N_6597,N_4803,N_4259);
nor U6598 (N_6598,N_1549,N_2560);
nor U6599 (N_6599,N_856,N_2915);
nand U6600 (N_6600,N_2705,N_3311);
nand U6601 (N_6601,N_3288,N_761);
nand U6602 (N_6602,N_4961,N_1226);
or U6603 (N_6603,N_4447,N_2039);
nand U6604 (N_6604,N_2179,N_4299);
nand U6605 (N_6605,N_2067,N_3113);
xnor U6606 (N_6606,N_1431,N_2105);
and U6607 (N_6607,N_2114,N_2564);
nand U6608 (N_6608,N_1944,N_3394);
and U6609 (N_6609,N_4491,N_3336);
nor U6610 (N_6610,N_245,N_1308);
or U6611 (N_6611,N_2621,N_4431);
and U6612 (N_6612,N_666,N_850);
nor U6613 (N_6613,N_415,N_3732);
nor U6614 (N_6614,N_59,N_1918);
and U6615 (N_6615,N_3597,N_2392);
or U6616 (N_6616,N_1966,N_675);
nor U6617 (N_6617,N_3498,N_907);
nand U6618 (N_6618,N_3581,N_102);
or U6619 (N_6619,N_3654,N_394);
and U6620 (N_6620,N_4171,N_4705);
nor U6621 (N_6621,N_3350,N_468);
nand U6622 (N_6622,N_146,N_365);
and U6623 (N_6623,N_4860,N_2559);
and U6624 (N_6624,N_3152,N_3170);
and U6625 (N_6625,N_939,N_4841);
xnor U6626 (N_6626,N_2986,N_848);
nor U6627 (N_6627,N_2184,N_1757);
nand U6628 (N_6628,N_3701,N_2606);
or U6629 (N_6629,N_1498,N_1484);
or U6630 (N_6630,N_3819,N_3648);
and U6631 (N_6631,N_3532,N_1688);
nor U6632 (N_6632,N_1874,N_1652);
nor U6633 (N_6633,N_1662,N_748);
and U6634 (N_6634,N_1477,N_4112);
and U6635 (N_6635,N_2363,N_1272);
and U6636 (N_6636,N_1041,N_3202);
or U6637 (N_6637,N_541,N_521);
nor U6638 (N_6638,N_1003,N_3495);
or U6639 (N_6639,N_1601,N_4828);
or U6640 (N_6640,N_2443,N_4328);
or U6641 (N_6641,N_2588,N_1882);
or U6642 (N_6642,N_948,N_518);
nor U6643 (N_6643,N_89,N_4753);
and U6644 (N_6644,N_4260,N_350);
and U6645 (N_6645,N_4110,N_3941);
or U6646 (N_6646,N_9,N_1176);
nand U6647 (N_6647,N_3490,N_3126);
nor U6648 (N_6648,N_424,N_3477);
nor U6649 (N_6649,N_3021,N_1406);
or U6650 (N_6650,N_1043,N_2934);
nand U6651 (N_6651,N_2404,N_3741);
or U6652 (N_6652,N_1899,N_2239);
nor U6653 (N_6653,N_1585,N_1980);
nor U6654 (N_6654,N_2304,N_4645);
nand U6655 (N_6655,N_1614,N_472);
or U6656 (N_6656,N_2148,N_3075);
xor U6657 (N_6657,N_708,N_3367);
and U6658 (N_6658,N_4024,N_946);
xor U6659 (N_6659,N_3469,N_4794);
nor U6660 (N_6660,N_4579,N_4734);
and U6661 (N_6661,N_1263,N_4314);
nand U6662 (N_6662,N_154,N_1144);
nor U6663 (N_6663,N_2449,N_2896);
nand U6664 (N_6664,N_299,N_794);
and U6665 (N_6665,N_3696,N_3731);
and U6666 (N_6666,N_777,N_4250);
nor U6667 (N_6667,N_3180,N_4859);
or U6668 (N_6668,N_2205,N_222);
nand U6669 (N_6669,N_2424,N_3123);
nand U6670 (N_6670,N_3584,N_3667);
or U6671 (N_6671,N_159,N_4532);
xnor U6672 (N_6672,N_1387,N_1286);
nor U6673 (N_6673,N_3963,N_2191);
and U6674 (N_6674,N_3888,N_1383);
nand U6675 (N_6675,N_1071,N_1559);
nor U6676 (N_6676,N_3092,N_145);
or U6677 (N_6677,N_1347,N_1087);
or U6678 (N_6678,N_3868,N_3921);
xor U6679 (N_6679,N_3063,N_3831);
or U6680 (N_6680,N_747,N_3127);
nand U6681 (N_6681,N_867,N_2929);
xnor U6682 (N_6682,N_4133,N_2353);
and U6683 (N_6683,N_972,N_773);
nor U6684 (N_6684,N_4144,N_445);
and U6685 (N_6685,N_2437,N_4480);
nor U6686 (N_6686,N_3137,N_4104);
nor U6687 (N_6687,N_4960,N_749);
nor U6688 (N_6688,N_4944,N_4057);
nor U6689 (N_6689,N_3928,N_3284);
or U6690 (N_6690,N_2028,N_98);
nand U6691 (N_6691,N_4815,N_1440);
nand U6692 (N_6692,N_1267,N_2372);
nor U6693 (N_6693,N_4418,N_3717);
nor U6694 (N_6694,N_1184,N_4698);
or U6695 (N_6695,N_1666,N_1846);
xnor U6696 (N_6696,N_1042,N_1519);
and U6697 (N_6697,N_3175,N_2445);
and U6698 (N_6698,N_1537,N_4777);
nor U6699 (N_6699,N_1663,N_4615);
xor U6700 (N_6700,N_3049,N_1718);
or U6701 (N_6701,N_3774,N_664);
and U6702 (N_6702,N_4335,N_534);
xor U6703 (N_6703,N_976,N_2632);
and U6704 (N_6704,N_298,N_2630);
and U6705 (N_6705,N_2185,N_3392);
nor U6706 (N_6706,N_775,N_4281);
or U6707 (N_6707,N_2870,N_718);
nand U6708 (N_6708,N_160,N_398);
nand U6709 (N_6709,N_4456,N_1936);
nand U6710 (N_6710,N_1278,N_880);
and U6711 (N_6711,N_722,N_1373);
and U6712 (N_6712,N_2786,N_3407);
and U6713 (N_6713,N_265,N_4772);
and U6714 (N_6714,N_4407,N_3980);
and U6715 (N_6715,N_3231,N_1642);
and U6716 (N_6716,N_4563,N_418);
or U6717 (N_6717,N_3144,N_2693);
and U6718 (N_6718,N_1982,N_2373);
nand U6719 (N_6719,N_294,N_1636);
nand U6720 (N_6720,N_2116,N_278);
nand U6721 (N_6721,N_3937,N_539);
nand U6722 (N_6722,N_4497,N_1027);
nor U6723 (N_6723,N_450,N_1912);
or U6724 (N_6724,N_2060,N_1678);
or U6725 (N_6725,N_2196,N_1389);
nor U6726 (N_6726,N_1361,N_2008);
or U6727 (N_6727,N_1271,N_2209);
nand U6728 (N_6728,N_348,N_3803);
nand U6729 (N_6729,N_319,N_1608);
nand U6730 (N_6730,N_942,N_2289);
nand U6731 (N_6731,N_207,N_921);
or U6732 (N_6732,N_2208,N_2673);
nor U6733 (N_6733,N_1627,N_490);
nor U6734 (N_6734,N_593,N_572);
nor U6735 (N_6735,N_4175,N_3223);
nand U6736 (N_6736,N_3518,N_3913);
nor U6737 (N_6737,N_3012,N_3133);
nor U6738 (N_6738,N_4056,N_1425);
and U6739 (N_6739,N_4786,N_1197);
nand U6740 (N_6740,N_19,N_4577);
and U6741 (N_6741,N_1748,N_3595);
nand U6742 (N_6742,N_3481,N_647);
nor U6743 (N_6743,N_1281,N_668);
and U6744 (N_6744,N_4473,N_331);
or U6745 (N_6745,N_835,N_1208);
nand U6746 (N_6746,N_4602,N_3520);
or U6747 (N_6747,N_4706,N_1172);
nor U6748 (N_6748,N_625,N_85);
or U6749 (N_6749,N_3303,N_3128);
nand U6750 (N_6750,N_3340,N_4050);
and U6751 (N_6751,N_4738,N_1037);
nand U6752 (N_6752,N_3177,N_3661);
nor U6753 (N_6753,N_3358,N_4164);
and U6754 (N_6754,N_853,N_4855);
nand U6755 (N_6755,N_4386,N_2323);
and U6756 (N_6756,N_3567,N_610);
or U6757 (N_6757,N_2243,N_3621);
xor U6758 (N_6758,N_898,N_2276);
and U6759 (N_6759,N_2640,N_789);
and U6760 (N_6760,N_3758,N_2641);
and U6761 (N_6761,N_4277,N_2652);
nand U6762 (N_6762,N_432,N_2409);
nand U6763 (N_6763,N_2011,N_3926);
or U6764 (N_6764,N_114,N_3299);
or U6765 (N_6765,N_1603,N_2326);
and U6766 (N_6766,N_3457,N_3594);
or U6767 (N_6767,N_4540,N_3100);
nand U6768 (N_6768,N_386,N_277);
nor U6769 (N_6769,N_3061,N_216);
nor U6770 (N_6770,N_2847,N_1563);
and U6771 (N_6771,N_3080,N_270);
and U6772 (N_6772,N_4915,N_2534);
nor U6773 (N_6773,N_806,N_601);
and U6774 (N_6774,N_2707,N_4748);
and U6775 (N_6775,N_2314,N_843);
nor U6776 (N_6776,N_1270,N_192);
nor U6777 (N_6777,N_3895,N_3319);
or U6778 (N_6778,N_2839,N_3224);
or U6779 (N_6779,N_1099,N_3391);
or U6780 (N_6780,N_1405,N_454);
nor U6781 (N_6781,N_644,N_1407);
and U6782 (N_6782,N_3591,N_2103);
and U6783 (N_6783,N_1556,N_4528);
nand U6784 (N_6784,N_4752,N_434);
nand U6785 (N_6785,N_1313,N_752);
or U6786 (N_6786,N_492,N_1159);
nor U6787 (N_6787,N_3417,N_774);
nand U6788 (N_6788,N_1434,N_1760);
nor U6789 (N_6789,N_132,N_4088);
and U6790 (N_6790,N_2689,N_4887);
or U6791 (N_6791,N_4247,N_4130);
nor U6792 (N_6792,N_3739,N_3812);
or U6793 (N_6793,N_886,N_887);
nor U6794 (N_6794,N_3529,N_3838);
or U6795 (N_6795,N_4682,N_683);
or U6796 (N_6796,N_1797,N_2434);
xor U6797 (N_6797,N_228,N_2578);
nor U6798 (N_6798,N_2238,N_3713);
nand U6799 (N_6799,N_2143,N_3932);
nor U6800 (N_6800,N_2398,N_4814);
and U6801 (N_6801,N_4973,N_4068);
and U6802 (N_6802,N_1442,N_3346);
nor U6803 (N_6803,N_14,N_22);
nand U6804 (N_6804,N_4503,N_2737);
nand U6805 (N_6805,N_2543,N_1301);
nor U6806 (N_6806,N_2822,N_2524);
and U6807 (N_6807,N_7,N_3398);
and U6808 (N_6808,N_4703,N_4599);
nand U6809 (N_6809,N_2061,N_2484);
and U6810 (N_6810,N_4048,N_382);
nand U6811 (N_6811,N_2871,N_2252);
nand U6812 (N_6812,N_239,N_2258);
xnor U6813 (N_6813,N_2310,N_2154);
xor U6814 (N_6814,N_3905,N_594);
and U6815 (N_6815,N_4716,N_1247);
xor U6816 (N_6816,N_1903,N_4785);
nor U6817 (N_6817,N_3599,N_2497);
or U6818 (N_6818,N_4346,N_2716);
xnor U6819 (N_6819,N_3743,N_1863);
nor U6820 (N_6820,N_4628,N_61);
xnor U6821 (N_6821,N_3159,N_2583);
or U6822 (N_6822,N_4419,N_1692);
xnor U6823 (N_6823,N_4797,N_3455);
xnor U6824 (N_6824,N_3034,N_1242);
nor U6825 (N_6825,N_1296,N_4861);
nand U6826 (N_6826,N_4825,N_4216);
nor U6827 (N_6827,N_778,N_4039);
nor U6828 (N_6828,N_3435,N_3780);
or U6829 (N_6829,N_3215,N_4001);
nor U6830 (N_6830,N_2571,N_3334);
or U6831 (N_6831,N_578,N_4019);
nand U6832 (N_6832,N_564,N_1525);
nor U6833 (N_6833,N_88,N_1460);
nand U6834 (N_6834,N_1592,N_4143);
nand U6835 (N_6835,N_4158,N_3420);
nor U6836 (N_6836,N_1992,N_3095);
and U6837 (N_6837,N_471,N_4922);
nor U6838 (N_6838,N_3652,N_4917);
and U6839 (N_6839,N_2614,N_1234);
nand U6840 (N_6840,N_4388,N_1629);
and U6841 (N_6841,N_2195,N_3283);
nand U6842 (N_6842,N_4100,N_1753);
and U6843 (N_6843,N_1561,N_1951);
and U6844 (N_6844,N_4710,N_3855);
or U6845 (N_6845,N_1342,N_2459);
nand U6846 (N_6846,N_3796,N_2019);
nand U6847 (N_6847,N_1949,N_4758);
and U6848 (N_6848,N_3678,N_2762);
or U6849 (N_6849,N_3147,N_1501);
or U6850 (N_6850,N_2050,N_4687);
nand U6851 (N_6851,N_3158,N_293);
or U6852 (N_6852,N_374,N_3339);
nand U6853 (N_6853,N_3521,N_3210);
nor U6854 (N_6854,N_4330,N_2069);
nor U6855 (N_6855,N_4747,N_695);
nand U6856 (N_6856,N_851,N_422);
or U6857 (N_6857,N_658,N_2228);
and U6858 (N_6858,N_1470,N_1493);
and U6859 (N_6859,N_448,N_3994);
nor U6860 (N_6860,N_1970,N_2033);
or U6861 (N_6861,N_4387,N_3873);
nor U6862 (N_6862,N_4238,N_655);
nor U6863 (N_6863,N_1279,N_3979);
and U6864 (N_6864,N_3784,N_52);
nand U6865 (N_6865,N_0,N_700);
xor U6866 (N_6866,N_1702,N_4719);
nand U6867 (N_6867,N_2340,N_4827);
nand U6868 (N_6868,N_1750,N_1283);
and U6869 (N_6869,N_1318,N_2530);
and U6870 (N_6870,N_2603,N_2088);
nor U6871 (N_6871,N_1833,N_1304);
or U6872 (N_6872,N_2594,N_4545);
nand U6873 (N_6873,N_3181,N_1170);
nor U6874 (N_6874,N_1822,N_3154);
or U6875 (N_6875,N_2361,N_1183);
nand U6876 (N_6876,N_4711,N_4082);
and U6877 (N_6877,N_4466,N_2201);
and U6878 (N_6878,N_2390,N_3120);
and U6879 (N_6879,N_3241,N_2375);
or U6880 (N_6880,N_2819,N_4680);
or U6881 (N_6881,N_2458,N_674);
nand U6882 (N_6882,N_4140,N_2845);
or U6883 (N_6883,N_2101,N_3116);
and U6884 (N_6884,N_4928,N_3315);
and U6885 (N_6885,N_935,N_4003);
and U6886 (N_6886,N_2100,N_3140);
or U6887 (N_6887,N_2967,N_4379);
nor U6888 (N_6888,N_4375,N_1002);
nor U6889 (N_6889,N_3124,N_1581);
and U6890 (N_6890,N_1443,N_4033);
and U6891 (N_6891,N_2187,N_1180);
or U6892 (N_6892,N_4364,N_2981);
and U6893 (N_6893,N_66,N_2226);
and U6894 (N_6894,N_3428,N_2405);
and U6895 (N_6895,N_2102,N_3513);
nor U6896 (N_6896,N_3547,N_2138);
xnor U6897 (N_6897,N_1437,N_4562);
or U6898 (N_6898,N_807,N_1914);
or U6899 (N_6899,N_2789,N_1462);
nand U6900 (N_6900,N_2153,N_2976);
nand U6901 (N_6901,N_3766,N_1643);
or U6902 (N_6902,N_2292,N_2874);
nor U6903 (N_6903,N_3545,N_4319);
or U6904 (N_6904,N_643,N_525);
nor U6905 (N_6905,N_1836,N_633);
nand U6906 (N_6906,N_380,N_4901);
nand U6907 (N_6907,N_938,N_2078);
or U6908 (N_6908,N_703,N_2700);
nand U6909 (N_6909,N_2406,N_649);
and U6910 (N_6910,N_4382,N_4078);
or U6911 (N_6911,N_2287,N_2009);
and U6912 (N_6912,N_4455,N_4321);
or U6913 (N_6913,N_1126,N_40);
nor U6914 (N_6914,N_1796,N_4173);
nand U6915 (N_6915,N_463,N_1331);
nor U6916 (N_6916,N_857,N_825);
nor U6917 (N_6917,N_3153,N_937);
and U6918 (N_6918,N_3281,N_2468);
nand U6919 (N_6919,N_2697,N_459);
nor U6920 (N_6920,N_378,N_2236);
and U6921 (N_6921,N_3410,N_250);
and U6922 (N_6922,N_3323,N_271);
or U6923 (N_6923,N_2761,N_1515);
nor U6924 (N_6924,N_3609,N_3419);
nand U6925 (N_6925,N_3787,N_4420);
or U6926 (N_6926,N_3261,N_4412);
or U6927 (N_6927,N_2683,N_3823);
nor U6928 (N_6928,N_122,N_302);
nand U6929 (N_6929,N_2687,N_2586);
nand U6930 (N_6930,N_4878,N_3801);
or U6931 (N_6931,N_45,N_989);
and U6932 (N_6932,N_949,N_17);
nand U6933 (N_6933,N_4009,N_2522);
nand U6934 (N_6934,N_3471,N_2022);
or U6935 (N_6935,N_3845,N_1022);
and U6936 (N_6936,N_1292,N_473);
or U6937 (N_6937,N_4231,N_2249);
xor U6938 (N_6938,N_980,N_480);
nand U6939 (N_6939,N_2334,N_4982);
xor U6940 (N_6940,N_4468,N_2556);
or U6941 (N_6941,N_2305,N_2480);
or U6942 (N_6942,N_495,N_403);
or U6943 (N_6943,N_295,N_3541);
nor U6944 (N_6944,N_1105,N_2865);
nor U6945 (N_6945,N_1193,N_2704);
nand U6946 (N_6946,N_2130,N_2777);
nand U6947 (N_6947,N_2407,N_1130);
and U6948 (N_6948,N_1919,N_1562);
nand U6949 (N_6949,N_4601,N_4519);
xnor U6950 (N_6950,N_1917,N_4607);
xor U6951 (N_6951,N_573,N_940);
nand U6952 (N_6952,N_2059,N_3854);
nand U6953 (N_6953,N_516,N_301);
nor U6954 (N_6954,N_325,N_3211);
or U6955 (N_6955,N_1384,N_4153);
and U6956 (N_6956,N_757,N_3506);
xnor U6957 (N_6957,N_399,N_3896);
nor U6958 (N_6958,N_4157,N_4598);
nor U6959 (N_6959,N_930,N_1866);
nor U6960 (N_6960,N_2956,N_3883);
and U6961 (N_6961,N_4195,N_2021);
and U6962 (N_6962,N_4262,N_4099);
nand U6963 (N_6963,N_342,N_4802);
nor U6964 (N_6964,N_1789,N_715);
or U6965 (N_6965,N_2042,N_2783);
nor U6966 (N_6966,N_3570,N_2759);
and U6967 (N_6967,N_1015,N_4539);
nor U6968 (N_6968,N_4461,N_4464);
and U6969 (N_6969,N_1205,N_4059);
or U6970 (N_6970,N_1641,N_2488);
and U6971 (N_6971,N_4744,N_1569);
xor U6972 (N_6972,N_65,N_559);
and U6973 (N_6973,N_393,N_2118);
xnor U6974 (N_6974,N_3981,N_871);
or U6975 (N_6975,N_1596,N_2419);
xor U6976 (N_6976,N_963,N_1163);
nor U6977 (N_6977,N_1250,N_3413);
or U6978 (N_6978,N_3655,N_4916);
or U6979 (N_6979,N_3556,N_478);
nor U6980 (N_6980,N_4543,N_2230);
nand U6981 (N_6981,N_766,N_1645);
nor U6982 (N_6982,N_4684,N_4207);
nand U6983 (N_6983,N_1736,N_3764);
or U6984 (N_6984,N_3761,N_2229);
nand U6985 (N_6985,N_3173,N_193);
or U6986 (N_6986,N_706,N_3071);
nand U6987 (N_6987,N_2602,N_1438);
or U6988 (N_6988,N_20,N_2852);
or U6989 (N_6989,N_1551,N_3268);
xnor U6990 (N_6990,N_2456,N_1621);
and U6991 (N_6991,N_1488,N_3099);
or U6992 (N_6992,N_4290,N_4268);
or U6993 (N_6993,N_2151,N_163);
and U6994 (N_6994,N_3645,N_1337);
or U6995 (N_6995,N_915,N_1639);
xor U6996 (N_6996,N_1155,N_801);
nor U6997 (N_6997,N_1466,N_1859);
xor U6998 (N_6998,N_1932,N_2075);
nor U6999 (N_6999,N_734,N_1574);
nor U7000 (N_7000,N_730,N_2876);
nor U7001 (N_7001,N_3492,N_3552);
xnor U7002 (N_7002,N_4799,N_1067);
and U7003 (N_7003,N_597,N_1465);
nor U7004 (N_7004,N_4937,N_4020);
nor U7005 (N_7005,N_3087,N_1187);
nor U7006 (N_7006,N_1976,N_3798);
or U7007 (N_7007,N_1216,N_3704);
nand U7008 (N_7008,N_1463,N_3025);
xor U7009 (N_7009,N_1265,N_1385);
nor U7010 (N_7010,N_1828,N_4363);
or U7011 (N_7011,N_1084,N_4779);
or U7012 (N_7012,N_2403,N_639);
nor U7013 (N_7013,N_4534,N_2838);
and U7014 (N_7014,N_1120,N_1553);
or U7015 (N_7015,N_3929,N_3414);
or U7016 (N_7016,N_2425,N_2076);
nand U7017 (N_7017,N_458,N_988);
or U7018 (N_7018,N_1957,N_3105);
nor U7019 (N_7019,N_1795,N_4115);
or U7020 (N_7020,N_4629,N_2978);
nor U7021 (N_7021,N_543,N_767);
and U7022 (N_7022,N_1036,N_3566);
or U7023 (N_7023,N_1701,N_841);
nand U7024 (N_7024,N_3786,N_1485);
nor U7025 (N_7025,N_3974,N_958);
nand U7026 (N_7026,N_3321,N_107);
and U7027 (N_7027,N_2928,N_1761);
and U7028 (N_7028,N_858,N_2082);
or U7029 (N_7029,N_161,N_2477);
or U7030 (N_7030,N_1030,N_552);
nor U7031 (N_7031,N_3059,N_4914);
nor U7032 (N_7032,N_3245,N_3923);
nor U7033 (N_7033,N_3860,N_1651);
nor U7034 (N_7034,N_990,N_2575);
and U7035 (N_7035,N_4189,N_1588);
xnor U7036 (N_7036,N_4836,N_2256);
xor U7037 (N_7037,N_4614,N_3810);
nor U7038 (N_7038,N_408,N_4211);
or U7039 (N_7039,N_3015,N_180);
and U7040 (N_7040,N_943,N_3685);
xor U7041 (N_7041,N_3510,N_1380);
or U7042 (N_7042,N_2399,N_961);
and U7043 (N_7043,N_3753,N_3991);
and U7044 (N_7044,N_4235,N_3165);
and U7045 (N_7045,N_2041,N_3446);
and U7046 (N_7046,N_1780,N_3110);
or U7047 (N_7047,N_407,N_1659);
nor U7048 (N_7048,N_2546,N_3914);
xnor U7049 (N_7049,N_4162,N_4463);
nor U7050 (N_7050,N_710,N_3613);
or U7051 (N_7051,N_1366,N_4864);
nand U7052 (N_7052,N_4323,N_3844);
nor U7053 (N_7053,N_1705,N_1369);
xnor U7054 (N_7054,N_4306,N_997);
xor U7055 (N_7055,N_2751,N_233);
and U7056 (N_7056,N_3053,N_4030);
and U7057 (N_7057,N_3965,N_476);
nor U7058 (N_7058,N_3546,N_4049);
nand U7059 (N_7059,N_3436,N_1376);
or U7060 (N_7060,N_4303,N_4837);
nand U7061 (N_7061,N_888,N_587);
or U7062 (N_7062,N_4408,N_210);
and U7063 (N_7063,N_2655,N_3849);
nand U7064 (N_7064,N_2346,N_1817);
and U7065 (N_7065,N_4862,N_4833);
and U7066 (N_7066,N_3583,N_1873);
and U7067 (N_7067,N_4044,N_2709);
xor U7068 (N_7068,N_4424,N_3755);
or U7069 (N_7069,N_528,N_1734);
nand U7070 (N_7070,N_4640,N_4955);
or U7071 (N_7071,N_1268,N_1876);
and U7072 (N_7072,N_1508,N_1153);
xnor U7073 (N_7073,N_3273,N_2662);
or U7074 (N_7074,N_1076,N_2825);
nor U7075 (N_7075,N_1694,N_2432);
xor U7076 (N_7076,N_2639,N_4821);
nor U7077 (N_7077,N_770,N_4462);
xnor U7078 (N_7078,N_4061,N_3919);
and U7079 (N_7079,N_2605,N_4017);
and U7080 (N_7080,N_2994,N_3174);
and U7081 (N_7081,N_546,N_763);
xnor U7082 (N_7082,N_1040,N_1023);
nor U7083 (N_7083,N_1628,N_3722);
xor U7084 (N_7084,N_3267,N_2417);
nor U7085 (N_7085,N_4776,N_3806);
xnor U7086 (N_7086,N_4945,N_1799);
and U7087 (N_7087,N_900,N_4108);
or U7088 (N_7088,N_4662,N_2046);
or U7089 (N_7089,N_2866,N_1258);
nand U7090 (N_7090,N_4967,N_1840);
xnor U7091 (N_7091,N_2186,N_735);
nand U7092 (N_7092,N_1518,N_3927);
nor U7093 (N_7093,N_347,N_1423);
or U7094 (N_7094,N_430,N_3775);
nor U7095 (N_7095,N_3320,N_1404);
or U7096 (N_7096,N_3542,N_4204);
nand U7097 (N_7097,N_698,N_2014);
or U7098 (N_7098,N_3307,N_164);
and U7099 (N_7099,N_2916,N_3925);
or U7100 (N_7100,N_1764,N_3139);
and U7101 (N_7101,N_4842,N_2653);
nand U7102 (N_7102,N_1552,N_3788);
or U7103 (N_7103,N_903,N_3274);
xnor U7104 (N_7104,N_3354,N_3001);
nand U7105 (N_7105,N_2266,N_4957);
nor U7106 (N_7106,N_1469,N_416);
and U7107 (N_7107,N_3192,N_3017);
and U7108 (N_7108,N_2336,N_2607);
and U7109 (N_7109,N_3674,N_3470);
nand U7110 (N_7110,N_218,N_3280);
and U7111 (N_7111,N_2755,N_2698);
or U7112 (N_7112,N_3644,N_4505);
or U7113 (N_7113,N_2089,N_2906);
or U7114 (N_7114,N_648,N_3387);
nand U7115 (N_7115,N_62,N_2725);
and U7116 (N_7116,N_3044,N_2302);
nor U7117 (N_7117,N_1411,N_4036);
nor U7118 (N_7118,N_2024,N_4288);
or U7119 (N_7119,N_3543,N_4275);
and U7120 (N_7120,N_3359,N_3408);
nor U7121 (N_7121,N_631,N_3377);
and U7122 (N_7122,N_822,N_4754);
nand U7123 (N_7123,N_3402,N_2265);
nand U7124 (N_7124,N_4434,N_1810);
nand U7125 (N_7125,N_1175,N_1011);
nor U7126 (N_7126,N_3876,N_4641);
nand U7127 (N_7127,N_1359,N_4771);
and U7128 (N_7128,N_395,N_2139);
nand U7129 (N_7129,N_479,N_2371);
xnor U7130 (N_7130,N_4089,N_3908);
nand U7131 (N_7131,N_2428,N_3000);
nand U7132 (N_7132,N_1875,N_4676);
and U7133 (N_7133,N_3893,N_595);
nand U7134 (N_7134,N_1305,N_3482);
or U7135 (N_7135,N_447,N_1971);
or U7136 (N_7136,N_1345,N_3088);
xnor U7137 (N_7137,N_4373,N_3055);
nor U7138 (N_7138,N_103,N_3324);
or U7139 (N_7139,N_626,N_3875);
or U7140 (N_7140,N_3964,N_3912);
or U7141 (N_7141,N_3629,N_2317);
or U7142 (N_7142,N_258,N_1339);
xnor U7143 (N_7143,N_51,N_762);
and U7144 (N_7144,N_3818,N_1512);
nand U7145 (N_7145,N_2962,N_2277);
nor U7146 (N_7146,N_2987,N_2473);
or U7147 (N_7147,N_2746,N_153);
nand U7148 (N_7148,N_1744,N_482);
or U7149 (N_7149,N_82,N_3051);
xor U7150 (N_7150,N_2891,N_3847);
or U7151 (N_7151,N_501,N_409);
nor U7152 (N_7152,N_3427,N_143);
and U7153 (N_7153,N_1605,N_4215);
and U7154 (N_7154,N_2222,N_2864);
nor U7155 (N_7155,N_2567,N_4526);
and U7156 (N_7156,N_1767,N_2260);
xor U7157 (N_7157,N_1322,N_353);
and U7158 (N_7158,N_669,N_1114);
nand U7159 (N_7159,N_4897,N_979);
and U7160 (N_7160,N_2732,N_1560);
and U7161 (N_7161,N_4835,N_3006);
or U7162 (N_7162,N_4034,N_3501);
xor U7163 (N_7163,N_4225,N_2160);
nor U7164 (N_7164,N_2850,N_2389);
xnor U7165 (N_7165,N_719,N_2232);
or U7166 (N_7166,N_3757,N_3353);
nand U7167 (N_7167,N_2853,N_3515);
nand U7168 (N_7168,N_3946,N_3702);
nand U7169 (N_7169,N_3449,N_2960);
nand U7170 (N_7170,N_315,N_2880);
nor U7171 (N_7171,N_4177,N_4092);
nand U7172 (N_7172,N_576,N_4075);
nand U7173 (N_7173,N_4782,N_3638);
nand U7174 (N_7174,N_4429,N_3330);
nand U7175 (N_7175,N_3076,N_1051);
nor U7176 (N_7176,N_3142,N_1274);
nand U7177 (N_7177,N_3719,N_1355);
nand U7178 (N_7178,N_2109,N_3641);
and U7179 (N_7179,N_177,N_3074);
and U7180 (N_7180,N_3565,N_2890);
and U7181 (N_7181,N_785,N_1800);
nor U7182 (N_7182,N_975,N_797);
nor U7183 (N_7183,N_227,N_2984);
nand U7184 (N_7184,N_697,N_2592);
and U7185 (N_7185,N_1075,N_201);
xor U7186 (N_7186,N_1623,N_4047);
and U7187 (N_7187,N_1947,N_4342);
nand U7188 (N_7188,N_2206,N_4846);
and U7189 (N_7189,N_2475,N_2422);
nand U7190 (N_7190,N_524,N_1093);
xor U7191 (N_7191,N_4438,N_4806);
nor U7192 (N_7192,N_3388,N_2823);
nor U7193 (N_7193,N_1019,N_4071);
xnor U7194 (N_7194,N_1238,N_1612);
nand U7195 (N_7195,N_1604,N_4696);
and U7196 (N_7196,N_3605,N_4712);
nand U7197 (N_7197,N_332,N_4226);
nand U7198 (N_7198,N_1915,N_884);
nand U7199 (N_7199,N_3694,N_1622);
nor U7200 (N_7200,N_2717,N_1746);
nand U7201 (N_7201,N_3822,N_3098);
and U7202 (N_7202,N_75,N_1445);
nand U7203 (N_7203,N_288,N_1334);
or U7204 (N_7204,N_795,N_4531);
or U7205 (N_7205,N_2827,N_3886);
nand U7206 (N_7206,N_451,N_4103);
nor U7207 (N_7207,N_2058,N_927);
or U7208 (N_7208,N_2923,N_467);
and U7209 (N_7209,N_3254,N_4472);
and U7210 (N_7210,N_4800,N_4646);
xnor U7211 (N_7211,N_1316,N_2344);
or U7212 (N_7212,N_1706,N_4196);
and U7213 (N_7213,N_2809,N_4818);
and U7214 (N_7214,N_4135,N_1935);
or U7215 (N_7215,N_3108,N_1740);
nor U7216 (N_7216,N_358,N_1928);
nor U7217 (N_7217,N_4469,N_832);
or U7218 (N_7218,N_126,N_1788);
or U7219 (N_7219,N_3500,N_917);
and U7220 (N_7220,N_282,N_1853);
nand U7221 (N_7221,N_229,N_3467);
and U7222 (N_7222,N_2207,N_2123);
and U7223 (N_7223,N_2053,N_4675);
nand U7224 (N_7224,N_4378,N_355);
nor U7225 (N_7225,N_2066,N_4251);
nor U7226 (N_7226,N_4895,N_1923);
nor U7227 (N_7227,N_705,N_2062);
and U7228 (N_7228,N_339,N_1835);
nand U7229 (N_7229,N_1118,N_2472);
nand U7230 (N_7230,N_2775,N_4022);
nand U7231 (N_7231,N_1547,N_3856);
or U7232 (N_7232,N_813,N_542);
and U7233 (N_7233,N_4991,N_3762);
and U7234 (N_7234,N_772,N_2032);
nor U7235 (N_7235,N_3951,N_1294);
nor U7236 (N_7236,N_291,N_3616);
nand U7237 (N_7237,N_1161,N_4938);
nand U7238 (N_7238,N_1900,N_2860);
nand U7239 (N_7239,N_2651,N_3296);
or U7240 (N_7240,N_3770,N_4784);
or U7241 (N_7241,N_4743,N_3548);
nor U7242 (N_7242,N_1964,N_4137);
or U7243 (N_7243,N_3897,N_583);
or U7244 (N_7244,N_1555,N_1479);
nor U7245 (N_7245,N_1657,N_4995);
nand U7246 (N_7246,N_4574,N_561);
nand U7247 (N_7247,N_1769,N_1262);
or U7248 (N_7248,N_3374,N_175);
nand U7249 (N_7249,N_4016,N_3072);
nand U7250 (N_7250,N_4863,N_2706);
and U7251 (N_7251,N_3935,N_3304);
or U7252 (N_7252,N_3356,N_4768);
and U7253 (N_7253,N_3817,N_2760);
nor U7254 (N_7254,N_1110,N_3114);
nor U7255 (N_7255,N_3836,N_2995);
xor U7256 (N_7256,N_3328,N_3289);
nor U7257 (N_7257,N_4120,N_76);
or U7258 (N_7258,N_234,N_2465);
nor U7259 (N_7259,N_3978,N_4446);
and U7260 (N_7260,N_4853,N_2914);
xor U7261 (N_7261,N_2931,N_466);
and U7262 (N_7262,N_2920,N_2817);
or U7263 (N_7263,N_465,N_3028);
and U7264 (N_7264,N_1032,N_4320);
or U7265 (N_7265,N_3089,N_4677);
nand U7266 (N_7266,N_2980,N_960);
and U7267 (N_7267,N_2442,N_3904);
nand U7268 (N_7268,N_4167,N_3841);
or U7269 (N_7269,N_1851,N_3636);
nand U7270 (N_7270,N_4309,N_2092);
xor U7271 (N_7271,N_4896,N_4084);
nor U7272 (N_7272,N_2338,N_1426);
xor U7273 (N_7273,N_4998,N_3437);
or U7274 (N_7274,N_3487,N_2620);
nor U7275 (N_7275,N_104,N_4774);
nand U7276 (N_7276,N_3830,N_654);
and U7277 (N_7277,N_326,N_3485);
nand U7278 (N_7278,N_3802,N_2541);
or U7279 (N_7279,N_1333,N_1046);
nand U7280 (N_7280,N_4936,N_1837);
and U7281 (N_7281,N_3958,N_3032);
or U7282 (N_7282,N_4749,N_4618);
and U7283 (N_7283,N_1719,N_1925);
nor U7284 (N_7284,N_1492,N_2793);
nor U7285 (N_7285,N_1691,N_3411);
nand U7286 (N_7286,N_3325,N_4222);
xnor U7287 (N_7287,N_46,N_1567);
and U7288 (N_7288,N_3474,N_3526);
and U7289 (N_7289,N_2912,N_3275);
nand U7290 (N_7290,N_3544,N_2841);
xnor U7291 (N_7291,N_2242,N_74);
xor U7292 (N_7292,N_4848,N_4055);
or U7293 (N_7293,N_3750,N_873);
nand U7294 (N_7294,N_993,N_4263);
nand U7295 (N_7295,N_2964,N_2937);
nand U7296 (N_7296,N_3475,N_4965);
or U7297 (N_7297,N_2999,N_1240);
or U7298 (N_7298,N_4376,N_1372);
nand U7299 (N_7299,N_4265,N_4344);
and U7300 (N_7300,N_3872,N_117);
or U7301 (N_7301,N_1531,N_4838);
nor U7302 (N_7302,N_1983,N_1722);
nand U7303 (N_7303,N_3318,N_338);
nor U7304 (N_7304,N_4819,N_2367);
and U7305 (N_7305,N_2878,N_4612);
xor U7306 (N_7306,N_4494,N_1707);
nand U7307 (N_7307,N_897,N_2935);
nor U7308 (N_7308,N_874,N_1248);
and U7309 (N_7309,N_12,N_4905);
nor U7310 (N_7310,N_300,N_4865);
and U7311 (N_7311,N_2359,N_485);
or U7312 (N_7312,N_3962,N_1490);
nor U7313 (N_7313,N_3257,N_953);
nor U7314 (N_7314,N_2090,N_3840);
or U7315 (N_7315,N_1616,N_38);
or U7316 (N_7316,N_3767,N_80);
nor U7317 (N_7317,N_2415,N_3360);
or U7318 (N_7318,N_590,N_1131);
nor U7319 (N_7319,N_2692,N_1080);
or U7320 (N_7320,N_640,N_4435);
nand U7321 (N_7321,N_1367,N_614);
xnor U7322 (N_7322,N_2966,N_3653);
and U7323 (N_7323,N_2385,N_3811);
or U7324 (N_7324,N_2537,N_2263);
nor U7325 (N_7325,N_3370,N_487);
nand U7326 (N_7326,N_3915,N_4510);
nor U7327 (N_7327,N_4843,N_4742);
or U7328 (N_7328,N_4780,N_2269);
or U7329 (N_7329,N_4483,N_2922);
or U7330 (N_7330,N_1808,N_3188);
and U7331 (N_7331,N_3642,N_1711);
and U7332 (N_7332,N_2382,N_4512);
or U7333 (N_7333,N_955,N_1483);
nand U7334 (N_7334,N_4355,N_3723);
nand U7335 (N_7335,N_3422,N_1625);
or U7336 (N_7336,N_1251,N_2366);
nor U7337 (N_7337,N_556,N_3715);
xnor U7338 (N_7338,N_58,N_4798);
nand U7339 (N_7339,N_924,N_4232);
nor U7340 (N_7340,N_457,N_2805);
or U7341 (N_7341,N_4000,N_3256);
xnor U7342 (N_7342,N_3918,N_1414);
nand U7343 (N_7343,N_4731,N_707);
nor U7344 (N_7344,N_1086,N_3081);
nor U7345 (N_7345,N_4987,N_3943);
nor U7346 (N_7346,N_4538,N_2098);
nor U7347 (N_7347,N_4552,N_1591);
nand U7348 (N_7348,N_1610,N_1768);
or U7349 (N_7349,N_3578,N_3659);
xnor U7350 (N_7350,N_4307,N_4630);
nor U7351 (N_7351,N_3016,N_3907);
xnor U7352 (N_7352,N_535,N_1038);
nor U7353 (N_7353,N_2535,N_3237);
and U7354 (N_7354,N_599,N_4691);
nand U7355 (N_7355,N_1536,N_2341);
or U7356 (N_7356,N_3442,N_4291);
nor U7357 (N_7357,N_4228,N_3011);
nor U7358 (N_7358,N_1459,N_4297);
nand U7359 (N_7359,N_1516,N_1390);
nor U7360 (N_7360,N_1696,N_3602);
nor U7361 (N_7361,N_4880,N_1698);
or U7362 (N_7362,N_1667,N_4983);
xnor U7363 (N_7363,N_400,N_2785);
or U7364 (N_7364,N_1177,N_3416);
nand U7365 (N_7365,N_1441,N_526);
or U7366 (N_7366,N_1497,N_1726);
nand U7367 (N_7367,N_1841,N_4511);
or U7368 (N_7368,N_384,N_3102);
nand U7369 (N_7369,N_629,N_3312);
and U7370 (N_7370,N_4638,N_3944);
and U7371 (N_7371,N_4093,N_4673);
and U7372 (N_7372,N_1195,N_3301);
nor U7373 (N_7373,N_1474,N_70);
or U7374 (N_7374,N_1429,N_4212);
or U7375 (N_7375,N_1381,N_4500);
or U7376 (N_7376,N_269,N_4432);
or U7377 (N_7377,N_2873,N_1770);
xnor U7378 (N_7378,N_3966,N_2126);
or U7379 (N_7379,N_1940,N_2331);
and U7380 (N_7380,N_657,N_1192);
nor U7381 (N_7381,N_167,N_3285);
nor U7382 (N_7382,N_4499,N_3310);
nor U7383 (N_7383,N_2561,N_1972);
xnor U7384 (N_7384,N_4174,N_1101);
nor U7385 (N_7385,N_1403,N_720);
nor U7386 (N_7386,N_4811,N_4188);
nand U7387 (N_7387,N_3582,N_2900);
nand U7388 (N_7388,N_1648,N_4805);
xnor U7389 (N_7389,N_489,N_820);
xnor U7390 (N_7390,N_3577,N_3431);
or U7391 (N_7391,N_4823,N_1545);
nor U7392 (N_7392,N_443,N_3754);
nor U7393 (N_7393,N_1122,N_1196);
nand U7394 (N_7394,N_1741,N_4289);
nor U7395 (N_7395,N_515,N_4595);
or U7396 (N_7396,N_1832,N_1654);
nand U7397 (N_7397,N_1491,N_4484);
and U7398 (N_7398,N_33,N_2144);
nor U7399 (N_7399,N_3535,N_2231);
nand U7400 (N_7400,N_3270,N_4150);
or U7401 (N_7401,N_3706,N_4183);
and U7402 (N_7402,N_56,N_2968);
or U7403 (N_7403,N_1535,N_2782);
nor U7404 (N_7404,N_1452,N_369);
or U7405 (N_7405,N_2623,N_1995);
or U7406 (N_7406,N_235,N_1529);
and U7407 (N_7407,N_642,N_381);
xnor U7408 (N_7408,N_41,N_3238);
and U7409 (N_7409,N_3078,N_257);
nand U7410 (N_7410,N_4452,N_442);
and U7411 (N_7411,N_2842,N_3036);
nor U7412 (N_7412,N_2194,N_2576);
xor U7413 (N_7413,N_4517,N_995);
nand U7414 (N_7414,N_4043,N_4537);
nand U7415 (N_7415,N_2376,N_4203);
and U7416 (N_7416,N_2461,N_3451);
nand U7417 (N_7417,N_3033,N_4350);
and U7418 (N_7418,N_1365,N_4481);
nand U7419 (N_7419,N_4726,N_63);
and U7420 (N_7420,N_4181,N_3975);
xor U7421 (N_7421,N_4513,N_328);
and U7422 (N_7422,N_1136,N_2552);
and U7423 (N_7423,N_3066,N_4358);
and U7424 (N_7424,N_1578,N_3726);
or U7425 (N_7425,N_165,N_1065);
or U7426 (N_7426,N_2244,N_3269);
nor U7427 (N_7427,N_3920,N_3197);
or U7428 (N_7428,N_519,N_3922);
nor U7429 (N_7429,N_2170,N_4608);
xor U7430 (N_7430,N_2237,N_2214);
and U7431 (N_7431,N_3533,N_2017);
and U7432 (N_7432,N_2026,N_1026);
nor U7433 (N_7433,N_1055,N_2932);
nor U7434 (N_7434,N_3610,N_985);
and U7435 (N_7435,N_827,N_3226);
or U7436 (N_7436,N_1930,N_4405);
nand U7437 (N_7437,N_2795,N_4421);
and U7438 (N_7438,N_3950,N_4243);
or U7439 (N_7439,N_2264,N_570);
or U7440 (N_7440,N_1758,N_1200);
and U7441 (N_7441,N_1241,N_892);
and U7442 (N_7442,N_1540,N_3186);
or U7443 (N_7443,N_768,N_1299);
nor U7444 (N_7444,N_881,N_219);
nand U7445 (N_7445,N_901,N_2202);
and U7446 (N_7446,N_925,N_2946);
and U7447 (N_7447,N_2365,N_702);
nand U7448 (N_7448,N_3264,N_2079);
and U7449 (N_7449,N_4559,N_3942);
nor U7450 (N_7450,N_2142,N_2613);
nand U7451 (N_7451,N_2551,N_4567);
or U7452 (N_7452,N_2001,N_1147);
or U7453 (N_7453,N_753,N_3572);
and U7454 (N_7454,N_1430,N_1784);
xor U7455 (N_7455,N_199,N_4672);
and U7456 (N_7456,N_1821,N_2496);
and U7457 (N_7457,N_1204,N_1979);
xnor U7458 (N_7458,N_3198,N_3825);
or U7459 (N_7459,N_998,N_2601);
nor U7460 (N_7460,N_3157,N_100);
or U7461 (N_7461,N_496,N_1968);
or U7462 (N_7462,N_1593,N_882);
and U7463 (N_7463,N_2002,N_2023);
nor U7464 (N_7464,N_2701,N_1864);
nand U7465 (N_7465,N_1803,N_4414);
nor U7466 (N_7466,N_4643,N_3117);
xor U7467 (N_7467,N_3984,N_1480);
nand U7468 (N_7468,N_4223,N_2925);
nor U7469 (N_7469,N_1888,N_4636);
and U7470 (N_7470,N_1317,N_4857);
nor U7471 (N_7471,N_3432,N_4479);
and U7472 (N_7472,N_2736,N_846);
and U7473 (N_7473,N_1880,N_329);
nor U7474 (N_7474,N_4184,N_3131);
nand U7475 (N_7475,N_3258,N_1806);
or U7476 (N_7476,N_2949,N_2115);
and U7477 (N_7477,N_3712,N_2985);
nor U7478 (N_7478,N_641,N_4582);
or U7479 (N_7479,N_3785,N_3472);
xor U7480 (N_7480,N_1021,N_2646);
nand U7481 (N_7481,N_304,N_838);
and U7482 (N_7482,N_2013,N_4227);
xor U7483 (N_7483,N_1024,N_728);
and U7484 (N_7484,N_2859,N_1773);
or U7485 (N_7485,N_2738,N_1778);
nand U7486 (N_7486,N_1341,N_2722);
or U7487 (N_7487,N_4546,N_1926);
and U7488 (N_7488,N_527,N_1291);
nand U7489 (N_7489,N_251,N_4467);
or U7490 (N_7490,N_2200,N_1156);
and U7491 (N_7491,N_475,N_4925);
and U7492 (N_7492,N_2503,N_1045);
or U7493 (N_7493,N_2799,N_3632);
and U7494 (N_7494,N_2812,N_290);
and U7495 (N_7495,N_4490,N_2293);
or U7496 (N_7496,N_4659,N_918);
xnor U7497 (N_7497,N_653,N_1724);
nand U7498 (N_7498,N_4096,N_3631);
or U7499 (N_7499,N_2837,N_1771);
and U7500 (N_7500,N_476,N_2988);
and U7501 (N_7501,N_138,N_3882);
nand U7502 (N_7502,N_3118,N_2368);
nand U7503 (N_7503,N_1627,N_1332);
nor U7504 (N_7504,N_4068,N_2742);
or U7505 (N_7505,N_3141,N_4823);
or U7506 (N_7506,N_3055,N_921);
or U7507 (N_7507,N_3398,N_4818);
and U7508 (N_7508,N_2298,N_4449);
nor U7509 (N_7509,N_2975,N_332);
or U7510 (N_7510,N_2803,N_2064);
xnor U7511 (N_7511,N_603,N_4408);
nor U7512 (N_7512,N_534,N_2639);
nand U7513 (N_7513,N_476,N_1027);
nand U7514 (N_7514,N_3853,N_3695);
xnor U7515 (N_7515,N_716,N_2469);
or U7516 (N_7516,N_1373,N_4182);
or U7517 (N_7517,N_801,N_4634);
and U7518 (N_7518,N_1570,N_3289);
or U7519 (N_7519,N_3852,N_2542);
or U7520 (N_7520,N_741,N_3955);
or U7521 (N_7521,N_1224,N_91);
nor U7522 (N_7522,N_2286,N_2812);
or U7523 (N_7523,N_2086,N_2541);
or U7524 (N_7524,N_2572,N_256);
or U7525 (N_7525,N_350,N_4877);
or U7526 (N_7526,N_935,N_2380);
nand U7527 (N_7527,N_933,N_6);
and U7528 (N_7528,N_3504,N_1633);
nand U7529 (N_7529,N_1278,N_4785);
or U7530 (N_7530,N_1261,N_3231);
or U7531 (N_7531,N_3203,N_3147);
xor U7532 (N_7532,N_3983,N_2723);
and U7533 (N_7533,N_4770,N_4434);
or U7534 (N_7534,N_1136,N_135);
nor U7535 (N_7535,N_1767,N_429);
and U7536 (N_7536,N_1798,N_3859);
and U7537 (N_7537,N_1475,N_883);
or U7538 (N_7538,N_3704,N_4025);
or U7539 (N_7539,N_2085,N_200);
xnor U7540 (N_7540,N_2625,N_2973);
and U7541 (N_7541,N_2061,N_1965);
nor U7542 (N_7542,N_1217,N_4139);
and U7543 (N_7543,N_4948,N_1815);
and U7544 (N_7544,N_4760,N_116);
nand U7545 (N_7545,N_2683,N_703);
nor U7546 (N_7546,N_1851,N_4306);
nand U7547 (N_7547,N_2033,N_2864);
nor U7548 (N_7548,N_3109,N_962);
and U7549 (N_7549,N_1273,N_3208);
xor U7550 (N_7550,N_1255,N_16);
nand U7551 (N_7551,N_1452,N_3942);
and U7552 (N_7552,N_1613,N_4899);
and U7553 (N_7553,N_4190,N_2459);
and U7554 (N_7554,N_4210,N_361);
xor U7555 (N_7555,N_2420,N_2137);
and U7556 (N_7556,N_815,N_2801);
nand U7557 (N_7557,N_1454,N_1133);
nor U7558 (N_7558,N_82,N_3757);
or U7559 (N_7559,N_1157,N_100);
and U7560 (N_7560,N_295,N_101);
nand U7561 (N_7561,N_1627,N_3174);
nand U7562 (N_7562,N_3743,N_1573);
and U7563 (N_7563,N_642,N_3879);
nor U7564 (N_7564,N_201,N_3705);
or U7565 (N_7565,N_1525,N_538);
nand U7566 (N_7566,N_4817,N_2418);
nor U7567 (N_7567,N_4591,N_2457);
or U7568 (N_7568,N_286,N_1341);
or U7569 (N_7569,N_4591,N_3030);
xor U7570 (N_7570,N_2382,N_1500);
and U7571 (N_7571,N_4260,N_459);
or U7572 (N_7572,N_4952,N_834);
nor U7573 (N_7573,N_4748,N_3757);
nand U7574 (N_7574,N_1708,N_1035);
nor U7575 (N_7575,N_3331,N_1602);
nor U7576 (N_7576,N_3707,N_1200);
nand U7577 (N_7577,N_2186,N_1679);
and U7578 (N_7578,N_1607,N_1816);
nand U7579 (N_7579,N_127,N_2195);
and U7580 (N_7580,N_4866,N_2078);
xnor U7581 (N_7581,N_3588,N_4060);
xor U7582 (N_7582,N_242,N_2160);
or U7583 (N_7583,N_4247,N_477);
nand U7584 (N_7584,N_4855,N_4427);
xor U7585 (N_7585,N_3781,N_3830);
or U7586 (N_7586,N_4877,N_1834);
xnor U7587 (N_7587,N_417,N_3588);
nand U7588 (N_7588,N_3440,N_2421);
or U7589 (N_7589,N_1183,N_2038);
nand U7590 (N_7590,N_2841,N_4230);
and U7591 (N_7591,N_4483,N_84);
nand U7592 (N_7592,N_743,N_3552);
or U7593 (N_7593,N_1991,N_535);
and U7594 (N_7594,N_4710,N_4085);
or U7595 (N_7595,N_808,N_90);
and U7596 (N_7596,N_1193,N_2045);
nor U7597 (N_7597,N_2555,N_1637);
or U7598 (N_7598,N_2490,N_2071);
and U7599 (N_7599,N_320,N_1519);
nand U7600 (N_7600,N_5,N_1367);
nand U7601 (N_7601,N_3506,N_827);
xor U7602 (N_7602,N_4112,N_3680);
nor U7603 (N_7603,N_1684,N_3049);
or U7604 (N_7604,N_4515,N_3253);
and U7605 (N_7605,N_2041,N_1587);
and U7606 (N_7606,N_3305,N_2061);
or U7607 (N_7607,N_4734,N_1480);
nand U7608 (N_7608,N_4649,N_3985);
nand U7609 (N_7609,N_2387,N_3625);
xnor U7610 (N_7610,N_4967,N_630);
or U7611 (N_7611,N_3709,N_1845);
and U7612 (N_7612,N_4314,N_2917);
and U7613 (N_7613,N_868,N_4259);
nor U7614 (N_7614,N_890,N_2809);
or U7615 (N_7615,N_4686,N_1267);
nor U7616 (N_7616,N_4828,N_3717);
xor U7617 (N_7617,N_2512,N_4106);
and U7618 (N_7618,N_2768,N_4312);
nand U7619 (N_7619,N_4555,N_4747);
nor U7620 (N_7620,N_4796,N_2402);
nand U7621 (N_7621,N_2540,N_95);
or U7622 (N_7622,N_3929,N_4248);
xor U7623 (N_7623,N_45,N_3649);
nor U7624 (N_7624,N_767,N_1062);
nand U7625 (N_7625,N_816,N_3552);
nor U7626 (N_7626,N_1594,N_3973);
and U7627 (N_7627,N_4587,N_4868);
or U7628 (N_7628,N_95,N_4759);
nand U7629 (N_7629,N_2513,N_295);
and U7630 (N_7630,N_271,N_336);
or U7631 (N_7631,N_4954,N_4253);
nor U7632 (N_7632,N_3018,N_9);
or U7633 (N_7633,N_3819,N_1886);
or U7634 (N_7634,N_2750,N_3945);
nor U7635 (N_7635,N_4425,N_4978);
xor U7636 (N_7636,N_1471,N_2377);
nand U7637 (N_7637,N_3703,N_573);
xnor U7638 (N_7638,N_466,N_1759);
nor U7639 (N_7639,N_2022,N_1661);
or U7640 (N_7640,N_3177,N_1634);
nand U7641 (N_7641,N_236,N_4174);
or U7642 (N_7642,N_2704,N_2753);
and U7643 (N_7643,N_291,N_1350);
nor U7644 (N_7644,N_1732,N_256);
or U7645 (N_7645,N_544,N_3390);
and U7646 (N_7646,N_805,N_1575);
and U7647 (N_7647,N_1477,N_168);
or U7648 (N_7648,N_2041,N_1117);
or U7649 (N_7649,N_2989,N_3504);
or U7650 (N_7650,N_1335,N_2795);
nor U7651 (N_7651,N_1084,N_1847);
and U7652 (N_7652,N_4129,N_332);
and U7653 (N_7653,N_2270,N_4373);
nand U7654 (N_7654,N_683,N_3019);
or U7655 (N_7655,N_2671,N_4333);
or U7656 (N_7656,N_862,N_2275);
nor U7657 (N_7657,N_1901,N_4046);
nor U7658 (N_7658,N_829,N_4596);
or U7659 (N_7659,N_534,N_1761);
nand U7660 (N_7660,N_2785,N_1995);
or U7661 (N_7661,N_4841,N_3257);
nor U7662 (N_7662,N_306,N_1202);
nor U7663 (N_7663,N_3316,N_4587);
nand U7664 (N_7664,N_2388,N_4325);
nand U7665 (N_7665,N_974,N_2197);
or U7666 (N_7666,N_382,N_3765);
or U7667 (N_7667,N_3732,N_2443);
nor U7668 (N_7668,N_811,N_260);
xor U7669 (N_7669,N_1514,N_2885);
nand U7670 (N_7670,N_4908,N_167);
and U7671 (N_7671,N_2649,N_2195);
or U7672 (N_7672,N_4692,N_2842);
nor U7673 (N_7673,N_4704,N_3824);
nor U7674 (N_7674,N_2098,N_414);
and U7675 (N_7675,N_4065,N_2287);
or U7676 (N_7676,N_4467,N_1260);
nor U7677 (N_7677,N_478,N_768);
or U7678 (N_7678,N_1366,N_127);
nor U7679 (N_7679,N_2644,N_323);
xor U7680 (N_7680,N_4242,N_4098);
nand U7681 (N_7681,N_3820,N_2016);
and U7682 (N_7682,N_1484,N_4236);
and U7683 (N_7683,N_4439,N_297);
nand U7684 (N_7684,N_2492,N_3829);
xnor U7685 (N_7685,N_1605,N_4217);
or U7686 (N_7686,N_2490,N_300);
or U7687 (N_7687,N_1393,N_3643);
nand U7688 (N_7688,N_181,N_3878);
nor U7689 (N_7689,N_3218,N_1735);
or U7690 (N_7690,N_3989,N_607);
xnor U7691 (N_7691,N_367,N_1259);
nor U7692 (N_7692,N_4050,N_1421);
nand U7693 (N_7693,N_602,N_1765);
nand U7694 (N_7694,N_339,N_609);
or U7695 (N_7695,N_1866,N_3658);
or U7696 (N_7696,N_2734,N_4798);
xnor U7697 (N_7697,N_2973,N_4451);
nor U7698 (N_7698,N_3400,N_4718);
and U7699 (N_7699,N_1737,N_162);
nor U7700 (N_7700,N_777,N_3463);
nand U7701 (N_7701,N_3353,N_4398);
xor U7702 (N_7702,N_986,N_931);
and U7703 (N_7703,N_1849,N_1823);
nand U7704 (N_7704,N_3847,N_2396);
nor U7705 (N_7705,N_601,N_4567);
nand U7706 (N_7706,N_3392,N_1059);
or U7707 (N_7707,N_3351,N_3641);
or U7708 (N_7708,N_2885,N_4581);
nand U7709 (N_7709,N_4630,N_3448);
nor U7710 (N_7710,N_3156,N_2083);
nor U7711 (N_7711,N_2271,N_727);
nor U7712 (N_7712,N_3683,N_1560);
nand U7713 (N_7713,N_4136,N_872);
nand U7714 (N_7714,N_3041,N_3575);
or U7715 (N_7715,N_1952,N_1116);
or U7716 (N_7716,N_2187,N_1951);
or U7717 (N_7717,N_4118,N_2053);
nand U7718 (N_7718,N_937,N_2189);
nor U7719 (N_7719,N_1347,N_4592);
xnor U7720 (N_7720,N_4689,N_2676);
or U7721 (N_7721,N_2280,N_4063);
nand U7722 (N_7722,N_3928,N_4778);
or U7723 (N_7723,N_4355,N_4400);
and U7724 (N_7724,N_3765,N_4310);
nor U7725 (N_7725,N_4389,N_583);
nand U7726 (N_7726,N_4631,N_2575);
nand U7727 (N_7727,N_4020,N_23);
nand U7728 (N_7728,N_1460,N_3368);
xor U7729 (N_7729,N_444,N_1500);
nor U7730 (N_7730,N_57,N_2715);
and U7731 (N_7731,N_1026,N_154);
and U7732 (N_7732,N_3757,N_3125);
nand U7733 (N_7733,N_2695,N_1346);
and U7734 (N_7734,N_1365,N_510);
nand U7735 (N_7735,N_4533,N_4650);
nand U7736 (N_7736,N_4189,N_4804);
and U7737 (N_7737,N_4238,N_2570);
and U7738 (N_7738,N_4196,N_4265);
nor U7739 (N_7739,N_4029,N_2255);
nand U7740 (N_7740,N_1159,N_1297);
xor U7741 (N_7741,N_3124,N_1441);
nand U7742 (N_7742,N_1365,N_4483);
or U7743 (N_7743,N_4276,N_4521);
nand U7744 (N_7744,N_4724,N_2749);
xnor U7745 (N_7745,N_847,N_4845);
or U7746 (N_7746,N_2113,N_4545);
and U7747 (N_7747,N_2989,N_617);
nor U7748 (N_7748,N_3955,N_69);
xor U7749 (N_7749,N_4398,N_280);
nand U7750 (N_7750,N_2028,N_1671);
and U7751 (N_7751,N_3708,N_4317);
or U7752 (N_7752,N_386,N_4328);
or U7753 (N_7753,N_1847,N_4757);
nor U7754 (N_7754,N_2956,N_2733);
nand U7755 (N_7755,N_1623,N_645);
or U7756 (N_7756,N_4976,N_2924);
nor U7757 (N_7757,N_1250,N_4197);
and U7758 (N_7758,N_3144,N_4098);
nand U7759 (N_7759,N_898,N_3196);
nor U7760 (N_7760,N_1382,N_2708);
and U7761 (N_7761,N_2078,N_4915);
nand U7762 (N_7762,N_2479,N_2138);
xor U7763 (N_7763,N_1849,N_1327);
nor U7764 (N_7764,N_2103,N_2588);
and U7765 (N_7765,N_3497,N_288);
or U7766 (N_7766,N_59,N_707);
nand U7767 (N_7767,N_1630,N_2532);
and U7768 (N_7768,N_4560,N_1955);
or U7769 (N_7769,N_4899,N_1100);
nand U7770 (N_7770,N_2127,N_1456);
and U7771 (N_7771,N_2820,N_4902);
nand U7772 (N_7772,N_2201,N_2791);
or U7773 (N_7773,N_3052,N_638);
xnor U7774 (N_7774,N_4973,N_524);
xnor U7775 (N_7775,N_3161,N_2482);
nand U7776 (N_7776,N_4636,N_2708);
nand U7777 (N_7777,N_4903,N_2466);
nand U7778 (N_7778,N_4332,N_4782);
and U7779 (N_7779,N_4246,N_706);
or U7780 (N_7780,N_943,N_3407);
and U7781 (N_7781,N_1988,N_691);
and U7782 (N_7782,N_1717,N_1217);
nand U7783 (N_7783,N_4510,N_4478);
and U7784 (N_7784,N_2575,N_4346);
xnor U7785 (N_7785,N_466,N_2838);
nor U7786 (N_7786,N_4206,N_860);
or U7787 (N_7787,N_3306,N_614);
and U7788 (N_7788,N_4105,N_1645);
nor U7789 (N_7789,N_3895,N_4761);
xor U7790 (N_7790,N_1197,N_1355);
and U7791 (N_7791,N_4833,N_4600);
and U7792 (N_7792,N_3272,N_4614);
and U7793 (N_7793,N_3692,N_3956);
nor U7794 (N_7794,N_288,N_110);
and U7795 (N_7795,N_768,N_1695);
xnor U7796 (N_7796,N_4247,N_886);
nand U7797 (N_7797,N_1181,N_510);
nor U7798 (N_7798,N_3337,N_1461);
or U7799 (N_7799,N_4544,N_4581);
nand U7800 (N_7800,N_2792,N_3532);
and U7801 (N_7801,N_1372,N_4540);
and U7802 (N_7802,N_749,N_1721);
and U7803 (N_7803,N_3503,N_2219);
nor U7804 (N_7804,N_1456,N_663);
nand U7805 (N_7805,N_3269,N_1159);
nand U7806 (N_7806,N_368,N_406);
nor U7807 (N_7807,N_4311,N_2126);
or U7808 (N_7808,N_4147,N_1572);
nand U7809 (N_7809,N_853,N_2346);
or U7810 (N_7810,N_138,N_327);
or U7811 (N_7811,N_2496,N_1559);
or U7812 (N_7812,N_2250,N_2827);
nand U7813 (N_7813,N_2716,N_1091);
nand U7814 (N_7814,N_2128,N_2479);
nand U7815 (N_7815,N_4831,N_3858);
and U7816 (N_7816,N_787,N_2637);
nor U7817 (N_7817,N_3937,N_2074);
or U7818 (N_7818,N_299,N_4687);
and U7819 (N_7819,N_2848,N_1962);
xor U7820 (N_7820,N_1738,N_4879);
nor U7821 (N_7821,N_2241,N_1018);
and U7822 (N_7822,N_2046,N_3388);
nor U7823 (N_7823,N_1090,N_4496);
or U7824 (N_7824,N_3710,N_2150);
nor U7825 (N_7825,N_4551,N_3179);
nor U7826 (N_7826,N_3378,N_446);
and U7827 (N_7827,N_2576,N_4648);
nand U7828 (N_7828,N_682,N_3586);
xnor U7829 (N_7829,N_2835,N_4765);
nand U7830 (N_7830,N_742,N_3931);
or U7831 (N_7831,N_818,N_3856);
or U7832 (N_7832,N_2012,N_2407);
nor U7833 (N_7833,N_2363,N_614);
nor U7834 (N_7834,N_1526,N_3246);
and U7835 (N_7835,N_1687,N_626);
or U7836 (N_7836,N_2634,N_3711);
nand U7837 (N_7837,N_2922,N_3106);
and U7838 (N_7838,N_932,N_3280);
nor U7839 (N_7839,N_2774,N_4884);
or U7840 (N_7840,N_4451,N_2128);
nand U7841 (N_7841,N_1538,N_828);
nand U7842 (N_7842,N_3756,N_4753);
xor U7843 (N_7843,N_2638,N_4818);
xor U7844 (N_7844,N_2216,N_1932);
nor U7845 (N_7845,N_1317,N_3236);
and U7846 (N_7846,N_1687,N_1690);
nand U7847 (N_7847,N_2488,N_4380);
nand U7848 (N_7848,N_4442,N_4414);
nor U7849 (N_7849,N_4449,N_2159);
and U7850 (N_7850,N_111,N_2159);
and U7851 (N_7851,N_1773,N_4612);
nand U7852 (N_7852,N_498,N_2134);
nand U7853 (N_7853,N_1968,N_4669);
nor U7854 (N_7854,N_1159,N_4874);
xor U7855 (N_7855,N_3323,N_2712);
or U7856 (N_7856,N_3112,N_2806);
xnor U7857 (N_7857,N_1287,N_645);
nand U7858 (N_7858,N_4925,N_3885);
or U7859 (N_7859,N_3221,N_544);
or U7860 (N_7860,N_3142,N_129);
and U7861 (N_7861,N_168,N_4890);
or U7862 (N_7862,N_2363,N_671);
and U7863 (N_7863,N_199,N_223);
and U7864 (N_7864,N_4648,N_1872);
and U7865 (N_7865,N_1319,N_3552);
and U7866 (N_7866,N_2248,N_3778);
nand U7867 (N_7867,N_2852,N_1981);
nor U7868 (N_7868,N_4586,N_1770);
and U7869 (N_7869,N_4453,N_52);
or U7870 (N_7870,N_3206,N_4659);
nand U7871 (N_7871,N_342,N_942);
and U7872 (N_7872,N_1150,N_2202);
nand U7873 (N_7873,N_2986,N_2506);
xor U7874 (N_7874,N_2739,N_66);
nor U7875 (N_7875,N_2080,N_4841);
and U7876 (N_7876,N_3409,N_1654);
or U7877 (N_7877,N_4396,N_2986);
nand U7878 (N_7878,N_2088,N_2641);
nor U7879 (N_7879,N_3470,N_132);
or U7880 (N_7880,N_1533,N_3686);
nand U7881 (N_7881,N_777,N_2155);
or U7882 (N_7882,N_445,N_1265);
xnor U7883 (N_7883,N_3917,N_617);
nor U7884 (N_7884,N_4510,N_796);
and U7885 (N_7885,N_1269,N_2039);
xnor U7886 (N_7886,N_52,N_561);
nor U7887 (N_7887,N_4014,N_2274);
nand U7888 (N_7888,N_85,N_4309);
or U7889 (N_7889,N_1100,N_1920);
nand U7890 (N_7890,N_3157,N_1040);
nand U7891 (N_7891,N_1230,N_4745);
and U7892 (N_7892,N_4199,N_2489);
nor U7893 (N_7893,N_3188,N_447);
nand U7894 (N_7894,N_3430,N_224);
nor U7895 (N_7895,N_2332,N_762);
nand U7896 (N_7896,N_3508,N_3499);
and U7897 (N_7897,N_406,N_4619);
or U7898 (N_7898,N_4263,N_3575);
or U7899 (N_7899,N_1701,N_484);
nand U7900 (N_7900,N_2601,N_2050);
or U7901 (N_7901,N_4713,N_4439);
nand U7902 (N_7902,N_1535,N_4841);
or U7903 (N_7903,N_3073,N_3230);
nand U7904 (N_7904,N_1054,N_617);
and U7905 (N_7905,N_2075,N_2452);
nor U7906 (N_7906,N_1457,N_3495);
nand U7907 (N_7907,N_262,N_4921);
or U7908 (N_7908,N_67,N_3423);
nor U7909 (N_7909,N_1995,N_310);
xor U7910 (N_7910,N_3515,N_635);
and U7911 (N_7911,N_305,N_2517);
nor U7912 (N_7912,N_4017,N_2949);
nand U7913 (N_7913,N_3250,N_2278);
or U7914 (N_7914,N_4209,N_1699);
xor U7915 (N_7915,N_4238,N_165);
and U7916 (N_7916,N_287,N_2191);
or U7917 (N_7917,N_2880,N_4124);
nor U7918 (N_7918,N_3705,N_1512);
nand U7919 (N_7919,N_1634,N_4791);
xor U7920 (N_7920,N_1888,N_3079);
nand U7921 (N_7921,N_467,N_3065);
nor U7922 (N_7922,N_2016,N_3349);
xor U7923 (N_7923,N_4404,N_4910);
or U7924 (N_7924,N_2101,N_887);
or U7925 (N_7925,N_2632,N_4524);
and U7926 (N_7926,N_4529,N_1911);
and U7927 (N_7927,N_4225,N_2550);
nor U7928 (N_7928,N_3763,N_4593);
nand U7929 (N_7929,N_1043,N_4406);
nand U7930 (N_7930,N_3919,N_4069);
and U7931 (N_7931,N_3876,N_684);
and U7932 (N_7932,N_633,N_990);
and U7933 (N_7933,N_850,N_1945);
nor U7934 (N_7934,N_1621,N_4877);
and U7935 (N_7935,N_4159,N_3695);
nand U7936 (N_7936,N_84,N_2641);
xor U7937 (N_7937,N_1985,N_1705);
or U7938 (N_7938,N_437,N_2641);
or U7939 (N_7939,N_3500,N_4339);
and U7940 (N_7940,N_2291,N_4650);
xnor U7941 (N_7941,N_3019,N_743);
xor U7942 (N_7942,N_1977,N_3774);
nor U7943 (N_7943,N_1959,N_2864);
and U7944 (N_7944,N_220,N_3171);
or U7945 (N_7945,N_2203,N_4707);
nand U7946 (N_7946,N_1320,N_4305);
or U7947 (N_7947,N_1385,N_673);
nand U7948 (N_7948,N_332,N_2340);
nand U7949 (N_7949,N_4556,N_548);
nor U7950 (N_7950,N_3963,N_1736);
nand U7951 (N_7951,N_4496,N_366);
nand U7952 (N_7952,N_3604,N_4643);
and U7953 (N_7953,N_1184,N_3037);
and U7954 (N_7954,N_1764,N_2639);
nand U7955 (N_7955,N_1285,N_280);
or U7956 (N_7956,N_2565,N_3280);
nand U7957 (N_7957,N_3327,N_1309);
and U7958 (N_7958,N_3816,N_867);
nand U7959 (N_7959,N_1993,N_3888);
nor U7960 (N_7960,N_3304,N_753);
and U7961 (N_7961,N_4680,N_3013);
or U7962 (N_7962,N_773,N_2229);
nand U7963 (N_7963,N_4657,N_4166);
or U7964 (N_7964,N_2772,N_2049);
nand U7965 (N_7965,N_1694,N_1887);
or U7966 (N_7966,N_1339,N_2258);
nor U7967 (N_7967,N_1857,N_4887);
nand U7968 (N_7968,N_2059,N_4332);
nand U7969 (N_7969,N_4681,N_1215);
nand U7970 (N_7970,N_1046,N_4080);
nand U7971 (N_7971,N_4286,N_4868);
or U7972 (N_7972,N_472,N_1876);
nand U7973 (N_7973,N_2422,N_4163);
and U7974 (N_7974,N_323,N_3172);
nand U7975 (N_7975,N_1781,N_283);
and U7976 (N_7976,N_3071,N_1657);
or U7977 (N_7977,N_2718,N_1359);
nor U7978 (N_7978,N_4617,N_3299);
or U7979 (N_7979,N_3318,N_3757);
or U7980 (N_7980,N_4750,N_3994);
xor U7981 (N_7981,N_1679,N_461);
or U7982 (N_7982,N_944,N_2777);
and U7983 (N_7983,N_4778,N_437);
or U7984 (N_7984,N_4864,N_1680);
and U7985 (N_7985,N_2695,N_318);
nor U7986 (N_7986,N_4350,N_2405);
nand U7987 (N_7987,N_3522,N_691);
or U7988 (N_7988,N_829,N_1113);
nor U7989 (N_7989,N_3077,N_1862);
xor U7990 (N_7990,N_4215,N_242);
nand U7991 (N_7991,N_1893,N_4206);
and U7992 (N_7992,N_1761,N_3368);
nand U7993 (N_7993,N_378,N_3902);
nor U7994 (N_7994,N_3514,N_3970);
nand U7995 (N_7995,N_2853,N_4741);
or U7996 (N_7996,N_1700,N_2249);
nor U7997 (N_7997,N_4000,N_177);
nand U7998 (N_7998,N_3606,N_2134);
nand U7999 (N_7999,N_920,N_4995);
nand U8000 (N_8000,N_3390,N_785);
nand U8001 (N_8001,N_4811,N_4125);
or U8002 (N_8002,N_3899,N_4877);
nor U8003 (N_8003,N_728,N_4923);
or U8004 (N_8004,N_2215,N_4733);
or U8005 (N_8005,N_104,N_2979);
and U8006 (N_8006,N_721,N_4897);
and U8007 (N_8007,N_4008,N_825);
and U8008 (N_8008,N_3194,N_4818);
nor U8009 (N_8009,N_227,N_1458);
nand U8010 (N_8010,N_3049,N_231);
or U8011 (N_8011,N_1304,N_3666);
and U8012 (N_8012,N_4096,N_1273);
and U8013 (N_8013,N_3142,N_4974);
and U8014 (N_8014,N_1945,N_594);
nand U8015 (N_8015,N_2331,N_4806);
and U8016 (N_8016,N_1172,N_2455);
and U8017 (N_8017,N_3064,N_1351);
nand U8018 (N_8018,N_1748,N_866);
nand U8019 (N_8019,N_4383,N_4728);
or U8020 (N_8020,N_1312,N_2875);
or U8021 (N_8021,N_780,N_1227);
and U8022 (N_8022,N_4340,N_3163);
xnor U8023 (N_8023,N_1370,N_1523);
xor U8024 (N_8024,N_420,N_786);
nor U8025 (N_8025,N_2960,N_4364);
nor U8026 (N_8026,N_3606,N_4662);
or U8027 (N_8027,N_1339,N_4615);
nor U8028 (N_8028,N_2056,N_1148);
nor U8029 (N_8029,N_1305,N_1439);
nor U8030 (N_8030,N_4855,N_793);
nand U8031 (N_8031,N_4149,N_1478);
xnor U8032 (N_8032,N_1345,N_2413);
nor U8033 (N_8033,N_2043,N_341);
and U8034 (N_8034,N_3614,N_3397);
or U8035 (N_8035,N_375,N_161);
or U8036 (N_8036,N_2884,N_4671);
xor U8037 (N_8037,N_2956,N_4348);
nand U8038 (N_8038,N_2642,N_297);
nand U8039 (N_8039,N_2503,N_4674);
or U8040 (N_8040,N_688,N_2796);
and U8041 (N_8041,N_3893,N_1367);
and U8042 (N_8042,N_404,N_4663);
nand U8043 (N_8043,N_2096,N_130);
or U8044 (N_8044,N_2367,N_2119);
xnor U8045 (N_8045,N_1884,N_3706);
or U8046 (N_8046,N_1300,N_1006);
nor U8047 (N_8047,N_1252,N_4729);
nor U8048 (N_8048,N_808,N_754);
and U8049 (N_8049,N_3703,N_3704);
nor U8050 (N_8050,N_3854,N_4754);
nand U8051 (N_8051,N_3713,N_2481);
and U8052 (N_8052,N_3452,N_2182);
and U8053 (N_8053,N_2197,N_4926);
or U8054 (N_8054,N_1722,N_1100);
nor U8055 (N_8055,N_396,N_1843);
or U8056 (N_8056,N_2128,N_183);
nand U8057 (N_8057,N_503,N_2881);
and U8058 (N_8058,N_3177,N_4499);
nand U8059 (N_8059,N_1249,N_3139);
nand U8060 (N_8060,N_1193,N_507);
nor U8061 (N_8061,N_1131,N_3018);
or U8062 (N_8062,N_4154,N_2029);
nand U8063 (N_8063,N_1722,N_1950);
and U8064 (N_8064,N_4029,N_1327);
and U8065 (N_8065,N_2956,N_4113);
nor U8066 (N_8066,N_1959,N_2576);
or U8067 (N_8067,N_289,N_4496);
nand U8068 (N_8068,N_807,N_1460);
nand U8069 (N_8069,N_382,N_1092);
and U8070 (N_8070,N_3940,N_2912);
and U8071 (N_8071,N_3854,N_4160);
and U8072 (N_8072,N_566,N_1697);
and U8073 (N_8073,N_2925,N_4353);
and U8074 (N_8074,N_1171,N_1298);
and U8075 (N_8075,N_3761,N_336);
or U8076 (N_8076,N_1244,N_1080);
nand U8077 (N_8077,N_387,N_2024);
xnor U8078 (N_8078,N_1235,N_3886);
or U8079 (N_8079,N_2204,N_1660);
xor U8080 (N_8080,N_901,N_2149);
and U8081 (N_8081,N_3983,N_1096);
nor U8082 (N_8082,N_1787,N_361);
or U8083 (N_8083,N_4422,N_2982);
nor U8084 (N_8084,N_1149,N_2050);
and U8085 (N_8085,N_117,N_1383);
and U8086 (N_8086,N_53,N_3501);
nor U8087 (N_8087,N_3241,N_1886);
or U8088 (N_8088,N_2509,N_4315);
xor U8089 (N_8089,N_127,N_626);
nor U8090 (N_8090,N_644,N_1828);
nor U8091 (N_8091,N_2873,N_32);
nand U8092 (N_8092,N_1285,N_691);
or U8093 (N_8093,N_1550,N_1834);
xnor U8094 (N_8094,N_338,N_1345);
and U8095 (N_8095,N_294,N_609);
nand U8096 (N_8096,N_4894,N_3565);
nor U8097 (N_8097,N_1707,N_3028);
nor U8098 (N_8098,N_1013,N_2654);
and U8099 (N_8099,N_3729,N_4645);
nand U8100 (N_8100,N_3386,N_1502);
nor U8101 (N_8101,N_4234,N_4723);
and U8102 (N_8102,N_2816,N_1003);
nor U8103 (N_8103,N_2070,N_4824);
nor U8104 (N_8104,N_4264,N_4135);
xnor U8105 (N_8105,N_1560,N_25);
nand U8106 (N_8106,N_4158,N_4940);
and U8107 (N_8107,N_4117,N_4788);
nand U8108 (N_8108,N_1390,N_2219);
xor U8109 (N_8109,N_4982,N_1751);
and U8110 (N_8110,N_967,N_2684);
or U8111 (N_8111,N_4534,N_395);
xnor U8112 (N_8112,N_3211,N_4640);
nand U8113 (N_8113,N_3262,N_237);
and U8114 (N_8114,N_3215,N_273);
nand U8115 (N_8115,N_1277,N_767);
nor U8116 (N_8116,N_2424,N_2259);
or U8117 (N_8117,N_3859,N_4355);
nor U8118 (N_8118,N_352,N_4228);
nor U8119 (N_8119,N_4963,N_1176);
and U8120 (N_8120,N_2792,N_268);
and U8121 (N_8121,N_2188,N_227);
and U8122 (N_8122,N_1250,N_1597);
nor U8123 (N_8123,N_3307,N_1826);
nand U8124 (N_8124,N_401,N_3885);
or U8125 (N_8125,N_2064,N_679);
or U8126 (N_8126,N_61,N_567);
nand U8127 (N_8127,N_1139,N_4608);
nand U8128 (N_8128,N_744,N_2999);
and U8129 (N_8129,N_4504,N_2257);
xor U8130 (N_8130,N_21,N_2034);
nor U8131 (N_8131,N_1564,N_2594);
and U8132 (N_8132,N_3892,N_3568);
nand U8133 (N_8133,N_1103,N_329);
or U8134 (N_8134,N_3959,N_1951);
and U8135 (N_8135,N_2679,N_4071);
or U8136 (N_8136,N_1875,N_3962);
nand U8137 (N_8137,N_2320,N_3723);
nor U8138 (N_8138,N_4612,N_1579);
and U8139 (N_8139,N_3982,N_2195);
xnor U8140 (N_8140,N_4826,N_1548);
nor U8141 (N_8141,N_4606,N_4441);
xnor U8142 (N_8142,N_1488,N_3688);
and U8143 (N_8143,N_1435,N_806);
and U8144 (N_8144,N_100,N_2695);
nand U8145 (N_8145,N_3624,N_4819);
nand U8146 (N_8146,N_3939,N_3674);
nor U8147 (N_8147,N_2806,N_4674);
or U8148 (N_8148,N_1710,N_3521);
nor U8149 (N_8149,N_3867,N_1);
or U8150 (N_8150,N_4409,N_1841);
or U8151 (N_8151,N_1089,N_3771);
nor U8152 (N_8152,N_4918,N_4015);
nor U8153 (N_8153,N_1708,N_555);
and U8154 (N_8154,N_3914,N_8);
and U8155 (N_8155,N_4131,N_4830);
and U8156 (N_8156,N_3632,N_3841);
nor U8157 (N_8157,N_3633,N_1171);
nand U8158 (N_8158,N_1746,N_3048);
nand U8159 (N_8159,N_1995,N_3191);
and U8160 (N_8160,N_3984,N_4341);
and U8161 (N_8161,N_2349,N_3992);
nand U8162 (N_8162,N_462,N_2390);
and U8163 (N_8163,N_1875,N_3192);
nor U8164 (N_8164,N_3446,N_2431);
and U8165 (N_8165,N_3125,N_3662);
nand U8166 (N_8166,N_1854,N_1337);
nor U8167 (N_8167,N_1665,N_4292);
nor U8168 (N_8168,N_950,N_3996);
nor U8169 (N_8169,N_359,N_4950);
nor U8170 (N_8170,N_4736,N_294);
nand U8171 (N_8171,N_984,N_549);
or U8172 (N_8172,N_4030,N_2401);
nand U8173 (N_8173,N_2917,N_4484);
nor U8174 (N_8174,N_808,N_4341);
and U8175 (N_8175,N_2474,N_977);
and U8176 (N_8176,N_105,N_342);
xor U8177 (N_8177,N_1008,N_1909);
nand U8178 (N_8178,N_4105,N_153);
nor U8179 (N_8179,N_1798,N_4311);
and U8180 (N_8180,N_2620,N_2156);
and U8181 (N_8181,N_419,N_4501);
nor U8182 (N_8182,N_1163,N_3478);
and U8183 (N_8183,N_685,N_1089);
or U8184 (N_8184,N_3138,N_3098);
xor U8185 (N_8185,N_2024,N_3618);
xnor U8186 (N_8186,N_3627,N_2452);
nor U8187 (N_8187,N_3897,N_3924);
and U8188 (N_8188,N_2410,N_4300);
nand U8189 (N_8189,N_2328,N_1254);
xnor U8190 (N_8190,N_3839,N_2625);
nand U8191 (N_8191,N_1914,N_2701);
xnor U8192 (N_8192,N_2061,N_3251);
nor U8193 (N_8193,N_4683,N_237);
xnor U8194 (N_8194,N_817,N_4027);
nor U8195 (N_8195,N_1108,N_358);
xnor U8196 (N_8196,N_3745,N_2055);
nor U8197 (N_8197,N_2325,N_2243);
nand U8198 (N_8198,N_2590,N_2714);
or U8199 (N_8199,N_2369,N_1185);
or U8200 (N_8200,N_1401,N_4732);
nor U8201 (N_8201,N_2106,N_4031);
xor U8202 (N_8202,N_2339,N_358);
and U8203 (N_8203,N_4099,N_4506);
and U8204 (N_8204,N_1099,N_3192);
nand U8205 (N_8205,N_4894,N_2625);
xor U8206 (N_8206,N_3208,N_1260);
nor U8207 (N_8207,N_4802,N_999);
nand U8208 (N_8208,N_1550,N_467);
or U8209 (N_8209,N_568,N_2642);
nor U8210 (N_8210,N_2628,N_1367);
nor U8211 (N_8211,N_2524,N_274);
xor U8212 (N_8212,N_2333,N_3476);
and U8213 (N_8213,N_4823,N_1840);
and U8214 (N_8214,N_2885,N_1981);
and U8215 (N_8215,N_1138,N_2295);
or U8216 (N_8216,N_61,N_816);
and U8217 (N_8217,N_4479,N_1830);
and U8218 (N_8218,N_4924,N_2351);
nand U8219 (N_8219,N_4849,N_4463);
and U8220 (N_8220,N_1018,N_643);
nand U8221 (N_8221,N_4040,N_3013);
and U8222 (N_8222,N_2686,N_3380);
xnor U8223 (N_8223,N_41,N_676);
nor U8224 (N_8224,N_517,N_474);
and U8225 (N_8225,N_2999,N_4380);
xor U8226 (N_8226,N_4960,N_890);
and U8227 (N_8227,N_36,N_3155);
nor U8228 (N_8228,N_3182,N_4414);
or U8229 (N_8229,N_963,N_1134);
nor U8230 (N_8230,N_3553,N_4723);
nor U8231 (N_8231,N_3432,N_2746);
or U8232 (N_8232,N_874,N_3441);
nor U8233 (N_8233,N_3569,N_4379);
or U8234 (N_8234,N_2031,N_4288);
nand U8235 (N_8235,N_4814,N_2439);
and U8236 (N_8236,N_648,N_132);
nand U8237 (N_8237,N_1661,N_2080);
or U8238 (N_8238,N_4667,N_4961);
or U8239 (N_8239,N_386,N_1052);
nor U8240 (N_8240,N_4921,N_2636);
nand U8241 (N_8241,N_2621,N_675);
nor U8242 (N_8242,N_1017,N_545);
and U8243 (N_8243,N_4466,N_3710);
or U8244 (N_8244,N_2002,N_4000);
nand U8245 (N_8245,N_4685,N_2425);
nor U8246 (N_8246,N_1244,N_1369);
or U8247 (N_8247,N_917,N_1660);
xor U8248 (N_8248,N_1464,N_1435);
nand U8249 (N_8249,N_4801,N_3750);
nand U8250 (N_8250,N_4142,N_2333);
nand U8251 (N_8251,N_1986,N_3317);
or U8252 (N_8252,N_1021,N_4074);
nand U8253 (N_8253,N_4108,N_1878);
nand U8254 (N_8254,N_291,N_4607);
xor U8255 (N_8255,N_66,N_2767);
xor U8256 (N_8256,N_1625,N_2970);
nand U8257 (N_8257,N_4199,N_4758);
and U8258 (N_8258,N_3365,N_1792);
and U8259 (N_8259,N_3643,N_660);
nor U8260 (N_8260,N_1253,N_4627);
and U8261 (N_8261,N_17,N_3636);
and U8262 (N_8262,N_2501,N_2335);
or U8263 (N_8263,N_3980,N_4671);
and U8264 (N_8264,N_2578,N_2065);
xor U8265 (N_8265,N_3283,N_3);
or U8266 (N_8266,N_1377,N_3173);
nand U8267 (N_8267,N_252,N_2776);
and U8268 (N_8268,N_1594,N_803);
and U8269 (N_8269,N_1459,N_3647);
nor U8270 (N_8270,N_4922,N_3937);
xnor U8271 (N_8271,N_4901,N_4507);
nand U8272 (N_8272,N_4651,N_3084);
nor U8273 (N_8273,N_2551,N_2513);
and U8274 (N_8274,N_4850,N_3252);
nor U8275 (N_8275,N_3741,N_2600);
and U8276 (N_8276,N_2284,N_4197);
nand U8277 (N_8277,N_1944,N_3366);
and U8278 (N_8278,N_2884,N_4375);
and U8279 (N_8279,N_1650,N_1851);
nor U8280 (N_8280,N_2446,N_1406);
xnor U8281 (N_8281,N_1510,N_4191);
nor U8282 (N_8282,N_1338,N_3554);
and U8283 (N_8283,N_1281,N_746);
nand U8284 (N_8284,N_394,N_438);
and U8285 (N_8285,N_3883,N_1289);
and U8286 (N_8286,N_1620,N_713);
and U8287 (N_8287,N_1588,N_468);
or U8288 (N_8288,N_4055,N_1901);
nand U8289 (N_8289,N_3123,N_4997);
nand U8290 (N_8290,N_2641,N_3270);
nor U8291 (N_8291,N_345,N_2022);
and U8292 (N_8292,N_913,N_4230);
nand U8293 (N_8293,N_2179,N_4115);
nor U8294 (N_8294,N_133,N_4614);
or U8295 (N_8295,N_771,N_4789);
nor U8296 (N_8296,N_808,N_1642);
and U8297 (N_8297,N_2789,N_2613);
and U8298 (N_8298,N_691,N_4673);
and U8299 (N_8299,N_875,N_3061);
and U8300 (N_8300,N_3466,N_3235);
nand U8301 (N_8301,N_380,N_4379);
nor U8302 (N_8302,N_2959,N_4938);
nand U8303 (N_8303,N_4454,N_1090);
nor U8304 (N_8304,N_789,N_545);
nand U8305 (N_8305,N_2095,N_4590);
nand U8306 (N_8306,N_2260,N_3350);
nor U8307 (N_8307,N_3928,N_2078);
nor U8308 (N_8308,N_3761,N_213);
nand U8309 (N_8309,N_3598,N_3627);
or U8310 (N_8310,N_407,N_2605);
or U8311 (N_8311,N_155,N_4757);
and U8312 (N_8312,N_368,N_3490);
or U8313 (N_8313,N_2907,N_4446);
or U8314 (N_8314,N_3079,N_2855);
and U8315 (N_8315,N_715,N_1315);
or U8316 (N_8316,N_4638,N_3029);
or U8317 (N_8317,N_580,N_3925);
or U8318 (N_8318,N_1180,N_930);
or U8319 (N_8319,N_65,N_2928);
nand U8320 (N_8320,N_4818,N_3917);
nor U8321 (N_8321,N_1263,N_106);
nand U8322 (N_8322,N_2962,N_4153);
and U8323 (N_8323,N_251,N_222);
nor U8324 (N_8324,N_2517,N_4392);
nand U8325 (N_8325,N_4673,N_2057);
and U8326 (N_8326,N_3840,N_1306);
or U8327 (N_8327,N_22,N_3880);
or U8328 (N_8328,N_4439,N_2552);
and U8329 (N_8329,N_3953,N_1445);
and U8330 (N_8330,N_102,N_457);
nor U8331 (N_8331,N_1959,N_3801);
or U8332 (N_8332,N_3005,N_1970);
nor U8333 (N_8333,N_3783,N_2068);
and U8334 (N_8334,N_1572,N_272);
nand U8335 (N_8335,N_4279,N_397);
nor U8336 (N_8336,N_472,N_1937);
nor U8337 (N_8337,N_3629,N_2408);
nand U8338 (N_8338,N_4033,N_2734);
xnor U8339 (N_8339,N_1827,N_4714);
xnor U8340 (N_8340,N_3720,N_1804);
and U8341 (N_8341,N_2239,N_1839);
nor U8342 (N_8342,N_3303,N_3053);
nand U8343 (N_8343,N_4862,N_3383);
xnor U8344 (N_8344,N_4766,N_4040);
and U8345 (N_8345,N_4995,N_837);
and U8346 (N_8346,N_4899,N_4901);
or U8347 (N_8347,N_4806,N_874);
nor U8348 (N_8348,N_4591,N_3121);
or U8349 (N_8349,N_528,N_2281);
nor U8350 (N_8350,N_1331,N_3790);
nand U8351 (N_8351,N_2059,N_2394);
and U8352 (N_8352,N_616,N_211);
xnor U8353 (N_8353,N_1547,N_376);
and U8354 (N_8354,N_1776,N_3946);
nand U8355 (N_8355,N_4511,N_4303);
xor U8356 (N_8356,N_2739,N_4348);
nor U8357 (N_8357,N_933,N_2500);
nand U8358 (N_8358,N_3420,N_2120);
and U8359 (N_8359,N_737,N_210);
nor U8360 (N_8360,N_4959,N_4873);
and U8361 (N_8361,N_2585,N_3715);
and U8362 (N_8362,N_23,N_607);
or U8363 (N_8363,N_3895,N_4305);
nand U8364 (N_8364,N_2849,N_573);
and U8365 (N_8365,N_2867,N_947);
or U8366 (N_8366,N_3644,N_2776);
nand U8367 (N_8367,N_4129,N_975);
and U8368 (N_8368,N_321,N_2019);
and U8369 (N_8369,N_345,N_1685);
nor U8370 (N_8370,N_3423,N_1669);
nand U8371 (N_8371,N_1201,N_3774);
or U8372 (N_8372,N_4607,N_2176);
or U8373 (N_8373,N_885,N_3117);
or U8374 (N_8374,N_1227,N_3014);
nand U8375 (N_8375,N_1362,N_2325);
nor U8376 (N_8376,N_2628,N_1381);
nand U8377 (N_8377,N_1649,N_1607);
and U8378 (N_8378,N_847,N_600);
nor U8379 (N_8379,N_1389,N_396);
xnor U8380 (N_8380,N_3709,N_1552);
and U8381 (N_8381,N_3201,N_1488);
and U8382 (N_8382,N_4523,N_3498);
or U8383 (N_8383,N_3309,N_3372);
xor U8384 (N_8384,N_2772,N_4768);
or U8385 (N_8385,N_1788,N_599);
nor U8386 (N_8386,N_1445,N_184);
nor U8387 (N_8387,N_3518,N_622);
or U8388 (N_8388,N_2285,N_1423);
and U8389 (N_8389,N_2747,N_4463);
or U8390 (N_8390,N_3811,N_3790);
nor U8391 (N_8391,N_490,N_1810);
or U8392 (N_8392,N_1731,N_182);
nand U8393 (N_8393,N_1168,N_2478);
and U8394 (N_8394,N_1640,N_660);
nor U8395 (N_8395,N_50,N_4201);
nand U8396 (N_8396,N_4386,N_3426);
nor U8397 (N_8397,N_73,N_387);
nor U8398 (N_8398,N_1650,N_3940);
or U8399 (N_8399,N_2353,N_1470);
xor U8400 (N_8400,N_1633,N_1771);
and U8401 (N_8401,N_4439,N_2398);
and U8402 (N_8402,N_1770,N_3954);
and U8403 (N_8403,N_1839,N_2031);
nand U8404 (N_8404,N_631,N_4281);
or U8405 (N_8405,N_1765,N_2034);
xnor U8406 (N_8406,N_4764,N_927);
or U8407 (N_8407,N_4571,N_3929);
nor U8408 (N_8408,N_339,N_1676);
nor U8409 (N_8409,N_4379,N_3687);
or U8410 (N_8410,N_3328,N_1630);
or U8411 (N_8411,N_4227,N_2899);
and U8412 (N_8412,N_695,N_2791);
xnor U8413 (N_8413,N_2605,N_2519);
or U8414 (N_8414,N_1189,N_1970);
and U8415 (N_8415,N_3312,N_1190);
and U8416 (N_8416,N_1452,N_3001);
nor U8417 (N_8417,N_2474,N_412);
and U8418 (N_8418,N_2739,N_2202);
and U8419 (N_8419,N_1965,N_2973);
nor U8420 (N_8420,N_80,N_4191);
or U8421 (N_8421,N_1972,N_2760);
nand U8422 (N_8422,N_651,N_2331);
and U8423 (N_8423,N_2047,N_1397);
or U8424 (N_8424,N_1696,N_3588);
or U8425 (N_8425,N_3052,N_2334);
or U8426 (N_8426,N_2275,N_1268);
nor U8427 (N_8427,N_3840,N_3279);
or U8428 (N_8428,N_524,N_1069);
or U8429 (N_8429,N_2090,N_4950);
nand U8430 (N_8430,N_2532,N_4016);
xnor U8431 (N_8431,N_4389,N_2644);
or U8432 (N_8432,N_4945,N_3016);
xnor U8433 (N_8433,N_348,N_2631);
nor U8434 (N_8434,N_1781,N_4775);
and U8435 (N_8435,N_3428,N_1909);
nor U8436 (N_8436,N_3085,N_3959);
and U8437 (N_8437,N_2406,N_1306);
or U8438 (N_8438,N_3332,N_462);
or U8439 (N_8439,N_1668,N_2038);
or U8440 (N_8440,N_1678,N_1882);
and U8441 (N_8441,N_436,N_883);
and U8442 (N_8442,N_1086,N_2721);
nand U8443 (N_8443,N_3094,N_893);
nor U8444 (N_8444,N_25,N_3826);
and U8445 (N_8445,N_1654,N_2311);
or U8446 (N_8446,N_3207,N_4221);
and U8447 (N_8447,N_3233,N_294);
and U8448 (N_8448,N_1813,N_4884);
and U8449 (N_8449,N_4143,N_937);
and U8450 (N_8450,N_3451,N_3708);
nor U8451 (N_8451,N_303,N_2052);
nor U8452 (N_8452,N_986,N_4542);
or U8453 (N_8453,N_115,N_2337);
nand U8454 (N_8454,N_3097,N_565);
or U8455 (N_8455,N_1841,N_1290);
nand U8456 (N_8456,N_3833,N_532);
or U8457 (N_8457,N_675,N_248);
nor U8458 (N_8458,N_2666,N_3530);
xnor U8459 (N_8459,N_3352,N_4875);
xnor U8460 (N_8460,N_3287,N_2951);
nand U8461 (N_8461,N_4122,N_639);
nor U8462 (N_8462,N_4163,N_4935);
nand U8463 (N_8463,N_4668,N_2090);
nor U8464 (N_8464,N_4981,N_4850);
nand U8465 (N_8465,N_1345,N_2734);
and U8466 (N_8466,N_1397,N_1517);
or U8467 (N_8467,N_3271,N_4583);
nor U8468 (N_8468,N_1838,N_1600);
or U8469 (N_8469,N_4693,N_4508);
xor U8470 (N_8470,N_4951,N_2315);
nor U8471 (N_8471,N_593,N_2671);
and U8472 (N_8472,N_790,N_750);
nor U8473 (N_8473,N_2235,N_4794);
nand U8474 (N_8474,N_2231,N_1515);
and U8475 (N_8475,N_4762,N_931);
nand U8476 (N_8476,N_4159,N_2377);
or U8477 (N_8477,N_1785,N_4710);
and U8478 (N_8478,N_480,N_2163);
and U8479 (N_8479,N_3434,N_4641);
nand U8480 (N_8480,N_4118,N_2469);
and U8481 (N_8481,N_2547,N_1902);
and U8482 (N_8482,N_4335,N_4860);
nand U8483 (N_8483,N_3877,N_2976);
or U8484 (N_8484,N_1240,N_1026);
and U8485 (N_8485,N_4719,N_81);
nor U8486 (N_8486,N_1635,N_134);
and U8487 (N_8487,N_1405,N_2665);
or U8488 (N_8488,N_725,N_4433);
nor U8489 (N_8489,N_858,N_110);
nand U8490 (N_8490,N_2130,N_2122);
or U8491 (N_8491,N_2013,N_146);
xor U8492 (N_8492,N_966,N_2451);
and U8493 (N_8493,N_4532,N_1827);
nand U8494 (N_8494,N_1567,N_2188);
nand U8495 (N_8495,N_1593,N_3150);
and U8496 (N_8496,N_1606,N_2413);
and U8497 (N_8497,N_2618,N_4334);
and U8498 (N_8498,N_4336,N_1240);
or U8499 (N_8499,N_2823,N_4790);
or U8500 (N_8500,N_3714,N_2998);
xor U8501 (N_8501,N_178,N_3129);
and U8502 (N_8502,N_2767,N_186);
nor U8503 (N_8503,N_2131,N_4181);
or U8504 (N_8504,N_147,N_4798);
nand U8505 (N_8505,N_817,N_3149);
nor U8506 (N_8506,N_3850,N_4055);
and U8507 (N_8507,N_181,N_2000);
nand U8508 (N_8508,N_710,N_2248);
or U8509 (N_8509,N_398,N_2661);
nand U8510 (N_8510,N_1533,N_3671);
or U8511 (N_8511,N_322,N_1085);
xor U8512 (N_8512,N_3735,N_2799);
xor U8513 (N_8513,N_3372,N_259);
or U8514 (N_8514,N_1187,N_1914);
or U8515 (N_8515,N_3780,N_2132);
and U8516 (N_8516,N_613,N_3954);
nor U8517 (N_8517,N_1915,N_2762);
and U8518 (N_8518,N_1213,N_4140);
or U8519 (N_8519,N_2010,N_3979);
nor U8520 (N_8520,N_3470,N_2873);
or U8521 (N_8521,N_1636,N_933);
nand U8522 (N_8522,N_1155,N_2479);
nand U8523 (N_8523,N_1646,N_3242);
nor U8524 (N_8524,N_432,N_461);
nor U8525 (N_8525,N_4100,N_2252);
nand U8526 (N_8526,N_2754,N_424);
nor U8527 (N_8527,N_4496,N_3992);
nor U8528 (N_8528,N_4917,N_289);
and U8529 (N_8529,N_246,N_988);
nand U8530 (N_8530,N_160,N_1139);
nor U8531 (N_8531,N_3368,N_553);
or U8532 (N_8532,N_3218,N_3671);
or U8533 (N_8533,N_1851,N_1845);
and U8534 (N_8534,N_1878,N_1344);
nand U8535 (N_8535,N_796,N_1942);
or U8536 (N_8536,N_2172,N_1303);
or U8537 (N_8537,N_1133,N_3225);
or U8538 (N_8538,N_1251,N_3016);
nand U8539 (N_8539,N_2155,N_3894);
and U8540 (N_8540,N_3447,N_1862);
and U8541 (N_8541,N_2204,N_2983);
xor U8542 (N_8542,N_3625,N_2312);
and U8543 (N_8543,N_4664,N_2208);
or U8544 (N_8544,N_2200,N_2167);
nand U8545 (N_8545,N_3161,N_4696);
nor U8546 (N_8546,N_1124,N_4343);
and U8547 (N_8547,N_2556,N_4053);
or U8548 (N_8548,N_2171,N_1135);
or U8549 (N_8549,N_804,N_2283);
nor U8550 (N_8550,N_1659,N_1045);
nor U8551 (N_8551,N_126,N_2819);
and U8552 (N_8552,N_2874,N_3689);
nor U8553 (N_8553,N_1051,N_780);
nor U8554 (N_8554,N_210,N_2437);
nor U8555 (N_8555,N_1017,N_4436);
nor U8556 (N_8556,N_4511,N_2538);
and U8557 (N_8557,N_3024,N_4618);
and U8558 (N_8558,N_3026,N_4369);
nor U8559 (N_8559,N_3052,N_4508);
nor U8560 (N_8560,N_2594,N_2167);
nand U8561 (N_8561,N_2162,N_1737);
nor U8562 (N_8562,N_3642,N_1858);
and U8563 (N_8563,N_1925,N_2678);
nand U8564 (N_8564,N_582,N_4449);
or U8565 (N_8565,N_2464,N_3693);
nor U8566 (N_8566,N_2838,N_624);
nor U8567 (N_8567,N_3178,N_1646);
and U8568 (N_8568,N_759,N_176);
nor U8569 (N_8569,N_4321,N_589);
or U8570 (N_8570,N_4064,N_4943);
or U8571 (N_8571,N_2296,N_3139);
and U8572 (N_8572,N_2627,N_326);
nor U8573 (N_8573,N_3859,N_4738);
nor U8574 (N_8574,N_3044,N_723);
xor U8575 (N_8575,N_332,N_4338);
or U8576 (N_8576,N_3767,N_1362);
nand U8577 (N_8577,N_4288,N_4621);
nor U8578 (N_8578,N_4457,N_2549);
nor U8579 (N_8579,N_3660,N_1484);
nor U8580 (N_8580,N_2900,N_419);
and U8581 (N_8581,N_4472,N_3505);
xnor U8582 (N_8582,N_1912,N_4960);
xor U8583 (N_8583,N_782,N_3024);
and U8584 (N_8584,N_4151,N_2789);
and U8585 (N_8585,N_358,N_244);
nor U8586 (N_8586,N_2086,N_3998);
or U8587 (N_8587,N_3563,N_1168);
and U8588 (N_8588,N_727,N_2717);
or U8589 (N_8589,N_1762,N_2608);
and U8590 (N_8590,N_3418,N_4629);
and U8591 (N_8591,N_26,N_3623);
xnor U8592 (N_8592,N_2570,N_3479);
and U8593 (N_8593,N_1787,N_2132);
nand U8594 (N_8594,N_1736,N_1145);
and U8595 (N_8595,N_13,N_297);
and U8596 (N_8596,N_3563,N_3781);
and U8597 (N_8597,N_4406,N_2293);
xor U8598 (N_8598,N_2787,N_2866);
or U8599 (N_8599,N_2416,N_2160);
nor U8600 (N_8600,N_4797,N_3154);
nor U8601 (N_8601,N_1910,N_3032);
or U8602 (N_8602,N_3862,N_3809);
or U8603 (N_8603,N_1834,N_2331);
nand U8604 (N_8604,N_2671,N_4235);
and U8605 (N_8605,N_4830,N_2445);
and U8606 (N_8606,N_478,N_1971);
nand U8607 (N_8607,N_2201,N_3528);
and U8608 (N_8608,N_2841,N_1862);
nand U8609 (N_8609,N_4952,N_220);
nor U8610 (N_8610,N_534,N_1436);
and U8611 (N_8611,N_4408,N_902);
nor U8612 (N_8612,N_3425,N_869);
and U8613 (N_8613,N_4696,N_2014);
and U8614 (N_8614,N_1978,N_487);
nor U8615 (N_8615,N_4269,N_982);
and U8616 (N_8616,N_2290,N_2715);
xnor U8617 (N_8617,N_373,N_4927);
or U8618 (N_8618,N_3096,N_4694);
and U8619 (N_8619,N_4863,N_4596);
nor U8620 (N_8620,N_3982,N_1163);
nand U8621 (N_8621,N_4992,N_4002);
nand U8622 (N_8622,N_1217,N_2704);
and U8623 (N_8623,N_3961,N_1400);
xnor U8624 (N_8624,N_1090,N_2108);
nor U8625 (N_8625,N_1442,N_4139);
nand U8626 (N_8626,N_802,N_1098);
xor U8627 (N_8627,N_1409,N_2812);
nand U8628 (N_8628,N_2457,N_3037);
nor U8629 (N_8629,N_3262,N_78);
nand U8630 (N_8630,N_1680,N_1075);
and U8631 (N_8631,N_1819,N_3586);
or U8632 (N_8632,N_1632,N_4992);
nor U8633 (N_8633,N_4630,N_1963);
xor U8634 (N_8634,N_472,N_3073);
and U8635 (N_8635,N_281,N_2611);
nand U8636 (N_8636,N_2549,N_4678);
nor U8637 (N_8637,N_4614,N_4679);
nand U8638 (N_8638,N_1599,N_1683);
and U8639 (N_8639,N_3825,N_1825);
and U8640 (N_8640,N_865,N_1221);
and U8641 (N_8641,N_1652,N_2020);
and U8642 (N_8642,N_3706,N_4155);
nor U8643 (N_8643,N_2956,N_3816);
nand U8644 (N_8644,N_1669,N_3848);
or U8645 (N_8645,N_2262,N_439);
or U8646 (N_8646,N_1469,N_4489);
nand U8647 (N_8647,N_3969,N_2106);
and U8648 (N_8648,N_1953,N_4335);
or U8649 (N_8649,N_2559,N_201);
xnor U8650 (N_8650,N_0,N_4624);
xor U8651 (N_8651,N_7,N_1822);
or U8652 (N_8652,N_2444,N_1542);
or U8653 (N_8653,N_2625,N_2618);
nor U8654 (N_8654,N_1850,N_4405);
and U8655 (N_8655,N_1302,N_836);
or U8656 (N_8656,N_2696,N_4802);
nand U8657 (N_8657,N_1316,N_618);
nand U8658 (N_8658,N_4752,N_311);
nor U8659 (N_8659,N_880,N_559);
or U8660 (N_8660,N_4604,N_4441);
or U8661 (N_8661,N_4466,N_2011);
or U8662 (N_8662,N_4861,N_0);
nand U8663 (N_8663,N_2017,N_2292);
or U8664 (N_8664,N_2482,N_495);
xor U8665 (N_8665,N_3898,N_123);
nor U8666 (N_8666,N_2821,N_4133);
and U8667 (N_8667,N_3945,N_4908);
xor U8668 (N_8668,N_902,N_3695);
nand U8669 (N_8669,N_3225,N_3938);
and U8670 (N_8670,N_1951,N_4301);
and U8671 (N_8671,N_3279,N_1790);
nor U8672 (N_8672,N_224,N_2120);
or U8673 (N_8673,N_3388,N_4068);
and U8674 (N_8674,N_4448,N_4584);
or U8675 (N_8675,N_2387,N_2793);
or U8676 (N_8676,N_4607,N_4076);
nor U8677 (N_8677,N_2282,N_523);
xor U8678 (N_8678,N_2252,N_855);
nor U8679 (N_8679,N_4420,N_672);
nor U8680 (N_8680,N_2956,N_1516);
nand U8681 (N_8681,N_4252,N_2434);
nor U8682 (N_8682,N_3378,N_3323);
or U8683 (N_8683,N_2727,N_693);
and U8684 (N_8684,N_2432,N_1557);
or U8685 (N_8685,N_3318,N_3332);
and U8686 (N_8686,N_4234,N_1065);
xor U8687 (N_8687,N_767,N_2864);
nor U8688 (N_8688,N_2193,N_4022);
and U8689 (N_8689,N_790,N_2920);
xnor U8690 (N_8690,N_4584,N_3578);
nand U8691 (N_8691,N_3079,N_590);
nor U8692 (N_8692,N_4976,N_2339);
nor U8693 (N_8693,N_4712,N_3063);
or U8694 (N_8694,N_3829,N_1259);
or U8695 (N_8695,N_878,N_2518);
nor U8696 (N_8696,N_64,N_3319);
and U8697 (N_8697,N_4608,N_465);
and U8698 (N_8698,N_4900,N_3228);
nand U8699 (N_8699,N_3336,N_3248);
and U8700 (N_8700,N_3051,N_3131);
and U8701 (N_8701,N_1410,N_4162);
nor U8702 (N_8702,N_2660,N_237);
and U8703 (N_8703,N_3311,N_317);
and U8704 (N_8704,N_3593,N_1113);
nor U8705 (N_8705,N_4392,N_3461);
or U8706 (N_8706,N_2021,N_3357);
or U8707 (N_8707,N_800,N_4099);
and U8708 (N_8708,N_612,N_4438);
and U8709 (N_8709,N_3516,N_225);
nor U8710 (N_8710,N_3985,N_2458);
nor U8711 (N_8711,N_4347,N_4294);
xnor U8712 (N_8712,N_3440,N_1618);
and U8713 (N_8713,N_1486,N_1011);
nand U8714 (N_8714,N_4738,N_2038);
or U8715 (N_8715,N_2606,N_336);
and U8716 (N_8716,N_3142,N_4238);
nand U8717 (N_8717,N_3815,N_3317);
or U8718 (N_8718,N_2333,N_4379);
or U8719 (N_8719,N_3562,N_3800);
nand U8720 (N_8720,N_1795,N_922);
nor U8721 (N_8721,N_2023,N_4042);
nand U8722 (N_8722,N_3260,N_1057);
or U8723 (N_8723,N_1472,N_2735);
nand U8724 (N_8724,N_4159,N_4203);
or U8725 (N_8725,N_3262,N_1806);
nand U8726 (N_8726,N_4575,N_3820);
nand U8727 (N_8727,N_1756,N_3870);
nand U8728 (N_8728,N_2280,N_3377);
or U8729 (N_8729,N_2347,N_2101);
or U8730 (N_8730,N_3422,N_3347);
nor U8731 (N_8731,N_2526,N_2737);
nor U8732 (N_8732,N_2067,N_497);
or U8733 (N_8733,N_4790,N_1314);
or U8734 (N_8734,N_4683,N_4999);
nand U8735 (N_8735,N_1978,N_4414);
nand U8736 (N_8736,N_1088,N_4788);
nand U8737 (N_8737,N_4312,N_4015);
and U8738 (N_8738,N_4785,N_2039);
nand U8739 (N_8739,N_129,N_4882);
xnor U8740 (N_8740,N_717,N_1567);
xnor U8741 (N_8741,N_833,N_51);
and U8742 (N_8742,N_3458,N_1722);
nand U8743 (N_8743,N_3032,N_4254);
or U8744 (N_8744,N_1180,N_1928);
nor U8745 (N_8745,N_1330,N_3714);
or U8746 (N_8746,N_176,N_2005);
nor U8747 (N_8747,N_2722,N_4971);
nand U8748 (N_8748,N_4298,N_4562);
or U8749 (N_8749,N_1261,N_3686);
xor U8750 (N_8750,N_1291,N_1691);
or U8751 (N_8751,N_1812,N_4957);
or U8752 (N_8752,N_377,N_4287);
and U8753 (N_8753,N_4196,N_3892);
nand U8754 (N_8754,N_4095,N_4878);
nand U8755 (N_8755,N_834,N_3101);
xnor U8756 (N_8756,N_407,N_3608);
nor U8757 (N_8757,N_452,N_4225);
and U8758 (N_8758,N_1084,N_4545);
nor U8759 (N_8759,N_2121,N_1033);
and U8760 (N_8760,N_841,N_3154);
xnor U8761 (N_8761,N_4711,N_1081);
and U8762 (N_8762,N_4241,N_2499);
nor U8763 (N_8763,N_495,N_3451);
nor U8764 (N_8764,N_593,N_4208);
or U8765 (N_8765,N_2071,N_2056);
nand U8766 (N_8766,N_1190,N_3445);
nand U8767 (N_8767,N_2324,N_2820);
xnor U8768 (N_8768,N_2852,N_4983);
and U8769 (N_8769,N_449,N_400);
nand U8770 (N_8770,N_2787,N_2471);
or U8771 (N_8771,N_1360,N_3569);
nor U8772 (N_8772,N_4686,N_1951);
nand U8773 (N_8773,N_2992,N_477);
and U8774 (N_8774,N_4363,N_3046);
and U8775 (N_8775,N_3022,N_2032);
nand U8776 (N_8776,N_2688,N_3856);
xor U8777 (N_8777,N_4255,N_3056);
nor U8778 (N_8778,N_4388,N_4804);
nand U8779 (N_8779,N_4420,N_1312);
nor U8780 (N_8780,N_4385,N_3135);
or U8781 (N_8781,N_3516,N_4461);
nor U8782 (N_8782,N_4172,N_1161);
or U8783 (N_8783,N_4666,N_3861);
nor U8784 (N_8784,N_3262,N_3066);
nor U8785 (N_8785,N_3209,N_3837);
nor U8786 (N_8786,N_1669,N_91);
nor U8787 (N_8787,N_4211,N_909);
nand U8788 (N_8788,N_1858,N_2874);
nor U8789 (N_8789,N_10,N_1891);
or U8790 (N_8790,N_3395,N_3581);
or U8791 (N_8791,N_2950,N_2609);
nand U8792 (N_8792,N_42,N_4176);
nand U8793 (N_8793,N_4967,N_4544);
nand U8794 (N_8794,N_4613,N_405);
and U8795 (N_8795,N_921,N_2200);
and U8796 (N_8796,N_2455,N_4108);
xnor U8797 (N_8797,N_2062,N_3258);
or U8798 (N_8798,N_3053,N_864);
nor U8799 (N_8799,N_3454,N_2293);
and U8800 (N_8800,N_2610,N_4871);
and U8801 (N_8801,N_490,N_4786);
or U8802 (N_8802,N_3409,N_4912);
and U8803 (N_8803,N_661,N_970);
and U8804 (N_8804,N_2012,N_2820);
nor U8805 (N_8805,N_4029,N_3220);
nand U8806 (N_8806,N_4566,N_1153);
xnor U8807 (N_8807,N_2419,N_396);
xnor U8808 (N_8808,N_132,N_3869);
xor U8809 (N_8809,N_4800,N_552);
xnor U8810 (N_8810,N_4723,N_2145);
and U8811 (N_8811,N_4966,N_3213);
and U8812 (N_8812,N_804,N_4915);
and U8813 (N_8813,N_1613,N_4876);
nand U8814 (N_8814,N_1177,N_3306);
and U8815 (N_8815,N_3550,N_3312);
nand U8816 (N_8816,N_3685,N_3181);
nor U8817 (N_8817,N_4019,N_476);
nor U8818 (N_8818,N_2371,N_3083);
nand U8819 (N_8819,N_3786,N_762);
nand U8820 (N_8820,N_202,N_2224);
nand U8821 (N_8821,N_630,N_1168);
or U8822 (N_8822,N_2932,N_2866);
or U8823 (N_8823,N_1241,N_2226);
nand U8824 (N_8824,N_442,N_4063);
nand U8825 (N_8825,N_1456,N_1674);
or U8826 (N_8826,N_1882,N_3167);
nand U8827 (N_8827,N_3685,N_222);
nor U8828 (N_8828,N_4943,N_4820);
xnor U8829 (N_8829,N_3955,N_2526);
nand U8830 (N_8830,N_4398,N_3836);
or U8831 (N_8831,N_3111,N_3464);
nand U8832 (N_8832,N_2940,N_4139);
xor U8833 (N_8833,N_2822,N_2479);
nor U8834 (N_8834,N_2257,N_2940);
xor U8835 (N_8835,N_1054,N_4006);
or U8836 (N_8836,N_1227,N_135);
or U8837 (N_8837,N_484,N_1366);
nor U8838 (N_8838,N_2373,N_562);
nand U8839 (N_8839,N_3579,N_4262);
or U8840 (N_8840,N_1570,N_3889);
xor U8841 (N_8841,N_4605,N_2815);
xnor U8842 (N_8842,N_3152,N_4990);
nor U8843 (N_8843,N_105,N_1831);
or U8844 (N_8844,N_2884,N_2589);
or U8845 (N_8845,N_1453,N_1841);
nand U8846 (N_8846,N_3085,N_230);
and U8847 (N_8847,N_317,N_398);
or U8848 (N_8848,N_2474,N_1029);
nor U8849 (N_8849,N_4604,N_3251);
nor U8850 (N_8850,N_4780,N_3590);
nand U8851 (N_8851,N_2547,N_3736);
nor U8852 (N_8852,N_3168,N_60);
and U8853 (N_8853,N_4245,N_2324);
or U8854 (N_8854,N_1550,N_2878);
or U8855 (N_8855,N_2941,N_4632);
and U8856 (N_8856,N_757,N_1403);
or U8857 (N_8857,N_975,N_1532);
nand U8858 (N_8858,N_1591,N_1992);
nand U8859 (N_8859,N_3381,N_46);
or U8860 (N_8860,N_3117,N_4087);
and U8861 (N_8861,N_1510,N_2425);
and U8862 (N_8862,N_4019,N_1550);
nand U8863 (N_8863,N_875,N_136);
or U8864 (N_8864,N_13,N_2098);
xnor U8865 (N_8865,N_1911,N_1006);
or U8866 (N_8866,N_771,N_4063);
xor U8867 (N_8867,N_3628,N_676);
or U8868 (N_8868,N_4754,N_1616);
and U8869 (N_8869,N_2962,N_2220);
nand U8870 (N_8870,N_1886,N_4558);
and U8871 (N_8871,N_3197,N_2420);
or U8872 (N_8872,N_3909,N_987);
xor U8873 (N_8873,N_2888,N_477);
or U8874 (N_8874,N_2096,N_2291);
nand U8875 (N_8875,N_2001,N_2156);
xnor U8876 (N_8876,N_3687,N_1110);
xnor U8877 (N_8877,N_81,N_2118);
and U8878 (N_8878,N_4814,N_51);
nor U8879 (N_8879,N_2131,N_3864);
and U8880 (N_8880,N_1309,N_648);
nand U8881 (N_8881,N_3496,N_3135);
or U8882 (N_8882,N_3899,N_4095);
nand U8883 (N_8883,N_2223,N_3319);
or U8884 (N_8884,N_493,N_4233);
or U8885 (N_8885,N_1564,N_371);
and U8886 (N_8886,N_136,N_462);
or U8887 (N_8887,N_3595,N_1906);
nand U8888 (N_8888,N_3505,N_1215);
nor U8889 (N_8889,N_516,N_3181);
nor U8890 (N_8890,N_3299,N_1555);
or U8891 (N_8891,N_1803,N_3864);
xor U8892 (N_8892,N_3676,N_297);
nor U8893 (N_8893,N_3855,N_4590);
and U8894 (N_8894,N_3708,N_2139);
nor U8895 (N_8895,N_789,N_1710);
xnor U8896 (N_8896,N_3759,N_16);
nor U8897 (N_8897,N_4449,N_1258);
nor U8898 (N_8898,N_4181,N_724);
or U8899 (N_8899,N_2821,N_4517);
or U8900 (N_8900,N_4637,N_1511);
nor U8901 (N_8901,N_1062,N_3597);
nor U8902 (N_8902,N_2259,N_2721);
or U8903 (N_8903,N_1917,N_2436);
nor U8904 (N_8904,N_3761,N_4766);
or U8905 (N_8905,N_4824,N_2717);
or U8906 (N_8906,N_2315,N_3213);
and U8907 (N_8907,N_3733,N_2335);
xor U8908 (N_8908,N_1835,N_216);
nor U8909 (N_8909,N_3188,N_1248);
nand U8910 (N_8910,N_3494,N_4944);
nor U8911 (N_8911,N_1176,N_2705);
nand U8912 (N_8912,N_4460,N_2234);
nor U8913 (N_8913,N_4996,N_1559);
nor U8914 (N_8914,N_733,N_2074);
nand U8915 (N_8915,N_4939,N_3537);
and U8916 (N_8916,N_4343,N_94);
and U8917 (N_8917,N_3057,N_2866);
or U8918 (N_8918,N_1686,N_4762);
nor U8919 (N_8919,N_3923,N_1646);
and U8920 (N_8920,N_2024,N_834);
nor U8921 (N_8921,N_4199,N_1709);
and U8922 (N_8922,N_4443,N_441);
nand U8923 (N_8923,N_3200,N_2065);
and U8924 (N_8924,N_1079,N_3509);
nor U8925 (N_8925,N_3202,N_574);
and U8926 (N_8926,N_3311,N_3959);
or U8927 (N_8927,N_712,N_1008);
or U8928 (N_8928,N_1726,N_3453);
nor U8929 (N_8929,N_1942,N_931);
nand U8930 (N_8930,N_4358,N_3609);
or U8931 (N_8931,N_3910,N_2191);
nor U8932 (N_8932,N_2393,N_2582);
nor U8933 (N_8933,N_1188,N_633);
nand U8934 (N_8934,N_114,N_864);
nand U8935 (N_8935,N_3545,N_4164);
nor U8936 (N_8936,N_2545,N_4230);
xor U8937 (N_8937,N_3631,N_3719);
nor U8938 (N_8938,N_4097,N_546);
and U8939 (N_8939,N_4182,N_1922);
or U8940 (N_8940,N_505,N_2077);
or U8941 (N_8941,N_2088,N_3103);
or U8942 (N_8942,N_1463,N_2264);
and U8943 (N_8943,N_3880,N_2429);
or U8944 (N_8944,N_3389,N_1049);
or U8945 (N_8945,N_579,N_376);
xnor U8946 (N_8946,N_4270,N_4080);
and U8947 (N_8947,N_3178,N_968);
and U8948 (N_8948,N_2691,N_3919);
or U8949 (N_8949,N_3302,N_2067);
and U8950 (N_8950,N_2968,N_3476);
nor U8951 (N_8951,N_4019,N_3048);
or U8952 (N_8952,N_2345,N_1522);
or U8953 (N_8953,N_2090,N_2346);
and U8954 (N_8954,N_2381,N_663);
nand U8955 (N_8955,N_881,N_4999);
nor U8956 (N_8956,N_2220,N_3141);
xnor U8957 (N_8957,N_4078,N_1914);
nor U8958 (N_8958,N_4011,N_2892);
nor U8959 (N_8959,N_1425,N_1450);
and U8960 (N_8960,N_62,N_3488);
nor U8961 (N_8961,N_2617,N_2586);
nand U8962 (N_8962,N_2225,N_3100);
or U8963 (N_8963,N_404,N_3638);
nand U8964 (N_8964,N_1298,N_163);
nor U8965 (N_8965,N_1133,N_1487);
nand U8966 (N_8966,N_1668,N_1430);
nand U8967 (N_8967,N_1615,N_3261);
nand U8968 (N_8968,N_3485,N_4184);
nand U8969 (N_8969,N_1963,N_852);
or U8970 (N_8970,N_1608,N_1692);
or U8971 (N_8971,N_154,N_2309);
nor U8972 (N_8972,N_593,N_3097);
and U8973 (N_8973,N_1252,N_3239);
and U8974 (N_8974,N_919,N_4249);
nand U8975 (N_8975,N_2575,N_740);
nor U8976 (N_8976,N_2681,N_3478);
or U8977 (N_8977,N_1984,N_1173);
or U8978 (N_8978,N_3942,N_2914);
or U8979 (N_8979,N_1501,N_2904);
nand U8980 (N_8980,N_4447,N_1353);
nand U8981 (N_8981,N_1112,N_2193);
nand U8982 (N_8982,N_3282,N_811);
nand U8983 (N_8983,N_4379,N_3675);
nand U8984 (N_8984,N_4156,N_485);
nand U8985 (N_8985,N_1595,N_401);
nand U8986 (N_8986,N_1483,N_266);
and U8987 (N_8987,N_1252,N_668);
or U8988 (N_8988,N_1871,N_2416);
nand U8989 (N_8989,N_1335,N_4010);
nor U8990 (N_8990,N_1637,N_3876);
and U8991 (N_8991,N_523,N_3186);
nor U8992 (N_8992,N_3397,N_1259);
or U8993 (N_8993,N_532,N_3345);
nor U8994 (N_8994,N_154,N_4660);
xor U8995 (N_8995,N_2164,N_4986);
nand U8996 (N_8996,N_1566,N_405);
or U8997 (N_8997,N_3490,N_310);
nand U8998 (N_8998,N_193,N_1609);
or U8999 (N_8999,N_2265,N_578);
nand U9000 (N_9000,N_1847,N_2498);
nor U9001 (N_9001,N_2282,N_698);
nor U9002 (N_9002,N_3905,N_3691);
nand U9003 (N_9003,N_4957,N_4842);
nand U9004 (N_9004,N_4616,N_4897);
or U9005 (N_9005,N_1579,N_2482);
or U9006 (N_9006,N_2864,N_4870);
nand U9007 (N_9007,N_3591,N_1868);
nor U9008 (N_9008,N_3636,N_1958);
or U9009 (N_9009,N_111,N_1629);
nand U9010 (N_9010,N_4754,N_2162);
and U9011 (N_9011,N_4441,N_4666);
and U9012 (N_9012,N_827,N_4169);
nand U9013 (N_9013,N_4960,N_4851);
and U9014 (N_9014,N_309,N_3975);
and U9015 (N_9015,N_1333,N_3605);
nand U9016 (N_9016,N_1019,N_1106);
or U9017 (N_9017,N_901,N_4521);
xnor U9018 (N_9018,N_2646,N_3301);
nor U9019 (N_9019,N_962,N_1428);
xor U9020 (N_9020,N_2667,N_4327);
nand U9021 (N_9021,N_4304,N_3877);
or U9022 (N_9022,N_1996,N_3876);
nor U9023 (N_9023,N_2987,N_2255);
nand U9024 (N_9024,N_4445,N_4427);
or U9025 (N_9025,N_723,N_1428);
xnor U9026 (N_9026,N_2796,N_440);
nor U9027 (N_9027,N_4989,N_1720);
nand U9028 (N_9028,N_3088,N_3354);
nand U9029 (N_9029,N_2179,N_3082);
nand U9030 (N_9030,N_3855,N_3713);
nor U9031 (N_9031,N_1279,N_4533);
or U9032 (N_9032,N_2939,N_299);
and U9033 (N_9033,N_3729,N_3396);
nand U9034 (N_9034,N_4321,N_1028);
nor U9035 (N_9035,N_2886,N_627);
xnor U9036 (N_9036,N_235,N_1788);
nor U9037 (N_9037,N_1806,N_4986);
and U9038 (N_9038,N_3255,N_3456);
or U9039 (N_9039,N_4033,N_455);
nand U9040 (N_9040,N_4457,N_3060);
nand U9041 (N_9041,N_3062,N_1375);
or U9042 (N_9042,N_798,N_1170);
nand U9043 (N_9043,N_4082,N_2490);
or U9044 (N_9044,N_3643,N_2468);
or U9045 (N_9045,N_1711,N_4011);
or U9046 (N_9046,N_578,N_2043);
and U9047 (N_9047,N_2536,N_3395);
and U9048 (N_9048,N_3418,N_562);
nor U9049 (N_9049,N_2335,N_2857);
and U9050 (N_9050,N_813,N_4224);
or U9051 (N_9051,N_4385,N_3754);
and U9052 (N_9052,N_2785,N_2932);
nor U9053 (N_9053,N_455,N_2819);
nor U9054 (N_9054,N_2055,N_2582);
or U9055 (N_9055,N_3829,N_2202);
nor U9056 (N_9056,N_4419,N_2797);
nor U9057 (N_9057,N_1599,N_3751);
nor U9058 (N_9058,N_4320,N_3580);
nor U9059 (N_9059,N_3716,N_1293);
nand U9060 (N_9060,N_4452,N_2523);
nor U9061 (N_9061,N_3727,N_3489);
and U9062 (N_9062,N_241,N_3942);
nand U9063 (N_9063,N_2573,N_2618);
and U9064 (N_9064,N_2355,N_3106);
or U9065 (N_9065,N_824,N_4829);
and U9066 (N_9066,N_4660,N_2507);
or U9067 (N_9067,N_2154,N_915);
and U9068 (N_9068,N_1759,N_1362);
and U9069 (N_9069,N_335,N_4301);
nor U9070 (N_9070,N_2115,N_1117);
nand U9071 (N_9071,N_2068,N_2117);
nand U9072 (N_9072,N_3122,N_1199);
xor U9073 (N_9073,N_4677,N_4390);
nor U9074 (N_9074,N_3137,N_1847);
or U9075 (N_9075,N_4084,N_4342);
and U9076 (N_9076,N_1853,N_1619);
nand U9077 (N_9077,N_3470,N_1734);
or U9078 (N_9078,N_2011,N_4257);
or U9079 (N_9079,N_4901,N_2608);
and U9080 (N_9080,N_4639,N_2165);
nor U9081 (N_9081,N_2999,N_3742);
or U9082 (N_9082,N_1837,N_4309);
and U9083 (N_9083,N_3838,N_150);
xor U9084 (N_9084,N_155,N_890);
or U9085 (N_9085,N_1373,N_4940);
nor U9086 (N_9086,N_1550,N_3115);
nand U9087 (N_9087,N_1148,N_1105);
nor U9088 (N_9088,N_1093,N_4300);
and U9089 (N_9089,N_2589,N_4049);
nor U9090 (N_9090,N_328,N_4085);
and U9091 (N_9091,N_3661,N_2363);
or U9092 (N_9092,N_3019,N_1660);
nor U9093 (N_9093,N_4022,N_3421);
nor U9094 (N_9094,N_2201,N_695);
and U9095 (N_9095,N_42,N_2771);
nor U9096 (N_9096,N_3636,N_2286);
and U9097 (N_9097,N_2485,N_3848);
and U9098 (N_9098,N_3972,N_1909);
and U9099 (N_9099,N_1056,N_664);
nand U9100 (N_9100,N_2616,N_2442);
xnor U9101 (N_9101,N_2411,N_946);
nor U9102 (N_9102,N_1157,N_385);
nor U9103 (N_9103,N_328,N_1406);
and U9104 (N_9104,N_904,N_3749);
or U9105 (N_9105,N_3459,N_72);
xnor U9106 (N_9106,N_4974,N_3946);
nand U9107 (N_9107,N_2462,N_2444);
nor U9108 (N_9108,N_1907,N_3705);
nor U9109 (N_9109,N_534,N_3788);
or U9110 (N_9110,N_4263,N_4552);
nor U9111 (N_9111,N_4749,N_4587);
nand U9112 (N_9112,N_2424,N_3162);
and U9113 (N_9113,N_1937,N_866);
or U9114 (N_9114,N_2651,N_3767);
or U9115 (N_9115,N_3225,N_2847);
nor U9116 (N_9116,N_2659,N_2261);
nand U9117 (N_9117,N_529,N_1808);
nor U9118 (N_9118,N_1087,N_1250);
nor U9119 (N_9119,N_693,N_4886);
or U9120 (N_9120,N_402,N_888);
nor U9121 (N_9121,N_2813,N_1715);
or U9122 (N_9122,N_930,N_1262);
and U9123 (N_9123,N_3739,N_3028);
nand U9124 (N_9124,N_4315,N_1062);
xor U9125 (N_9125,N_1352,N_2938);
nand U9126 (N_9126,N_4225,N_1458);
nand U9127 (N_9127,N_3538,N_796);
nand U9128 (N_9128,N_1408,N_4911);
and U9129 (N_9129,N_555,N_3882);
nor U9130 (N_9130,N_3667,N_1157);
or U9131 (N_9131,N_1145,N_4167);
and U9132 (N_9132,N_2561,N_862);
and U9133 (N_9133,N_4609,N_1171);
or U9134 (N_9134,N_4654,N_4731);
or U9135 (N_9135,N_2328,N_1712);
nand U9136 (N_9136,N_1452,N_4318);
nand U9137 (N_9137,N_4518,N_3459);
nor U9138 (N_9138,N_21,N_4413);
or U9139 (N_9139,N_4556,N_4172);
xor U9140 (N_9140,N_2621,N_2011);
xor U9141 (N_9141,N_4266,N_4798);
and U9142 (N_9142,N_2340,N_1159);
nor U9143 (N_9143,N_3531,N_1230);
xor U9144 (N_9144,N_1623,N_3988);
or U9145 (N_9145,N_654,N_4050);
nor U9146 (N_9146,N_2231,N_2686);
xnor U9147 (N_9147,N_4548,N_3567);
or U9148 (N_9148,N_921,N_4059);
or U9149 (N_9149,N_3254,N_4342);
and U9150 (N_9150,N_4176,N_1618);
and U9151 (N_9151,N_4984,N_1230);
nand U9152 (N_9152,N_2258,N_1397);
nand U9153 (N_9153,N_2389,N_4705);
xor U9154 (N_9154,N_1106,N_346);
or U9155 (N_9155,N_4346,N_886);
or U9156 (N_9156,N_1819,N_4035);
nand U9157 (N_9157,N_2945,N_3999);
nand U9158 (N_9158,N_4322,N_1715);
nand U9159 (N_9159,N_2433,N_606);
nor U9160 (N_9160,N_2339,N_961);
nor U9161 (N_9161,N_1128,N_2081);
xnor U9162 (N_9162,N_3296,N_4600);
and U9163 (N_9163,N_4373,N_2822);
nand U9164 (N_9164,N_1603,N_880);
nand U9165 (N_9165,N_2448,N_4674);
nand U9166 (N_9166,N_312,N_326);
or U9167 (N_9167,N_3208,N_2880);
and U9168 (N_9168,N_2754,N_681);
and U9169 (N_9169,N_287,N_1191);
nand U9170 (N_9170,N_4238,N_2567);
nor U9171 (N_9171,N_148,N_2864);
and U9172 (N_9172,N_771,N_2550);
or U9173 (N_9173,N_348,N_2931);
nor U9174 (N_9174,N_4407,N_3522);
nor U9175 (N_9175,N_2150,N_575);
and U9176 (N_9176,N_753,N_1362);
nand U9177 (N_9177,N_825,N_1696);
nor U9178 (N_9178,N_1467,N_3442);
xor U9179 (N_9179,N_876,N_4703);
nand U9180 (N_9180,N_2366,N_1698);
nor U9181 (N_9181,N_873,N_4673);
nor U9182 (N_9182,N_721,N_1877);
and U9183 (N_9183,N_1829,N_1481);
nand U9184 (N_9184,N_4625,N_2902);
nand U9185 (N_9185,N_3585,N_4525);
xor U9186 (N_9186,N_3758,N_2271);
and U9187 (N_9187,N_3230,N_3534);
nand U9188 (N_9188,N_547,N_293);
nand U9189 (N_9189,N_379,N_2067);
nand U9190 (N_9190,N_3186,N_3192);
or U9191 (N_9191,N_4569,N_2156);
or U9192 (N_9192,N_358,N_3106);
or U9193 (N_9193,N_3105,N_3902);
and U9194 (N_9194,N_3609,N_4204);
or U9195 (N_9195,N_1062,N_4928);
and U9196 (N_9196,N_595,N_1939);
nand U9197 (N_9197,N_3619,N_1138);
or U9198 (N_9198,N_306,N_111);
and U9199 (N_9199,N_2700,N_4779);
and U9200 (N_9200,N_912,N_4003);
or U9201 (N_9201,N_1780,N_2694);
nor U9202 (N_9202,N_789,N_4354);
or U9203 (N_9203,N_1244,N_1756);
or U9204 (N_9204,N_2886,N_1304);
and U9205 (N_9205,N_4461,N_4376);
or U9206 (N_9206,N_3832,N_1090);
xor U9207 (N_9207,N_2594,N_4410);
and U9208 (N_9208,N_2901,N_4067);
nor U9209 (N_9209,N_3975,N_717);
nand U9210 (N_9210,N_3399,N_1983);
nand U9211 (N_9211,N_4708,N_2146);
nor U9212 (N_9212,N_4517,N_3524);
xnor U9213 (N_9213,N_2501,N_4894);
nor U9214 (N_9214,N_1259,N_1475);
nor U9215 (N_9215,N_1557,N_1792);
and U9216 (N_9216,N_4321,N_2865);
nor U9217 (N_9217,N_993,N_1515);
nor U9218 (N_9218,N_471,N_896);
nand U9219 (N_9219,N_3159,N_811);
nand U9220 (N_9220,N_2720,N_4745);
and U9221 (N_9221,N_140,N_2436);
nand U9222 (N_9222,N_2170,N_2948);
or U9223 (N_9223,N_3224,N_120);
or U9224 (N_9224,N_3558,N_3449);
nand U9225 (N_9225,N_232,N_1028);
nand U9226 (N_9226,N_4631,N_1759);
and U9227 (N_9227,N_546,N_2081);
xor U9228 (N_9228,N_1522,N_380);
nand U9229 (N_9229,N_715,N_4053);
xnor U9230 (N_9230,N_4857,N_2137);
and U9231 (N_9231,N_2583,N_1577);
nand U9232 (N_9232,N_2031,N_4099);
nand U9233 (N_9233,N_4638,N_4924);
xnor U9234 (N_9234,N_4472,N_66);
nand U9235 (N_9235,N_3353,N_3346);
and U9236 (N_9236,N_3098,N_4477);
and U9237 (N_9237,N_4133,N_3);
or U9238 (N_9238,N_91,N_1125);
or U9239 (N_9239,N_1088,N_1009);
and U9240 (N_9240,N_4109,N_3371);
or U9241 (N_9241,N_3276,N_3988);
or U9242 (N_9242,N_4518,N_3952);
or U9243 (N_9243,N_3970,N_2864);
and U9244 (N_9244,N_4629,N_4620);
nor U9245 (N_9245,N_467,N_2157);
and U9246 (N_9246,N_982,N_1922);
and U9247 (N_9247,N_4661,N_977);
nor U9248 (N_9248,N_2907,N_4436);
nor U9249 (N_9249,N_1297,N_53);
or U9250 (N_9250,N_2058,N_1700);
nand U9251 (N_9251,N_4634,N_2168);
nor U9252 (N_9252,N_3765,N_356);
nor U9253 (N_9253,N_1030,N_981);
or U9254 (N_9254,N_150,N_2647);
and U9255 (N_9255,N_3847,N_4005);
nand U9256 (N_9256,N_1933,N_4172);
nor U9257 (N_9257,N_4869,N_4794);
nand U9258 (N_9258,N_1420,N_2496);
xor U9259 (N_9259,N_3915,N_1569);
and U9260 (N_9260,N_2632,N_814);
and U9261 (N_9261,N_3212,N_4688);
xor U9262 (N_9262,N_2630,N_3877);
nor U9263 (N_9263,N_3431,N_4893);
nor U9264 (N_9264,N_508,N_3929);
nor U9265 (N_9265,N_2922,N_3477);
or U9266 (N_9266,N_2175,N_446);
nand U9267 (N_9267,N_1278,N_3026);
nor U9268 (N_9268,N_2802,N_2800);
nand U9269 (N_9269,N_4819,N_4072);
nor U9270 (N_9270,N_3060,N_2900);
nand U9271 (N_9271,N_1468,N_6);
nand U9272 (N_9272,N_4859,N_3465);
and U9273 (N_9273,N_4859,N_4927);
nor U9274 (N_9274,N_1044,N_3665);
nand U9275 (N_9275,N_3896,N_1667);
xnor U9276 (N_9276,N_3137,N_4749);
or U9277 (N_9277,N_311,N_4278);
nor U9278 (N_9278,N_2172,N_4165);
and U9279 (N_9279,N_4985,N_2071);
nor U9280 (N_9280,N_4634,N_1169);
nor U9281 (N_9281,N_1840,N_213);
xnor U9282 (N_9282,N_427,N_1638);
nand U9283 (N_9283,N_1863,N_1843);
or U9284 (N_9284,N_4706,N_872);
nor U9285 (N_9285,N_1934,N_434);
nand U9286 (N_9286,N_4222,N_1285);
or U9287 (N_9287,N_4308,N_2477);
nor U9288 (N_9288,N_3769,N_1605);
nand U9289 (N_9289,N_3723,N_2422);
or U9290 (N_9290,N_628,N_969);
nor U9291 (N_9291,N_2945,N_411);
and U9292 (N_9292,N_259,N_644);
and U9293 (N_9293,N_3685,N_3867);
nand U9294 (N_9294,N_44,N_3069);
xor U9295 (N_9295,N_4884,N_112);
xor U9296 (N_9296,N_1458,N_4617);
nand U9297 (N_9297,N_1505,N_768);
nand U9298 (N_9298,N_3158,N_460);
and U9299 (N_9299,N_4451,N_573);
xnor U9300 (N_9300,N_845,N_2183);
and U9301 (N_9301,N_3759,N_1308);
or U9302 (N_9302,N_2958,N_864);
xor U9303 (N_9303,N_2628,N_4200);
xor U9304 (N_9304,N_3888,N_3613);
nand U9305 (N_9305,N_4458,N_1034);
and U9306 (N_9306,N_4213,N_4840);
nand U9307 (N_9307,N_1764,N_2015);
and U9308 (N_9308,N_4342,N_2468);
or U9309 (N_9309,N_1848,N_2143);
or U9310 (N_9310,N_367,N_2304);
xor U9311 (N_9311,N_335,N_2007);
or U9312 (N_9312,N_4364,N_3794);
and U9313 (N_9313,N_3188,N_345);
and U9314 (N_9314,N_1407,N_3851);
xor U9315 (N_9315,N_3182,N_4146);
nor U9316 (N_9316,N_2641,N_4576);
xnor U9317 (N_9317,N_408,N_4155);
or U9318 (N_9318,N_161,N_1027);
xnor U9319 (N_9319,N_4176,N_2256);
or U9320 (N_9320,N_4805,N_1070);
nand U9321 (N_9321,N_3153,N_2525);
nor U9322 (N_9322,N_1570,N_3730);
xnor U9323 (N_9323,N_2297,N_160);
and U9324 (N_9324,N_2853,N_2510);
or U9325 (N_9325,N_4325,N_4545);
nor U9326 (N_9326,N_4720,N_2015);
and U9327 (N_9327,N_4597,N_3195);
nor U9328 (N_9328,N_1166,N_314);
nor U9329 (N_9329,N_1207,N_2475);
nand U9330 (N_9330,N_853,N_130);
nand U9331 (N_9331,N_452,N_4674);
nand U9332 (N_9332,N_2156,N_2901);
or U9333 (N_9333,N_4299,N_1572);
or U9334 (N_9334,N_4234,N_2530);
and U9335 (N_9335,N_1296,N_866);
nor U9336 (N_9336,N_2271,N_3846);
nand U9337 (N_9337,N_4429,N_4866);
and U9338 (N_9338,N_2880,N_4080);
and U9339 (N_9339,N_630,N_4376);
nor U9340 (N_9340,N_3223,N_4737);
or U9341 (N_9341,N_2706,N_4027);
nor U9342 (N_9342,N_4444,N_85);
or U9343 (N_9343,N_2127,N_89);
and U9344 (N_9344,N_4357,N_985);
nand U9345 (N_9345,N_1729,N_2279);
nor U9346 (N_9346,N_1392,N_3757);
xnor U9347 (N_9347,N_741,N_3228);
nor U9348 (N_9348,N_1862,N_1951);
or U9349 (N_9349,N_3217,N_4114);
and U9350 (N_9350,N_546,N_1433);
nand U9351 (N_9351,N_1667,N_4157);
nand U9352 (N_9352,N_3318,N_3174);
nor U9353 (N_9353,N_4535,N_433);
nand U9354 (N_9354,N_2337,N_2256);
and U9355 (N_9355,N_4794,N_3002);
nand U9356 (N_9356,N_3563,N_1025);
and U9357 (N_9357,N_3508,N_185);
nor U9358 (N_9358,N_3805,N_4367);
xnor U9359 (N_9359,N_2351,N_1467);
nor U9360 (N_9360,N_2701,N_2901);
nand U9361 (N_9361,N_2928,N_3928);
and U9362 (N_9362,N_1340,N_1733);
nand U9363 (N_9363,N_3613,N_2180);
nand U9364 (N_9364,N_3073,N_4866);
or U9365 (N_9365,N_1861,N_1049);
nor U9366 (N_9366,N_1476,N_3022);
and U9367 (N_9367,N_2108,N_4977);
nor U9368 (N_9368,N_3302,N_2806);
or U9369 (N_9369,N_3101,N_4295);
nand U9370 (N_9370,N_600,N_4691);
or U9371 (N_9371,N_352,N_2802);
or U9372 (N_9372,N_2968,N_2468);
nand U9373 (N_9373,N_4472,N_1883);
nor U9374 (N_9374,N_4872,N_4028);
xnor U9375 (N_9375,N_4996,N_3474);
xor U9376 (N_9376,N_2123,N_41);
and U9377 (N_9377,N_227,N_4732);
xnor U9378 (N_9378,N_416,N_3125);
and U9379 (N_9379,N_4771,N_1908);
nand U9380 (N_9380,N_104,N_2587);
xor U9381 (N_9381,N_4436,N_2840);
or U9382 (N_9382,N_2475,N_2063);
nor U9383 (N_9383,N_2544,N_699);
xor U9384 (N_9384,N_1846,N_4538);
and U9385 (N_9385,N_4037,N_3546);
nand U9386 (N_9386,N_4881,N_4231);
or U9387 (N_9387,N_978,N_2156);
or U9388 (N_9388,N_1103,N_201);
nand U9389 (N_9389,N_3748,N_1877);
or U9390 (N_9390,N_4719,N_150);
or U9391 (N_9391,N_3991,N_4973);
or U9392 (N_9392,N_3788,N_3231);
or U9393 (N_9393,N_3978,N_2504);
nand U9394 (N_9394,N_4467,N_2319);
xnor U9395 (N_9395,N_4135,N_3479);
xor U9396 (N_9396,N_1119,N_1955);
nor U9397 (N_9397,N_1646,N_4406);
and U9398 (N_9398,N_3433,N_1905);
or U9399 (N_9399,N_773,N_4170);
or U9400 (N_9400,N_537,N_3297);
and U9401 (N_9401,N_1587,N_2205);
xor U9402 (N_9402,N_3490,N_4958);
or U9403 (N_9403,N_2214,N_3261);
or U9404 (N_9404,N_555,N_2533);
xnor U9405 (N_9405,N_4847,N_3388);
nor U9406 (N_9406,N_1574,N_3790);
or U9407 (N_9407,N_2036,N_4039);
xnor U9408 (N_9408,N_3617,N_2408);
or U9409 (N_9409,N_813,N_4842);
nor U9410 (N_9410,N_3264,N_271);
nor U9411 (N_9411,N_1345,N_2056);
and U9412 (N_9412,N_1052,N_1123);
nor U9413 (N_9413,N_4445,N_1879);
nor U9414 (N_9414,N_4429,N_3134);
nand U9415 (N_9415,N_4742,N_4879);
or U9416 (N_9416,N_619,N_2881);
and U9417 (N_9417,N_2779,N_325);
nor U9418 (N_9418,N_2195,N_2645);
and U9419 (N_9419,N_949,N_3971);
nand U9420 (N_9420,N_997,N_667);
or U9421 (N_9421,N_583,N_3024);
xnor U9422 (N_9422,N_3010,N_3626);
or U9423 (N_9423,N_319,N_4123);
nand U9424 (N_9424,N_3998,N_1334);
nor U9425 (N_9425,N_3209,N_2310);
nor U9426 (N_9426,N_1901,N_1283);
nand U9427 (N_9427,N_167,N_4902);
or U9428 (N_9428,N_1560,N_591);
nand U9429 (N_9429,N_2005,N_1617);
or U9430 (N_9430,N_1427,N_876);
and U9431 (N_9431,N_3251,N_2378);
nor U9432 (N_9432,N_543,N_1240);
nor U9433 (N_9433,N_2229,N_4929);
nor U9434 (N_9434,N_2646,N_3436);
nand U9435 (N_9435,N_2339,N_41);
and U9436 (N_9436,N_3570,N_1065);
nor U9437 (N_9437,N_4566,N_930);
nor U9438 (N_9438,N_4360,N_3686);
nand U9439 (N_9439,N_3736,N_1909);
xnor U9440 (N_9440,N_221,N_2232);
or U9441 (N_9441,N_3727,N_4534);
nand U9442 (N_9442,N_1646,N_112);
or U9443 (N_9443,N_1461,N_590);
or U9444 (N_9444,N_2681,N_2703);
nor U9445 (N_9445,N_3402,N_3274);
nor U9446 (N_9446,N_2277,N_440);
and U9447 (N_9447,N_2714,N_3143);
nor U9448 (N_9448,N_1188,N_443);
nand U9449 (N_9449,N_1553,N_2384);
xnor U9450 (N_9450,N_1523,N_3345);
nor U9451 (N_9451,N_3957,N_2801);
or U9452 (N_9452,N_936,N_4139);
and U9453 (N_9453,N_1415,N_4092);
nand U9454 (N_9454,N_1953,N_1560);
nand U9455 (N_9455,N_4346,N_268);
nor U9456 (N_9456,N_509,N_1635);
or U9457 (N_9457,N_2296,N_951);
or U9458 (N_9458,N_1209,N_2724);
nand U9459 (N_9459,N_4600,N_3634);
nand U9460 (N_9460,N_1700,N_314);
nor U9461 (N_9461,N_4928,N_3053);
nor U9462 (N_9462,N_2239,N_3147);
xor U9463 (N_9463,N_606,N_3293);
and U9464 (N_9464,N_3323,N_3977);
or U9465 (N_9465,N_4997,N_1857);
or U9466 (N_9466,N_131,N_3712);
nand U9467 (N_9467,N_4347,N_3320);
nand U9468 (N_9468,N_3865,N_4539);
and U9469 (N_9469,N_3993,N_2788);
xor U9470 (N_9470,N_1930,N_2093);
nor U9471 (N_9471,N_4648,N_3373);
nand U9472 (N_9472,N_4331,N_4337);
nand U9473 (N_9473,N_2639,N_395);
nor U9474 (N_9474,N_820,N_1658);
and U9475 (N_9475,N_2762,N_4749);
nand U9476 (N_9476,N_3454,N_1961);
xor U9477 (N_9477,N_2696,N_1911);
nor U9478 (N_9478,N_4331,N_1742);
and U9479 (N_9479,N_108,N_2811);
and U9480 (N_9480,N_2717,N_3442);
or U9481 (N_9481,N_463,N_492);
xnor U9482 (N_9482,N_3826,N_3252);
or U9483 (N_9483,N_4217,N_4353);
nor U9484 (N_9484,N_1306,N_3832);
nand U9485 (N_9485,N_4100,N_203);
and U9486 (N_9486,N_1889,N_3062);
nand U9487 (N_9487,N_170,N_2263);
and U9488 (N_9488,N_3982,N_2058);
nand U9489 (N_9489,N_497,N_1219);
and U9490 (N_9490,N_1680,N_790);
and U9491 (N_9491,N_3836,N_3779);
and U9492 (N_9492,N_4734,N_3516);
or U9493 (N_9493,N_3598,N_4294);
xor U9494 (N_9494,N_689,N_1350);
and U9495 (N_9495,N_2570,N_223);
nand U9496 (N_9496,N_3010,N_2344);
and U9497 (N_9497,N_1517,N_4189);
nor U9498 (N_9498,N_259,N_862);
or U9499 (N_9499,N_619,N_558);
or U9500 (N_9500,N_781,N_1647);
or U9501 (N_9501,N_2957,N_499);
nor U9502 (N_9502,N_2695,N_3802);
nor U9503 (N_9503,N_1967,N_4502);
and U9504 (N_9504,N_4336,N_4866);
and U9505 (N_9505,N_3340,N_3234);
and U9506 (N_9506,N_1543,N_852);
and U9507 (N_9507,N_648,N_1317);
nor U9508 (N_9508,N_1947,N_437);
nor U9509 (N_9509,N_4995,N_1025);
or U9510 (N_9510,N_4779,N_403);
nand U9511 (N_9511,N_3622,N_1702);
nor U9512 (N_9512,N_1425,N_1475);
xor U9513 (N_9513,N_4538,N_4077);
or U9514 (N_9514,N_2556,N_2757);
and U9515 (N_9515,N_73,N_1236);
xor U9516 (N_9516,N_452,N_4098);
or U9517 (N_9517,N_3738,N_727);
and U9518 (N_9518,N_4182,N_1558);
nor U9519 (N_9519,N_1002,N_1027);
or U9520 (N_9520,N_3771,N_2051);
or U9521 (N_9521,N_2566,N_365);
or U9522 (N_9522,N_2837,N_906);
nand U9523 (N_9523,N_943,N_1308);
and U9524 (N_9524,N_412,N_926);
nor U9525 (N_9525,N_1479,N_504);
or U9526 (N_9526,N_1584,N_3044);
or U9527 (N_9527,N_367,N_866);
nand U9528 (N_9528,N_3038,N_2988);
or U9529 (N_9529,N_3564,N_4591);
nor U9530 (N_9530,N_2154,N_2121);
nor U9531 (N_9531,N_4178,N_666);
or U9532 (N_9532,N_2159,N_46);
nor U9533 (N_9533,N_1578,N_500);
xor U9534 (N_9534,N_2758,N_1);
nor U9535 (N_9535,N_3437,N_2981);
and U9536 (N_9536,N_3162,N_987);
and U9537 (N_9537,N_4192,N_4841);
or U9538 (N_9538,N_2662,N_3013);
and U9539 (N_9539,N_2685,N_975);
xor U9540 (N_9540,N_1286,N_2359);
xor U9541 (N_9541,N_4307,N_4596);
nor U9542 (N_9542,N_459,N_2098);
nor U9543 (N_9543,N_2834,N_222);
nand U9544 (N_9544,N_353,N_4611);
nand U9545 (N_9545,N_3523,N_1000);
or U9546 (N_9546,N_2757,N_2638);
and U9547 (N_9547,N_1638,N_741);
nor U9548 (N_9548,N_4287,N_4820);
or U9549 (N_9549,N_4943,N_4767);
or U9550 (N_9550,N_1896,N_3581);
or U9551 (N_9551,N_307,N_2246);
nor U9552 (N_9552,N_979,N_1370);
nand U9553 (N_9553,N_2505,N_833);
nand U9554 (N_9554,N_4272,N_2148);
xor U9555 (N_9555,N_3847,N_3418);
and U9556 (N_9556,N_3572,N_177);
xor U9557 (N_9557,N_4014,N_2997);
or U9558 (N_9558,N_2527,N_109);
nor U9559 (N_9559,N_4496,N_1659);
and U9560 (N_9560,N_4171,N_705);
nor U9561 (N_9561,N_768,N_1615);
nor U9562 (N_9562,N_3355,N_886);
nand U9563 (N_9563,N_2284,N_2119);
and U9564 (N_9564,N_4245,N_2812);
nor U9565 (N_9565,N_1980,N_1027);
or U9566 (N_9566,N_2716,N_3983);
xor U9567 (N_9567,N_2376,N_1349);
or U9568 (N_9568,N_253,N_3589);
nor U9569 (N_9569,N_2725,N_4952);
nand U9570 (N_9570,N_3440,N_4870);
nand U9571 (N_9571,N_3681,N_2965);
xnor U9572 (N_9572,N_1897,N_2380);
or U9573 (N_9573,N_1259,N_2476);
or U9574 (N_9574,N_4434,N_162);
nand U9575 (N_9575,N_484,N_347);
nor U9576 (N_9576,N_4130,N_4838);
nor U9577 (N_9577,N_2317,N_2477);
or U9578 (N_9578,N_1744,N_2797);
nor U9579 (N_9579,N_2459,N_1434);
and U9580 (N_9580,N_3400,N_3854);
and U9581 (N_9581,N_362,N_4943);
and U9582 (N_9582,N_2444,N_2467);
nand U9583 (N_9583,N_1853,N_3751);
nor U9584 (N_9584,N_3860,N_4446);
xor U9585 (N_9585,N_3788,N_2869);
nand U9586 (N_9586,N_3077,N_1398);
xnor U9587 (N_9587,N_3999,N_3777);
or U9588 (N_9588,N_4546,N_4660);
and U9589 (N_9589,N_3114,N_1715);
or U9590 (N_9590,N_366,N_4117);
and U9591 (N_9591,N_846,N_1872);
nand U9592 (N_9592,N_3598,N_4418);
nor U9593 (N_9593,N_3410,N_1502);
nand U9594 (N_9594,N_1001,N_4386);
or U9595 (N_9595,N_1750,N_796);
and U9596 (N_9596,N_1543,N_1309);
or U9597 (N_9597,N_2878,N_3844);
and U9598 (N_9598,N_3677,N_1204);
or U9599 (N_9599,N_1393,N_2448);
xnor U9600 (N_9600,N_3046,N_1219);
or U9601 (N_9601,N_1838,N_1590);
nand U9602 (N_9602,N_470,N_2644);
or U9603 (N_9603,N_4788,N_1011);
xor U9604 (N_9604,N_1426,N_489);
or U9605 (N_9605,N_1570,N_2546);
nand U9606 (N_9606,N_2109,N_1911);
nand U9607 (N_9607,N_1241,N_3267);
nand U9608 (N_9608,N_1579,N_2850);
xnor U9609 (N_9609,N_4310,N_3616);
or U9610 (N_9610,N_1633,N_4524);
or U9611 (N_9611,N_4486,N_3287);
nand U9612 (N_9612,N_3693,N_4310);
nand U9613 (N_9613,N_4209,N_941);
and U9614 (N_9614,N_3199,N_410);
and U9615 (N_9615,N_63,N_3355);
and U9616 (N_9616,N_837,N_4138);
and U9617 (N_9617,N_3320,N_4678);
nor U9618 (N_9618,N_2923,N_4243);
and U9619 (N_9619,N_2204,N_2180);
and U9620 (N_9620,N_1413,N_1066);
and U9621 (N_9621,N_2345,N_2325);
or U9622 (N_9622,N_2781,N_828);
and U9623 (N_9623,N_4305,N_2818);
nand U9624 (N_9624,N_2813,N_4391);
or U9625 (N_9625,N_3449,N_297);
nand U9626 (N_9626,N_3171,N_1576);
and U9627 (N_9627,N_1864,N_873);
nor U9628 (N_9628,N_1631,N_120);
nor U9629 (N_9629,N_213,N_3307);
nand U9630 (N_9630,N_1515,N_4393);
nand U9631 (N_9631,N_2270,N_3180);
nor U9632 (N_9632,N_1562,N_1515);
nand U9633 (N_9633,N_323,N_3175);
and U9634 (N_9634,N_3498,N_4675);
nand U9635 (N_9635,N_958,N_47);
and U9636 (N_9636,N_2552,N_2317);
or U9637 (N_9637,N_982,N_763);
or U9638 (N_9638,N_1983,N_2267);
nand U9639 (N_9639,N_3380,N_2421);
nor U9640 (N_9640,N_4248,N_865);
nor U9641 (N_9641,N_4678,N_4067);
nand U9642 (N_9642,N_3685,N_3802);
nand U9643 (N_9643,N_1373,N_15);
nor U9644 (N_9644,N_3065,N_680);
or U9645 (N_9645,N_2397,N_269);
nor U9646 (N_9646,N_937,N_3338);
nand U9647 (N_9647,N_3854,N_2579);
nor U9648 (N_9648,N_2185,N_1416);
nand U9649 (N_9649,N_352,N_1570);
nand U9650 (N_9650,N_537,N_2376);
nor U9651 (N_9651,N_2589,N_2821);
and U9652 (N_9652,N_3432,N_887);
or U9653 (N_9653,N_1806,N_568);
and U9654 (N_9654,N_1961,N_1837);
nand U9655 (N_9655,N_1566,N_883);
nand U9656 (N_9656,N_1462,N_3143);
xor U9657 (N_9657,N_1171,N_1633);
and U9658 (N_9658,N_3250,N_3685);
nor U9659 (N_9659,N_4490,N_3747);
xor U9660 (N_9660,N_4029,N_3030);
nand U9661 (N_9661,N_1993,N_441);
or U9662 (N_9662,N_1690,N_3883);
xnor U9663 (N_9663,N_4660,N_1675);
nor U9664 (N_9664,N_1628,N_2582);
or U9665 (N_9665,N_2596,N_1898);
nand U9666 (N_9666,N_3483,N_429);
xor U9667 (N_9667,N_970,N_4059);
and U9668 (N_9668,N_761,N_1287);
or U9669 (N_9669,N_4098,N_2562);
xnor U9670 (N_9670,N_926,N_2071);
nand U9671 (N_9671,N_2740,N_206);
nor U9672 (N_9672,N_1475,N_2073);
nor U9673 (N_9673,N_1357,N_855);
and U9674 (N_9674,N_3526,N_430);
nor U9675 (N_9675,N_2271,N_2771);
and U9676 (N_9676,N_4139,N_2791);
or U9677 (N_9677,N_3750,N_4514);
and U9678 (N_9678,N_4982,N_4543);
nand U9679 (N_9679,N_914,N_3210);
nand U9680 (N_9680,N_909,N_4077);
or U9681 (N_9681,N_314,N_4732);
nand U9682 (N_9682,N_2963,N_1453);
nand U9683 (N_9683,N_1262,N_903);
and U9684 (N_9684,N_1727,N_991);
nor U9685 (N_9685,N_4045,N_4796);
nor U9686 (N_9686,N_4179,N_825);
and U9687 (N_9687,N_4445,N_4993);
or U9688 (N_9688,N_4048,N_1020);
and U9689 (N_9689,N_1245,N_1389);
and U9690 (N_9690,N_3092,N_4272);
nor U9691 (N_9691,N_3111,N_2599);
and U9692 (N_9692,N_1486,N_2173);
or U9693 (N_9693,N_1557,N_2369);
or U9694 (N_9694,N_480,N_1166);
or U9695 (N_9695,N_3442,N_3599);
nand U9696 (N_9696,N_4851,N_1221);
and U9697 (N_9697,N_2498,N_1443);
or U9698 (N_9698,N_4623,N_713);
nand U9699 (N_9699,N_4724,N_3067);
nor U9700 (N_9700,N_1994,N_4449);
nor U9701 (N_9701,N_1283,N_2426);
nor U9702 (N_9702,N_3325,N_4397);
nor U9703 (N_9703,N_2253,N_2147);
and U9704 (N_9704,N_72,N_4704);
nand U9705 (N_9705,N_4940,N_1882);
nand U9706 (N_9706,N_4821,N_2431);
nor U9707 (N_9707,N_1701,N_3770);
and U9708 (N_9708,N_1701,N_4446);
nor U9709 (N_9709,N_2925,N_4359);
or U9710 (N_9710,N_2331,N_218);
or U9711 (N_9711,N_109,N_4549);
nor U9712 (N_9712,N_2689,N_368);
or U9713 (N_9713,N_2233,N_4127);
nand U9714 (N_9714,N_1257,N_1872);
or U9715 (N_9715,N_4317,N_861);
and U9716 (N_9716,N_3436,N_1034);
or U9717 (N_9717,N_4986,N_2378);
or U9718 (N_9718,N_2040,N_1128);
nand U9719 (N_9719,N_942,N_2442);
and U9720 (N_9720,N_785,N_148);
nor U9721 (N_9721,N_3667,N_4926);
nand U9722 (N_9722,N_2877,N_879);
nand U9723 (N_9723,N_4600,N_1363);
nor U9724 (N_9724,N_43,N_3897);
and U9725 (N_9725,N_3488,N_2253);
and U9726 (N_9726,N_4125,N_2506);
nand U9727 (N_9727,N_240,N_3220);
or U9728 (N_9728,N_1833,N_3324);
nand U9729 (N_9729,N_2948,N_805);
and U9730 (N_9730,N_1895,N_3550);
and U9731 (N_9731,N_2153,N_489);
xnor U9732 (N_9732,N_32,N_1831);
and U9733 (N_9733,N_1615,N_1826);
nand U9734 (N_9734,N_4963,N_4533);
and U9735 (N_9735,N_4854,N_2082);
and U9736 (N_9736,N_4573,N_3449);
nor U9737 (N_9737,N_2300,N_3831);
or U9738 (N_9738,N_4878,N_977);
or U9739 (N_9739,N_530,N_1550);
or U9740 (N_9740,N_3367,N_1398);
and U9741 (N_9741,N_2578,N_1452);
or U9742 (N_9742,N_4525,N_774);
nor U9743 (N_9743,N_2378,N_2510);
nor U9744 (N_9744,N_73,N_2253);
and U9745 (N_9745,N_4111,N_4749);
nand U9746 (N_9746,N_963,N_1122);
xnor U9747 (N_9747,N_976,N_2021);
nor U9748 (N_9748,N_2799,N_4766);
and U9749 (N_9749,N_1745,N_2239);
or U9750 (N_9750,N_2586,N_2824);
or U9751 (N_9751,N_393,N_363);
nor U9752 (N_9752,N_864,N_4864);
nor U9753 (N_9753,N_1876,N_3193);
nand U9754 (N_9754,N_1830,N_2238);
nor U9755 (N_9755,N_3469,N_3564);
nor U9756 (N_9756,N_1764,N_384);
and U9757 (N_9757,N_2279,N_3571);
and U9758 (N_9758,N_2490,N_3259);
or U9759 (N_9759,N_2039,N_4072);
nor U9760 (N_9760,N_3713,N_4069);
xnor U9761 (N_9761,N_3232,N_1766);
nand U9762 (N_9762,N_4994,N_470);
nand U9763 (N_9763,N_2084,N_2496);
nand U9764 (N_9764,N_3275,N_947);
or U9765 (N_9765,N_4878,N_1327);
nor U9766 (N_9766,N_4636,N_2617);
and U9767 (N_9767,N_4077,N_1000);
nand U9768 (N_9768,N_3459,N_1488);
or U9769 (N_9769,N_2841,N_1210);
and U9770 (N_9770,N_1037,N_4575);
or U9771 (N_9771,N_1810,N_3704);
or U9772 (N_9772,N_2328,N_3921);
nand U9773 (N_9773,N_3473,N_2986);
xor U9774 (N_9774,N_384,N_3921);
or U9775 (N_9775,N_955,N_3393);
nor U9776 (N_9776,N_3944,N_4992);
xor U9777 (N_9777,N_4674,N_1737);
or U9778 (N_9778,N_3843,N_950);
or U9779 (N_9779,N_4458,N_3200);
nand U9780 (N_9780,N_1975,N_237);
nor U9781 (N_9781,N_2947,N_720);
nor U9782 (N_9782,N_3919,N_1267);
and U9783 (N_9783,N_355,N_1456);
nand U9784 (N_9784,N_3942,N_1910);
xor U9785 (N_9785,N_4989,N_863);
nand U9786 (N_9786,N_3534,N_4258);
xor U9787 (N_9787,N_3612,N_4021);
nor U9788 (N_9788,N_4043,N_2337);
or U9789 (N_9789,N_4424,N_281);
nor U9790 (N_9790,N_623,N_4672);
or U9791 (N_9791,N_3328,N_1055);
nand U9792 (N_9792,N_3913,N_2469);
and U9793 (N_9793,N_3709,N_1755);
and U9794 (N_9794,N_813,N_4629);
nor U9795 (N_9795,N_3748,N_338);
nand U9796 (N_9796,N_4871,N_3710);
nand U9797 (N_9797,N_4027,N_1795);
xnor U9798 (N_9798,N_4690,N_1415);
xor U9799 (N_9799,N_1772,N_3202);
xor U9800 (N_9800,N_2880,N_1273);
or U9801 (N_9801,N_3690,N_1693);
nor U9802 (N_9802,N_2716,N_2944);
nand U9803 (N_9803,N_2411,N_1347);
or U9804 (N_9804,N_638,N_4848);
nor U9805 (N_9805,N_2385,N_4190);
nor U9806 (N_9806,N_2414,N_344);
xnor U9807 (N_9807,N_1701,N_2588);
nand U9808 (N_9808,N_3645,N_4125);
or U9809 (N_9809,N_3074,N_4566);
nand U9810 (N_9810,N_2775,N_1751);
nor U9811 (N_9811,N_4228,N_3367);
and U9812 (N_9812,N_3269,N_1269);
or U9813 (N_9813,N_4397,N_950);
or U9814 (N_9814,N_4077,N_1692);
xnor U9815 (N_9815,N_3364,N_2343);
nand U9816 (N_9816,N_4066,N_1047);
nand U9817 (N_9817,N_4260,N_3886);
or U9818 (N_9818,N_4697,N_2116);
or U9819 (N_9819,N_4647,N_3623);
nor U9820 (N_9820,N_3405,N_4487);
nand U9821 (N_9821,N_3450,N_4301);
or U9822 (N_9822,N_3393,N_968);
and U9823 (N_9823,N_422,N_914);
xor U9824 (N_9824,N_224,N_628);
or U9825 (N_9825,N_4171,N_4680);
xor U9826 (N_9826,N_2626,N_2218);
or U9827 (N_9827,N_2888,N_886);
nand U9828 (N_9828,N_3025,N_4187);
or U9829 (N_9829,N_1674,N_3061);
nor U9830 (N_9830,N_4428,N_2743);
nor U9831 (N_9831,N_444,N_777);
xnor U9832 (N_9832,N_4269,N_1469);
or U9833 (N_9833,N_3647,N_904);
nor U9834 (N_9834,N_3680,N_554);
nand U9835 (N_9835,N_538,N_680);
or U9836 (N_9836,N_2441,N_569);
or U9837 (N_9837,N_3555,N_1473);
or U9838 (N_9838,N_2878,N_3633);
or U9839 (N_9839,N_4356,N_598);
xor U9840 (N_9840,N_832,N_2396);
xnor U9841 (N_9841,N_4599,N_3132);
nand U9842 (N_9842,N_4675,N_4107);
xnor U9843 (N_9843,N_3357,N_2810);
nand U9844 (N_9844,N_2620,N_3347);
nand U9845 (N_9845,N_4673,N_4298);
nor U9846 (N_9846,N_274,N_4294);
nand U9847 (N_9847,N_708,N_3649);
and U9848 (N_9848,N_2173,N_3282);
nor U9849 (N_9849,N_1920,N_4317);
xor U9850 (N_9850,N_2211,N_4841);
xnor U9851 (N_9851,N_1837,N_2894);
and U9852 (N_9852,N_2636,N_4365);
and U9853 (N_9853,N_4604,N_4329);
or U9854 (N_9854,N_2784,N_3377);
nand U9855 (N_9855,N_3843,N_1111);
nand U9856 (N_9856,N_1470,N_206);
and U9857 (N_9857,N_3611,N_3445);
xor U9858 (N_9858,N_1971,N_4788);
nand U9859 (N_9859,N_3895,N_2238);
nand U9860 (N_9860,N_603,N_483);
or U9861 (N_9861,N_4400,N_3936);
nand U9862 (N_9862,N_26,N_818);
nand U9863 (N_9863,N_2141,N_1304);
xnor U9864 (N_9864,N_4701,N_4554);
and U9865 (N_9865,N_415,N_1500);
or U9866 (N_9866,N_1388,N_2685);
or U9867 (N_9867,N_3951,N_2960);
xnor U9868 (N_9868,N_4481,N_1749);
nand U9869 (N_9869,N_3894,N_3998);
xnor U9870 (N_9870,N_223,N_566);
nand U9871 (N_9871,N_2962,N_3866);
and U9872 (N_9872,N_1641,N_1525);
and U9873 (N_9873,N_1406,N_3214);
xnor U9874 (N_9874,N_4776,N_2693);
nor U9875 (N_9875,N_1458,N_304);
and U9876 (N_9876,N_1195,N_4152);
and U9877 (N_9877,N_131,N_694);
nand U9878 (N_9878,N_4227,N_2310);
and U9879 (N_9879,N_3785,N_4968);
or U9880 (N_9880,N_3243,N_4133);
and U9881 (N_9881,N_1035,N_6);
or U9882 (N_9882,N_1774,N_1435);
nor U9883 (N_9883,N_413,N_2262);
nand U9884 (N_9884,N_1082,N_3823);
and U9885 (N_9885,N_2923,N_3642);
and U9886 (N_9886,N_827,N_1151);
nand U9887 (N_9887,N_1486,N_4616);
and U9888 (N_9888,N_335,N_2560);
or U9889 (N_9889,N_2325,N_2615);
or U9890 (N_9890,N_3819,N_2543);
or U9891 (N_9891,N_657,N_826);
nor U9892 (N_9892,N_4463,N_1365);
nand U9893 (N_9893,N_1314,N_3098);
nand U9894 (N_9894,N_182,N_1624);
or U9895 (N_9895,N_1166,N_3798);
nor U9896 (N_9896,N_4711,N_4206);
or U9897 (N_9897,N_2132,N_4075);
nor U9898 (N_9898,N_4626,N_1016);
xnor U9899 (N_9899,N_2152,N_3622);
or U9900 (N_9900,N_3882,N_3431);
and U9901 (N_9901,N_2177,N_1419);
nor U9902 (N_9902,N_2355,N_1194);
and U9903 (N_9903,N_104,N_1714);
xor U9904 (N_9904,N_86,N_497);
nor U9905 (N_9905,N_388,N_1814);
or U9906 (N_9906,N_375,N_2125);
or U9907 (N_9907,N_341,N_4978);
nor U9908 (N_9908,N_2272,N_641);
or U9909 (N_9909,N_4474,N_1828);
nand U9910 (N_9910,N_904,N_4461);
or U9911 (N_9911,N_2806,N_1512);
and U9912 (N_9912,N_4218,N_3612);
or U9913 (N_9913,N_1877,N_1799);
xnor U9914 (N_9914,N_4682,N_4963);
or U9915 (N_9915,N_187,N_2525);
and U9916 (N_9916,N_1591,N_2575);
nor U9917 (N_9917,N_3069,N_4663);
nor U9918 (N_9918,N_1610,N_1220);
or U9919 (N_9919,N_1875,N_3025);
and U9920 (N_9920,N_3579,N_3035);
xor U9921 (N_9921,N_147,N_1540);
nand U9922 (N_9922,N_2607,N_1023);
and U9923 (N_9923,N_4719,N_3803);
nor U9924 (N_9924,N_1049,N_3456);
nor U9925 (N_9925,N_3904,N_3371);
and U9926 (N_9926,N_4038,N_3266);
nor U9927 (N_9927,N_3308,N_114);
or U9928 (N_9928,N_4150,N_2204);
nand U9929 (N_9929,N_3259,N_239);
or U9930 (N_9930,N_1886,N_4274);
or U9931 (N_9931,N_1253,N_2060);
or U9932 (N_9932,N_1156,N_4634);
or U9933 (N_9933,N_1353,N_3066);
nor U9934 (N_9934,N_265,N_2195);
nand U9935 (N_9935,N_3723,N_4515);
nor U9936 (N_9936,N_3836,N_1891);
or U9937 (N_9937,N_1998,N_1241);
xnor U9938 (N_9938,N_4679,N_171);
or U9939 (N_9939,N_2211,N_1819);
nand U9940 (N_9940,N_3542,N_2266);
nor U9941 (N_9941,N_1555,N_448);
xnor U9942 (N_9942,N_4886,N_1627);
nor U9943 (N_9943,N_2383,N_4044);
or U9944 (N_9944,N_4153,N_2230);
nor U9945 (N_9945,N_4781,N_2326);
nor U9946 (N_9946,N_2176,N_1796);
and U9947 (N_9947,N_1684,N_4795);
and U9948 (N_9948,N_4085,N_1650);
nor U9949 (N_9949,N_4692,N_4356);
nor U9950 (N_9950,N_3455,N_3669);
and U9951 (N_9951,N_4111,N_2360);
nor U9952 (N_9952,N_4424,N_4912);
nor U9953 (N_9953,N_1271,N_2820);
or U9954 (N_9954,N_2996,N_378);
nand U9955 (N_9955,N_2589,N_3042);
or U9956 (N_9956,N_2069,N_3872);
nor U9957 (N_9957,N_2456,N_1726);
nor U9958 (N_9958,N_1331,N_2914);
nor U9959 (N_9959,N_27,N_4404);
and U9960 (N_9960,N_4415,N_2484);
and U9961 (N_9961,N_3309,N_1061);
nor U9962 (N_9962,N_917,N_2713);
and U9963 (N_9963,N_1073,N_722);
and U9964 (N_9964,N_4423,N_3722);
nand U9965 (N_9965,N_4404,N_720);
nor U9966 (N_9966,N_2041,N_2891);
xor U9967 (N_9967,N_555,N_2295);
and U9968 (N_9968,N_2901,N_2191);
nor U9969 (N_9969,N_3430,N_4478);
nand U9970 (N_9970,N_4258,N_3193);
or U9971 (N_9971,N_4990,N_1018);
or U9972 (N_9972,N_352,N_3011);
or U9973 (N_9973,N_2392,N_1928);
and U9974 (N_9974,N_2547,N_3829);
nand U9975 (N_9975,N_4224,N_2916);
nand U9976 (N_9976,N_4918,N_2806);
nor U9977 (N_9977,N_2518,N_1077);
or U9978 (N_9978,N_2624,N_2968);
nor U9979 (N_9979,N_4020,N_3592);
nand U9980 (N_9980,N_1539,N_1267);
or U9981 (N_9981,N_52,N_3162);
nand U9982 (N_9982,N_2884,N_2448);
nor U9983 (N_9983,N_4737,N_3433);
or U9984 (N_9984,N_4768,N_3377);
and U9985 (N_9985,N_3869,N_294);
and U9986 (N_9986,N_1749,N_1934);
and U9987 (N_9987,N_2157,N_1513);
and U9988 (N_9988,N_4045,N_400);
nor U9989 (N_9989,N_3268,N_269);
and U9990 (N_9990,N_3632,N_3285);
or U9991 (N_9991,N_2751,N_4711);
or U9992 (N_9992,N_3824,N_4995);
or U9993 (N_9993,N_1897,N_33);
nand U9994 (N_9994,N_3472,N_926);
nor U9995 (N_9995,N_3974,N_1645);
and U9996 (N_9996,N_4934,N_484);
or U9997 (N_9997,N_1493,N_2877);
nand U9998 (N_9998,N_618,N_4698);
nand U9999 (N_9999,N_3084,N_4818);
and UO_0 (O_0,N_8012,N_7879);
or UO_1 (O_1,N_9356,N_7024);
nor UO_2 (O_2,N_7588,N_9414);
nand UO_3 (O_3,N_5782,N_8070);
nand UO_4 (O_4,N_6378,N_7292);
xor UO_5 (O_5,N_8405,N_7304);
and UO_6 (O_6,N_9489,N_5308);
or UO_7 (O_7,N_9315,N_9484);
nand UO_8 (O_8,N_7964,N_8426);
and UO_9 (O_9,N_9550,N_6549);
and UO_10 (O_10,N_7667,N_6930);
nor UO_11 (O_11,N_5894,N_8158);
xnor UO_12 (O_12,N_7689,N_8984);
or UO_13 (O_13,N_8679,N_9420);
nand UO_14 (O_14,N_8791,N_7945);
nand UO_15 (O_15,N_5649,N_6904);
nor UO_16 (O_16,N_6103,N_6403);
nor UO_17 (O_17,N_5364,N_7697);
and UO_18 (O_18,N_5487,N_5985);
or UO_19 (O_19,N_8120,N_5087);
nand UO_20 (O_20,N_9344,N_9435);
xor UO_21 (O_21,N_8360,N_8275);
nor UO_22 (O_22,N_6501,N_9505);
nand UO_23 (O_23,N_5523,N_7212);
or UO_24 (O_24,N_7156,N_8589);
nand UO_25 (O_25,N_5441,N_5241);
nor UO_26 (O_26,N_5422,N_7260);
and UO_27 (O_27,N_6025,N_8184);
nor UO_28 (O_28,N_8137,N_9201);
nor UO_29 (O_29,N_8031,N_7977);
and UO_30 (O_30,N_5993,N_9273);
and UO_31 (O_31,N_5330,N_5553);
nor UO_32 (O_32,N_6147,N_9860);
nand UO_33 (O_33,N_6674,N_5948);
nor UO_34 (O_34,N_9079,N_8785);
or UO_35 (O_35,N_7190,N_8923);
nor UO_36 (O_36,N_6543,N_7957);
and UO_37 (O_37,N_7046,N_5511);
or UO_38 (O_38,N_8382,N_8332);
and UO_39 (O_39,N_7493,N_7405);
nor UO_40 (O_40,N_8840,N_6879);
and UO_41 (O_41,N_5306,N_5675);
xor UO_42 (O_42,N_6503,N_9164);
and UO_43 (O_43,N_6089,N_7911);
and UO_44 (O_44,N_8674,N_6706);
or UO_45 (O_45,N_9274,N_5050);
and UO_46 (O_46,N_9293,N_6291);
nand UO_47 (O_47,N_6481,N_9297);
nand UO_48 (O_48,N_5752,N_9999);
nor UO_49 (O_49,N_8523,N_6317);
or UO_50 (O_50,N_8395,N_5869);
or UO_51 (O_51,N_8810,N_8000);
nand UO_52 (O_52,N_6387,N_9669);
nand UO_53 (O_53,N_8466,N_9354);
and UO_54 (O_54,N_5578,N_9869);
xor UO_55 (O_55,N_6487,N_8677);
nand UO_56 (O_56,N_8009,N_7927);
and UO_57 (O_57,N_9843,N_7522);
nand UO_58 (O_58,N_8565,N_9893);
nand UO_59 (O_59,N_8051,N_7648);
xnor UO_60 (O_60,N_7814,N_7258);
nand UO_61 (O_61,N_9982,N_9705);
nor UO_62 (O_62,N_8135,N_5100);
nor UO_63 (O_63,N_6705,N_5359);
or UO_64 (O_64,N_7221,N_8680);
nor UO_65 (O_65,N_9124,N_7103);
nand UO_66 (O_66,N_7871,N_8584);
or UO_67 (O_67,N_7775,N_7607);
nand UO_68 (O_68,N_8261,N_6167);
nor UO_69 (O_69,N_8488,N_9346);
nand UO_70 (O_70,N_7651,N_6539);
nand UO_71 (O_71,N_5824,N_5611);
nand UO_72 (O_72,N_7072,N_9062);
or UO_73 (O_73,N_6914,N_8111);
xor UO_74 (O_74,N_8618,N_6348);
or UO_75 (O_75,N_5607,N_6073);
or UO_76 (O_76,N_5692,N_9761);
nor UO_77 (O_77,N_9562,N_9607);
or UO_78 (O_78,N_9267,N_7666);
xnor UO_79 (O_79,N_8231,N_6666);
nor UO_80 (O_80,N_8781,N_9280);
xor UO_81 (O_81,N_6012,N_7891);
or UO_82 (O_82,N_6793,N_8538);
and UO_83 (O_83,N_9087,N_6280);
and UO_84 (O_84,N_6301,N_6082);
and UO_85 (O_85,N_7739,N_5632);
nor UO_86 (O_86,N_8559,N_6765);
or UO_87 (O_87,N_5189,N_5490);
nand UO_88 (O_88,N_7947,N_9865);
nand UO_89 (O_89,N_9196,N_5619);
nor UO_90 (O_90,N_7201,N_9624);
xor UO_91 (O_91,N_7662,N_8516);
xor UO_92 (O_92,N_8826,N_6965);
xnor UO_93 (O_93,N_9149,N_7468);
nand UO_94 (O_94,N_8703,N_5146);
nor UO_95 (O_95,N_9492,N_5081);
and UO_96 (O_96,N_9334,N_8470);
nand UO_97 (O_97,N_7723,N_5900);
nor UO_98 (O_98,N_7997,N_7823);
and UO_99 (O_99,N_9677,N_9307);
nor UO_100 (O_100,N_7913,N_8918);
nand UO_101 (O_101,N_5999,N_6847);
nand UO_102 (O_102,N_5449,N_6294);
nand UO_103 (O_103,N_9911,N_5740);
or UO_104 (O_104,N_5854,N_9218);
nand UO_105 (O_105,N_5056,N_8448);
and UO_106 (O_106,N_5135,N_7722);
nor UO_107 (O_107,N_9833,N_8525);
xor UO_108 (O_108,N_9212,N_8153);
nand UO_109 (O_109,N_9424,N_9173);
or UO_110 (O_110,N_9324,N_7684);
nand UO_111 (O_111,N_8287,N_8601);
and UO_112 (O_112,N_5904,N_9389);
or UO_113 (O_113,N_5398,N_6766);
nor UO_114 (O_114,N_7294,N_6232);
nor UO_115 (O_115,N_6165,N_6296);
and UO_116 (O_116,N_6537,N_6621);
xnor UO_117 (O_117,N_8002,N_7115);
or UO_118 (O_118,N_5925,N_8654);
xor UO_119 (O_119,N_5386,N_7415);
nand UO_120 (O_120,N_8539,N_5152);
or UO_121 (O_121,N_9581,N_6821);
or UO_122 (O_122,N_5097,N_7291);
nand UO_123 (O_123,N_9082,N_6480);
and UO_124 (O_124,N_8181,N_5975);
xor UO_125 (O_125,N_9836,N_8316);
and UO_126 (O_126,N_7381,N_8972);
and UO_127 (O_127,N_8229,N_8859);
or UO_128 (O_128,N_5158,N_5917);
and UO_129 (O_129,N_5745,N_5022);
nand UO_130 (O_130,N_9073,N_7113);
or UO_131 (O_131,N_6519,N_6863);
or UO_132 (O_132,N_8459,N_9875);
and UO_133 (O_133,N_9491,N_6606);
nand UO_134 (O_134,N_6907,N_8354);
or UO_135 (O_135,N_5210,N_7051);
and UO_136 (O_136,N_7663,N_6397);
or UO_137 (O_137,N_7540,N_7021);
xnor UO_138 (O_138,N_9631,N_6069);
nand UO_139 (O_139,N_5508,N_9286);
or UO_140 (O_140,N_8088,N_7626);
nor UO_141 (O_141,N_9125,N_7009);
and UO_142 (O_142,N_7066,N_7138);
nand UO_143 (O_143,N_6625,N_7821);
or UO_144 (O_144,N_5857,N_5633);
xor UO_145 (O_145,N_6675,N_6919);
and UO_146 (O_146,N_9377,N_8886);
and UO_147 (O_147,N_9907,N_9681);
nand UO_148 (O_148,N_5264,N_8064);
or UO_149 (O_149,N_7223,N_5242);
or UO_150 (O_150,N_8312,N_5101);
nor UO_151 (O_151,N_9158,N_6399);
nor UO_152 (O_152,N_5763,N_6521);
nand UO_153 (O_153,N_9202,N_5911);
or UO_154 (O_154,N_9449,N_8049);
xor UO_155 (O_155,N_8204,N_7316);
or UO_156 (O_156,N_6588,N_6080);
or UO_157 (O_157,N_7197,N_9983);
and UO_158 (O_158,N_9779,N_7311);
xnor UO_159 (O_159,N_7279,N_5122);
and UO_160 (O_160,N_8683,N_9830);
and UO_161 (O_161,N_9567,N_7457);
nand UO_162 (O_162,N_6159,N_7720);
nor UO_163 (O_163,N_9471,N_6191);
nor UO_164 (O_164,N_7153,N_8334);
nand UO_165 (O_165,N_6573,N_7685);
nor UO_166 (O_166,N_8369,N_9322);
xor UO_167 (O_167,N_8582,N_5301);
nor UO_168 (O_168,N_7826,N_8074);
and UO_169 (O_169,N_6457,N_7097);
and UO_170 (O_170,N_8082,N_8945);
nor UO_171 (O_171,N_8879,N_9966);
and UO_172 (O_172,N_8185,N_7025);
nor UO_173 (O_173,N_6314,N_9332);
or UO_174 (O_174,N_7375,N_8608);
and UO_175 (O_175,N_6175,N_8401);
xnor UO_176 (O_176,N_9994,N_5232);
or UO_177 (O_177,N_9885,N_9849);
or UO_178 (O_178,N_7598,N_7608);
or UO_179 (O_179,N_6100,N_6818);
and UO_180 (O_180,N_5378,N_5401);
nand UO_181 (O_181,N_5945,N_6297);
nor UO_182 (O_182,N_9047,N_7317);
or UO_183 (O_183,N_6926,N_7376);
nor UO_184 (O_184,N_6584,N_7277);
nor UO_185 (O_185,N_8750,N_9415);
nor UO_186 (O_186,N_9832,N_6307);
xnor UO_187 (O_187,N_9984,N_6791);
and UO_188 (O_188,N_9673,N_6047);
nand UO_189 (O_189,N_9752,N_8414);
nand UO_190 (O_190,N_9805,N_6023);
nand UO_191 (O_191,N_7170,N_9243);
xor UO_192 (O_192,N_5247,N_6347);
and UO_193 (O_193,N_8642,N_6238);
nand UO_194 (O_194,N_7090,N_8048);
nor UO_195 (O_195,N_8682,N_8764);
nand UO_196 (O_196,N_5551,N_7484);
xor UO_197 (O_197,N_7721,N_9958);
or UO_198 (O_198,N_9376,N_6439);
nor UO_199 (O_199,N_5762,N_7248);
or UO_200 (O_200,N_9373,N_5329);
and UO_201 (O_201,N_6361,N_9383);
or UO_202 (O_202,N_7851,N_8259);
and UO_203 (O_203,N_8991,N_5534);
or UO_204 (O_204,N_5557,N_6144);
and UO_205 (O_205,N_8609,N_6553);
nand UO_206 (O_206,N_5216,N_7318);
or UO_207 (O_207,N_5229,N_5750);
or UO_208 (O_208,N_5839,N_7654);
or UO_209 (O_209,N_9992,N_5093);
nand UO_210 (O_210,N_8001,N_5270);
nor UO_211 (O_211,N_5843,N_6933);
and UO_212 (O_212,N_5631,N_8892);
and UO_213 (O_213,N_6349,N_7265);
nand UO_214 (O_214,N_9342,N_6586);
nor UO_215 (O_215,N_8819,N_7218);
or UO_216 (O_216,N_7434,N_7994);
and UO_217 (O_217,N_7032,N_6611);
and UO_218 (O_218,N_5005,N_7554);
and UO_219 (O_219,N_8078,N_9565);
nor UO_220 (O_220,N_5908,N_6078);
and UO_221 (O_221,N_6613,N_5676);
nand UO_222 (O_222,N_8960,N_9181);
xor UO_223 (O_223,N_7022,N_5182);
and UO_224 (O_224,N_6287,N_6729);
nand UO_225 (O_225,N_5032,N_7846);
and UO_226 (O_226,N_7491,N_8822);
and UO_227 (O_227,N_8770,N_5126);
and UO_228 (O_228,N_9209,N_7233);
nor UO_229 (O_229,N_7623,N_6653);
or UO_230 (O_230,N_8508,N_5261);
or UO_231 (O_231,N_6156,N_6394);
nand UO_232 (O_232,N_5590,N_7989);
or UO_233 (O_233,N_8878,N_8604);
and UO_234 (O_234,N_7732,N_6043);
nor UO_235 (O_235,N_9458,N_9750);
or UO_236 (O_236,N_9936,N_7769);
nor UO_237 (O_237,N_8762,N_7409);
and UO_238 (O_238,N_5118,N_6900);
nor UO_239 (O_239,N_9846,N_9213);
nand UO_240 (O_240,N_9236,N_7859);
nor UO_241 (O_241,N_8710,N_7149);
xnor UO_242 (O_242,N_6090,N_5473);
or UO_243 (O_243,N_8147,N_5340);
nand UO_244 (O_244,N_5956,N_5098);
nor UO_245 (O_245,N_8748,N_8966);
nand UO_246 (O_246,N_6430,N_7668);
nand UO_247 (O_247,N_9066,N_6801);
and UO_248 (O_248,N_7637,N_5923);
and UO_249 (O_249,N_9039,N_7771);
nand UO_250 (O_250,N_9152,N_6035);
nor UO_251 (O_251,N_5655,N_7580);
and UO_252 (O_252,N_7781,N_5510);
xnor UO_253 (O_253,N_9440,N_6490);
nor UO_254 (O_254,N_6467,N_7041);
nor UO_255 (O_255,N_6970,N_5028);
nor UO_256 (O_256,N_7404,N_6835);
and UO_257 (O_257,N_5464,N_7935);
and UO_258 (O_258,N_9061,N_7897);
nor UO_259 (O_259,N_8653,N_7185);
and UO_260 (O_260,N_7147,N_5552);
nand UO_261 (O_261,N_5223,N_9818);
xor UO_262 (O_262,N_7225,N_6071);
xnor UO_263 (O_263,N_7787,N_7130);
nand UO_264 (O_264,N_7240,N_9520);
and UO_265 (O_265,N_7517,N_9538);
and UO_266 (O_266,N_6255,N_9452);
and UO_267 (O_267,N_5714,N_8665);
nand UO_268 (O_268,N_8694,N_6104);
or UO_269 (O_269,N_9000,N_6101);
nor UO_270 (O_270,N_8925,N_7282);
nand UO_271 (O_271,N_9593,N_6760);
and UO_272 (O_272,N_8747,N_7649);
nand UO_273 (O_273,N_8457,N_8243);
nor UO_274 (O_274,N_6665,N_7333);
or UO_275 (O_275,N_5379,N_8474);
and UO_276 (O_276,N_6817,N_7813);
xor UO_277 (O_277,N_9464,N_9825);
and UO_278 (O_278,N_7498,N_6527);
nand UO_279 (O_279,N_5339,N_6293);
and UO_280 (O_280,N_9877,N_7569);
nand UO_281 (O_281,N_8257,N_9914);
nand UO_282 (O_282,N_8323,N_9572);
nand UO_283 (O_283,N_6376,N_5990);
nand UO_284 (O_284,N_9627,N_7374);
xor UO_285 (O_285,N_7716,N_9518);
or UO_286 (O_286,N_8080,N_8828);
nor UO_287 (O_287,N_5610,N_7344);
or UO_288 (O_288,N_9549,N_6891);
or UO_289 (O_289,N_5479,N_5297);
nand UO_290 (O_290,N_8728,N_5801);
or UO_291 (O_291,N_8499,N_6044);
or UO_292 (O_292,N_8143,N_8417);
or UO_293 (O_293,N_8571,N_9569);
and UO_294 (O_294,N_6433,N_8362);
and UO_295 (O_295,N_9775,N_6806);
or UO_296 (O_296,N_6559,N_8438);
and UO_297 (O_297,N_5153,N_7572);
and UO_298 (O_298,N_9288,N_5370);
nor UO_299 (O_299,N_9205,N_7263);
nor UO_300 (O_300,N_7255,N_6846);
nor UO_301 (O_301,N_8739,N_7319);
nand UO_302 (O_302,N_6964,N_9887);
nand UO_303 (O_303,N_9544,N_7169);
nand UO_304 (O_304,N_7981,N_5157);
xor UO_305 (O_305,N_7208,N_9166);
nor UO_306 (O_306,N_5667,N_8979);
nand UO_307 (O_307,N_8733,N_9862);
nand UO_308 (O_308,N_7116,N_9847);
xnor UO_309 (O_309,N_7929,N_7015);
and UO_310 (O_310,N_7873,N_7872);
or UO_311 (O_311,N_6404,N_6188);
nor UO_312 (O_312,N_9309,N_9462);
nor UO_313 (O_313,N_8042,N_5391);
and UO_314 (O_314,N_9511,N_5731);
xnor UO_315 (O_315,N_7342,N_7520);
and UO_316 (O_316,N_6524,N_8037);
and UO_317 (O_317,N_5049,N_8795);
nor UO_318 (O_318,N_5568,N_6381);
nand UO_319 (O_319,N_7373,N_6673);
or UO_320 (O_320,N_7785,N_7980);
nand UO_321 (O_321,N_9400,N_8305);
and UO_322 (O_322,N_8114,N_6644);
xor UO_323 (O_323,N_5389,N_9519);
or UO_324 (O_324,N_7705,N_5325);
nand UO_325 (O_325,N_7958,N_8197);
and UO_326 (O_326,N_7386,N_8841);
and UO_327 (O_327,N_8377,N_9379);
and UO_328 (O_328,N_8522,N_8512);
nand UO_329 (O_329,N_6340,N_5285);
nor UO_330 (O_330,N_7952,N_7106);
or UO_331 (O_331,N_9251,N_8552);
or UO_332 (O_332,N_7600,N_6580);
nand UO_333 (O_333,N_5035,N_5616);
xnor UO_334 (O_334,N_6030,N_5503);
nor UO_335 (O_335,N_5711,N_9003);
or UO_336 (O_336,N_8328,N_5856);
nand UO_337 (O_337,N_9231,N_9408);
and UO_338 (O_338,N_5546,N_8357);
xor UO_339 (O_339,N_7121,N_9754);
and UO_340 (O_340,N_8329,N_5099);
nor UO_341 (O_341,N_8948,N_5674);
and UO_342 (O_342,N_9814,N_8232);
nor UO_343 (O_343,N_7440,N_7102);
xor UO_344 (O_344,N_8730,N_8929);
nor UO_345 (O_345,N_8743,N_8006);
nor UO_346 (O_346,N_7759,N_9405);
or UO_347 (O_347,N_9207,N_8560);
nand UO_348 (O_348,N_7647,N_5996);
and UO_349 (O_349,N_8515,N_7724);
or UO_350 (O_350,N_5978,N_7987);
and UO_351 (O_351,N_6802,N_8039);
and UO_352 (O_352,N_5159,N_7899);
nand UO_353 (O_353,N_9927,N_7533);
or UO_354 (O_354,N_8221,N_6018);
nand UO_355 (O_355,N_8806,N_5496);
and UO_356 (O_356,N_8524,N_8630);
and UO_357 (O_357,N_6852,N_8490);
nand UO_358 (O_358,N_7754,N_9160);
xor UO_359 (O_359,N_6230,N_6909);
or UO_360 (O_360,N_6257,N_9855);
nand UO_361 (O_361,N_5341,N_5226);
nor UO_362 (O_362,N_5424,N_9022);
nand UO_363 (O_363,N_5961,N_9823);
nor UO_364 (O_364,N_6488,N_6845);
nand UO_365 (O_365,N_5320,N_8430);
or UO_366 (O_366,N_5791,N_6321);
nor UO_367 (O_367,N_7207,N_7001);
and UO_368 (O_368,N_9745,N_9476);
nor UO_369 (O_369,N_6552,N_5295);
nor UO_370 (O_370,N_5236,N_7603);
or UO_371 (O_371,N_7486,N_6084);
and UO_372 (O_372,N_7108,N_6342);
and UO_373 (O_373,N_8635,N_6508);
or UO_374 (O_374,N_8327,N_5840);
or UO_375 (O_375,N_5031,N_7433);
and UO_376 (O_376,N_9521,N_8790);
nand UO_377 (O_377,N_9600,N_6911);
nor UO_378 (O_378,N_7313,N_8473);
and UO_379 (O_379,N_9672,N_6384);
nand UO_380 (O_380,N_9660,N_9465);
nand UO_381 (O_381,N_6708,N_6790);
nor UO_382 (O_382,N_5872,N_9799);
xor UO_383 (O_383,N_8077,N_6452);
nor UO_384 (O_384,N_5986,N_7003);
nand UO_385 (O_385,N_9555,N_6235);
or UO_386 (O_386,N_8541,N_8353);
and UO_387 (O_387,N_7475,N_8533);
xor UO_388 (O_388,N_8372,N_8534);
nand UO_389 (O_389,N_8390,N_7379);
nor UO_390 (O_390,N_6867,N_8659);
nor UO_391 (O_391,N_8449,N_6076);
nor UO_392 (O_392,N_6936,N_9014);
nand UO_393 (O_393,N_8977,N_6612);
nand UO_394 (O_394,N_7271,N_8947);
or UO_395 (O_395,N_7918,N_5882);
nand UO_396 (O_396,N_5994,N_9157);
nand UO_397 (O_397,N_9616,N_5493);
or UO_398 (O_398,N_9528,N_5151);
nand UO_399 (O_399,N_6008,N_6792);
nor UO_400 (O_400,N_6669,N_5432);
or UO_401 (O_401,N_6141,N_5058);
nor UO_402 (O_402,N_7079,N_9599);
or UO_403 (O_403,N_6724,N_9902);
nand UO_404 (O_404,N_7252,N_5434);
xor UO_405 (O_405,N_5304,N_9123);
nand UO_406 (O_406,N_6335,N_8707);
nand UO_407 (O_407,N_6275,N_9618);
nor UO_408 (O_408,N_6231,N_8939);
or UO_409 (O_409,N_8628,N_7880);
or UO_410 (O_410,N_6822,N_8647);
and UO_411 (O_411,N_9208,N_6465);
and UO_412 (O_412,N_6979,N_8375);
nor UO_413 (O_413,N_6341,N_8563);
nor UO_414 (O_414,N_9192,N_7237);
and UO_415 (O_415,N_6954,N_6574);
xnor UO_416 (O_416,N_7842,N_6594);
xnor UO_417 (O_417,N_8152,N_5959);
nand UO_418 (O_418,N_7591,N_6619);
and UO_419 (O_419,N_6661,N_5154);
or UO_420 (O_420,N_7866,N_5573);
nand UO_421 (O_421,N_7920,N_5516);
nand UO_422 (O_422,N_9988,N_6422);
nor UO_423 (O_423,N_9726,N_8467);
nand UO_424 (O_424,N_5417,N_7828);
or UO_425 (O_425,N_8548,N_7992);
and UO_426 (O_426,N_7464,N_9674);
nand UO_427 (O_427,N_9821,N_5439);
nor UO_428 (O_428,N_5597,N_6203);
and UO_429 (O_429,N_5561,N_7298);
nor UO_430 (O_430,N_5698,N_6648);
or UO_431 (O_431,N_8667,N_8050);
or UO_432 (O_432,N_6726,N_5070);
or UO_433 (O_433,N_6504,N_5788);
and UO_434 (O_434,N_6624,N_7861);
and UO_435 (O_435,N_7548,N_9502);
and UO_436 (O_436,N_9333,N_8897);
and UO_437 (O_437,N_9900,N_6310);
or UO_438 (O_438,N_8833,N_6476);
nand UO_439 (O_439,N_7395,N_8864);
and UO_440 (O_440,N_8767,N_8115);
or UO_441 (O_441,N_7951,N_8163);
and UO_442 (O_442,N_9883,N_9904);
and UO_443 (O_443,N_7605,N_9856);
nand UO_444 (O_444,N_5409,N_7299);
and UO_445 (O_445,N_8165,N_9220);
nor UO_446 (O_446,N_9179,N_9638);
and UO_447 (O_447,N_8471,N_8429);
and UO_448 (O_448,N_6785,N_8520);
and UO_449 (O_449,N_9522,N_7758);
or UO_450 (O_450,N_8567,N_8496);
nor UO_451 (O_451,N_9937,N_8260);
and UO_452 (O_452,N_6860,N_7076);
nand UO_453 (O_453,N_5292,N_6639);
or UO_454 (O_454,N_5583,N_8801);
and UO_455 (O_455,N_9276,N_5451);
or UO_456 (O_456,N_7061,N_8361);
nor UO_457 (O_457,N_6000,N_5746);
or UO_458 (O_458,N_7488,N_7806);
and UO_459 (O_459,N_5614,N_5928);
nand UO_460 (O_460,N_5890,N_9968);
or UO_461 (O_461,N_7627,N_9970);
and UO_462 (O_462,N_6782,N_5785);
and UO_463 (O_463,N_7753,N_8262);
and UO_464 (O_464,N_8451,N_7365);
or UO_465 (O_465,N_9174,N_8835);
nor UO_466 (O_466,N_8343,N_9253);
nand UO_467 (O_467,N_8445,N_6542);
nand UO_468 (O_468,N_9585,N_9788);
or UO_469 (O_469,N_8936,N_7583);
nand UO_470 (O_470,N_8107,N_7565);
and UO_471 (O_471,N_6991,N_9853);
xnor UO_472 (O_472,N_6289,N_6385);
nand UO_473 (O_473,N_9278,N_5663);
and UO_474 (O_474,N_7742,N_7619);
and UO_475 (O_475,N_9425,N_9637);
xnor UO_476 (O_476,N_6771,N_8681);
or UO_477 (O_477,N_5274,N_6416);
and UO_478 (O_478,N_9249,N_6239);
and UO_479 (O_479,N_5064,N_8128);
and UO_480 (O_480,N_7820,N_9026);
or UO_481 (O_481,N_9978,N_6053);
nor UO_482 (O_482,N_9738,N_5351);
or UO_483 (O_483,N_9765,N_6725);
xnor UO_484 (O_484,N_7681,N_7220);
xor UO_485 (O_485,N_6920,N_9995);
nand UO_486 (O_486,N_6005,N_7751);
xnor UO_487 (O_487,N_9359,N_7242);
nand UO_488 (O_488,N_5887,N_9271);
and UO_489 (O_489,N_6330,N_8792);
or UO_490 (O_490,N_5954,N_5574);
nor UO_491 (O_491,N_9279,N_5211);
nor UO_492 (O_492,N_9812,N_5388);
nand UO_493 (O_493,N_9153,N_8493);
nor UO_494 (O_494,N_9163,N_7043);
nand UO_495 (O_495,N_9496,N_7084);
nor UO_496 (O_496,N_5580,N_9686);
or UO_497 (O_497,N_9735,N_6253);
nand UO_498 (O_498,N_6987,N_6898);
or UO_499 (O_499,N_9041,N_8962);
nand UO_500 (O_500,N_9685,N_5278);
or UO_501 (O_501,N_5661,N_5565);
and UO_502 (O_502,N_9935,N_7564);
or UO_503 (O_503,N_6058,N_5832);
or UO_504 (O_504,N_9250,N_7161);
and UO_505 (O_505,N_8245,N_5068);
and UO_506 (O_506,N_7912,N_7810);
nand UO_507 (O_507,N_5541,N_5302);
or UO_508 (O_508,N_5192,N_6198);
and UO_509 (O_509,N_5767,N_7538);
and UO_510 (O_510,N_6016,N_9943);
nor UO_511 (O_511,N_5776,N_6704);
or UO_512 (O_512,N_8901,N_5392);
nand UO_513 (O_513,N_5199,N_5831);
nor UO_514 (O_514,N_5988,N_6595);
nor UO_515 (O_515,N_8469,N_7546);
or UO_516 (O_516,N_9967,N_8041);
and UO_517 (O_517,N_5443,N_5253);
or UO_518 (O_518,N_8823,N_9058);
nor UO_519 (O_519,N_7574,N_7216);
nand UO_520 (O_520,N_8514,N_9277);
and UO_521 (O_521,N_9859,N_5613);
or UO_522 (O_522,N_5455,N_6883);
xor UO_523 (O_523,N_8210,N_7111);
nor UO_524 (O_524,N_7808,N_6528);
xor UO_525 (O_525,N_8408,N_8834);
nor UO_526 (O_526,N_9177,N_6414);
nand UO_527 (O_527,N_5570,N_5132);
nand UO_528 (O_528,N_7518,N_9634);
and UO_529 (O_529,N_9070,N_5266);
or UO_530 (O_530,N_8862,N_9027);
nor UO_531 (O_531,N_7280,N_7482);
nand UO_532 (O_532,N_5437,N_8558);
nor UO_533 (O_533,N_6710,N_6662);
nor UO_534 (O_534,N_5425,N_6276);
or UO_535 (O_535,N_9835,N_8723);
nand UO_536 (O_536,N_8371,N_7057);
xnor UO_537 (O_537,N_5717,N_5082);
or UO_538 (O_538,N_9787,N_8176);
xnor UO_539 (O_539,N_5369,N_7359);
xor UO_540 (O_540,N_7228,N_6172);
nor UO_541 (O_541,N_6734,N_8004);
nor UO_542 (O_542,N_8922,N_6789);
nand UO_543 (O_543,N_7187,N_7809);
or UO_544 (O_544,N_8934,N_5463);
nor UO_545 (O_545,N_9341,N_9751);
nor UO_546 (O_546,N_6153,N_6855);
nor UO_547 (O_547,N_7701,N_8793);
nor UO_548 (O_548,N_8554,N_8017);
or UO_549 (O_549,N_8727,N_6748);
and UO_550 (O_550,N_8637,N_8249);
nor UO_551 (O_551,N_9078,N_7544);
nand UO_552 (O_552,N_6998,N_5271);
nand UO_553 (O_553,N_9168,N_6472);
and UO_554 (O_554,N_9770,N_8098);
nor UO_555 (O_555,N_6168,N_6819);
and UO_556 (O_556,N_9361,N_7174);
nand UO_557 (O_557,N_8660,N_8954);
or UO_558 (O_558,N_6677,N_6333);
nor UO_559 (O_559,N_9928,N_9199);
or UO_560 (O_560,N_8706,N_7983);
or UO_561 (O_561,N_5979,N_9116);
nand UO_562 (O_562,N_9328,N_9001);
and UO_563 (O_563,N_5920,N_6927);
nand UO_564 (O_564,N_5466,N_8950);
nand UO_565 (O_565,N_6383,N_9556);
nand UO_566 (O_566,N_7117,N_8842);
or UO_567 (O_567,N_9048,N_5595);
nand UO_568 (O_568,N_7528,N_5096);
nor UO_569 (O_569,N_6718,N_7553);
and UO_570 (O_570,N_7211,N_7924);
xor UO_571 (O_571,N_8942,N_9065);
nor UO_572 (O_572,N_6807,N_5348);
xnor UO_573 (O_573,N_6872,N_5310);
and UO_574 (O_574,N_6532,N_6423);
nand UO_575 (O_575,N_7587,N_7841);
nand UO_576 (O_576,N_8182,N_9470);
or UO_577 (O_577,N_6805,N_8865);
nand UO_578 (O_578,N_8695,N_6626);
nor UO_579 (O_579,N_8010,N_6854);
nand UO_580 (O_580,N_9789,N_8378);
and UO_581 (O_581,N_7016,N_5078);
nand UO_582 (O_582,N_6477,N_6114);
nand UO_583 (O_583,N_9986,N_6720);
or UO_584 (O_584,N_5475,N_9617);
or UO_585 (O_585,N_8588,N_7129);
nand UO_586 (O_586,N_5855,N_9386);
and UO_587 (O_587,N_7728,N_6795);
nand UO_588 (O_588,N_7214,N_5156);
and UO_589 (O_589,N_6269,N_6831);
nand UO_590 (O_590,N_6312,N_7290);
nor UO_591 (O_591,N_7243,N_9535);
nor UO_592 (O_592,N_9760,N_7633);
nor UO_593 (O_593,N_6097,N_6756);
nand UO_594 (O_594,N_6796,N_9284);
nor UO_595 (O_595,N_5799,N_5780);
or UO_596 (O_596,N_6794,N_7542);
and UO_597 (O_597,N_6956,N_6306);
or UO_598 (O_598,N_9411,N_9302);
nor UO_599 (O_599,N_5103,N_8626);
or UO_600 (O_600,N_9863,N_7960);
nand UO_601 (O_601,N_8495,N_5826);
and UO_602 (O_602,N_8265,N_7505);
nand UO_603 (O_603,N_9387,N_6451);
or UO_604 (O_604,N_6684,N_8745);
nand UO_605 (O_605,N_6489,N_6021);
nor UO_606 (O_606,N_5877,N_8113);
xnor UO_607 (O_607,N_8634,N_9238);
nor UO_608 (O_608,N_8215,N_8423);
xor UO_609 (O_609,N_5693,N_7549);
and UO_610 (O_610,N_8068,N_6195);
nor UO_611 (O_611,N_6632,N_6164);
nand UO_612 (O_612,N_6109,N_5336);
and UO_613 (O_613,N_5536,N_5940);
nor UO_614 (O_614,N_9711,N_9077);
and UO_615 (O_615,N_7232,N_7135);
nand UO_616 (O_616,N_5659,N_8851);
nand UO_617 (O_617,N_6246,N_8052);
nor UO_618 (O_618,N_6870,N_7105);
nor UO_619 (O_619,N_7641,N_9005);
and UO_620 (O_620,N_9852,N_7532);
and UO_621 (O_621,N_8536,N_7454);
nor UO_622 (O_622,N_5423,N_9382);
or UO_623 (O_623,N_7329,N_8132);
nor UO_624 (O_624,N_8839,N_7699);
and UO_625 (O_625,N_9296,N_6303);
nand UO_626 (O_626,N_6408,N_9203);
and UO_627 (O_627,N_9217,N_6514);
xnor UO_628 (O_628,N_5963,N_7350);
or UO_629 (O_629,N_8200,N_6120);
or UO_630 (O_630,N_8621,N_9460);
xnor UO_631 (O_631,N_5327,N_5520);
or UO_632 (O_632,N_7182,N_8765);
xnor UO_633 (O_633,N_8302,N_9102);
or UO_634 (O_634,N_8482,N_9719);
xor UO_635 (O_635,N_9628,N_9891);
and UO_636 (O_636,N_8615,N_8870);
nand UO_637 (O_637,N_6770,N_9827);
and UO_638 (O_638,N_5939,N_6407);
nand UO_639 (O_639,N_6150,N_6739);
nand UO_640 (O_640,N_6960,N_7602);
and UO_641 (O_641,N_6056,N_9432);
or UO_642 (O_642,N_5326,N_5203);
nand UO_643 (O_643,N_5006,N_5172);
nand UO_644 (O_644,N_7644,N_5059);
or UO_645 (O_645,N_6179,N_7177);
nand UO_646 (O_646,N_8250,N_9076);
nand UO_647 (O_647,N_6228,N_7403);
or UO_648 (O_648,N_9997,N_7217);
and UO_649 (O_649,N_6252,N_9498);
nor UO_650 (O_650,N_5964,N_9796);
xnor UO_651 (O_651,N_5499,N_5219);
nand UO_652 (O_652,N_6603,N_5491);
or UO_653 (O_653,N_6969,N_9870);
or UO_654 (O_654,N_9345,N_8148);
or UO_655 (O_655,N_6279,N_5615);
or UO_656 (O_656,N_5664,N_6903);
nand UO_657 (O_657,N_8638,N_8772);
and UO_658 (O_658,N_5640,N_7919);
and UO_659 (O_659,N_8097,N_6875);
nor UO_660 (O_660,N_7412,N_7870);
nor UO_661 (O_661,N_7539,N_9444);
and UO_662 (O_662,N_9579,N_9504);
and UO_663 (O_663,N_6941,N_6479);
or UO_664 (O_664,N_9819,N_6737);
xor UO_665 (O_665,N_6049,N_6997);
nand UO_666 (O_666,N_8829,N_5275);
nand UO_667 (O_667,N_5795,N_8072);
and UO_668 (O_668,N_5571,N_5248);
or UO_669 (O_669,N_9979,N_7736);
nor UO_670 (O_670,N_6157,N_6170);
or UO_671 (O_671,N_7334,N_9006);
or UO_672 (O_672,N_8217,N_9586);
and UO_673 (O_673,N_7816,N_5531);
nand UO_674 (O_674,N_5930,N_9558);
and UO_675 (O_675,N_8228,N_7713);
and UO_676 (O_676,N_8898,N_7002);
or UO_677 (O_677,N_5170,N_5629);
nand UO_678 (O_678,N_8356,N_7036);
nor UO_679 (O_679,N_5283,N_7708);
and UO_680 (O_680,N_8914,N_6572);
nand UO_681 (O_681,N_6251,N_6133);
nor UO_682 (O_682,N_6245,N_9588);
nor UO_683 (O_683,N_9723,N_6562);
nor UO_684 (O_684,N_9537,N_8941);
or UO_685 (O_685,N_5662,N_9516);
nand UO_686 (O_686,N_9268,N_8569);
or UO_687 (O_687,N_8059,N_7202);
and UO_688 (O_688,N_8754,N_7867);
xor UO_689 (O_689,N_9214,N_8347);
and UO_690 (O_690,N_5209,N_9539);
nor UO_691 (O_691,N_7402,N_9013);
and UO_692 (O_692,N_7896,N_6130);
nor UO_693 (O_693,N_8020,N_5608);
or UO_694 (O_694,N_8606,N_7140);
and UO_695 (O_695,N_5148,N_6469);
or UO_696 (O_696,N_7749,N_9120);
and UO_697 (O_697,N_5944,N_9225);
nor UO_698 (O_698,N_5272,N_7073);
or UO_699 (O_699,N_5017,N_9057);
nand UO_700 (O_700,N_9155,N_7577);
or UO_701 (O_701,N_8420,N_7288);
nand UO_702 (O_702,N_7437,N_6592);
xor UO_703 (O_703,N_8285,N_9461);
or UO_704 (O_704,N_8444,N_9651);
xor UO_705 (O_705,N_6216,N_6305);
nor UO_706 (O_706,N_5770,N_8439);
xnor UO_707 (O_707,N_5892,N_9305);
nor UO_708 (O_708,N_5651,N_6261);
nand UO_709 (O_709,N_5559,N_8752);
nor UO_710 (O_710,N_8857,N_6601);
xor UO_711 (O_711,N_8090,N_7895);
nand UO_712 (O_712,N_6171,N_5034);
nand UO_713 (O_713,N_6328,N_6531);
or UO_714 (O_714,N_8394,N_8882);
nand UO_715 (O_715,N_8597,N_7483);
or UO_716 (O_716,N_8106,N_8624);
and UO_717 (O_717,N_5803,N_7536);
or UO_718 (O_718,N_5815,N_6547);
and UO_719 (O_719,N_9609,N_7825);
and UO_720 (O_720,N_9533,N_9912);
xor UO_721 (O_721,N_5710,N_6703);
or UO_722 (O_722,N_7432,N_7698);
nand UO_723 (O_723,N_7527,N_6596);
and UO_724 (O_724,N_5102,N_7776);
and UO_725 (O_725,N_8478,N_8040);
nor UO_726 (O_726,N_7007,N_5263);
xor UO_727 (O_727,N_7339,N_7492);
nand UO_728 (O_728,N_8159,N_7890);
nand UO_729 (O_729,N_8226,N_6302);
nor UO_730 (O_730,N_8888,N_6869);
nand UO_731 (O_731,N_8413,N_8021);
or UO_732 (O_732,N_5588,N_6123);
nor UO_733 (O_733,N_7283,N_5941);
nor UO_734 (O_734,N_6513,N_7206);
or UO_735 (O_735,N_8374,N_7345);
nand UO_736 (O_736,N_8958,N_9500);
and UO_737 (O_737,N_5367,N_9285);
and UO_738 (O_738,N_9584,N_6735);
and UO_739 (O_739,N_8808,N_7620);
or UO_740 (O_740,N_6116,N_5528);
nand UO_741 (O_741,N_8251,N_5594);
and UO_742 (O_742,N_7418,N_5526);
nand UO_743 (O_743,N_9131,N_9097);
and UO_744 (O_744,N_6557,N_9699);
and UO_745 (O_745,N_6685,N_9525);
and UO_746 (O_746,N_6893,N_6282);
or UO_747 (O_747,N_8591,N_7253);
or UO_748 (O_748,N_9838,N_6811);
xor UO_749 (O_749,N_6316,N_9443);
nor UO_750 (O_750,N_9655,N_5609);
nand UO_751 (O_751,N_6740,N_8732);
or UO_752 (O_752,N_9230,N_9559);
and UO_753 (O_753,N_9729,N_5544);
nor UO_754 (O_754,N_6712,N_5547);
and UO_755 (O_755,N_8996,N_9955);
and UO_756 (O_756,N_8242,N_8345);
and UO_757 (O_757,N_8131,N_5349);
or UO_758 (O_758,N_9216,N_5634);
nor UO_759 (O_759,N_7609,N_9431);
xor UO_760 (O_760,N_8805,N_9032);
nand UO_761 (O_761,N_5952,N_9824);
nor UO_762 (O_762,N_7894,N_8561);
and UO_763 (O_763,N_6486,N_8944);
and UO_764 (O_764,N_5759,N_6299);
and UO_765 (O_765,N_7974,N_8649);
or UO_766 (O_766,N_8166,N_9036);
and UO_767 (O_767,N_6615,N_9241);
nand UO_768 (O_768,N_6077,N_6323);
nor UO_769 (O_769,N_6112,N_8341);
or UO_770 (O_770,N_6764,N_8288);
or UO_771 (O_771,N_6800,N_8056);
and UO_772 (O_772,N_5403,N_5808);
or UO_773 (O_773,N_9879,N_5060);
and UO_774 (O_774,N_5361,N_5042);
and UO_775 (O_775,N_9882,N_9138);
and UO_776 (O_776,N_6346,N_8081);
nand UO_777 (O_777,N_8593,N_9899);
nand UO_778 (O_778,N_5620,N_9365);
nor UO_779 (O_779,N_9394,N_9896);
and UO_780 (O_780,N_6787,N_8721);
or UO_781 (O_781,N_8435,N_5691);
and UO_782 (O_782,N_8156,N_6885);
nor UO_783 (O_783,N_9031,N_7822);
nand UO_784 (O_784,N_8779,N_7467);
xor UO_785 (O_785,N_9054,N_6931);
and UO_786 (O_786,N_7314,N_5053);
or UO_787 (O_787,N_9552,N_7931);
and UO_788 (O_788,N_9551,N_6442);
or UO_789 (O_789,N_9290,N_8183);
nand UO_790 (O_790,N_5935,N_6045);
nor UO_791 (O_791,N_6953,N_8136);
and UO_792 (O_792,N_7511,N_7428);
and UO_793 (O_793,N_7686,N_6410);
and UO_794 (O_794,N_7986,N_8544);
nor UO_795 (O_795,N_7165,N_6522);
xnor UO_796 (O_796,N_6618,N_8218);
nand UO_797 (O_797,N_7709,N_6236);
xor UO_798 (O_798,N_7738,N_6429);
or UO_799 (O_799,N_6695,N_8904);
nor UO_800 (O_800,N_8079,N_5566);
and UO_801 (O_801,N_7887,N_5690);
nor UO_802 (O_802,N_7932,N_6224);
nor UO_803 (O_803,N_7297,N_7677);
nor UO_804 (O_804,N_6354,N_7955);
nand UO_805 (O_805,N_9759,N_7599);
nor UO_806 (O_806,N_9646,N_7541);
nand UO_807 (O_807,N_7782,N_5769);
and UO_808 (O_808,N_7714,N_9619);
nand UO_809 (O_809,N_9156,N_7238);
or UO_810 (O_810,N_8246,N_7452);
nand UO_811 (O_811,N_7307,N_9954);
nor UO_812 (O_812,N_6446,N_7059);
or UO_813 (O_813,N_5593,N_9690);
xnor UO_814 (O_814,N_7864,N_8928);
nand UO_815 (O_815,N_8850,N_5864);
nand UO_816 (O_816,N_6448,N_5841);
and UO_817 (O_817,N_5467,N_5246);
xnor UO_818 (O_818,N_5825,N_6778);
nand UO_819 (O_819,N_6366,N_7293);
and UO_820 (O_820,N_7366,N_7547);
nand UO_821 (O_821,N_5265,N_5524);
nand UO_822 (O_822,N_7671,N_5813);
and UO_823 (O_823,N_7456,N_9680);
and UO_824 (O_824,N_8670,N_7400);
and UO_825 (O_825,N_8930,N_9985);
nand UO_826 (O_826,N_9917,N_7000);
nor UO_827 (O_827,N_5279,N_7323);
or UO_828 (O_828,N_7352,N_5572);
or UO_829 (O_829,N_7210,N_7680);
and UO_830 (O_830,N_7438,N_7306);
nand UO_831 (O_831,N_5471,N_7086);
and UO_832 (O_832,N_9959,N_8126);
xor UO_833 (O_833,N_9219,N_8669);
or UO_834 (O_834,N_6395,N_9033);
nand UO_835 (O_835,N_8428,N_8633);
nor UO_836 (O_836,N_8276,N_5281);
nand UO_837 (O_837,N_8980,N_7854);
xor UO_838 (O_838,N_7552,N_8932);
or UO_839 (O_839,N_5149,N_8555);
xnor UO_840 (O_840,N_5497,N_9380);
and UO_841 (O_841,N_8299,N_9069);
nor UO_842 (O_842,N_7038,N_8146);
nand UO_843 (O_843,N_5141,N_7606);
nand UO_844 (O_844,N_5238,N_9194);
or UO_845 (O_845,N_8281,N_5345);
or UO_846 (O_846,N_7683,N_9398);
and UO_847 (O_847,N_9118,N_6373);
xnor UO_848 (O_848,N_6836,N_6491);
and UO_849 (O_849,N_6754,N_7712);
and UO_850 (O_850,N_7089,N_7512);
and UO_851 (O_851,N_8691,N_6001);
nand UO_852 (O_852,N_8716,N_9121);
xnor UO_853 (O_853,N_9112,N_5637);
nor UO_854 (O_854,N_5987,N_9951);
nand UO_855 (O_855,N_5910,N_8172);
nand UO_856 (O_856,N_5657,N_9407);
or UO_857 (O_857,N_7407,N_9582);
and UO_858 (O_858,N_7324,N_9210);
nand UO_859 (O_859,N_5205,N_6474);
or UO_860 (O_860,N_5732,N_8998);
and UO_861 (O_861,N_5313,N_8383);
nor UO_862 (O_862,N_5137,N_6550);
nor UO_863 (O_863,N_5131,N_6088);
nor UO_864 (O_864,N_5718,N_9682);
or UO_865 (O_865,N_8603,N_8213);
or UO_866 (O_866,N_8013,N_5811);
and UO_867 (O_867,N_5445,N_8178);
nor UO_868 (O_868,N_8324,N_9601);
nor UO_869 (O_869,N_8844,N_8300);
and UO_870 (O_870,N_5668,N_7581);
or UO_871 (O_871,N_7151,N_5673);
or UO_872 (O_872,N_6617,N_7786);
and UO_873 (O_873,N_9109,N_6155);
or UO_874 (O_874,N_6738,N_6650);
or UO_875 (O_875,N_6105,N_5227);
nand UO_876 (O_876,N_8110,N_9509);
nor UO_877 (O_877,N_9010,N_6460);
and UO_878 (O_878,N_9529,N_9141);
nor UO_879 (O_879,N_5380,N_8786);
or UO_880 (O_880,N_5478,N_5560);
nor UO_881 (O_881,N_6176,N_9547);
and UO_882 (O_882,N_8751,N_5061);
nand UO_883 (O_883,N_6379,N_6694);
and UO_884 (O_884,N_9629,N_5778);
xnor UO_885 (O_885,N_6285,N_9137);
nor UO_886 (O_886,N_8812,N_7515);
xor UO_887 (O_887,N_9772,N_8935);
nor UO_888 (O_888,N_5418,N_5530);
nor UO_889 (O_889,N_7504,N_9244);
nor UO_890 (O_890,N_6402,N_5726);
or UO_891 (O_891,N_8891,N_9732);
and UO_892 (O_892,N_9517,N_8546);
and UO_893 (O_893,N_5228,N_8673);
or UO_894 (O_894,N_5666,N_8198);
and UO_895 (O_895,N_7408,N_5214);
nand UO_896 (O_896,N_6700,N_7907);
or UO_897 (O_897,N_7019,N_5067);
or UO_898 (O_898,N_7534,N_6343);
nor UO_899 (O_899,N_5243,N_9133);
and UO_900 (O_900,N_6946,N_8376);
or UO_901 (O_901,N_5372,N_8173);
nor UO_902 (O_902,N_6040,N_8067);
xnor UO_903 (O_903,N_8921,N_5175);
and UO_904 (O_904,N_7179,N_5876);
nand UO_905 (O_905,N_6751,N_8900);
nor UO_906 (O_906,N_9866,N_8130);
and UO_907 (O_907,N_8370,N_6918);
and UO_908 (O_908,N_6136,N_7362);
and UO_909 (O_909,N_7453,N_6362);
nor UO_910 (O_910,N_8650,N_6072);
nor UO_911 (O_911,N_6731,N_9915);
nand UO_912 (O_912,N_9266,N_6593);
nand UO_913 (O_913,N_7088,N_9466);
nor UO_914 (O_914,N_8581,N_8971);
and UO_915 (O_915,N_8885,N_9864);
nand UO_916 (O_916,N_6124,N_8510);
nor UO_917 (O_917,N_8322,N_6352);
xnor UO_918 (O_918,N_8392,N_9597);
and UO_919 (O_919,N_6019,N_8045);
nor UO_920 (O_920,N_7254,N_5089);
xor UO_921 (O_921,N_6221,N_8540);
xnor UO_922 (O_922,N_9508,N_5121);
and UO_923 (O_923,N_9294,N_5207);
or UO_924 (O_924,N_5092,N_5260);
and UO_925 (O_925,N_7249,N_5342);
or UO_926 (O_926,N_7118,N_8399);
xor UO_927 (O_927,N_8911,N_8254);
nand UO_928 (O_928,N_6672,N_5013);
xor UO_929 (O_929,N_7799,N_8709);
nor UO_930 (O_930,N_5991,N_6616);
nor UO_931 (O_931,N_9353,N_9176);
or UO_932 (O_932,N_8737,N_8044);
nor UO_933 (O_933,N_6767,N_9311);
nor UO_934 (O_934,N_8071,N_7031);
nand UO_935 (O_935,N_9226,N_7660);
nor UO_936 (O_936,N_5428,N_7327);
xor UO_937 (O_937,N_7604,N_6113);
nor UO_938 (O_938,N_7767,N_8600);
and UO_939 (O_939,N_9541,N_5922);
nor UO_940 (O_940,N_6281,N_5881);
nor UO_941 (O_941,N_5200,N_8297);
and UO_942 (O_942,N_7235,N_5343);
nand UO_943 (O_943,N_6733,N_5239);
xor UO_944 (O_944,N_7442,N_7150);
nor UO_945 (O_945,N_7910,N_8869);
nand UO_946 (O_946,N_6727,N_6545);
nor UO_947 (O_947,N_8411,N_6741);
nand UO_948 (O_948,N_6215,N_9991);
nor UO_949 (O_949,N_5179,N_7917);
nor UO_950 (O_950,N_9295,N_6719);
or UO_951 (O_951,N_5867,N_5875);
nand UO_952 (O_952,N_8389,N_6443);
nand UO_953 (O_953,N_8402,N_5617);
nor UO_954 (O_954,N_8759,N_6322);
and UO_955 (O_955,N_8675,N_8994);
nor UO_956 (O_956,N_9648,N_9423);
nand UO_957 (O_957,N_8872,N_5712);
or UO_958 (O_958,N_8827,N_8022);
nand UO_959 (O_959,N_7296,N_5899);
or UO_960 (O_960,N_8967,N_5076);
nor UO_961 (O_961,N_8734,N_5596);
nor UO_962 (O_962,N_5628,N_9797);
and UO_963 (O_963,N_6115,N_8269);
and UO_964 (O_964,N_7970,N_7494);
or UO_965 (O_965,N_5976,N_5115);
and UO_966 (O_966,N_5123,N_5772);
nand UO_967 (O_967,N_6320,N_8503);
nand UO_968 (O_968,N_9668,N_7501);
and UO_969 (O_969,N_9185,N_7968);
xnor UO_970 (O_970,N_9287,N_6538);
nand UO_971 (O_971,N_5249,N_9740);
or UO_972 (O_972,N_8122,N_5397);
nor UO_973 (O_973,N_8161,N_6938);
nor UO_974 (O_974,N_5702,N_8899);
or UO_975 (O_975,N_6478,N_7830);
and UO_976 (O_976,N_6081,N_8566);
or UO_977 (O_977,N_5684,N_9052);
xnor UO_978 (O_978,N_7940,N_9445);
or UO_979 (O_979,N_8489,N_6509);
nand UO_980 (O_980,N_6589,N_9884);
or UO_981 (O_981,N_5066,N_5010);
or UO_982 (O_982,N_9136,N_7083);
nand UO_983 (O_983,N_8460,N_6229);
or UO_984 (O_984,N_8019,N_9447);
nand UO_985 (O_985,N_8193,N_9110);
and UO_986 (O_986,N_6265,N_6959);
or UO_987 (O_987,N_6656,N_9753);
and UO_988 (O_988,N_7490,N_8738);
or UO_989 (O_989,N_7790,N_8203);
nand UO_990 (O_990,N_9612,N_7590);
and UO_991 (O_991,N_6696,N_7531);
nand UO_992 (O_992,N_9304,N_6249);
nand UO_993 (O_993,N_6412,N_9375);
or UO_994 (O_994,N_6313,N_5480);
and UO_995 (O_995,N_9437,N_7398);
xnor UO_996 (O_996,N_5290,N_8307);
nand UO_997 (O_997,N_5884,N_6850);
nand UO_998 (O_998,N_5233,N_9774);
or UO_999 (O_999,N_7636,N_7886);
nand UO_1000 (O_1000,N_7725,N_5395);
nor UO_1001 (O_1001,N_9029,N_7449);
nand UO_1002 (O_1002,N_9813,N_6512);
or UO_1003 (O_1003,N_6978,N_7503);
or UO_1004 (O_1004,N_8336,N_8645);
and UO_1005 (O_1005,N_8333,N_7812);
nand UO_1006 (O_1006,N_6406,N_6670);
nor UO_1007 (O_1007,N_7159,N_5055);
nand UO_1008 (O_1008,N_9457,N_9858);
and UO_1009 (O_1009,N_9749,N_8016);
and UO_1010 (O_1010,N_7330,N_5810);
nand UO_1011 (O_1011,N_9630,N_9564);
and UO_1012 (O_1012,N_5734,N_6463);
and UO_1013 (O_1013,N_7937,N_5408);
xnor UO_1014 (O_1014,N_7340,N_9190);
and UO_1015 (O_1015,N_5412,N_9247);
nand UO_1016 (O_1016,N_5833,N_6638);
or UO_1017 (O_1017,N_7014,N_8223);
nor UO_1018 (O_1018,N_8104,N_7961);
or UO_1019 (O_1019,N_5934,N_9596);
and UO_1020 (O_1020,N_9370,N_8112);
nand UO_1021 (O_1021,N_9794,N_9910);
and UO_1022 (O_1022,N_8816,N_6319);
nor UO_1023 (O_1023,N_7509,N_8623);
or UO_1024 (O_1024,N_6210,N_7514);
xnor UO_1025 (O_1025,N_6747,N_9901);
nor UO_1026 (O_1026,N_7848,N_6989);
and UO_1027 (O_1027,N_7261,N_7704);
and UO_1028 (O_1028,N_9283,N_8700);
and UO_1029 (O_1029,N_8303,N_7227);
or UO_1030 (O_1030,N_9675,N_9234);
nor UO_1031 (O_1031,N_9084,N_5779);
xor UO_1032 (O_1032,N_5143,N_6563);
nand UO_1033 (O_1033,N_5430,N_7757);
or UO_1034 (O_1034,N_8946,N_9422);
or UO_1035 (O_1035,N_6126,N_9117);
or UO_1036 (O_1036,N_5235,N_6915);
nand UO_1037 (O_1037,N_9925,N_5728);
or UO_1038 (O_1038,N_7476,N_9687);
nand UO_1039 (O_1039,N_6022,N_7657);
and UO_1040 (O_1040,N_6091,N_6240);
and UO_1041 (O_1041,N_5784,N_5998);
or UO_1042 (O_1042,N_9256,N_9946);
or UO_1043 (O_1043,N_6011,N_7752);
nand UO_1044 (O_1044,N_9200,N_5024);
or UO_1045 (O_1045,N_8629,N_6732);
xor UO_1046 (O_1046,N_5394,N_5802);
nor UO_1047 (O_1047,N_8556,N_7811);
nor UO_1048 (O_1048,N_9568,N_7141);
xor UO_1049 (O_1049,N_8290,N_8252);
or UO_1050 (O_1050,N_5470,N_5871);
nor UO_1051 (O_1051,N_6119,N_5468);
xor UO_1052 (O_1052,N_8848,N_5618);
nor UO_1053 (O_1053,N_7463,N_7908);
and UO_1054 (O_1054,N_8093,N_7764);
xnor UO_1055 (O_1055,N_5315,N_9867);
and UO_1056 (O_1056,N_5981,N_9493);
or UO_1057 (O_1057,N_6565,N_6174);
xor UO_1058 (O_1058,N_8121,N_7301);
and UO_1059 (O_1059,N_8598,N_5015);
xor UO_1060 (O_1060,N_7702,N_8442);
nor UO_1061 (O_1061,N_7624,N_9714);
or UO_1062 (O_1062,N_6635,N_9576);
xnor UO_1063 (O_1063,N_6728,N_8953);
nor UO_1064 (O_1064,N_8403,N_7585);
nor UO_1065 (O_1065,N_5707,N_5704);
xnor UO_1066 (O_1066,N_5870,N_5020);
nor UO_1067 (O_1067,N_7963,N_6367);
or UO_1068 (O_1068,N_6623,N_8368);
nand UO_1069 (O_1069,N_6986,N_8513);
nand UO_1070 (O_1070,N_6908,N_9105);
nand UO_1071 (O_1071,N_7341,N_8418);
nor UO_1072 (O_1072,N_6715,N_6878);
xnor UO_1073 (O_1073,N_8458,N_5919);
xor UO_1074 (O_1074,N_5517,N_9888);
and UO_1075 (O_1075,N_8219,N_9480);
nor UO_1076 (O_1076,N_5012,N_5742);
nor UO_1077 (O_1077,N_5626,N_7448);
or UO_1078 (O_1078,N_6304,N_7137);
xor UO_1079 (O_1079,N_8247,N_8970);
or UO_1080 (O_1080,N_8761,N_6212);
nand UO_1081 (O_1081,N_9183,N_6597);
nand UO_1082 (O_1082,N_9654,N_6816);
and UO_1083 (O_1083,N_5585,N_7838);
nand UO_1084 (O_1084,N_9543,N_6382);
nor UO_1085 (O_1085,N_5562,N_5116);
nand UO_1086 (O_1086,N_9920,N_5088);
and UO_1087 (O_1087,N_8625,N_5836);
nor UO_1088 (O_1088,N_9874,N_5601);
nand UO_1089 (O_1089,N_6516,N_7257);
nor UO_1090 (O_1090,N_8139,N_6350);
nand UO_1091 (O_1091,N_5931,N_6922);
and UO_1092 (O_1092,N_5624,N_9499);
xor UO_1093 (O_1093,N_5474,N_8572);
nor UO_1094 (O_1094,N_9237,N_8701);
xor UO_1095 (O_1095,N_9291,N_9347);
and UO_1096 (O_1096,N_7406,N_6431);
and UO_1097 (O_1097,N_6605,N_8472);
nand UO_1098 (O_1098,N_9459,N_6128);
nand UO_1099 (O_1099,N_8594,N_7507);
nand UO_1100 (O_1100,N_9303,N_6132);
nand UO_1101 (O_1101,N_6500,N_9456);
nor UO_1102 (O_1102,N_9695,N_8986);
nand UO_1103 (O_1103,N_7401,N_8893);
or UO_1104 (O_1104,N_9756,N_7364);
nand UO_1105 (O_1105,N_9418,N_9402);
nor UO_1106 (O_1106,N_7082,N_8811);
xnor UO_1107 (O_1107,N_9088,N_8500);
nand UO_1108 (O_1108,N_7093,N_9232);
xor UO_1109 (O_1109,N_7302,N_7100);
nor UO_1110 (O_1110,N_6571,N_6889);
nand UO_1111 (O_1111,N_9395,N_8735);
nor UO_1112 (O_1112,N_9790,N_9734);
nor UO_1113 (O_1113,N_6540,N_9656);
or UO_1114 (O_1114,N_5507,N_5830);
xor UO_1115 (O_1115,N_6561,N_7524);
and UO_1116 (O_1116,N_8545,N_9728);
nand UO_1117 (O_1117,N_5777,N_7010);
and UO_1118 (O_1118,N_9339,N_8306);
and UO_1119 (O_1119,N_9692,N_9242);
and UO_1120 (O_1120,N_7696,N_8272);
nor UO_1121 (O_1121,N_5706,N_9330);
or UO_1122 (O_1122,N_7993,N_6214);
nand UO_1123 (O_1123,N_7441,N_8446);
nand UO_1124 (O_1124,N_7560,N_5307);
xnor UO_1125 (O_1125,N_6055,N_6495);
or UO_1126 (O_1126,N_5007,N_5927);
nand UO_1127 (O_1127,N_6375,N_6812);
and UO_1128 (O_1128,N_5030,N_9906);
and UO_1129 (O_1129,N_5178,N_6928);
nand UO_1130 (O_1130,N_9049,N_7295);
and UO_1131 (O_1131,N_5077,N_6668);
xor UO_1132 (O_1132,N_8501,N_5110);
and UO_1133 (O_1133,N_9299,N_9557);
nor UO_1134 (O_1134,N_8641,N_9987);
nand UO_1135 (O_1135,N_6716,N_9355);
nand UO_1136 (O_1136,N_9260,N_5686);
nor UO_1137 (O_1137,N_5689,N_9406);
nand UO_1138 (O_1138,N_9050,N_5936);
nand UO_1139 (O_1139,N_7431,N_5817);
nand UO_1140 (O_1140,N_7516,N_9632);
nand UO_1141 (O_1141,N_6558,N_5730);
nor UO_1142 (O_1142,N_5206,N_6332);
or UO_1143 (O_1143,N_6149,N_6475);
nand UO_1144 (O_1144,N_9223,N_5323);
nor UO_1145 (O_1145,N_5735,N_9658);
nor UO_1146 (O_1146,N_9313,N_8729);
nand UO_1147 (O_1147,N_5965,N_8463);
and UO_1148 (O_1148,N_9793,N_9096);
and UO_1149 (O_1149,N_5317,N_6698);
and UO_1150 (O_1150,N_9327,N_6966);
nand UO_1151 (O_1151,N_6948,N_5368);
nand UO_1152 (O_1152,N_6493,N_6154);
and UO_1153 (O_1153,N_8613,N_7972);
and UO_1154 (O_1154,N_5184,N_7006);
xnor UO_1155 (O_1155,N_9715,N_6338);
nor UO_1156 (O_1156,N_6396,N_6197);
or UO_1157 (O_1157,N_9602,N_9055);
xnor UO_1158 (O_1158,N_6166,N_5130);
nor UO_1159 (O_1159,N_9886,N_8875);
or UO_1160 (O_1160,N_8617,N_5812);
xor UO_1161 (O_1161,N_5245,N_7726);
and UO_1162 (O_1162,N_7916,N_5043);
nand UO_1163 (O_1163,N_7101,N_7933);
and UO_1164 (O_1164,N_6692,N_8321);
nor UO_1165 (O_1165,N_7898,N_8101);
or UO_1166 (O_1166,N_5764,N_8917);
and UO_1167 (O_1167,N_8646,N_5041);
nand UO_1168 (O_1168,N_6848,N_7109);
nand UO_1169 (O_1169,N_5254,N_9645);
and UO_1170 (O_1170,N_6148,N_5191);
nor UO_1171 (O_1171,N_6746,N_5697);
nor UO_1172 (O_1172,N_5521,N_5344);
or UO_1173 (O_1173,N_8054,N_6193);
nor UO_1174 (O_1174,N_9495,N_8105);
nand UO_1175 (O_1175,N_9932,N_7763);
and UO_1176 (O_1176,N_9028,N_7966);
nor UO_1177 (O_1177,N_6939,N_7959);
nand UO_1178 (O_1178,N_5164,N_5682);
nand UO_1179 (O_1179,N_7578,N_5739);
xnor UO_1180 (O_1180,N_8244,N_6851);
or UO_1181 (O_1181,N_9965,N_6814);
nor UO_1182 (O_1182,N_7856,N_8926);
nor UO_1183 (O_1183,N_6940,N_7652);
and UO_1184 (O_1184,N_6651,N_6877);
xnor UO_1185 (O_1185,N_6074,N_8845);
xnor UO_1186 (O_1186,N_8990,N_5250);
nor UO_1187 (O_1187,N_8066,N_7419);
and UO_1188 (O_1188,N_7991,N_8631);
and UO_1189 (O_1189,N_8662,N_9701);
xnor UO_1190 (O_1190,N_8796,N_6730);
and UO_1191 (O_1191,N_6654,N_8313);
nor UO_1192 (O_1192,N_7774,N_6523);
nor UO_1193 (O_1193,N_8274,N_9366);
and UO_1194 (O_1194,N_7695,N_7436);
nand UO_1195 (O_1195,N_6952,N_5376);
or UO_1196 (O_1196,N_9016,N_9861);
nor UO_1197 (O_1197,N_5873,N_6094);
or UO_1198 (O_1198,N_6834,N_8578);
nand UO_1199 (O_1199,N_8949,N_5314);
or UO_1200 (O_1200,N_7416,N_9144);
or UO_1201 (O_1201,N_6688,N_6020);
and UO_1202 (O_1202,N_7278,N_7360);
and UO_1203 (O_1203,N_6582,N_6780);
nor UO_1204 (O_1204,N_7745,N_9506);
nand UO_1205 (O_1205,N_5069,N_7348);
nand UO_1206 (O_1206,N_9368,N_6690);
nor UO_1207 (O_1207,N_8083,N_5252);
nor UO_1208 (O_1208,N_8407,N_7017);
or UO_1209 (O_1209,N_9950,N_8763);
and UO_1210 (O_1210,N_9744,N_8492);
nor UO_1211 (O_1211,N_9684,N_9042);
nand UO_1212 (O_1212,N_9191,N_6983);
xnor UO_1213 (O_1213,N_8119,N_7178);
nor UO_1214 (O_1214,N_7794,N_9815);
nor UO_1215 (O_1215,N_9776,N_6614);
and UO_1216 (O_1216,N_6608,N_6426);
nor UO_1217 (O_1217,N_9222,N_5809);
or UO_1218 (O_1218,N_5371,N_8087);
or UO_1219 (O_1219,N_7584,N_9289);
and UO_1220 (O_1220,N_8852,N_5084);
or UO_1221 (O_1221,N_6896,N_7568);
or UO_1222 (O_1222,N_6947,N_5492);
or UO_1223 (O_1223,N_9448,N_5033);
nor UO_1224 (O_1224,N_7902,N_7901);
and UO_1225 (O_1225,N_8557,N_8861);
or UO_1226 (O_1226,N_5901,N_6925);
and UO_1227 (O_1227,N_7706,N_6336);
nand UO_1228 (O_1228,N_8672,N_6645);
xor UO_1229 (O_1229,N_8927,N_5258);
or UO_1230 (O_1230,N_8335,N_9074);
xnor UO_1231 (O_1231,N_7936,N_6386);
nand UO_1232 (O_1232,N_7616,N_5112);
xnor UO_1233 (O_1233,N_7239,N_7874);
or UO_1234 (O_1234,N_5083,N_8393);
and UO_1235 (O_1235,N_5193,N_5483);
xnor UO_1236 (O_1236,N_5003,N_9993);
or UO_1237 (O_1237,N_5280,N_5477);
nand UO_1238 (O_1238,N_6284,N_7458);
nor UO_1239 (O_1239,N_5955,N_7204);
or UO_1240 (O_1240,N_9007,N_6363);
or UO_1241 (O_1241,N_7250,N_8605);
xor UO_1242 (O_1242,N_5273,N_8652);
nand UO_1243 (O_1243,N_5602,N_7589);
nand UO_1244 (O_1244,N_8753,N_8397);
and UO_1245 (O_1245,N_5599,N_8693);
and UO_1246 (O_1246,N_7803,N_8337);
and UO_1247 (O_1247,N_9561,N_6248);
nor UO_1248 (O_1248,N_6663,N_7184);
or UO_1249 (O_1249,N_6808,N_8982);
xor UO_1250 (O_1250,N_9892,N_7573);
or UO_1251 (O_1251,N_6187,N_8883);
nor UO_1252 (O_1252,N_9479,N_6205);
nand UO_1253 (O_1253,N_8502,N_7367);
xnor UO_1254 (O_1254,N_7535,N_7331);
nor UO_1255 (O_1255,N_9030,N_7122);
nand UO_1256 (O_1256,N_7148,N_5969);
xor UO_1257 (O_1257,N_8619,N_8933);
nor UO_1258 (O_1258,N_6583,N_9246);
or UO_1259 (O_1259,N_7954,N_7067);
and UO_1260 (O_1260,N_9777,N_6950);
xnor UO_1261 (O_1261,N_6497,N_5548);
nand UO_1262 (O_1262,N_7496,N_9108);
or UO_1263 (O_1263,N_5074,N_9349);
or UO_1264 (O_1264,N_7643,N_6138);
nand UO_1265 (O_1265,N_9947,N_8585);
nor UO_1266 (O_1266,N_6459,N_6353);
nor UO_1267 (O_1267,N_9635,N_8993);
nor UO_1268 (O_1268,N_6994,N_8046);
nand UO_1269 (O_1269,N_6181,N_6200);
nand UO_1270 (O_1270,N_8359,N_6995);
nand UO_1271 (O_1271,N_8351,N_6518);
nor UO_1272 (O_1272,N_9807,N_7888);
and UO_1273 (O_1273,N_6036,N_8096);
and UO_1274 (O_1274,N_9075,N_7310);
and UO_1275 (O_1275,N_8778,N_8511);
nor UO_1276 (O_1276,N_9708,N_7850);
and UO_1277 (O_1277,N_5505,N_8133);
nand UO_1278 (O_1278,N_6420,N_7112);
and UO_1279 (O_1279,N_5563,N_8702);
nand UO_1280 (O_1280,N_6828,N_9688);
or UO_1281 (O_1281,N_6772,N_8699);
or UO_1282 (O_1282,N_6085,N_8705);
nand UO_1283 (O_1283,N_5150,N_9340);
nand UO_1284 (O_1284,N_9707,N_8849);
nand UO_1285 (O_1285,N_5090,N_7788);
xnor UO_1286 (O_1286,N_5180,N_7012);
and UO_1287 (O_1287,N_6419,N_7139);
xor UO_1288 (O_1288,N_7921,N_6371);
or UO_1289 (O_1289,N_5793,N_7925);
or UO_1290 (O_1290,N_9098,N_9727);
nand UO_1291 (O_1291,N_6267,N_8866);
or UO_1292 (O_1292,N_7962,N_5512);
xnor UO_1293 (O_1293,N_5377,N_7656);
nor UO_1294 (O_1294,N_8915,N_9921);
nor UO_1295 (O_1295,N_5120,N_7114);
nor UO_1296 (O_1296,N_5094,N_6699);
nor UO_1297 (O_1297,N_9828,N_8168);
nor UO_1298 (O_1298,N_7876,N_8570);
or UO_1299 (O_1299,N_6629,N_7559);
nand UO_1300 (O_1300,N_9512,N_5768);
or UO_1301 (O_1301,N_9961,N_6059);
nand UO_1302 (O_1302,N_7186,N_5582);
or UO_1303 (O_1303,N_8684,N_8815);
and UO_1304 (O_1304,N_5765,N_9417);
and UO_1305 (O_1305,N_8154,N_6517);
and UO_1306 (O_1306,N_8931,N_9964);
or UO_1307 (O_1307,N_8367,N_8187);
nor UO_1308 (O_1308,N_9890,N_5622);
nand UO_1309 (O_1309,N_5754,N_7832);
nor UO_1310 (O_1310,N_7383,N_6884);
and UO_1311 (O_1311,N_7368,N_5095);
nor UO_1312 (O_1312,N_8831,N_6041);
or UO_1313 (O_1313,N_8867,N_6681);
nor UO_1314 (O_1314,N_9487,N_8380);
or UO_1315 (O_1315,N_5289,N_5167);
or UO_1316 (O_1316,N_7965,N_5973);
nand UO_1317 (O_1317,N_9306,N_9169);
nand UO_1318 (O_1318,N_5845,N_5419);
or UO_1319 (O_1319,N_9595,N_5896);
xor UO_1320 (O_1320,N_7029,N_9298);
or UO_1321 (O_1321,N_6466,N_9165);
nor UO_1322 (O_1322,N_8595,N_7703);
and UO_1323 (O_1323,N_9996,N_5185);
or UO_1324 (O_1324,N_6849,N_8688);
xor UO_1325 (O_1325,N_6010,N_5106);
xor UO_1326 (O_1326,N_7414,N_8951);
nor UO_1327 (O_1327,N_6525,N_7661);
or UO_1328 (O_1328,N_8814,N_9107);
nand UO_1329 (O_1329,N_6207,N_9046);
xor UO_1330 (O_1330,N_7889,N_9570);
nor UO_1331 (O_1331,N_5677,N_5790);
xor UO_1332 (O_1332,N_9369,N_7551);
nor UO_1333 (O_1333,N_8836,N_5775);
nor UO_1334 (O_1334,N_8326,N_8320);
or UO_1335 (O_1335,N_6510,N_5481);
nand UO_1336 (O_1336,N_5781,N_6209);
nor UO_1337 (O_1337,N_9626,N_7869);
and UO_1338 (O_1338,N_8599,N_7731);
and UO_1339 (O_1339,N_7939,N_9515);
nand UO_1340 (O_1340,N_9248,N_6968);
nor UO_1341 (O_1341,N_8527,N_8301);
or UO_1342 (O_1342,N_5650,N_9257);
nor UO_1343 (O_1343,N_6024,N_8592);
nand UO_1344 (O_1344,N_8685,N_5733);
nand UO_1345 (O_1345,N_6689,N_7510);
and UO_1346 (O_1346,N_9497,N_9633);
and UO_1347 (O_1347,N_8784,N_5414);
nand UO_1348 (O_1348,N_9122,N_9566);
or UO_1349 (O_1349,N_5018,N_7506);
nand UO_1350 (O_1350,N_6658,N_8725);
nand UO_1351 (O_1351,N_9605,N_7091);
and UO_1352 (O_1352,N_8517,N_5286);
nor UO_1353 (O_1353,N_8476,N_5537);
nand UO_1354 (O_1354,N_7944,N_8271);
and UO_1355 (O_1355,N_5128,N_8464);
nor UO_1356 (O_1356,N_8129,N_5163);
or UO_1357 (O_1357,N_9371,N_6308);
and UO_1358 (O_1358,N_9020,N_6759);
and UO_1359 (O_1359,N_7740,N_7439);
and UO_1360 (O_1360,N_8887,N_9221);
nand UO_1361 (O_1361,N_6325,N_8535);
or UO_1362 (O_1362,N_6507,N_5144);
and UO_1363 (O_1363,N_5863,N_5267);
or UO_1364 (O_1364,N_7132,N_8206);
or UO_1365 (O_1365,N_7166,N_5555);
nand UO_1366 (O_1366,N_8782,N_7023);
or UO_1367 (O_1367,N_8043,N_9554);
nand UO_1368 (O_1368,N_6068,N_7312);
or UO_1369 (O_1369,N_6569,N_8192);
nand UO_1370 (O_1370,N_7030,N_8622);
and UO_1371 (O_1371,N_8212,N_7099);
and UO_1372 (O_1372,N_5783,N_5047);
nand UO_1373 (O_1373,N_9783,N_8719);
and UO_1374 (O_1374,N_9483,N_8919);
nand UO_1375 (O_1375,N_5457,N_6868);
nand UO_1376 (O_1376,N_8964,N_7026);
nor UO_1377 (O_1377,N_7477,N_9769);
and UO_1378 (O_1378,N_5079,N_5543);
nand UO_1379 (O_1379,N_5554,N_8029);
or UO_1380 (O_1380,N_9321,N_8712);
nand UO_1381 (O_1381,N_9140,N_8607);
nor UO_1382 (O_1382,N_7707,N_8698);
or UO_1383 (O_1383,N_8279,N_5623);
or UO_1384 (O_1384,N_9101,N_5950);
and UO_1385 (O_1385,N_7829,N_5436);
xnor UO_1386 (O_1386,N_6520,N_8880);
nand UO_1387 (O_1387,N_8663,N_7495);
xor UO_1388 (O_1388,N_6671,N_6473);
nand UO_1389 (O_1389,N_8053,N_8789);
or UO_1390 (O_1390,N_5381,N_9663);
nor UO_1391 (O_1391,N_5641,N_7796);
xor UO_1392 (O_1392,N_6173,N_7593);
xnor UO_1393 (O_1393,N_9530,N_9068);
nand UO_1394 (O_1394,N_8874,N_5316);
and UO_1395 (O_1395,N_8364,N_5652);
nand UO_1396 (O_1396,N_7679,N_9312);
nor UO_1397 (O_1397,N_7682,N_5413);
and UO_1398 (O_1398,N_6087,N_7048);
and UO_1399 (O_1399,N_8820,N_7575);
nor UO_1400 (O_1400,N_6392,N_6013);
nand UO_1401 (O_1401,N_6856,N_7783);
or UO_1402 (O_1402,N_7499,N_7044);
nand UO_1403 (O_1403,N_6762,N_8824);
or UO_1404 (O_1404,N_8963,N_6372);
xnor UO_1405 (O_1405,N_7556,N_9972);
nor UO_1406 (O_1406,N_5926,N_7284);
and UO_1407 (O_1407,N_7969,N_9782);
or UO_1408 (O_1408,N_9011,N_6761);
or UO_1409 (O_1409,N_9409,N_5814);
xor UO_1410 (O_1410,N_6060,N_8855);
or UO_1411 (O_1411,N_7286,N_6389);
xnor UO_1412 (O_1412,N_7934,N_8987);
nor UO_1413 (O_1413,N_8817,N_6934);
and UO_1414 (O_1414,N_9842,N_7473);
or UO_1415 (O_1415,N_5244,N_5410);
nand UO_1416 (O_1416,N_8975,N_5962);
and UO_1417 (O_1417,N_5194,N_8358);
and UO_1418 (O_1418,N_9857,N_8452);
and UO_1419 (O_1419,N_8258,N_6530);
xor UO_1420 (O_1420,N_5288,N_5635);
nor UO_1421 (O_1421,N_9531,N_9338);
and UO_1422 (O_1422,N_9002,N_7191);
or UO_1423 (O_1423,N_9012,N_6365);
and UO_1424 (O_1424,N_7802,N_7868);
nor UO_1425 (O_1425,N_7700,N_5037);
or UO_1426 (O_1426,N_8214,N_6286);
nand UO_1427 (O_1427,N_9167,N_5188);
nand UO_1428 (O_1428,N_7126,N_8768);
and UO_1429 (O_1429,N_6570,N_8758);
nand UO_1430 (O_1430,N_9942,N_8099);
and UO_1431 (O_1431,N_7343,N_9826);
and UO_1432 (O_1432,N_6401,N_5362);
xor UO_1433 (O_1433,N_9494,N_8117);
xor UO_1434 (O_1434,N_8190,N_6062);
or UO_1435 (O_1435,N_5044,N_7865);
nor UO_1436 (O_1436,N_6837,N_8575);
or UO_1437 (O_1437,N_7729,N_7640);
nand UO_1438 (O_1438,N_8286,N_5460);
or UO_1439 (O_1439,N_8632,N_8803);
or UO_1440 (O_1440,N_7194,N_7058);
nand UO_1441 (O_1441,N_5405,N_6418);
nand UO_1442 (O_1442,N_6070,N_6895);
nor UO_1443 (O_1443,N_9388,N_9733);
nor UO_1444 (O_1444,N_6981,N_6086);
nor UO_1445 (O_1445,N_7107,N_9913);
xnor UO_1446 (O_1446,N_8475,N_6498);
nor UO_1447 (O_1447,N_7630,N_7154);
nand UO_1448 (O_1448,N_5792,N_9233);
or UO_1449 (O_1449,N_9015,N_9004);
or UO_1450 (O_1450,N_6254,N_6295);
nand UO_1451 (O_1451,N_7338,N_9956);
nor UO_1452 (O_1452,N_5915,N_8248);
nand UO_1453 (O_1453,N_5045,N_5456);
or UO_1454 (O_1454,N_5485,N_7755);
or UO_1455 (O_1455,N_6106,N_5612);
nand UO_1456 (O_1456,N_6976,N_9809);
nor UO_1457 (O_1457,N_8027,N_5929);
and UO_1458 (O_1458,N_5171,N_6607);
nand UO_1459 (O_1459,N_8847,N_9706);
nor UO_1460 (O_1460,N_9503,N_7566);
and UO_1461 (O_1461,N_9329,N_8744);
nor UO_1462 (O_1462,N_6888,N_5458);
and UO_1463 (O_1463,N_8453,N_5119);
and UO_1464 (O_1464,N_6006,N_7843);
or UO_1465 (O_1465,N_6204,N_9712);
nand UO_1466 (O_1466,N_5197,N_7180);
nor UO_1467 (O_1467,N_9608,N_8868);
nand UO_1468 (O_1468,N_5721,N_5539);
or UO_1469 (O_1469,N_8381,N_9510);
xnor UO_1470 (O_1470,N_7673,N_9182);
nor UO_1471 (O_1471,N_9604,N_5909);
or UO_1472 (O_1472,N_6646,N_7160);
and UO_1473 (O_1473,N_5234,N_5838);
nor UO_1474 (O_1474,N_6554,N_9264);
nor UO_1475 (O_1475,N_5705,N_7144);
nor UO_1476 (O_1476,N_9700,N_9114);
or UO_1477 (O_1477,N_7904,N_6897);
or UO_1478 (O_1478,N_7845,N_7737);
and UO_1479 (O_1479,N_5658,N_9969);
nand UO_1480 (O_1480,N_7950,N_6456);
and UO_1481 (O_1481,N_5004,N_5751);
and UO_1482 (O_1482,N_7309,N_7760);
nand UO_1483 (O_1483,N_9594,N_5305);
and UO_1484 (O_1484,N_9081,N_6955);
nand UO_1485 (O_1485,N_6485,N_6225);
or UO_1486 (O_1486,N_5352,N_8689);
nor UO_1487 (O_1487,N_7055,N_6999);
nand UO_1488 (O_1488,N_7878,N_5186);
nor UO_1489 (O_1489,N_8195,N_8415);
nor UO_1490 (O_1490,N_8292,N_6827);
or UO_1491 (O_1491,N_8235,N_9650);
or UO_1492 (O_1492,N_8379,N_7519);
xnor UO_1493 (O_1493,N_9142,N_7040);
or UO_1494 (O_1494,N_9403,N_9957);
nor UO_1495 (O_1495,N_6315,N_9868);
or UO_1496 (O_1496,N_9154,N_5787);
nand UO_1497 (O_1497,N_9477,N_7267);
nand UO_1498 (O_1498,N_6327,N_7353);
nor UO_1499 (O_1499,N_5852,N_7857);
endmodule