module basic_750_5000_1000_5_levels_2xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
and U0 (N_0,In_92,In_707);
nor U1 (N_1,In_533,In_10);
or U2 (N_2,In_221,In_82);
nand U3 (N_3,In_376,In_634);
and U4 (N_4,In_66,In_249);
nor U5 (N_5,In_475,In_541);
and U6 (N_6,In_470,In_420);
or U7 (N_7,In_64,In_318);
nor U8 (N_8,In_214,In_642);
and U9 (N_9,In_286,In_621);
nand U10 (N_10,In_463,In_731);
and U11 (N_11,In_582,In_629);
nand U12 (N_12,In_122,In_157);
xor U13 (N_13,In_315,In_572);
nor U14 (N_14,In_511,In_303);
nand U15 (N_15,In_189,In_15);
nand U16 (N_16,In_253,In_4);
and U17 (N_17,In_121,In_523);
nor U18 (N_18,In_34,In_412);
nand U19 (N_19,In_273,In_219);
and U20 (N_20,In_738,In_123);
and U21 (N_21,In_696,In_9);
or U22 (N_22,In_468,In_643);
nor U23 (N_23,In_521,In_218);
nor U24 (N_24,In_649,In_314);
nand U25 (N_25,In_651,In_519);
nand U26 (N_26,In_40,In_14);
nand U27 (N_27,In_363,In_619);
and U28 (N_28,In_403,In_602);
or U29 (N_29,In_276,In_479);
nand U30 (N_30,In_236,In_311);
and U31 (N_31,In_383,In_553);
nor U32 (N_32,In_549,In_170);
and U33 (N_33,In_335,In_667);
and U34 (N_34,In_52,In_243);
and U35 (N_35,In_749,In_486);
nor U36 (N_36,In_517,In_647);
nand U37 (N_37,In_145,In_228);
or U38 (N_38,In_490,In_153);
nand U39 (N_39,In_510,In_319);
and U40 (N_40,In_63,In_266);
or U41 (N_41,In_258,In_560);
nor U42 (N_42,In_265,In_493);
nor U43 (N_43,In_155,In_718);
nor U44 (N_44,In_116,In_86);
or U45 (N_45,In_309,In_341);
nand U46 (N_46,In_618,In_728);
nor U47 (N_47,In_435,In_692);
nor U48 (N_48,In_178,In_736);
nand U49 (N_49,In_416,In_409);
xor U50 (N_50,In_543,In_106);
xor U51 (N_51,In_180,In_331);
and U52 (N_52,In_23,In_604);
and U53 (N_53,In_184,In_352);
or U54 (N_54,In_661,In_307);
and U55 (N_55,In_635,In_550);
and U56 (N_56,In_62,In_535);
and U57 (N_57,In_606,In_584);
or U58 (N_58,In_638,In_141);
nor U59 (N_59,In_93,In_520);
nor U60 (N_60,In_652,In_187);
nand U61 (N_61,In_77,In_226);
and U62 (N_62,In_353,In_746);
and U63 (N_63,In_298,In_264);
nand U64 (N_64,In_225,In_117);
and U65 (N_65,In_588,In_338);
nand U66 (N_66,In_300,In_85);
nand U67 (N_67,In_312,In_175);
nand U68 (N_68,In_415,In_748);
nor U69 (N_69,In_671,In_502);
and U70 (N_70,In_81,In_382);
nand U71 (N_71,In_613,In_1);
nor U72 (N_72,In_306,In_21);
nand U73 (N_73,In_43,In_135);
nand U74 (N_74,In_712,In_5);
nor U75 (N_75,In_204,In_200);
and U76 (N_76,In_326,In_385);
or U77 (N_77,In_744,In_125);
nand U78 (N_78,In_473,In_413);
nand U79 (N_79,In_102,In_609);
nor U80 (N_80,In_632,In_657);
nand U81 (N_81,In_732,In_239);
nor U82 (N_82,In_79,In_587);
nor U83 (N_83,In_656,In_626);
nor U84 (N_84,In_71,In_118);
and U85 (N_85,In_571,In_317);
and U86 (N_86,In_721,In_430);
nand U87 (N_87,In_710,In_150);
or U88 (N_88,In_148,In_589);
nor U89 (N_89,In_539,In_347);
and U90 (N_90,In_574,In_737);
or U91 (N_91,In_185,In_612);
nor U92 (N_92,In_288,In_97);
nor U93 (N_93,In_723,In_599);
nor U94 (N_94,In_50,In_408);
nand U95 (N_95,In_561,In_320);
or U96 (N_96,In_45,In_223);
xnor U97 (N_97,In_215,In_531);
or U98 (N_98,In_143,In_73);
or U99 (N_99,In_583,In_396);
nand U100 (N_100,In_480,In_322);
nor U101 (N_101,In_190,In_354);
or U102 (N_102,In_450,In_299);
or U103 (N_103,In_244,In_260);
nand U104 (N_104,In_358,In_467);
nand U105 (N_105,In_72,In_133);
nor U106 (N_106,In_270,In_384);
and U107 (N_107,In_329,In_207);
and U108 (N_108,In_213,In_351);
nand U109 (N_109,In_713,In_8);
nor U110 (N_110,In_41,In_459);
and U111 (N_111,In_679,In_705);
and U112 (N_112,In_30,In_147);
nand U113 (N_113,In_130,In_503);
and U114 (N_114,In_423,In_137);
xnor U115 (N_115,In_78,In_665);
nand U116 (N_116,In_367,In_378);
nor U117 (N_117,In_648,In_88);
nor U118 (N_118,In_287,In_685);
xnor U119 (N_119,In_110,In_578);
nand U120 (N_120,In_688,In_442);
nor U121 (N_121,In_682,In_53);
nor U122 (N_122,In_440,In_591);
or U123 (N_123,In_182,In_417);
nand U124 (N_124,In_24,In_340);
or U125 (N_125,In_568,In_527);
and U126 (N_126,In_162,In_74);
and U127 (N_127,In_172,In_136);
nand U128 (N_128,In_488,In_304);
and U129 (N_129,In_348,In_402);
nand U130 (N_130,In_538,In_603);
or U131 (N_131,In_144,In_212);
or U132 (N_132,In_485,In_529);
or U133 (N_133,In_70,In_58);
or U134 (N_134,In_637,In_103);
nor U135 (N_135,In_120,In_261);
nand U136 (N_136,In_158,In_372);
nor U137 (N_137,In_272,In_129);
nor U138 (N_138,In_366,In_727);
nor U139 (N_139,In_17,In_722);
or U140 (N_140,In_343,In_466);
nor U141 (N_141,In_641,In_655);
or U142 (N_142,In_391,In_188);
and U143 (N_143,In_499,In_166);
and U144 (N_144,In_460,In_379);
nand U145 (N_145,In_666,In_684);
and U146 (N_146,In_742,In_636);
and U147 (N_147,In_559,In_484);
and U148 (N_148,In_487,In_720);
nor U149 (N_149,In_428,In_482);
nor U150 (N_150,In_247,In_594);
or U151 (N_151,In_142,In_83);
nor U152 (N_152,In_154,In_336);
or U153 (N_153,In_210,In_557);
and U154 (N_154,In_234,In_191);
or U155 (N_155,In_169,In_13);
or U156 (N_156,In_699,In_427);
or U157 (N_157,In_80,In_414);
or U158 (N_158,In_230,In_76);
nand U159 (N_159,In_232,In_410);
nand U160 (N_160,In_168,In_434);
nand U161 (N_161,In_429,In_250);
or U162 (N_162,In_149,In_316);
and U163 (N_163,In_530,In_203);
and U164 (N_164,In_278,In_222);
nand U165 (N_165,In_703,In_217);
and U166 (N_166,In_548,In_674);
nor U167 (N_167,In_708,In_245);
and U168 (N_168,In_725,In_438);
nor U169 (N_169,In_262,In_202);
nor U170 (N_170,In_194,In_181);
or U171 (N_171,In_139,In_516);
nand U172 (N_172,In_44,In_60);
and U173 (N_173,In_160,In_254);
nand U174 (N_174,In_498,In_356);
and U175 (N_175,In_573,In_421);
nand U176 (N_176,In_663,In_151);
and U177 (N_177,In_330,In_6);
and U178 (N_178,In_595,In_325);
nand U179 (N_179,In_392,In_186);
and U180 (N_180,In_395,In_569);
or U181 (N_181,In_741,In_443);
or U182 (N_182,In_669,In_100);
and U183 (N_183,In_631,In_360);
nor U184 (N_184,In_528,In_394);
or U185 (N_185,In_419,In_49);
nand U186 (N_186,In_38,In_237);
and U187 (N_187,In_639,In_552);
nor U188 (N_188,In_259,In_592);
nor U189 (N_189,In_115,In_478);
nand U190 (N_190,In_282,In_422);
or U191 (N_191,In_747,In_471);
nor U192 (N_192,In_441,In_537);
or U193 (N_193,In_565,In_567);
nand U194 (N_194,In_193,In_179);
or U195 (N_195,In_691,In_579);
or U196 (N_196,In_233,In_167);
or U197 (N_197,In_20,In_701);
nor U198 (N_198,In_593,In_295);
or U199 (N_199,In_515,In_323);
and U200 (N_200,In_645,In_54);
or U201 (N_201,In_114,In_362);
or U202 (N_202,In_706,In_398);
nand U203 (N_203,In_28,In_365);
and U204 (N_204,In_0,In_644);
or U205 (N_205,In_159,In_534);
or U206 (N_206,In_183,In_390);
or U207 (N_207,In_346,In_19);
or U208 (N_208,In_623,In_734);
nor U209 (N_209,In_472,In_581);
nor U210 (N_210,In_280,In_281);
nand U211 (N_211,In_717,In_733);
nor U212 (N_212,In_451,In_289);
or U213 (N_213,In_205,In_715);
nor U214 (N_214,In_585,In_698);
and U215 (N_215,In_545,In_33);
nor U216 (N_216,In_640,In_206);
and U217 (N_217,In_681,In_524);
or U218 (N_218,In_597,In_37);
and U219 (N_219,In_628,In_601);
nand U220 (N_220,In_377,In_489);
nand U221 (N_221,In_658,In_55);
or U222 (N_222,In_461,In_405);
nand U223 (N_223,In_285,In_105);
or U224 (N_224,In_293,In_231);
nand U225 (N_225,In_453,In_371);
nand U226 (N_226,In_369,In_337);
and U227 (N_227,In_702,In_542);
and U228 (N_228,In_400,In_174);
or U229 (N_229,In_22,In_477);
and U230 (N_230,In_364,In_101);
or U231 (N_231,In_586,In_576);
or U232 (N_232,In_241,In_406);
nand U233 (N_233,In_263,In_610);
nor U234 (N_234,In_454,In_659);
and U235 (N_235,In_596,In_127);
or U236 (N_236,In_305,In_399);
or U237 (N_237,In_615,In_670);
nand U238 (N_238,In_693,In_124);
and U239 (N_239,In_455,In_495);
and U240 (N_240,In_598,In_558);
nor U241 (N_241,In_284,In_397);
and U242 (N_242,In_171,In_426);
or U243 (N_243,In_554,In_32);
or U244 (N_244,In_192,In_290);
nor U245 (N_245,In_474,In_374);
or U246 (N_246,In_302,In_238);
nor U247 (N_247,In_446,In_199);
or U248 (N_248,In_69,In_308);
or U249 (N_249,In_381,In_3);
nor U250 (N_250,In_68,In_506);
or U251 (N_251,In_507,In_126);
or U252 (N_252,In_458,In_313);
or U253 (N_253,In_449,In_673);
nor U254 (N_254,In_18,In_177);
xnor U255 (N_255,In_294,In_35);
and U256 (N_256,In_119,In_418);
nor U257 (N_257,In_107,In_140);
nand U258 (N_258,In_432,In_57);
or U259 (N_259,In_26,In_690);
and U260 (N_260,In_389,In_457);
nor U261 (N_261,In_512,In_252);
nand U262 (N_262,In_156,In_536);
or U263 (N_263,In_321,In_729);
nor U264 (N_264,In_227,In_689);
nor U265 (N_265,In_11,In_248);
nand U266 (N_266,In_653,In_7);
nor U267 (N_267,In_201,In_128);
nor U268 (N_268,In_445,In_256);
nand U269 (N_269,In_697,In_387);
nor U270 (N_270,In_431,In_373);
and U271 (N_271,In_494,In_739);
and U272 (N_272,In_476,In_611);
nor U273 (N_273,In_350,In_138);
and U274 (N_274,In_709,In_349);
and U275 (N_275,In_283,In_687);
xnor U276 (N_276,In_25,In_65);
nand U277 (N_277,In_555,In_633);
or U278 (N_278,In_163,In_492);
nand U279 (N_279,In_683,In_59);
or U280 (N_280,In_75,In_46);
or U281 (N_281,In_716,In_532);
nand U282 (N_282,In_452,In_447);
and U283 (N_283,In_342,In_2);
nand U284 (N_284,In_566,In_355);
nand U285 (N_285,In_570,In_575);
nor U286 (N_286,In_91,In_99);
nand U287 (N_287,In_745,In_562);
or U288 (N_288,In_161,In_146);
or U289 (N_289,In_109,In_401);
and U290 (N_290,In_513,In_439);
nor U291 (N_291,In_424,In_497);
and U292 (N_292,In_345,In_500);
nand U293 (N_293,In_84,In_607);
nand U294 (N_294,In_616,In_664);
and U295 (N_295,In_268,In_301);
or U296 (N_296,In_481,In_310);
xnor U297 (N_297,In_197,In_580);
or U298 (N_298,In_505,In_134);
xor U299 (N_299,In_334,In_87);
or U300 (N_300,In_292,In_235);
or U301 (N_301,In_208,In_333);
nand U302 (N_302,In_271,In_646);
nand U303 (N_303,In_164,In_483);
nor U304 (N_304,In_522,In_269);
nand U305 (N_305,In_242,In_98);
and U306 (N_306,In_388,In_393);
nor U307 (N_307,In_456,In_700);
and U308 (N_308,In_714,In_67);
nand U309 (N_309,In_719,In_686);
nand U310 (N_310,In_48,In_370);
xnor U311 (N_311,In_209,In_12);
nor U312 (N_312,In_496,In_332);
and U313 (N_313,In_614,In_678);
nand U314 (N_314,In_694,In_625);
nor U315 (N_315,In_743,In_407);
nor U316 (N_316,In_672,In_198);
and U317 (N_317,In_255,In_27);
nand U318 (N_318,In_469,In_267);
nand U319 (N_319,In_627,In_677);
nand U320 (N_320,In_246,In_726);
or U321 (N_321,In_95,In_375);
and U322 (N_322,In_96,In_131);
and U323 (N_323,In_108,In_257);
or U324 (N_324,In_29,In_444);
or U325 (N_325,In_104,In_176);
nand U326 (N_326,In_433,In_504);
nand U327 (N_327,In_508,In_386);
and U328 (N_328,In_622,In_16);
nor U329 (N_329,In_740,In_224);
nand U330 (N_330,In_425,In_617);
or U331 (N_331,In_89,In_251);
or U332 (N_332,In_296,In_509);
or U333 (N_333,In_695,In_112);
nor U334 (N_334,In_563,In_411);
nor U335 (N_335,In_436,In_540);
and U336 (N_336,In_380,In_464);
or U337 (N_337,In_547,In_546);
nor U338 (N_338,In_630,In_368);
or U339 (N_339,In_240,In_544);
nor U340 (N_340,In_551,In_195);
nor U341 (N_341,In_165,In_600);
nor U342 (N_342,In_624,In_36);
or U343 (N_343,In_277,In_650);
nor U344 (N_344,In_216,In_501);
or U345 (N_345,In_211,In_605);
or U346 (N_346,In_654,In_196);
nor U347 (N_347,In_327,In_404);
or U348 (N_348,In_357,In_339);
and U349 (N_349,In_608,In_39);
nor U350 (N_350,In_279,In_220);
xor U351 (N_351,In_324,In_675);
nor U352 (N_352,In_94,In_735);
xnor U353 (N_353,In_526,In_491);
nand U354 (N_354,In_361,In_328);
nor U355 (N_355,In_514,In_437);
nand U356 (N_356,In_152,In_56);
or U357 (N_357,In_132,In_42);
and U358 (N_358,In_711,In_462);
and U359 (N_359,In_518,In_676);
nor U360 (N_360,In_525,In_275);
nand U361 (N_361,In_31,In_448);
and U362 (N_362,In_577,In_47);
nor U363 (N_363,In_274,In_173);
nand U364 (N_364,In_359,In_730);
nand U365 (N_365,In_724,In_465);
and U366 (N_366,In_90,In_660);
and U367 (N_367,In_291,In_113);
nand U368 (N_368,In_297,In_564);
and U369 (N_369,In_556,In_668);
and U370 (N_370,In_61,In_51);
xnor U371 (N_371,In_229,In_111);
or U372 (N_372,In_680,In_344);
nor U373 (N_373,In_590,In_620);
and U374 (N_374,In_662,In_704);
nand U375 (N_375,In_448,In_423);
and U376 (N_376,In_356,In_541);
or U377 (N_377,In_594,In_292);
nor U378 (N_378,In_528,In_598);
or U379 (N_379,In_607,In_444);
or U380 (N_380,In_297,In_693);
or U381 (N_381,In_458,In_357);
nor U382 (N_382,In_695,In_636);
or U383 (N_383,In_27,In_588);
nand U384 (N_384,In_573,In_613);
or U385 (N_385,In_620,In_206);
or U386 (N_386,In_18,In_333);
nor U387 (N_387,In_649,In_670);
nor U388 (N_388,In_167,In_436);
or U389 (N_389,In_452,In_324);
or U390 (N_390,In_734,In_251);
xnor U391 (N_391,In_638,In_529);
and U392 (N_392,In_585,In_322);
and U393 (N_393,In_226,In_354);
and U394 (N_394,In_452,In_17);
nand U395 (N_395,In_34,In_274);
nor U396 (N_396,In_69,In_734);
nand U397 (N_397,In_150,In_249);
and U398 (N_398,In_471,In_389);
or U399 (N_399,In_620,In_540);
nor U400 (N_400,In_156,In_624);
and U401 (N_401,In_703,In_440);
nand U402 (N_402,In_348,In_454);
and U403 (N_403,In_671,In_599);
nor U404 (N_404,In_601,In_404);
and U405 (N_405,In_620,In_660);
and U406 (N_406,In_415,In_290);
and U407 (N_407,In_409,In_605);
nand U408 (N_408,In_514,In_398);
nor U409 (N_409,In_560,In_580);
xnor U410 (N_410,In_58,In_267);
nor U411 (N_411,In_258,In_281);
nor U412 (N_412,In_484,In_634);
or U413 (N_413,In_22,In_746);
or U414 (N_414,In_17,In_662);
or U415 (N_415,In_454,In_364);
and U416 (N_416,In_303,In_102);
or U417 (N_417,In_632,In_429);
and U418 (N_418,In_600,In_193);
nor U419 (N_419,In_646,In_617);
nand U420 (N_420,In_523,In_53);
nor U421 (N_421,In_108,In_112);
nand U422 (N_422,In_555,In_663);
nor U423 (N_423,In_291,In_211);
nor U424 (N_424,In_243,In_339);
or U425 (N_425,In_424,In_227);
or U426 (N_426,In_448,In_235);
and U427 (N_427,In_165,In_319);
and U428 (N_428,In_697,In_80);
or U429 (N_429,In_529,In_175);
nor U430 (N_430,In_647,In_505);
nor U431 (N_431,In_135,In_517);
and U432 (N_432,In_466,In_42);
nand U433 (N_433,In_218,In_487);
or U434 (N_434,In_701,In_327);
nor U435 (N_435,In_74,In_133);
or U436 (N_436,In_491,In_732);
nand U437 (N_437,In_155,In_300);
and U438 (N_438,In_661,In_697);
nand U439 (N_439,In_395,In_333);
and U440 (N_440,In_728,In_1);
or U441 (N_441,In_568,In_565);
nand U442 (N_442,In_638,In_184);
or U443 (N_443,In_539,In_372);
or U444 (N_444,In_96,In_246);
and U445 (N_445,In_275,In_257);
nand U446 (N_446,In_401,In_397);
and U447 (N_447,In_71,In_682);
or U448 (N_448,In_168,In_721);
nand U449 (N_449,In_307,In_371);
and U450 (N_450,In_564,In_552);
xnor U451 (N_451,In_459,In_267);
xor U452 (N_452,In_713,In_497);
or U453 (N_453,In_184,In_681);
nor U454 (N_454,In_350,In_724);
nor U455 (N_455,In_507,In_467);
and U456 (N_456,In_14,In_520);
and U457 (N_457,In_329,In_647);
nor U458 (N_458,In_722,In_745);
nor U459 (N_459,In_491,In_642);
nor U460 (N_460,In_370,In_123);
or U461 (N_461,In_101,In_703);
and U462 (N_462,In_542,In_168);
or U463 (N_463,In_664,In_498);
nand U464 (N_464,In_366,In_363);
nand U465 (N_465,In_355,In_337);
and U466 (N_466,In_687,In_35);
nor U467 (N_467,In_104,In_12);
nand U468 (N_468,In_133,In_187);
or U469 (N_469,In_547,In_544);
nand U470 (N_470,In_183,In_251);
nand U471 (N_471,In_60,In_511);
nand U472 (N_472,In_665,In_487);
nor U473 (N_473,In_538,In_410);
nand U474 (N_474,In_72,In_658);
nor U475 (N_475,In_279,In_213);
or U476 (N_476,In_679,In_462);
or U477 (N_477,In_659,In_658);
nand U478 (N_478,In_164,In_466);
nand U479 (N_479,In_462,In_574);
and U480 (N_480,In_307,In_422);
and U481 (N_481,In_522,In_110);
nand U482 (N_482,In_683,In_302);
nor U483 (N_483,In_302,In_300);
or U484 (N_484,In_35,In_306);
nor U485 (N_485,In_748,In_616);
nor U486 (N_486,In_394,In_538);
nand U487 (N_487,In_148,In_119);
nand U488 (N_488,In_278,In_353);
nor U489 (N_489,In_474,In_370);
nand U490 (N_490,In_111,In_563);
nor U491 (N_491,In_215,In_237);
nor U492 (N_492,In_68,In_533);
and U493 (N_493,In_109,In_204);
and U494 (N_494,In_560,In_328);
nor U495 (N_495,In_367,In_694);
or U496 (N_496,In_482,In_495);
and U497 (N_497,In_358,In_705);
xor U498 (N_498,In_735,In_563);
nor U499 (N_499,In_63,In_707);
nand U500 (N_500,In_440,In_114);
and U501 (N_501,In_238,In_61);
nor U502 (N_502,In_90,In_471);
or U503 (N_503,In_276,In_728);
nand U504 (N_504,In_542,In_104);
and U505 (N_505,In_675,In_426);
and U506 (N_506,In_640,In_103);
nand U507 (N_507,In_64,In_273);
or U508 (N_508,In_214,In_294);
or U509 (N_509,In_440,In_17);
nor U510 (N_510,In_387,In_653);
nor U511 (N_511,In_411,In_173);
or U512 (N_512,In_209,In_564);
and U513 (N_513,In_107,In_25);
nor U514 (N_514,In_287,In_438);
nor U515 (N_515,In_70,In_71);
and U516 (N_516,In_302,In_505);
or U517 (N_517,In_72,In_466);
nor U518 (N_518,In_79,In_438);
nand U519 (N_519,In_245,In_93);
or U520 (N_520,In_748,In_412);
nor U521 (N_521,In_277,In_395);
nor U522 (N_522,In_83,In_379);
xnor U523 (N_523,In_705,In_315);
nand U524 (N_524,In_400,In_618);
and U525 (N_525,In_544,In_74);
nor U526 (N_526,In_393,In_544);
or U527 (N_527,In_137,In_313);
nor U528 (N_528,In_284,In_544);
or U529 (N_529,In_672,In_492);
or U530 (N_530,In_85,In_69);
and U531 (N_531,In_352,In_667);
xor U532 (N_532,In_118,In_605);
nor U533 (N_533,In_304,In_700);
nor U534 (N_534,In_164,In_330);
and U535 (N_535,In_344,In_537);
nor U536 (N_536,In_747,In_68);
or U537 (N_537,In_554,In_568);
or U538 (N_538,In_439,In_679);
nor U539 (N_539,In_312,In_476);
nor U540 (N_540,In_58,In_533);
nand U541 (N_541,In_157,In_75);
nand U542 (N_542,In_675,In_563);
or U543 (N_543,In_524,In_37);
or U544 (N_544,In_129,In_693);
and U545 (N_545,In_452,In_134);
nand U546 (N_546,In_233,In_173);
or U547 (N_547,In_511,In_278);
or U548 (N_548,In_691,In_725);
nand U549 (N_549,In_530,In_385);
and U550 (N_550,In_303,In_130);
nor U551 (N_551,In_685,In_558);
or U552 (N_552,In_184,In_644);
nand U553 (N_553,In_654,In_568);
nand U554 (N_554,In_601,In_95);
nor U555 (N_555,In_649,In_326);
nor U556 (N_556,In_241,In_738);
nor U557 (N_557,In_656,In_389);
nand U558 (N_558,In_715,In_561);
nand U559 (N_559,In_116,In_642);
nand U560 (N_560,In_182,In_312);
and U561 (N_561,In_475,In_681);
nor U562 (N_562,In_560,In_738);
or U563 (N_563,In_41,In_498);
xnor U564 (N_564,In_579,In_21);
or U565 (N_565,In_661,In_442);
nand U566 (N_566,In_204,In_6);
nand U567 (N_567,In_439,In_49);
or U568 (N_568,In_343,In_572);
and U569 (N_569,In_365,In_540);
and U570 (N_570,In_663,In_461);
nor U571 (N_571,In_522,In_502);
xnor U572 (N_572,In_630,In_69);
nor U573 (N_573,In_92,In_408);
nor U574 (N_574,In_612,In_709);
nand U575 (N_575,In_273,In_34);
and U576 (N_576,In_201,In_665);
xor U577 (N_577,In_12,In_339);
xor U578 (N_578,In_274,In_709);
nand U579 (N_579,In_381,In_484);
nand U580 (N_580,In_375,In_630);
and U581 (N_581,In_138,In_39);
and U582 (N_582,In_460,In_66);
or U583 (N_583,In_206,In_271);
nor U584 (N_584,In_379,In_667);
nand U585 (N_585,In_281,In_82);
nand U586 (N_586,In_273,In_515);
nand U587 (N_587,In_479,In_217);
nor U588 (N_588,In_407,In_396);
and U589 (N_589,In_317,In_347);
nor U590 (N_590,In_350,In_92);
and U591 (N_591,In_430,In_329);
nand U592 (N_592,In_391,In_675);
nand U593 (N_593,In_299,In_97);
or U594 (N_594,In_567,In_595);
or U595 (N_595,In_488,In_82);
and U596 (N_596,In_634,In_710);
and U597 (N_597,In_33,In_360);
nand U598 (N_598,In_745,In_117);
and U599 (N_599,In_102,In_387);
or U600 (N_600,In_224,In_220);
or U601 (N_601,In_177,In_133);
nand U602 (N_602,In_122,In_71);
and U603 (N_603,In_273,In_201);
or U604 (N_604,In_15,In_646);
nand U605 (N_605,In_428,In_719);
nand U606 (N_606,In_40,In_155);
and U607 (N_607,In_361,In_441);
or U608 (N_608,In_519,In_244);
xor U609 (N_609,In_286,In_63);
or U610 (N_610,In_198,In_42);
and U611 (N_611,In_480,In_509);
or U612 (N_612,In_484,In_343);
or U613 (N_613,In_73,In_270);
and U614 (N_614,In_4,In_546);
nand U615 (N_615,In_404,In_488);
nor U616 (N_616,In_267,In_716);
nor U617 (N_617,In_397,In_380);
nor U618 (N_618,In_594,In_487);
nor U619 (N_619,In_423,In_175);
nor U620 (N_620,In_209,In_353);
or U621 (N_621,In_170,In_516);
nand U622 (N_622,In_495,In_367);
and U623 (N_623,In_226,In_595);
and U624 (N_624,In_609,In_516);
nand U625 (N_625,In_312,In_403);
and U626 (N_626,In_278,In_643);
nand U627 (N_627,In_747,In_27);
nand U628 (N_628,In_108,In_236);
nand U629 (N_629,In_278,In_597);
or U630 (N_630,In_228,In_395);
nor U631 (N_631,In_607,In_506);
nand U632 (N_632,In_31,In_130);
and U633 (N_633,In_419,In_542);
or U634 (N_634,In_282,In_303);
or U635 (N_635,In_164,In_193);
nand U636 (N_636,In_197,In_195);
and U637 (N_637,In_367,In_639);
nand U638 (N_638,In_469,In_204);
nand U639 (N_639,In_499,In_474);
xnor U640 (N_640,In_518,In_235);
nand U641 (N_641,In_599,In_241);
or U642 (N_642,In_79,In_106);
nand U643 (N_643,In_458,In_15);
nor U644 (N_644,In_603,In_111);
nor U645 (N_645,In_673,In_623);
nor U646 (N_646,In_225,In_384);
nand U647 (N_647,In_63,In_422);
or U648 (N_648,In_466,In_69);
and U649 (N_649,In_322,In_657);
and U650 (N_650,In_650,In_693);
nand U651 (N_651,In_385,In_397);
and U652 (N_652,In_494,In_422);
nor U653 (N_653,In_86,In_6);
and U654 (N_654,In_374,In_398);
and U655 (N_655,In_53,In_61);
nor U656 (N_656,In_646,In_451);
xnor U657 (N_657,In_17,In_468);
and U658 (N_658,In_514,In_419);
and U659 (N_659,In_389,In_403);
nand U660 (N_660,In_273,In_360);
or U661 (N_661,In_544,In_603);
or U662 (N_662,In_451,In_142);
nor U663 (N_663,In_745,In_68);
or U664 (N_664,In_237,In_274);
and U665 (N_665,In_243,In_284);
nor U666 (N_666,In_651,In_367);
nor U667 (N_667,In_230,In_533);
and U668 (N_668,In_610,In_666);
or U669 (N_669,In_79,In_426);
nand U670 (N_670,In_725,In_614);
and U671 (N_671,In_251,In_287);
nand U672 (N_672,In_552,In_371);
or U673 (N_673,In_234,In_608);
or U674 (N_674,In_646,In_687);
or U675 (N_675,In_518,In_10);
and U676 (N_676,In_28,In_18);
or U677 (N_677,In_54,In_494);
nand U678 (N_678,In_438,In_529);
or U679 (N_679,In_569,In_671);
nand U680 (N_680,In_178,In_22);
nand U681 (N_681,In_658,In_587);
and U682 (N_682,In_435,In_726);
and U683 (N_683,In_269,In_377);
and U684 (N_684,In_53,In_319);
nor U685 (N_685,In_460,In_355);
or U686 (N_686,In_232,In_326);
nor U687 (N_687,In_530,In_295);
or U688 (N_688,In_488,In_425);
nand U689 (N_689,In_490,In_744);
nor U690 (N_690,In_350,In_625);
nor U691 (N_691,In_114,In_232);
and U692 (N_692,In_613,In_506);
nor U693 (N_693,In_114,In_82);
or U694 (N_694,In_19,In_50);
nor U695 (N_695,In_581,In_474);
and U696 (N_696,In_207,In_103);
nand U697 (N_697,In_58,In_341);
or U698 (N_698,In_694,In_636);
nor U699 (N_699,In_35,In_411);
or U700 (N_700,In_58,In_562);
nor U701 (N_701,In_648,In_294);
or U702 (N_702,In_422,In_365);
nand U703 (N_703,In_2,In_190);
or U704 (N_704,In_572,In_254);
or U705 (N_705,In_284,In_440);
or U706 (N_706,In_123,In_143);
nor U707 (N_707,In_20,In_261);
or U708 (N_708,In_186,In_72);
nor U709 (N_709,In_23,In_460);
and U710 (N_710,In_39,In_190);
nor U711 (N_711,In_707,In_620);
or U712 (N_712,In_545,In_358);
xor U713 (N_713,In_624,In_505);
nor U714 (N_714,In_394,In_283);
and U715 (N_715,In_735,In_78);
nor U716 (N_716,In_446,In_40);
nor U717 (N_717,In_606,In_704);
nand U718 (N_718,In_222,In_62);
or U719 (N_719,In_659,In_494);
or U720 (N_720,In_181,In_655);
nor U721 (N_721,In_125,In_22);
and U722 (N_722,In_372,In_665);
nand U723 (N_723,In_267,In_386);
and U724 (N_724,In_245,In_517);
xor U725 (N_725,In_565,In_109);
and U726 (N_726,In_479,In_262);
nor U727 (N_727,In_443,In_744);
or U728 (N_728,In_517,In_364);
or U729 (N_729,In_588,In_507);
nand U730 (N_730,In_492,In_679);
nand U731 (N_731,In_607,In_579);
nand U732 (N_732,In_171,In_49);
nand U733 (N_733,In_701,In_636);
nand U734 (N_734,In_151,In_324);
and U735 (N_735,In_749,In_197);
nor U736 (N_736,In_278,In_365);
or U737 (N_737,In_119,In_25);
and U738 (N_738,In_60,In_139);
nand U739 (N_739,In_119,In_273);
nand U740 (N_740,In_271,In_98);
nor U741 (N_741,In_92,In_199);
and U742 (N_742,In_136,In_482);
nand U743 (N_743,In_524,In_440);
and U744 (N_744,In_21,In_696);
and U745 (N_745,In_691,In_243);
nor U746 (N_746,In_50,In_383);
or U747 (N_747,In_522,In_476);
or U748 (N_748,In_629,In_492);
nand U749 (N_749,In_171,In_518);
nor U750 (N_750,In_109,In_93);
nand U751 (N_751,In_543,In_421);
or U752 (N_752,In_411,In_49);
or U753 (N_753,In_551,In_587);
and U754 (N_754,In_3,In_663);
and U755 (N_755,In_110,In_638);
and U756 (N_756,In_587,In_271);
nand U757 (N_757,In_74,In_256);
nand U758 (N_758,In_415,In_602);
or U759 (N_759,In_17,In_612);
nand U760 (N_760,In_667,In_93);
and U761 (N_761,In_373,In_592);
nand U762 (N_762,In_576,In_47);
or U763 (N_763,In_604,In_458);
or U764 (N_764,In_721,In_710);
nor U765 (N_765,In_105,In_539);
nand U766 (N_766,In_432,In_437);
nand U767 (N_767,In_307,In_114);
or U768 (N_768,In_583,In_586);
nor U769 (N_769,In_65,In_351);
nand U770 (N_770,In_624,In_528);
and U771 (N_771,In_165,In_349);
and U772 (N_772,In_543,In_264);
nand U773 (N_773,In_352,In_600);
xnor U774 (N_774,In_602,In_684);
or U775 (N_775,In_290,In_604);
and U776 (N_776,In_579,In_222);
nor U777 (N_777,In_204,In_196);
and U778 (N_778,In_374,In_566);
xnor U779 (N_779,In_428,In_64);
nand U780 (N_780,In_122,In_420);
and U781 (N_781,In_81,In_122);
or U782 (N_782,In_122,In_221);
and U783 (N_783,In_41,In_476);
nand U784 (N_784,In_171,In_727);
nor U785 (N_785,In_726,In_14);
nand U786 (N_786,In_447,In_512);
and U787 (N_787,In_585,In_434);
or U788 (N_788,In_465,In_210);
nand U789 (N_789,In_186,In_350);
or U790 (N_790,In_522,In_701);
and U791 (N_791,In_447,In_733);
xnor U792 (N_792,In_554,In_428);
and U793 (N_793,In_93,In_114);
nor U794 (N_794,In_412,In_578);
nand U795 (N_795,In_457,In_275);
nor U796 (N_796,In_463,In_633);
or U797 (N_797,In_255,In_64);
nor U798 (N_798,In_522,In_445);
nor U799 (N_799,In_152,In_219);
nor U800 (N_800,In_590,In_200);
nand U801 (N_801,In_551,In_201);
and U802 (N_802,In_281,In_129);
nor U803 (N_803,In_16,In_535);
nand U804 (N_804,In_108,In_538);
nor U805 (N_805,In_211,In_229);
and U806 (N_806,In_250,In_747);
nand U807 (N_807,In_319,In_459);
xor U808 (N_808,In_586,In_620);
and U809 (N_809,In_707,In_725);
and U810 (N_810,In_539,In_178);
and U811 (N_811,In_710,In_706);
and U812 (N_812,In_202,In_206);
nor U813 (N_813,In_460,In_435);
nand U814 (N_814,In_167,In_666);
nand U815 (N_815,In_312,In_146);
nor U816 (N_816,In_189,In_374);
or U817 (N_817,In_426,In_609);
nor U818 (N_818,In_396,In_593);
nand U819 (N_819,In_397,In_416);
nor U820 (N_820,In_518,In_80);
and U821 (N_821,In_213,In_547);
nand U822 (N_822,In_100,In_332);
or U823 (N_823,In_638,In_601);
xnor U824 (N_824,In_397,In_619);
xnor U825 (N_825,In_169,In_476);
and U826 (N_826,In_544,In_566);
or U827 (N_827,In_642,In_288);
nor U828 (N_828,In_702,In_85);
and U829 (N_829,In_30,In_1);
nand U830 (N_830,In_42,In_600);
or U831 (N_831,In_260,In_676);
nand U832 (N_832,In_393,In_82);
and U833 (N_833,In_24,In_154);
or U834 (N_834,In_315,In_172);
and U835 (N_835,In_628,In_28);
nand U836 (N_836,In_209,In_442);
nand U837 (N_837,In_22,In_623);
and U838 (N_838,In_79,In_612);
nand U839 (N_839,In_290,In_449);
nand U840 (N_840,In_415,In_388);
nand U841 (N_841,In_135,In_229);
or U842 (N_842,In_81,In_467);
nand U843 (N_843,In_99,In_249);
or U844 (N_844,In_121,In_98);
or U845 (N_845,In_725,In_454);
nor U846 (N_846,In_643,In_388);
or U847 (N_847,In_662,In_263);
and U848 (N_848,In_162,In_231);
or U849 (N_849,In_242,In_103);
or U850 (N_850,In_646,In_338);
and U851 (N_851,In_11,In_2);
or U852 (N_852,In_194,In_674);
and U853 (N_853,In_33,In_671);
or U854 (N_854,In_45,In_573);
nor U855 (N_855,In_380,In_722);
nor U856 (N_856,In_689,In_192);
or U857 (N_857,In_501,In_252);
nand U858 (N_858,In_329,In_652);
and U859 (N_859,In_326,In_393);
or U860 (N_860,In_305,In_346);
and U861 (N_861,In_269,In_340);
nand U862 (N_862,In_380,In_694);
nor U863 (N_863,In_245,In_59);
nor U864 (N_864,In_516,In_385);
or U865 (N_865,In_333,In_361);
and U866 (N_866,In_317,In_726);
nand U867 (N_867,In_59,In_4);
nand U868 (N_868,In_416,In_151);
nor U869 (N_869,In_700,In_143);
nor U870 (N_870,In_617,In_620);
and U871 (N_871,In_31,In_322);
nand U872 (N_872,In_326,In_311);
or U873 (N_873,In_545,In_389);
nor U874 (N_874,In_307,In_692);
nor U875 (N_875,In_645,In_226);
nor U876 (N_876,In_277,In_291);
nor U877 (N_877,In_558,In_352);
or U878 (N_878,In_660,In_506);
and U879 (N_879,In_678,In_151);
nor U880 (N_880,In_661,In_104);
nand U881 (N_881,In_345,In_740);
and U882 (N_882,In_316,In_256);
nor U883 (N_883,In_531,In_640);
nand U884 (N_884,In_328,In_545);
or U885 (N_885,In_381,In_67);
nor U886 (N_886,In_230,In_745);
nor U887 (N_887,In_281,In_347);
and U888 (N_888,In_529,In_610);
nand U889 (N_889,In_701,In_247);
nor U890 (N_890,In_640,In_493);
nor U891 (N_891,In_398,In_748);
or U892 (N_892,In_391,In_548);
or U893 (N_893,In_681,In_453);
nor U894 (N_894,In_430,In_711);
nand U895 (N_895,In_564,In_578);
or U896 (N_896,In_194,In_336);
and U897 (N_897,In_686,In_202);
and U898 (N_898,In_479,In_310);
or U899 (N_899,In_745,In_484);
and U900 (N_900,In_184,In_405);
nor U901 (N_901,In_442,In_572);
nand U902 (N_902,In_49,In_679);
nor U903 (N_903,In_11,In_73);
nand U904 (N_904,In_450,In_494);
and U905 (N_905,In_548,In_93);
or U906 (N_906,In_16,In_304);
and U907 (N_907,In_194,In_264);
nand U908 (N_908,In_456,In_723);
nand U909 (N_909,In_688,In_713);
or U910 (N_910,In_656,In_294);
nand U911 (N_911,In_236,In_61);
nor U912 (N_912,In_374,In_468);
nand U913 (N_913,In_156,In_561);
and U914 (N_914,In_208,In_382);
nand U915 (N_915,In_629,In_657);
nor U916 (N_916,In_138,In_430);
and U917 (N_917,In_431,In_653);
nand U918 (N_918,In_311,In_657);
and U919 (N_919,In_209,In_565);
or U920 (N_920,In_247,In_476);
nor U921 (N_921,In_726,In_704);
nand U922 (N_922,In_394,In_351);
nand U923 (N_923,In_114,In_273);
nor U924 (N_924,In_317,In_480);
nor U925 (N_925,In_251,In_246);
xnor U926 (N_926,In_233,In_356);
and U927 (N_927,In_676,In_278);
or U928 (N_928,In_167,In_735);
nor U929 (N_929,In_133,In_685);
and U930 (N_930,In_304,In_150);
or U931 (N_931,In_244,In_691);
nand U932 (N_932,In_648,In_297);
xor U933 (N_933,In_427,In_428);
nand U934 (N_934,In_66,In_207);
or U935 (N_935,In_408,In_418);
and U936 (N_936,In_405,In_23);
nor U937 (N_937,In_67,In_478);
or U938 (N_938,In_166,In_285);
and U939 (N_939,In_432,In_146);
nand U940 (N_940,In_123,In_102);
and U941 (N_941,In_552,In_217);
nand U942 (N_942,In_573,In_348);
nand U943 (N_943,In_49,In_354);
or U944 (N_944,In_607,In_517);
or U945 (N_945,In_5,In_428);
or U946 (N_946,In_140,In_47);
or U947 (N_947,In_643,In_180);
nor U948 (N_948,In_83,In_430);
and U949 (N_949,In_417,In_10);
and U950 (N_950,In_308,In_454);
or U951 (N_951,In_25,In_392);
and U952 (N_952,In_587,In_584);
nor U953 (N_953,In_86,In_240);
and U954 (N_954,In_119,In_615);
or U955 (N_955,In_490,In_472);
nor U956 (N_956,In_235,In_109);
or U957 (N_957,In_118,In_562);
nand U958 (N_958,In_361,In_18);
and U959 (N_959,In_312,In_27);
and U960 (N_960,In_168,In_658);
and U961 (N_961,In_474,In_571);
and U962 (N_962,In_619,In_375);
and U963 (N_963,In_107,In_621);
or U964 (N_964,In_739,In_370);
nand U965 (N_965,In_127,In_156);
nor U966 (N_966,In_215,In_695);
nor U967 (N_967,In_400,In_120);
nand U968 (N_968,In_631,In_46);
or U969 (N_969,In_308,In_583);
nand U970 (N_970,In_724,In_331);
nor U971 (N_971,In_365,In_697);
or U972 (N_972,In_300,In_77);
nand U973 (N_973,In_238,In_603);
or U974 (N_974,In_705,In_493);
and U975 (N_975,In_41,In_22);
nand U976 (N_976,In_347,In_328);
nor U977 (N_977,In_372,In_145);
nand U978 (N_978,In_528,In_244);
and U979 (N_979,In_279,In_657);
nor U980 (N_980,In_77,In_244);
or U981 (N_981,In_319,In_710);
or U982 (N_982,In_83,In_468);
and U983 (N_983,In_660,In_477);
nor U984 (N_984,In_299,In_83);
and U985 (N_985,In_596,In_364);
and U986 (N_986,In_449,In_341);
nor U987 (N_987,In_276,In_726);
nor U988 (N_988,In_271,In_27);
nor U989 (N_989,In_329,In_567);
or U990 (N_990,In_8,In_142);
nor U991 (N_991,In_692,In_470);
or U992 (N_992,In_508,In_446);
or U993 (N_993,In_500,In_136);
nor U994 (N_994,In_386,In_530);
nand U995 (N_995,In_1,In_228);
and U996 (N_996,In_565,In_517);
and U997 (N_997,In_126,In_51);
and U998 (N_998,In_728,In_738);
and U999 (N_999,In_257,In_292);
and U1000 (N_1000,N_246,N_423);
nor U1001 (N_1001,N_128,N_85);
or U1002 (N_1002,N_655,N_244);
or U1003 (N_1003,N_776,N_406);
or U1004 (N_1004,N_898,N_508);
and U1005 (N_1005,N_855,N_391);
xor U1006 (N_1006,N_999,N_226);
or U1007 (N_1007,N_453,N_537);
nand U1008 (N_1008,N_117,N_507);
nor U1009 (N_1009,N_615,N_430);
or U1010 (N_1010,N_256,N_198);
and U1011 (N_1011,N_635,N_730);
and U1012 (N_1012,N_355,N_70);
or U1013 (N_1013,N_264,N_853);
nand U1014 (N_1014,N_598,N_161);
and U1015 (N_1015,N_762,N_57);
nor U1016 (N_1016,N_27,N_720);
nor U1017 (N_1017,N_540,N_463);
or U1018 (N_1018,N_620,N_62);
or U1019 (N_1019,N_634,N_392);
nor U1020 (N_1020,N_409,N_407);
nand U1021 (N_1021,N_848,N_412);
or U1022 (N_1022,N_528,N_433);
or U1023 (N_1023,N_492,N_530);
xnor U1024 (N_1024,N_954,N_243);
and U1025 (N_1025,N_488,N_214);
nor U1026 (N_1026,N_34,N_60);
nor U1027 (N_1027,N_516,N_440);
and U1028 (N_1028,N_472,N_342);
and U1029 (N_1029,N_520,N_344);
nand U1030 (N_1030,N_926,N_651);
nor U1031 (N_1031,N_144,N_394);
nor U1032 (N_1032,N_638,N_676);
nor U1033 (N_1033,N_712,N_928);
nand U1034 (N_1034,N_580,N_308);
nand U1035 (N_1035,N_663,N_19);
nand U1036 (N_1036,N_944,N_22);
nand U1037 (N_1037,N_704,N_485);
nor U1038 (N_1038,N_556,N_671);
or U1039 (N_1039,N_672,N_310);
or U1040 (N_1040,N_827,N_583);
or U1041 (N_1041,N_187,N_319);
nand U1042 (N_1042,N_260,N_825);
or U1043 (N_1043,N_362,N_466);
nor U1044 (N_1044,N_545,N_765);
nand U1045 (N_1045,N_31,N_670);
nand U1046 (N_1046,N_872,N_821);
and U1047 (N_1047,N_114,N_504);
nor U1048 (N_1048,N_986,N_330);
or U1049 (N_1049,N_212,N_905);
nand U1050 (N_1050,N_102,N_633);
nand U1051 (N_1051,N_305,N_118);
nand U1052 (N_1052,N_541,N_293);
xnor U1053 (N_1053,N_259,N_797);
or U1054 (N_1054,N_434,N_796);
nor U1055 (N_1055,N_242,N_735);
nor U1056 (N_1056,N_913,N_549);
and U1057 (N_1057,N_405,N_594);
or U1058 (N_1058,N_511,N_533);
nand U1059 (N_1059,N_744,N_6);
and U1060 (N_1060,N_439,N_650);
or U1061 (N_1061,N_452,N_250);
and U1062 (N_1062,N_331,N_457);
nand U1063 (N_1063,N_172,N_194);
xor U1064 (N_1064,N_982,N_639);
and U1065 (N_1065,N_678,N_625);
nor U1066 (N_1066,N_358,N_177);
and U1067 (N_1067,N_658,N_205);
or U1068 (N_1068,N_654,N_980);
nor U1069 (N_1069,N_686,N_660);
nor U1070 (N_1070,N_858,N_952);
or U1071 (N_1071,N_554,N_182);
nand U1072 (N_1072,N_421,N_737);
or U1073 (N_1073,N_499,N_691);
nand U1074 (N_1074,N_725,N_352);
and U1075 (N_1075,N_469,N_422);
nor U1076 (N_1076,N_224,N_346);
nand U1077 (N_1077,N_402,N_397);
or U1078 (N_1078,N_763,N_360);
nand U1079 (N_1079,N_673,N_496);
nor U1080 (N_1080,N_335,N_839);
or U1081 (N_1081,N_950,N_122);
and U1082 (N_1082,N_637,N_404);
and U1083 (N_1083,N_602,N_771);
and U1084 (N_1084,N_486,N_150);
and U1085 (N_1085,N_241,N_699);
nor U1086 (N_1086,N_661,N_413);
or U1087 (N_1087,N_851,N_290);
or U1088 (N_1088,N_875,N_896);
nand U1089 (N_1089,N_399,N_687);
nor U1090 (N_1090,N_774,N_832);
and U1091 (N_1091,N_199,N_201);
nor U1092 (N_1092,N_403,N_436);
nor U1093 (N_1093,N_990,N_417);
or U1094 (N_1094,N_757,N_36);
or U1095 (N_1095,N_566,N_525);
nand U1096 (N_1096,N_804,N_273);
and U1097 (N_1097,N_18,N_746);
or U1098 (N_1098,N_121,N_674);
nor U1099 (N_1099,N_960,N_828);
and U1100 (N_1100,N_315,N_572);
and U1101 (N_1101,N_592,N_595);
nand U1102 (N_1102,N_79,N_279);
nor U1103 (N_1103,N_14,N_450);
or U1104 (N_1104,N_265,N_612);
nor U1105 (N_1105,N_175,N_39);
xor U1106 (N_1106,N_603,N_419);
nand U1107 (N_1107,N_732,N_274);
and U1108 (N_1108,N_788,N_963);
nor U1109 (N_1109,N_679,N_321);
nor U1110 (N_1110,N_123,N_956);
nand U1111 (N_1111,N_316,N_747);
and U1112 (N_1112,N_333,N_569);
and U1113 (N_1113,N_743,N_465);
or U1114 (N_1114,N_48,N_613);
and U1115 (N_1115,N_824,N_716);
nand U1116 (N_1116,N_728,N_325);
and U1117 (N_1117,N_695,N_131);
nand U1118 (N_1118,N_561,N_113);
nand U1119 (N_1119,N_411,N_285);
nor U1120 (N_1120,N_912,N_476);
nand U1121 (N_1121,N_631,N_281);
or U1122 (N_1122,N_366,N_13);
nand U1123 (N_1123,N_854,N_234);
or U1124 (N_1124,N_731,N_745);
nor U1125 (N_1125,N_455,N_587);
or U1126 (N_1126,N_862,N_334);
or U1127 (N_1127,N_618,N_213);
and U1128 (N_1128,N_675,N_899);
nor U1129 (N_1129,N_599,N_664);
nand U1130 (N_1130,N_207,N_245);
and U1131 (N_1131,N_130,N_152);
nand U1132 (N_1132,N_420,N_965);
nor U1133 (N_1133,N_864,N_221);
nand U1134 (N_1134,N_662,N_966);
nor U1135 (N_1135,N_361,N_880);
or U1136 (N_1136,N_877,N_665);
or U1137 (N_1137,N_647,N_840);
and U1138 (N_1138,N_90,N_992);
nand U1139 (N_1139,N_483,N_159);
and U1140 (N_1140,N_61,N_365);
and U1141 (N_1141,N_685,N_987);
and U1142 (N_1142,N_425,N_581);
nor U1143 (N_1143,N_138,N_734);
and U1144 (N_1144,N_69,N_444);
nor U1145 (N_1145,N_43,N_805);
nand U1146 (N_1146,N_560,N_641);
or U1147 (N_1147,N_148,N_220);
or U1148 (N_1148,N_773,N_823);
nand U1149 (N_1149,N_309,N_286);
nand U1150 (N_1150,N_521,N_21);
or U1151 (N_1151,N_793,N_844);
nand U1152 (N_1152,N_544,N_99);
nor U1153 (N_1153,N_188,N_870);
and U1154 (N_1154,N_555,N_733);
nor U1155 (N_1155,N_291,N_523);
nor U1156 (N_1156,N_971,N_551);
or U1157 (N_1157,N_814,N_863);
nor U1158 (N_1158,N_389,N_761);
nand U1159 (N_1159,N_922,N_866);
or U1160 (N_1160,N_856,N_363);
and U1161 (N_1161,N_408,N_74);
nand U1162 (N_1162,N_697,N_101);
nor U1163 (N_1163,N_652,N_106);
nand U1164 (N_1164,N_77,N_609);
or U1165 (N_1165,N_681,N_626);
or U1166 (N_1166,N_881,N_775);
or U1167 (N_1167,N_559,N_54);
xnor U1168 (N_1168,N_147,N_103);
or U1169 (N_1169,N_183,N_885);
nor U1170 (N_1170,N_842,N_482);
and U1171 (N_1171,N_341,N_715);
nor U1172 (N_1172,N_888,N_228);
nand U1173 (N_1173,N_480,N_63);
and U1174 (N_1174,N_962,N_170);
and U1175 (N_1175,N_98,N_158);
or U1176 (N_1176,N_445,N_15);
nand U1177 (N_1177,N_340,N_543);
nor U1178 (N_1178,N_314,N_958);
nor U1179 (N_1179,N_865,N_656);
nor U1180 (N_1180,N_126,N_738);
and U1181 (N_1181,N_822,N_235);
or U1182 (N_1182,N_81,N_969);
nor U1183 (N_1183,N_336,N_993);
or U1184 (N_1184,N_88,N_169);
nand U1185 (N_1185,N_184,N_818);
or U1186 (N_1186,N_945,N_350);
nor U1187 (N_1187,N_49,N_813);
nand U1188 (N_1188,N_367,N_616);
nor U1189 (N_1189,N_550,N_902);
nand U1190 (N_1190,N_186,N_448);
nand U1191 (N_1191,N_710,N_299);
nor U1192 (N_1192,N_884,N_381);
nor U1193 (N_1193,N_754,N_109);
and U1194 (N_1194,N_531,N_949);
nand U1195 (N_1195,N_32,N_203);
or U1196 (N_1196,N_611,N_921);
or U1197 (N_1197,N_302,N_23);
nand U1198 (N_1198,N_933,N_134);
nor U1199 (N_1199,N_727,N_629);
nand U1200 (N_1200,N_906,N_370);
nor U1201 (N_1201,N_558,N_957);
and U1202 (N_1202,N_972,N_11);
xnor U1203 (N_1203,N_92,N_240);
and U1204 (N_1204,N_160,N_740);
nand U1205 (N_1205,N_810,N_816);
or U1206 (N_1206,N_619,N_964);
and U1207 (N_1207,N_239,N_939);
and U1208 (N_1208,N_287,N_108);
nor U1209 (N_1209,N_791,N_717);
nand U1210 (N_1210,N_565,N_874);
or U1211 (N_1211,N_783,N_12);
and U1212 (N_1212,N_850,N_137);
or U1213 (N_1213,N_838,N_871);
or U1214 (N_1214,N_522,N_597);
or U1215 (N_1215,N_383,N_371);
nor U1216 (N_1216,N_223,N_538);
nor U1217 (N_1217,N_50,N_171);
and U1218 (N_1218,N_772,N_56);
and U1219 (N_1219,N_111,N_86);
nand U1220 (N_1220,N_849,N_846);
nor U1221 (N_1221,N_973,N_192);
and U1222 (N_1222,N_571,N_802);
xnor U1223 (N_1223,N_459,N_836);
nand U1224 (N_1224,N_104,N_512);
and U1225 (N_1225,N_454,N_696);
or U1226 (N_1226,N_28,N_364);
or U1227 (N_1227,N_276,N_238);
nor U1228 (N_1228,N_369,N_372);
and U1229 (N_1229,N_494,N_644);
or U1230 (N_1230,N_280,N_173);
or U1231 (N_1231,N_792,N_518);
and U1232 (N_1232,N_298,N_932);
and U1233 (N_1233,N_296,N_557);
or U1234 (N_1234,N_384,N_534);
nor U1235 (N_1235,N_112,N_261);
nand U1236 (N_1236,N_831,N_924);
or U1237 (N_1237,N_536,N_105);
and U1238 (N_1238,N_795,N_861);
nand U1239 (N_1239,N_3,N_843);
and U1240 (N_1240,N_711,N_984);
and U1241 (N_1241,N_708,N_784);
xnor U1242 (N_1242,N_432,N_329);
nand U1243 (N_1243,N_236,N_202);
nor U1244 (N_1244,N_567,N_812);
nor U1245 (N_1245,N_232,N_251);
and U1246 (N_1246,N_596,N_777);
nor U1247 (N_1247,N_785,N_501);
and U1248 (N_1248,N_584,N_903);
and U1249 (N_1249,N_217,N_778);
or U1250 (N_1250,N_263,N_841);
nand U1251 (N_1251,N_200,N_829);
nand U1252 (N_1252,N_67,N_487);
and U1253 (N_1253,N_312,N_72);
xnor U1254 (N_1254,N_506,N_484);
or U1255 (N_1255,N_124,N_968);
nand U1256 (N_1256,N_497,N_573);
and U1257 (N_1257,N_955,N_689);
nand U1258 (N_1258,N_272,N_490);
nor U1259 (N_1259,N_868,N_229);
nand U1260 (N_1260,N_2,N_890);
or U1261 (N_1261,N_996,N_210);
xnor U1262 (N_1262,N_677,N_624);
nor U1263 (N_1263,N_395,N_377);
nand U1264 (N_1264,N_800,N_789);
or U1265 (N_1265,N_292,N_943);
xnor U1266 (N_1266,N_517,N_166);
nor U1267 (N_1267,N_748,N_713);
nand U1268 (N_1268,N_750,N_378);
nor U1269 (N_1269,N_542,N_847);
or U1270 (N_1270,N_925,N_353);
nor U1271 (N_1271,N_266,N_967);
nor U1272 (N_1272,N_979,N_191);
nand U1273 (N_1273,N_337,N_535);
or U1274 (N_1274,N_931,N_119);
nand U1275 (N_1275,N_895,N_857);
nand U1276 (N_1276,N_278,N_723);
nand U1277 (N_1277,N_458,N_424);
and U1278 (N_1278,N_593,N_219);
or U1279 (N_1279,N_41,N_129);
nor U1280 (N_1280,N_927,N_891);
and U1281 (N_1281,N_961,N_782);
and U1282 (N_1282,N_837,N_657);
nand U1283 (N_1283,N_684,N_869);
nand U1284 (N_1284,N_268,N_151);
or U1285 (N_1285,N_703,N_87);
nor U1286 (N_1286,N_375,N_338);
and U1287 (N_1287,N_820,N_948);
xor U1288 (N_1288,N_909,N_649);
xor U1289 (N_1289,N_718,N_461);
nand U1290 (N_1290,N_576,N_179);
nand U1291 (N_1291,N_97,N_288);
or U1292 (N_1292,N_254,N_387);
nand U1293 (N_1293,N_892,N_82);
and U1294 (N_1294,N_887,N_59);
nor U1295 (N_1295,N_653,N_93);
or U1296 (N_1296,N_47,N_883);
nand U1297 (N_1297,N_33,N_359);
nor U1298 (N_1298,N_867,N_323);
nor U1299 (N_1299,N_798,N_271);
and U1300 (N_1300,N_766,N_78);
nor U1301 (N_1301,N_357,N_30);
or U1302 (N_1302,N_218,N_683);
nor U1303 (N_1303,N_894,N_908);
and U1304 (N_1304,N_35,N_132);
nand U1305 (N_1305,N_449,N_468);
nor U1306 (N_1306,N_590,N_705);
nand U1307 (N_1307,N_267,N_206);
and U1308 (N_1308,N_473,N_456);
xnor U1309 (N_1309,N_435,N_324);
nand U1310 (N_1310,N_991,N_736);
or U1311 (N_1311,N_859,N_493);
xnor U1312 (N_1312,N_978,N_115);
and U1313 (N_1313,N_441,N_724);
and U1314 (N_1314,N_349,N_601);
and U1315 (N_1315,N_694,N_89);
nor U1316 (N_1316,N_668,N_167);
and U1317 (N_1317,N_415,N_416);
nor U1318 (N_1318,N_91,N_873);
nor U1319 (N_1319,N_320,N_510);
and U1320 (N_1320,N_742,N_429);
nand U1321 (N_1321,N_768,N_769);
nand U1322 (N_1322,N_692,N_505);
and U1323 (N_1323,N_38,N_513);
and U1324 (N_1324,N_693,N_632);
and U1325 (N_1325,N_10,N_636);
or U1326 (N_1326,N_879,N_646);
nor U1327 (N_1327,N_749,N_42);
nor U1328 (N_1328,N_889,N_446);
nand U1329 (N_1329,N_110,N_878);
nand U1330 (N_1330,N_1,N_529);
nor U1331 (N_1331,N_781,N_168);
nor U1332 (N_1332,N_174,N_640);
nand U1333 (N_1333,N_706,N_20);
nand U1334 (N_1334,N_589,N_503);
nand U1335 (N_1335,N_339,N_295);
nor U1336 (N_1336,N_382,N_294);
or U1337 (N_1337,N_139,N_356);
or U1338 (N_1338,N_477,N_585);
nor U1339 (N_1339,N_193,N_519);
nand U1340 (N_1340,N_751,N_208);
nor U1341 (N_1341,N_71,N_227);
or U1342 (N_1342,N_489,N_709);
nor U1343 (N_1343,N_438,N_153);
nand U1344 (N_1344,N_630,N_396);
or U1345 (N_1345,N_666,N_915);
xor U1346 (N_1346,N_714,N_24);
nand U1347 (N_1347,N_907,N_68);
nand U1348 (N_1348,N_17,N_373);
nor U1349 (N_1349,N_989,N_526);
xor U1350 (N_1350,N_547,N_269);
and U1351 (N_1351,N_195,N_176);
nand U1352 (N_1352,N_920,N_4);
and U1353 (N_1353,N_985,N_918);
and U1354 (N_1354,N_995,N_591);
nand U1355 (N_1355,N_946,N_46);
or U1356 (N_1356,N_600,N_189);
xor U1357 (N_1357,N_418,N_552);
and U1358 (N_1358,N_579,N_690);
nand U1359 (N_1359,N_318,N_940);
nor U1360 (N_1360,N_313,N_947);
nand U1361 (N_1361,N_351,N_233);
nand U1362 (N_1362,N_532,N_45);
and U1363 (N_1363,N_911,N_648);
or U1364 (N_1364,N_155,N_474);
nor U1365 (N_1365,N_426,N_451);
and U1366 (N_1366,N_852,N_688);
nand U1367 (N_1367,N_142,N_794);
nand U1368 (N_1368,N_211,N_760);
nand U1369 (N_1369,N_916,N_919);
xor U1370 (N_1370,N_860,N_431);
and U1371 (N_1371,N_178,N_209);
nand U1372 (N_1372,N_51,N_467);
nand U1373 (N_1373,N_64,N_133);
nor U1374 (N_1374,N_143,N_475);
nor U1375 (N_1375,N_617,N_0);
or U1376 (N_1376,N_698,N_524);
nand U1377 (N_1377,N_937,N_498);
or U1378 (N_1378,N_442,N_154);
nand U1379 (N_1379,N_196,N_669);
nor U1380 (N_1380,N_317,N_819);
nand U1381 (N_1381,N_759,N_876);
nor U1382 (N_1382,N_258,N_328);
and U1383 (N_1383,N_970,N_185);
and U1384 (N_1384,N_343,N_808);
and U1385 (N_1385,N_398,N_502);
nand U1386 (N_1386,N_753,N_462);
or U1387 (N_1387,N_807,N_180);
nor U1388 (N_1388,N_247,N_300);
or U1389 (N_1389,N_306,N_826);
nor U1390 (N_1390,N_479,N_135);
nand U1391 (N_1391,N_301,N_741);
nor U1392 (N_1392,N_53,N_307);
nand U1393 (N_1393,N_929,N_7);
nor U1394 (N_1394,N_9,N_553);
and U1395 (N_1395,N_156,N_707);
or U1396 (N_1396,N_495,N_146);
and U1397 (N_1397,N_275,N_739);
or U1398 (N_1398,N_73,N_815);
nand U1399 (N_1399,N_835,N_368);
nor U1400 (N_1400,N_29,N_8);
xnor U1401 (N_1401,N_787,N_722);
or U1402 (N_1402,N_354,N_181);
nor U1403 (N_1403,N_562,N_780);
and U1404 (N_1404,N_622,N_437);
or U1405 (N_1405,N_515,N_447);
nand U1406 (N_1406,N_95,N_262);
nor U1407 (N_1407,N_882,N_910);
or U1408 (N_1408,N_44,N_975);
or U1409 (N_1409,N_701,N_120);
nand U1410 (N_1410,N_248,N_577);
nand U1411 (N_1411,N_570,N_470);
nor U1412 (N_1412,N_141,N_627);
and U1413 (N_1413,N_659,N_26);
nand U1414 (N_1414,N_427,N_164);
nor U1415 (N_1415,N_374,N_162);
or U1416 (N_1416,N_610,N_500);
nand U1417 (N_1417,N_755,N_886);
and U1418 (N_1418,N_282,N_326);
and U1419 (N_1419,N_941,N_222);
and U1420 (N_1420,N_230,N_255);
nand U1421 (N_1421,N_586,N_322);
nor U1422 (N_1422,N_237,N_817);
nor U1423 (N_1423,N_700,N_327);
or U1424 (N_1424,N_252,N_983);
or U1425 (N_1425,N_388,N_994);
and U1426 (N_1426,N_758,N_803);
nand U1427 (N_1427,N_702,N_464);
or U1428 (N_1428,N_284,N_893);
nand U1429 (N_1429,N_953,N_231);
and U1430 (N_1430,N_645,N_767);
nor U1431 (N_1431,N_951,N_348);
nor U1432 (N_1432,N_605,N_478);
or U1433 (N_1433,N_136,N_347);
or U1434 (N_1434,N_998,N_80);
and U1435 (N_1435,N_834,N_410);
or U1436 (N_1436,N_215,N_157);
or U1437 (N_1437,N_786,N_604);
nand U1438 (N_1438,N_623,N_52);
and U1439 (N_1439,N_277,N_667);
or U1440 (N_1440,N_303,N_390);
and U1441 (N_1441,N_311,N_682);
nor U1442 (N_1442,N_997,N_116);
nand U1443 (N_1443,N_165,N_582);
and U1444 (N_1444,N_935,N_400);
nor U1445 (N_1445,N_332,N_801);
nor U1446 (N_1446,N_901,N_934);
nor U1447 (N_1447,N_756,N_83);
nand U1448 (N_1448,N_642,N_16);
nand U1449 (N_1449,N_471,N_5);
xnor U1450 (N_1450,N_25,N_65);
nand U1451 (N_1451,N_270,N_614);
and U1452 (N_1452,N_140,N_621);
nand U1453 (N_1453,N_345,N_799);
nand U1454 (N_1454,N_607,N_574);
nand U1455 (N_1455,N_564,N_546);
nand U1456 (N_1456,N_900,N_833);
nand U1457 (N_1457,N_930,N_379);
nor U1458 (N_1458,N_790,N_40);
nand U1459 (N_1459,N_145,N_988);
nor U1460 (N_1460,N_401,N_385);
nor U1461 (N_1461,N_163,N_514);
and U1462 (N_1462,N_58,N_414);
and U1463 (N_1463,N_289,N_225);
nand U1464 (N_1464,N_460,N_197);
and U1465 (N_1465,N_37,N_914);
nor U1466 (N_1466,N_539,N_393);
nor U1467 (N_1467,N_845,N_923);
xor U1468 (N_1468,N_107,N_376);
or U1469 (N_1469,N_304,N_897);
nor U1470 (N_1470,N_568,N_55);
and U1471 (N_1471,N_643,N_976);
nand U1472 (N_1472,N_149,N_719);
and U1473 (N_1473,N_588,N_386);
or U1474 (N_1474,N_100,N_628);
and U1475 (N_1475,N_606,N_66);
or U1476 (N_1476,N_125,N_481);
or U1477 (N_1477,N_938,N_578);
nor U1478 (N_1478,N_936,N_726);
nor U1479 (N_1479,N_917,N_811);
nand U1480 (N_1480,N_84,N_548);
nor U1481 (N_1481,N_216,N_257);
and U1482 (N_1482,N_721,N_729);
and U1483 (N_1483,N_563,N_76);
or U1484 (N_1484,N_443,N_491);
nand U1485 (N_1485,N_959,N_608);
or U1486 (N_1486,N_283,N_830);
xnor U1487 (N_1487,N_527,N_809);
nand U1488 (N_1488,N_770,N_253);
or U1489 (N_1489,N_806,N_249);
or U1490 (N_1490,N_96,N_127);
nor U1491 (N_1491,N_904,N_680);
or U1492 (N_1492,N_575,N_297);
or U1493 (N_1493,N_75,N_981);
nor U1494 (N_1494,N_94,N_974);
nand U1495 (N_1495,N_942,N_204);
and U1496 (N_1496,N_752,N_509);
nor U1497 (N_1497,N_428,N_764);
nor U1498 (N_1498,N_779,N_977);
and U1499 (N_1499,N_380,N_190);
nor U1500 (N_1500,N_734,N_812);
nor U1501 (N_1501,N_407,N_397);
nor U1502 (N_1502,N_951,N_550);
and U1503 (N_1503,N_530,N_756);
nor U1504 (N_1504,N_651,N_223);
and U1505 (N_1505,N_878,N_139);
and U1506 (N_1506,N_313,N_750);
nand U1507 (N_1507,N_223,N_404);
nor U1508 (N_1508,N_698,N_116);
and U1509 (N_1509,N_567,N_828);
nor U1510 (N_1510,N_234,N_326);
nand U1511 (N_1511,N_773,N_887);
xnor U1512 (N_1512,N_317,N_720);
nor U1513 (N_1513,N_885,N_312);
nand U1514 (N_1514,N_163,N_360);
nand U1515 (N_1515,N_373,N_684);
nand U1516 (N_1516,N_199,N_740);
xnor U1517 (N_1517,N_849,N_24);
nand U1518 (N_1518,N_58,N_606);
nor U1519 (N_1519,N_386,N_873);
nand U1520 (N_1520,N_647,N_462);
nor U1521 (N_1521,N_820,N_199);
nor U1522 (N_1522,N_5,N_186);
or U1523 (N_1523,N_832,N_942);
nor U1524 (N_1524,N_747,N_911);
and U1525 (N_1525,N_676,N_484);
nor U1526 (N_1526,N_613,N_815);
or U1527 (N_1527,N_15,N_282);
and U1528 (N_1528,N_621,N_832);
or U1529 (N_1529,N_623,N_72);
nor U1530 (N_1530,N_605,N_501);
nor U1531 (N_1531,N_321,N_778);
nand U1532 (N_1532,N_953,N_719);
nand U1533 (N_1533,N_930,N_662);
and U1534 (N_1534,N_954,N_8);
nand U1535 (N_1535,N_501,N_540);
nor U1536 (N_1536,N_804,N_599);
nor U1537 (N_1537,N_279,N_947);
xnor U1538 (N_1538,N_255,N_843);
nor U1539 (N_1539,N_91,N_437);
nand U1540 (N_1540,N_877,N_469);
or U1541 (N_1541,N_536,N_277);
or U1542 (N_1542,N_958,N_225);
and U1543 (N_1543,N_570,N_307);
xnor U1544 (N_1544,N_632,N_102);
nor U1545 (N_1545,N_239,N_654);
or U1546 (N_1546,N_590,N_401);
nor U1547 (N_1547,N_407,N_799);
or U1548 (N_1548,N_521,N_634);
xor U1549 (N_1549,N_845,N_17);
and U1550 (N_1550,N_139,N_240);
and U1551 (N_1551,N_253,N_749);
and U1552 (N_1552,N_240,N_744);
or U1553 (N_1553,N_169,N_527);
or U1554 (N_1554,N_129,N_653);
nor U1555 (N_1555,N_950,N_275);
or U1556 (N_1556,N_810,N_949);
nor U1557 (N_1557,N_505,N_948);
nor U1558 (N_1558,N_302,N_464);
or U1559 (N_1559,N_16,N_259);
and U1560 (N_1560,N_701,N_806);
nand U1561 (N_1561,N_973,N_464);
or U1562 (N_1562,N_12,N_553);
or U1563 (N_1563,N_266,N_955);
or U1564 (N_1564,N_48,N_418);
or U1565 (N_1565,N_439,N_635);
and U1566 (N_1566,N_940,N_562);
nor U1567 (N_1567,N_970,N_774);
and U1568 (N_1568,N_484,N_164);
and U1569 (N_1569,N_626,N_995);
and U1570 (N_1570,N_134,N_351);
nor U1571 (N_1571,N_404,N_782);
nand U1572 (N_1572,N_2,N_409);
or U1573 (N_1573,N_813,N_128);
nor U1574 (N_1574,N_282,N_415);
or U1575 (N_1575,N_54,N_422);
and U1576 (N_1576,N_209,N_918);
nor U1577 (N_1577,N_773,N_189);
nor U1578 (N_1578,N_851,N_159);
nand U1579 (N_1579,N_142,N_136);
nand U1580 (N_1580,N_385,N_973);
or U1581 (N_1581,N_10,N_553);
nand U1582 (N_1582,N_891,N_705);
nand U1583 (N_1583,N_752,N_453);
or U1584 (N_1584,N_287,N_385);
and U1585 (N_1585,N_941,N_436);
and U1586 (N_1586,N_665,N_822);
nand U1587 (N_1587,N_702,N_916);
or U1588 (N_1588,N_506,N_463);
and U1589 (N_1589,N_638,N_164);
nor U1590 (N_1590,N_771,N_511);
or U1591 (N_1591,N_339,N_16);
nand U1592 (N_1592,N_296,N_593);
or U1593 (N_1593,N_846,N_52);
or U1594 (N_1594,N_45,N_4);
nor U1595 (N_1595,N_745,N_806);
and U1596 (N_1596,N_168,N_441);
nand U1597 (N_1597,N_883,N_12);
and U1598 (N_1598,N_257,N_558);
nor U1599 (N_1599,N_112,N_958);
nand U1600 (N_1600,N_913,N_171);
and U1601 (N_1601,N_279,N_493);
nand U1602 (N_1602,N_417,N_718);
nand U1603 (N_1603,N_678,N_250);
or U1604 (N_1604,N_863,N_234);
nor U1605 (N_1605,N_453,N_507);
or U1606 (N_1606,N_291,N_381);
or U1607 (N_1607,N_652,N_635);
nor U1608 (N_1608,N_570,N_818);
and U1609 (N_1609,N_381,N_196);
nor U1610 (N_1610,N_102,N_508);
nand U1611 (N_1611,N_458,N_671);
xnor U1612 (N_1612,N_445,N_737);
or U1613 (N_1613,N_961,N_395);
nor U1614 (N_1614,N_649,N_598);
and U1615 (N_1615,N_359,N_604);
or U1616 (N_1616,N_218,N_74);
or U1617 (N_1617,N_283,N_176);
nor U1618 (N_1618,N_795,N_811);
nor U1619 (N_1619,N_961,N_702);
and U1620 (N_1620,N_387,N_823);
or U1621 (N_1621,N_901,N_410);
or U1622 (N_1622,N_2,N_378);
or U1623 (N_1623,N_297,N_707);
nor U1624 (N_1624,N_724,N_128);
nor U1625 (N_1625,N_320,N_991);
or U1626 (N_1626,N_441,N_31);
nand U1627 (N_1627,N_406,N_966);
nand U1628 (N_1628,N_808,N_120);
nand U1629 (N_1629,N_681,N_110);
nand U1630 (N_1630,N_181,N_925);
nor U1631 (N_1631,N_486,N_186);
nor U1632 (N_1632,N_391,N_674);
or U1633 (N_1633,N_573,N_418);
nand U1634 (N_1634,N_890,N_652);
nor U1635 (N_1635,N_871,N_471);
and U1636 (N_1636,N_840,N_191);
nor U1637 (N_1637,N_857,N_896);
nor U1638 (N_1638,N_234,N_594);
or U1639 (N_1639,N_726,N_948);
or U1640 (N_1640,N_500,N_160);
nor U1641 (N_1641,N_584,N_894);
nor U1642 (N_1642,N_600,N_874);
xor U1643 (N_1643,N_800,N_136);
nor U1644 (N_1644,N_448,N_88);
xor U1645 (N_1645,N_719,N_384);
nand U1646 (N_1646,N_125,N_432);
nand U1647 (N_1647,N_395,N_223);
or U1648 (N_1648,N_145,N_929);
and U1649 (N_1649,N_122,N_581);
and U1650 (N_1650,N_125,N_667);
or U1651 (N_1651,N_861,N_501);
nor U1652 (N_1652,N_52,N_605);
nor U1653 (N_1653,N_811,N_792);
and U1654 (N_1654,N_960,N_469);
nand U1655 (N_1655,N_422,N_415);
nor U1656 (N_1656,N_904,N_793);
or U1657 (N_1657,N_6,N_948);
or U1658 (N_1658,N_603,N_963);
or U1659 (N_1659,N_390,N_203);
and U1660 (N_1660,N_599,N_159);
or U1661 (N_1661,N_700,N_38);
and U1662 (N_1662,N_680,N_576);
nand U1663 (N_1663,N_801,N_361);
or U1664 (N_1664,N_687,N_765);
nand U1665 (N_1665,N_733,N_776);
and U1666 (N_1666,N_518,N_623);
nor U1667 (N_1667,N_153,N_849);
xnor U1668 (N_1668,N_894,N_128);
and U1669 (N_1669,N_116,N_236);
or U1670 (N_1670,N_781,N_543);
nand U1671 (N_1671,N_924,N_910);
and U1672 (N_1672,N_754,N_61);
or U1673 (N_1673,N_156,N_590);
nor U1674 (N_1674,N_941,N_519);
nand U1675 (N_1675,N_56,N_63);
and U1676 (N_1676,N_680,N_957);
or U1677 (N_1677,N_272,N_263);
nor U1678 (N_1678,N_516,N_925);
or U1679 (N_1679,N_714,N_707);
nand U1680 (N_1680,N_633,N_116);
nand U1681 (N_1681,N_589,N_425);
nor U1682 (N_1682,N_263,N_645);
nor U1683 (N_1683,N_570,N_167);
nor U1684 (N_1684,N_944,N_360);
nand U1685 (N_1685,N_915,N_125);
nor U1686 (N_1686,N_624,N_992);
nor U1687 (N_1687,N_861,N_855);
or U1688 (N_1688,N_623,N_442);
nor U1689 (N_1689,N_172,N_412);
or U1690 (N_1690,N_441,N_377);
or U1691 (N_1691,N_516,N_333);
nor U1692 (N_1692,N_251,N_894);
and U1693 (N_1693,N_971,N_534);
or U1694 (N_1694,N_280,N_304);
nand U1695 (N_1695,N_44,N_920);
nor U1696 (N_1696,N_862,N_600);
and U1697 (N_1697,N_426,N_8);
nor U1698 (N_1698,N_109,N_257);
nand U1699 (N_1699,N_593,N_33);
and U1700 (N_1700,N_657,N_925);
nand U1701 (N_1701,N_1,N_774);
or U1702 (N_1702,N_400,N_503);
or U1703 (N_1703,N_96,N_101);
nor U1704 (N_1704,N_135,N_231);
nand U1705 (N_1705,N_673,N_717);
xnor U1706 (N_1706,N_437,N_140);
xnor U1707 (N_1707,N_306,N_6);
nor U1708 (N_1708,N_670,N_674);
nor U1709 (N_1709,N_319,N_987);
and U1710 (N_1710,N_391,N_244);
nand U1711 (N_1711,N_888,N_271);
nand U1712 (N_1712,N_490,N_635);
nand U1713 (N_1713,N_273,N_207);
and U1714 (N_1714,N_268,N_461);
nor U1715 (N_1715,N_915,N_872);
nor U1716 (N_1716,N_179,N_421);
and U1717 (N_1717,N_971,N_954);
and U1718 (N_1718,N_745,N_779);
nand U1719 (N_1719,N_600,N_230);
or U1720 (N_1720,N_994,N_881);
and U1721 (N_1721,N_255,N_702);
nor U1722 (N_1722,N_308,N_330);
nand U1723 (N_1723,N_368,N_654);
xnor U1724 (N_1724,N_260,N_452);
or U1725 (N_1725,N_656,N_726);
nor U1726 (N_1726,N_981,N_286);
or U1727 (N_1727,N_722,N_805);
or U1728 (N_1728,N_819,N_309);
or U1729 (N_1729,N_970,N_630);
and U1730 (N_1730,N_77,N_592);
and U1731 (N_1731,N_601,N_168);
nand U1732 (N_1732,N_89,N_350);
nand U1733 (N_1733,N_504,N_244);
nor U1734 (N_1734,N_889,N_805);
nor U1735 (N_1735,N_859,N_181);
nand U1736 (N_1736,N_835,N_771);
nor U1737 (N_1737,N_0,N_10);
nor U1738 (N_1738,N_51,N_106);
nand U1739 (N_1739,N_628,N_903);
nor U1740 (N_1740,N_229,N_356);
or U1741 (N_1741,N_85,N_441);
and U1742 (N_1742,N_334,N_547);
nand U1743 (N_1743,N_866,N_429);
and U1744 (N_1744,N_411,N_948);
and U1745 (N_1745,N_348,N_347);
nor U1746 (N_1746,N_297,N_553);
nand U1747 (N_1747,N_846,N_966);
or U1748 (N_1748,N_923,N_932);
nor U1749 (N_1749,N_628,N_673);
nor U1750 (N_1750,N_532,N_782);
nor U1751 (N_1751,N_477,N_263);
nand U1752 (N_1752,N_392,N_767);
nand U1753 (N_1753,N_629,N_393);
nor U1754 (N_1754,N_582,N_554);
nor U1755 (N_1755,N_55,N_206);
or U1756 (N_1756,N_931,N_275);
nand U1757 (N_1757,N_826,N_165);
or U1758 (N_1758,N_715,N_967);
or U1759 (N_1759,N_214,N_169);
and U1760 (N_1760,N_620,N_150);
and U1761 (N_1761,N_937,N_18);
nand U1762 (N_1762,N_611,N_990);
or U1763 (N_1763,N_997,N_895);
and U1764 (N_1764,N_526,N_679);
nor U1765 (N_1765,N_405,N_729);
nor U1766 (N_1766,N_290,N_596);
and U1767 (N_1767,N_440,N_380);
and U1768 (N_1768,N_695,N_920);
and U1769 (N_1769,N_802,N_339);
or U1770 (N_1770,N_417,N_379);
xor U1771 (N_1771,N_864,N_182);
nor U1772 (N_1772,N_909,N_270);
nand U1773 (N_1773,N_580,N_136);
nand U1774 (N_1774,N_276,N_943);
and U1775 (N_1775,N_983,N_124);
and U1776 (N_1776,N_119,N_677);
or U1777 (N_1777,N_173,N_279);
nor U1778 (N_1778,N_444,N_191);
and U1779 (N_1779,N_962,N_951);
and U1780 (N_1780,N_898,N_464);
and U1781 (N_1781,N_251,N_170);
or U1782 (N_1782,N_424,N_542);
nor U1783 (N_1783,N_400,N_162);
or U1784 (N_1784,N_516,N_644);
and U1785 (N_1785,N_593,N_922);
nor U1786 (N_1786,N_504,N_623);
nor U1787 (N_1787,N_390,N_509);
nor U1788 (N_1788,N_304,N_988);
or U1789 (N_1789,N_11,N_164);
nand U1790 (N_1790,N_763,N_862);
and U1791 (N_1791,N_488,N_179);
nor U1792 (N_1792,N_733,N_778);
nor U1793 (N_1793,N_396,N_185);
nand U1794 (N_1794,N_592,N_579);
and U1795 (N_1795,N_781,N_90);
nand U1796 (N_1796,N_178,N_915);
or U1797 (N_1797,N_490,N_119);
and U1798 (N_1798,N_665,N_827);
and U1799 (N_1799,N_418,N_600);
and U1800 (N_1800,N_502,N_104);
or U1801 (N_1801,N_809,N_638);
and U1802 (N_1802,N_383,N_328);
and U1803 (N_1803,N_363,N_644);
nor U1804 (N_1804,N_799,N_203);
and U1805 (N_1805,N_617,N_291);
nand U1806 (N_1806,N_730,N_294);
and U1807 (N_1807,N_507,N_9);
nand U1808 (N_1808,N_58,N_259);
nand U1809 (N_1809,N_526,N_869);
or U1810 (N_1810,N_258,N_0);
and U1811 (N_1811,N_647,N_99);
and U1812 (N_1812,N_426,N_952);
nand U1813 (N_1813,N_696,N_695);
and U1814 (N_1814,N_237,N_555);
and U1815 (N_1815,N_720,N_358);
nor U1816 (N_1816,N_567,N_308);
or U1817 (N_1817,N_845,N_215);
nand U1818 (N_1818,N_365,N_645);
nand U1819 (N_1819,N_970,N_9);
or U1820 (N_1820,N_962,N_532);
or U1821 (N_1821,N_39,N_959);
nor U1822 (N_1822,N_326,N_302);
nor U1823 (N_1823,N_87,N_45);
and U1824 (N_1824,N_172,N_267);
or U1825 (N_1825,N_832,N_184);
xor U1826 (N_1826,N_887,N_29);
nand U1827 (N_1827,N_125,N_828);
nand U1828 (N_1828,N_75,N_156);
nor U1829 (N_1829,N_531,N_552);
or U1830 (N_1830,N_809,N_695);
and U1831 (N_1831,N_262,N_520);
or U1832 (N_1832,N_603,N_410);
nand U1833 (N_1833,N_273,N_593);
nor U1834 (N_1834,N_969,N_172);
and U1835 (N_1835,N_863,N_287);
or U1836 (N_1836,N_896,N_251);
or U1837 (N_1837,N_919,N_198);
nor U1838 (N_1838,N_853,N_203);
and U1839 (N_1839,N_618,N_302);
and U1840 (N_1840,N_1,N_302);
nor U1841 (N_1841,N_886,N_935);
nand U1842 (N_1842,N_945,N_65);
and U1843 (N_1843,N_571,N_288);
nand U1844 (N_1844,N_322,N_837);
xor U1845 (N_1845,N_558,N_903);
nand U1846 (N_1846,N_253,N_267);
nor U1847 (N_1847,N_17,N_344);
and U1848 (N_1848,N_22,N_719);
or U1849 (N_1849,N_524,N_10);
or U1850 (N_1850,N_709,N_514);
nor U1851 (N_1851,N_840,N_701);
and U1852 (N_1852,N_323,N_328);
and U1853 (N_1853,N_379,N_21);
nand U1854 (N_1854,N_325,N_295);
and U1855 (N_1855,N_455,N_582);
and U1856 (N_1856,N_373,N_769);
xor U1857 (N_1857,N_344,N_713);
and U1858 (N_1858,N_620,N_57);
and U1859 (N_1859,N_143,N_177);
nor U1860 (N_1860,N_695,N_932);
nor U1861 (N_1861,N_181,N_661);
nor U1862 (N_1862,N_968,N_204);
nor U1863 (N_1863,N_16,N_942);
nand U1864 (N_1864,N_267,N_769);
or U1865 (N_1865,N_667,N_856);
or U1866 (N_1866,N_518,N_8);
nand U1867 (N_1867,N_807,N_726);
and U1868 (N_1868,N_569,N_45);
nand U1869 (N_1869,N_957,N_959);
and U1870 (N_1870,N_94,N_420);
and U1871 (N_1871,N_224,N_634);
nand U1872 (N_1872,N_595,N_141);
nor U1873 (N_1873,N_905,N_33);
nor U1874 (N_1874,N_619,N_645);
or U1875 (N_1875,N_318,N_958);
nor U1876 (N_1876,N_617,N_75);
nand U1877 (N_1877,N_681,N_489);
or U1878 (N_1878,N_85,N_623);
nor U1879 (N_1879,N_153,N_850);
and U1880 (N_1880,N_374,N_132);
nor U1881 (N_1881,N_724,N_108);
nand U1882 (N_1882,N_338,N_968);
nor U1883 (N_1883,N_685,N_938);
and U1884 (N_1884,N_792,N_141);
nand U1885 (N_1885,N_943,N_315);
nand U1886 (N_1886,N_156,N_190);
nand U1887 (N_1887,N_884,N_779);
nand U1888 (N_1888,N_30,N_299);
nor U1889 (N_1889,N_993,N_788);
nor U1890 (N_1890,N_867,N_434);
nor U1891 (N_1891,N_729,N_215);
nand U1892 (N_1892,N_779,N_105);
or U1893 (N_1893,N_582,N_332);
or U1894 (N_1894,N_762,N_996);
nand U1895 (N_1895,N_330,N_608);
and U1896 (N_1896,N_463,N_581);
xor U1897 (N_1897,N_891,N_136);
and U1898 (N_1898,N_71,N_673);
and U1899 (N_1899,N_524,N_343);
or U1900 (N_1900,N_494,N_867);
and U1901 (N_1901,N_843,N_646);
nor U1902 (N_1902,N_668,N_136);
nand U1903 (N_1903,N_601,N_768);
or U1904 (N_1904,N_795,N_78);
nor U1905 (N_1905,N_800,N_653);
nor U1906 (N_1906,N_854,N_548);
nand U1907 (N_1907,N_603,N_540);
nand U1908 (N_1908,N_887,N_700);
nand U1909 (N_1909,N_608,N_631);
nand U1910 (N_1910,N_837,N_143);
nor U1911 (N_1911,N_986,N_196);
nor U1912 (N_1912,N_237,N_397);
or U1913 (N_1913,N_617,N_205);
nor U1914 (N_1914,N_377,N_122);
or U1915 (N_1915,N_92,N_955);
and U1916 (N_1916,N_300,N_168);
and U1917 (N_1917,N_147,N_446);
and U1918 (N_1918,N_978,N_859);
and U1919 (N_1919,N_61,N_223);
or U1920 (N_1920,N_410,N_565);
and U1921 (N_1921,N_792,N_45);
or U1922 (N_1922,N_246,N_333);
nand U1923 (N_1923,N_477,N_145);
and U1924 (N_1924,N_449,N_635);
and U1925 (N_1925,N_400,N_770);
and U1926 (N_1926,N_895,N_84);
and U1927 (N_1927,N_712,N_574);
and U1928 (N_1928,N_924,N_391);
and U1929 (N_1929,N_7,N_396);
nor U1930 (N_1930,N_414,N_759);
and U1931 (N_1931,N_516,N_240);
or U1932 (N_1932,N_740,N_744);
and U1933 (N_1933,N_349,N_169);
nor U1934 (N_1934,N_134,N_962);
nor U1935 (N_1935,N_293,N_891);
nor U1936 (N_1936,N_53,N_492);
nor U1937 (N_1937,N_81,N_807);
or U1938 (N_1938,N_237,N_57);
nor U1939 (N_1939,N_867,N_767);
nand U1940 (N_1940,N_667,N_454);
or U1941 (N_1941,N_774,N_405);
nand U1942 (N_1942,N_415,N_575);
and U1943 (N_1943,N_162,N_907);
or U1944 (N_1944,N_35,N_400);
nand U1945 (N_1945,N_868,N_874);
or U1946 (N_1946,N_164,N_978);
or U1947 (N_1947,N_977,N_340);
nor U1948 (N_1948,N_935,N_56);
or U1949 (N_1949,N_160,N_829);
and U1950 (N_1950,N_84,N_280);
and U1951 (N_1951,N_575,N_926);
or U1952 (N_1952,N_345,N_792);
or U1953 (N_1953,N_513,N_338);
and U1954 (N_1954,N_301,N_155);
nand U1955 (N_1955,N_393,N_505);
nor U1956 (N_1956,N_522,N_806);
nor U1957 (N_1957,N_774,N_764);
or U1958 (N_1958,N_412,N_915);
and U1959 (N_1959,N_426,N_658);
or U1960 (N_1960,N_891,N_693);
nor U1961 (N_1961,N_929,N_16);
nor U1962 (N_1962,N_357,N_467);
nor U1963 (N_1963,N_824,N_673);
or U1964 (N_1964,N_201,N_391);
nor U1965 (N_1965,N_228,N_282);
nor U1966 (N_1966,N_149,N_738);
nor U1967 (N_1967,N_128,N_776);
or U1968 (N_1968,N_572,N_399);
xnor U1969 (N_1969,N_161,N_706);
nor U1970 (N_1970,N_326,N_627);
or U1971 (N_1971,N_517,N_999);
nand U1972 (N_1972,N_699,N_568);
or U1973 (N_1973,N_519,N_96);
nand U1974 (N_1974,N_888,N_765);
nor U1975 (N_1975,N_946,N_404);
nand U1976 (N_1976,N_598,N_874);
and U1977 (N_1977,N_944,N_279);
nor U1978 (N_1978,N_960,N_930);
and U1979 (N_1979,N_296,N_914);
xnor U1980 (N_1980,N_101,N_361);
and U1981 (N_1981,N_922,N_647);
and U1982 (N_1982,N_157,N_750);
and U1983 (N_1983,N_120,N_820);
nand U1984 (N_1984,N_976,N_279);
nor U1985 (N_1985,N_520,N_165);
or U1986 (N_1986,N_349,N_874);
nand U1987 (N_1987,N_856,N_806);
nand U1988 (N_1988,N_562,N_902);
nor U1989 (N_1989,N_703,N_531);
and U1990 (N_1990,N_238,N_875);
or U1991 (N_1991,N_130,N_248);
and U1992 (N_1992,N_274,N_326);
nand U1993 (N_1993,N_162,N_127);
and U1994 (N_1994,N_891,N_830);
or U1995 (N_1995,N_353,N_960);
nor U1996 (N_1996,N_277,N_528);
or U1997 (N_1997,N_353,N_837);
or U1998 (N_1998,N_197,N_4);
nand U1999 (N_1999,N_802,N_859);
nor U2000 (N_2000,N_1776,N_1996);
and U2001 (N_2001,N_1139,N_1701);
and U2002 (N_2002,N_1081,N_1619);
nand U2003 (N_2003,N_1568,N_1461);
or U2004 (N_2004,N_1625,N_1954);
and U2005 (N_2005,N_1246,N_1698);
nor U2006 (N_2006,N_1407,N_1831);
or U2007 (N_2007,N_1021,N_1880);
or U2008 (N_2008,N_1377,N_1800);
nor U2009 (N_2009,N_1828,N_1593);
or U2010 (N_2010,N_1662,N_1026);
and U2011 (N_2011,N_1840,N_1463);
nor U2012 (N_2012,N_1218,N_1849);
or U2013 (N_2013,N_1865,N_1882);
nor U2014 (N_2014,N_1319,N_1522);
and U2015 (N_2015,N_1303,N_1755);
and U2016 (N_2016,N_1567,N_1757);
or U2017 (N_2017,N_1200,N_1771);
and U2018 (N_2018,N_1358,N_1927);
and U2019 (N_2019,N_1342,N_1496);
and U2020 (N_2020,N_1846,N_1607);
and U2021 (N_2021,N_1029,N_1844);
xor U2022 (N_2022,N_1613,N_1042);
or U2023 (N_2023,N_1624,N_1862);
and U2024 (N_2024,N_1864,N_1942);
nor U2025 (N_2025,N_1122,N_1648);
nand U2026 (N_2026,N_1052,N_1403);
nor U2027 (N_2027,N_1657,N_1529);
nand U2028 (N_2028,N_1451,N_1684);
nand U2029 (N_2029,N_1580,N_1136);
or U2030 (N_2030,N_1510,N_1527);
nand U2031 (N_2031,N_1813,N_1804);
nor U2032 (N_2032,N_1105,N_1413);
nor U2033 (N_2033,N_1353,N_1266);
nor U2034 (N_2034,N_1815,N_1896);
or U2035 (N_2035,N_1868,N_1752);
nand U2036 (N_2036,N_1202,N_1082);
nor U2037 (N_2037,N_1298,N_1090);
nand U2038 (N_2038,N_1273,N_1396);
nor U2039 (N_2039,N_1857,N_1229);
or U2040 (N_2040,N_1208,N_1498);
xor U2041 (N_2041,N_1426,N_1751);
nor U2042 (N_2042,N_1159,N_1723);
and U2043 (N_2043,N_1276,N_1732);
nand U2044 (N_2044,N_1677,N_1025);
nand U2045 (N_2045,N_1274,N_1913);
nor U2046 (N_2046,N_1307,N_1700);
nand U2047 (N_2047,N_1577,N_1295);
and U2048 (N_2048,N_1111,N_1656);
nor U2049 (N_2049,N_1950,N_1576);
nand U2050 (N_2050,N_1489,N_1121);
and U2051 (N_2051,N_1057,N_1412);
nor U2052 (N_2052,N_1243,N_1308);
and U2053 (N_2053,N_1022,N_1038);
nand U2054 (N_2054,N_1615,N_1690);
nand U2055 (N_2055,N_1141,N_1346);
and U2056 (N_2056,N_1311,N_1907);
xor U2057 (N_2057,N_1670,N_1309);
nor U2058 (N_2058,N_1058,N_1877);
nand U2059 (N_2059,N_1505,N_1742);
nor U2060 (N_2060,N_1124,N_1545);
and U2061 (N_2061,N_1419,N_1211);
nor U2062 (N_2062,N_1939,N_1334);
and U2063 (N_2063,N_1088,N_1083);
nand U2064 (N_2064,N_1245,N_1989);
nand U2065 (N_2065,N_1251,N_1078);
and U2066 (N_2066,N_1934,N_1736);
or U2067 (N_2067,N_1340,N_1036);
or U2068 (N_2068,N_1630,N_1447);
nor U2069 (N_2069,N_1195,N_1129);
nor U2070 (N_2070,N_1649,N_1578);
or U2071 (N_2071,N_1914,N_1949);
or U2072 (N_2072,N_1360,N_1879);
nand U2073 (N_2073,N_1370,N_1720);
and U2074 (N_2074,N_1957,N_1571);
nand U2075 (N_2075,N_1374,N_1287);
nand U2076 (N_2076,N_1014,N_1724);
or U2077 (N_2077,N_1620,N_1401);
xnor U2078 (N_2078,N_1556,N_1661);
nor U2079 (N_2079,N_1803,N_1119);
or U2080 (N_2080,N_1151,N_1910);
or U2081 (N_2081,N_1772,N_1693);
nor U2082 (N_2082,N_1970,N_1676);
xnor U2083 (N_2083,N_1532,N_1156);
nor U2084 (N_2084,N_1063,N_1850);
and U2085 (N_2085,N_1509,N_1232);
or U2086 (N_2086,N_1688,N_1660);
nand U2087 (N_2087,N_1092,N_1691);
nor U2088 (N_2088,N_1219,N_1833);
nand U2089 (N_2089,N_1912,N_1060);
nor U2090 (N_2090,N_1521,N_1854);
nand U2091 (N_2091,N_1997,N_1591);
and U2092 (N_2092,N_1381,N_1956);
or U2093 (N_2093,N_1250,N_1982);
nand U2094 (N_2094,N_1196,N_1668);
and U2095 (N_2095,N_1429,N_1127);
and U2096 (N_2096,N_1427,N_1493);
nand U2097 (N_2097,N_1476,N_1100);
or U2098 (N_2098,N_1260,N_1599);
and U2099 (N_2099,N_1174,N_1801);
or U2100 (N_2100,N_1045,N_1627);
nand U2101 (N_2101,N_1074,N_1255);
nor U2102 (N_2102,N_1711,N_1290);
and U2103 (N_2103,N_1695,N_1072);
nand U2104 (N_2104,N_1399,N_1992);
nor U2105 (N_2105,N_1550,N_1442);
nor U2106 (N_2106,N_1935,N_1456);
nand U2107 (N_2107,N_1023,N_1838);
and U2108 (N_2108,N_1604,N_1589);
and U2109 (N_2109,N_1969,N_1796);
or U2110 (N_2110,N_1972,N_1728);
nor U2111 (N_2111,N_1408,N_1157);
nand U2112 (N_2112,N_1533,N_1280);
nand U2113 (N_2113,N_1183,N_1528);
or U2114 (N_2114,N_1192,N_1165);
nand U2115 (N_2115,N_1128,N_1512);
or U2116 (N_2116,N_1397,N_1486);
nand U2117 (N_2117,N_1337,N_1973);
and U2118 (N_2118,N_1712,N_1046);
nand U2119 (N_2119,N_1786,N_1194);
nor U2120 (N_2120,N_1393,N_1453);
or U2121 (N_2121,N_1106,N_1985);
nor U2122 (N_2122,N_1988,N_1908);
and U2123 (N_2123,N_1836,N_1123);
nand U2124 (N_2124,N_1548,N_1080);
or U2125 (N_2125,N_1653,N_1125);
nand U2126 (N_2126,N_1317,N_1481);
and U2127 (N_2127,N_1318,N_1924);
nor U2128 (N_2128,N_1071,N_1717);
or U2129 (N_2129,N_1714,N_1707);
or U2130 (N_2130,N_1416,N_1859);
nor U2131 (N_2131,N_1806,N_1050);
or U2132 (N_2132,N_1437,N_1704);
or U2133 (N_2133,N_1542,N_1596);
and U2134 (N_2134,N_1323,N_1254);
or U2135 (N_2135,N_1076,N_1172);
nor U2136 (N_2136,N_1055,N_1637);
or U2137 (N_2137,N_1602,N_1301);
nor U2138 (N_2138,N_1696,N_1663);
nand U2139 (N_2139,N_1733,N_1978);
nor U2140 (N_2140,N_1465,N_1600);
nor U2141 (N_2141,N_1686,N_1976);
and U2142 (N_2142,N_1802,N_1356);
nor U2143 (N_2143,N_1858,N_1009);
nor U2144 (N_2144,N_1333,N_1573);
nor U2145 (N_2145,N_1418,N_1530);
and U2146 (N_2146,N_1570,N_1007);
nand U2147 (N_2147,N_1537,N_1645);
nor U2148 (N_2148,N_1448,N_1561);
nor U2149 (N_2149,N_1146,N_1765);
and U2150 (N_2150,N_1424,N_1513);
nand U2151 (N_2151,N_1264,N_1906);
or U2152 (N_2152,N_1584,N_1843);
nor U2153 (N_2153,N_1227,N_1807);
and U2154 (N_2154,N_1117,N_1108);
nor U2155 (N_2155,N_1061,N_1926);
or U2156 (N_2156,N_1147,N_1197);
nor U2157 (N_2157,N_1998,N_1873);
nor U2158 (N_2158,N_1932,N_1839);
or U2159 (N_2159,N_1856,N_1727);
nand U2160 (N_2160,N_1500,N_1352);
or U2161 (N_2161,N_1047,N_1341);
nor U2162 (N_2162,N_1737,N_1034);
and U2163 (N_2163,N_1310,N_1626);
nor U2164 (N_2164,N_1654,N_1941);
and U2165 (N_2165,N_1595,N_1415);
and U2166 (N_2166,N_1820,N_1169);
nor U2167 (N_2167,N_1256,N_1778);
and U2168 (N_2168,N_1889,N_1581);
nand U2169 (N_2169,N_1716,N_1709);
or U2170 (N_2170,N_1164,N_1937);
nor U2171 (N_2171,N_1344,N_1763);
and U2172 (N_2172,N_1443,N_1073);
nor U2173 (N_2173,N_1488,N_1919);
xor U2174 (N_2174,N_1313,N_1735);
nand U2175 (N_2175,N_1261,N_1475);
and U2176 (N_2176,N_1592,N_1790);
nor U2177 (N_2177,N_1621,N_1940);
or U2178 (N_2178,N_1903,N_1553);
and U2179 (N_2179,N_1634,N_1491);
nor U2180 (N_2180,N_1968,N_1039);
or U2181 (N_2181,N_1909,N_1470);
xnor U2182 (N_2182,N_1462,N_1137);
nand U2183 (N_2183,N_1205,N_1135);
or U2184 (N_2184,N_1030,N_1984);
nor U2185 (N_2185,N_1086,N_1417);
nand U2186 (N_2186,N_1430,N_1093);
nor U2187 (N_2187,N_1354,N_1361);
and U2188 (N_2188,N_1198,N_1872);
nor U2189 (N_2189,N_1239,N_1874);
or U2190 (N_2190,N_1345,N_1897);
and U2191 (N_2191,N_1925,N_1841);
nand U2192 (N_2192,N_1569,N_1871);
and U2193 (N_2193,N_1945,N_1678);
and U2194 (N_2194,N_1446,N_1331);
nand U2195 (N_2195,N_1726,N_1444);
nor U2196 (N_2196,N_1632,N_1975);
xnor U2197 (N_2197,N_1506,N_1845);
nor U2198 (N_2198,N_1638,N_1441);
nor U2199 (N_2199,N_1699,N_1233);
or U2200 (N_2200,N_1702,N_1269);
nand U2201 (N_2201,N_1517,N_1759);
or U2202 (N_2202,N_1368,N_1881);
nand U2203 (N_2203,N_1162,N_1473);
nand U2204 (N_2204,N_1785,N_1990);
or U2205 (N_2205,N_1434,N_1915);
nor U2206 (N_2206,N_1618,N_1911);
or U2207 (N_2207,N_1155,N_1284);
and U2208 (N_2208,N_1019,N_1952);
nor U2209 (N_2209,N_1375,N_1750);
and U2210 (N_2210,N_1962,N_1249);
nor U2211 (N_2211,N_1706,N_1546);
and U2212 (N_2212,N_1214,N_1758);
or U2213 (N_2213,N_1431,N_1031);
nor U2214 (N_2214,N_1224,N_1003);
nand U2215 (N_2215,N_1543,N_1824);
and U2216 (N_2216,N_1299,N_1348);
and U2217 (N_2217,N_1501,N_1275);
and U2218 (N_2218,N_1979,N_1540);
and U2219 (N_2219,N_1539,N_1390);
and U2220 (N_2220,N_1821,N_1452);
and U2221 (N_2221,N_1837,N_1760);
nand U2222 (N_2222,N_1715,N_1414);
and U2223 (N_2223,N_1213,N_1876);
nand U2224 (N_2224,N_1102,N_1667);
nor U2225 (N_2225,N_1575,N_1536);
nor U2226 (N_2226,N_1328,N_1458);
nand U2227 (N_2227,N_1015,N_1885);
nand U2228 (N_2228,N_1633,N_1469);
or U2229 (N_2229,N_1244,N_1349);
or U2230 (N_2230,N_1054,N_1705);
or U2231 (N_2231,N_1495,N_1296);
xor U2232 (N_2232,N_1499,N_1114);
xnor U2233 (N_2233,N_1207,N_1566);
xor U2234 (N_2234,N_1916,N_1432);
nand U2235 (N_2235,N_1297,N_1226);
nor U2236 (N_2236,N_1142,N_1177);
nand U2237 (N_2237,N_1825,N_1248);
or U2238 (N_2238,N_1423,N_1107);
nand U2239 (N_2239,N_1235,N_1692);
nor U2240 (N_2240,N_1209,N_1930);
nor U2241 (N_2241,N_1904,N_1756);
nand U2242 (N_2242,N_1380,N_1372);
nor U2243 (N_2243,N_1049,N_1267);
nor U2244 (N_2244,N_1861,N_1109);
nor U2245 (N_2245,N_1336,N_1797);
and U2246 (N_2246,N_1193,N_1999);
nor U2247 (N_2247,N_1587,N_1258);
nand U2248 (N_2248,N_1449,N_1293);
and U2249 (N_2249,N_1572,N_1020);
and U2250 (N_2250,N_1236,N_1199);
nand U2251 (N_2251,N_1640,N_1314);
or U2252 (N_2252,N_1222,N_1161);
and U2253 (N_2253,N_1382,N_1819);
and U2254 (N_2254,N_1697,N_1773);
nand U2255 (N_2255,N_1673,N_1075);
and U2256 (N_2256,N_1775,N_1933);
nand U2257 (N_2257,N_1315,N_1321);
nand U2258 (N_2258,N_1094,N_1977);
nor U2259 (N_2259,N_1270,N_1748);
nand U2260 (N_2260,N_1731,N_1863);
nand U2261 (N_2261,N_1464,N_1835);
or U2262 (N_2262,N_1466,N_1823);
or U2263 (N_2263,N_1410,N_1579);
or U2264 (N_2264,N_1585,N_1622);
nor U2265 (N_2265,N_1987,N_1379);
and U2266 (N_2266,N_1671,N_1631);
or U2267 (N_2267,N_1886,N_1791);
and U2268 (N_2268,N_1703,N_1520);
xor U2269 (N_2269,N_1069,N_1212);
nand U2270 (N_2270,N_1822,N_1883);
or U2271 (N_2271,N_1383,N_1118);
nand U2272 (N_2272,N_1544,N_1641);
nand U2273 (N_2273,N_1422,N_1669);
or U2274 (N_2274,N_1944,N_1901);
nand U2275 (N_2275,N_1629,N_1253);
and U2276 (N_2276,N_1203,N_1611);
nand U2277 (N_2277,N_1095,N_1289);
or U2278 (N_2278,N_1384,N_1689);
nand U2279 (N_2279,N_1001,N_1190);
and U2280 (N_2280,N_1482,N_1044);
or U2281 (N_2281,N_1325,N_1508);
nand U2282 (N_2282,N_1767,N_1875);
nand U2283 (N_2283,N_1666,N_1206);
nand U2284 (N_2284,N_1744,N_1980);
or U2285 (N_2285,N_1518,N_1048);
nand U2286 (N_2286,N_1745,N_1394);
or U2287 (N_2287,N_1981,N_1598);
or U2288 (N_2288,N_1826,N_1175);
nor U2289 (N_2289,N_1217,N_1739);
or U2290 (N_2290,N_1718,N_1000);
nor U2291 (N_2291,N_1643,N_1163);
nand U2292 (N_2292,N_1268,N_1525);
nand U2293 (N_2293,N_1597,N_1035);
and U2294 (N_2294,N_1582,N_1339);
nor U2295 (N_2295,N_1409,N_1762);
nor U2296 (N_2296,N_1898,N_1178);
and U2297 (N_2297,N_1832,N_1016);
and U2298 (N_2298,N_1490,N_1818);
nand U2299 (N_2299,N_1960,N_1257);
nor U2300 (N_2300,N_1247,N_1497);
nor U2301 (N_2301,N_1829,N_1893);
or U2302 (N_2302,N_1590,N_1112);
or U2303 (N_2303,N_1355,N_1167);
and U2304 (N_2304,N_1869,N_1552);
and U2305 (N_2305,N_1316,N_1535);
and U2306 (N_2306,N_1168,N_1768);
and U2307 (N_2307,N_1900,N_1974);
or U2308 (N_2308,N_1387,N_1385);
or U2309 (N_2309,N_1359,N_1655);
nor U2310 (N_2310,N_1555,N_1665);
nand U2311 (N_2311,N_1004,N_1067);
and U2312 (N_2312,N_1484,N_1089);
or U2313 (N_2313,N_1428,N_1779);
nor U2314 (N_2314,N_1805,N_1281);
nor U2315 (N_2315,N_1378,N_1398);
and U2316 (N_2316,N_1616,N_1842);
nand U2317 (N_2317,N_1240,N_1799);
or U2318 (N_2318,N_1764,N_1460);
and U2319 (N_2319,N_1005,N_1526);
nor U2320 (N_2320,N_1445,N_1320);
or U2321 (N_2321,N_1734,N_1792);
nand U2322 (N_2322,N_1766,N_1562);
or U2323 (N_2323,N_1636,N_1483);
xnor U2324 (N_2324,N_1391,N_1965);
or U2325 (N_2325,N_1010,N_1524);
nor U2326 (N_2326,N_1187,N_1614);
and U2327 (N_2327,N_1955,N_1514);
and U2328 (N_2328,N_1130,N_1652);
or U2329 (N_2329,N_1606,N_1215);
nand U2330 (N_2330,N_1586,N_1938);
or U2331 (N_2331,N_1326,N_1783);
nand U2332 (N_2332,N_1558,N_1182);
nand U2333 (N_2333,N_1721,N_1420);
or U2334 (N_2334,N_1923,N_1347);
or U2335 (N_2335,N_1583,N_1888);
nor U2336 (N_2336,N_1120,N_1116);
or U2337 (N_2337,N_1811,N_1302);
xor U2338 (N_2338,N_1389,N_1180);
or U2339 (N_2339,N_1421,N_1395);
nand U2340 (N_2340,N_1551,N_1033);
nor U2341 (N_2341,N_1787,N_1133);
or U2342 (N_2342,N_1097,N_1754);
nor U2343 (N_2343,N_1158,N_1131);
nor U2344 (N_2344,N_1574,N_1740);
or U2345 (N_2345,N_1966,N_1563);
and U2346 (N_2346,N_1793,N_1292);
nand U2347 (N_2347,N_1467,N_1230);
nor U2348 (N_2348,N_1436,N_1639);
nand U2349 (N_2349,N_1152,N_1515);
and U2350 (N_2350,N_1892,N_1931);
or U2351 (N_2351,N_1221,N_1210);
and U2352 (N_2352,N_1189,N_1332);
and U2353 (N_2353,N_1376,N_1134);
and U2354 (N_2354,N_1145,N_1810);
nor U2355 (N_2355,N_1008,N_1993);
and U2356 (N_2356,N_1343,N_1392);
nor U2357 (N_2357,N_1659,N_1995);
and U2358 (N_2358,N_1565,N_1983);
or U2359 (N_2359,N_1024,N_1674);
nor U2360 (N_2360,N_1743,N_1738);
nor U2361 (N_2361,N_1181,N_1357);
nor U2362 (N_2362,N_1781,N_1150);
and U2363 (N_2363,N_1948,N_1223);
or U2364 (N_2364,N_1782,N_1367);
or U2365 (N_2365,N_1459,N_1784);
or U2366 (N_2366,N_1064,N_1710);
nor U2367 (N_2367,N_1531,N_1472);
nand U2368 (N_2368,N_1478,N_1511);
or U2369 (N_2369,N_1241,N_1557);
or U2370 (N_2370,N_1288,N_1364);
or U2371 (N_2371,N_1032,N_1306);
nor U2372 (N_2372,N_1283,N_1770);
and U2373 (N_2373,N_1808,N_1730);
or U2374 (N_2374,N_1612,N_1855);
and U2375 (N_2375,N_1884,N_1679);
and U2376 (N_2376,N_1794,N_1062);
nand U2377 (N_2377,N_1848,N_1642);
nand U2378 (N_2378,N_1780,N_1680);
nand U2379 (N_2379,N_1827,N_1438);
nand U2380 (N_2380,N_1650,N_1601);
nand U2381 (N_2381,N_1503,N_1646);
or U2382 (N_2382,N_1485,N_1265);
nor U2383 (N_2383,N_1366,N_1994);
and U2384 (N_2384,N_1166,N_1946);
or U2385 (N_2385,N_1917,N_1492);
and U2386 (N_2386,N_1891,N_1285);
and U2387 (N_2387,N_1788,N_1371);
nand U2388 (N_2388,N_1160,N_1789);
nor U2389 (N_2389,N_1683,N_1623);
nor U2390 (N_2390,N_1746,N_1365);
or U2391 (N_2391,N_1282,N_1439);
nand U2392 (N_2392,N_1713,N_1651);
or U2393 (N_2393,N_1608,N_1610);
nor U2394 (N_2394,N_1675,N_1929);
nor U2395 (N_2395,N_1991,N_1184);
nand U2396 (N_2396,N_1435,N_1402);
nor U2397 (N_2397,N_1362,N_1400);
nor U2398 (N_2398,N_1644,N_1238);
nor U2399 (N_2399,N_1635,N_1018);
nand U2400 (N_2400,N_1959,N_1369);
nor U2401 (N_2401,N_1101,N_1685);
and U2402 (N_2402,N_1534,N_1936);
nor U2403 (N_2403,N_1065,N_1201);
nor U2404 (N_2404,N_1852,N_1719);
and U2405 (N_2405,N_1404,N_1263);
nor U2406 (N_2406,N_1068,N_1037);
or U2407 (N_2407,N_1087,N_1126);
nor U2408 (N_2408,N_1560,N_1279);
and U2409 (N_2409,N_1028,N_1363);
or U2410 (N_2410,N_1870,N_1468);
and U2411 (N_2411,N_1658,N_1225);
nor U2412 (N_2412,N_1457,N_1928);
or U2413 (N_2413,N_1853,N_1041);
and U2414 (N_2414,N_1694,N_1559);
and U2415 (N_2415,N_1887,N_1305);
or U2416 (N_2416,N_1110,N_1188);
nor U2417 (N_2417,N_1103,N_1216);
and U2418 (N_2418,N_1964,N_1958);
xor U2419 (N_2419,N_1170,N_1153);
nand U2420 (N_2420,N_1300,N_1228);
nor U2421 (N_2421,N_1741,N_1617);
nand U2422 (N_2422,N_1798,N_1549);
nand U2423 (N_2423,N_1091,N_1851);
or U2424 (N_2424,N_1040,N_1176);
and U2425 (N_2425,N_1605,N_1471);
and U2426 (N_2426,N_1053,N_1479);
and U2427 (N_2427,N_1132,N_1777);
nand U2428 (N_2428,N_1523,N_1272);
nor U2429 (N_2429,N_1330,N_1480);
nor U2430 (N_2430,N_1947,N_1507);
nand U2431 (N_2431,N_1011,N_1077);
nor U2432 (N_2432,N_1312,N_1830);
and U2433 (N_2433,N_1322,N_1753);
or U2434 (N_2434,N_1905,N_1749);
nand U2435 (N_2435,N_1259,N_1816);
nor U2436 (N_2436,N_1017,N_1277);
nor U2437 (N_2437,N_1411,N_1173);
nor U2438 (N_2438,N_1866,N_1204);
nand U2439 (N_2439,N_1477,N_1681);
xnor U2440 (N_2440,N_1234,N_1494);
and U2441 (N_2441,N_1943,N_1405);
or U2442 (N_2442,N_1388,N_1812);
and U2443 (N_2443,N_1725,N_1795);
nand U2444 (N_2444,N_1406,N_1327);
nor U2445 (N_2445,N_1487,N_1335);
or U2446 (N_2446,N_1350,N_1474);
nand U2447 (N_2447,N_1220,N_1847);
and U2448 (N_2448,N_1425,N_1967);
nand U2449 (N_2449,N_1971,N_1554);
nor U2450 (N_2450,N_1027,N_1113);
and U2451 (N_2451,N_1143,N_1538);
or U2452 (N_2452,N_1098,N_1304);
and U2453 (N_2453,N_1953,N_1099);
nor U2454 (N_2454,N_1138,N_1231);
and U2455 (N_2455,N_1179,N_1329);
and U2456 (N_2456,N_1096,N_1294);
nand U2457 (N_2457,N_1951,N_1729);
nor U2458 (N_2458,N_1708,N_1006);
nand U2459 (N_2459,N_1386,N_1252);
or U2460 (N_2460,N_1547,N_1070);
and U2461 (N_2461,N_1059,N_1051);
and U2462 (N_2462,N_1519,N_1043);
or U2463 (N_2463,N_1922,N_1056);
nand U2464 (N_2464,N_1154,N_1271);
nand U2465 (N_2465,N_1140,N_1085);
and U2466 (N_2466,N_1104,N_1440);
or U2467 (N_2467,N_1286,N_1687);
or U2468 (N_2468,N_1237,N_1373);
nand U2469 (N_2469,N_1594,N_1963);
and U2470 (N_2470,N_1867,N_1890);
xor U2471 (N_2471,N_1278,N_1920);
nor U2472 (N_2472,N_1609,N_1878);
or U2473 (N_2473,N_1860,N_1191);
and U2474 (N_2474,N_1986,N_1899);
nor U2475 (N_2475,N_1761,N_1809);
nor U2476 (N_2476,N_1291,N_1672);
nand U2477 (N_2477,N_1902,N_1682);
and U2478 (N_2478,N_1324,N_1894);
nor U2479 (N_2479,N_1262,N_1149);
nor U2480 (N_2480,N_1564,N_1171);
nand U2481 (N_2481,N_1603,N_1148);
and U2482 (N_2482,N_1013,N_1664);
nand U2483 (N_2483,N_1834,N_1921);
or U2484 (N_2484,N_1918,N_1186);
or U2485 (N_2485,N_1588,N_1079);
xor U2486 (N_2486,N_1454,N_1351);
nor U2487 (N_2487,N_1747,N_1455);
or U2488 (N_2488,N_1002,N_1722);
and U2489 (N_2489,N_1895,N_1433);
or U2490 (N_2490,N_1647,N_1450);
and U2491 (N_2491,N_1541,N_1012);
nor U2492 (N_2492,N_1504,N_1502);
or U2493 (N_2493,N_1144,N_1084);
and U2494 (N_2494,N_1185,N_1066);
or U2495 (N_2495,N_1516,N_1961);
or U2496 (N_2496,N_1628,N_1774);
nor U2497 (N_2497,N_1769,N_1242);
or U2498 (N_2498,N_1115,N_1338);
nor U2499 (N_2499,N_1814,N_1817);
nand U2500 (N_2500,N_1578,N_1225);
or U2501 (N_2501,N_1978,N_1349);
nor U2502 (N_2502,N_1598,N_1398);
nand U2503 (N_2503,N_1898,N_1272);
and U2504 (N_2504,N_1027,N_1335);
nand U2505 (N_2505,N_1993,N_1738);
nor U2506 (N_2506,N_1266,N_1036);
nand U2507 (N_2507,N_1101,N_1750);
and U2508 (N_2508,N_1034,N_1104);
nor U2509 (N_2509,N_1246,N_1460);
nor U2510 (N_2510,N_1184,N_1177);
or U2511 (N_2511,N_1808,N_1732);
or U2512 (N_2512,N_1397,N_1750);
or U2513 (N_2513,N_1163,N_1711);
nand U2514 (N_2514,N_1742,N_1250);
nand U2515 (N_2515,N_1864,N_1334);
nand U2516 (N_2516,N_1774,N_1808);
and U2517 (N_2517,N_1524,N_1518);
and U2518 (N_2518,N_1806,N_1180);
nand U2519 (N_2519,N_1710,N_1017);
nor U2520 (N_2520,N_1917,N_1330);
nor U2521 (N_2521,N_1484,N_1016);
and U2522 (N_2522,N_1691,N_1996);
and U2523 (N_2523,N_1508,N_1291);
nor U2524 (N_2524,N_1309,N_1567);
nand U2525 (N_2525,N_1049,N_1726);
or U2526 (N_2526,N_1773,N_1821);
nand U2527 (N_2527,N_1029,N_1817);
nand U2528 (N_2528,N_1267,N_1705);
and U2529 (N_2529,N_1245,N_1831);
nor U2530 (N_2530,N_1845,N_1062);
nor U2531 (N_2531,N_1290,N_1002);
and U2532 (N_2532,N_1569,N_1313);
nor U2533 (N_2533,N_1157,N_1101);
nor U2534 (N_2534,N_1231,N_1150);
nor U2535 (N_2535,N_1825,N_1765);
and U2536 (N_2536,N_1606,N_1976);
or U2537 (N_2537,N_1288,N_1159);
or U2538 (N_2538,N_1073,N_1659);
or U2539 (N_2539,N_1803,N_1027);
and U2540 (N_2540,N_1270,N_1040);
nand U2541 (N_2541,N_1614,N_1041);
xnor U2542 (N_2542,N_1664,N_1008);
nor U2543 (N_2543,N_1633,N_1001);
or U2544 (N_2544,N_1651,N_1456);
nand U2545 (N_2545,N_1230,N_1963);
nor U2546 (N_2546,N_1911,N_1607);
nor U2547 (N_2547,N_1172,N_1680);
and U2548 (N_2548,N_1517,N_1346);
nor U2549 (N_2549,N_1577,N_1551);
or U2550 (N_2550,N_1658,N_1670);
and U2551 (N_2551,N_1052,N_1298);
nand U2552 (N_2552,N_1707,N_1748);
or U2553 (N_2553,N_1463,N_1460);
nand U2554 (N_2554,N_1285,N_1518);
or U2555 (N_2555,N_1636,N_1906);
nor U2556 (N_2556,N_1449,N_1104);
nand U2557 (N_2557,N_1085,N_1230);
nand U2558 (N_2558,N_1767,N_1733);
or U2559 (N_2559,N_1137,N_1983);
nor U2560 (N_2560,N_1142,N_1466);
and U2561 (N_2561,N_1403,N_1774);
or U2562 (N_2562,N_1687,N_1519);
or U2563 (N_2563,N_1303,N_1778);
or U2564 (N_2564,N_1016,N_1960);
xor U2565 (N_2565,N_1681,N_1493);
or U2566 (N_2566,N_1903,N_1179);
nor U2567 (N_2567,N_1662,N_1802);
nor U2568 (N_2568,N_1646,N_1342);
nor U2569 (N_2569,N_1172,N_1242);
nor U2570 (N_2570,N_1896,N_1724);
nand U2571 (N_2571,N_1176,N_1456);
nand U2572 (N_2572,N_1779,N_1098);
nand U2573 (N_2573,N_1464,N_1969);
or U2574 (N_2574,N_1373,N_1242);
nand U2575 (N_2575,N_1173,N_1262);
and U2576 (N_2576,N_1342,N_1796);
nor U2577 (N_2577,N_1143,N_1261);
and U2578 (N_2578,N_1006,N_1024);
nand U2579 (N_2579,N_1132,N_1274);
or U2580 (N_2580,N_1800,N_1556);
nand U2581 (N_2581,N_1702,N_1030);
nand U2582 (N_2582,N_1502,N_1529);
and U2583 (N_2583,N_1701,N_1686);
nand U2584 (N_2584,N_1133,N_1337);
or U2585 (N_2585,N_1698,N_1588);
nor U2586 (N_2586,N_1142,N_1738);
nor U2587 (N_2587,N_1578,N_1895);
or U2588 (N_2588,N_1767,N_1446);
and U2589 (N_2589,N_1328,N_1024);
xor U2590 (N_2590,N_1781,N_1232);
nor U2591 (N_2591,N_1908,N_1564);
xor U2592 (N_2592,N_1853,N_1746);
xor U2593 (N_2593,N_1272,N_1337);
and U2594 (N_2594,N_1708,N_1139);
nor U2595 (N_2595,N_1374,N_1415);
nand U2596 (N_2596,N_1087,N_1111);
nor U2597 (N_2597,N_1783,N_1317);
nand U2598 (N_2598,N_1156,N_1426);
nand U2599 (N_2599,N_1374,N_1617);
nand U2600 (N_2600,N_1601,N_1768);
and U2601 (N_2601,N_1607,N_1815);
and U2602 (N_2602,N_1615,N_1819);
or U2603 (N_2603,N_1274,N_1903);
nand U2604 (N_2604,N_1027,N_1891);
nor U2605 (N_2605,N_1395,N_1760);
or U2606 (N_2606,N_1239,N_1553);
and U2607 (N_2607,N_1627,N_1484);
nor U2608 (N_2608,N_1737,N_1305);
nand U2609 (N_2609,N_1937,N_1228);
nor U2610 (N_2610,N_1625,N_1159);
or U2611 (N_2611,N_1843,N_1880);
nor U2612 (N_2612,N_1521,N_1225);
xor U2613 (N_2613,N_1686,N_1681);
nor U2614 (N_2614,N_1061,N_1618);
and U2615 (N_2615,N_1212,N_1766);
and U2616 (N_2616,N_1783,N_1759);
nand U2617 (N_2617,N_1182,N_1804);
nor U2618 (N_2618,N_1980,N_1728);
or U2619 (N_2619,N_1440,N_1410);
nand U2620 (N_2620,N_1611,N_1151);
and U2621 (N_2621,N_1850,N_1658);
or U2622 (N_2622,N_1848,N_1456);
or U2623 (N_2623,N_1190,N_1031);
or U2624 (N_2624,N_1626,N_1869);
nor U2625 (N_2625,N_1208,N_1995);
or U2626 (N_2626,N_1058,N_1113);
nor U2627 (N_2627,N_1276,N_1082);
or U2628 (N_2628,N_1545,N_1797);
nor U2629 (N_2629,N_1893,N_1090);
or U2630 (N_2630,N_1493,N_1834);
xor U2631 (N_2631,N_1370,N_1445);
or U2632 (N_2632,N_1530,N_1104);
nand U2633 (N_2633,N_1920,N_1015);
nand U2634 (N_2634,N_1315,N_1958);
nor U2635 (N_2635,N_1565,N_1201);
or U2636 (N_2636,N_1127,N_1627);
or U2637 (N_2637,N_1476,N_1432);
nand U2638 (N_2638,N_1577,N_1985);
nand U2639 (N_2639,N_1434,N_1075);
or U2640 (N_2640,N_1568,N_1435);
nand U2641 (N_2641,N_1869,N_1842);
nand U2642 (N_2642,N_1767,N_1615);
or U2643 (N_2643,N_1560,N_1148);
or U2644 (N_2644,N_1737,N_1772);
nand U2645 (N_2645,N_1360,N_1744);
nand U2646 (N_2646,N_1157,N_1819);
nor U2647 (N_2647,N_1518,N_1521);
xor U2648 (N_2648,N_1225,N_1758);
or U2649 (N_2649,N_1385,N_1287);
or U2650 (N_2650,N_1627,N_1008);
or U2651 (N_2651,N_1815,N_1155);
and U2652 (N_2652,N_1353,N_1099);
or U2653 (N_2653,N_1388,N_1883);
and U2654 (N_2654,N_1600,N_1647);
nand U2655 (N_2655,N_1210,N_1603);
nor U2656 (N_2656,N_1439,N_1427);
nor U2657 (N_2657,N_1677,N_1705);
or U2658 (N_2658,N_1808,N_1270);
and U2659 (N_2659,N_1126,N_1458);
nor U2660 (N_2660,N_1389,N_1759);
or U2661 (N_2661,N_1387,N_1960);
nor U2662 (N_2662,N_1890,N_1321);
nor U2663 (N_2663,N_1562,N_1711);
or U2664 (N_2664,N_1612,N_1994);
or U2665 (N_2665,N_1295,N_1066);
and U2666 (N_2666,N_1087,N_1179);
nor U2667 (N_2667,N_1467,N_1955);
nor U2668 (N_2668,N_1022,N_1891);
and U2669 (N_2669,N_1539,N_1511);
or U2670 (N_2670,N_1546,N_1885);
nor U2671 (N_2671,N_1712,N_1460);
and U2672 (N_2672,N_1170,N_1800);
and U2673 (N_2673,N_1055,N_1442);
and U2674 (N_2674,N_1072,N_1911);
or U2675 (N_2675,N_1198,N_1015);
or U2676 (N_2676,N_1567,N_1029);
nand U2677 (N_2677,N_1174,N_1912);
nor U2678 (N_2678,N_1673,N_1641);
nor U2679 (N_2679,N_1130,N_1646);
and U2680 (N_2680,N_1582,N_1026);
and U2681 (N_2681,N_1628,N_1915);
nor U2682 (N_2682,N_1717,N_1769);
and U2683 (N_2683,N_1154,N_1112);
and U2684 (N_2684,N_1716,N_1474);
nor U2685 (N_2685,N_1521,N_1404);
or U2686 (N_2686,N_1011,N_1440);
or U2687 (N_2687,N_1941,N_1921);
nand U2688 (N_2688,N_1833,N_1403);
or U2689 (N_2689,N_1411,N_1753);
and U2690 (N_2690,N_1772,N_1363);
nor U2691 (N_2691,N_1146,N_1027);
nor U2692 (N_2692,N_1205,N_1250);
nor U2693 (N_2693,N_1114,N_1567);
and U2694 (N_2694,N_1855,N_1295);
and U2695 (N_2695,N_1008,N_1066);
nor U2696 (N_2696,N_1555,N_1187);
nor U2697 (N_2697,N_1438,N_1809);
nor U2698 (N_2698,N_1523,N_1408);
or U2699 (N_2699,N_1922,N_1201);
nor U2700 (N_2700,N_1782,N_1740);
or U2701 (N_2701,N_1510,N_1095);
nor U2702 (N_2702,N_1661,N_1834);
nand U2703 (N_2703,N_1829,N_1045);
nand U2704 (N_2704,N_1096,N_1181);
nor U2705 (N_2705,N_1524,N_1647);
or U2706 (N_2706,N_1220,N_1735);
nand U2707 (N_2707,N_1477,N_1363);
nand U2708 (N_2708,N_1096,N_1143);
or U2709 (N_2709,N_1806,N_1027);
and U2710 (N_2710,N_1055,N_1859);
nor U2711 (N_2711,N_1048,N_1938);
nor U2712 (N_2712,N_1930,N_1618);
nand U2713 (N_2713,N_1569,N_1761);
or U2714 (N_2714,N_1208,N_1794);
and U2715 (N_2715,N_1354,N_1122);
and U2716 (N_2716,N_1882,N_1675);
nor U2717 (N_2717,N_1665,N_1757);
nor U2718 (N_2718,N_1434,N_1467);
or U2719 (N_2719,N_1708,N_1244);
nand U2720 (N_2720,N_1596,N_1011);
nor U2721 (N_2721,N_1452,N_1516);
or U2722 (N_2722,N_1047,N_1945);
or U2723 (N_2723,N_1935,N_1707);
or U2724 (N_2724,N_1380,N_1327);
or U2725 (N_2725,N_1559,N_1295);
and U2726 (N_2726,N_1436,N_1756);
or U2727 (N_2727,N_1000,N_1174);
nand U2728 (N_2728,N_1178,N_1417);
nand U2729 (N_2729,N_1109,N_1883);
or U2730 (N_2730,N_1751,N_1869);
nor U2731 (N_2731,N_1741,N_1447);
and U2732 (N_2732,N_1055,N_1606);
nand U2733 (N_2733,N_1125,N_1971);
nand U2734 (N_2734,N_1836,N_1594);
or U2735 (N_2735,N_1700,N_1663);
nor U2736 (N_2736,N_1143,N_1486);
nor U2737 (N_2737,N_1635,N_1110);
or U2738 (N_2738,N_1995,N_1090);
or U2739 (N_2739,N_1220,N_1681);
or U2740 (N_2740,N_1762,N_1255);
or U2741 (N_2741,N_1417,N_1583);
nor U2742 (N_2742,N_1559,N_1681);
and U2743 (N_2743,N_1585,N_1088);
nand U2744 (N_2744,N_1978,N_1890);
nand U2745 (N_2745,N_1185,N_1109);
or U2746 (N_2746,N_1452,N_1759);
and U2747 (N_2747,N_1443,N_1662);
and U2748 (N_2748,N_1676,N_1076);
or U2749 (N_2749,N_1858,N_1115);
and U2750 (N_2750,N_1312,N_1418);
nand U2751 (N_2751,N_1623,N_1343);
nand U2752 (N_2752,N_1117,N_1302);
nand U2753 (N_2753,N_1712,N_1035);
and U2754 (N_2754,N_1006,N_1409);
and U2755 (N_2755,N_1330,N_1293);
or U2756 (N_2756,N_1495,N_1681);
and U2757 (N_2757,N_1914,N_1873);
nor U2758 (N_2758,N_1602,N_1005);
or U2759 (N_2759,N_1989,N_1544);
or U2760 (N_2760,N_1524,N_1517);
or U2761 (N_2761,N_1747,N_1807);
nor U2762 (N_2762,N_1497,N_1267);
nor U2763 (N_2763,N_1783,N_1260);
and U2764 (N_2764,N_1221,N_1805);
nand U2765 (N_2765,N_1914,N_1468);
nor U2766 (N_2766,N_1177,N_1941);
nand U2767 (N_2767,N_1110,N_1764);
and U2768 (N_2768,N_1431,N_1958);
or U2769 (N_2769,N_1906,N_1519);
nor U2770 (N_2770,N_1657,N_1709);
nand U2771 (N_2771,N_1500,N_1820);
nand U2772 (N_2772,N_1522,N_1447);
or U2773 (N_2773,N_1588,N_1188);
nor U2774 (N_2774,N_1092,N_1058);
nor U2775 (N_2775,N_1848,N_1730);
and U2776 (N_2776,N_1414,N_1989);
nor U2777 (N_2777,N_1119,N_1749);
nor U2778 (N_2778,N_1653,N_1242);
and U2779 (N_2779,N_1102,N_1022);
nor U2780 (N_2780,N_1378,N_1640);
nand U2781 (N_2781,N_1645,N_1352);
and U2782 (N_2782,N_1567,N_1279);
nand U2783 (N_2783,N_1902,N_1357);
or U2784 (N_2784,N_1327,N_1565);
nand U2785 (N_2785,N_1875,N_1741);
nand U2786 (N_2786,N_1688,N_1060);
nand U2787 (N_2787,N_1182,N_1328);
nor U2788 (N_2788,N_1954,N_1660);
xnor U2789 (N_2789,N_1531,N_1088);
nor U2790 (N_2790,N_1112,N_1855);
or U2791 (N_2791,N_1665,N_1451);
nand U2792 (N_2792,N_1925,N_1592);
nand U2793 (N_2793,N_1280,N_1717);
nand U2794 (N_2794,N_1195,N_1786);
nor U2795 (N_2795,N_1820,N_1236);
and U2796 (N_2796,N_1325,N_1331);
nor U2797 (N_2797,N_1153,N_1044);
or U2798 (N_2798,N_1063,N_1901);
nor U2799 (N_2799,N_1286,N_1049);
nor U2800 (N_2800,N_1991,N_1557);
or U2801 (N_2801,N_1073,N_1593);
nor U2802 (N_2802,N_1333,N_1947);
nand U2803 (N_2803,N_1780,N_1038);
or U2804 (N_2804,N_1095,N_1961);
and U2805 (N_2805,N_1935,N_1533);
or U2806 (N_2806,N_1593,N_1610);
nand U2807 (N_2807,N_1021,N_1491);
or U2808 (N_2808,N_1164,N_1957);
or U2809 (N_2809,N_1378,N_1481);
nor U2810 (N_2810,N_1939,N_1213);
or U2811 (N_2811,N_1359,N_1469);
or U2812 (N_2812,N_1236,N_1149);
nand U2813 (N_2813,N_1520,N_1791);
or U2814 (N_2814,N_1221,N_1165);
xor U2815 (N_2815,N_1913,N_1956);
or U2816 (N_2816,N_1720,N_1571);
xnor U2817 (N_2817,N_1838,N_1233);
and U2818 (N_2818,N_1012,N_1493);
or U2819 (N_2819,N_1315,N_1093);
or U2820 (N_2820,N_1951,N_1144);
nand U2821 (N_2821,N_1691,N_1962);
nand U2822 (N_2822,N_1570,N_1003);
nor U2823 (N_2823,N_1394,N_1817);
nand U2824 (N_2824,N_1289,N_1859);
or U2825 (N_2825,N_1615,N_1115);
or U2826 (N_2826,N_1866,N_1617);
or U2827 (N_2827,N_1991,N_1312);
nand U2828 (N_2828,N_1043,N_1482);
nor U2829 (N_2829,N_1673,N_1896);
or U2830 (N_2830,N_1791,N_1556);
nand U2831 (N_2831,N_1292,N_1843);
nand U2832 (N_2832,N_1362,N_1398);
and U2833 (N_2833,N_1466,N_1712);
nand U2834 (N_2834,N_1596,N_1660);
nand U2835 (N_2835,N_1692,N_1216);
nor U2836 (N_2836,N_1942,N_1401);
nand U2837 (N_2837,N_1494,N_1644);
nor U2838 (N_2838,N_1230,N_1742);
nand U2839 (N_2839,N_1299,N_1902);
nand U2840 (N_2840,N_1114,N_1364);
nor U2841 (N_2841,N_1308,N_1364);
nand U2842 (N_2842,N_1349,N_1114);
nand U2843 (N_2843,N_1317,N_1327);
nand U2844 (N_2844,N_1480,N_1155);
and U2845 (N_2845,N_1312,N_1355);
nand U2846 (N_2846,N_1368,N_1228);
nand U2847 (N_2847,N_1436,N_1458);
nand U2848 (N_2848,N_1198,N_1551);
nand U2849 (N_2849,N_1267,N_1481);
nand U2850 (N_2850,N_1537,N_1945);
and U2851 (N_2851,N_1045,N_1738);
or U2852 (N_2852,N_1526,N_1436);
or U2853 (N_2853,N_1154,N_1601);
and U2854 (N_2854,N_1886,N_1719);
xnor U2855 (N_2855,N_1436,N_1336);
nand U2856 (N_2856,N_1547,N_1191);
and U2857 (N_2857,N_1967,N_1504);
nor U2858 (N_2858,N_1310,N_1363);
xnor U2859 (N_2859,N_1284,N_1472);
or U2860 (N_2860,N_1202,N_1963);
or U2861 (N_2861,N_1311,N_1246);
and U2862 (N_2862,N_1604,N_1152);
or U2863 (N_2863,N_1389,N_1833);
nor U2864 (N_2864,N_1373,N_1200);
xnor U2865 (N_2865,N_1722,N_1715);
or U2866 (N_2866,N_1391,N_1029);
and U2867 (N_2867,N_1098,N_1706);
or U2868 (N_2868,N_1259,N_1966);
or U2869 (N_2869,N_1206,N_1612);
and U2870 (N_2870,N_1124,N_1998);
and U2871 (N_2871,N_1713,N_1642);
nand U2872 (N_2872,N_1962,N_1394);
nand U2873 (N_2873,N_1278,N_1850);
xor U2874 (N_2874,N_1371,N_1339);
nand U2875 (N_2875,N_1176,N_1174);
and U2876 (N_2876,N_1462,N_1700);
nor U2877 (N_2877,N_1210,N_1402);
or U2878 (N_2878,N_1688,N_1232);
nor U2879 (N_2879,N_1918,N_1104);
and U2880 (N_2880,N_1104,N_1226);
or U2881 (N_2881,N_1346,N_1955);
and U2882 (N_2882,N_1259,N_1328);
and U2883 (N_2883,N_1229,N_1895);
nand U2884 (N_2884,N_1226,N_1220);
or U2885 (N_2885,N_1824,N_1370);
nand U2886 (N_2886,N_1681,N_1589);
nand U2887 (N_2887,N_1106,N_1144);
and U2888 (N_2888,N_1439,N_1534);
nand U2889 (N_2889,N_1781,N_1649);
nor U2890 (N_2890,N_1934,N_1541);
and U2891 (N_2891,N_1991,N_1922);
nor U2892 (N_2892,N_1421,N_1934);
or U2893 (N_2893,N_1409,N_1227);
nor U2894 (N_2894,N_1435,N_1060);
or U2895 (N_2895,N_1165,N_1525);
or U2896 (N_2896,N_1610,N_1633);
and U2897 (N_2897,N_1687,N_1660);
and U2898 (N_2898,N_1791,N_1349);
nand U2899 (N_2899,N_1104,N_1125);
nand U2900 (N_2900,N_1820,N_1610);
and U2901 (N_2901,N_1546,N_1048);
nor U2902 (N_2902,N_1446,N_1591);
nand U2903 (N_2903,N_1058,N_1662);
nand U2904 (N_2904,N_1299,N_1681);
nand U2905 (N_2905,N_1473,N_1250);
nand U2906 (N_2906,N_1039,N_1060);
and U2907 (N_2907,N_1554,N_1710);
nand U2908 (N_2908,N_1287,N_1513);
and U2909 (N_2909,N_1452,N_1830);
nor U2910 (N_2910,N_1468,N_1345);
nor U2911 (N_2911,N_1686,N_1867);
or U2912 (N_2912,N_1008,N_1721);
nor U2913 (N_2913,N_1429,N_1109);
nand U2914 (N_2914,N_1305,N_1070);
nand U2915 (N_2915,N_1433,N_1948);
or U2916 (N_2916,N_1358,N_1868);
or U2917 (N_2917,N_1045,N_1826);
and U2918 (N_2918,N_1015,N_1880);
nand U2919 (N_2919,N_1703,N_1606);
or U2920 (N_2920,N_1438,N_1284);
or U2921 (N_2921,N_1702,N_1048);
nor U2922 (N_2922,N_1587,N_1726);
nand U2923 (N_2923,N_1699,N_1150);
nand U2924 (N_2924,N_1084,N_1537);
or U2925 (N_2925,N_1060,N_1272);
nand U2926 (N_2926,N_1365,N_1682);
nor U2927 (N_2927,N_1997,N_1055);
and U2928 (N_2928,N_1234,N_1805);
and U2929 (N_2929,N_1570,N_1381);
or U2930 (N_2930,N_1622,N_1384);
or U2931 (N_2931,N_1260,N_1312);
nor U2932 (N_2932,N_1046,N_1787);
nand U2933 (N_2933,N_1634,N_1149);
or U2934 (N_2934,N_1012,N_1936);
and U2935 (N_2935,N_1770,N_1727);
nand U2936 (N_2936,N_1710,N_1488);
or U2937 (N_2937,N_1656,N_1337);
and U2938 (N_2938,N_1434,N_1229);
xor U2939 (N_2939,N_1604,N_1878);
or U2940 (N_2940,N_1674,N_1526);
or U2941 (N_2941,N_1882,N_1989);
nor U2942 (N_2942,N_1517,N_1641);
nor U2943 (N_2943,N_1342,N_1597);
nand U2944 (N_2944,N_1604,N_1705);
or U2945 (N_2945,N_1468,N_1991);
and U2946 (N_2946,N_1925,N_1494);
nand U2947 (N_2947,N_1624,N_1837);
or U2948 (N_2948,N_1285,N_1909);
and U2949 (N_2949,N_1576,N_1384);
nand U2950 (N_2950,N_1720,N_1870);
nor U2951 (N_2951,N_1330,N_1312);
nor U2952 (N_2952,N_1818,N_1340);
nand U2953 (N_2953,N_1856,N_1301);
nand U2954 (N_2954,N_1242,N_1659);
nand U2955 (N_2955,N_1573,N_1946);
and U2956 (N_2956,N_1631,N_1883);
and U2957 (N_2957,N_1409,N_1631);
nor U2958 (N_2958,N_1164,N_1786);
or U2959 (N_2959,N_1322,N_1572);
xnor U2960 (N_2960,N_1678,N_1734);
nor U2961 (N_2961,N_1476,N_1912);
nor U2962 (N_2962,N_1454,N_1291);
nand U2963 (N_2963,N_1826,N_1368);
or U2964 (N_2964,N_1826,N_1800);
and U2965 (N_2965,N_1974,N_1574);
or U2966 (N_2966,N_1261,N_1607);
or U2967 (N_2967,N_1976,N_1523);
nand U2968 (N_2968,N_1604,N_1835);
or U2969 (N_2969,N_1216,N_1568);
nor U2970 (N_2970,N_1812,N_1065);
or U2971 (N_2971,N_1925,N_1766);
and U2972 (N_2972,N_1629,N_1795);
and U2973 (N_2973,N_1529,N_1864);
nor U2974 (N_2974,N_1502,N_1617);
and U2975 (N_2975,N_1692,N_1412);
and U2976 (N_2976,N_1510,N_1767);
nor U2977 (N_2977,N_1998,N_1354);
nor U2978 (N_2978,N_1523,N_1036);
and U2979 (N_2979,N_1471,N_1493);
or U2980 (N_2980,N_1401,N_1509);
nor U2981 (N_2981,N_1913,N_1808);
or U2982 (N_2982,N_1201,N_1443);
xor U2983 (N_2983,N_1081,N_1394);
and U2984 (N_2984,N_1167,N_1579);
nand U2985 (N_2985,N_1223,N_1171);
xnor U2986 (N_2986,N_1909,N_1969);
and U2987 (N_2987,N_1901,N_1954);
and U2988 (N_2988,N_1458,N_1544);
or U2989 (N_2989,N_1141,N_1058);
and U2990 (N_2990,N_1213,N_1886);
nor U2991 (N_2991,N_1862,N_1422);
and U2992 (N_2992,N_1093,N_1844);
or U2993 (N_2993,N_1261,N_1827);
or U2994 (N_2994,N_1619,N_1386);
xnor U2995 (N_2995,N_1008,N_1700);
and U2996 (N_2996,N_1065,N_1197);
or U2997 (N_2997,N_1311,N_1815);
nand U2998 (N_2998,N_1241,N_1622);
and U2999 (N_2999,N_1272,N_1650);
nor U3000 (N_3000,N_2927,N_2665);
xnor U3001 (N_3001,N_2422,N_2751);
or U3002 (N_3002,N_2877,N_2532);
or U3003 (N_3003,N_2447,N_2712);
xor U3004 (N_3004,N_2896,N_2918);
nand U3005 (N_3005,N_2948,N_2146);
nor U3006 (N_3006,N_2546,N_2084);
and U3007 (N_3007,N_2080,N_2800);
nand U3008 (N_3008,N_2108,N_2318);
nor U3009 (N_3009,N_2079,N_2273);
or U3010 (N_3010,N_2162,N_2207);
or U3011 (N_3011,N_2405,N_2563);
and U3012 (N_3012,N_2886,N_2304);
nand U3013 (N_3013,N_2820,N_2005);
and U3014 (N_3014,N_2627,N_2115);
or U3015 (N_3015,N_2061,N_2917);
nand U3016 (N_3016,N_2314,N_2349);
or U3017 (N_3017,N_2694,N_2029);
nor U3018 (N_3018,N_2122,N_2338);
nand U3019 (N_3019,N_2899,N_2865);
nand U3020 (N_3020,N_2515,N_2517);
nor U3021 (N_3021,N_2726,N_2850);
nand U3022 (N_3022,N_2325,N_2017);
nand U3023 (N_3023,N_2804,N_2764);
nor U3024 (N_3024,N_2600,N_2097);
nand U3025 (N_3025,N_2553,N_2842);
nor U3026 (N_3026,N_2872,N_2632);
nand U3027 (N_3027,N_2169,N_2659);
and U3028 (N_3028,N_2026,N_2720);
nand U3029 (N_3029,N_2759,N_2147);
and U3030 (N_3030,N_2004,N_2956);
or U3031 (N_3031,N_2824,N_2721);
nor U3032 (N_3032,N_2643,N_2934);
and U3033 (N_3033,N_2062,N_2581);
nand U3034 (N_3034,N_2569,N_2438);
nor U3035 (N_3035,N_2460,N_2173);
xnor U3036 (N_3036,N_2662,N_2033);
and U3037 (N_3037,N_2675,N_2595);
nand U3038 (N_3038,N_2398,N_2365);
and U3039 (N_3039,N_2091,N_2280);
nand U3040 (N_3040,N_2845,N_2477);
and U3041 (N_3041,N_2100,N_2673);
nor U3042 (N_3042,N_2219,N_2233);
xnor U3043 (N_3043,N_2691,N_2040);
nor U3044 (N_3044,N_2582,N_2035);
nand U3045 (N_3045,N_2578,N_2819);
nand U3046 (N_3046,N_2024,N_2735);
and U3047 (N_3047,N_2323,N_2959);
nor U3048 (N_3048,N_2602,N_2401);
and U3049 (N_3049,N_2473,N_2944);
nand U3050 (N_3050,N_2381,N_2901);
nand U3051 (N_3051,N_2980,N_2468);
nor U3052 (N_3052,N_2536,N_2808);
or U3053 (N_3053,N_2623,N_2277);
nor U3054 (N_3054,N_2175,N_2640);
and U3055 (N_3055,N_2109,N_2199);
nand U3056 (N_3056,N_2107,N_2612);
and U3057 (N_3057,N_2394,N_2737);
or U3058 (N_3058,N_2063,N_2526);
nand U3059 (N_3059,N_2562,N_2121);
or U3060 (N_3060,N_2119,N_2060);
nand U3061 (N_3061,N_2204,N_2789);
xnor U3062 (N_3062,N_2476,N_2603);
or U3063 (N_3063,N_2150,N_2670);
xnor U3064 (N_3064,N_2876,N_2149);
or U3065 (N_3065,N_2625,N_2963);
or U3066 (N_3066,N_2888,N_2651);
and U3067 (N_3067,N_2009,N_2893);
nor U3068 (N_3068,N_2818,N_2940);
nand U3069 (N_3069,N_2458,N_2406);
nand U3070 (N_3070,N_2211,N_2125);
or U3071 (N_3071,N_2978,N_2561);
nand U3072 (N_3072,N_2027,N_2259);
nor U3073 (N_3073,N_2585,N_2501);
and U3074 (N_3074,N_2250,N_2282);
or U3075 (N_3075,N_2565,N_2191);
or U3076 (N_3076,N_2500,N_2567);
or U3077 (N_3077,N_2400,N_2674);
and U3078 (N_3078,N_2984,N_2853);
and U3079 (N_3079,N_2439,N_2622);
nand U3080 (N_3080,N_2426,N_2195);
nor U3081 (N_3081,N_2791,N_2159);
nand U3082 (N_3082,N_2520,N_2237);
nor U3083 (N_3083,N_2152,N_2472);
nor U3084 (N_3084,N_2895,N_2758);
and U3085 (N_3085,N_2849,N_2385);
or U3086 (N_3086,N_2444,N_2114);
xor U3087 (N_3087,N_2188,N_2315);
nor U3088 (N_3088,N_2573,N_2559);
nand U3089 (N_3089,N_2189,N_2930);
nor U3090 (N_3090,N_2187,N_2792);
or U3091 (N_3091,N_2781,N_2794);
nor U3092 (N_3092,N_2018,N_2424);
or U3093 (N_3093,N_2652,N_2692);
nand U3094 (N_3094,N_2656,N_2760);
nand U3095 (N_3095,N_2240,N_2540);
nand U3096 (N_3096,N_2265,N_2176);
and U3097 (N_3097,N_2958,N_2545);
xnor U3098 (N_3098,N_2441,N_2373);
nor U3099 (N_3099,N_2293,N_2783);
or U3100 (N_3100,N_2952,N_2671);
nand U3101 (N_3101,N_2619,N_2345);
nand U3102 (N_3102,N_2482,N_2977);
or U3103 (N_3103,N_2010,N_2423);
nand U3104 (N_3104,N_2587,N_2555);
nor U3105 (N_3105,N_2890,N_2833);
or U3106 (N_3106,N_2341,N_2511);
nor U3107 (N_3107,N_2052,N_2283);
nor U3108 (N_3108,N_2081,N_2658);
and U3109 (N_3109,N_2596,N_2795);
or U3110 (N_3110,N_2230,N_2856);
nor U3111 (N_3111,N_2408,N_2007);
and U3112 (N_3112,N_2298,N_2731);
nor U3113 (N_3113,N_2593,N_2928);
or U3114 (N_3114,N_2547,N_2364);
nand U3115 (N_3115,N_2861,N_2413);
nand U3116 (N_3116,N_2252,N_2055);
and U3117 (N_3117,N_2586,N_2975);
nand U3118 (N_3118,N_2769,N_2317);
nor U3119 (N_3119,N_2755,N_2809);
or U3120 (N_3120,N_2701,N_2677);
nor U3121 (N_3121,N_2069,N_2261);
or U3122 (N_3122,N_2267,N_2331);
and U3123 (N_3123,N_2418,N_2234);
nand U3124 (N_3124,N_2799,N_2183);
or U3125 (N_3125,N_2527,N_2370);
nand U3126 (N_3126,N_2908,N_2151);
xor U3127 (N_3127,N_2772,N_2648);
nand U3128 (N_3128,N_2947,N_2128);
nand U3129 (N_3129,N_2059,N_2112);
and U3130 (N_3130,N_2208,N_2368);
nand U3131 (N_3131,N_2480,N_2232);
nand U3132 (N_3132,N_2556,N_2613);
and U3133 (N_3133,N_2636,N_2218);
xnor U3134 (N_3134,N_2324,N_2165);
nor U3135 (N_3135,N_2919,N_2431);
or U3136 (N_3136,N_2181,N_2481);
nor U3137 (N_3137,N_2038,N_2154);
nand U3138 (N_3138,N_2634,N_2668);
or U3139 (N_3139,N_2488,N_2521);
xor U3140 (N_3140,N_2493,N_2678);
and U3141 (N_3141,N_2570,N_2744);
and U3142 (N_3142,N_2649,N_2163);
and U3143 (N_3143,N_2516,N_2666);
and U3144 (N_3144,N_2369,N_2443);
nand U3145 (N_3145,N_2885,N_2492);
nand U3146 (N_3146,N_2319,N_2736);
and U3147 (N_3147,N_2343,N_2839);
nor U3148 (N_3148,N_2860,N_2358);
or U3149 (N_3149,N_2387,N_2311);
or U3150 (N_3150,N_2136,N_2822);
nor U3151 (N_3151,N_2337,N_2415);
nor U3152 (N_3152,N_2044,N_2339);
or U3153 (N_3153,N_2479,N_2523);
nand U3154 (N_3154,N_2435,N_2372);
and U3155 (N_3155,N_2272,N_2457);
and U3156 (N_3156,N_2243,N_2245);
nand U3157 (N_3157,N_2498,N_2275);
or U3158 (N_3158,N_2157,N_2747);
nand U3159 (N_3159,N_2085,N_2912);
and U3160 (N_3160,N_2786,N_2306);
nand U3161 (N_3161,N_2777,N_2655);
nor U3162 (N_3162,N_2143,N_2420);
and U3163 (N_3163,N_2212,N_2548);
or U3164 (N_3164,N_2192,N_2834);
and U3165 (N_3165,N_2766,N_2838);
nand U3166 (N_3166,N_2994,N_2524);
and U3167 (N_3167,N_2813,N_2057);
and U3168 (N_3168,N_2979,N_2981);
and U3169 (N_3169,N_2003,N_2268);
and U3170 (N_3170,N_2032,N_2653);
nor U3171 (N_3171,N_2502,N_2434);
nand U3172 (N_3172,N_2762,N_2993);
nor U3173 (N_3173,N_2048,N_2088);
nand U3174 (N_3174,N_2106,N_2437);
or U3175 (N_3175,N_2637,N_2359);
and U3176 (N_3176,N_2043,N_2560);
and U3177 (N_3177,N_2130,N_2104);
and U3178 (N_3178,N_2054,N_2904);
or U3179 (N_3179,N_2356,N_2870);
or U3180 (N_3180,N_2598,N_2973);
and U3181 (N_3181,N_2278,N_2740);
nor U3182 (N_3182,N_2328,N_2411);
nand U3183 (N_3183,N_2310,N_2951);
or U3184 (N_3184,N_2654,N_2168);
nor U3185 (N_3185,N_2857,N_2214);
or U3186 (N_3186,N_2894,N_2663);
nand U3187 (N_3187,N_2787,N_2138);
nor U3188 (N_3188,N_2463,N_2594);
and U3189 (N_3189,N_2021,N_2153);
nand U3190 (N_3190,N_2983,N_2825);
nand U3191 (N_3191,N_2164,N_2148);
and U3192 (N_3192,N_2262,N_2361);
and U3193 (N_3193,N_2402,N_2134);
nor U3194 (N_3194,N_2638,N_2390);
nand U3195 (N_3195,N_2068,N_2236);
nand U3196 (N_3196,N_2699,N_2051);
xor U3197 (N_3197,N_2704,N_2986);
nand U3198 (N_3198,N_2946,N_2353);
nand U3199 (N_3199,N_2116,N_2913);
or U3200 (N_3200,N_2806,N_2377);
or U3201 (N_3201,N_2635,N_2810);
or U3202 (N_3202,N_2182,N_2681);
nor U3203 (N_3203,N_2185,N_2626);
nor U3204 (N_3204,N_2248,N_2803);
or U3205 (N_3205,N_2030,N_2728);
or U3206 (N_3206,N_2417,N_2333);
nor U3207 (N_3207,N_2875,N_2644);
or U3208 (N_3208,N_2891,N_2924);
and U3209 (N_3209,N_2916,N_2225);
or U3210 (N_3210,N_2290,N_2628);
or U3211 (N_3211,N_2879,N_2525);
and U3212 (N_3212,N_2244,N_2831);
and U3213 (N_3213,N_2892,N_2193);
xor U3214 (N_3214,N_2601,N_2882);
and U3215 (N_3215,N_2969,N_2773);
nor U3216 (N_3216,N_2025,N_2884);
or U3217 (N_3217,N_2748,N_2949);
nand U3218 (N_3218,N_2036,N_2095);
and U3219 (N_3219,N_2579,N_2445);
nor U3220 (N_3220,N_2887,N_2485);
nand U3221 (N_3221,N_2935,N_2826);
nor U3222 (N_3222,N_2023,N_2451);
or U3223 (N_3223,N_2931,N_2287);
xnor U3224 (N_3224,N_2780,N_2862);
nor U3225 (N_3225,N_2906,N_2231);
nor U3226 (N_3226,N_2194,N_2126);
or U3227 (N_3227,N_2782,N_2607);
nor U3228 (N_3228,N_2442,N_2732);
nor U3229 (N_3229,N_2551,N_2767);
or U3230 (N_3230,N_2065,N_2289);
nor U3231 (N_3231,N_2915,N_2332);
and U3232 (N_3232,N_2945,N_2371);
nor U3233 (N_3233,N_2630,N_2690);
and U3234 (N_3234,N_2874,N_2123);
nor U3235 (N_3235,N_2611,N_2170);
nand U3236 (N_3236,N_2615,N_2467);
and U3237 (N_3237,N_2995,N_2939);
nor U3238 (N_3238,N_2297,N_2774);
and U3239 (N_3239,N_2409,N_2974);
nand U3240 (N_3240,N_2403,N_2491);
and U3241 (N_3241,N_2851,N_2881);
nor U3242 (N_3242,N_2399,N_2698);
nand U3243 (N_3243,N_2037,N_2733);
or U3244 (N_3244,N_2592,N_2226);
or U3245 (N_3245,N_2041,N_2835);
nand U3246 (N_3246,N_2763,N_2537);
or U3247 (N_3247,N_2669,N_2001);
nand U3248 (N_3248,N_2689,N_2105);
and U3249 (N_3249,N_2840,N_2535);
or U3250 (N_3250,N_2599,N_2957);
or U3251 (N_3251,N_2329,N_2542);
nand U3252 (N_3252,N_2484,N_2990);
nand U3253 (N_3253,N_2206,N_2190);
and U3254 (N_3254,N_2889,N_2518);
or U3255 (N_3255,N_2013,N_2513);
nor U3256 (N_3256,N_2528,N_2871);
or U3257 (N_3257,N_2305,N_2503);
nor U3258 (N_3258,N_2910,N_2450);
nand U3259 (N_3259,N_2827,N_2785);
nand U3260 (N_3260,N_2717,N_2281);
nand U3261 (N_3261,N_2247,N_2486);
nor U3262 (N_3262,N_2459,N_2430);
nand U3263 (N_3263,N_2960,N_2858);
nand U3264 (N_3264,N_2776,N_2779);
or U3265 (N_3265,N_2446,N_2351);
nand U3266 (N_3266,N_2530,N_2710);
nand U3267 (N_3267,N_2274,N_2843);
and U3268 (N_3268,N_2461,N_2129);
or U3269 (N_3269,N_2000,N_2257);
nor U3270 (N_3270,N_2696,N_2046);
or U3271 (N_3271,N_2380,N_2719);
or U3272 (N_3272,N_2067,N_2264);
xor U3273 (N_3273,N_2155,N_2284);
nor U3274 (N_3274,N_2954,N_2475);
nor U3275 (N_3275,N_2179,N_2522);
nand U3276 (N_3276,N_2543,N_2166);
or U3277 (N_3277,N_2308,N_2558);
nor U3278 (N_3278,N_2404,N_2897);
and U3279 (N_3279,N_2629,N_2743);
nand U3280 (N_3280,N_2647,N_2823);
or U3281 (N_3281,N_2702,N_2241);
or U3282 (N_3282,N_2448,N_2086);
or U3283 (N_3283,N_2002,N_2873);
or U3284 (N_3284,N_2577,N_2504);
or U3285 (N_3285,N_2180,N_2145);
and U3286 (N_3286,N_2837,N_2258);
nand U3287 (N_3287,N_2078,N_2898);
and U3288 (N_3288,N_2367,N_2650);
nand U3289 (N_3289,N_2900,N_2660);
or U3290 (N_3290,N_2961,N_2374);
and U3291 (N_3291,N_2074,N_2830);
nor U3292 (N_3292,N_2713,N_2962);
nor U3293 (N_3293,N_2757,N_2684);
nand U3294 (N_3294,N_2178,N_2727);
nor U3295 (N_3295,N_2802,N_2070);
and U3296 (N_3296,N_2715,N_2083);
nand U3297 (N_3297,N_2346,N_2964);
or U3298 (N_3298,N_2421,N_2902);
nor U3299 (N_3299,N_2829,N_2514);
or U3300 (N_3300,N_2925,N_2807);
and U3301 (N_3301,N_2470,N_2923);
nand U3302 (N_3302,N_2242,N_2756);
or U3303 (N_3303,N_2541,N_2686);
nor U3304 (N_3304,N_2303,N_2695);
nor U3305 (N_3305,N_2202,N_2836);
nor U3306 (N_3306,N_2749,N_2464);
and U3307 (N_3307,N_2156,N_2921);
or U3308 (N_3308,N_2734,N_2133);
and U3309 (N_3309,N_2288,N_2429);
and U3310 (N_3310,N_2936,N_2433);
xor U3311 (N_3311,N_2127,N_2869);
and U3312 (N_3312,N_2985,N_2215);
or U3313 (N_3313,N_2844,N_2082);
and U3314 (N_3314,N_2455,N_2942);
or U3315 (N_3315,N_2066,N_2224);
nand U3316 (N_3316,N_2922,N_2494);
or U3317 (N_3317,N_2222,N_2999);
nand U3318 (N_3318,N_2752,N_2014);
nor U3319 (N_3319,N_2938,N_2087);
and U3320 (N_3320,N_2746,N_2775);
or U3321 (N_3321,N_2911,N_2131);
and U3322 (N_3322,N_2863,N_2711);
and U3323 (N_3323,N_2584,N_2933);
and U3324 (N_3324,N_2828,N_2209);
nor U3325 (N_3325,N_2379,N_2680);
or U3326 (N_3326,N_2296,N_2425);
nand U3327 (N_3327,N_2177,N_2534);
or U3328 (N_3328,N_2142,N_2572);
nor U3329 (N_3329,N_2076,N_2172);
nor U3330 (N_3330,N_2801,N_2707);
nand U3331 (N_3331,N_2639,N_2382);
and U3332 (N_3332,N_2723,N_2693);
nand U3333 (N_3333,N_2706,N_2388);
nor U3334 (N_3334,N_2965,N_2340);
and U3335 (N_3335,N_2633,N_2507);
and U3336 (N_3336,N_2725,N_2805);
nor U3337 (N_3337,N_2821,N_2575);
nand U3338 (N_3338,N_2090,N_2047);
xnor U3339 (N_3339,N_2302,N_2606);
nand U3340 (N_3340,N_2327,N_2483);
or U3341 (N_3341,N_2407,N_2101);
nor U3342 (N_3342,N_2389,N_2583);
nor U3343 (N_3343,N_2118,N_2393);
and U3344 (N_3344,N_2102,N_2249);
or U3345 (N_3345,N_2641,N_2217);
or U3346 (N_3346,N_2270,N_2811);
and U3347 (N_3347,N_2347,N_2741);
and U3348 (N_3348,N_2624,N_2096);
nor U3349 (N_3349,N_2926,N_2714);
and U3350 (N_3350,N_2589,N_2852);
nor U3351 (N_3351,N_2378,N_2784);
or U3352 (N_3352,N_2238,N_2631);
nor U3353 (N_3353,N_2220,N_2255);
xor U3354 (N_3354,N_2730,N_2729);
nor U3355 (N_3355,N_2508,N_2228);
nor U3356 (N_3356,N_2914,N_2449);
or U3357 (N_3357,N_2621,N_2754);
or U3358 (N_3358,N_2456,N_2618);
or U3359 (N_3359,N_2436,N_2867);
nor U3360 (N_3360,N_2197,N_2011);
xnor U3361 (N_3361,N_2972,N_2552);
or U3362 (N_3362,N_2943,N_2509);
or U3363 (N_3363,N_2571,N_2383);
nand U3364 (N_3364,N_2793,N_2765);
nand U3365 (N_3365,N_2309,N_2519);
nor U3366 (N_3366,N_2617,N_2254);
and U3367 (N_3367,N_2098,N_2742);
nand U3368 (N_3368,N_2110,N_2750);
nand U3369 (N_3369,N_2761,N_2778);
nand U3370 (N_3370,N_2276,N_2466);
and U3371 (N_3371,N_2841,N_2609);
and U3372 (N_3372,N_2512,N_2201);
nand U3373 (N_3373,N_2072,N_2683);
nand U3374 (N_3374,N_2161,N_2770);
and U3375 (N_3375,N_2529,N_2988);
and U3376 (N_3376,N_2815,N_2616);
nor U3377 (N_3377,N_2141,N_2094);
nand U3378 (N_3378,N_2416,N_2132);
nor U3379 (N_3379,N_2847,N_2566);
and U3380 (N_3380,N_2907,N_2903);
and U3381 (N_3381,N_2395,N_2544);
nand U3382 (N_3382,N_2967,N_2321);
and U3383 (N_3383,N_2798,N_2075);
xor U3384 (N_3384,N_2200,N_2039);
xnor U3385 (N_3385,N_2474,N_2608);
nand U3386 (N_3386,N_2160,N_2223);
and U3387 (N_3387,N_2657,N_2452);
nand U3388 (N_3388,N_2266,N_2968);
nand U3389 (N_3389,N_2745,N_2316);
or U3390 (N_3390,N_2256,N_2950);
or U3391 (N_3391,N_2554,N_2661);
or U3392 (N_3392,N_2991,N_2300);
xnor U3393 (N_3393,N_2855,N_2989);
or U3394 (N_3394,N_2490,N_2953);
and U3395 (N_3395,N_2064,N_2350);
nor U3396 (N_3396,N_2056,N_2428);
and U3397 (N_3397,N_2357,N_2006);
or U3398 (N_3398,N_2307,N_2103);
nor U3399 (N_3399,N_2868,N_2697);
and U3400 (N_3400,N_2614,N_2050);
and U3401 (N_3401,N_2753,N_2344);
and U3402 (N_3402,N_2471,N_2120);
and U3403 (N_3403,N_2342,N_2920);
nand U3404 (N_3404,N_2709,N_2679);
or U3405 (N_3405,N_2576,N_2998);
nand U3406 (N_3406,N_2135,N_2588);
and U3407 (N_3407,N_2929,N_2111);
and U3408 (N_3408,N_2883,N_2049);
nand U3409 (N_3409,N_2672,N_2077);
or U3410 (N_3410,N_2976,N_2597);
or U3411 (N_3411,N_2788,N_2814);
nor U3412 (N_3412,N_2687,N_2997);
or U3413 (N_3413,N_2604,N_2724);
nand U3414 (N_3414,N_2499,N_2591);
nor U3415 (N_3415,N_2042,N_2700);
nor U3416 (N_3416,N_2642,N_2229);
nor U3417 (N_3417,N_2859,N_2538);
or U3418 (N_3418,N_2722,N_2966);
nand U3419 (N_3419,N_2440,N_2295);
or U3420 (N_3420,N_2366,N_2140);
nand U3421 (N_3421,N_2396,N_2184);
and U3422 (N_3422,N_2996,N_2866);
or U3423 (N_3423,N_2375,N_2221);
and U3424 (N_3424,N_2213,N_2391);
nor U3425 (N_3425,N_2708,N_2971);
or U3426 (N_3426,N_2326,N_2139);
nand U3427 (N_3427,N_2313,N_2646);
or U3428 (N_3428,N_2320,N_2019);
and U3429 (N_3429,N_2093,N_2469);
nand U3430 (N_3430,N_2012,N_2427);
and U3431 (N_3431,N_2292,N_2992);
nand U3432 (N_3432,N_2932,N_2239);
and U3433 (N_3433,N_2196,N_2846);
and U3434 (N_3434,N_2113,N_2330);
and U3435 (N_3435,N_2269,N_2271);
nor U3436 (N_3436,N_2716,N_2352);
or U3437 (N_3437,N_2738,N_2557);
nor U3438 (N_3438,N_2880,N_2854);
or U3439 (N_3439,N_2620,N_2015);
nand U3440 (N_3440,N_2263,N_2970);
nor U3441 (N_3441,N_2279,N_2260);
or U3442 (N_3442,N_2465,N_2246);
nand U3443 (N_3443,N_2685,N_2909);
nor U3444 (N_3444,N_2487,N_2092);
and U3445 (N_3445,N_2137,N_2531);
nand U3446 (N_3446,N_2376,N_2354);
or U3447 (N_3447,N_2412,N_2505);
nand U3448 (N_3448,N_2568,N_2334);
or U3449 (N_3449,N_2878,N_2158);
and U3450 (N_3450,N_2506,N_2363);
nor U3451 (N_3451,N_2312,N_2058);
nor U3452 (N_3452,N_2941,N_2982);
and U3453 (N_3453,N_2099,N_2020);
or U3454 (N_3454,N_2034,N_2253);
nor U3455 (N_3455,N_2495,N_2790);
nor U3456 (N_3456,N_2605,N_2905);
and U3457 (N_3457,N_2028,N_2235);
or U3458 (N_3458,N_2386,N_2718);
nor U3459 (N_3459,N_2144,N_2392);
and U3460 (N_3460,N_2031,N_2073);
nand U3461 (N_3461,N_2414,N_2216);
nand U3462 (N_3462,N_2682,N_2688);
or U3463 (N_3463,N_2590,N_2348);
or U3464 (N_3464,N_2739,N_2564);
and U3465 (N_3465,N_2384,N_2768);
nand U3466 (N_3466,N_2489,N_2053);
nand U3467 (N_3467,N_2322,N_2171);
xnor U3468 (N_3468,N_2533,N_2397);
nand U3469 (N_3469,N_2008,N_2987);
nand U3470 (N_3470,N_2574,N_2203);
nand U3471 (N_3471,N_2771,N_2335);
and U3472 (N_3472,N_2453,N_2497);
nor U3473 (N_3473,N_2432,N_2955);
or U3474 (N_3474,N_2832,N_2462);
or U3475 (N_3475,N_2362,N_2454);
or U3476 (N_3476,N_2089,N_2117);
or U3477 (N_3477,N_2285,N_2703);
nor U3478 (N_3478,N_2167,N_2705);
or U3479 (N_3479,N_2174,N_2360);
nand U3480 (N_3480,N_2210,N_2291);
xor U3481 (N_3481,N_2510,N_2022);
nor U3482 (N_3482,N_2549,N_2645);
or U3483 (N_3483,N_2251,N_2797);
nor U3484 (N_3484,N_2336,N_2610);
nand U3485 (N_3485,N_2796,N_2227);
or U3486 (N_3486,N_2186,N_2817);
nor U3487 (N_3487,N_2124,N_2676);
and U3488 (N_3488,N_2301,N_2419);
nor U3489 (N_3489,N_2286,N_2580);
or U3490 (N_3490,N_2496,N_2478);
or U3491 (N_3491,N_2294,N_2045);
nor U3492 (N_3492,N_2816,N_2205);
or U3493 (N_3493,N_2198,N_2667);
xor U3494 (N_3494,N_2016,N_2664);
xor U3495 (N_3495,N_2848,N_2071);
nor U3496 (N_3496,N_2299,N_2937);
nand U3497 (N_3497,N_2550,N_2812);
nor U3498 (N_3498,N_2355,N_2410);
nand U3499 (N_3499,N_2864,N_2539);
nand U3500 (N_3500,N_2136,N_2517);
nand U3501 (N_3501,N_2708,N_2630);
nor U3502 (N_3502,N_2351,N_2546);
nand U3503 (N_3503,N_2473,N_2823);
or U3504 (N_3504,N_2915,N_2301);
nand U3505 (N_3505,N_2037,N_2194);
nor U3506 (N_3506,N_2007,N_2305);
or U3507 (N_3507,N_2655,N_2272);
or U3508 (N_3508,N_2210,N_2420);
nor U3509 (N_3509,N_2123,N_2087);
nand U3510 (N_3510,N_2924,N_2610);
nand U3511 (N_3511,N_2632,N_2328);
nand U3512 (N_3512,N_2169,N_2163);
nand U3513 (N_3513,N_2471,N_2427);
and U3514 (N_3514,N_2645,N_2599);
and U3515 (N_3515,N_2220,N_2762);
nand U3516 (N_3516,N_2587,N_2647);
nand U3517 (N_3517,N_2376,N_2146);
or U3518 (N_3518,N_2411,N_2597);
and U3519 (N_3519,N_2197,N_2697);
nand U3520 (N_3520,N_2065,N_2931);
and U3521 (N_3521,N_2075,N_2122);
and U3522 (N_3522,N_2264,N_2471);
and U3523 (N_3523,N_2224,N_2731);
nor U3524 (N_3524,N_2047,N_2279);
xor U3525 (N_3525,N_2832,N_2841);
nand U3526 (N_3526,N_2193,N_2674);
nand U3527 (N_3527,N_2788,N_2162);
nand U3528 (N_3528,N_2540,N_2572);
or U3529 (N_3529,N_2950,N_2543);
nand U3530 (N_3530,N_2995,N_2556);
or U3531 (N_3531,N_2872,N_2198);
nor U3532 (N_3532,N_2073,N_2626);
and U3533 (N_3533,N_2795,N_2581);
or U3534 (N_3534,N_2776,N_2533);
nand U3535 (N_3535,N_2594,N_2784);
xor U3536 (N_3536,N_2951,N_2507);
nand U3537 (N_3537,N_2976,N_2134);
nor U3538 (N_3538,N_2925,N_2847);
nand U3539 (N_3539,N_2581,N_2794);
xnor U3540 (N_3540,N_2630,N_2226);
or U3541 (N_3541,N_2245,N_2053);
and U3542 (N_3542,N_2572,N_2208);
or U3543 (N_3543,N_2868,N_2208);
nor U3544 (N_3544,N_2018,N_2486);
nand U3545 (N_3545,N_2531,N_2159);
and U3546 (N_3546,N_2437,N_2680);
nand U3547 (N_3547,N_2919,N_2266);
and U3548 (N_3548,N_2799,N_2679);
or U3549 (N_3549,N_2840,N_2192);
or U3550 (N_3550,N_2954,N_2466);
or U3551 (N_3551,N_2355,N_2356);
nor U3552 (N_3552,N_2301,N_2063);
nand U3553 (N_3553,N_2582,N_2764);
or U3554 (N_3554,N_2503,N_2047);
or U3555 (N_3555,N_2302,N_2747);
nor U3556 (N_3556,N_2736,N_2030);
nor U3557 (N_3557,N_2314,N_2113);
and U3558 (N_3558,N_2750,N_2051);
or U3559 (N_3559,N_2388,N_2536);
nand U3560 (N_3560,N_2111,N_2899);
nand U3561 (N_3561,N_2057,N_2594);
or U3562 (N_3562,N_2105,N_2247);
and U3563 (N_3563,N_2835,N_2749);
and U3564 (N_3564,N_2916,N_2420);
nor U3565 (N_3565,N_2928,N_2582);
xor U3566 (N_3566,N_2063,N_2431);
or U3567 (N_3567,N_2723,N_2701);
nor U3568 (N_3568,N_2188,N_2876);
nor U3569 (N_3569,N_2372,N_2035);
nand U3570 (N_3570,N_2898,N_2643);
nand U3571 (N_3571,N_2299,N_2935);
nor U3572 (N_3572,N_2134,N_2477);
xnor U3573 (N_3573,N_2692,N_2689);
or U3574 (N_3574,N_2134,N_2653);
nand U3575 (N_3575,N_2345,N_2008);
xnor U3576 (N_3576,N_2825,N_2424);
nor U3577 (N_3577,N_2108,N_2940);
or U3578 (N_3578,N_2096,N_2072);
nor U3579 (N_3579,N_2466,N_2713);
and U3580 (N_3580,N_2295,N_2706);
or U3581 (N_3581,N_2135,N_2012);
or U3582 (N_3582,N_2520,N_2003);
nand U3583 (N_3583,N_2497,N_2012);
or U3584 (N_3584,N_2862,N_2637);
and U3585 (N_3585,N_2377,N_2315);
nor U3586 (N_3586,N_2933,N_2516);
and U3587 (N_3587,N_2732,N_2630);
and U3588 (N_3588,N_2169,N_2342);
and U3589 (N_3589,N_2930,N_2478);
or U3590 (N_3590,N_2291,N_2273);
nand U3591 (N_3591,N_2876,N_2125);
nor U3592 (N_3592,N_2180,N_2945);
or U3593 (N_3593,N_2130,N_2129);
nor U3594 (N_3594,N_2496,N_2888);
nor U3595 (N_3595,N_2884,N_2574);
and U3596 (N_3596,N_2887,N_2577);
nor U3597 (N_3597,N_2573,N_2933);
and U3598 (N_3598,N_2140,N_2202);
or U3599 (N_3599,N_2038,N_2919);
nor U3600 (N_3600,N_2203,N_2467);
and U3601 (N_3601,N_2331,N_2107);
nand U3602 (N_3602,N_2898,N_2583);
or U3603 (N_3603,N_2347,N_2875);
and U3604 (N_3604,N_2154,N_2622);
xor U3605 (N_3605,N_2116,N_2988);
nor U3606 (N_3606,N_2065,N_2333);
nand U3607 (N_3607,N_2378,N_2100);
nor U3608 (N_3608,N_2497,N_2883);
nor U3609 (N_3609,N_2227,N_2397);
nand U3610 (N_3610,N_2329,N_2725);
or U3611 (N_3611,N_2457,N_2678);
nand U3612 (N_3612,N_2505,N_2557);
nand U3613 (N_3613,N_2547,N_2017);
and U3614 (N_3614,N_2160,N_2112);
nand U3615 (N_3615,N_2903,N_2037);
nor U3616 (N_3616,N_2073,N_2523);
nor U3617 (N_3617,N_2626,N_2149);
and U3618 (N_3618,N_2784,N_2080);
nor U3619 (N_3619,N_2027,N_2391);
nand U3620 (N_3620,N_2552,N_2032);
or U3621 (N_3621,N_2748,N_2523);
or U3622 (N_3622,N_2643,N_2415);
nor U3623 (N_3623,N_2334,N_2532);
nand U3624 (N_3624,N_2668,N_2780);
or U3625 (N_3625,N_2988,N_2947);
or U3626 (N_3626,N_2130,N_2439);
nor U3627 (N_3627,N_2737,N_2534);
and U3628 (N_3628,N_2469,N_2941);
nor U3629 (N_3629,N_2954,N_2177);
and U3630 (N_3630,N_2055,N_2072);
nand U3631 (N_3631,N_2320,N_2818);
nand U3632 (N_3632,N_2161,N_2149);
nand U3633 (N_3633,N_2365,N_2498);
and U3634 (N_3634,N_2805,N_2125);
or U3635 (N_3635,N_2169,N_2485);
nor U3636 (N_3636,N_2371,N_2564);
nand U3637 (N_3637,N_2772,N_2063);
or U3638 (N_3638,N_2465,N_2183);
nand U3639 (N_3639,N_2499,N_2996);
nor U3640 (N_3640,N_2508,N_2234);
and U3641 (N_3641,N_2962,N_2380);
nand U3642 (N_3642,N_2742,N_2575);
nand U3643 (N_3643,N_2874,N_2926);
nand U3644 (N_3644,N_2277,N_2243);
nor U3645 (N_3645,N_2732,N_2992);
nand U3646 (N_3646,N_2620,N_2229);
and U3647 (N_3647,N_2754,N_2507);
and U3648 (N_3648,N_2785,N_2856);
nand U3649 (N_3649,N_2239,N_2820);
or U3650 (N_3650,N_2578,N_2990);
and U3651 (N_3651,N_2801,N_2257);
and U3652 (N_3652,N_2656,N_2369);
nand U3653 (N_3653,N_2632,N_2741);
nor U3654 (N_3654,N_2851,N_2333);
and U3655 (N_3655,N_2018,N_2812);
or U3656 (N_3656,N_2160,N_2395);
or U3657 (N_3657,N_2757,N_2131);
and U3658 (N_3658,N_2571,N_2069);
and U3659 (N_3659,N_2388,N_2646);
nand U3660 (N_3660,N_2101,N_2998);
or U3661 (N_3661,N_2983,N_2504);
or U3662 (N_3662,N_2863,N_2679);
nand U3663 (N_3663,N_2737,N_2304);
and U3664 (N_3664,N_2133,N_2517);
nand U3665 (N_3665,N_2356,N_2149);
nor U3666 (N_3666,N_2377,N_2470);
nand U3667 (N_3667,N_2219,N_2589);
nor U3668 (N_3668,N_2972,N_2709);
nand U3669 (N_3669,N_2573,N_2744);
nor U3670 (N_3670,N_2972,N_2590);
nor U3671 (N_3671,N_2843,N_2643);
or U3672 (N_3672,N_2163,N_2174);
nor U3673 (N_3673,N_2809,N_2795);
or U3674 (N_3674,N_2799,N_2728);
or U3675 (N_3675,N_2705,N_2365);
nand U3676 (N_3676,N_2892,N_2272);
nor U3677 (N_3677,N_2791,N_2592);
nand U3678 (N_3678,N_2771,N_2641);
or U3679 (N_3679,N_2672,N_2308);
and U3680 (N_3680,N_2185,N_2800);
or U3681 (N_3681,N_2147,N_2893);
nand U3682 (N_3682,N_2841,N_2033);
nor U3683 (N_3683,N_2827,N_2430);
nand U3684 (N_3684,N_2898,N_2957);
nand U3685 (N_3685,N_2655,N_2398);
or U3686 (N_3686,N_2074,N_2431);
nand U3687 (N_3687,N_2739,N_2231);
or U3688 (N_3688,N_2544,N_2136);
nand U3689 (N_3689,N_2738,N_2502);
or U3690 (N_3690,N_2375,N_2693);
or U3691 (N_3691,N_2642,N_2729);
nor U3692 (N_3692,N_2748,N_2176);
nor U3693 (N_3693,N_2188,N_2276);
and U3694 (N_3694,N_2127,N_2059);
or U3695 (N_3695,N_2207,N_2252);
nor U3696 (N_3696,N_2173,N_2215);
or U3697 (N_3697,N_2786,N_2190);
nor U3698 (N_3698,N_2516,N_2585);
nand U3699 (N_3699,N_2949,N_2098);
or U3700 (N_3700,N_2611,N_2407);
nor U3701 (N_3701,N_2073,N_2484);
or U3702 (N_3702,N_2884,N_2424);
or U3703 (N_3703,N_2714,N_2454);
and U3704 (N_3704,N_2734,N_2120);
nand U3705 (N_3705,N_2748,N_2633);
and U3706 (N_3706,N_2377,N_2719);
or U3707 (N_3707,N_2285,N_2942);
and U3708 (N_3708,N_2250,N_2652);
and U3709 (N_3709,N_2207,N_2343);
nor U3710 (N_3710,N_2571,N_2969);
or U3711 (N_3711,N_2634,N_2826);
nor U3712 (N_3712,N_2961,N_2033);
and U3713 (N_3713,N_2679,N_2827);
and U3714 (N_3714,N_2720,N_2410);
or U3715 (N_3715,N_2509,N_2338);
or U3716 (N_3716,N_2239,N_2512);
and U3717 (N_3717,N_2127,N_2577);
or U3718 (N_3718,N_2033,N_2234);
and U3719 (N_3719,N_2387,N_2649);
and U3720 (N_3720,N_2176,N_2240);
and U3721 (N_3721,N_2453,N_2061);
nor U3722 (N_3722,N_2470,N_2830);
and U3723 (N_3723,N_2385,N_2214);
and U3724 (N_3724,N_2967,N_2538);
or U3725 (N_3725,N_2577,N_2518);
nand U3726 (N_3726,N_2746,N_2619);
nand U3727 (N_3727,N_2467,N_2611);
or U3728 (N_3728,N_2098,N_2443);
nand U3729 (N_3729,N_2844,N_2169);
or U3730 (N_3730,N_2039,N_2516);
nor U3731 (N_3731,N_2438,N_2330);
nand U3732 (N_3732,N_2070,N_2814);
and U3733 (N_3733,N_2960,N_2958);
nor U3734 (N_3734,N_2263,N_2750);
nor U3735 (N_3735,N_2530,N_2294);
nor U3736 (N_3736,N_2160,N_2693);
nand U3737 (N_3737,N_2874,N_2818);
nand U3738 (N_3738,N_2447,N_2994);
nand U3739 (N_3739,N_2507,N_2925);
nand U3740 (N_3740,N_2382,N_2347);
nor U3741 (N_3741,N_2807,N_2420);
nand U3742 (N_3742,N_2779,N_2800);
and U3743 (N_3743,N_2660,N_2111);
nor U3744 (N_3744,N_2232,N_2622);
and U3745 (N_3745,N_2792,N_2256);
and U3746 (N_3746,N_2603,N_2833);
and U3747 (N_3747,N_2241,N_2695);
nor U3748 (N_3748,N_2232,N_2653);
and U3749 (N_3749,N_2823,N_2271);
or U3750 (N_3750,N_2304,N_2085);
or U3751 (N_3751,N_2584,N_2222);
nor U3752 (N_3752,N_2289,N_2960);
nand U3753 (N_3753,N_2831,N_2596);
nor U3754 (N_3754,N_2524,N_2794);
nand U3755 (N_3755,N_2823,N_2431);
nor U3756 (N_3756,N_2500,N_2290);
and U3757 (N_3757,N_2845,N_2643);
nand U3758 (N_3758,N_2435,N_2289);
nand U3759 (N_3759,N_2083,N_2349);
nor U3760 (N_3760,N_2336,N_2257);
nor U3761 (N_3761,N_2587,N_2907);
nor U3762 (N_3762,N_2779,N_2026);
nand U3763 (N_3763,N_2551,N_2071);
nand U3764 (N_3764,N_2589,N_2748);
or U3765 (N_3765,N_2127,N_2209);
or U3766 (N_3766,N_2109,N_2695);
and U3767 (N_3767,N_2477,N_2796);
and U3768 (N_3768,N_2646,N_2998);
nand U3769 (N_3769,N_2574,N_2491);
nand U3770 (N_3770,N_2621,N_2297);
or U3771 (N_3771,N_2151,N_2779);
nor U3772 (N_3772,N_2858,N_2670);
nand U3773 (N_3773,N_2403,N_2257);
and U3774 (N_3774,N_2606,N_2685);
or U3775 (N_3775,N_2700,N_2633);
or U3776 (N_3776,N_2098,N_2638);
and U3777 (N_3777,N_2532,N_2400);
nand U3778 (N_3778,N_2344,N_2423);
and U3779 (N_3779,N_2519,N_2105);
nand U3780 (N_3780,N_2426,N_2963);
nand U3781 (N_3781,N_2504,N_2209);
and U3782 (N_3782,N_2853,N_2119);
or U3783 (N_3783,N_2325,N_2971);
or U3784 (N_3784,N_2602,N_2079);
nand U3785 (N_3785,N_2445,N_2873);
or U3786 (N_3786,N_2344,N_2177);
and U3787 (N_3787,N_2362,N_2154);
xnor U3788 (N_3788,N_2124,N_2371);
nor U3789 (N_3789,N_2602,N_2419);
or U3790 (N_3790,N_2868,N_2615);
nand U3791 (N_3791,N_2690,N_2216);
and U3792 (N_3792,N_2513,N_2920);
and U3793 (N_3793,N_2823,N_2573);
nor U3794 (N_3794,N_2413,N_2858);
or U3795 (N_3795,N_2011,N_2394);
nor U3796 (N_3796,N_2467,N_2139);
or U3797 (N_3797,N_2375,N_2513);
nand U3798 (N_3798,N_2741,N_2978);
or U3799 (N_3799,N_2560,N_2871);
nand U3800 (N_3800,N_2627,N_2840);
nand U3801 (N_3801,N_2436,N_2804);
nor U3802 (N_3802,N_2843,N_2051);
nor U3803 (N_3803,N_2909,N_2911);
nand U3804 (N_3804,N_2323,N_2135);
nor U3805 (N_3805,N_2339,N_2364);
and U3806 (N_3806,N_2819,N_2015);
nand U3807 (N_3807,N_2126,N_2887);
nand U3808 (N_3808,N_2444,N_2482);
and U3809 (N_3809,N_2266,N_2225);
and U3810 (N_3810,N_2164,N_2693);
or U3811 (N_3811,N_2541,N_2201);
nor U3812 (N_3812,N_2138,N_2607);
nand U3813 (N_3813,N_2423,N_2291);
nand U3814 (N_3814,N_2197,N_2031);
nor U3815 (N_3815,N_2417,N_2749);
nor U3816 (N_3816,N_2898,N_2779);
and U3817 (N_3817,N_2780,N_2237);
and U3818 (N_3818,N_2116,N_2373);
and U3819 (N_3819,N_2916,N_2735);
nor U3820 (N_3820,N_2922,N_2844);
and U3821 (N_3821,N_2760,N_2629);
nor U3822 (N_3822,N_2747,N_2593);
and U3823 (N_3823,N_2324,N_2772);
or U3824 (N_3824,N_2771,N_2591);
nor U3825 (N_3825,N_2698,N_2453);
and U3826 (N_3826,N_2145,N_2128);
nand U3827 (N_3827,N_2735,N_2198);
and U3828 (N_3828,N_2621,N_2321);
or U3829 (N_3829,N_2624,N_2786);
nor U3830 (N_3830,N_2178,N_2869);
or U3831 (N_3831,N_2474,N_2352);
nor U3832 (N_3832,N_2041,N_2621);
nand U3833 (N_3833,N_2506,N_2478);
and U3834 (N_3834,N_2138,N_2249);
and U3835 (N_3835,N_2961,N_2258);
nor U3836 (N_3836,N_2014,N_2205);
nand U3837 (N_3837,N_2330,N_2695);
nor U3838 (N_3838,N_2860,N_2689);
nand U3839 (N_3839,N_2727,N_2244);
or U3840 (N_3840,N_2825,N_2551);
nand U3841 (N_3841,N_2495,N_2689);
nor U3842 (N_3842,N_2756,N_2921);
and U3843 (N_3843,N_2008,N_2044);
or U3844 (N_3844,N_2415,N_2427);
nor U3845 (N_3845,N_2404,N_2271);
nand U3846 (N_3846,N_2852,N_2685);
or U3847 (N_3847,N_2339,N_2849);
nor U3848 (N_3848,N_2708,N_2266);
or U3849 (N_3849,N_2399,N_2426);
nand U3850 (N_3850,N_2631,N_2448);
nor U3851 (N_3851,N_2248,N_2106);
and U3852 (N_3852,N_2526,N_2166);
or U3853 (N_3853,N_2306,N_2684);
nor U3854 (N_3854,N_2825,N_2542);
xnor U3855 (N_3855,N_2455,N_2326);
and U3856 (N_3856,N_2898,N_2686);
nor U3857 (N_3857,N_2659,N_2254);
xor U3858 (N_3858,N_2635,N_2600);
nand U3859 (N_3859,N_2268,N_2288);
and U3860 (N_3860,N_2616,N_2673);
nand U3861 (N_3861,N_2214,N_2575);
and U3862 (N_3862,N_2919,N_2564);
or U3863 (N_3863,N_2251,N_2603);
or U3864 (N_3864,N_2762,N_2377);
nand U3865 (N_3865,N_2811,N_2486);
nand U3866 (N_3866,N_2693,N_2363);
or U3867 (N_3867,N_2666,N_2584);
nor U3868 (N_3868,N_2190,N_2143);
and U3869 (N_3869,N_2470,N_2698);
and U3870 (N_3870,N_2011,N_2261);
and U3871 (N_3871,N_2208,N_2687);
nor U3872 (N_3872,N_2161,N_2071);
or U3873 (N_3873,N_2970,N_2139);
or U3874 (N_3874,N_2303,N_2374);
or U3875 (N_3875,N_2155,N_2665);
nor U3876 (N_3876,N_2158,N_2138);
or U3877 (N_3877,N_2954,N_2355);
nand U3878 (N_3878,N_2597,N_2925);
and U3879 (N_3879,N_2498,N_2516);
or U3880 (N_3880,N_2310,N_2140);
nor U3881 (N_3881,N_2490,N_2704);
or U3882 (N_3882,N_2522,N_2353);
or U3883 (N_3883,N_2343,N_2306);
or U3884 (N_3884,N_2563,N_2872);
and U3885 (N_3885,N_2503,N_2540);
nor U3886 (N_3886,N_2567,N_2319);
and U3887 (N_3887,N_2719,N_2909);
xor U3888 (N_3888,N_2493,N_2896);
nand U3889 (N_3889,N_2420,N_2862);
nor U3890 (N_3890,N_2458,N_2229);
nor U3891 (N_3891,N_2657,N_2256);
nand U3892 (N_3892,N_2986,N_2563);
or U3893 (N_3893,N_2562,N_2459);
nand U3894 (N_3894,N_2633,N_2403);
nand U3895 (N_3895,N_2085,N_2041);
or U3896 (N_3896,N_2375,N_2873);
nor U3897 (N_3897,N_2738,N_2477);
nor U3898 (N_3898,N_2160,N_2834);
nand U3899 (N_3899,N_2002,N_2029);
or U3900 (N_3900,N_2317,N_2304);
and U3901 (N_3901,N_2018,N_2152);
nor U3902 (N_3902,N_2156,N_2773);
nand U3903 (N_3903,N_2293,N_2192);
nand U3904 (N_3904,N_2004,N_2521);
or U3905 (N_3905,N_2687,N_2085);
and U3906 (N_3906,N_2808,N_2855);
and U3907 (N_3907,N_2663,N_2176);
or U3908 (N_3908,N_2833,N_2765);
nand U3909 (N_3909,N_2376,N_2202);
nor U3910 (N_3910,N_2646,N_2929);
and U3911 (N_3911,N_2580,N_2101);
nor U3912 (N_3912,N_2336,N_2467);
nand U3913 (N_3913,N_2079,N_2574);
and U3914 (N_3914,N_2971,N_2833);
and U3915 (N_3915,N_2936,N_2216);
nand U3916 (N_3916,N_2762,N_2847);
nand U3917 (N_3917,N_2667,N_2897);
nand U3918 (N_3918,N_2205,N_2501);
and U3919 (N_3919,N_2567,N_2317);
nor U3920 (N_3920,N_2237,N_2151);
nor U3921 (N_3921,N_2987,N_2717);
nor U3922 (N_3922,N_2439,N_2019);
nand U3923 (N_3923,N_2730,N_2566);
or U3924 (N_3924,N_2734,N_2812);
xor U3925 (N_3925,N_2397,N_2366);
or U3926 (N_3926,N_2346,N_2309);
nand U3927 (N_3927,N_2254,N_2662);
or U3928 (N_3928,N_2532,N_2020);
and U3929 (N_3929,N_2622,N_2353);
nand U3930 (N_3930,N_2523,N_2407);
nor U3931 (N_3931,N_2676,N_2766);
or U3932 (N_3932,N_2118,N_2407);
nand U3933 (N_3933,N_2511,N_2668);
and U3934 (N_3934,N_2448,N_2859);
nand U3935 (N_3935,N_2169,N_2309);
nor U3936 (N_3936,N_2401,N_2121);
nand U3937 (N_3937,N_2877,N_2695);
nor U3938 (N_3938,N_2748,N_2025);
nand U3939 (N_3939,N_2973,N_2250);
and U3940 (N_3940,N_2715,N_2820);
nand U3941 (N_3941,N_2514,N_2980);
and U3942 (N_3942,N_2582,N_2306);
nand U3943 (N_3943,N_2859,N_2202);
nor U3944 (N_3944,N_2222,N_2738);
nand U3945 (N_3945,N_2283,N_2184);
and U3946 (N_3946,N_2798,N_2953);
nand U3947 (N_3947,N_2820,N_2513);
nor U3948 (N_3948,N_2231,N_2829);
and U3949 (N_3949,N_2540,N_2147);
nor U3950 (N_3950,N_2810,N_2369);
or U3951 (N_3951,N_2452,N_2379);
nand U3952 (N_3952,N_2402,N_2118);
nand U3953 (N_3953,N_2253,N_2839);
nor U3954 (N_3954,N_2844,N_2656);
and U3955 (N_3955,N_2615,N_2168);
nand U3956 (N_3956,N_2605,N_2137);
nand U3957 (N_3957,N_2515,N_2224);
and U3958 (N_3958,N_2497,N_2969);
and U3959 (N_3959,N_2212,N_2440);
or U3960 (N_3960,N_2735,N_2027);
or U3961 (N_3961,N_2603,N_2614);
and U3962 (N_3962,N_2772,N_2515);
nor U3963 (N_3963,N_2108,N_2645);
nand U3964 (N_3964,N_2597,N_2076);
and U3965 (N_3965,N_2031,N_2218);
nor U3966 (N_3966,N_2488,N_2134);
or U3967 (N_3967,N_2301,N_2056);
nand U3968 (N_3968,N_2461,N_2130);
and U3969 (N_3969,N_2639,N_2391);
and U3970 (N_3970,N_2063,N_2261);
xor U3971 (N_3971,N_2127,N_2855);
nor U3972 (N_3972,N_2958,N_2351);
nand U3973 (N_3973,N_2877,N_2709);
nand U3974 (N_3974,N_2224,N_2885);
nor U3975 (N_3975,N_2567,N_2836);
and U3976 (N_3976,N_2863,N_2489);
and U3977 (N_3977,N_2569,N_2738);
and U3978 (N_3978,N_2580,N_2609);
and U3979 (N_3979,N_2460,N_2637);
nand U3980 (N_3980,N_2875,N_2728);
nand U3981 (N_3981,N_2585,N_2853);
and U3982 (N_3982,N_2371,N_2803);
or U3983 (N_3983,N_2356,N_2055);
nor U3984 (N_3984,N_2019,N_2971);
and U3985 (N_3985,N_2171,N_2471);
or U3986 (N_3986,N_2336,N_2171);
and U3987 (N_3987,N_2490,N_2832);
nand U3988 (N_3988,N_2099,N_2745);
nand U3989 (N_3989,N_2059,N_2997);
and U3990 (N_3990,N_2734,N_2212);
and U3991 (N_3991,N_2102,N_2229);
and U3992 (N_3992,N_2921,N_2805);
and U3993 (N_3993,N_2141,N_2482);
and U3994 (N_3994,N_2682,N_2711);
nand U3995 (N_3995,N_2753,N_2237);
nor U3996 (N_3996,N_2138,N_2572);
xnor U3997 (N_3997,N_2699,N_2166);
or U3998 (N_3998,N_2227,N_2001);
and U3999 (N_3999,N_2596,N_2248);
or U4000 (N_4000,N_3676,N_3065);
or U4001 (N_4001,N_3947,N_3636);
or U4002 (N_4002,N_3954,N_3935);
nand U4003 (N_4003,N_3920,N_3200);
and U4004 (N_4004,N_3258,N_3378);
or U4005 (N_4005,N_3777,N_3529);
nor U4006 (N_4006,N_3774,N_3376);
nand U4007 (N_4007,N_3907,N_3773);
and U4008 (N_4008,N_3639,N_3230);
or U4009 (N_4009,N_3135,N_3081);
nor U4010 (N_4010,N_3006,N_3345);
or U4011 (N_4011,N_3027,N_3609);
or U4012 (N_4012,N_3829,N_3956);
nand U4013 (N_4013,N_3674,N_3323);
nor U4014 (N_4014,N_3998,N_3790);
xor U4015 (N_4015,N_3978,N_3382);
or U4016 (N_4016,N_3386,N_3291);
nand U4017 (N_4017,N_3955,N_3061);
xor U4018 (N_4018,N_3976,N_3002);
nor U4019 (N_4019,N_3940,N_3595);
nor U4020 (N_4020,N_3614,N_3255);
xnor U4021 (N_4021,N_3422,N_3951);
and U4022 (N_4022,N_3884,N_3821);
and U4023 (N_4023,N_3154,N_3669);
nand U4024 (N_4024,N_3311,N_3656);
and U4025 (N_4025,N_3764,N_3279);
nand U4026 (N_4026,N_3041,N_3072);
nor U4027 (N_4027,N_3520,N_3138);
nand U4028 (N_4028,N_3387,N_3144);
nand U4029 (N_4029,N_3148,N_3496);
nor U4030 (N_4030,N_3872,N_3199);
and U4031 (N_4031,N_3886,N_3342);
xor U4032 (N_4032,N_3729,N_3835);
and U4033 (N_4033,N_3441,N_3557);
and U4034 (N_4034,N_3256,N_3352);
nor U4035 (N_4035,N_3048,N_3592);
or U4036 (N_4036,N_3681,N_3887);
and U4037 (N_4037,N_3848,N_3085);
and U4038 (N_4038,N_3899,N_3815);
or U4039 (N_4039,N_3314,N_3984);
nor U4040 (N_4040,N_3634,N_3379);
nand U4041 (N_4041,N_3110,N_3745);
nand U4042 (N_4042,N_3056,N_3626);
xor U4043 (N_4043,N_3740,N_3555);
nor U4044 (N_4044,N_3938,N_3748);
or U4045 (N_4045,N_3599,N_3414);
nor U4046 (N_4046,N_3469,N_3466);
nand U4047 (N_4047,N_3299,N_3460);
and U4048 (N_4048,N_3807,N_3753);
nor U4049 (N_4049,N_3127,N_3250);
and U4050 (N_4050,N_3217,N_3194);
or U4051 (N_4051,N_3670,N_3131);
nand U4052 (N_4052,N_3475,N_3703);
and U4053 (N_4053,N_3248,N_3343);
nor U4054 (N_4054,N_3123,N_3071);
nor U4055 (N_4055,N_3948,N_3627);
or U4056 (N_4056,N_3915,N_3397);
and U4057 (N_4057,N_3846,N_3814);
or U4058 (N_4058,N_3507,N_3327);
and U4059 (N_4059,N_3488,N_3827);
and U4060 (N_4060,N_3518,N_3996);
and U4061 (N_4061,N_3730,N_3832);
or U4062 (N_4062,N_3057,N_3362);
or U4063 (N_4063,N_3128,N_3042);
and U4064 (N_4064,N_3452,N_3541);
and U4065 (N_4065,N_3337,N_3544);
and U4066 (N_4066,N_3623,N_3186);
and U4067 (N_4067,N_3543,N_3432);
nand U4068 (N_4068,N_3744,N_3310);
nor U4069 (N_4069,N_3263,N_3140);
and U4070 (N_4070,N_3408,N_3303);
nand U4071 (N_4071,N_3980,N_3563);
or U4072 (N_4072,N_3179,N_3741);
nor U4073 (N_4073,N_3137,N_3019);
nand U4074 (N_4074,N_3348,N_3715);
or U4075 (N_4075,N_3638,N_3000);
and U4076 (N_4076,N_3463,N_3569);
and U4077 (N_4077,N_3244,N_3805);
and U4078 (N_4078,N_3582,N_3806);
nand U4079 (N_4079,N_3032,N_3702);
and U4080 (N_4080,N_3666,N_3124);
and U4081 (N_4081,N_3210,N_3995);
or U4082 (N_4082,N_3714,N_3163);
xor U4083 (N_4083,N_3937,N_3840);
nand U4084 (N_4084,N_3024,N_3005);
and U4085 (N_4085,N_3369,N_3487);
and U4086 (N_4086,N_3690,N_3107);
and U4087 (N_4087,N_3063,N_3738);
nor U4088 (N_4088,N_3377,N_3685);
and U4089 (N_4089,N_3007,N_3578);
nor U4090 (N_4090,N_3853,N_3062);
or U4091 (N_4091,N_3818,N_3118);
nor U4092 (N_4092,N_3917,N_3500);
nor U4093 (N_4093,N_3657,N_3608);
xnor U4094 (N_4094,N_3304,N_3012);
or U4095 (N_4095,N_3939,N_3548);
nand U4096 (N_4096,N_3338,N_3420);
and U4097 (N_4097,N_3506,N_3227);
and U4098 (N_4098,N_3981,N_3439);
nand U4099 (N_4099,N_3510,N_3795);
or U4100 (N_4100,N_3659,N_3859);
or U4101 (N_4101,N_3589,N_3178);
or U4102 (N_4102,N_3016,N_3476);
nand U4103 (N_4103,N_3285,N_3246);
nor U4104 (N_4104,N_3698,N_3363);
or U4105 (N_4105,N_3169,N_3885);
nor U4106 (N_4106,N_3394,N_3473);
and U4107 (N_4107,N_3551,N_3992);
or U4108 (N_4108,N_3413,N_3309);
nand U4109 (N_4109,N_3326,N_3407);
nor U4110 (N_4110,N_3001,N_3538);
nor U4111 (N_4111,N_3882,N_3651);
or U4112 (N_4112,N_3416,N_3811);
nand U4113 (N_4113,N_3950,N_3347);
nor U4114 (N_4114,N_3521,N_3874);
and U4115 (N_4115,N_3236,N_3550);
nand U4116 (N_4116,N_3704,N_3328);
nor U4117 (N_4117,N_3017,N_3505);
and U4118 (N_4118,N_3008,N_3504);
nor U4119 (N_4119,N_3812,N_3214);
nor U4120 (N_4120,N_3604,N_3332);
and U4121 (N_4121,N_3393,N_3883);
nor U4122 (N_4122,N_3784,N_3875);
xor U4123 (N_4123,N_3161,N_3442);
nor U4124 (N_4124,N_3316,N_3096);
xnor U4125 (N_4125,N_3403,N_3864);
or U4126 (N_4126,N_3440,N_3453);
nand U4127 (N_4127,N_3406,N_3173);
nor U4128 (N_4128,N_3726,N_3512);
nor U4129 (N_4129,N_3216,N_3919);
and U4130 (N_4130,N_3121,N_3423);
and U4131 (N_4131,N_3014,N_3390);
or U4132 (N_4132,N_3411,N_3464);
nand U4133 (N_4133,N_3459,N_3513);
nor U4134 (N_4134,N_3725,N_3718);
nor U4135 (N_4135,N_3974,N_3064);
nand U4136 (N_4136,N_3040,N_3828);
and U4137 (N_4137,N_3241,N_3486);
or U4138 (N_4138,N_3191,N_3755);
and U4139 (N_4139,N_3136,N_3746);
or U4140 (N_4140,N_3896,N_3462);
or U4141 (N_4141,N_3372,N_3943);
or U4142 (N_4142,N_3203,N_3713);
or U4143 (N_4143,N_3108,N_3759);
nor U4144 (N_4144,N_3038,N_3105);
nand U4145 (N_4145,N_3461,N_3305);
nor U4146 (N_4146,N_3170,N_3498);
and U4147 (N_4147,N_3426,N_3590);
or U4148 (N_4148,N_3101,N_3801);
nand U4149 (N_4149,N_3654,N_3572);
and U4150 (N_4150,N_3830,N_3100);
and U4151 (N_4151,N_3259,N_3571);
nor U4152 (N_4152,N_3116,N_3990);
nor U4153 (N_4153,N_3458,N_3554);
nor U4154 (N_4154,N_3999,N_3152);
nor U4155 (N_4155,N_3942,N_3301);
nor U4156 (N_4156,N_3257,N_3562);
or U4157 (N_4157,N_3192,N_3252);
and U4158 (N_4158,N_3953,N_3810);
nor U4159 (N_4159,N_3537,N_3854);
and U4160 (N_4160,N_3766,N_3941);
nand U4161 (N_4161,N_3059,N_3535);
or U4162 (N_4162,N_3679,N_3353);
and U4163 (N_4163,N_3763,N_3392);
nor U4164 (N_4164,N_3606,N_3313);
and U4165 (N_4165,N_3825,N_3682);
nor U4166 (N_4166,N_3662,N_3644);
and U4167 (N_4167,N_3208,N_3479);
nand U4168 (N_4168,N_3201,N_3404);
and U4169 (N_4169,N_3616,N_3568);
and U4170 (N_4170,N_3261,N_3972);
or U4171 (N_4171,N_3735,N_3325);
and U4172 (N_4172,N_3482,N_3477);
nand U4173 (N_4173,N_3388,N_3402);
nor U4174 (N_4174,N_3286,N_3333);
and U4175 (N_4175,N_3485,N_3354);
or U4176 (N_4176,N_3078,N_3904);
nor U4177 (N_4177,N_3962,N_3558);
and U4178 (N_4178,N_3223,N_3357);
xnor U4179 (N_4179,N_3076,N_3973);
xor U4180 (N_4180,N_3794,N_3142);
and U4181 (N_4181,N_3160,N_3130);
or U4182 (N_4182,N_3033,N_3364);
or U4183 (N_4183,N_3637,N_3080);
nor U4184 (N_4184,N_3119,N_3916);
nand U4185 (N_4185,N_3022,N_3028);
and U4186 (N_4186,N_3985,N_3923);
and U4187 (N_4187,N_3297,N_3360);
nor U4188 (N_4188,N_3232,N_3576);
and U4189 (N_4189,N_3909,N_3092);
nand U4190 (N_4190,N_3594,N_3046);
and U4191 (N_4191,N_3172,N_3819);
or U4192 (N_4192,N_3969,N_3077);
and U4193 (N_4193,N_3340,N_3591);
or U4194 (N_4194,N_3205,N_3266);
and U4195 (N_4195,N_3444,N_3876);
or U4196 (N_4196,N_3391,N_3873);
or U4197 (N_4197,N_3727,N_3243);
or U4198 (N_4198,N_3113,N_3858);
nor U4199 (N_4199,N_3752,N_3798);
or U4200 (N_4200,N_3700,N_3621);
or U4201 (N_4201,N_3739,N_3385);
nand U4202 (N_4202,N_3175,N_3435);
and U4203 (N_4203,N_3561,N_3312);
and U4204 (N_4204,N_3754,N_3074);
and U4205 (N_4205,N_3067,N_3914);
and U4206 (N_4206,N_3447,N_3536);
or U4207 (N_4207,N_3660,N_3375);
xnor U4208 (N_4208,N_3911,N_3011);
nor U4209 (N_4209,N_3736,N_3630);
nor U4210 (N_4210,N_3125,N_3839);
or U4211 (N_4211,N_3415,N_3893);
nor U4212 (N_4212,N_3991,N_3283);
or U4213 (N_4213,N_3090,N_3862);
nor U4214 (N_4214,N_3384,N_3800);
nand U4215 (N_4215,N_3281,N_3617);
or U4216 (N_4216,N_3018,N_3901);
nor U4217 (N_4217,N_3029,N_3499);
and U4218 (N_4218,N_3857,N_3946);
nand U4219 (N_4219,N_3716,N_3260);
nor U4220 (N_4220,N_3117,N_3721);
nand U4221 (N_4221,N_3497,N_3525);
nand U4222 (N_4222,N_3982,N_3437);
nand U4223 (N_4223,N_3855,N_3769);
and U4224 (N_4224,N_3928,N_3383);
and U4225 (N_4225,N_3418,N_3091);
or U4226 (N_4226,N_3409,N_3796);
nor U4227 (N_4227,N_3603,N_3026);
or U4228 (N_4228,N_3146,N_3234);
or U4229 (N_4229,N_3547,N_3593);
and U4230 (N_4230,N_3215,N_3239);
nor U4231 (N_4231,N_3710,N_3844);
and U4232 (N_4232,N_3824,N_3468);
or U4233 (N_4233,N_3629,N_3997);
or U4234 (N_4234,N_3517,N_3833);
and U4235 (N_4235,N_3035,N_3190);
and U4236 (N_4236,N_3988,N_3270);
nand U4237 (N_4237,N_3979,N_3867);
nor U4238 (N_4238,N_3424,N_3324);
and U4239 (N_4239,N_3095,N_3293);
or U4240 (N_4240,N_3799,N_3361);
nand U4241 (N_4241,N_3374,N_3860);
and U4242 (N_4242,N_3359,N_3778);
xnor U4243 (N_4243,N_3273,N_3193);
nor U4244 (N_4244,N_3141,N_3701);
or U4245 (N_4245,N_3083,N_3159);
or U4246 (N_4246,N_3856,N_3331);
and U4247 (N_4247,N_3456,N_3508);
and U4248 (N_4248,N_3284,N_3612);
nand U4249 (N_4249,N_3134,N_3419);
and U4250 (N_4250,N_3212,N_3177);
nand U4251 (N_4251,N_3445,N_3964);
nor U4252 (N_4252,N_3672,N_3319);
nor U4253 (N_4253,N_3601,N_3921);
nand U4254 (N_4254,N_3278,N_3647);
xor U4255 (N_4255,N_3610,N_3747);
nor U4256 (N_4256,N_3852,N_3157);
or U4257 (N_4257,N_3724,N_3924);
or U4258 (N_4258,N_3358,N_3483);
nand U4259 (N_4259,N_3533,N_3254);
nor U4260 (N_4260,N_3756,N_3720);
nor U4261 (N_4261,N_3549,N_3066);
nand U4262 (N_4262,N_3474,N_3514);
or U4263 (N_4263,N_3761,N_3966);
and U4264 (N_4264,N_3993,N_3607);
nand U4265 (N_4265,N_3280,N_3509);
nand U4266 (N_4266,N_3155,N_3088);
nand U4267 (N_4267,N_3102,N_3793);
nor U4268 (N_4268,N_3129,N_3597);
or U4269 (N_4269,N_3526,N_3282);
nor U4270 (N_4270,N_3399,N_3771);
nand U4271 (N_4271,N_3013,N_3534);
and U4272 (N_4272,N_3398,N_3455);
nand U4273 (N_4273,N_3895,N_3706);
nor U4274 (N_4274,N_3838,N_3523);
or U4275 (N_4275,N_3245,N_3344);
and U4276 (N_4276,N_3448,N_3868);
nand U4277 (N_4277,N_3936,N_3635);
and U4278 (N_4278,N_3196,N_3320);
nand U4279 (N_4279,N_3182,N_3410);
nand U4280 (N_4280,N_3668,N_3037);
or U4281 (N_4281,N_3350,N_3652);
nand U4282 (N_4282,N_3139,N_3371);
and U4283 (N_4283,N_3339,N_3622);
nor U4284 (N_4284,N_3841,N_3454);
nand U4285 (N_4285,N_3765,N_3808);
nand U4286 (N_4286,N_3020,N_3315);
nor U4287 (N_4287,N_3039,N_3705);
nand U4288 (N_4288,N_3691,N_3202);
nand U4289 (N_4289,N_3831,N_3187);
nand U4290 (N_4290,N_3251,N_3145);
nand U4291 (N_4291,N_3213,N_3658);
or U4292 (N_4292,N_3913,N_3197);
or U4293 (N_4293,N_3249,N_3242);
and U4294 (N_4294,N_3697,N_3625);
nand U4295 (N_4295,N_3478,N_3493);
nand U4296 (N_4296,N_3269,N_3122);
or U4297 (N_4297,N_3211,N_3489);
and U4298 (N_4298,N_3184,N_3926);
nand U4299 (N_4299,N_3758,N_3958);
or U4300 (N_4300,N_3322,N_3743);
and U4301 (N_4301,N_3871,N_3708);
nor U4302 (N_4302,N_3823,N_3929);
nor U4303 (N_4303,N_3089,N_3598);
or U4304 (N_4304,N_3772,N_3431);
xor U4305 (N_4305,N_3695,N_3428);
xor U4306 (N_4306,N_3055,N_3174);
nor U4307 (N_4307,N_3646,N_3709);
nand U4308 (N_4308,N_3539,N_3680);
or U4309 (N_4309,N_3043,N_3495);
nand U4310 (N_4310,N_3683,N_3932);
nor U4311 (N_4311,N_3849,N_3559);
nor U4312 (N_4312,N_3734,N_3265);
nand U4313 (N_4313,N_3093,N_3579);
nor U4314 (N_4314,N_3959,N_3696);
nand U4315 (N_4315,N_3933,N_3677);
nor U4316 (N_4316,N_3775,N_3963);
or U4317 (N_4317,N_3619,N_3570);
nor U4318 (N_4318,N_3780,N_3845);
nor U4319 (N_4319,N_3438,N_3180);
nand U4320 (N_4320,N_3471,N_3803);
and U4321 (N_4321,N_3588,N_3132);
or U4322 (N_4322,N_3381,N_3684);
or U4323 (N_4323,N_3010,N_3181);
or U4324 (N_4324,N_3268,N_3667);
nor U4325 (N_4325,N_3224,N_3298);
or U4326 (N_4326,N_3288,N_3994);
nand U4327 (N_4327,N_3531,N_3870);
and U4328 (N_4328,N_3087,N_3490);
or U4329 (N_4329,N_3425,N_3968);
nor U4330 (N_4330,N_3401,N_3600);
nand U4331 (N_4331,N_3967,N_3267);
or U4332 (N_4332,N_3156,N_3031);
or U4333 (N_4333,N_3296,N_3183);
xor U4334 (N_4334,N_3306,N_3430);
nor U4335 (N_4335,N_3501,N_3712);
nand U4336 (N_4336,N_3120,N_3717);
nand U4337 (N_4337,N_3908,N_3516);
or U4338 (N_4338,N_3198,N_3025);
nor U4339 (N_4339,N_3052,N_3931);
or U4340 (N_4340,N_3813,N_3098);
and U4341 (N_4341,N_3235,N_3961);
nand U4342 (N_4342,N_3069,N_3433);
and U4343 (N_4343,N_3004,N_3613);
and U4344 (N_4344,N_3511,N_3620);
or U4345 (N_4345,N_3728,N_3757);
nand U4346 (N_4346,N_3826,N_3166);
nor U4347 (N_4347,N_3515,N_3564);
nor U4348 (N_4348,N_3986,N_3176);
nand U4349 (N_4349,N_3566,N_3545);
nor U4350 (N_4350,N_3611,N_3204);
or U4351 (N_4351,N_3643,N_3834);
nor U4352 (N_4352,N_3733,N_3552);
nand U4353 (N_4353,N_3480,N_3195);
or U4354 (N_4354,N_3335,N_3165);
nor U4355 (N_4355,N_3290,N_3632);
or U4356 (N_4356,N_3112,N_3889);
or U4357 (N_4357,N_3631,N_3400);
nand U4358 (N_4358,N_3115,N_3084);
and U4359 (N_4359,N_3070,N_3542);
nor U4360 (N_4360,N_3302,N_3692);
nor U4361 (N_4361,N_3952,N_3779);
and U4362 (N_4362,N_3228,N_3355);
nand U4363 (N_4363,N_3786,N_3295);
nand U4364 (N_4364,N_3068,N_3427);
xnor U4365 (N_4365,N_3143,N_3731);
and U4366 (N_4366,N_3292,N_3220);
and U4367 (N_4367,N_3751,N_3104);
and U4368 (N_4368,N_3106,N_3365);
nor U4369 (N_4369,N_3879,N_3346);
and U4370 (N_4370,N_3412,N_3587);
nor U4371 (N_4371,N_3686,N_3737);
or U4372 (N_4372,N_3417,N_3949);
nor U4373 (N_4373,N_3484,N_3527);
and U4374 (N_4374,N_3149,N_3470);
nor U4375 (N_4375,N_3642,N_3503);
nor U4376 (N_4376,N_3318,N_3894);
or U4377 (N_4377,N_3274,N_3097);
nand U4378 (N_4378,N_3837,N_3624);
or U4379 (N_4379,N_3050,N_3082);
nor U4380 (N_4380,N_3049,N_3164);
and U4381 (N_4381,N_3767,N_3863);
or U4382 (N_4382,N_3902,N_3645);
or U4383 (N_4383,N_3054,N_3878);
nor U4384 (N_4384,N_3553,N_3294);
nand U4385 (N_4385,N_3804,N_3491);
nand U4386 (N_4386,N_3877,N_3262);
and U4387 (N_4387,N_3836,N_3649);
and U4388 (N_4388,N_3922,N_3207);
nor U4389 (N_4389,N_3802,N_3276);
and U4390 (N_4390,N_3694,N_3605);
nand U4391 (N_4391,N_3396,N_3866);
nor U4392 (N_4392,N_3436,N_3168);
nand U4393 (N_4393,N_3618,N_3334);
or U4394 (N_4394,N_3927,N_3231);
nor U4395 (N_4395,N_3861,N_3073);
nand U4396 (N_4396,N_3047,N_3842);
nor U4397 (N_4397,N_3865,N_3580);
nand U4398 (N_4398,N_3114,N_3308);
and U4399 (N_4399,N_3051,N_3633);
or U4400 (N_4400,N_3060,N_3015);
and U4401 (N_4401,N_3944,N_3405);
nor U4402 (N_4402,N_3188,N_3675);
and U4403 (N_4403,N_3222,N_3965);
or U4404 (N_4404,N_3891,N_3912);
xnor U4405 (N_4405,N_3264,N_3380);
xnor U4406 (N_4406,N_3307,N_3467);
or U4407 (N_4407,N_3820,N_3465);
or U4408 (N_4408,N_3030,N_3653);
or U4409 (N_4409,N_3881,N_3109);
or U4410 (N_4410,N_3975,N_3434);
and U4411 (N_4411,N_3443,N_3206);
or U4412 (N_4412,N_3905,N_3707);
or U4413 (N_4413,N_3532,N_3540);
nand U4414 (N_4414,N_3451,N_3989);
or U4415 (N_4415,N_3577,N_3225);
nor U4416 (N_4416,N_3776,N_3167);
or U4417 (N_4417,N_3583,N_3171);
or U4418 (N_4418,N_3678,N_3762);
xor U4419 (N_4419,N_3351,N_3584);
or U4420 (N_4420,N_3151,N_3356);
and U4421 (N_4421,N_3519,N_3218);
and U4422 (N_4422,N_3693,N_3768);
nor U4423 (N_4423,N_3329,N_3655);
nor U4424 (N_4424,N_3229,N_3722);
or U4425 (N_4425,N_3341,N_3492);
nor U4426 (N_4426,N_3481,N_3664);
and U4427 (N_4427,N_3079,N_3147);
nand U4428 (N_4428,N_3153,N_3970);
and U4429 (N_4429,N_3321,N_3809);
or U4430 (N_4430,N_3233,N_3058);
or U4431 (N_4431,N_3869,N_3971);
or U4432 (N_4432,N_3472,N_3546);
or U4433 (N_4433,N_3628,N_3792);
nor U4434 (N_4434,N_3045,N_3781);
xor U4435 (N_4435,N_3150,N_3945);
or U4436 (N_4436,N_3910,N_3036);
or U4437 (N_4437,N_3900,N_3585);
or U4438 (N_4438,N_3671,N_3934);
and U4439 (N_4439,N_3395,N_3663);
xnor U4440 (N_4440,N_3851,N_3850);
nor U4441 (N_4441,N_3287,N_3641);
nand U4442 (N_4442,N_3960,N_3918);
xor U4443 (N_4443,N_3898,N_3892);
nor U4444 (N_4444,N_3797,N_3665);
nor U4445 (N_4445,N_3111,N_3300);
nand U4446 (N_4446,N_3791,N_3750);
nand U4447 (N_4447,N_3373,N_3502);
or U4448 (N_4448,N_3573,N_3277);
nand U4449 (N_4449,N_3247,N_3565);
or U4450 (N_4450,N_3732,N_3788);
or U4451 (N_4451,N_3560,N_3789);
nand U4452 (N_4452,N_3034,N_3987);
nand U4453 (N_4453,N_3185,N_3330);
nand U4454 (N_4454,N_3086,N_3389);
or U4455 (N_4455,N_3237,N_3782);
nand U4456 (N_4456,N_3003,N_3673);
nand U4457 (N_4457,N_3366,N_3289);
nor U4458 (N_4458,N_3370,N_3524);
or U4459 (N_4459,N_3661,N_3760);
nand U4460 (N_4460,N_3770,N_3890);
or U4461 (N_4461,N_3699,N_3581);
nand U4462 (N_4462,N_3897,N_3421);
or U4463 (N_4463,N_3240,N_3189);
nor U4464 (N_4464,N_3023,N_3977);
nand U4465 (N_4465,N_3880,N_3723);
and U4466 (N_4466,N_3640,N_3816);
or U4467 (N_4467,N_3528,N_3783);
nor U4468 (N_4468,N_3530,N_3162);
and U4469 (N_4469,N_3888,N_3336);
or U4470 (N_4470,N_3449,N_3368);
xnor U4471 (N_4471,N_3648,N_3817);
nor U4472 (N_4472,N_3785,N_3567);
nand U4473 (N_4473,N_3615,N_3787);
xnor U4474 (N_4474,N_3158,N_3219);
and U4475 (N_4475,N_3094,N_3742);
or U4476 (N_4476,N_3226,N_3494);
and U4477 (N_4477,N_3429,N_3209);
or U4478 (N_4478,N_3689,N_3556);
nand U4479 (N_4479,N_3847,N_3749);
and U4480 (N_4480,N_3925,N_3650);
and U4481 (N_4481,N_3075,N_3317);
nand U4482 (N_4482,N_3719,N_3586);
nor U4483 (N_4483,N_3271,N_3367);
or U4484 (N_4484,N_3575,N_3906);
nor U4485 (N_4485,N_3596,N_3957);
and U4486 (N_4486,N_3930,N_3688);
nor U4487 (N_4487,N_3522,N_3238);
and U4488 (N_4488,N_3126,N_3133);
xnor U4489 (N_4489,N_3103,N_3021);
nand U4490 (N_4490,N_3450,N_3099);
nor U4491 (N_4491,N_3687,N_3446);
nor U4492 (N_4492,N_3711,N_3253);
and U4493 (N_4493,N_3602,N_3457);
and U4494 (N_4494,N_3574,N_3221);
nor U4495 (N_4495,N_3349,N_3822);
and U4496 (N_4496,N_3903,N_3053);
and U4497 (N_4497,N_3009,N_3843);
nor U4498 (N_4498,N_3983,N_3044);
or U4499 (N_4499,N_3275,N_3272);
nor U4500 (N_4500,N_3195,N_3291);
or U4501 (N_4501,N_3882,N_3683);
or U4502 (N_4502,N_3418,N_3498);
nand U4503 (N_4503,N_3777,N_3420);
nor U4504 (N_4504,N_3720,N_3618);
and U4505 (N_4505,N_3322,N_3764);
nand U4506 (N_4506,N_3885,N_3518);
or U4507 (N_4507,N_3629,N_3153);
nor U4508 (N_4508,N_3325,N_3298);
and U4509 (N_4509,N_3834,N_3414);
nor U4510 (N_4510,N_3928,N_3778);
or U4511 (N_4511,N_3479,N_3884);
or U4512 (N_4512,N_3599,N_3875);
or U4513 (N_4513,N_3578,N_3038);
or U4514 (N_4514,N_3707,N_3979);
or U4515 (N_4515,N_3494,N_3111);
nor U4516 (N_4516,N_3178,N_3639);
nor U4517 (N_4517,N_3726,N_3693);
nand U4518 (N_4518,N_3778,N_3473);
or U4519 (N_4519,N_3877,N_3835);
nand U4520 (N_4520,N_3180,N_3651);
nand U4521 (N_4521,N_3189,N_3482);
xnor U4522 (N_4522,N_3098,N_3748);
nand U4523 (N_4523,N_3617,N_3406);
or U4524 (N_4524,N_3176,N_3108);
or U4525 (N_4525,N_3442,N_3619);
nor U4526 (N_4526,N_3905,N_3904);
nor U4527 (N_4527,N_3133,N_3197);
or U4528 (N_4528,N_3093,N_3495);
or U4529 (N_4529,N_3604,N_3147);
or U4530 (N_4530,N_3745,N_3140);
nand U4531 (N_4531,N_3260,N_3237);
and U4532 (N_4532,N_3119,N_3231);
nor U4533 (N_4533,N_3797,N_3474);
and U4534 (N_4534,N_3211,N_3907);
xnor U4535 (N_4535,N_3165,N_3976);
nor U4536 (N_4536,N_3658,N_3531);
and U4537 (N_4537,N_3149,N_3992);
or U4538 (N_4538,N_3256,N_3588);
nand U4539 (N_4539,N_3604,N_3111);
or U4540 (N_4540,N_3354,N_3342);
nor U4541 (N_4541,N_3115,N_3734);
xor U4542 (N_4542,N_3479,N_3379);
or U4543 (N_4543,N_3631,N_3258);
or U4544 (N_4544,N_3898,N_3782);
nor U4545 (N_4545,N_3478,N_3961);
or U4546 (N_4546,N_3561,N_3233);
and U4547 (N_4547,N_3914,N_3545);
nor U4548 (N_4548,N_3602,N_3478);
or U4549 (N_4549,N_3246,N_3617);
and U4550 (N_4550,N_3438,N_3668);
nand U4551 (N_4551,N_3001,N_3885);
nand U4552 (N_4552,N_3431,N_3906);
nand U4553 (N_4553,N_3606,N_3511);
and U4554 (N_4554,N_3196,N_3293);
nand U4555 (N_4555,N_3790,N_3290);
or U4556 (N_4556,N_3691,N_3721);
and U4557 (N_4557,N_3218,N_3904);
and U4558 (N_4558,N_3119,N_3292);
nand U4559 (N_4559,N_3345,N_3916);
or U4560 (N_4560,N_3090,N_3139);
nand U4561 (N_4561,N_3364,N_3592);
and U4562 (N_4562,N_3048,N_3264);
nor U4563 (N_4563,N_3773,N_3402);
or U4564 (N_4564,N_3988,N_3084);
nand U4565 (N_4565,N_3503,N_3576);
and U4566 (N_4566,N_3164,N_3436);
or U4567 (N_4567,N_3854,N_3560);
nand U4568 (N_4568,N_3415,N_3335);
or U4569 (N_4569,N_3941,N_3213);
and U4570 (N_4570,N_3150,N_3276);
or U4571 (N_4571,N_3792,N_3076);
nor U4572 (N_4572,N_3439,N_3595);
or U4573 (N_4573,N_3081,N_3738);
or U4574 (N_4574,N_3347,N_3343);
nor U4575 (N_4575,N_3212,N_3218);
nor U4576 (N_4576,N_3568,N_3154);
and U4577 (N_4577,N_3067,N_3345);
or U4578 (N_4578,N_3561,N_3151);
and U4579 (N_4579,N_3474,N_3429);
and U4580 (N_4580,N_3617,N_3471);
and U4581 (N_4581,N_3715,N_3085);
nor U4582 (N_4582,N_3631,N_3499);
nor U4583 (N_4583,N_3262,N_3496);
nand U4584 (N_4584,N_3845,N_3131);
nand U4585 (N_4585,N_3111,N_3951);
xnor U4586 (N_4586,N_3000,N_3387);
and U4587 (N_4587,N_3779,N_3221);
nor U4588 (N_4588,N_3358,N_3417);
and U4589 (N_4589,N_3527,N_3958);
and U4590 (N_4590,N_3436,N_3826);
nand U4591 (N_4591,N_3574,N_3861);
or U4592 (N_4592,N_3351,N_3393);
nor U4593 (N_4593,N_3363,N_3073);
and U4594 (N_4594,N_3710,N_3787);
nor U4595 (N_4595,N_3590,N_3342);
nand U4596 (N_4596,N_3692,N_3805);
or U4597 (N_4597,N_3453,N_3654);
nand U4598 (N_4598,N_3506,N_3335);
nand U4599 (N_4599,N_3927,N_3913);
or U4600 (N_4600,N_3255,N_3364);
and U4601 (N_4601,N_3480,N_3529);
nand U4602 (N_4602,N_3566,N_3955);
nor U4603 (N_4603,N_3799,N_3834);
or U4604 (N_4604,N_3723,N_3381);
nor U4605 (N_4605,N_3926,N_3079);
and U4606 (N_4606,N_3740,N_3390);
or U4607 (N_4607,N_3368,N_3533);
and U4608 (N_4608,N_3241,N_3019);
nand U4609 (N_4609,N_3793,N_3702);
nor U4610 (N_4610,N_3804,N_3814);
and U4611 (N_4611,N_3263,N_3641);
and U4612 (N_4612,N_3153,N_3630);
nand U4613 (N_4613,N_3206,N_3573);
or U4614 (N_4614,N_3717,N_3538);
and U4615 (N_4615,N_3089,N_3143);
or U4616 (N_4616,N_3211,N_3954);
nand U4617 (N_4617,N_3000,N_3983);
nor U4618 (N_4618,N_3319,N_3255);
or U4619 (N_4619,N_3397,N_3016);
nand U4620 (N_4620,N_3874,N_3682);
nor U4621 (N_4621,N_3272,N_3457);
or U4622 (N_4622,N_3490,N_3273);
or U4623 (N_4623,N_3515,N_3386);
nor U4624 (N_4624,N_3393,N_3177);
and U4625 (N_4625,N_3030,N_3120);
or U4626 (N_4626,N_3019,N_3276);
nor U4627 (N_4627,N_3184,N_3682);
and U4628 (N_4628,N_3549,N_3337);
or U4629 (N_4629,N_3213,N_3437);
nand U4630 (N_4630,N_3237,N_3717);
nor U4631 (N_4631,N_3104,N_3510);
nor U4632 (N_4632,N_3078,N_3862);
nand U4633 (N_4633,N_3879,N_3440);
nor U4634 (N_4634,N_3854,N_3528);
xor U4635 (N_4635,N_3716,N_3060);
or U4636 (N_4636,N_3982,N_3054);
or U4637 (N_4637,N_3867,N_3358);
nor U4638 (N_4638,N_3295,N_3859);
and U4639 (N_4639,N_3648,N_3295);
and U4640 (N_4640,N_3840,N_3422);
nand U4641 (N_4641,N_3993,N_3529);
nor U4642 (N_4642,N_3014,N_3916);
and U4643 (N_4643,N_3206,N_3093);
or U4644 (N_4644,N_3068,N_3752);
nor U4645 (N_4645,N_3801,N_3772);
or U4646 (N_4646,N_3760,N_3001);
or U4647 (N_4647,N_3334,N_3316);
and U4648 (N_4648,N_3900,N_3496);
nor U4649 (N_4649,N_3188,N_3027);
nand U4650 (N_4650,N_3859,N_3170);
and U4651 (N_4651,N_3230,N_3801);
xor U4652 (N_4652,N_3802,N_3538);
or U4653 (N_4653,N_3184,N_3592);
nand U4654 (N_4654,N_3267,N_3339);
or U4655 (N_4655,N_3699,N_3637);
and U4656 (N_4656,N_3651,N_3465);
and U4657 (N_4657,N_3011,N_3805);
nand U4658 (N_4658,N_3614,N_3967);
nand U4659 (N_4659,N_3213,N_3027);
and U4660 (N_4660,N_3151,N_3895);
or U4661 (N_4661,N_3117,N_3453);
and U4662 (N_4662,N_3539,N_3129);
and U4663 (N_4663,N_3238,N_3511);
nand U4664 (N_4664,N_3188,N_3171);
or U4665 (N_4665,N_3820,N_3882);
or U4666 (N_4666,N_3690,N_3890);
and U4667 (N_4667,N_3057,N_3734);
and U4668 (N_4668,N_3564,N_3483);
nand U4669 (N_4669,N_3951,N_3480);
or U4670 (N_4670,N_3189,N_3902);
and U4671 (N_4671,N_3804,N_3367);
nor U4672 (N_4672,N_3538,N_3625);
or U4673 (N_4673,N_3933,N_3508);
or U4674 (N_4674,N_3681,N_3465);
nand U4675 (N_4675,N_3814,N_3293);
or U4676 (N_4676,N_3670,N_3227);
nand U4677 (N_4677,N_3294,N_3307);
and U4678 (N_4678,N_3023,N_3069);
or U4679 (N_4679,N_3822,N_3663);
xnor U4680 (N_4680,N_3949,N_3854);
nand U4681 (N_4681,N_3222,N_3396);
nor U4682 (N_4682,N_3694,N_3349);
or U4683 (N_4683,N_3048,N_3804);
or U4684 (N_4684,N_3710,N_3488);
nor U4685 (N_4685,N_3984,N_3972);
nor U4686 (N_4686,N_3594,N_3429);
and U4687 (N_4687,N_3434,N_3423);
or U4688 (N_4688,N_3689,N_3500);
or U4689 (N_4689,N_3095,N_3989);
or U4690 (N_4690,N_3153,N_3062);
or U4691 (N_4691,N_3943,N_3053);
and U4692 (N_4692,N_3209,N_3234);
nor U4693 (N_4693,N_3323,N_3495);
nand U4694 (N_4694,N_3227,N_3075);
nor U4695 (N_4695,N_3715,N_3691);
nor U4696 (N_4696,N_3124,N_3182);
xor U4697 (N_4697,N_3930,N_3368);
nand U4698 (N_4698,N_3588,N_3768);
or U4699 (N_4699,N_3358,N_3070);
nor U4700 (N_4700,N_3933,N_3867);
and U4701 (N_4701,N_3377,N_3236);
nand U4702 (N_4702,N_3425,N_3562);
nor U4703 (N_4703,N_3242,N_3676);
nor U4704 (N_4704,N_3674,N_3946);
nand U4705 (N_4705,N_3608,N_3264);
nor U4706 (N_4706,N_3017,N_3081);
nor U4707 (N_4707,N_3653,N_3555);
nor U4708 (N_4708,N_3117,N_3025);
nor U4709 (N_4709,N_3800,N_3005);
or U4710 (N_4710,N_3945,N_3170);
or U4711 (N_4711,N_3464,N_3572);
nor U4712 (N_4712,N_3158,N_3431);
and U4713 (N_4713,N_3198,N_3646);
nor U4714 (N_4714,N_3880,N_3556);
xnor U4715 (N_4715,N_3119,N_3332);
and U4716 (N_4716,N_3820,N_3719);
or U4717 (N_4717,N_3984,N_3640);
or U4718 (N_4718,N_3891,N_3752);
nand U4719 (N_4719,N_3111,N_3933);
nand U4720 (N_4720,N_3954,N_3205);
nand U4721 (N_4721,N_3940,N_3640);
and U4722 (N_4722,N_3387,N_3623);
nor U4723 (N_4723,N_3872,N_3325);
nand U4724 (N_4724,N_3291,N_3723);
or U4725 (N_4725,N_3917,N_3608);
nor U4726 (N_4726,N_3426,N_3126);
nor U4727 (N_4727,N_3089,N_3086);
or U4728 (N_4728,N_3532,N_3725);
or U4729 (N_4729,N_3373,N_3493);
or U4730 (N_4730,N_3808,N_3260);
nand U4731 (N_4731,N_3824,N_3715);
and U4732 (N_4732,N_3631,N_3629);
nor U4733 (N_4733,N_3084,N_3302);
or U4734 (N_4734,N_3026,N_3855);
nand U4735 (N_4735,N_3402,N_3014);
and U4736 (N_4736,N_3375,N_3152);
or U4737 (N_4737,N_3746,N_3513);
nand U4738 (N_4738,N_3409,N_3113);
nor U4739 (N_4739,N_3390,N_3399);
or U4740 (N_4740,N_3774,N_3995);
or U4741 (N_4741,N_3235,N_3929);
nor U4742 (N_4742,N_3973,N_3583);
xnor U4743 (N_4743,N_3941,N_3569);
nor U4744 (N_4744,N_3411,N_3522);
nor U4745 (N_4745,N_3928,N_3477);
or U4746 (N_4746,N_3504,N_3943);
nand U4747 (N_4747,N_3767,N_3630);
nand U4748 (N_4748,N_3673,N_3191);
xnor U4749 (N_4749,N_3335,N_3575);
nand U4750 (N_4750,N_3521,N_3016);
or U4751 (N_4751,N_3995,N_3992);
or U4752 (N_4752,N_3039,N_3849);
nand U4753 (N_4753,N_3080,N_3068);
and U4754 (N_4754,N_3441,N_3079);
nand U4755 (N_4755,N_3986,N_3838);
nor U4756 (N_4756,N_3243,N_3696);
nand U4757 (N_4757,N_3031,N_3241);
and U4758 (N_4758,N_3358,N_3945);
xnor U4759 (N_4759,N_3254,N_3203);
nor U4760 (N_4760,N_3143,N_3225);
and U4761 (N_4761,N_3384,N_3225);
and U4762 (N_4762,N_3044,N_3003);
or U4763 (N_4763,N_3313,N_3288);
nor U4764 (N_4764,N_3612,N_3919);
or U4765 (N_4765,N_3034,N_3904);
or U4766 (N_4766,N_3470,N_3600);
nand U4767 (N_4767,N_3995,N_3221);
or U4768 (N_4768,N_3220,N_3327);
and U4769 (N_4769,N_3686,N_3397);
and U4770 (N_4770,N_3841,N_3173);
nand U4771 (N_4771,N_3204,N_3380);
and U4772 (N_4772,N_3152,N_3442);
and U4773 (N_4773,N_3934,N_3806);
xnor U4774 (N_4774,N_3854,N_3895);
or U4775 (N_4775,N_3968,N_3447);
or U4776 (N_4776,N_3962,N_3660);
or U4777 (N_4777,N_3743,N_3890);
nand U4778 (N_4778,N_3123,N_3782);
or U4779 (N_4779,N_3255,N_3175);
nor U4780 (N_4780,N_3969,N_3251);
or U4781 (N_4781,N_3858,N_3104);
and U4782 (N_4782,N_3374,N_3843);
or U4783 (N_4783,N_3789,N_3779);
xor U4784 (N_4784,N_3715,N_3899);
nor U4785 (N_4785,N_3477,N_3208);
nand U4786 (N_4786,N_3706,N_3928);
xor U4787 (N_4787,N_3576,N_3655);
nand U4788 (N_4788,N_3614,N_3776);
nand U4789 (N_4789,N_3209,N_3464);
and U4790 (N_4790,N_3927,N_3687);
or U4791 (N_4791,N_3332,N_3475);
and U4792 (N_4792,N_3003,N_3536);
or U4793 (N_4793,N_3137,N_3011);
nor U4794 (N_4794,N_3454,N_3704);
and U4795 (N_4795,N_3500,N_3905);
nand U4796 (N_4796,N_3364,N_3186);
and U4797 (N_4797,N_3646,N_3730);
or U4798 (N_4798,N_3012,N_3720);
or U4799 (N_4799,N_3662,N_3462);
nand U4800 (N_4800,N_3097,N_3899);
or U4801 (N_4801,N_3647,N_3578);
or U4802 (N_4802,N_3318,N_3329);
nand U4803 (N_4803,N_3168,N_3336);
nor U4804 (N_4804,N_3243,N_3315);
nor U4805 (N_4805,N_3138,N_3238);
nand U4806 (N_4806,N_3783,N_3989);
nor U4807 (N_4807,N_3290,N_3899);
nand U4808 (N_4808,N_3467,N_3823);
and U4809 (N_4809,N_3385,N_3641);
nor U4810 (N_4810,N_3249,N_3082);
and U4811 (N_4811,N_3812,N_3025);
nor U4812 (N_4812,N_3117,N_3941);
or U4813 (N_4813,N_3107,N_3027);
nand U4814 (N_4814,N_3979,N_3785);
nor U4815 (N_4815,N_3693,N_3782);
nor U4816 (N_4816,N_3981,N_3602);
or U4817 (N_4817,N_3527,N_3761);
nand U4818 (N_4818,N_3234,N_3916);
and U4819 (N_4819,N_3397,N_3843);
or U4820 (N_4820,N_3728,N_3407);
or U4821 (N_4821,N_3547,N_3317);
nor U4822 (N_4822,N_3187,N_3546);
or U4823 (N_4823,N_3451,N_3328);
or U4824 (N_4824,N_3851,N_3748);
nand U4825 (N_4825,N_3461,N_3943);
and U4826 (N_4826,N_3860,N_3305);
nor U4827 (N_4827,N_3584,N_3426);
or U4828 (N_4828,N_3553,N_3833);
nor U4829 (N_4829,N_3627,N_3349);
nor U4830 (N_4830,N_3860,N_3538);
or U4831 (N_4831,N_3109,N_3903);
nand U4832 (N_4832,N_3692,N_3325);
nor U4833 (N_4833,N_3585,N_3080);
and U4834 (N_4834,N_3503,N_3127);
or U4835 (N_4835,N_3322,N_3240);
nand U4836 (N_4836,N_3870,N_3566);
or U4837 (N_4837,N_3278,N_3558);
and U4838 (N_4838,N_3159,N_3106);
and U4839 (N_4839,N_3861,N_3558);
and U4840 (N_4840,N_3709,N_3983);
nand U4841 (N_4841,N_3928,N_3569);
nor U4842 (N_4842,N_3182,N_3372);
and U4843 (N_4843,N_3585,N_3337);
nand U4844 (N_4844,N_3562,N_3285);
and U4845 (N_4845,N_3255,N_3421);
or U4846 (N_4846,N_3391,N_3522);
nor U4847 (N_4847,N_3848,N_3611);
or U4848 (N_4848,N_3592,N_3291);
or U4849 (N_4849,N_3497,N_3152);
nand U4850 (N_4850,N_3172,N_3833);
and U4851 (N_4851,N_3373,N_3314);
and U4852 (N_4852,N_3705,N_3159);
and U4853 (N_4853,N_3649,N_3901);
and U4854 (N_4854,N_3115,N_3231);
nor U4855 (N_4855,N_3461,N_3135);
and U4856 (N_4856,N_3789,N_3885);
nor U4857 (N_4857,N_3841,N_3075);
nand U4858 (N_4858,N_3374,N_3508);
nor U4859 (N_4859,N_3537,N_3665);
and U4860 (N_4860,N_3285,N_3174);
nand U4861 (N_4861,N_3363,N_3301);
xnor U4862 (N_4862,N_3799,N_3878);
nand U4863 (N_4863,N_3544,N_3276);
or U4864 (N_4864,N_3079,N_3065);
and U4865 (N_4865,N_3416,N_3667);
and U4866 (N_4866,N_3844,N_3946);
nor U4867 (N_4867,N_3868,N_3759);
xor U4868 (N_4868,N_3535,N_3434);
nand U4869 (N_4869,N_3749,N_3413);
and U4870 (N_4870,N_3621,N_3090);
or U4871 (N_4871,N_3488,N_3327);
nand U4872 (N_4872,N_3658,N_3588);
nor U4873 (N_4873,N_3238,N_3697);
nand U4874 (N_4874,N_3779,N_3974);
and U4875 (N_4875,N_3718,N_3736);
or U4876 (N_4876,N_3607,N_3007);
and U4877 (N_4877,N_3731,N_3850);
nand U4878 (N_4878,N_3877,N_3064);
or U4879 (N_4879,N_3669,N_3274);
nand U4880 (N_4880,N_3946,N_3177);
or U4881 (N_4881,N_3236,N_3237);
and U4882 (N_4882,N_3718,N_3000);
nor U4883 (N_4883,N_3268,N_3067);
nor U4884 (N_4884,N_3441,N_3767);
and U4885 (N_4885,N_3649,N_3071);
xnor U4886 (N_4886,N_3872,N_3885);
nor U4887 (N_4887,N_3573,N_3463);
and U4888 (N_4888,N_3379,N_3042);
nand U4889 (N_4889,N_3987,N_3543);
or U4890 (N_4890,N_3616,N_3491);
xnor U4891 (N_4891,N_3988,N_3804);
nand U4892 (N_4892,N_3472,N_3132);
and U4893 (N_4893,N_3272,N_3724);
nor U4894 (N_4894,N_3241,N_3186);
nor U4895 (N_4895,N_3428,N_3006);
nand U4896 (N_4896,N_3837,N_3879);
nor U4897 (N_4897,N_3954,N_3500);
nor U4898 (N_4898,N_3991,N_3350);
nand U4899 (N_4899,N_3083,N_3347);
nand U4900 (N_4900,N_3494,N_3870);
and U4901 (N_4901,N_3868,N_3289);
nand U4902 (N_4902,N_3770,N_3247);
nand U4903 (N_4903,N_3012,N_3695);
or U4904 (N_4904,N_3489,N_3724);
nand U4905 (N_4905,N_3731,N_3021);
or U4906 (N_4906,N_3637,N_3003);
nand U4907 (N_4907,N_3279,N_3389);
nor U4908 (N_4908,N_3578,N_3226);
nand U4909 (N_4909,N_3452,N_3749);
nor U4910 (N_4910,N_3106,N_3029);
and U4911 (N_4911,N_3433,N_3664);
nor U4912 (N_4912,N_3955,N_3488);
or U4913 (N_4913,N_3553,N_3339);
nor U4914 (N_4914,N_3668,N_3629);
nand U4915 (N_4915,N_3633,N_3289);
or U4916 (N_4916,N_3984,N_3584);
or U4917 (N_4917,N_3387,N_3138);
and U4918 (N_4918,N_3192,N_3553);
or U4919 (N_4919,N_3535,N_3146);
nand U4920 (N_4920,N_3474,N_3253);
nor U4921 (N_4921,N_3878,N_3506);
and U4922 (N_4922,N_3839,N_3911);
or U4923 (N_4923,N_3701,N_3190);
and U4924 (N_4924,N_3687,N_3451);
nor U4925 (N_4925,N_3147,N_3323);
nor U4926 (N_4926,N_3689,N_3935);
and U4927 (N_4927,N_3643,N_3411);
nand U4928 (N_4928,N_3382,N_3923);
nor U4929 (N_4929,N_3822,N_3905);
nand U4930 (N_4930,N_3666,N_3235);
xnor U4931 (N_4931,N_3243,N_3011);
nor U4932 (N_4932,N_3786,N_3664);
and U4933 (N_4933,N_3504,N_3908);
and U4934 (N_4934,N_3842,N_3456);
xnor U4935 (N_4935,N_3444,N_3721);
nand U4936 (N_4936,N_3174,N_3272);
nor U4937 (N_4937,N_3606,N_3826);
xor U4938 (N_4938,N_3181,N_3966);
or U4939 (N_4939,N_3263,N_3976);
and U4940 (N_4940,N_3821,N_3152);
nand U4941 (N_4941,N_3470,N_3444);
nand U4942 (N_4942,N_3588,N_3983);
or U4943 (N_4943,N_3908,N_3019);
and U4944 (N_4944,N_3992,N_3776);
and U4945 (N_4945,N_3165,N_3924);
xnor U4946 (N_4946,N_3653,N_3151);
nand U4947 (N_4947,N_3687,N_3593);
and U4948 (N_4948,N_3623,N_3863);
or U4949 (N_4949,N_3635,N_3169);
nand U4950 (N_4950,N_3464,N_3002);
and U4951 (N_4951,N_3657,N_3006);
nand U4952 (N_4952,N_3893,N_3494);
and U4953 (N_4953,N_3347,N_3401);
nand U4954 (N_4954,N_3522,N_3176);
and U4955 (N_4955,N_3940,N_3259);
and U4956 (N_4956,N_3167,N_3884);
or U4957 (N_4957,N_3264,N_3248);
or U4958 (N_4958,N_3825,N_3795);
nand U4959 (N_4959,N_3246,N_3495);
and U4960 (N_4960,N_3399,N_3731);
nor U4961 (N_4961,N_3785,N_3909);
or U4962 (N_4962,N_3595,N_3801);
nor U4963 (N_4963,N_3308,N_3379);
nand U4964 (N_4964,N_3769,N_3825);
nand U4965 (N_4965,N_3576,N_3501);
nor U4966 (N_4966,N_3835,N_3424);
and U4967 (N_4967,N_3641,N_3090);
or U4968 (N_4968,N_3817,N_3789);
and U4969 (N_4969,N_3419,N_3914);
xnor U4970 (N_4970,N_3589,N_3566);
nor U4971 (N_4971,N_3958,N_3448);
nand U4972 (N_4972,N_3372,N_3625);
nand U4973 (N_4973,N_3331,N_3289);
nor U4974 (N_4974,N_3393,N_3871);
and U4975 (N_4975,N_3701,N_3936);
nand U4976 (N_4976,N_3293,N_3412);
or U4977 (N_4977,N_3531,N_3134);
or U4978 (N_4978,N_3194,N_3674);
or U4979 (N_4979,N_3052,N_3623);
nand U4980 (N_4980,N_3109,N_3451);
and U4981 (N_4981,N_3364,N_3406);
nand U4982 (N_4982,N_3233,N_3326);
and U4983 (N_4983,N_3623,N_3464);
or U4984 (N_4984,N_3400,N_3310);
nand U4985 (N_4985,N_3723,N_3477);
nor U4986 (N_4986,N_3282,N_3359);
nor U4987 (N_4987,N_3188,N_3107);
or U4988 (N_4988,N_3501,N_3856);
and U4989 (N_4989,N_3457,N_3395);
or U4990 (N_4990,N_3843,N_3889);
nor U4991 (N_4991,N_3950,N_3307);
nor U4992 (N_4992,N_3343,N_3679);
nand U4993 (N_4993,N_3183,N_3841);
or U4994 (N_4994,N_3858,N_3254);
nor U4995 (N_4995,N_3181,N_3676);
or U4996 (N_4996,N_3548,N_3969);
and U4997 (N_4997,N_3189,N_3298);
nand U4998 (N_4998,N_3644,N_3304);
and U4999 (N_4999,N_3766,N_3787);
nand UO_0 (O_0,N_4724,N_4628);
nand UO_1 (O_1,N_4579,N_4929);
nand UO_2 (O_2,N_4896,N_4084);
and UO_3 (O_3,N_4024,N_4610);
nor UO_4 (O_4,N_4709,N_4815);
nand UO_5 (O_5,N_4745,N_4742);
nand UO_6 (O_6,N_4324,N_4766);
and UO_7 (O_7,N_4274,N_4032);
and UO_8 (O_8,N_4966,N_4314);
or UO_9 (O_9,N_4465,N_4591);
and UO_10 (O_10,N_4356,N_4537);
nor UO_11 (O_11,N_4076,N_4752);
nand UO_12 (O_12,N_4082,N_4222);
and UO_13 (O_13,N_4906,N_4697);
nand UO_14 (O_14,N_4204,N_4051);
nor UO_15 (O_15,N_4480,N_4382);
nand UO_16 (O_16,N_4509,N_4535);
or UO_17 (O_17,N_4443,N_4009);
and UO_18 (O_18,N_4106,N_4780);
nor UO_19 (O_19,N_4171,N_4835);
and UO_20 (O_20,N_4963,N_4000);
or UO_21 (O_21,N_4345,N_4773);
nand UO_22 (O_22,N_4375,N_4998);
nor UO_23 (O_23,N_4332,N_4034);
nand UO_24 (O_24,N_4823,N_4467);
nand UO_25 (O_25,N_4486,N_4093);
or UO_26 (O_26,N_4978,N_4696);
or UO_27 (O_27,N_4269,N_4042);
nor UO_28 (O_28,N_4622,N_4168);
nand UO_29 (O_29,N_4016,N_4405);
and UO_30 (O_30,N_4525,N_4540);
and UO_31 (O_31,N_4598,N_4720);
nand UO_32 (O_32,N_4897,N_4834);
and UO_33 (O_33,N_4441,N_4312);
nand UO_34 (O_34,N_4526,N_4144);
and UO_35 (O_35,N_4921,N_4840);
xnor UO_36 (O_36,N_4175,N_4505);
nor UO_37 (O_37,N_4160,N_4620);
nand UO_38 (O_38,N_4881,N_4374);
nor UO_39 (O_39,N_4096,N_4939);
nor UO_40 (O_40,N_4006,N_4759);
nand UO_41 (O_41,N_4733,N_4249);
nand UO_42 (O_42,N_4098,N_4933);
and UO_43 (O_43,N_4767,N_4466);
nor UO_44 (O_44,N_4729,N_4296);
or UO_45 (O_45,N_4196,N_4458);
and UO_46 (O_46,N_4420,N_4687);
xnor UO_47 (O_47,N_4642,N_4242);
or UO_48 (O_48,N_4992,N_4271);
and UO_49 (O_49,N_4521,N_4412);
nand UO_50 (O_50,N_4248,N_4627);
or UO_51 (O_51,N_4472,N_4692);
or UO_52 (O_52,N_4967,N_4250);
nand UO_53 (O_53,N_4445,N_4712);
and UO_54 (O_54,N_4119,N_4007);
or UO_55 (O_55,N_4124,N_4403);
and UO_56 (O_56,N_4303,N_4878);
nand UO_57 (O_57,N_4576,N_4865);
nand UO_58 (O_58,N_4680,N_4112);
nand UO_59 (O_59,N_4961,N_4725);
nand UO_60 (O_60,N_4636,N_4109);
nor UO_61 (O_61,N_4859,N_4281);
nor UO_62 (O_62,N_4284,N_4651);
or UO_63 (O_63,N_4463,N_4397);
or UO_64 (O_64,N_4900,N_4727);
xor UO_65 (O_65,N_4691,N_4718);
or UO_66 (O_66,N_4979,N_4965);
or UO_67 (O_67,N_4208,N_4563);
and UO_68 (O_68,N_4512,N_4682);
and UO_69 (O_69,N_4842,N_4765);
nor UO_70 (O_70,N_4056,N_4819);
or UO_71 (O_71,N_4990,N_4442);
nor UO_72 (O_72,N_4934,N_4582);
nor UO_73 (O_73,N_4418,N_4552);
or UO_74 (O_74,N_4581,N_4524);
or UO_75 (O_75,N_4212,N_4510);
and UO_76 (O_76,N_4080,N_4519);
and UO_77 (O_77,N_4241,N_4750);
or UO_78 (O_78,N_4782,N_4984);
nor UO_79 (O_79,N_4050,N_4055);
nand UO_80 (O_80,N_4101,N_4430);
nand UO_81 (O_81,N_4272,N_4370);
nor UO_82 (O_82,N_4203,N_4390);
or UO_83 (O_83,N_4955,N_4327);
nand UO_84 (O_84,N_4191,N_4159);
or UO_85 (O_85,N_4623,N_4536);
and UO_86 (O_86,N_4330,N_4090);
or UO_87 (O_87,N_4947,N_4791);
nor UO_88 (O_88,N_4980,N_4502);
and UO_89 (O_89,N_4679,N_4898);
and UO_90 (O_90,N_4422,N_4528);
or UO_91 (O_91,N_4776,N_4589);
and UO_92 (O_92,N_4221,N_4796);
xnor UO_93 (O_93,N_4938,N_4937);
nand UO_94 (O_94,N_4243,N_4608);
and UO_95 (O_95,N_4460,N_4849);
or UO_96 (O_96,N_4348,N_4760);
and UO_97 (O_97,N_4671,N_4981);
nor UO_98 (O_98,N_4943,N_4029);
nor UO_99 (O_99,N_4038,N_4232);
nor UO_100 (O_100,N_4276,N_4614);
nand UO_101 (O_101,N_4832,N_4468);
or UO_102 (O_102,N_4104,N_4383);
nand UO_103 (O_103,N_4064,N_4654);
or UO_104 (O_104,N_4987,N_4067);
nor UO_105 (O_105,N_4137,N_4360);
nand UO_106 (O_106,N_4731,N_4532);
nand UO_107 (O_107,N_4223,N_4735);
nor UO_108 (O_108,N_4787,N_4806);
and UO_109 (O_109,N_4923,N_4944);
nor UO_110 (O_110,N_4503,N_4349);
nor UO_111 (O_111,N_4863,N_4037);
nor UO_112 (O_112,N_4198,N_4613);
and UO_113 (O_113,N_4170,N_4774);
or UO_114 (O_114,N_4634,N_4117);
and UO_115 (O_115,N_4027,N_4932);
or UO_116 (O_116,N_4139,N_4111);
or UO_117 (O_117,N_4775,N_4376);
nand UO_118 (O_118,N_4647,N_4909);
nand UO_119 (O_119,N_4695,N_4630);
or UO_120 (O_120,N_4877,N_4290);
and UO_121 (O_121,N_4044,N_4131);
or UO_122 (O_122,N_4008,N_4311);
and UO_123 (O_123,N_4942,N_4551);
and UO_124 (O_124,N_4631,N_4533);
and UO_125 (O_125,N_4690,N_4656);
and UO_126 (O_126,N_4761,N_4425);
nor UO_127 (O_127,N_4428,N_4378);
nand UO_128 (O_128,N_4520,N_4740);
nand UO_129 (O_129,N_4141,N_4398);
nor UO_130 (O_130,N_4570,N_4496);
nor UO_131 (O_131,N_4818,N_4910);
nor UO_132 (O_132,N_4522,N_4237);
nor UO_133 (O_133,N_4143,N_4833);
nor UO_134 (O_134,N_4280,N_4188);
or UO_135 (O_135,N_4785,N_4150);
nor UO_136 (O_136,N_4149,N_4229);
and UO_137 (O_137,N_4781,N_4263);
nor UO_138 (O_138,N_4368,N_4297);
and UO_139 (O_139,N_4172,N_4322);
and UO_140 (O_140,N_4798,N_4115);
and UO_141 (O_141,N_4672,N_4257);
or UO_142 (O_142,N_4244,N_4895);
nor UO_143 (O_143,N_4371,N_4077);
and UO_144 (O_144,N_4769,N_4092);
nand UO_145 (O_145,N_4924,N_4635);
nand UO_146 (O_146,N_4207,N_4220);
nor UO_147 (O_147,N_4662,N_4238);
nand UO_148 (O_148,N_4091,N_4005);
nand UO_149 (O_149,N_4351,N_4639);
and UO_150 (O_150,N_4476,N_4268);
nand UO_151 (O_151,N_4538,N_4316);
nor UO_152 (O_152,N_4726,N_4844);
nor UO_153 (O_153,N_4911,N_4231);
or UO_154 (O_154,N_4040,N_4068);
or UO_155 (O_155,N_4811,N_4414);
nor UO_156 (O_156,N_4266,N_4105);
nor UO_157 (O_157,N_4971,N_4621);
and UO_158 (O_158,N_4048,N_4035);
nor UO_159 (O_159,N_4440,N_4797);
nor UO_160 (O_160,N_4617,N_4454);
and UO_161 (O_161,N_4583,N_4573);
and UO_162 (O_162,N_4857,N_4347);
or UO_163 (O_163,N_4210,N_4022);
and UO_164 (O_164,N_4547,N_4683);
nand UO_165 (O_165,N_4291,N_4013);
and UO_166 (O_166,N_4564,N_4380);
and UO_167 (O_167,N_4163,N_4571);
and UO_168 (O_168,N_4194,N_4179);
nand UO_169 (O_169,N_4861,N_4429);
or UO_170 (O_170,N_4883,N_4918);
nor UO_171 (O_171,N_4789,N_4286);
nand UO_172 (O_172,N_4600,N_4173);
and UO_173 (O_173,N_4065,N_4338);
and UO_174 (O_174,N_4554,N_4164);
nor UO_175 (O_175,N_4001,N_4640);
nand UO_176 (O_176,N_4419,N_4036);
or UO_177 (O_177,N_4511,N_4189);
nor UO_178 (O_178,N_4985,N_4255);
nand UO_179 (O_179,N_4523,N_4957);
nand UO_180 (O_180,N_4219,N_4950);
or UO_181 (O_181,N_4206,N_4886);
or UO_182 (O_182,N_4461,N_4108);
and UO_183 (O_183,N_4434,N_4501);
xnor UO_184 (O_184,N_4299,N_4153);
nor UO_185 (O_185,N_4996,N_4282);
and UO_186 (O_186,N_4860,N_4308);
and UO_187 (O_187,N_4756,N_4549);
and UO_188 (O_188,N_4305,N_4795);
and UO_189 (O_189,N_4655,N_4363);
or UO_190 (O_190,N_4328,N_4905);
and UO_191 (O_191,N_4930,N_4026);
or UO_192 (O_192,N_4839,N_4644);
or UO_193 (O_193,N_4748,N_4874);
nor UO_194 (O_194,N_4675,N_4660);
nand UO_195 (O_195,N_4320,N_4753);
or UO_196 (O_196,N_4964,N_4872);
nand UO_197 (O_197,N_4273,N_4416);
nand UO_198 (O_198,N_4894,N_4122);
or UO_199 (O_199,N_4217,N_4252);
nor UO_200 (O_200,N_4135,N_4653);
nor UO_201 (O_201,N_4258,N_4459);
nor UO_202 (O_202,N_4094,N_4670);
xor UO_203 (O_203,N_4875,N_4666);
and UO_204 (O_204,N_4784,N_4293);
or UO_205 (O_205,N_4783,N_4058);
nor UO_206 (O_206,N_4810,N_4855);
and UO_207 (O_207,N_4542,N_4728);
or UO_208 (O_208,N_4490,N_4593);
and UO_209 (O_209,N_4663,N_4306);
or UO_210 (O_210,N_4086,N_4764);
and UO_211 (O_211,N_4071,N_4821);
or UO_212 (O_212,N_4128,N_4605);
or UO_213 (O_213,N_4344,N_4073);
nor UO_214 (O_214,N_4667,N_4464);
and UO_215 (O_215,N_4471,N_4134);
nand UO_216 (O_216,N_4313,N_4919);
or UO_217 (O_217,N_4214,N_4566);
nand UO_218 (O_218,N_4688,N_4657);
nand UO_219 (O_219,N_4121,N_4130);
nor UO_220 (O_220,N_4396,N_4705);
or UO_221 (O_221,N_4394,N_4226);
nor UO_222 (O_222,N_4972,N_4952);
nand UO_223 (O_223,N_4777,N_4719);
nand UO_224 (O_224,N_4014,N_4550);
nor UO_225 (O_225,N_4018,N_4908);
nor UO_226 (O_226,N_4711,N_4125);
and UO_227 (O_227,N_4145,N_4643);
nor UO_228 (O_228,N_4493,N_4674);
nand UO_229 (O_229,N_4668,N_4235);
and UO_230 (O_230,N_4133,N_4562);
nor UO_231 (O_231,N_4424,N_4456);
nand UO_232 (O_232,N_4354,N_4224);
nand UO_233 (O_233,N_4702,N_4066);
nand UO_234 (O_234,N_4181,N_4358);
and UO_235 (O_235,N_4070,N_4295);
and UO_236 (O_236,N_4063,N_4757);
and UO_237 (O_237,N_4178,N_4127);
or UO_238 (O_238,N_4515,N_4176);
nand UO_239 (O_239,N_4514,N_4028);
nand UO_240 (O_240,N_4236,N_4954);
or UO_241 (O_241,N_4402,N_4030);
nand UO_242 (O_242,N_4645,N_4555);
and UO_243 (O_243,N_4851,N_4078);
nor UO_244 (O_244,N_4548,N_4021);
nand UO_245 (O_245,N_4300,N_4880);
nand UO_246 (O_246,N_4734,N_4342);
and UO_247 (O_247,N_4132,N_4033);
nand UO_248 (O_248,N_4110,N_4816);
nor UO_249 (O_249,N_4543,N_4218);
or UO_250 (O_250,N_4448,N_4357);
nand UO_251 (O_251,N_4853,N_4199);
or UO_252 (O_252,N_4262,N_4335);
nor UO_253 (O_253,N_4969,N_4618);
or UO_254 (O_254,N_4499,N_4343);
nor UO_255 (O_255,N_4365,N_4407);
or UO_256 (O_256,N_4722,N_4304);
nor UO_257 (O_257,N_4432,N_4917);
and UO_258 (O_258,N_4158,N_4808);
nor UO_259 (O_259,N_4129,N_4891);
nor UO_260 (O_260,N_4567,N_4513);
nand UO_261 (O_261,N_4253,N_4156);
nand UO_262 (O_262,N_4377,N_4935);
xnor UO_263 (O_263,N_4632,N_4928);
nand UO_264 (O_264,N_4245,N_4045);
or UO_265 (O_265,N_4444,N_4417);
nand UO_266 (O_266,N_4557,N_4053);
or UO_267 (O_267,N_4556,N_4439);
and UO_268 (O_268,N_4638,N_4577);
nor UO_269 (O_269,N_4041,N_4624);
nand UO_270 (O_270,N_4813,N_4062);
nand UO_271 (O_271,N_4807,N_4915);
nand UO_272 (O_272,N_4707,N_4400);
nand UO_273 (O_273,N_4546,N_4019);
nor UO_274 (O_274,N_4677,N_4060);
nor UO_275 (O_275,N_4958,N_4993);
and UO_276 (O_276,N_4267,N_4912);
nor UO_277 (O_277,N_4604,N_4580);
and UO_278 (O_278,N_4177,N_4081);
nand UO_279 (O_279,N_4749,N_4870);
and UO_280 (O_280,N_4612,N_4658);
xor UO_281 (O_281,N_4633,N_4146);
or UO_282 (O_282,N_4113,N_4003);
nor UO_283 (O_283,N_4353,N_4446);
xor UO_284 (O_284,N_4778,N_4002);
or UO_285 (O_285,N_4453,N_4820);
and UO_286 (O_286,N_4824,N_4099);
or UO_287 (O_287,N_4061,N_4369);
or UO_288 (O_288,N_4350,N_4504);
nor UO_289 (O_289,N_4879,N_4885);
and UO_290 (O_290,N_4602,N_4846);
and UO_291 (O_291,N_4721,N_4495);
and UO_292 (O_292,N_4799,N_4559);
nor UO_293 (O_293,N_4346,N_4333);
nand UO_294 (O_294,N_4867,N_4619);
nand UO_295 (O_295,N_4603,N_4661);
or UO_296 (O_296,N_4126,N_4020);
or UO_297 (O_297,N_4531,N_4743);
nor UO_298 (O_298,N_4801,N_4052);
or UO_299 (O_299,N_4287,N_4072);
nor UO_300 (O_300,N_4039,N_4926);
nor UO_301 (O_301,N_4664,N_4195);
xor UO_302 (O_302,N_4057,N_4481);
nand UO_303 (O_303,N_4334,N_4574);
and UO_304 (O_304,N_4936,N_4366);
and UO_305 (O_305,N_4254,N_4873);
nand UO_306 (O_306,N_4046,N_4482);
nand UO_307 (O_307,N_4889,N_4234);
xnor UO_308 (O_308,N_4951,N_4578);
nand UO_309 (O_309,N_4478,N_4585);
nor UO_310 (O_310,N_4829,N_4703);
or UO_311 (O_311,N_4892,N_4152);
or UO_312 (O_312,N_4116,N_4771);
or UO_313 (O_313,N_4595,N_4858);
and UO_314 (O_314,N_4736,N_4922);
nand UO_315 (O_315,N_4491,N_4364);
nor UO_316 (O_316,N_4059,N_4800);
and UO_317 (O_317,N_4148,N_4315);
nand UO_318 (O_318,N_4341,N_4541);
and UO_319 (O_319,N_4848,N_4601);
nand UO_320 (O_320,N_4261,N_4278);
nor UO_321 (O_321,N_4869,N_4715);
or UO_322 (O_322,N_4893,N_4864);
xor UO_323 (O_323,N_4385,N_4592);
xnor UO_324 (O_324,N_4372,N_4903);
or UO_325 (O_325,N_4450,N_4588);
nand UO_326 (O_326,N_4686,N_4292);
or UO_327 (O_327,N_4830,N_4714);
nand UO_328 (O_328,N_4770,N_4568);
and UO_329 (O_329,N_4850,N_4483);
and UO_330 (O_330,N_4427,N_4455);
and UO_331 (O_331,N_4960,N_4545);
and UO_332 (O_332,N_4404,N_4659);
nor UO_333 (O_333,N_4976,N_4590);
nand UO_334 (O_334,N_4862,N_4747);
nor UO_335 (O_335,N_4899,N_4594);
and UO_336 (O_336,N_4946,N_4596);
nor UO_337 (O_337,N_4275,N_4890);
nand UO_338 (O_338,N_4487,N_4136);
nand UO_339 (O_339,N_4488,N_4956);
or UO_340 (O_340,N_4948,N_4805);
or UO_341 (O_341,N_4560,N_4393);
and UO_342 (O_342,N_4907,N_4211);
nand UO_343 (O_343,N_4768,N_4251);
and UO_344 (O_344,N_4216,N_4866);
or UO_345 (O_345,N_4277,N_4240);
nand UO_346 (O_346,N_4561,N_4831);
or UO_347 (O_347,N_4569,N_4423);
and UO_348 (O_348,N_4401,N_4916);
nor UO_349 (O_349,N_4882,N_4751);
nor UO_350 (O_350,N_4421,N_4438);
xor UO_351 (O_351,N_4264,N_4436);
or UO_352 (O_352,N_4607,N_4288);
or UO_353 (O_353,N_4959,N_4147);
or UO_354 (O_354,N_4205,N_4140);
and UO_355 (O_355,N_4270,N_4534);
nor UO_356 (O_356,N_4498,N_4888);
nand UO_357 (O_357,N_4553,N_4279);
xor UO_358 (O_358,N_4854,N_4973);
nand UO_359 (O_359,N_4856,N_4694);
and UO_360 (O_360,N_4706,N_4361);
nor UO_361 (O_361,N_4507,N_4399);
or UO_362 (O_362,N_4689,N_4744);
nand UO_363 (O_363,N_4256,N_4452);
and UO_364 (O_364,N_4167,N_4516);
or UO_365 (O_365,N_4822,N_4247);
xnor UO_366 (O_366,N_4010,N_4544);
and UO_367 (O_367,N_4506,N_4762);
and UO_368 (O_368,N_4118,N_4625);
nand UO_369 (O_369,N_4319,N_4629);
or UO_370 (O_370,N_4225,N_4852);
nor UO_371 (O_371,N_4913,N_4166);
nor UO_372 (O_372,N_4192,N_4395);
and UO_373 (O_373,N_4406,N_4165);
and UO_374 (O_374,N_4355,N_4678);
nand UO_375 (O_375,N_4161,N_4047);
and UO_376 (O_376,N_4457,N_4102);
or UO_377 (O_377,N_4887,N_4107);
nor UO_378 (O_378,N_4758,N_4381);
nor UO_379 (O_379,N_4904,N_4215);
or UO_380 (O_380,N_4435,N_4565);
or UO_381 (O_381,N_4704,N_4710);
or UO_382 (O_382,N_4527,N_4982);
nor UO_383 (O_383,N_4684,N_4763);
or UO_384 (O_384,N_4317,N_4283);
nor UO_385 (O_385,N_4074,N_4925);
or UO_386 (O_386,N_4410,N_4517);
or UO_387 (O_387,N_4814,N_4847);
or UO_388 (O_388,N_4871,N_4841);
nor UO_389 (O_389,N_4530,N_4572);
or UO_390 (O_390,N_4097,N_4362);
nand UO_391 (O_391,N_4100,N_4477);
and UO_392 (O_392,N_4339,N_4186);
nor UO_393 (O_393,N_4717,N_4323);
or UO_394 (O_394,N_4389,N_4431);
nor UO_395 (O_395,N_4716,N_4451);
nor UO_396 (O_396,N_4983,N_4485);
nand UO_397 (O_397,N_4386,N_4652);
xnor UO_398 (O_398,N_4193,N_4648);
and UO_399 (O_399,N_4079,N_4794);
nand UO_400 (O_400,N_4968,N_4447);
xnor UO_401 (O_401,N_4804,N_4575);
nand UO_402 (O_402,N_4433,N_4470);
or UO_403 (O_403,N_4387,N_4754);
and UO_404 (O_404,N_4646,N_4779);
nand UO_405 (O_405,N_4508,N_4138);
and UO_406 (O_406,N_4584,N_4310);
nor UO_407 (O_407,N_4184,N_4991);
or UO_408 (O_408,N_4408,N_4285);
or UO_409 (O_409,N_4474,N_4325);
or UO_410 (O_410,N_4793,N_4114);
or UO_411 (O_411,N_4201,N_4817);
and UO_412 (O_412,N_4352,N_4988);
nor UO_413 (O_413,N_4384,N_4187);
and UO_414 (O_414,N_4017,N_4239);
nand UO_415 (O_415,N_4200,N_4202);
or UO_416 (O_416,N_4977,N_4949);
and UO_417 (O_417,N_4786,N_4597);
nand UO_418 (O_418,N_4994,N_4230);
or UO_419 (O_419,N_4708,N_4700);
nand UO_420 (O_420,N_4737,N_4012);
and UO_421 (O_421,N_4876,N_4741);
or UO_422 (O_422,N_4391,N_4120);
nor UO_423 (O_423,N_4185,N_4169);
nand UO_424 (O_424,N_4974,N_4437);
and UO_425 (O_425,N_4868,N_4837);
and UO_426 (O_426,N_4825,N_4411);
or UO_427 (O_427,N_4023,N_4790);
and UO_428 (O_428,N_4154,N_4331);
or UO_429 (O_429,N_4970,N_4902);
nand UO_430 (O_430,N_4157,N_4479);
nor UO_431 (O_431,N_4043,N_4845);
nand UO_432 (O_432,N_4123,N_4698);
nand UO_433 (O_433,N_4836,N_4739);
or UO_434 (O_434,N_4388,N_4586);
or UO_435 (O_435,N_4755,N_4415);
nand UO_436 (O_436,N_4473,N_4927);
or UO_437 (O_437,N_4497,N_4986);
nand UO_438 (O_438,N_4318,N_4180);
and UO_439 (O_439,N_4103,N_4945);
nand UO_440 (O_440,N_4500,N_4259);
or UO_441 (O_441,N_4373,N_4233);
nor UO_442 (O_442,N_4197,N_4997);
or UO_443 (O_443,N_4260,N_4587);
and UO_444 (O_444,N_4518,N_4529);
nand UO_445 (O_445,N_4183,N_4392);
or UO_446 (O_446,N_4151,N_4174);
nor UO_447 (O_447,N_4641,N_4539);
or UO_448 (O_448,N_4075,N_4302);
nand UO_449 (O_449,N_4379,N_4609);
nand UO_450 (O_450,N_4413,N_4142);
and UO_451 (O_451,N_4746,N_4321);
and UO_452 (O_452,N_4307,N_4699);
and UO_453 (O_453,N_4329,N_4289);
or UO_454 (O_454,N_4265,N_4637);
nand UO_455 (O_455,N_4326,N_4301);
nor UO_456 (O_456,N_4409,N_4920);
nor UO_457 (O_457,N_4901,N_4962);
nor UO_458 (O_458,N_4995,N_4931);
and UO_459 (O_459,N_4676,N_4827);
nand UO_460 (O_460,N_4788,N_4941);
and UO_461 (O_461,N_4031,N_4828);
nor UO_462 (O_462,N_4089,N_4838);
nor UO_463 (O_463,N_4809,N_4182);
or UO_464 (O_464,N_4693,N_4701);
or UO_465 (O_465,N_4953,N_4475);
and UO_466 (O_466,N_4227,N_4611);
or UO_467 (O_467,N_4989,N_4802);
and UO_468 (O_468,N_4616,N_4649);
and UO_469 (O_469,N_4738,N_4213);
or UO_470 (O_470,N_4015,N_4914);
and UO_471 (O_471,N_4812,N_4462);
or UO_472 (O_472,N_4054,N_4049);
nand UO_473 (O_473,N_4309,N_4665);
or UO_474 (O_474,N_4732,N_4772);
or UO_475 (O_475,N_4803,N_4884);
or UO_476 (O_476,N_4088,N_4246);
or UO_477 (O_477,N_4673,N_4999);
nor UO_478 (O_478,N_4626,N_4162);
and UO_479 (O_479,N_4484,N_4025);
nor UO_480 (O_480,N_4449,N_4336);
nand UO_481 (O_481,N_4426,N_4843);
nor UO_482 (O_482,N_4826,N_4155);
nor UO_483 (O_483,N_4599,N_4940);
or UO_484 (O_484,N_4792,N_4095);
nor UO_485 (O_485,N_4469,N_4087);
nand UO_486 (O_486,N_4298,N_4558);
nand UO_487 (O_487,N_4011,N_4615);
nor UO_488 (O_488,N_4367,N_4489);
nand UO_489 (O_489,N_4685,N_4340);
nor UO_490 (O_490,N_4681,N_4723);
xor UO_491 (O_491,N_4650,N_4359);
or UO_492 (O_492,N_4492,N_4190);
and UO_493 (O_493,N_4606,N_4975);
and UO_494 (O_494,N_4713,N_4730);
nor UO_495 (O_495,N_4494,N_4004);
nor UO_496 (O_496,N_4209,N_4069);
and UO_497 (O_497,N_4337,N_4228);
xor UO_498 (O_498,N_4669,N_4294);
and UO_499 (O_499,N_4083,N_4085);
nand UO_500 (O_500,N_4907,N_4201);
or UO_501 (O_501,N_4664,N_4009);
nand UO_502 (O_502,N_4299,N_4361);
or UO_503 (O_503,N_4891,N_4542);
and UO_504 (O_504,N_4147,N_4195);
nand UO_505 (O_505,N_4308,N_4562);
nor UO_506 (O_506,N_4107,N_4350);
nor UO_507 (O_507,N_4904,N_4303);
and UO_508 (O_508,N_4402,N_4345);
and UO_509 (O_509,N_4909,N_4745);
nor UO_510 (O_510,N_4829,N_4496);
nand UO_511 (O_511,N_4297,N_4287);
nand UO_512 (O_512,N_4723,N_4576);
or UO_513 (O_513,N_4585,N_4164);
nor UO_514 (O_514,N_4428,N_4978);
and UO_515 (O_515,N_4278,N_4348);
nand UO_516 (O_516,N_4080,N_4220);
and UO_517 (O_517,N_4656,N_4284);
nor UO_518 (O_518,N_4464,N_4303);
and UO_519 (O_519,N_4468,N_4250);
nand UO_520 (O_520,N_4706,N_4809);
nor UO_521 (O_521,N_4068,N_4856);
or UO_522 (O_522,N_4254,N_4321);
nand UO_523 (O_523,N_4080,N_4669);
and UO_524 (O_524,N_4147,N_4013);
xnor UO_525 (O_525,N_4238,N_4487);
or UO_526 (O_526,N_4059,N_4766);
and UO_527 (O_527,N_4148,N_4428);
nand UO_528 (O_528,N_4668,N_4873);
nor UO_529 (O_529,N_4491,N_4588);
nor UO_530 (O_530,N_4288,N_4046);
nand UO_531 (O_531,N_4310,N_4518);
and UO_532 (O_532,N_4278,N_4591);
xor UO_533 (O_533,N_4288,N_4532);
or UO_534 (O_534,N_4681,N_4166);
and UO_535 (O_535,N_4643,N_4062);
and UO_536 (O_536,N_4211,N_4437);
nand UO_537 (O_537,N_4042,N_4765);
and UO_538 (O_538,N_4887,N_4830);
nor UO_539 (O_539,N_4735,N_4026);
and UO_540 (O_540,N_4573,N_4822);
or UO_541 (O_541,N_4038,N_4873);
nand UO_542 (O_542,N_4560,N_4229);
or UO_543 (O_543,N_4879,N_4660);
or UO_544 (O_544,N_4956,N_4814);
nand UO_545 (O_545,N_4330,N_4604);
nor UO_546 (O_546,N_4740,N_4581);
or UO_547 (O_547,N_4761,N_4918);
or UO_548 (O_548,N_4760,N_4452);
nor UO_549 (O_549,N_4039,N_4680);
nand UO_550 (O_550,N_4051,N_4017);
or UO_551 (O_551,N_4457,N_4257);
nand UO_552 (O_552,N_4122,N_4909);
nor UO_553 (O_553,N_4811,N_4581);
nor UO_554 (O_554,N_4764,N_4829);
nor UO_555 (O_555,N_4987,N_4511);
nor UO_556 (O_556,N_4321,N_4022);
and UO_557 (O_557,N_4786,N_4691);
or UO_558 (O_558,N_4138,N_4236);
and UO_559 (O_559,N_4800,N_4781);
or UO_560 (O_560,N_4387,N_4217);
and UO_561 (O_561,N_4808,N_4012);
xor UO_562 (O_562,N_4973,N_4804);
nand UO_563 (O_563,N_4772,N_4636);
nand UO_564 (O_564,N_4946,N_4680);
or UO_565 (O_565,N_4505,N_4552);
nor UO_566 (O_566,N_4401,N_4730);
nor UO_567 (O_567,N_4807,N_4816);
and UO_568 (O_568,N_4419,N_4831);
and UO_569 (O_569,N_4870,N_4401);
and UO_570 (O_570,N_4848,N_4763);
nor UO_571 (O_571,N_4726,N_4474);
and UO_572 (O_572,N_4542,N_4049);
nor UO_573 (O_573,N_4136,N_4003);
and UO_574 (O_574,N_4678,N_4549);
and UO_575 (O_575,N_4110,N_4465);
and UO_576 (O_576,N_4173,N_4680);
nand UO_577 (O_577,N_4406,N_4259);
nor UO_578 (O_578,N_4391,N_4896);
or UO_579 (O_579,N_4988,N_4738);
nand UO_580 (O_580,N_4091,N_4709);
nor UO_581 (O_581,N_4553,N_4863);
and UO_582 (O_582,N_4347,N_4274);
nor UO_583 (O_583,N_4437,N_4629);
and UO_584 (O_584,N_4475,N_4423);
nand UO_585 (O_585,N_4561,N_4902);
nor UO_586 (O_586,N_4351,N_4123);
nor UO_587 (O_587,N_4298,N_4676);
nor UO_588 (O_588,N_4700,N_4612);
and UO_589 (O_589,N_4442,N_4674);
nor UO_590 (O_590,N_4071,N_4055);
or UO_591 (O_591,N_4266,N_4087);
and UO_592 (O_592,N_4414,N_4445);
nor UO_593 (O_593,N_4203,N_4882);
nand UO_594 (O_594,N_4181,N_4047);
and UO_595 (O_595,N_4537,N_4758);
or UO_596 (O_596,N_4747,N_4912);
nand UO_597 (O_597,N_4037,N_4345);
or UO_598 (O_598,N_4750,N_4021);
and UO_599 (O_599,N_4985,N_4279);
nand UO_600 (O_600,N_4050,N_4759);
or UO_601 (O_601,N_4970,N_4587);
nor UO_602 (O_602,N_4218,N_4739);
and UO_603 (O_603,N_4735,N_4442);
nand UO_604 (O_604,N_4430,N_4578);
nand UO_605 (O_605,N_4480,N_4334);
nand UO_606 (O_606,N_4667,N_4664);
nor UO_607 (O_607,N_4032,N_4803);
nor UO_608 (O_608,N_4034,N_4584);
or UO_609 (O_609,N_4148,N_4262);
and UO_610 (O_610,N_4142,N_4050);
and UO_611 (O_611,N_4200,N_4438);
nand UO_612 (O_612,N_4608,N_4826);
or UO_613 (O_613,N_4947,N_4014);
and UO_614 (O_614,N_4961,N_4603);
or UO_615 (O_615,N_4997,N_4634);
nand UO_616 (O_616,N_4345,N_4862);
or UO_617 (O_617,N_4472,N_4270);
nor UO_618 (O_618,N_4930,N_4892);
nor UO_619 (O_619,N_4716,N_4978);
nor UO_620 (O_620,N_4359,N_4467);
and UO_621 (O_621,N_4777,N_4789);
nor UO_622 (O_622,N_4723,N_4535);
and UO_623 (O_623,N_4001,N_4499);
nor UO_624 (O_624,N_4463,N_4422);
nor UO_625 (O_625,N_4728,N_4328);
nor UO_626 (O_626,N_4901,N_4206);
nand UO_627 (O_627,N_4946,N_4106);
or UO_628 (O_628,N_4067,N_4976);
xnor UO_629 (O_629,N_4754,N_4163);
nor UO_630 (O_630,N_4865,N_4585);
or UO_631 (O_631,N_4716,N_4665);
xor UO_632 (O_632,N_4723,N_4229);
nor UO_633 (O_633,N_4287,N_4096);
nand UO_634 (O_634,N_4450,N_4700);
and UO_635 (O_635,N_4757,N_4073);
or UO_636 (O_636,N_4106,N_4333);
nand UO_637 (O_637,N_4312,N_4808);
nor UO_638 (O_638,N_4132,N_4960);
or UO_639 (O_639,N_4948,N_4287);
or UO_640 (O_640,N_4715,N_4074);
nand UO_641 (O_641,N_4022,N_4324);
and UO_642 (O_642,N_4884,N_4500);
nand UO_643 (O_643,N_4228,N_4993);
and UO_644 (O_644,N_4955,N_4087);
or UO_645 (O_645,N_4382,N_4202);
or UO_646 (O_646,N_4988,N_4954);
nor UO_647 (O_647,N_4339,N_4357);
and UO_648 (O_648,N_4514,N_4671);
and UO_649 (O_649,N_4931,N_4089);
nor UO_650 (O_650,N_4928,N_4877);
and UO_651 (O_651,N_4069,N_4968);
nor UO_652 (O_652,N_4920,N_4786);
nor UO_653 (O_653,N_4472,N_4887);
or UO_654 (O_654,N_4731,N_4234);
or UO_655 (O_655,N_4459,N_4824);
or UO_656 (O_656,N_4827,N_4595);
nand UO_657 (O_657,N_4843,N_4723);
or UO_658 (O_658,N_4731,N_4956);
nor UO_659 (O_659,N_4373,N_4985);
and UO_660 (O_660,N_4965,N_4117);
nand UO_661 (O_661,N_4254,N_4021);
or UO_662 (O_662,N_4122,N_4386);
nor UO_663 (O_663,N_4023,N_4676);
and UO_664 (O_664,N_4366,N_4238);
nand UO_665 (O_665,N_4319,N_4385);
and UO_666 (O_666,N_4218,N_4664);
nand UO_667 (O_667,N_4908,N_4639);
and UO_668 (O_668,N_4627,N_4207);
nand UO_669 (O_669,N_4957,N_4087);
nor UO_670 (O_670,N_4783,N_4415);
nor UO_671 (O_671,N_4919,N_4195);
nand UO_672 (O_672,N_4737,N_4408);
nor UO_673 (O_673,N_4205,N_4720);
nand UO_674 (O_674,N_4289,N_4310);
and UO_675 (O_675,N_4021,N_4834);
nand UO_676 (O_676,N_4282,N_4449);
and UO_677 (O_677,N_4145,N_4120);
nor UO_678 (O_678,N_4063,N_4432);
and UO_679 (O_679,N_4731,N_4383);
nand UO_680 (O_680,N_4082,N_4145);
or UO_681 (O_681,N_4819,N_4262);
and UO_682 (O_682,N_4272,N_4144);
nor UO_683 (O_683,N_4269,N_4615);
xnor UO_684 (O_684,N_4069,N_4887);
nand UO_685 (O_685,N_4670,N_4984);
nor UO_686 (O_686,N_4523,N_4959);
nand UO_687 (O_687,N_4597,N_4314);
nand UO_688 (O_688,N_4068,N_4227);
nand UO_689 (O_689,N_4518,N_4952);
and UO_690 (O_690,N_4274,N_4226);
and UO_691 (O_691,N_4535,N_4948);
and UO_692 (O_692,N_4595,N_4027);
or UO_693 (O_693,N_4881,N_4500);
and UO_694 (O_694,N_4124,N_4092);
or UO_695 (O_695,N_4253,N_4464);
nor UO_696 (O_696,N_4893,N_4992);
nand UO_697 (O_697,N_4723,N_4503);
nand UO_698 (O_698,N_4665,N_4815);
nand UO_699 (O_699,N_4999,N_4562);
and UO_700 (O_700,N_4268,N_4827);
and UO_701 (O_701,N_4108,N_4297);
or UO_702 (O_702,N_4402,N_4881);
nand UO_703 (O_703,N_4758,N_4363);
or UO_704 (O_704,N_4344,N_4070);
or UO_705 (O_705,N_4012,N_4133);
nand UO_706 (O_706,N_4895,N_4750);
nor UO_707 (O_707,N_4403,N_4107);
nor UO_708 (O_708,N_4131,N_4283);
and UO_709 (O_709,N_4958,N_4687);
and UO_710 (O_710,N_4361,N_4659);
nand UO_711 (O_711,N_4787,N_4638);
nand UO_712 (O_712,N_4323,N_4265);
xnor UO_713 (O_713,N_4685,N_4529);
nor UO_714 (O_714,N_4561,N_4398);
nand UO_715 (O_715,N_4679,N_4254);
nand UO_716 (O_716,N_4798,N_4976);
or UO_717 (O_717,N_4691,N_4983);
nand UO_718 (O_718,N_4158,N_4722);
or UO_719 (O_719,N_4022,N_4637);
or UO_720 (O_720,N_4871,N_4040);
and UO_721 (O_721,N_4338,N_4099);
nand UO_722 (O_722,N_4638,N_4232);
and UO_723 (O_723,N_4515,N_4320);
nand UO_724 (O_724,N_4175,N_4326);
nand UO_725 (O_725,N_4871,N_4973);
nand UO_726 (O_726,N_4413,N_4062);
nand UO_727 (O_727,N_4911,N_4783);
or UO_728 (O_728,N_4386,N_4811);
nand UO_729 (O_729,N_4561,N_4989);
or UO_730 (O_730,N_4211,N_4488);
nand UO_731 (O_731,N_4303,N_4654);
nand UO_732 (O_732,N_4955,N_4460);
nand UO_733 (O_733,N_4854,N_4425);
nor UO_734 (O_734,N_4937,N_4965);
nand UO_735 (O_735,N_4449,N_4173);
nor UO_736 (O_736,N_4305,N_4932);
nand UO_737 (O_737,N_4299,N_4374);
and UO_738 (O_738,N_4152,N_4678);
nor UO_739 (O_739,N_4278,N_4879);
and UO_740 (O_740,N_4413,N_4398);
or UO_741 (O_741,N_4213,N_4882);
or UO_742 (O_742,N_4760,N_4704);
nor UO_743 (O_743,N_4134,N_4869);
and UO_744 (O_744,N_4739,N_4095);
and UO_745 (O_745,N_4396,N_4016);
nand UO_746 (O_746,N_4656,N_4208);
nand UO_747 (O_747,N_4990,N_4004);
nand UO_748 (O_748,N_4504,N_4115);
nand UO_749 (O_749,N_4609,N_4184);
nor UO_750 (O_750,N_4168,N_4539);
nand UO_751 (O_751,N_4243,N_4424);
or UO_752 (O_752,N_4005,N_4500);
and UO_753 (O_753,N_4142,N_4279);
nand UO_754 (O_754,N_4951,N_4403);
nor UO_755 (O_755,N_4608,N_4796);
and UO_756 (O_756,N_4833,N_4771);
nand UO_757 (O_757,N_4893,N_4539);
nand UO_758 (O_758,N_4977,N_4342);
nand UO_759 (O_759,N_4626,N_4018);
and UO_760 (O_760,N_4152,N_4358);
or UO_761 (O_761,N_4866,N_4338);
or UO_762 (O_762,N_4780,N_4002);
nor UO_763 (O_763,N_4118,N_4010);
nor UO_764 (O_764,N_4126,N_4110);
or UO_765 (O_765,N_4505,N_4036);
or UO_766 (O_766,N_4776,N_4984);
or UO_767 (O_767,N_4306,N_4118);
nand UO_768 (O_768,N_4597,N_4785);
nor UO_769 (O_769,N_4589,N_4186);
or UO_770 (O_770,N_4425,N_4259);
or UO_771 (O_771,N_4915,N_4064);
and UO_772 (O_772,N_4391,N_4959);
or UO_773 (O_773,N_4765,N_4328);
nor UO_774 (O_774,N_4680,N_4827);
nor UO_775 (O_775,N_4105,N_4843);
nor UO_776 (O_776,N_4604,N_4612);
and UO_777 (O_777,N_4597,N_4682);
nor UO_778 (O_778,N_4607,N_4672);
xor UO_779 (O_779,N_4974,N_4065);
or UO_780 (O_780,N_4245,N_4031);
nor UO_781 (O_781,N_4251,N_4161);
xnor UO_782 (O_782,N_4854,N_4411);
or UO_783 (O_783,N_4636,N_4103);
and UO_784 (O_784,N_4173,N_4987);
nor UO_785 (O_785,N_4591,N_4063);
or UO_786 (O_786,N_4203,N_4854);
and UO_787 (O_787,N_4767,N_4235);
nand UO_788 (O_788,N_4077,N_4196);
nor UO_789 (O_789,N_4172,N_4486);
nand UO_790 (O_790,N_4831,N_4213);
and UO_791 (O_791,N_4908,N_4286);
nor UO_792 (O_792,N_4590,N_4355);
nor UO_793 (O_793,N_4564,N_4544);
nor UO_794 (O_794,N_4302,N_4568);
or UO_795 (O_795,N_4536,N_4585);
and UO_796 (O_796,N_4015,N_4824);
nor UO_797 (O_797,N_4463,N_4840);
and UO_798 (O_798,N_4040,N_4862);
nor UO_799 (O_799,N_4327,N_4709);
nand UO_800 (O_800,N_4172,N_4313);
or UO_801 (O_801,N_4380,N_4955);
or UO_802 (O_802,N_4804,N_4023);
or UO_803 (O_803,N_4244,N_4784);
or UO_804 (O_804,N_4094,N_4132);
and UO_805 (O_805,N_4623,N_4569);
nor UO_806 (O_806,N_4721,N_4364);
nor UO_807 (O_807,N_4028,N_4208);
nand UO_808 (O_808,N_4938,N_4578);
and UO_809 (O_809,N_4411,N_4253);
and UO_810 (O_810,N_4998,N_4333);
nor UO_811 (O_811,N_4060,N_4132);
nor UO_812 (O_812,N_4583,N_4428);
nor UO_813 (O_813,N_4964,N_4322);
nor UO_814 (O_814,N_4462,N_4737);
or UO_815 (O_815,N_4847,N_4576);
nand UO_816 (O_816,N_4718,N_4037);
xnor UO_817 (O_817,N_4931,N_4346);
and UO_818 (O_818,N_4557,N_4992);
and UO_819 (O_819,N_4705,N_4488);
nor UO_820 (O_820,N_4721,N_4654);
or UO_821 (O_821,N_4520,N_4727);
nor UO_822 (O_822,N_4864,N_4929);
nor UO_823 (O_823,N_4784,N_4298);
and UO_824 (O_824,N_4902,N_4213);
nand UO_825 (O_825,N_4826,N_4974);
nand UO_826 (O_826,N_4333,N_4929);
nor UO_827 (O_827,N_4375,N_4855);
or UO_828 (O_828,N_4136,N_4995);
or UO_829 (O_829,N_4491,N_4141);
nor UO_830 (O_830,N_4198,N_4420);
nor UO_831 (O_831,N_4596,N_4372);
or UO_832 (O_832,N_4114,N_4779);
nand UO_833 (O_833,N_4672,N_4315);
and UO_834 (O_834,N_4922,N_4645);
and UO_835 (O_835,N_4936,N_4045);
nor UO_836 (O_836,N_4469,N_4474);
nor UO_837 (O_837,N_4180,N_4423);
nand UO_838 (O_838,N_4851,N_4902);
nor UO_839 (O_839,N_4802,N_4366);
or UO_840 (O_840,N_4138,N_4421);
nor UO_841 (O_841,N_4414,N_4762);
nor UO_842 (O_842,N_4347,N_4791);
nand UO_843 (O_843,N_4862,N_4161);
nor UO_844 (O_844,N_4956,N_4602);
and UO_845 (O_845,N_4156,N_4061);
or UO_846 (O_846,N_4816,N_4812);
or UO_847 (O_847,N_4915,N_4745);
or UO_848 (O_848,N_4628,N_4175);
or UO_849 (O_849,N_4303,N_4051);
or UO_850 (O_850,N_4771,N_4008);
and UO_851 (O_851,N_4638,N_4047);
and UO_852 (O_852,N_4974,N_4393);
and UO_853 (O_853,N_4959,N_4209);
nand UO_854 (O_854,N_4445,N_4748);
or UO_855 (O_855,N_4447,N_4406);
nor UO_856 (O_856,N_4036,N_4411);
nand UO_857 (O_857,N_4905,N_4113);
nor UO_858 (O_858,N_4391,N_4392);
nand UO_859 (O_859,N_4828,N_4265);
nor UO_860 (O_860,N_4071,N_4809);
or UO_861 (O_861,N_4231,N_4882);
xor UO_862 (O_862,N_4243,N_4756);
and UO_863 (O_863,N_4085,N_4240);
and UO_864 (O_864,N_4023,N_4743);
nand UO_865 (O_865,N_4407,N_4839);
nand UO_866 (O_866,N_4407,N_4380);
and UO_867 (O_867,N_4365,N_4660);
nor UO_868 (O_868,N_4185,N_4563);
nand UO_869 (O_869,N_4010,N_4040);
or UO_870 (O_870,N_4499,N_4969);
or UO_871 (O_871,N_4636,N_4165);
nand UO_872 (O_872,N_4465,N_4150);
nor UO_873 (O_873,N_4583,N_4912);
and UO_874 (O_874,N_4349,N_4397);
or UO_875 (O_875,N_4793,N_4578);
and UO_876 (O_876,N_4815,N_4779);
nor UO_877 (O_877,N_4097,N_4866);
or UO_878 (O_878,N_4222,N_4987);
nand UO_879 (O_879,N_4867,N_4925);
nand UO_880 (O_880,N_4953,N_4489);
nor UO_881 (O_881,N_4067,N_4740);
or UO_882 (O_882,N_4308,N_4921);
and UO_883 (O_883,N_4977,N_4401);
nand UO_884 (O_884,N_4094,N_4093);
xnor UO_885 (O_885,N_4647,N_4561);
or UO_886 (O_886,N_4361,N_4967);
nand UO_887 (O_887,N_4226,N_4206);
and UO_888 (O_888,N_4840,N_4959);
or UO_889 (O_889,N_4170,N_4911);
nand UO_890 (O_890,N_4538,N_4024);
nand UO_891 (O_891,N_4104,N_4808);
and UO_892 (O_892,N_4413,N_4912);
nor UO_893 (O_893,N_4550,N_4969);
nor UO_894 (O_894,N_4217,N_4094);
nor UO_895 (O_895,N_4464,N_4166);
nand UO_896 (O_896,N_4824,N_4162);
nand UO_897 (O_897,N_4481,N_4393);
nand UO_898 (O_898,N_4646,N_4257);
or UO_899 (O_899,N_4113,N_4618);
nand UO_900 (O_900,N_4254,N_4358);
nand UO_901 (O_901,N_4643,N_4654);
and UO_902 (O_902,N_4448,N_4441);
and UO_903 (O_903,N_4085,N_4441);
nand UO_904 (O_904,N_4361,N_4985);
nand UO_905 (O_905,N_4787,N_4942);
and UO_906 (O_906,N_4762,N_4299);
and UO_907 (O_907,N_4603,N_4760);
nand UO_908 (O_908,N_4424,N_4772);
nand UO_909 (O_909,N_4102,N_4776);
and UO_910 (O_910,N_4996,N_4257);
nand UO_911 (O_911,N_4545,N_4598);
nand UO_912 (O_912,N_4652,N_4625);
xnor UO_913 (O_913,N_4378,N_4495);
or UO_914 (O_914,N_4325,N_4871);
and UO_915 (O_915,N_4819,N_4399);
or UO_916 (O_916,N_4158,N_4485);
nand UO_917 (O_917,N_4834,N_4496);
and UO_918 (O_918,N_4929,N_4837);
or UO_919 (O_919,N_4562,N_4020);
or UO_920 (O_920,N_4684,N_4601);
nand UO_921 (O_921,N_4897,N_4128);
nor UO_922 (O_922,N_4573,N_4253);
nor UO_923 (O_923,N_4950,N_4926);
nor UO_924 (O_924,N_4452,N_4521);
nor UO_925 (O_925,N_4694,N_4166);
nor UO_926 (O_926,N_4094,N_4633);
nand UO_927 (O_927,N_4054,N_4913);
nand UO_928 (O_928,N_4202,N_4587);
nand UO_929 (O_929,N_4219,N_4839);
nor UO_930 (O_930,N_4983,N_4475);
nand UO_931 (O_931,N_4828,N_4621);
nand UO_932 (O_932,N_4671,N_4825);
and UO_933 (O_933,N_4839,N_4273);
and UO_934 (O_934,N_4317,N_4004);
nor UO_935 (O_935,N_4254,N_4572);
nand UO_936 (O_936,N_4537,N_4381);
nand UO_937 (O_937,N_4716,N_4293);
or UO_938 (O_938,N_4306,N_4178);
or UO_939 (O_939,N_4994,N_4941);
nor UO_940 (O_940,N_4023,N_4587);
and UO_941 (O_941,N_4088,N_4593);
or UO_942 (O_942,N_4634,N_4432);
nand UO_943 (O_943,N_4778,N_4304);
or UO_944 (O_944,N_4468,N_4802);
or UO_945 (O_945,N_4705,N_4293);
or UO_946 (O_946,N_4890,N_4864);
or UO_947 (O_947,N_4466,N_4861);
nand UO_948 (O_948,N_4406,N_4523);
and UO_949 (O_949,N_4016,N_4932);
or UO_950 (O_950,N_4965,N_4623);
and UO_951 (O_951,N_4800,N_4581);
nor UO_952 (O_952,N_4169,N_4282);
or UO_953 (O_953,N_4013,N_4164);
nand UO_954 (O_954,N_4964,N_4179);
nand UO_955 (O_955,N_4411,N_4237);
or UO_956 (O_956,N_4917,N_4813);
or UO_957 (O_957,N_4651,N_4401);
and UO_958 (O_958,N_4208,N_4716);
and UO_959 (O_959,N_4822,N_4665);
or UO_960 (O_960,N_4837,N_4478);
and UO_961 (O_961,N_4572,N_4742);
nor UO_962 (O_962,N_4340,N_4328);
nand UO_963 (O_963,N_4832,N_4059);
or UO_964 (O_964,N_4194,N_4985);
and UO_965 (O_965,N_4980,N_4255);
nor UO_966 (O_966,N_4402,N_4511);
or UO_967 (O_967,N_4860,N_4104);
nor UO_968 (O_968,N_4098,N_4642);
or UO_969 (O_969,N_4967,N_4652);
or UO_970 (O_970,N_4945,N_4109);
nor UO_971 (O_971,N_4000,N_4112);
or UO_972 (O_972,N_4348,N_4464);
nand UO_973 (O_973,N_4894,N_4625);
and UO_974 (O_974,N_4892,N_4498);
nand UO_975 (O_975,N_4254,N_4239);
nand UO_976 (O_976,N_4466,N_4923);
nand UO_977 (O_977,N_4765,N_4986);
or UO_978 (O_978,N_4755,N_4186);
nor UO_979 (O_979,N_4760,N_4566);
nor UO_980 (O_980,N_4762,N_4794);
or UO_981 (O_981,N_4299,N_4460);
nor UO_982 (O_982,N_4828,N_4941);
and UO_983 (O_983,N_4914,N_4377);
nand UO_984 (O_984,N_4577,N_4297);
nand UO_985 (O_985,N_4164,N_4206);
nand UO_986 (O_986,N_4276,N_4264);
nor UO_987 (O_987,N_4867,N_4074);
nor UO_988 (O_988,N_4590,N_4374);
nand UO_989 (O_989,N_4060,N_4369);
and UO_990 (O_990,N_4492,N_4632);
or UO_991 (O_991,N_4695,N_4803);
nor UO_992 (O_992,N_4680,N_4440);
nor UO_993 (O_993,N_4416,N_4558);
and UO_994 (O_994,N_4776,N_4513);
nand UO_995 (O_995,N_4029,N_4428);
and UO_996 (O_996,N_4020,N_4775);
or UO_997 (O_997,N_4197,N_4824);
or UO_998 (O_998,N_4637,N_4025);
nor UO_999 (O_999,N_4792,N_4816);
endmodule