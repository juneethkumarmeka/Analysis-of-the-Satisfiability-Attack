module basic_1000_10000_1500_20_levels_5xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
and U0 (N_0,In_969,In_200);
or U1 (N_1,In_361,In_173);
or U2 (N_2,In_378,In_911);
or U3 (N_3,In_269,In_219);
nor U4 (N_4,In_474,In_608);
or U5 (N_5,In_424,In_923);
and U6 (N_6,In_304,In_501);
nand U7 (N_7,In_3,In_636);
nand U8 (N_8,In_646,In_189);
or U9 (N_9,In_399,In_791);
nor U10 (N_10,In_752,In_210);
nand U11 (N_11,In_951,In_881);
or U12 (N_12,In_92,In_75);
and U13 (N_13,In_63,In_740);
or U14 (N_14,In_476,In_701);
nand U15 (N_15,In_493,In_97);
xnor U16 (N_16,In_855,In_820);
and U17 (N_17,In_345,In_296);
and U18 (N_18,In_594,In_109);
nor U19 (N_19,In_366,In_674);
xor U20 (N_20,In_813,In_984);
and U21 (N_21,In_913,In_599);
nand U22 (N_22,In_277,In_801);
or U23 (N_23,In_145,In_498);
nand U24 (N_24,In_255,In_153);
and U25 (N_25,In_922,In_696);
and U26 (N_26,In_241,In_449);
nand U27 (N_27,In_440,In_879);
or U28 (N_28,In_218,In_300);
nor U29 (N_29,In_460,In_726);
nor U30 (N_30,In_978,In_874);
nand U31 (N_31,In_258,In_687);
nand U32 (N_32,In_216,In_78);
nand U33 (N_33,In_810,In_187);
or U34 (N_34,In_166,In_179);
or U35 (N_35,In_254,In_172);
or U36 (N_36,In_120,In_30);
nand U37 (N_37,In_47,In_953);
nor U38 (N_38,In_665,In_682);
and U39 (N_39,In_483,In_621);
nand U40 (N_40,In_264,In_683);
and U41 (N_41,In_783,In_5);
and U42 (N_42,In_212,In_634);
nand U43 (N_43,In_662,In_418);
nand U44 (N_44,In_247,In_628);
nand U45 (N_45,In_561,In_133);
nor U46 (N_46,In_986,In_273);
nand U47 (N_47,In_523,In_387);
or U48 (N_48,In_585,In_68);
or U49 (N_49,In_147,In_142);
nand U50 (N_50,In_306,In_640);
and U51 (N_51,In_582,In_780);
xor U52 (N_52,In_240,In_528);
nand U53 (N_53,In_265,In_898);
and U54 (N_54,In_131,In_949);
nor U55 (N_55,In_948,In_360);
and U56 (N_56,In_473,In_482);
nor U57 (N_57,In_393,In_124);
nor U58 (N_58,In_759,In_128);
nor U59 (N_59,In_650,In_436);
or U60 (N_60,In_495,In_556);
nor U61 (N_61,In_91,In_417);
nor U62 (N_62,In_450,In_137);
nand U63 (N_63,In_257,In_467);
and U64 (N_64,In_283,In_485);
nor U65 (N_65,In_244,In_851);
or U66 (N_66,In_666,In_975);
nor U67 (N_67,In_544,In_633);
nand U68 (N_68,In_135,In_382);
or U69 (N_69,In_602,In_815);
nor U70 (N_70,In_617,In_769);
nand U71 (N_71,In_676,In_688);
and U72 (N_72,In_199,In_65);
nand U73 (N_73,In_644,In_822);
nor U74 (N_74,In_645,In_170);
or U75 (N_75,In_966,In_190);
and U76 (N_76,In_49,In_321);
nand U77 (N_77,In_282,In_13);
or U78 (N_78,In_936,In_336);
or U79 (N_79,In_253,In_99);
or U80 (N_80,In_712,In_389);
or U81 (N_81,In_568,In_339);
and U82 (N_82,In_130,In_7);
nand U83 (N_83,In_191,In_108);
nor U84 (N_84,In_977,In_895);
nor U85 (N_85,In_235,In_295);
nor U86 (N_86,In_20,In_880);
and U87 (N_87,In_243,In_517);
or U88 (N_88,In_165,In_454);
and U89 (N_89,In_394,In_654);
nor U90 (N_90,In_819,In_431);
nor U91 (N_91,In_846,In_349);
or U92 (N_92,In_765,In_148);
nor U93 (N_93,In_11,In_693);
and U94 (N_94,In_175,In_578);
and U95 (N_95,In_136,In_955);
nand U96 (N_96,In_756,In_45);
nor U97 (N_97,In_263,In_420);
and U98 (N_98,In_824,In_967);
nor U99 (N_99,In_694,In_525);
nor U100 (N_100,In_285,In_533);
or U101 (N_101,In_188,In_311);
and U102 (N_102,In_81,In_500);
nor U103 (N_103,In_419,In_248);
and U104 (N_104,In_267,In_299);
or U105 (N_105,In_384,In_62);
nor U106 (N_106,In_102,In_412);
nand U107 (N_107,In_660,In_875);
and U108 (N_108,In_841,In_176);
nand U109 (N_109,In_747,In_268);
nand U110 (N_110,In_853,In_798);
xor U111 (N_111,In_994,In_479);
nor U112 (N_112,In_509,In_208);
xnor U113 (N_113,In_987,In_775);
nor U114 (N_114,In_433,In_658);
nand U115 (N_115,In_404,In_900);
or U116 (N_116,In_941,In_596);
nand U117 (N_117,In_709,In_601);
nand U118 (N_118,In_335,In_564);
nand U119 (N_119,In_558,In_19);
nand U120 (N_120,In_0,In_885);
nand U121 (N_121,In_28,In_587);
xnor U122 (N_122,In_639,In_209);
and U123 (N_123,In_231,In_878);
nand U124 (N_124,In_860,In_100);
or U125 (N_125,In_274,In_475);
or U126 (N_126,In_921,In_678);
nor U127 (N_127,In_849,In_746);
xor U128 (N_128,In_591,In_757);
nand U129 (N_129,In_332,In_362);
xor U130 (N_130,In_615,In_252);
or U131 (N_131,In_43,In_391);
nand U132 (N_132,In_699,In_232);
nor U133 (N_133,In_272,In_991);
xor U134 (N_134,In_18,In_121);
nor U135 (N_135,In_831,In_426);
nand U136 (N_136,In_333,In_408);
nor U137 (N_137,In_446,In_88);
or U138 (N_138,In_799,In_227);
nor U139 (N_139,In_869,In_185);
nand U140 (N_140,In_320,In_623);
and U141 (N_141,In_286,In_718);
and U142 (N_142,In_432,In_888);
and U143 (N_143,In_551,In_992);
or U144 (N_144,In_341,In_547);
or U145 (N_145,In_23,In_787);
nand U146 (N_146,In_716,In_157);
nand U147 (N_147,In_85,In_89);
xor U148 (N_148,In_742,In_359);
nor U149 (N_149,In_723,In_939);
nand U150 (N_150,In_893,In_803);
and U151 (N_151,In_972,In_926);
nor U152 (N_152,In_53,In_552);
nor U153 (N_153,In_684,In_714);
or U154 (N_154,In_868,In_655);
nor U155 (N_155,In_260,In_220);
or U156 (N_156,In_537,In_996);
nand U157 (N_157,In_863,In_312);
nor U158 (N_158,In_764,In_445);
and U159 (N_159,In_94,In_961);
xor U160 (N_160,In_510,In_751);
or U161 (N_161,In_163,In_541);
xnor U162 (N_162,In_720,In_129);
xnor U163 (N_163,In_343,In_211);
xor U164 (N_164,In_183,In_298);
nand U165 (N_165,In_266,In_228);
nor U166 (N_166,In_581,In_867);
nor U167 (N_167,In_758,In_622);
nand U168 (N_168,In_203,In_937);
nor U169 (N_169,In_364,In_837);
nand U170 (N_170,In_207,In_838);
and U171 (N_171,In_318,In_125);
nand U172 (N_172,In_155,In_372);
and U173 (N_173,In_229,In_910);
nor U174 (N_174,In_308,In_821);
nand U175 (N_175,In_536,In_854);
or U176 (N_176,In_999,In_39);
or U177 (N_177,In_952,In_648);
xnor U178 (N_178,In_883,In_671);
or U179 (N_179,In_668,In_123);
nand U180 (N_180,In_721,In_584);
nor U181 (N_181,In_466,In_402);
and U182 (N_182,In_10,In_638);
and U183 (N_183,In_370,In_899);
nor U184 (N_184,In_83,In_386);
nor U185 (N_185,In_346,In_672);
nand U186 (N_186,In_256,In_985);
or U187 (N_187,In_470,In_856);
xnor U188 (N_188,In_105,In_70);
and U189 (N_189,In_670,In_988);
or U190 (N_190,In_158,In_713);
nand U191 (N_191,In_468,In_462);
or U192 (N_192,In_598,In_606);
or U193 (N_193,In_511,In_794);
and U194 (N_194,In_781,In_276);
or U195 (N_195,In_58,In_589);
or U196 (N_196,In_278,In_724);
nor U197 (N_197,In_873,In_326);
nand U198 (N_198,In_572,In_44);
xnor U199 (N_199,In_383,In_110);
or U200 (N_200,In_496,In_358);
or U201 (N_201,In_438,In_437);
xor U202 (N_202,In_945,In_61);
nand U203 (N_203,In_772,In_620);
or U204 (N_204,In_592,In_281);
nor U205 (N_205,In_486,In_681);
and U206 (N_206,In_652,In_882);
and U207 (N_207,In_48,In_98);
nor U208 (N_208,In_365,In_237);
and U209 (N_209,In_839,In_770);
nand U210 (N_210,In_653,In_962);
or U211 (N_211,In_421,In_569);
nor U212 (N_212,In_637,In_927);
or U213 (N_213,In_351,In_983);
nor U214 (N_214,In_330,In_609);
nor U215 (N_215,In_194,In_149);
nand U216 (N_216,In_524,In_643);
nand U217 (N_217,In_503,In_982);
nand U218 (N_218,In_980,In_892);
and U219 (N_219,In_776,In_215);
nand U220 (N_220,In_886,In_8);
or U221 (N_221,In_738,In_377);
or U222 (N_222,In_347,In_401);
nor U223 (N_223,In_754,In_21);
and U224 (N_224,In_12,In_192);
nand U225 (N_225,In_379,In_403);
or U226 (N_226,In_795,In_659);
or U227 (N_227,In_167,In_549);
and U228 (N_228,In_958,In_139);
nor U229 (N_229,In_57,In_559);
and U230 (N_230,In_107,In_706);
or U231 (N_231,In_641,In_857);
nor U232 (N_232,In_827,In_14);
and U233 (N_233,In_24,In_571);
nor U234 (N_234,In_531,In_150);
or U235 (N_235,In_118,In_848);
or U236 (N_236,In_270,In_891);
and U237 (N_237,In_380,In_538);
or U238 (N_238,In_146,In_381);
nor U239 (N_239,In_447,In_518);
or U240 (N_240,In_164,In_297);
nor U241 (N_241,In_522,In_334);
nand U242 (N_242,In_680,In_465);
nand U243 (N_243,In_292,In_793);
nand U244 (N_244,In_675,In_287);
or U245 (N_245,In_938,In_542);
xnor U246 (N_246,In_603,In_736);
and U247 (N_247,In_202,In_489);
nor U248 (N_248,In_656,In_710);
nor U249 (N_249,In_317,In_931);
nand U250 (N_250,In_233,In_245);
nand U251 (N_251,In_797,In_575);
or U252 (N_252,In_168,In_979);
nand U253 (N_253,In_872,In_457);
nor U254 (N_254,In_916,In_612);
and U255 (N_255,In_814,In_520);
and U256 (N_256,In_217,In_302);
and U257 (N_257,In_152,In_904);
or U258 (N_258,In_181,In_570);
nor U259 (N_259,In_458,In_186);
nor U260 (N_260,In_852,In_647);
or U261 (N_261,In_305,In_588);
and U262 (N_262,In_37,In_293);
and U263 (N_263,In_902,In_735);
nand U264 (N_264,In_722,In_204);
nor U265 (N_265,In_777,In_817);
xnor U266 (N_266,In_2,In_845);
and U267 (N_267,In_95,In_562);
or U268 (N_268,In_909,In_36);
nor U269 (N_269,In_77,In_87);
xnor U270 (N_270,In_64,In_411);
or U271 (N_271,In_41,In_823);
and U272 (N_272,In_935,In_870);
and U273 (N_273,In_516,In_160);
nand U274 (N_274,In_995,In_230);
or U275 (N_275,In_322,In_356);
and U276 (N_276,In_560,In_613);
nor U277 (N_277,In_513,In_239);
nor U278 (N_278,In_444,In_546);
and U279 (N_279,In_527,In_428);
nand U280 (N_280,In_597,In_861);
xor U281 (N_281,In_469,In_405);
xnor U282 (N_282,In_353,In_989);
and U283 (N_283,In_491,In_112);
nand U284 (N_284,In_236,In_455);
nor U285 (N_285,In_786,In_830);
or U286 (N_286,In_117,In_246);
xor U287 (N_287,In_906,In_126);
or U288 (N_288,In_315,In_692);
nor U289 (N_289,In_410,In_79);
xor U290 (N_290,In_630,In_748);
or U291 (N_291,In_607,In_708);
nand U292 (N_292,In_313,In_555);
and U293 (N_293,In_80,In_414);
or U294 (N_294,In_106,In_141);
nand U295 (N_295,In_526,In_506);
or U296 (N_296,In_456,In_583);
nand U297 (N_297,In_423,In_779);
and U298 (N_298,In_279,In_642);
and U299 (N_299,In_836,In_981);
or U300 (N_300,In_512,In_725);
and U301 (N_301,In_38,In_625);
nor U302 (N_302,In_529,In_327);
nand U303 (N_303,In_771,In_565);
nand U304 (N_304,In_956,In_734);
or U305 (N_305,In_632,In_811);
or U306 (N_306,In_543,In_805);
nor U307 (N_307,In_943,In_416);
nand U308 (N_308,In_908,In_354);
and U309 (N_309,In_844,In_34);
nor U310 (N_310,In_877,In_840);
and U311 (N_311,In_90,In_717);
xnor U312 (N_312,In_371,In_395);
nor U313 (N_313,In_990,In_871);
xor U314 (N_314,In_553,In_993);
and U315 (N_315,In_829,In_251);
or U316 (N_316,In_507,In_971);
and U317 (N_317,In_413,In_842);
xor U318 (N_318,In_422,In_288);
nand U319 (N_319,In_342,In_887);
nand U320 (N_320,In_812,In_225);
nor U321 (N_321,In_930,In_226);
or U322 (N_322,In_119,In_114);
and U323 (N_323,In_17,In_439);
nand U324 (N_324,In_732,In_605);
xnor U325 (N_325,In_69,In_750);
xnor U326 (N_326,In_729,In_785);
xnor U327 (N_327,In_790,In_250);
nor U328 (N_328,In_586,In_657);
or U329 (N_329,In_73,In_959);
nand U330 (N_330,In_914,In_976);
xnor U331 (N_331,In_700,In_213);
or U332 (N_332,In_784,In_957);
and U333 (N_333,In_649,In_540);
or U334 (N_334,In_398,In_545);
nor U335 (N_335,In_463,In_71);
nand U336 (N_336,In_532,In_651);
xnor U337 (N_337,In_397,In_374);
nor U338 (N_338,In_331,In_903);
nor U339 (N_339,In_610,In_530);
or U340 (N_340,In_698,In_385);
nand U341 (N_341,In_242,In_800);
xnor U342 (N_342,In_850,In_448);
or U343 (N_343,In_376,In_284);
nor U344 (N_344,In_72,In_677);
nor U345 (N_345,In_143,In_162);
xnor U346 (N_346,In_280,In_50);
or U347 (N_347,In_942,In_429);
or U348 (N_348,In_487,In_974);
and U349 (N_349,In_328,In_884);
and U350 (N_350,In_375,In_177);
xor U351 (N_351,In_940,In_773);
and U352 (N_352,In_593,In_6);
nor U353 (N_353,In_324,In_929);
and U354 (N_354,In_234,In_329);
nor U355 (N_355,In_392,In_352);
nand U356 (N_356,In_464,In_806);
nor U357 (N_357,In_290,In_944);
or U358 (N_358,In_196,In_25);
nor U359 (N_359,In_481,In_103);
or U360 (N_360,In_737,In_629);
and U361 (N_361,In_604,In_138);
nand U362 (N_362,In_753,In_802);
and U363 (N_363,In_847,In_340);
or U364 (N_364,In_499,In_865);
and U365 (N_365,In_521,In_685);
xor U366 (N_366,In_539,In_744);
nand U367 (N_367,In_453,In_368);
or U368 (N_368,In_127,In_901);
or U369 (N_369,In_719,In_249);
or U370 (N_370,In_833,In_259);
and U371 (N_371,In_894,In_862);
and U372 (N_372,In_1,In_74);
nand U373 (N_373,In_932,In_184);
nor U374 (N_374,In_82,In_434);
nand U375 (N_375,In_223,In_919);
nand U376 (N_376,In_858,In_174);
nor U377 (N_377,In_702,In_310);
nand U378 (N_378,In_101,In_579);
nand U379 (N_379,In_508,In_828);
nor U380 (N_380,In_774,In_93);
nor U381 (N_381,In_915,In_704);
nor U382 (N_382,In_425,In_182);
and U383 (N_383,In_221,In_535);
or U384 (N_384,In_195,In_925);
nand U385 (N_385,In_859,In_618);
or U386 (N_386,In_261,In_614);
nand U387 (N_387,In_111,In_789);
nand U388 (N_388,In_494,In_369);
xor U389 (N_389,In_122,In_954);
nor U390 (N_390,In_407,In_224);
or U391 (N_391,In_33,In_695);
nor U392 (N_392,In_619,In_350);
and U393 (N_393,In_924,In_554);
and U394 (N_394,In_627,In_154);
or U395 (N_395,In_534,In_205);
or U396 (N_396,In_960,In_970);
and U397 (N_397,In_178,In_161);
and U398 (N_398,In_262,In_950);
and U399 (N_399,In_400,In_762);
and U400 (N_400,In_749,In_663);
nor U401 (N_401,In_825,In_782);
or U402 (N_402,In_727,In_180);
and U403 (N_403,In_140,In_104);
nor U404 (N_404,In_733,In_889);
xnor U405 (N_405,In_519,In_731);
or U406 (N_406,In_67,In_406);
nor U407 (N_407,In_920,In_743);
and U408 (N_408,In_275,In_624);
or U409 (N_409,In_590,In_835);
and U410 (N_410,In_905,In_32);
nand U411 (N_411,In_344,In_761);
and U412 (N_412,In_661,In_132);
and U413 (N_413,In_357,In_301);
or U414 (N_414,In_818,In_928);
nor U415 (N_415,In_918,In_42);
and U416 (N_416,In_319,In_595);
and U417 (N_417,In_728,In_550);
or U418 (N_418,In_409,In_866);
nor U419 (N_419,In_576,In_973);
nor U420 (N_420,In_755,In_669);
xor U421 (N_421,In_964,In_480);
nand U422 (N_422,In_484,In_778);
nand U423 (N_423,In_271,In_16);
and U424 (N_424,In_631,In_86);
or U425 (N_425,In_745,In_768);
xor U426 (N_426,In_348,In_963);
nor U427 (N_427,In_567,In_689);
or U428 (N_428,In_415,In_76);
or U429 (N_429,In_673,In_763);
nand U430 (N_430,In_451,In_363);
xnor U431 (N_431,In_947,In_697);
xor U432 (N_432,In_144,In_705);
and U433 (N_433,In_291,In_316);
nor U434 (N_434,In_309,In_832);
or U435 (N_435,In_15,In_390);
and U436 (N_436,In_917,In_40);
and U437 (N_437,In_325,In_563);
nor U438 (N_438,In_711,In_998);
and U439 (N_439,In_134,In_514);
nand U440 (N_440,In_193,In_505);
and U441 (N_441,In_373,In_907);
xor U442 (N_442,In_767,In_478);
or U443 (N_443,In_876,In_314);
xnor U444 (N_444,In_515,In_826);
nand U445 (N_445,In_84,In_703);
or U446 (N_446,In_816,In_502);
and U447 (N_447,In_611,In_635);
and U448 (N_448,In_864,In_214);
nor U449 (N_449,In_804,In_54);
or U450 (N_450,In_490,In_488);
or U451 (N_451,In_443,In_337);
and U452 (N_452,In_809,In_834);
nand U453 (N_453,In_796,In_548);
xor U454 (N_454,In_739,In_52);
nor U455 (N_455,In_808,In_55);
and U456 (N_456,In_557,In_113);
and U457 (N_457,In_664,In_461);
or U458 (N_458,In_679,In_934);
and U459 (N_459,In_367,In_22);
nor U460 (N_460,In_497,In_51);
xnor U461 (N_461,In_788,In_4);
and U462 (N_462,In_427,In_715);
nor U463 (N_463,In_59,In_600);
xnor U464 (N_464,In_843,In_396);
or U465 (N_465,In_388,In_303);
or U466 (N_466,In_760,In_151);
and U467 (N_467,In_580,In_430);
nor U468 (N_468,In_616,In_471);
nor U469 (N_469,In_477,In_169);
xor U470 (N_470,In_472,In_222);
xnor U471 (N_471,In_115,In_890);
xor U472 (N_472,In_933,In_441);
nor U473 (N_473,In_946,In_691);
nand U474 (N_474,In_504,In_573);
nor U475 (N_475,In_159,In_31);
or U476 (N_476,In_435,In_338);
nor U477 (N_477,In_626,In_26);
nand U478 (N_478,In_289,In_792);
or U479 (N_479,In_577,In_323);
nand U480 (N_480,In_201,In_566);
nor U481 (N_481,In_912,In_238);
or U482 (N_482,In_492,In_686);
xor U483 (N_483,In_452,In_807);
and U484 (N_484,In_442,In_968);
nor U485 (N_485,In_9,In_741);
and U486 (N_486,In_707,In_96);
nor U487 (N_487,In_997,In_355);
or U488 (N_488,In_171,In_56);
nor U489 (N_489,In_206,In_690);
xor U490 (N_490,In_66,In_116);
or U491 (N_491,In_197,In_667);
nor U492 (N_492,In_766,In_730);
or U493 (N_493,In_897,In_27);
nor U494 (N_494,In_896,In_294);
and U495 (N_495,In_459,In_35);
nand U496 (N_496,In_198,In_574);
nand U497 (N_497,In_29,In_60);
nand U498 (N_498,In_46,In_965);
or U499 (N_499,In_156,In_307);
or U500 (N_500,N_470,N_423);
nand U501 (N_501,N_38,N_124);
nand U502 (N_502,N_33,N_342);
nor U503 (N_503,N_94,N_223);
or U504 (N_504,N_491,N_200);
and U505 (N_505,N_61,N_156);
nand U506 (N_506,N_9,N_145);
and U507 (N_507,N_62,N_332);
and U508 (N_508,N_224,N_231);
and U509 (N_509,N_250,N_482);
and U510 (N_510,N_316,N_195);
or U511 (N_511,N_322,N_15);
and U512 (N_512,N_424,N_209);
nand U513 (N_513,N_432,N_306);
or U514 (N_514,N_259,N_274);
and U515 (N_515,N_139,N_166);
nor U516 (N_516,N_90,N_17);
or U517 (N_517,N_283,N_268);
and U518 (N_518,N_159,N_435);
and U519 (N_519,N_386,N_304);
nand U520 (N_520,N_144,N_468);
nor U521 (N_521,N_295,N_51);
or U522 (N_522,N_175,N_112);
or U523 (N_523,N_221,N_81);
or U524 (N_524,N_93,N_192);
nand U525 (N_525,N_198,N_457);
and U526 (N_526,N_392,N_31);
or U527 (N_527,N_217,N_148);
nand U528 (N_528,N_25,N_430);
and U529 (N_529,N_155,N_262);
nand U530 (N_530,N_480,N_187);
nand U531 (N_531,N_450,N_301);
xnor U532 (N_532,N_417,N_201);
and U533 (N_533,N_368,N_100);
nor U534 (N_534,N_47,N_460);
and U535 (N_535,N_142,N_133);
nor U536 (N_536,N_334,N_356);
nand U537 (N_537,N_179,N_22);
and U538 (N_538,N_205,N_70);
or U539 (N_539,N_140,N_255);
or U540 (N_540,N_481,N_411);
and U541 (N_541,N_445,N_13);
nor U542 (N_542,N_494,N_208);
xnor U543 (N_543,N_202,N_71);
nand U544 (N_544,N_357,N_349);
and U545 (N_545,N_110,N_354);
or U546 (N_546,N_26,N_101);
or U547 (N_547,N_266,N_163);
and U548 (N_548,N_92,N_136);
nor U549 (N_549,N_241,N_353);
or U550 (N_550,N_390,N_171);
nor U551 (N_551,N_331,N_337);
nand U552 (N_552,N_242,N_399);
or U553 (N_553,N_251,N_376);
nand U554 (N_554,N_203,N_225);
and U555 (N_555,N_279,N_77);
nor U556 (N_556,N_18,N_169);
nor U557 (N_557,N_496,N_109);
nor U558 (N_558,N_24,N_311);
nor U559 (N_559,N_436,N_219);
xor U560 (N_560,N_85,N_21);
and U561 (N_561,N_486,N_260);
or U562 (N_562,N_95,N_474);
xnor U563 (N_563,N_264,N_49);
nand U564 (N_564,N_74,N_405);
or U565 (N_565,N_455,N_389);
or U566 (N_566,N_193,N_267);
nand U567 (N_567,N_400,N_14);
nand U568 (N_568,N_104,N_382);
xnor U569 (N_569,N_226,N_106);
and U570 (N_570,N_293,N_84);
nand U571 (N_571,N_281,N_287);
or U572 (N_572,N_72,N_384);
and U573 (N_573,N_347,N_29);
nor U574 (N_574,N_157,N_324);
or U575 (N_575,N_8,N_442);
nand U576 (N_576,N_403,N_7);
nor U577 (N_577,N_477,N_20);
or U578 (N_578,N_387,N_302);
nor U579 (N_579,N_487,N_42);
and U580 (N_580,N_10,N_365);
and U581 (N_581,N_286,N_414);
nor U582 (N_582,N_359,N_53);
nor U583 (N_583,N_214,N_488);
or U584 (N_584,N_151,N_440);
and U585 (N_585,N_122,N_204);
nor U586 (N_586,N_495,N_48);
nor U587 (N_587,N_375,N_149);
nor U588 (N_588,N_63,N_235);
and U589 (N_589,N_465,N_352);
and U590 (N_590,N_1,N_383);
and U591 (N_591,N_165,N_75);
xor U592 (N_592,N_355,N_238);
nor U593 (N_593,N_314,N_37);
or U594 (N_594,N_11,N_466);
nand U595 (N_595,N_420,N_50);
and U596 (N_596,N_111,N_278);
nand U597 (N_597,N_248,N_408);
or U598 (N_598,N_303,N_164);
nor U599 (N_599,N_102,N_99);
and U600 (N_600,N_30,N_67);
and U601 (N_601,N_360,N_275);
nor U602 (N_602,N_190,N_391);
nand U603 (N_603,N_45,N_167);
and U604 (N_604,N_153,N_176);
nor U605 (N_605,N_98,N_146);
xnor U606 (N_606,N_451,N_59);
nand U607 (N_607,N_441,N_254);
or U608 (N_608,N_426,N_128);
nor U609 (N_609,N_103,N_310);
and U610 (N_610,N_173,N_464);
or U611 (N_611,N_458,N_229);
nor U612 (N_612,N_317,N_401);
nand U613 (N_613,N_256,N_177);
nor U614 (N_614,N_215,N_207);
nor U615 (N_615,N_479,N_340);
and U616 (N_616,N_107,N_449);
and U617 (N_617,N_294,N_469);
and U618 (N_618,N_498,N_291);
or U619 (N_619,N_427,N_380);
and U620 (N_620,N_315,N_454);
nor U621 (N_621,N_80,N_227);
and U622 (N_622,N_330,N_258);
nand U623 (N_623,N_65,N_213);
nand U624 (N_624,N_196,N_237);
and U625 (N_625,N_188,N_409);
or U626 (N_626,N_270,N_467);
and U627 (N_627,N_378,N_485);
and U628 (N_628,N_448,N_497);
and U629 (N_629,N_117,N_152);
nand U630 (N_630,N_41,N_350);
nor U631 (N_631,N_232,N_483);
nor U632 (N_632,N_446,N_170);
or U633 (N_633,N_406,N_425);
nand U634 (N_634,N_431,N_174);
or U635 (N_635,N_141,N_361);
nand U636 (N_636,N_397,N_318);
xor U637 (N_637,N_341,N_396);
or U638 (N_638,N_308,N_12);
or U639 (N_639,N_381,N_277);
or U640 (N_640,N_407,N_27);
nor U641 (N_641,N_273,N_116);
nand U642 (N_642,N_313,N_57);
nand U643 (N_643,N_476,N_276);
nor U644 (N_644,N_16,N_183);
or U645 (N_645,N_484,N_364);
and U646 (N_646,N_39,N_210);
and U647 (N_647,N_97,N_66);
xnor U648 (N_648,N_3,N_114);
xnor U649 (N_649,N_121,N_263);
or U650 (N_650,N_249,N_125);
xnor U651 (N_651,N_108,N_394);
nor U652 (N_652,N_373,N_312);
or U653 (N_653,N_76,N_447);
xnor U654 (N_654,N_158,N_300);
nor U655 (N_655,N_351,N_46);
or U656 (N_656,N_393,N_118);
nor U657 (N_657,N_82,N_284);
nor U658 (N_658,N_43,N_191);
and U659 (N_659,N_410,N_135);
or U660 (N_660,N_490,N_309);
nor U661 (N_661,N_197,N_4);
nor U662 (N_662,N_105,N_222);
nand U663 (N_663,N_182,N_216);
and U664 (N_664,N_186,N_147);
nor U665 (N_665,N_272,N_325);
nand U666 (N_666,N_280,N_64);
and U667 (N_667,N_385,N_126);
nand U668 (N_668,N_473,N_32);
or U669 (N_669,N_138,N_185);
nand U670 (N_670,N_419,N_23);
nand U671 (N_671,N_434,N_245);
nor U672 (N_672,N_438,N_194);
nor U673 (N_673,N_437,N_404);
nor U674 (N_674,N_86,N_132);
or U675 (N_675,N_478,N_181);
xor U676 (N_676,N_444,N_292);
or U677 (N_677,N_492,N_162);
nand U678 (N_678,N_69,N_243);
and U679 (N_679,N_459,N_150);
nor U680 (N_680,N_5,N_338);
and U681 (N_681,N_246,N_367);
or U682 (N_682,N_297,N_344);
or U683 (N_683,N_79,N_180);
nor U684 (N_684,N_346,N_253);
and U685 (N_685,N_233,N_199);
or U686 (N_686,N_78,N_35);
xor U687 (N_687,N_339,N_115);
or U688 (N_688,N_230,N_168);
or U689 (N_689,N_271,N_240);
nor U690 (N_690,N_19,N_370);
xnor U691 (N_691,N_36,N_265);
nor U692 (N_692,N_299,N_44);
nand U693 (N_693,N_113,N_239);
xnor U694 (N_694,N_307,N_73);
and U695 (N_695,N_369,N_212);
nor U696 (N_696,N_422,N_456);
or U697 (N_697,N_261,N_91);
nand U698 (N_698,N_320,N_285);
or U699 (N_699,N_123,N_358);
nor U700 (N_700,N_362,N_34);
and U701 (N_701,N_96,N_333);
or U702 (N_702,N_211,N_402);
or U703 (N_703,N_429,N_335);
and U704 (N_704,N_366,N_178);
nand U705 (N_705,N_433,N_160);
and U706 (N_706,N_374,N_323);
nor U707 (N_707,N_257,N_372);
nor U708 (N_708,N_28,N_119);
xor U709 (N_709,N_172,N_443);
xnor U710 (N_710,N_412,N_290);
xor U711 (N_711,N_413,N_415);
nand U712 (N_712,N_418,N_54);
and U713 (N_713,N_252,N_471);
nand U714 (N_714,N_439,N_452);
or U715 (N_715,N_56,N_234);
or U716 (N_716,N_395,N_2);
nor U717 (N_717,N_329,N_0);
nor U718 (N_718,N_120,N_220);
and U719 (N_719,N_282,N_428);
or U720 (N_720,N_89,N_298);
or U721 (N_721,N_244,N_377);
nor U722 (N_722,N_60,N_83);
nand U723 (N_723,N_475,N_247);
or U724 (N_724,N_345,N_453);
or U725 (N_725,N_462,N_161);
and U726 (N_726,N_489,N_130);
or U727 (N_727,N_305,N_236);
nor U728 (N_728,N_371,N_6);
or U729 (N_729,N_58,N_319);
or U730 (N_730,N_87,N_134);
nor U731 (N_731,N_137,N_129);
nand U732 (N_732,N_52,N_55);
and U733 (N_733,N_228,N_421);
nor U734 (N_734,N_326,N_68);
nor U735 (N_735,N_184,N_321);
or U736 (N_736,N_363,N_461);
nand U737 (N_737,N_398,N_343);
or U738 (N_738,N_388,N_288);
nand U739 (N_739,N_88,N_206);
and U740 (N_740,N_493,N_499);
nor U741 (N_741,N_472,N_269);
nor U742 (N_742,N_336,N_328);
nand U743 (N_743,N_379,N_218);
xnor U744 (N_744,N_289,N_127);
and U745 (N_745,N_327,N_189);
or U746 (N_746,N_143,N_296);
nor U747 (N_747,N_348,N_154);
or U748 (N_748,N_463,N_416);
nand U749 (N_749,N_131,N_40);
nand U750 (N_750,N_427,N_374);
or U751 (N_751,N_309,N_117);
or U752 (N_752,N_442,N_23);
nand U753 (N_753,N_398,N_16);
nand U754 (N_754,N_285,N_356);
nor U755 (N_755,N_278,N_323);
and U756 (N_756,N_136,N_488);
nor U757 (N_757,N_337,N_131);
nor U758 (N_758,N_348,N_400);
xor U759 (N_759,N_423,N_414);
and U760 (N_760,N_181,N_138);
nor U761 (N_761,N_208,N_499);
or U762 (N_762,N_66,N_31);
or U763 (N_763,N_105,N_330);
nor U764 (N_764,N_481,N_382);
nor U765 (N_765,N_64,N_461);
nor U766 (N_766,N_357,N_322);
and U767 (N_767,N_100,N_485);
or U768 (N_768,N_389,N_346);
nor U769 (N_769,N_454,N_249);
or U770 (N_770,N_403,N_118);
or U771 (N_771,N_120,N_169);
and U772 (N_772,N_259,N_449);
and U773 (N_773,N_384,N_252);
nor U774 (N_774,N_40,N_95);
or U775 (N_775,N_71,N_447);
nand U776 (N_776,N_413,N_339);
and U777 (N_777,N_72,N_190);
and U778 (N_778,N_79,N_213);
and U779 (N_779,N_102,N_184);
nand U780 (N_780,N_458,N_392);
nand U781 (N_781,N_471,N_419);
or U782 (N_782,N_440,N_289);
nor U783 (N_783,N_207,N_481);
and U784 (N_784,N_194,N_300);
or U785 (N_785,N_393,N_141);
nand U786 (N_786,N_298,N_354);
or U787 (N_787,N_109,N_280);
and U788 (N_788,N_333,N_111);
nor U789 (N_789,N_341,N_215);
nor U790 (N_790,N_428,N_223);
and U791 (N_791,N_234,N_132);
xor U792 (N_792,N_48,N_139);
nor U793 (N_793,N_365,N_368);
and U794 (N_794,N_212,N_320);
nor U795 (N_795,N_199,N_472);
and U796 (N_796,N_139,N_271);
xor U797 (N_797,N_452,N_133);
xor U798 (N_798,N_401,N_125);
or U799 (N_799,N_92,N_83);
and U800 (N_800,N_287,N_104);
nor U801 (N_801,N_347,N_295);
xnor U802 (N_802,N_399,N_96);
xnor U803 (N_803,N_465,N_208);
xor U804 (N_804,N_290,N_79);
or U805 (N_805,N_408,N_16);
nand U806 (N_806,N_1,N_124);
nand U807 (N_807,N_292,N_61);
xnor U808 (N_808,N_35,N_86);
and U809 (N_809,N_296,N_18);
xnor U810 (N_810,N_447,N_260);
or U811 (N_811,N_210,N_154);
xnor U812 (N_812,N_381,N_78);
nor U813 (N_813,N_228,N_441);
nor U814 (N_814,N_12,N_49);
or U815 (N_815,N_478,N_414);
nand U816 (N_816,N_140,N_213);
and U817 (N_817,N_287,N_397);
nand U818 (N_818,N_348,N_143);
and U819 (N_819,N_485,N_429);
and U820 (N_820,N_112,N_405);
or U821 (N_821,N_377,N_449);
or U822 (N_822,N_166,N_263);
and U823 (N_823,N_438,N_165);
nor U824 (N_824,N_183,N_107);
and U825 (N_825,N_17,N_162);
and U826 (N_826,N_404,N_386);
nand U827 (N_827,N_203,N_71);
and U828 (N_828,N_182,N_283);
nor U829 (N_829,N_486,N_213);
and U830 (N_830,N_96,N_227);
or U831 (N_831,N_261,N_434);
or U832 (N_832,N_206,N_55);
xor U833 (N_833,N_212,N_172);
and U834 (N_834,N_376,N_446);
nor U835 (N_835,N_88,N_111);
nor U836 (N_836,N_323,N_327);
or U837 (N_837,N_236,N_13);
nand U838 (N_838,N_70,N_159);
nor U839 (N_839,N_419,N_104);
or U840 (N_840,N_64,N_482);
nor U841 (N_841,N_411,N_463);
or U842 (N_842,N_361,N_203);
or U843 (N_843,N_478,N_410);
xor U844 (N_844,N_190,N_266);
nand U845 (N_845,N_439,N_300);
and U846 (N_846,N_221,N_252);
and U847 (N_847,N_334,N_253);
and U848 (N_848,N_290,N_11);
or U849 (N_849,N_381,N_170);
or U850 (N_850,N_370,N_122);
or U851 (N_851,N_299,N_319);
and U852 (N_852,N_373,N_383);
and U853 (N_853,N_102,N_273);
nor U854 (N_854,N_77,N_416);
or U855 (N_855,N_477,N_378);
and U856 (N_856,N_171,N_5);
nor U857 (N_857,N_381,N_416);
and U858 (N_858,N_448,N_246);
nand U859 (N_859,N_325,N_263);
nor U860 (N_860,N_274,N_413);
or U861 (N_861,N_278,N_191);
nor U862 (N_862,N_206,N_195);
and U863 (N_863,N_144,N_110);
nand U864 (N_864,N_4,N_473);
and U865 (N_865,N_475,N_471);
xor U866 (N_866,N_445,N_357);
nand U867 (N_867,N_330,N_312);
nand U868 (N_868,N_254,N_53);
nor U869 (N_869,N_50,N_107);
and U870 (N_870,N_485,N_83);
and U871 (N_871,N_353,N_196);
nor U872 (N_872,N_421,N_403);
and U873 (N_873,N_481,N_206);
or U874 (N_874,N_249,N_132);
nand U875 (N_875,N_331,N_416);
nand U876 (N_876,N_483,N_394);
nor U877 (N_877,N_347,N_350);
and U878 (N_878,N_384,N_374);
or U879 (N_879,N_38,N_240);
xor U880 (N_880,N_447,N_125);
or U881 (N_881,N_316,N_258);
or U882 (N_882,N_419,N_264);
or U883 (N_883,N_136,N_385);
or U884 (N_884,N_476,N_149);
and U885 (N_885,N_164,N_113);
and U886 (N_886,N_323,N_315);
and U887 (N_887,N_65,N_230);
nor U888 (N_888,N_226,N_492);
and U889 (N_889,N_264,N_278);
nor U890 (N_890,N_402,N_461);
or U891 (N_891,N_38,N_27);
xnor U892 (N_892,N_160,N_314);
nand U893 (N_893,N_269,N_283);
or U894 (N_894,N_344,N_286);
nor U895 (N_895,N_470,N_455);
nor U896 (N_896,N_426,N_149);
xnor U897 (N_897,N_425,N_80);
nand U898 (N_898,N_441,N_65);
and U899 (N_899,N_322,N_405);
xor U900 (N_900,N_26,N_412);
nand U901 (N_901,N_192,N_472);
or U902 (N_902,N_26,N_252);
or U903 (N_903,N_228,N_265);
nand U904 (N_904,N_266,N_7);
and U905 (N_905,N_141,N_434);
and U906 (N_906,N_144,N_56);
or U907 (N_907,N_268,N_412);
and U908 (N_908,N_219,N_310);
and U909 (N_909,N_275,N_451);
nor U910 (N_910,N_117,N_3);
xor U911 (N_911,N_453,N_480);
xor U912 (N_912,N_304,N_336);
and U913 (N_913,N_469,N_349);
or U914 (N_914,N_198,N_101);
nor U915 (N_915,N_72,N_36);
and U916 (N_916,N_327,N_264);
or U917 (N_917,N_83,N_367);
or U918 (N_918,N_352,N_275);
nor U919 (N_919,N_40,N_402);
or U920 (N_920,N_409,N_266);
nand U921 (N_921,N_399,N_168);
nor U922 (N_922,N_349,N_245);
nor U923 (N_923,N_332,N_82);
nand U924 (N_924,N_233,N_485);
or U925 (N_925,N_355,N_394);
nor U926 (N_926,N_401,N_283);
and U927 (N_927,N_344,N_16);
nand U928 (N_928,N_423,N_438);
nor U929 (N_929,N_219,N_396);
and U930 (N_930,N_271,N_396);
or U931 (N_931,N_398,N_331);
nand U932 (N_932,N_232,N_83);
and U933 (N_933,N_258,N_95);
nand U934 (N_934,N_366,N_243);
nand U935 (N_935,N_318,N_165);
nand U936 (N_936,N_58,N_228);
nor U937 (N_937,N_227,N_220);
or U938 (N_938,N_133,N_316);
or U939 (N_939,N_198,N_37);
nand U940 (N_940,N_44,N_406);
nand U941 (N_941,N_417,N_432);
or U942 (N_942,N_130,N_160);
nand U943 (N_943,N_125,N_320);
nand U944 (N_944,N_3,N_156);
nand U945 (N_945,N_248,N_415);
and U946 (N_946,N_213,N_47);
and U947 (N_947,N_89,N_421);
nor U948 (N_948,N_246,N_284);
nand U949 (N_949,N_272,N_25);
or U950 (N_950,N_443,N_62);
or U951 (N_951,N_189,N_9);
nor U952 (N_952,N_54,N_203);
and U953 (N_953,N_59,N_211);
or U954 (N_954,N_340,N_186);
nand U955 (N_955,N_225,N_191);
or U956 (N_956,N_462,N_100);
or U957 (N_957,N_124,N_444);
and U958 (N_958,N_217,N_9);
nand U959 (N_959,N_188,N_258);
or U960 (N_960,N_224,N_436);
or U961 (N_961,N_183,N_491);
xnor U962 (N_962,N_281,N_400);
nand U963 (N_963,N_242,N_186);
and U964 (N_964,N_21,N_86);
or U965 (N_965,N_227,N_477);
nand U966 (N_966,N_480,N_110);
nor U967 (N_967,N_300,N_221);
and U968 (N_968,N_246,N_345);
nor U969 (N_969,N_491,N_107);
xnor U970 (N_970,N_354,N_174);
and U971 (N_971,N_177,N_267);
nand U972 (N_972,N_192,N_273);
or U973 (N_973,N_279,N_343);
nor U974 (N_974,N_380,N_445);
and U975 (N_975,N_453,N_438);
nand U976 (N_976,N_154,N_88);
nand U977 (N_977,N_255,N_246);
xor U978 (N_978,N_226,N_387);
xnor U979 (N_979,N_454,N_442);
nor U980 (N_980,N_344,N_293);
nor U981 (N_981,N_220,N_311);
nor U982 (N_982,N_81,N_167);
and U983 (N_983,N_129,N_152);
nand U984 (N_984,N_137,N_69);
and U985 (N_985,N_483,N_244);
nand U986 (N_986,N_392,N_107);
nand U987 (N_987,N_125,N_109);
nor U988 (N_988,N_130,N_231);
or U989 (N_989,N_69,N_172);
or U990 (N_990,N_439,N_19);
nand U991 (N_991,N_250,N_193);
nand U992 (N_992,N_111,N_328);
nor U993 (N_993,N_264,N_416);
nand U994 (N_994,N_239,N_192);
or U995 (N_995,N_85,N_290);
and U996 (N_996,N_467,N_116);
and U997 (N_997,N_315,N_56);
and U998 (N_998,N_97,N_258);
nand U999 (N_999,N_342,N_176);
nand U1000 (N_1000,N_724,N_863);
nor U1001 (N_1001,N_791,N_541);
and U1002 (N_1002,N_554,N_900);
xnor U1003 (N_1003,N_779,N_747);
and U1004 (N_1004,N_611,N_607);
or U1005 (N_1005,N_754,N_620);
nor U1006 (N_1006,N_929,N_512);
or U1007 (N_1007,N_557,N_540);
or U1008 (N_1008,N_957,N_521);
nand U1009 (N_1009,N_684,N_789);
or U1010 (N_1010,N_768,N_725);
and U1011 (N_1011,N_567,N_928);
and U1012 (N_1012,N_905,N_907);
nand U1013 (N_1013,N_654,N_617);
or U1014 (N_1014,N_920,N_822);
and U1015 (N_1015,N_819,N_872);
nor U1016 (N_1016,N_689,N_665);
xnor U1017 (N_1017,N_785,N_629);
or U1018 (N_1018,N_733,N_579);
or U1019 (N_1019,N_535,N_896);
and U1020 (N_1020,N_833,N_519);
and U1021 (N_1021,N_530,N_534);
xor U1022 (N_1022,N_693,N_569);
and U1023 (N_1023,N_542,N_827);
xnor U1024 (N_1024,N_606,N_637);
nor U1025 (N_1025,N_808,N_630);
or U1026 (N_1026,N_628,N_998);
nand U1027 (N_1027,N_784,N_953);
and U1028 (N_1028,N_644,N_758);
or U1029 (N_1029,N_986,N_802);
and U1030 (N_1030,N_522,N_775);
nand U1031 (N_1031,N_846,N_858);
xnor U1032 (N_1032,N_767,N_887);
xor U1033 (N_1033,N_918,N_824);
nand U1034 (N_1034,N_925,N_742);
nor U1035 (N_1035,N_596,N_837);
xnor U1036 (N_1036,N_520,N_993);
nor U1037 (N_1037,N_972,N_695);
nor U1038 (N_1038,N_717,N_729);
and U1039 (N_1039,N_648,N_865);
and U1040 (N_1040,N_773,N_755);
nand U1041 (N_1041,N_726,N_781);
nor U1042 (N_1042,N_828,N_801);
or U1043 (N_1043,N_966,N_978);
and U1044 (N_1044,N_680,N_658);
and U1045 (N_1045,N_963,N_983);
and U1046 (N_1046,N_692,N_585);
or U1047 (N_1047,N_832,N_575);
nand U1048 (N_1048,N_533,N_503);
nor U1049 (N_1049,N_732,N_968);
nor U1050 (N_1050,N_964,N_634);
nor U1051 (N_1051,N_645,N_715);
nor U1052 (N_1052,N_514,N_669);
and U1053 (N_1053,N_656,N_593);
and U1054 (N_1054,N_804,N_947);
or U1055 (N_1055,N_690,N_805);
nand U1056 (N_1056,N_627,N_948);
and U1057 (N_1057,N_753,N_651);
nand U1058 (N_1058,N_867,N_763);
nand U1059 (N_1059,N_639,N_696);
xor U1060 (N_1060,N_967,N_549);
nor U1061 (N_1061,N_958,N_675);
nor U1062 (N_1062,N_803,N_756);
nor U1063 (N_1063,N_746,N_860);
and U1064 (N_1064,N_699,N_547);
nor U1065 (N_1065,N_550,N_952);
xnor U1066 (N_1066,N_762,N_788);
or U1067 (N_1067,N_727,N_838);
and U1068 (N_1068,N_839,N_577);
or U1069 (N_1069,N_818,N_647);
or U1070 (N_1070,N_600,N_940);
or U1071 (N_1071,N_643,N_590);
xor U1072 (N_1072,N_605,N_594);
nor U1073 (N_1073,N_744,N_899);
xnor U1074 (N_1074,N_850,N_633);
or U1075 (N_1075,N_677,N_506);
nand U1076 (N_1076,N_661,N_795);
xnor U1077 (N_1077,N_987,N_570);
nand U1078 (N_1078,N_636,N_553);
or U1079 (N_1079,N_708,N_868);
nand U1080 (N_1080,N_923,N_769);
and U1081 (N_1081,N_843,N_602);
or U1082 (N_1082,N_613,N_668);
and U1083 (N_1083,N_616,N_556);
or U1084 (N_1084,N_826,N_861);
xor U1085 (N_1085,N_965,N_780);
and U1086 (N_1086,N_580,N_676);
xor U1087 (N_1087,N_825,N_912);
or U1088 (N_1088,N_854,N_943);
nor U1089 (N_1089,N_956,N_815);
or U1090 (N_1090,N_977,N_621);
nor U1091 (N_1091,N_908,N_848);
and U1092 (N_1092,N_700,N_578);
nor U1093 (N_1093,N_904,N_510);
and U1094 (N_1094,N_862,N_745);
nand U1095 (N_1095,N_853,N_683);
nor U1096 (N_1096,N_612,N_897);
xnor U1097 (N_1097,N_845,N_710);
nor U1098 (N_1098,N_945,N_551);
and U1099 (N_1099,N_974,N_513);
nor U1100 (N_1100,N_697,N_875);
nor U1101 (N_1101,N_632,N_841);
nand U1102 (N_1102,N_794,N_990);
or U1103 (N_1103,N_873,N_704);
nand U1104 (N_1104,N_735,N_609);
or U1105 (N_1105,N_691,N_881);
nor U1106 (N_1106,N_852,N_524);
and U1107 (N_1107,N_812,N_979);
nand U1108 (N_1108,N_538,N_976);
or U1109 (N_1109,N_561,N_576);
nand U1110 (N_1110,N_910,N_663);
xor U1111 (N_1111,N_688,N_523);
xnor U1112 (N_1112,N_934,N_572);
or U1113 (N_1113,N_831,N_619);
nand U1114 (N_1114,N_568,N_529);
nor U1115 (N_1115,N_664,N_526);
and U1116 (N_1116,N_652,N_624);
nand U1117 (N_1117,N_749,N_674);
nor U1118 (N_1118,N_807,N_936);
xnor U1119 (N_1119,N_573,N_728);
nand U1120 (N_1120,N_716,N_844);
and U1121 (N_1121,N_703,N_739);
and U1122 (N_1122,N_618,N_882);
and U1123 (N_1123,N_558,N_653);
or U1124 (N_1124,N_518,N_545);
nand U1125 (N_1125,N_913,N_714);
nand U1126 (N_1126,N_811,N_723);
nor U1127 (N_1127,N_750,N_552);
or U1128 (N_1128,N_614,N_893);
nor U1129 (N_1129,N_991,N_537);
and U1130 (N_1130,N_751,N_973);
nand U1131 (N_1131,N_597,N_820);
nor U1132 (N_1132,N_625,N_851);
nor U1133 (N_1133,N_626,N_711);
nor U1134 (N_1134,N_980,N_766);
or U1135 (N_1135,N_996,N_919);
or U1136 (N_1136,N_989,N_702);
nor U1137 (N_1137,N_588,N_984);
nand U1138 (N_1138,N_835,N_640);
xor U1139 (N_1139,N_603,N_836);
nand U1140 (N_1140,N_884,N_687);
nor U1141 (N_1141,N_581,N_760);
or U1142 (N_1142,N_938,N_536);
and U1143 (N_1143,N_571,N_840);
or U1144 (N_1144,N_981,N_604);
nand U1145 (N_1145,N_685,N_796);
and U1146 (N_1146,N_646,N_810);
or U1147 (N_1147,N_608,N_902);
or U1148 (N_1148,N_871,N_511);
nor U1149 (N_1149,N_829,N_988);
nor U1150 (N_1150,N_741,N_515);
nor U1151 (N_1151,N_666,N_921);
or U1152 (N_1152,N_670,N_889);
and U1153 (N_1153,N_731,N_813);
xnor U1154 (N_1154,N_774,N_792);
nand U1155 (N_1155,N_587,N_894);
and U1156 (N_1156,N_941,N_713);
or U1157 (N_1157,N_926,N_525);
or U1158 (N_1158,N_888,N_939);
nor U1159 (N_1159,N_660,N_992);
nor U1160 (N_1160,N_857,N_761);
and U1161 (N_1161,N_599,N_673);
nor U1162 (N_1162,N_771,N_949);
and U1163 (N_1163,N_903,N_916);
nand U1164 (N_1164,N_517,N_866);
nor U1165 (N_1165,N_583,N_759);
nand U1166 (N_1166,N_917,N_950);
nand U1167 (N_1167,N_649,N_642);
nand U1168 (N_1168,N_961,N_969);
nand U1169 (N_1169,N_707,N_922);
and U1170 (N_1170,N_622,N_722);
nand U1171 (N_1171,N_999,N_730);
nand U1172 (N_1172,N_752,N_705);
or U1173 (N_1173,N_584,N_864);
and U1174 (N_1174,N_712,N_778);
nor U1175 (N_1175,N_890,N_662);
nand U1176 (N_1176,N_507,N_698);
or U1177 (N_1177,N_994,N_772);
or U1178 (N_1178,N_886,N_876);
xor U1179 (N_1179,N_847,N_859);
or U1180 (N_1180,N_738,N_586);
nor U1181 (N_1181,N_931,N_709);
or U1182 (N_1182,N_532,N_719);
and U1183 (N_1183,N_849,N_798);
and U1184 (N_1184,N_623,N_564);
nor U1185 (N_1185,N_869,N_959);
or U1186 (N_1186,N_935,N_615);
xnor U1187 (N_1187,N_874,N_898);
nor U1188 (N_1188,N_951,N_982);
nor U1189 (N_1189,N_560,N_672);
or U1190 (N_1190,N_901,N_782);
nor U1191 (N_1191,N_544,N_933);
xnor U1192 (N_1192,N_659,N_793);
or U1193 (N_1193,N_679,N_914);
or U1194 (N_1194,N_591,N_505);
or U1195 (N_1195,N_770,N_531);
or U1196 (N_1196,N_806,N_800);
nand U1197 (N_1197,N_955,N_944);
and U1198 (N_1198,N_790,N_574);
nor U1199 (N_1199,N_543,N_870);
and U1200 (N_1200,N_765,N_721);
and U1201 (N_1201,N_821,N_786);
nor U1202 (N_1202,N_635,N_878);
nor U1203 (N_1203,N_816,N_509);
nor U1204 (N_1204,N_809,N_682);
nand U1205 (N_1205,N_971,N_641);
or U1206 (N_1206,N_748,N_823);
nand U1207 (N_1207,N_880,N_592);
or U1208 (N_1208,N_962,N_678);
and U1209 (N_1209,N_527,N_906);
nand U1210 (N_1210,N_638,N_909);
and U1211 (N_1211,N_559,N_814);
or U1212 (N_1212,N_856,N_565);
nor U1213 (N_1213,N_997,N_650);
xor U1214 (N_1214,N_501,N_667);
nand U1215 (N_1215,N_671,N_582);
or U1216 (N_1216,N_927,N_995);
or U1217 (N_1217,N_891,N_942);
nor U1218 (N_1218,N_970,N_508);
and U1219 (N_1219,N_743,N_783);
xor U1220 (N_1220,N_842,N_734);
nand U1221 (N_1221,N_694,N_706);
nand U1222 (N_1222,N_776,N_657);
nand U1223 (N_1223,N_548,N_937);
or U1224 (N_1224,N_855,N_892);
nand U1225 (N_1225,N_566,N_834);
xor U1226 (N_1226,N_879,N_830);
xor U1227 (N_1227,N_777,N_799);
nor U1228 (N_1228,N_562,N_817);
nor U1229 (N_1229,N_504,N_655);
nand U1230 (N_1230,N_555,N_764);
or U1231 (N_1231,N_500,N_895);
and U1232 (N_1232,N_701,N_502);
nand U1233 (N_1233,N_631,N_610);
and U1234 (N_1234,N_930,N_954);
and U1235 (N_1235,N_528,N_563);
and U1236 (N_1236,N_595,N_681);
nor U1237 (N_1237,N_598,N_546);
nand U1238 (N_1238,N_985,N_975);
xnor U1239 (N_1239,N_757,N_797);
and U1240 (N_1240,N_883,N_946);
and U1241 (N_1241,N_911,N_877);
nand U1242 (N_1242,N_924,N_686);
nand U1243 (N_1243,N_539,N_601);
nand U1244 (N_1244,N_740,N_915);
nand U1245 (N_1245,N_885,N_589);
nor U1246 (N_1246,N_787,N_736);
nor U1247 (N_1247,N_737,N_516);
nor U1248 (N_1248,N_720,N_718);
or U1249 (N_1249,N_932,N_960);
nor U1250 (N_1250,N_595,N_661);
and U1251 (N_1251,N_556,N_784);
nor U1252 (N_1252,N_669,N_946);
or U1253 (N_1253,N_636,N_843);
nand U1254 (N_1254,N_517,N_547);
and U1255 (N_1255,N_781,N_836);
or U1256 (N_1256,N_731,N_710);
nand U1257 (N_1257,N_752,N_519);
and U1258 (N_1258,N_878,N_632);
nor U1259 (N_1259,N_845,N_708);
nand U1260 (N_1260,N_643,N_945);
and U1261 (N_1261,N_510,N_963);
and U1262 (N_1262,N_605,N_892);
xnor U1263 (N_1263,N_990,N_703);
nand U1264 (N_1264,N_761,N_851);
or U1265 (N_1265,N_967,N_921);
nand U1266 (N_1266,N_755,N_625);
nand U1267 (N_1267,N_661,N_966);
nand U1268 (N_1268,N_803,N_833);
or U1269 (N_1269,N_744,N_727);
or U1270 (N_1270,N_545,N_899);
and U1271 (N_1271,N_626,N_873);
and U1272 (N_1272,N_663,N_658);
or U1273 (N_1273,N_766,N_718);
nand U1274 (N_1274,N_752,N_731);
and U1275 (N_1275,N_550,N_601);
nand U1276 (N_1276,N_702,N_874);
nand U1277 (N_1277,N_816,N_580);
nand U1278 (N_1278,N_819,N_793);
or U1279 (N_1279,N_814,N_890);
or U1280 (N_1280,N_965,N_575);
xnor U1281 (N_1281,N_914,N_778);
nand U1282 (N_1282,N_590,N_551);
nand U1283 (N_1283,N_955,N_961);
or U1284 (N_1284,N_585,N_673);
nand U1285 (N_1285,N_756,N_677);
and U1286 (N_1286,N_751,N_675);
nor U1287 (N_1287,N_715,N_523);
and U1288 (N_1288,N_723,N_745);
and U1289 (N_1289,N_749,N_967);
nor U1290 (N_1290,N_999,N_676);
and U1291 (N_1291,N_791,N_770);
nor U1292 (N_1292,N_930,N_908);
and U1293 (N_1293,N_579,N_939);
and U1294 (N_1294,N_689,N_925);
nand U1295 (N_1295,N_935,N_910);
nand U1296 (N_1296,N_811,N_842);
nand U1297 (N_1297,N_581,N_880);
xor U1298 (N_1298,N_835,N_904);
nor U1299 (N_1299,N_929,N_554);
and U1300 (N_1300,N_755,N_731);
nor U1301 (N_1301,N_966,N_544);
and U1302 (N_1302,N_753,N_927);
xnor U1303 (N_1303,N_942,N_902);
nand U1304 (N_1304,N_706,N_968);
nand U1305 (N_1305,N_730,N_848);
or U1306 (N_1306,N_932,N_921);
or U1307 (N_1307,N_962,N_681);
nand U1308 (N_1308,N_731,N_505);
and U1309 (N_1309,N_750,N_824);
nor U1310 (N_1310,N_748,N_816);
and U1311 (N_1311,N_984,N_986);
xor U1312 (N_1312,N_948,N_942);
and U1313 (N_1313,N_747,N_626);
and U1314 (N_1314,N_753,N_551);
or U1315 (N_1315,N_520,N_981);
nor U1316 (N_1316,N_790,N_874);
nand U1317 (N_1317,N_512,N_607);
or U1318 (N_1318,N_659,N_877);
nor U1319 (N_1319,N_669,N_535);
and U1320 (N_1320,N_962,N_851);
nand U1321 (N_1321,N_549,N_921);
nand U1322 (N_1322,N_924,N_834);
xor U1323 (N_1323,N_795,N_543);
nor U1324 (N_1324,N_961,N_844);
nor U1325 (N_1325,N_989,N_877);
nand U1326 (N_1326,N_997,N_582);
or U1327 (N_1327,N_903,N_582);
and U1328 (N_1328,N_652,N_889);
nand U1329 (N_1329,N_967,N_702);
and U1330 (N_1330,N_691,N_833);
xnor U1331 (N_1331,N_972,N_648);
nand U1332 (N_1332,N_727,N_628);
or U1333 (N_1333,N_669,N_628);
xor U1334 (N_1334,N_856,N_744);
or U1335 (N_1335,N_773,N_850);
nand U1336 (N_1336,N_617,N_866);
and U1337 (N_1337,N_661,N_897);
nor U1338 (N_1338,N_794,N_638);
and U1339 (N_1339,N_863,N_752);
xnor U1340 (N_1340,N_699,N_608);
nor U1341 (N_1341,N_871,N_994);
nor U1342 (N_1342,N_992,N_784);
nor U1343 (N_1343,N_606,N_561);
xor U1344 (N_1344,N_973,N_502);
nand U1345 (N_1345,N_922,N_663);
and U1346 (N_1346,N_574,N_575);
or U1347 (N_1347,N_587,N_688);
or U1348 (N_1348,N_906,N_944);
and U1349 (N_1349,N_987,N_821);
nand U1350 (N_1350,N_613,N_954);
nor U1351 (N_1351,N_998,N_891);
nand U1352 (N_1352,N_648,N_615);
and U1353 (N_1353,N_904,N_936);
or U1354 (N_1354,N_652,N_816);
or U1355 (N_1355,N_533,N_884);
nand U1356 (N_1356,N_538,N_884);
xnor U1357 (N_1357,N_917,N_610);
and U1358 (N_1358,N_875,N_587);
xor U1359 (N_1359,N_532,N_511);
or U1360 (N_1360,N_895,N_878);
and U1361 (N_1361,N_994,N_604);
nand U1362 (N_1362,N_578,N_905);
or U1363 (N_1363,N_907,N_780);
nor U1364 (N_1364,N_518,N_891);
xor U1365 (N_1365,N_745,N_567);
or U1366 (N_1366,N_965,N_805);
or U1367 (N_1367,N_657,N_717);
and U1368 (N_1368,N_713,N_507);
nand U1369 (N_1369,N_546,N_783);
nor U1370 (N_1370,N_627,N_962);
and U1371 (N_1371,N_586,N_516);
xnor U1372 (N_1372,N_868,N_982);
nor U1373 (N_1373,N_563,N_577);
and U1374 (N_1374,N_640,N_563);
or U1375 (N_1375,N_953,N_840);
or U1376 (N_1376,N_684,N_918);
nor U1377 (N_1377,N_701,N_797);
nand U1378 (N_1378,N_704,N_653);
or U1379 (N_1379,N_824,N_683);
and U1380 (N_1380,N_586,N_841);
or U1381 (N_1381,N_572,N_893);
nand U1382 (N_1382,N_787,N_802);
nand U1383 (N_1383,N_782,N_551);
or U1384 (N_1384,N_974,N_782);
or U1385 (N_1385,N_697,N_676);
and U1386 (N_1386,N_703,N_870);
xnor U1387 (N_1387,N_533,N_622);
nand U1388 (N_1388,N_842,N_973);
nand U1389 (N_1389,N_596,N_834);
or U1390 (N_1390,N_654,N_979);
nand U1391 (N_1391,N_877,N_907);
nand U1392 (N_1392,N_708,N_680);
nor U1393 (N_1393,N_578,N_546);
nand U1394 (N_1394,N_892,N_548);
and U1395 (N_1395,N_659,N_530);
nor U1396 (N_1396,N_814,N_813);
and U1397 (N_1397,N_640,N_972);
or U1398 (N_1398,N_618,N_711);
nor U1399 (N_1399,N_800,N_823);
and U1400 (N_1400,N_725,N_689);
nand U1401 (N_1401,N_716,N_962);
nor U1402 (N_1402,N_911,N_591);
or U1403 (N_1403,N_525,N_803);
nand U1404 (N_1404,N_656,N_881);
nand U1405 (N_1405,N_951,N_749);
or U1406 (N_1406,N_744,N_858);
nor U1407 (N_1407,N_733,N_672);
or U1408 (N_1408,N_965,N_833);
or U1409 (N_1409,N_987,N_957);
or U1410 (N_1410,N_667,N_642);
nor U1411 (N_1411,N_747,N_738);
xor U1412 (N_1412,N_529,N_970);
nand U1413 (N_1413,N_721,N_619);
or U1414 (N_1414,N_700,N_858);
or U1415 (N_1415,N_811,N_668);
nand U1416 (N_1416,N_617,N_726);
nor U1417 (N_1417,N_516,N_680);
nand U1418 (N_1418,N_968,N_841);
nand U1419 (N_1419,N_984,N_743);
or U1420 (N_1420,N_726,N_820);
nand U1421 (N_1421,N_590,N_539);
nand U1422 (N_1422,N_836,N_659);
nor U1423 (N_1423,N_870,N_536);
nor U1424 (N_1424,N_877,N_910);
or U1425 (N_1425,N_653,N_829);
nor U1426 (N_1426,N_548,N_528);
nand U1427 (N_1427,N_751,N_521);
nor U1428 (N_1428,N_945,N_663);
nor U1429 (N_1429,N_945,N_908);
or U1430 (N_1430,N_984,N_747);
and U1431 (N_1431,N_969,N_595);
xor U1432 (N_1432,N_944,N_615);
or U1433 (N_1433,N_904,N_733);
or U1434 (N_1434,N_568,N_685);
and U1435 (N_1435,N_635,N_993);
nand U1436 (N_1436,N_609,N_947);
and U1437 (N_1437,N_699,N_669);
or U1438 (N_1438,N_587,N_961);
nand U1439 (N_1439,N_731,N_733);
or U1440 (N_1440,N_633,N_934);
or U1441 (N_1441,N_693,N_541);
or U1442 (N_1442,N_978,N_664);
and U1443 (N_1443,N_758,N_809);
nand U1444 (N_1444,N_542,N_909);
and U1445 (N_1445,N_823,N_852);
and U1446 (N_1446,N_890,N_725);
xnor U1447 (N_1447,N_897,N_775);
and U1448 (N_1448,N_980,N_990);
nand U1449 (N_1449,N_732,N_915);
or U1450 (N_1450,N_906,N_888);
nand U1451 (N_1451,N_738,N_892);
or U1452 (N_1452,N_969,N_666);
nand U1453 (N_1453,N_614,N_573);
nor U1454 (N_1454,N_530,N_845);
xor U1455 (N_1455,N_683,N_675);
and U1456 (N_1456,N_917,N_783);
nor U1457 (N_1457,N_542,N_847);
nand U1458 (N_1458,N_799,N_881);
or U1459 (N_1459,N_686,N_919);
and U1460 (N_1460,N_623,N_909);
nand U1461 (N_1461,N_654,N_799);
nand U1462 (N_1462,N_800,N_511);
nor U1463 (N_1463,N_799,N_706);
or U1464 (N_1464,N_900,N_959);
and U1465 (N_1465,N_634,N_807);
nand U1466 (N_1466,N_520,N_827);
nor U1467 (N_1467,N_537,N_770);
nor U1468 (N_1468,N_840,N_648);
or U1469 (N_1469,N_947,N_781);
nand U1470 (N_1470,N_728,N_624);
and U1471 (N_1471,N_906,N_678);
nor U1472 (N_1472,N_712,N_554);
and U1473 (N_1473,N_615,N_873);
nor U1474 (N_1474,N_519,N_957);
nor U1475 (N_1475,N_855,N_732);
and U1476 (N_1476,N_514,N_509);
nand U1477 (N_1477,N_914,N_810);
or U1478 (N_1478,N_614,N_613);
nor U1479 (N_1479,N_948,N_739);
nand U1480 (N_1480,N_981,N_724);
nand U1481 (N_1481,N_848,N_537);
nor U1482 (N_1482,N_668,N_551);
and U1483 (N_1483,N_851,N_679);
nor U1484 (N_1484,N_952,N_672);
and U1485 (N_1485,N_656,N_511);
nor U1486 (N_1486,N_645,N_890);
and U1487 (N_1487,N_642,N_504);
nor U1488 (N_1488,N_847,N_705);
nor U1489 (N_1489,N_853,N_822);
nor U1490 (N_1490,N_501,N_857);
nor U1491 (N_1491,N_875,N_639);
and U1492 (N_1492,N_658,N_850);
and U1493 (N_1493,N_650,N_805);
and U1494 (N_1494,N_511,N_999);
or U1495 (N_1495,N_817,N_863);
or U1496 (N_1496,N_923,N_670);
or U1497 (N_1497,N_694,N_794);
nor U1498 (N_1498,N_875,N_627);
xnor U1499 (N_1499,N_971,N_819);
nand U1500 (N_1500,N_1427,N_1116);
nand U1501 (N_1501,N_1097,N_1246);
nand U1502 (N_1502,N_1403,N_1347);
and U1503 (N_1503,N_1496,N_1122);
and U1504 (N_1504,N_1060,N_1324);
and U1505 (N_1505,N_1467,N_1183);
nor U1506 (N_1506,N_1284,N_1181);
nor U1507 (N_1507,N_1411,N_1409);
and U1508 (N_1508,N_1092,N_1260);
xor U1509 (N_1509,N_1369,N_1441);
xnor U1510 (N_1510,N_1215,N_1152);
and U1511 (N_1511,N_1387,N_1451);
nor U1512 (N_1512,N_1459,N_1254);
and U1513 (N_1513,N_1013,N_1455);
nand U1514 (N_1514,N_1435,N_1279);
and U1515 (N_1515,N_1296,N_1188);
or U1516 (N_1516,N_1359,N_1253);
and U1517 (N_1517,N_1381,N_1492);
xnor U1518 (N_1518,N_1130,N_1065);
and U1519 (N_1519,N_1024,N_1317);
nand U1520 (N_1520,N_1225,N_1049);
or U1521 (N_1521,N_1154,N_1452);
and U1522 (N_1522,N_1098,N_1410);
or U1523 (N_1523,N_1119,N_1444);
nor U1524 (N_1524,N_1132,N_1101);
or U1525 (N_1525,N_1175,N_1153);
nand U1526 (N_1526,N_1430,N_1045);
nor U1527 (N_1527,N_1377,N_1449);
or U1528 (N_1528,N_1012,N_1137);
and U1529 (N_1529,N_1165,N_1257);
nand U1530 (N_1530,N_1345,N_1431);
xnor U1531 (N_1531,N_1035,N_1498);
and U1532 (N_1532,N_1242,N_1251);
nor U1533 (N_1533,N_1308,N_1182);
nand U1534 (N_1534,N_1143,N_1115);
nor U1535 (N_1535,N_1314,N_1147);
or U1536 (N_1536,N_1059,N_1159);
nor U1537 (N_1537,N_1234,N_1231);
or U1538 (N_1538,N_1198,N_1287);
nand U1539 (N_1539,N_1322,N_1004);
xnor U1540 (N_1540,N_1332,N_1155);
nor U1541 (N_1541,N_1385,N_1108);
or U1542 (N_1542,N_1388,N_1457);
or U1543 (N_1543,N_1080,N_1245);
nand U1544 (N_1544,N_1306,N_1187);
or U1545 (N_1545,N_1437,N_1463);
xnor U1546 (N_1546,N_1407,N_1432);
xnor U1547 (N_1547,N_1190,N_1267);
nand U1548 (N_1548,N_1297,N_1301);
nor U1549 (N_1549,N_1302,N_1408);
nand U1550 (N_1550,N_1447,N_1094);
nand U1551 (N_1551,N_1125,N_1037);
xnor U1552 (N_1552,N_1250,N_1391);
xnor U1553 (N_1553,N_1362,N_1400);
xor U1554 (N_1554,N_1394,N_1346);
nor U1555 (N_1555,N_1247,N_1028);
and U1556 (N_1556,N_1007,N_1095);
nor U1557 (N_1557,N_1390,N_1173);
and U1558 (N_1558,N_1236,N_1000);
xnor U1559 (N_1559,N_1376,N_1468);
and U1560 (N_1560,N_1353,N_1233);
and U1561 (N_1561,N_1490,N_1047);
nand U1562 (N_1562,N_1365,N_1050);
xor U1563 (N_1563,N_1210,N_1189);
xnor U1564 (N_1564,N_1494,N_1232);
xor U1565 (N_1565,N_1421,N_1099);
or U1566 (N_1566,N_1240,N_1171);
or U1567 (N_1567,N_1100,N_1052);
or U1568 (N_1568,N_1244,N_1022);
and U1569 (N_1569,N_1126,N_1285);
or U1570 (N_1570,N_1368,N_1396);
nand U1571 (N_1571,N_1361,N_1489);
xnor U1572 (N_1572,N_1383,N_1281);
nand U1573 (N_1573,N_1273,N_1061);
xnor U1574 (N_1574,N_1056,N_1062);
and U1575 (N_1575,N_1434,N_1337);
or U1576 (N_1576,N_1350,N_1406);
and U1577 (N_1577,N_1142,N_1033);
or U1578 (N_1578,N_1135,N_1224);
or U1579 (N_1579,N_1470,N_1200);
and U1580 (N_1580,N_1123,N_1323);
nand U1581 (N_1581,N_1292,N_1196);
nand U1582 (N_1582,N_1456,N_1386);
and U1583 (N_1583,N_1016,N_1029);
nor U1584 (N_1584,N_1229,N_1072);
nor U1585 (N_1585,N_1417,N_1472);
nor U1586 (N_1586,N_1248,N_1355);
and U1587 (N_1587,N_1474,N_1172);
nor U1588 (N_1588,N_1082,N_1473);
or U1589 (N_1589,N_1338,N_1063);
nor U1590 (N_1590,N_1151,N_1379);
or U1591 (N_1591,N_1136,N_1039);
and U1592 (N_1592,N_1331,N_1107);
nand U1593 (N_1593,N_1375,N_1429);
or U1594 (N_1594,N_1436,N_1483);
nand U1595 (N_1595,N_1318,N_1401);
nand U1596 (N_1596,N_1186,N_1184);
nand U1597 (N_1597,N_1077,N_1216);
nor U1598 (N_1598,N_1486,N_1048);
nor U1599 (N_1599,N_1488,N_1319);
or U1600 (N_1600,N_1040,N_1315);
nand U1601 (N_1601,N_1289,N_1178);
or U1602 (N_1602,N_1036,N_1360);
nand U1603 (N_1603,N_1144,N_1102);
or U1604 (N_1604,N_1085,N_1294);
nor U1605 (N_1605,N_1084,N_1027);
nand U1606 (N_1606,N_1433,N_1440);
and U1607 (N_1607,N_1237,N_1015);
and U1608 (N_1608,N_1316,N_1127);
and U1609 (N_1609,N_1073,N_1087);
xnor U1610 (N_1610,N_1380,N_1399);
and U1611 (N_1611,N_1480,N_1005);
nand U1612 (N_1612,N_1167,N_1482);
or U1613 (N_1613,N_1145,N_1255);
nor U1614 (N_1614,N_1259,N_1484);
xor U1615 (N_1615,N_1180,N_1169);
and U1616 (N_1616,N_1276,N_1348);
nor U1617 (N_1617,N_1081,N_1046);
nor U1618 (N_1618,N_1330,N_1031);
and U1619 (N_1619,N_1124,N_1105);
or U1620 (N_1620,N_1106,N_1032);
and U1621 (N_1621,N_1053,N_1193);
and U1622 (N_1622,N_1009,N_1358);
or U1623 (N_1623,N_1133,N_1389);
nor U1624 (N_1624,N_1371,N_1453);
nand U1625 (N_1625,N_1150,N_1382);
nand U1626 (N_1626,N_1208,N_1218);
nor U1627 (N_1627,N_1363,N_1228);
xnor U1628 (N_1628,N_1010,N_1089);
and U1629 (N_1629,N_1264,N_1286);
nor U1630 (N_1630,N_1272,N_1270);
and U1631 (N_1631,N_1282,N_1139);
nand U1632 (N_1632,N_1464,N_1177);
xor U1633 (N_1633,N_1034,N_1425);
xnor U1634 (N_1634,N_1422,N_1020);
and U1635 (N_1635,N_1161,N_1288);
and U1636 (N_1636,N_1026,N_1280);
nand U1637 (N_1637,N_1258,N_1131);
or U1638 (N_1638,N_1352,N_1088);
or U1639 (N_1639,N_1398,N_1068);
nor U1640 (N_1640,N_1491,N_1493);
and U1641 (N_1641,N_1460,N_1293);
nand U1642 (N_1642,N_1412,N_1327);
nor U1643 (N_1643,N_1156,N_1373);
xor U1644 (N_1644,N_1030,N_1235);
and U1645 (N_1645,N_1450,N_1148);
or U1646 (N_1646,N_1393,N_1214);
and U1647 (N_1647,N_1138,N_1220);
nand U1648 (N_1648,N_1207,N_1485);
or U1649 (N_1649,N_1415,N_1090);
nor U1650 (N_1650,N_1397,N_1356);
and U1651 (N_1651,N_1096,N_1149);
nor U1652 (N_1652,N_1023,N_1320);
or U1653 (N_1653,N_1203,N_1014);
nand U1654 (N_1654,N_1043,N_1075);
or U1655 (N_1655,N_1179,N_1185);
and U1656 (N_1656,N_1140,N_1176);
nor U1657 (N_1657,N_1295,N_1310);
nand U1658 (N_1658,N_1174,N_1249);
or U1659 (N_1659,N_1104,N_1219);
or U1660 (N_1660,N_1213,N_1299);
nor U1661 (N_1661,N_1458,N_1217);
nand U1662 (N_1662,N_1334,N_1262);
nand U1663 (N_1663,N_1162,N_1305);
nand U1664 (N_1664,N_1069,N_1274);
or U1665 (N_1665,N_1093,N_1277);
nor U1666 (N_1666,N_1495,N_1384);
and U1667 (N_1667,N_1357,N_1445);
or U1668 (N_1668,N_1311,N_1111);
or U1669 (N_1669,N_1477,N_1335);
nor U1670 (N_1670,N_1416,N_1168);
and U1671 (N_1671,N_1354,N_1476);
or U1672 (N_1672,N_1191,N_1443);
or U1673 (N_1673,N_1336,N_1160);
or U1674 (N_1674,N_1423,N_1146);
nand U1675 (N_1675,N_1304,N_1471);
xor U1676 (N_1676,N_1481,N_1438);
or U1677 (N_1677,N_1487,N_1011);
nor U1678 (N_1678,N_1239,N_1326);
and U1679 (N_1679,N_1309,N_1499);
or U1680 (N_1680,N_1117,N_1479);
nand U1681 (N_1681,N_1192,N_1018);
nor U1682 (N_1682,N_1298,N_1070);
nor U1683 (N_1683,N_1414,N_1238);
nor U1684 (N_1684,N_1266,N_1462);
or U1685 (N_1685,N_1428,N_1256);
nand U1686 (N_1686,N_1157,N_1340);
or U1687 (N_1687,N_1418,N_1426);
or U1688 (N_1688,N_1342,N_1103);
nand U1689 (N_1689,N_1121,N_1017);
nor U1690 (N_1690,N_1001,N_1392);
and U1691 (N_1691,N_1395,N_1170);
and U1692 (N_1692,N_1008,N_1067);
and U1693 (N_1693,N_1006,N_1497);
nor U1694 (N_1694,N_1263,N_1051);
or U1695 (N_1695,N_1404,N_1261);
and U1696 (N_1696,N_1372,N_1164);
nor U1697 (N_1697,N_1303,N_1044);
nand U1698 (N_1698,N_1118,N_1113);
or U1699 (N_1699,N_1064,N_1019);
and U1700 (N_1700,N_1448,N_1076);
and U1701 (N_1701,N_1413,N_1109);
nand U1702 (N_1702,N_1402,N_1041);
nand U1703 (N_1703,N_1405,N_1378);
nand U1704 (N_1704,N_1243,N_1025);
xor U1705 (N_1705,N_1110,N_1227);
or U1706 (N_1706,N_1209,N_1211);
and U1707 (N_1707,N_1078,N_1199);
and U1708 (N_1708,N_1283,N_1002);
nand U1709 (N_1709,N_1349,N_1204);
nand U1710 (N_1710,N_1275,N_1252);
nand U1711 (N_1711,N_1128,N_1112);
and U1712 (N_1712,N_1230,N_1313);
or U1713 (N_1713,N_1300,N_1222);
or U1714 (N_1714,N_1057,N_1158);
nand U1715 (N_1715,N_1439,N_1344);
or U1716 (N_1716,N_1091,N_1226);
nor U1717 (N_1717,N_1478,N_1333);
and U1718 (N_1718,N_1241,N_1291);
xor U1719 (N_1719,N_1454,N_1003);
or U1720 (N_1720,N_1466,N_1074);
nor U1721 (N_1721,N_1475,N_1021);
nand U1722 (N_1722,N_1329,N_1442);
or U1723 (N_1723,N_1079,N_1071);
and U1724 (N_1724,N_1205,N_1058);
or U1725 (N_1725,N_1163,N_1364);
or U1726 (N_1726,N_1202,N_1325);
nor U1727 (N_1727,N_1055,N_1461);
and U1728 (N_1728,N_1268,N_1201);
xnor U1729 (N_1729,N_1465,N_1351);
nand U1730 (N_1730,N_1206,N_1366);
nor U1731 (N_1731,N_1054,N_1278);
nand U1732 (N_1732,N_1194,N_1114);
nand U1733 (N_1733,N_1042,N_1419);
or U1734 (N_1734,N_1374,N_1038);
or U1735 (N_1735,N_1420,N_1424);
nand U1736 (N_1736,N_1328,N_1446);
nand U1737 (N_1737,N_1343,N_1370);
xnor U1738 (N_1738,N_1120,N_1312);
nand U1739 (N_1739,N_1341,N_1221);
nand U1740 (N_1740,N_1339,N_1134);
nor U1741 (N_1741,N_1321,N_1195);
and U1742 (N_1742,N_1307,N_1367);
nand U1743 (N_1743,N_1066,N_1469);
nand U1744 (N_1744,N_1166,N_1086);
nand U1745 (N_1745,N_1271,N_1223);
and U1746 (N_1746,N_1265,N_1141);
nor U1747 (N_1747,N_1269,N_1083);
nand U1748 (N_1748,N_1197,N_1129);
nor U1749 (N_1749,N_1290,N_1212);
nor U1750 (N_1750,N_1347,N_1011);
and U1751 (N_1751,N_1140,N_1051);
xor U1752 (N_1752,N_1181,N_1170);
xor U1753 (N_1753,N_1034,N_1322);
or U1754 (N_1754,N_1215,N_1236);
nor U1755 (N_1755,N_1322,N_1491);
nand U1756 (N_1756,N_1006,N_1121);
nand U1757 (N_1757,N_1090,N_1307);
nor U1758 (N_1758,N_1241,N_1268);
and U1759 (N_1759,N_1168,N_1159);
or U1760 (N_1760,N_1116,N_1310);
nand U1761 (N_1761,N_1465,N_1291);
or U1762 (N_1762,N_1481,N_1346);
nor U1763 (N_1763,N_1334,N_1217);
and U1764 (N_1764,N_1059,N_1491);
nand U1765 (N_1765,N_1017,N_1348);
nand U1766 (N_1766,N_1238,N_1003);
or U1767 (N_1767,N_1106,N_1224);
nand U1768 (N_1768,N_1346,N_1366);
and U1769 (N_1769,N_1009,N_1319);
or U1770 (N_1770,N_1259,N_1395);
and U1771 (N_1771,N_1161,N_1431);
or U1772 (N_1772,N_1111,N_1194);
xor U1773 (N_1773,N_1078,N_1306);
and U1774 (N_1774,N_1495,N_1346);
nor U1775 (N_1775,N_1223,N_1067);
or U1776 (N_1776,N_1036,N_1286);
nor U1777 (N_1777,N_1158,N_1428);
nand U1778 (N_1778,N_1017,N_1176);
or U1779 (N_1779,N_1175,N_1179);
nor U1780 (N_1780,N_1320,N_1376);
nand U1781 (N_1781,N_1095,N_1338);
or U1782 (N_1782,N_1472,N_1312);
or U1783 (N_1783,N_1455,N_1111);
and U1784 (N_1784,N_1307,N_1408);
nor U1785 (N_1785,N_1007,N_1011);
and U1786 (N_1786,N_1259,N_1285);
nand U1787 (N_1787,N_1408,N_1187);
nor U1788 (N_1788,N_1101,N_1011);
nor U1789 (N_1789,N_1194,N_1166);
nor U1790 (N_1790,N_1219,N_1000);
nor U1791 (N_1791,N_1458,N_1349);
or U1792 (N_1792,N_1248,N_1282);
or U1793 (N_1793,N_1028,N_1172);
or U1794 (N_1794,N_1076,N_1442);
or U1795 (N_1795,N_1477,N_1365);
nand U1796 (N_1796,N_1463,N_1116);
or U1797 (N_1797,N_1460,N_1318);
or U1798 (N_1798,N_1361,N_1177);
nor U1799 (N_1799,N_1078,N_1396);
and U1800 (N_1800,N_1221,N_1430);
nor U1801 (N_1801,N_1335,N_1223);
nand U1802 (N_1802,N_1250,N_1068);
nand U1803 (N_1803,N_1129,N_1167);
nor U1804 (N_1804,N_1031,N_1006);
nor U1805 (N_1805,N_1334,N_1291);
nor U1806 (N_1806,N_1221,N_1178);
and U1807 (N_1807,N_1228,N_1018);
nand U1808 (N_1808,N_1242,N_1356);
nor U1809 (N_1809,N_1156,N_1307);
nor U1810 (N_1810,N_1240,N_1043);
and U1811 (N_1811,N_1287,N_1286);
nand U1812 (N_1812,N_1160,N_1462);
and U1813 (N_1813,N_1487,N_1257);
and U1814 (N_1814,N_1152,N_1079);
nand U1815 (N_1815,N_1196,N_1347);
nand U1816 (N_1816,N_1229,N_1164);
xor U1817 (N_1817,N_1063,N_1227);
nor U1818 (N_1818,N_1142,N_1392);
nand U1819 (N_1819,N_1244,N_1069);
xor U1820 (N_1820,N_1295,N_1202);
nand U1821 (N_1821,N_1080,N_1445);
xnor U1822 (N_1822,N_1359,N_1176);
nand U1823 (N_1823,N_1359,N_1420);
or U1824 (N_1824,N_1276,N_1177);
nor U1825 (N_1825,N_1423,N_1227);
and U1826 (N_1826,N_1434,N_1308);
nand U1827 (N_1827,N_1190,N_1323);
and U1828 (N_1828,N_1078,N_1280);
nor U1829 (N_1829,N_1419,N_1018);
and U1830 (N_1830,N_1275,N_1316);
nor U1831 (N_1831,N_1035,N_1061);
nor U1832 (N_1832,N_1298,N_1149);
nand U1833 (N_1833,N_1444,N_1363);
nand U1834 (N_1834,N_1222,N_1206);
nand U1835 (N_1835,N_1095,N_1468);
nor U1836 (N_1836,N_1096,N_1249);
nand U1837 (N_1837,N_1482,N_1453);
nand U1838 (N_1838,N_1315,N_1160);
nand U1839 (N_1839,N_1472,N_1272);
or U1840 (N_1840,N_1228,N_1061);
xnor U1841 (N_1841,N_1377,N_1224);
or U1842 (N_1842,N_1174,N_1231);
nor U1843 (N_1843,N_1153,N_1381);
nand U1844 (N_1844,N_1439,N_1094);
and U1845 (N_1845,N_1011,N_1314);
nand U1846 (N_1846,N_1417,N_1038);
xnor U1847 (N_1847,N_1159,N_1043);
nand U1848 (N_1848,N_1351,N_1362);
nand U1849 (N_1849,N_1273,N_1306);
and U1850 (N_1850,N_1337,N_1010);
nand U1851 (N_1851,N_1358,N_1459);
and U1852 (N_1852,N_1191,N_1148);
or U1853 (N_1853,N_1298,N_1297);
nor U1854 (N_1854,N_1431,N_1478);
nor U1855 (N_1855,N_1379,N_1143);
or U1856 (N_1856,N_1225,N_1150);
nand U1857 (N_1857,N_1327,N_1244);
nand U1858 (N_1858,N_1474,N_1351);
and U1859 (N_1859,N_1151,N_1083);
nand U1860 (N_1860,N_1463,N_1400);
and U1861 (N_1861,N_1031,N_1097);
nand U1862 (N_1862,N_1224,N_1128);
nor U1863 (N_1863,N_1124,N_1201);
nor U1864 (N_1864,N_1188,N_1425);
nand U1865 (N_1865,N_1329,N_1357);
nor U1866 (N_1866,N_1443,N_1106);
and U1867 (N_1867,N_1038,N_1267);
or U1868 (N_1868,N_1219,N_1440);
nor U1869 (N_1869,N_1285,N_1391);
nor U1870 (N_1870,N_1386,N_1139);
or U1871 (N_1871,N_1484,N_1319);
nand U1872 (N_1872,N_1460,N_1301);
nor U1873 (N_1873,N_1345,N_1075);
nand U1874 (N_1874,N_1188,N_1244);
nand U1875 (N_1875,N_1359,N_1427);
nor U1876 (N_1876,N_1286,N_1260);
and U1877 (N_1877,N_1110,N_1470);
nor U1878 (N_1878,N_1071,N_1082);
xnor U1879 (N_1879,N_1018,N_1467);
or U1880 (N_1880,N_1206,N_1476);
or U1881 (N_1881,N_1285,N_1015);
or U1882 (N_1882,N_1301,N_1212);
nor U1883 (N_1883,N_1188,N_1414);
nand U1884 (N_1884,N_1325,N_1300);
xor U1885 (N_1885,N_1180,N_1159);
xor U1886 (N_1886,N_1266,N_1205);
xor U1887 (N_1887,N_1277,N_1279);
and U1888 (N_1888,N_1006,N_1159);
nand U1889 (N_1889,N_1428,N_1461);
nand U1890 (N_1890,N_1375,N_1196);
nand U1891 (N_1891,N_1356,N_1366);
and U1892 (N_1892,N_1282,N_1402);
xnor U1893 (N_1893,N_1304,N_1436);
nand U1894 (N_1894,N_1323,N_1022);
nand U1895 (N_1895,N_1140,N_1195);
or U1896 (N_1896,N_1078,N_1053);
nor U1897 (N_1897,N_1403,N_1208);
xor U1898 (N_1898,N_1270,N_1369);
nand U1899 (N_1899,N_1364,N_1456);
nand U1900 (N_1900,N_1393,N_1375);
nand U1901 (N_1901,N_1129,N_1420);
nor U1902 (N_1902,N_1048,N_1205);
nand U1903 (N_1903,N_1137,N_1154);
or U1904 (N_1904,N_1163,N_1231);
and U1905 (N_1905,N_1464,N_1293);
and U1906 (N_1906,N_1359,N_1221);
and U1907 (N_1907,N_1284,N_1003);
xor U1908 (N_1908,N_1124,N_1065);
and U1909 (N_1909,N_1038,N_1482);
xnor U1910 (N_1910,N_1416,N_1441);
or U1911 (N_1911,N_1465,N_1339);
or U1912 (N_1912,N_1029,N_1225);
xnor U1913 (N_1913,N_1062,N_1349);
xor U1914 (N_1914,N_1237,N_1202);
nor U1915 (N_1915,N_1059,N_1022);
nand U1916 (N_1916,N_1436,N_1264);
or U1917 (N_1917,N_1461,N_1423);
xor U1918 (N_1918,N_1133,N_1205);
nor U1919 (N_1919,N_1424,N_1146);
xor U1920 (N_1920,N_1408,N_1105);
nor U1921 (N_1921,N_1499,N_1361);
nor U1922 (N_1922,N_1015,N_1051);
nand U1923 (N_1923,N_1486,N_1090);
xor U1924 (N_1924,N_1053,N_1013);
nor U1925 (N_1925,N_1072,N_1064);
xor U1926 (N_1926,N_1311,N_1124);
nand U1927 (N_1927,N_1072,N_1154);
or U1928 (N_1928,N_1342,N_1184);
nand U1929 (N_1929,N_1234,N_1367);
or U1930 (N_1930,N_1118,N_1447);
nand U1931 (N_1931,N_1445,N_1040);
xnor U1932 (N_1932,N_1478,N_1207);
and U1933 (N_1933,N_1133,N_1019);
or U1934 (N_1934,N_1019,N_1283);
or U1935 (N_1935,N_1382,N_1292);
nor U1936 (N_1936,N_1238,N_1482);
or U1937 (N_1937,N_1431,N_1341);
nor U1938 (N_1938,N_1137,N_1445);
or U1939 (N_1939,N_1299,N_1441);
nand U1940 (N_1940,N_1097,N_1242);
nor U1941 (N_1941,N_1375,N_1268);
or U1942 (N_1942,N_1031,N_1073);
or U1943 (N_1943,N_1264,N_1406);
nor U1944 (N_1944,N_1392,N_1486);
nand U1945 (N_1945,N_1373,N_1334);
or U1946 (N_1946,N_1270,N_1257);
nand U1947 (N_1947,N_1465,N_1490);
and U1948 (N_1948,N_1011,N_1133);
xnor U1949 (N_1949,N_1212,N_1015);
nor U1950 (N_1950,N_1432,N_1015);
or U1951 (N_1951,N_1290,N_1260);
nor U1952 (N_1952,N_1391,N_1261);
nand U1953 (N_1953,N_1205,N_1300);
nor U1954 (N_1954,N_1407,N_1393);
and U1955 (N_1955,N_1352,N_1417);
or U1956 (N_1956,N_1296,N_1170);
or U1957 (N_1957,N_1142,N_1280);
and U1958 (N_1958,N_1181,N_1291);
nor U1959 (N_1959,N_1277,N_1220);
nor U1960 (N_1960,N_1098,N_1376);
nand U1961 (N_1961,N_1094,N_1175);
and U1962 (N_1962,N_1393,N_1370);
nor U1963 (N_1963,N_1088,N_1196);
nand U1964 (N_1964,N_1166,N_1491);
nand U1965 (N_1965,N_1380,N_1403);
nand U1966 (N_1966,N_1117,N_1008);
or U1967 (N_1967,N_1113,N_1316);
nand U1968 (N_1968,N_1274,N_1266);
and U1969 (N_1969,N_1022,N_1122);
or U1970 (N_1970,N_1301,N_1302);
nor U1971 (N_1971,N_1113,N_1451);
nor U1972 (N_1972,N_1022,N_1458);
or U1973 (N_1973,N_1301,N_1328);
or U1974 (N_1974,N_1442,N_1041);
nand U1975 (N_1975,N_1411,N_1137);
or U1976 (N_1976,N_1009,N_1067);
and U1977 (N_1977,N_1226,N_1247);
or U1978 (N_1978,N_1241,N_1380);
and U1979 (N_1979,N_1474,N_1234);
or U1980 (N_1980,N_1361,N_1396);
or U1981 (N_1981,N_1344,N_1320);
nor U1982 (N_1982,N_1020,N_1116);
and U1983 (N_1983,N_1460,N_1187);
nor U1984 (N_1984,N_1248,N_1181);
or U1985 (N_1985,N_1379,N_1287);
nor U1986 (N_1986,N_1169,N_1287);
nand U1987 (N_1987,N_1288,N_1106);
or U1988 (N_1988,N_1187,N_1107);
and U1989 (N_1989,N_1482,N_1485);
nor U1990 (N_1990,N_1185,N_1207);
nor U1991 (N_1991,N_1013,N_1293);
and U1992 (N_1992,N_1370,N_1284);
nor U1993 (N_1993,N_1373,N_1223);
nor U1994 (N_1994,N_1082,N_1115);
and U1995 (N_1995,N_1449,N_1152);
or U1996 (N_1996,N_1067,N_1494);
nor U1997 (N_1997,N_1047,N_1308);
or U1998 (N_1998,N_1237,N_1033);
nor U1999 (N_1999,N_1365,N_1229);
nand U2000 (N_2000,N_1527,N_1624);
or U2001 (N_2001,N_1875,N_1569);
nand U2002 (N_2002,N_1966,N_1621);
xnor U2003 (N_2003,N_1656,N_1899);
nor U2004 (N_2004,N_1914,N_1629);
nor U2005 (N_2005,N_1730,N_1913);
or U2006 (N_2006,N_1865,N_1771);
nand U2007 (N_2007,N_1874,N_1995);
nor U2008 (N_2008,N_1711,N_1563);
nand U2009 (N_2009,N_1727,N_1681);
xor U2010 (N_2010,N_1941,N_1674);
and U2011 (N_2011,N_1637,N_1816);
nor U2012 (N_2012,N_1792,N_1873);
nor U2013 (N_2013,N_1587,N_1748);
and U2014 (N_2014,N_1779,N_1616);
nor U2015 (N_2015,N_1612,N_1581);
or U2016 (N_2016,N_1946,N_1660);
or U2017 (N_2017,N_1859,N_1920);
or U2018 (N_2018,N_1867,N_1952);
nand U2019 (N_2019,N_1757,N_1762);
and U2020 (N_2020,N_1718,N_1615);
or U2021 (N_2021,N_1922,N_1566);
nand U2022 (N_2022,N_1672,N_1526);
nand U2023 (N_2023,N_1697,N_1901);
nand U2024 (N_2024,N_1758,N_1579);
nand U2025 (N_2025,N_1554,N_1676);
nor U2026 (N_2026,N_1880,N_1667);
and U2027 (N_2027,N_1845,N_1775);
nand U2028 (N_2028,N_1801,N_1693);
or U2029 (N_2029,N_1850,N_1887);
and U2030 (N_2030,N_1954,N_1720);
nand U2031 (N_2031,N_1906,N_1971);
and U2032 (N_2032,N_1630,N_1878);
and U2033 (N_2033,N_1766,N_1543);
and U2034 (N_2034,N_1652,N_1739);
nand U2035 (N_2035,N_1896,N_1552);
nand U2036 (N_2036,N_1602,N_1596);
and U2037 (N_2037,N_1951,N_1796);
or U2038 (N_2038,N_1839,N_1823);
and U2039 (N_2039,N_1789,N_1717);
nand U2040 (N_2040,N_1950,N_1933);
or U2041 (N_2041,N_1538,N_1648);
nand U2042 (N_2042,N_1734,N_1871);
nand U2043 (N_2043,N_1562,N_1611);
or U2044 (N_2044,N_1726,N_1858);
nand U2045 (N_2045,N_1740,N_1813);
and U2046 (N_2046,N_1561,N_1908);
or U2047 (N_2047,N_1668,N_1780);
and U2048 (N_2048,N_1550,N_1575);
or U2049 (N_2049,N_1683,N_1515);
nand U2050 (N_2050,N_1774,N_1591);
nor U2051 (N_2051,N_1653,N_1974);
and U2052 (N_2052,N_1745,N_1544);
nand U2053 (N_2053,N_1754,N_1853);
nand U2054 (N_2054,N_1905,N_1626);
or U2055 (N_2055,N_1585,N_1699);
nand U2056 (N_2056,N_1628,N_1953);
nor U2057 (N_2057,N_1959,N_1751);
and U2058 (N_2058,N_1589,N_1650);
or U2059 (N_2059,N_1507,N_1891);
nor U2060 (N_2060,N_1576,N_1996);
and U2061 (N_2061,N_1753,N_1578);
nor U2062 (N_2062,N_1925,N_1688);
nand U2063 (N_2063,N_1862,N_1743);
xor U2064 (N_2064,N_1814,N_1930);
or U2065 (N_2065,N_1980,N_1512);
nor U2066 (N_2066,N_1738,N_1705);
xnor U2067 (N_2067,N_1655,N_1898);
and U2068 (N_2068,N_1509,N_1877);
and U2069 (N_2069,N_1881,N_1784);
nand U2070 (N_2070,N_1694,N_1866);
and U2071 (N_2071,N_1894,N_1572);
nand U2072 (N_2072,N_1541,N_1943);
nor U2073 (N_2073,N_1764,N_1564);
or U2074 (N_2074,N_1610,N_1776);
or U2075 (N_2075,N_1768,N_1787);
xor U2076 (N_2076,N_1640,N_1670);
xnor U2077 (N_2077,N_1909,N_1742);
or U2078 (N_2078,N_1545,N_1584);
and U2079 (N_2079,N_1686,N_1879);
or U2080 (N_2080,N_1810,N_1707);
or U2081 (N_2081,N_1645,N_1781);
nor U2082 (N_2082,N_1857,N_1567);
nor U2083 (N_2083,N_1647,N_1838);
or U2084 (N_2084,N_1919,N_1613);
nor U2085 (N_2085,N_1662,N_1828);
and U2086 (N_2086,N_1945,N_1836);
nor U2087 (N_2087,N_1514,N_1590);
nor U2088 (N_2088,N_1593,N_1799);
nand U2089 (N_2089,N_1932,N_1682);
and U2090 (N_2090,N_1967,N_1884);
or U2091 (N_2091,N_1956,N_1605);
nand U2092 (N_2092,N_1599,N_1638);
or U2093 (N_2093,N_1634,N_1529);
or U2094 (N_2094,N_1820,N_1982);
nand U2095 (N_2095,N_1876,N_1825);
nand U2096 (N_2096,N_1870,N_1657);
and U2097 (N_2097,N_1993,N_1635);
xor U2098 (N_2098,N_1687,N_1869);
nor U2099 (N_2099,N_1724,N_1888);
nor U2100 (N_2100,N_1972,N_1614);
nand U2101 (N_2101,N_1903,N_1573);
nand U2102 (N_2102,N_1643,N_1934);
or U2103 (N_2103,N_1746,N_1520);
nand U2104 (N_2104,N_1555,N_1918);
and U2105 (N_2105,N_1793,N_1513);
nand U2106 (N_2106,N_1700,N_1607);
or U2107 (N_2107,N_1936,N_1958);
or U2108 (N_2108,N_1617,N_1533);
and U2109 (N_2109,N_1570,N_1594);
nor U2110 (N_2110,N_1651,N_1604);
nand U2111 (N_2111,N_1856,N_1991);
or U2112 (N_2112,N_1846,N_1890);
nand U2113 (N_2113,N_1981,N_1633);
nand U2114 (N_2114,N_1709,N_1534);
and U2115 (N_2115,N_1665,N_1802);
and U2116 (N_2116,N_1760,N_1818);
or U2117 (N_2117,N_1791,N_1864);
and U2118 (N_2118,N_1518,N_1904);
or U2119 (N_2119,N_1510,N_1749);
xor U2120 (N_2120,N_1938,N_1990);
nor U2121 (N_2121,N_1553,N_1924);
nor U2122 (N_2122,N_1897,N_1580);
or U2123 (N_2123,N_1639,N_1755);
xnor U2124 (N_2124,N_1900,N_1808);
and U2125 (N_2125,N_1636,N_1644);
and U2126 (N_2126,N_1911,N_1883);
nor U2127 (N_2127,N_1809,N_1855);
xor U2128 (N_2128,N_1673,N_1677);
or U2129 (N_2129,N_1765,N_1654);
nand U2130 (N_2130,N_1842,N_1916);
and U2131 (N_2131,N_1931,N_1992);
or U2132 (N_2132,N_1912,N_1804);
or U2133 (N_2133,N_1763,N_1568);
nor U2134 (N_2134,N_1747,N_1817);
nor U2135 (N_2135,N_1500,N_1935);
xnor U2136 (N_2136,N_1803,N_1625);
or U2137 (N_2137,N_1915,N_1968);
nand U2138 (N_2138,N_1664,N_1829);
nor U2139 (N_2139,N_1606,N_1841);
xnor U2140 (N_2140,N_1537,N_1986);
and U2141 (N_2141,N_1558,N_1790);
or U2142 (N_2142,N_1861,N_1752);
nor U2143 (N_2143,N_1511,N_1895);
nand U2144 (N_2144,N_1595,N_1600);
and U2145 (N_2145,N_1821,N_1522);
and U2146 (N_2146,N_1704,N_1994);
and U2147 (N_2147,N_1960,N_1588);
nand U2148 (N_2148,N_1977,N_1947);
xnor U2149 (N_2149,N_1530,N_1549);
nor U2150 (N_2150,N_1840,N_1517);
xor U2151 (N_2151,N_1571,N_1937);
nand U2152 (N_2152,N_1706,N_1532);
and U2153 (N_2153,N_1770,N_1921);
and U2154 (N_2154,N_1631,N_1548);
nand U2155 (N_2155,N_1948,N_1975);
nand U2156 (N_2156,N_1502,N_1761);
or U2157 (N_2157,N_1723,N_1939);
or U2158 (N_2158,N_1698,N_1988);
or U2159 (N_2159,N_1843,N_1715);
or U2160 (N_2160,N_1557,N_1852);
nor U2161 (N_2161,N_1811,N_1623);
and U2162 (N_2162,N_1849,N_1831);
nor U2163 (N_2163,N_1744,N_1620);
nand U2164 (N_2164,N_1642,N_1539);
nor U2165 (N_2165,N_1927,N_1970);
nand U2166 (N_2166,N_1999,N_1547);
nor U2167 (N_2167,N_1834,N_1710);
and U2168 (N_2168,N_1978,N_1926);
xnor U2169 (N_2169,N_1832,N_1504);
and U2170 (N_2170,N_1756,N_1783);
xnor U2171 (N_2171,N_1506,N_1782);
nand U2172 (N_2172,N_1528,N_1603);
and U2173 (N_2173,N_1684,N_1955);
and U2174 (N_2174,N_1679,N_1666);
nand U2175 (N_2175,N_1680,N_1508);
or U2176 (N_2176,N_1728,N_1722);
nor U2177 (N_2177,N_1767,N_1619);
xor U2178 (N_2178,N_1979,N_1860);
nor U2179 (N_2179,N_1586,N_1826);
nand U2180 (N_2180,N_1902,N_1797);
and U2181 (N_2181,N_1805,N_1523);
nor U2182 (N_2182,N_1659,N_1708);
and U2183 (N_2183,N_1917,N_1985);
or U2184 (N_2184,N_1889,N_1516);
and U2185 (N_2185,N_1886,N_1872);
nor U2186 (N_2186,N_1702,N_1844);
and U2187 (N_2187,N_1721,N_1536);
and U2188 (N_2188,N_1940,N_1689);
or U2189 (N_2189,N_1663,N_1546);
or U2190 (N_2190,N_1851,N_1713);
xnor U2191 (N_2191,N_1863,N_1559);
xor U2192 (N_2192,N_1929,N_1519);
nor U2193 (N_2193,N_1695,N_1618);
or U2194 (N_2194,N_1551,N_1535);
xnor U2195 (N_2195,N_1854,N_1669);
and U2196 (N_2196,N_1737,N_1983);
xor U2197 (N_2197,N_1691,N_1592);
nor U2198 (N_2198,N_1701,N_1641);
nand U2199 (N_2199,N_1984,N_1964);
nor U2200 (N_2200,N_1798,N_1907);
nor U2201 (N_2201,N_1976,N_1729);
nor U2202 (N_2202,N_1969,N_1703);
and U2203 (N_2203,N_1815,N_1735);
xnor U2204 (N_2204,N_1827,N_1957);
nor U2205 (N_2205,N_1675,N_1524);
xor U2206 (N_2206,N_1788,N_1690);
nor U2207 (N_2207,N_1685,N_1778);
or U2208 (N_2208,N_1893,N_1949);
xnor U2209 (N_2209,N_1733,N_1795);
or U2210 (N_2210,N_1830,N_1608);
and U2211 (N_2211,N_1998,N_1732);
or U2212 (N_2212,N_1773,N_1646);
or U2213 (N_2213,N_1824,N_1963);
nand U2214 (N_2214,N_1501,N_1598);
nand U2215 (N_2215,N_1583,N_1785);
and U2216 (N_2216,N_1885,N_1714);
xnor U2217 (N_2217,N_1772,N_1609);
or U2218 (N_2218,N_1835,N_1819);
nor U2219 (N_2219,N_1601,N_1868);
nor U2220 (N_2220,N_1961,N_1627);
and U2221 (N_2221,N_1622,N_1928);
and U2222 (N_2222,N_1837,N_1741);
xor U2223 (N_2223,N_1692,N_1987);
and U2224 (N_2224,N_1800,N_1989);
nor U2225 (N_2225,N_1719,N_1597);
xnor U2226 (N_2226,N_1574,N_1736);
or U2227 (N_2227,N_1503,N_1521);
xnor U2228 (N_2228,N_1716,N_1794);
and U2229 (N_2229,N_1833,N_1525);
and U2230 (N_2230,N_1965,N_1556);
or U2231 (N_2231,N_1696,N_1786);
or U2232 (N_2232,N_1658,N_1807);
or U2233 (N_2233,N_1632,N_1531);
nand U2234 (N_2234,N_1582,N_1560);
nand U2235 (N_2235,N_1910,N_1540);
nor U2236 (N_2236,N_1577,N_1882);
or U2237 (N_2237,N_1769,N_1973);
and U2238 (N_2238,N_1712,N_1671);
xor U2239 (N_2239,N_1731,N_1923);
or U2240 (N_2240,N_1962,N_1806);
or U2241 (N_2241,N_1759,N_1725);
xnor U2242 (N_2242,N_1997,N_1848);
nor U2243 (N_2243,N_1565,N_1678);
or U2244 (N_2244,N_1944,N_1505);
xor U2245 (N_2245,N_1892,N_1542);
nand U2246 (N_2246,N_1812,N_1942);
xnor U2247 (N_2247,N_1750,N_1777);
nor U2248 (N_2248,N_1822,N_1661);
or U2249 (N_2249,N_1847,N_1649);
xnor U2250 (N_2250,N_1912,N_1578);
or U2251 (N_2251,N_1878,N_1974);
or U2252 (N_2252,N_1663,N_1728);
or U2253 (N_2253,N_1733,N_1573);
and U2254 (N_2254,N_1816,N_1590);
and U2255 (N_2255,N_1620,N_1661);
and U2256 (N_2256,N_1865,N_1718);
nand U2257 (N_2257,N_1909,N_1500);
nor U2258 (N_2258,N_1916,N_1775);
nand U2259 (N_2259,N_1804,N_1806);
nor U2260 (N_2260,N_1593,N_1548);
or U2261 (N_2261,N_1762,N_1954);
xnor U2262 (N_2262,N_1888,N_1603);
or U2263 (N_2263,N_1673,N_1841);
nand U2264 (N_2264,N_1541,N_1864);
and U2265 (N_2265,N_1660,N_1715);
and U2266 (N_2266,N_1655,N_1555);
nor U2267 (N_2267,N_1831,N_1802);
nor U2268 (N_2268,N_1621,N_1632);
or U2269 (N_2269,N_1818,N_1805);
and U2270 (N_2270,N_1679,N_1857);
or U2271 (N_2271,N_1741,N_1986);
nor U2272 (N_2272,N_1890,N_1771);
or U2273 (N_2273,N_1836,N_1535);
or U2274 (N_2274,N_1607,N_1660);
nor U2275 (N_2275,N_1934,N_1835);
or U2276 (N_2276,N_1969,N_1647);
and U2277 (N_2277,N_1713,N_1575);
and U2278 (N_2278,N_1829,N_1966);
nor U2279 (N_2279,N_1962,N_1625);
or U2280 (N_2280,N_1665,N_1725);
nor U2281 (N_2281,N_1746,N_1587);
and U2282 (N_2282,N_1789,N_1749);
or U2283 (N_2283,N_1900,N_1994);
nor U2284 (N_2284,N_1783,N_1517);
nor U2285 (N_2285,N_1625,N_1864);
or U2286 (N_2286,N_1535,N_1743);
or U2287 (N_2287,N_1604,N_1996);
nand U2288 (N_2288,N_1577,N_1768);
and U2289 (N_2289,N_1588,N_1561);
nand U2290 (N_2290,N_1946,N_1929);
and U2291 (N_2291,N_1718,N_1776);
or U2292 (N_2292,N_1880,N_1547);
and U2293 (N_2293,N_1796,N_1761);
xor U2294 (N_2294,N_1641,N_1989);
nand U2295 (N_2295,N_1899,N_1959);
nor U2296 (N_2296,N_1640,N_1901);
and U2297 (N_2297,N_1721,N_1843);
nor U2298 (N_2298,N_1625,N_1563);
nand U2299 (N_2299,N_1857,N_1569);
nor U2300 (N_2300,N_1901,N_1906);
nand U2301 (N_2301,N_1757,N_1634);
xor U2302 (N_2302,N_1973,N_1685);
nand U2303 (N_2303,N_1659,N_1809);
nand U2304 (N_2304,N_1847,N_1838);
nor U2305 (N_2305,N_1552,N_1649);
nor U2306 (N_2306,N_1812,N_1749);
or U2307 (N_2307,N_1511,N_1640);
nand U2308 (N_2308,N_1893,N_1969);
or U2309 (N_2309,N_1845,N_1569);
nand U2310 (N_2310,N_1842,N_1972);
xor U2311 (N_2311,N_1728,N_1787);
nand U2312 (N_2312,N_1598,N_1804);
and U2313 (N_2313,N_1994,N_1764);
and U2314 (N_2314,N_1673,N_1500);
nand U2315 (N_2315,N_1575,N_1507);
nor U2316 (N_2316,N_1956,N_1501);
and U2317 (N_2317,N_1612,N_1828);
or U2318 (N_2318,N_1877,N_1783);
nor U2319 (N_2319,N_1665,N_1767);
and U2320 (N_2320,N_1572,N_1680);
nor U2321 (N_2321,N_1752,N_1528);
or U2322 (N_2322,N_1728,N_1769);
nand U2323 (N_2323,N_1949,N_1897);
or U2324 (N_2324,N_1684,N_1775);
or U2325 (N_2325,N_1904,N_1627);
or U2326 (N_2326,N_1616,N_1900);
nand U2327 (N_2327,N_1646,N_1655);
and U2328 (N_2328,N_1504,N_1547);
nand U2329 (N_2329,N_1896,N_1887);
or U2330 (N_2330,N_1778,N_1934);
or U2331 (N_2331,N_1607,N_1545);
nor U2332 (N_2332,N_1614,N_1558);
nor U2333 (N_2333,N_1793,N_1921);
and U2334 (N_2334,N_1683,N_1997);
and U2335 (N_2335,N_1877,N_1736);
nor U2336 (N_2336,N_1984,N_1612);
nand U2337 (N_2337,N_1928,N_1716);
or U2338 (N_2338,N_1621,N_1637);
and U2339 (N_2339,N_1703,N_1578);
and U2340 (N_2340,N_1791,N_1660);
and U2341 (N_2341,N_1856,N_1788);
nor U2342 (N_2342,N_1603,N_1670);
nor U2343 (N_2343,N_1842,N_1852);
nand U2344 (N_2344,N_1693,N_1969);
and U2345 (N_2345,N_1875,N_1632);
and U2346 (N_2346,N_1520,N_1551);
and U2347 (N_2347,N_1799,N_1821);
or U2348 (N_2348,N_1974,N_1909);
or U2349 (N_2349,N_1950,N_1576);
or U2350 (N_2350,N_1901,N_1503);
or U2351 (N_2351,N_1757,N_1571);
and U2352 (N_2352,N_1542,N_1506);
or U2353 (N_2353,N_1682,N_1964);
xor U2354 (N_2354,N_1730,N_1898);
nor U2355 (N_2355,N_1572,N_1863);
nand U2356 (N_2356,N_1978,N_1621);
nand U2357 (N_2357,N_1623,N_1793);
xnor U2358 (N_2358,N_1550,N_1897);
nand U2359 (N_2359,N_1706,N_1955);
nor U2360 (N_2360,N_1761,N_1565);
and U2361 (N_2361,N_1943,N_1921);
or U2362 (N_2362,N_1663,N_1628);
xnor U2363 (N_2363,N_1636,N_1818);
or U2364 (N_2364,N_1813,N_1869);
nor U2365 (N_2365,N_1770,N_1734);
and U2366 (N_2366,N_1857,N_1600);
or U2367 (N_2367,N_1804,N_1557);
and U2368 (N_2368,N_1863,N_1685);
or U2369 (N_2369,N_1702,N_1676);
and U2370 (N_2370,N_1744,N_1951);
and U2371 (N_2371,N_1838,N_1644);
or U2372 (N_2372,N_1666,N_1619);
nor U2373 (N_2373,N_1514,N_1696);
and U2374 (N_2374,N_1714,N_1906);
or U2375 (N_2375,N_1956,N_1898);
xnor U2376 (N_2376,N_1648,N_1630);
and U2377 (N_2377,N_1872,N_1673);
or U2378 (N_2378,N_1780,N_1757);
nand U2379 (N_2379,N_1754,N_1959);
or U2380 (N_2380,N_1920,N_1902);
or U2381 (N_2381,N_1858,N_1604);
xnor U2382 (N_2382,N_1734,N_1726);
xor U2383 (N_2383,N_1796,N_1558);
nand U2384 (N_2384,N_1716,N_1816);
or U2385 (N_2385,N_1984,N_1956);
or U2386 (N_2386,N_1818,N_1873);
nor U2387 (N_2387,N_1818,N_1843);
nand U2388 (N_2388,N_1822,N_1735);
nand U2389 (N_2389,N_1613,N_1708);
nor U2390 (N_2390,N_1867,N_1928);
and U2391 (N_2391,N_1511,N_1586);
and U2392 (N_2392,N_1814,N_1932);
and U2393 (N_2393,N_1860,N_1708);
and U2394 (N_2394,N_1696,N_1532);
or U2395 (N_2395,N_1908,N_1668);
and U2396 (N_2396,N_1514,N_1864);
or U2397 (N_2397,N_1556,N_1701);
nand U2398 (N_2398,N_1895,N_1858);
and U2399 (N_2399,N_1569,N_1961);
xnor U2400 (N_2400,N_1962,N_1736);
nor U2401 (N_2401,N_1787,N_1972);
nand U2402 (N_2402,N_1845,N_1542);
nor U2403 (N_2403,N_1582,N_1576);
and U2404 (N_2404,N_1991,N_1872);
nand U2405 (N_2405,N_1864,N_1937);
or U2406 (N_2406,N_1711,N_1986);
and U2407 (N_2407,N_1631,N_1657);
nor U2408 (N_2408,N_1785,N_1664);
or U2409 (N_2409,N_1500,N_1573);
or U2410 (N_2410,N_1650,N_1938);
nor U2411 (N_2411,N_1734,N_1710);
or U2412 (N_2412,N_1829,N_1707);
and U2413 (N_2413,N_1853,N_1718);
nor U2414 (N_2414,N_1803,N_1716);
and U2415 (N_2415,N_1813,N_1733);
nand U2416 (N_2416,N_1722,N_1891);
and U2417 (N_2417,N_1926,N_1733);
or U2418 (N_2418,N_1589,N_1835);
nor U2419 (N_2419,N_1825,N_1594);
nor U2420 (N_2420,N_1518,N_1854);
nand U2421 (N_2421,N_1751,N_1608);
or U2422 (N_2422,N_1642,N_1501);
and U2423 (N_2423,N_1690,N_1978);
and U2424 (N_2424,N_1676,N_1862);
nand U2425 (N_2425,N_1573,N_1713);
or U2426 (N_2426,N_1546,N_1653);
nand U2427 (N_2427,N_1705,N_1595);
nand U2428 (N_2428,N_1677,N_1710);
or U2429 (N_2429,N_1897,N_1695);
or U2430 (N_2430,N_1883,N_1649);
nor U2431 (N_2431,N_1766,N_1935);
nor U2432 (N_2432,N_1779,N_1944);
and U2433 (N_2433,N_1526,N_1777);
nand U2434 (N_2434,N_1584,N_1662);
nor U2435 (N_2435,N_1708,N_1561);
nand U2436 (N_2436,N_1591,N_1607);
nand U2437 (N_2437,N_1819,N_1898);
or U2438 (N_2438,N_1677,N_1569);
and U2439 (N_2439,N_1540,N_1803);
and U2440 (N_2440,N_1963,N_1874);
or U2441 (N_2441,N_1742,N_1759);
nor U2442 (N_2442,N_1725,N_1537);
nand U2443 (N_2443,N_1982,N_1601);
nor U2444 (N_2444,N_1719,N_1676);
nor U2445 (N_2445,N_1691,N_1530);
nand U2446 (N_2446,N_1920,N_1863);
and U2447 (N_2447,N_1869,N_1793);
nor U2448 (N_2448,N_1690,N_1518);
nand U2449 (N_2449,N_1929,N_1511);
nor U2450 (N_2450,N_1533,N_1550);
xnor U2451 (N_2451,N_1788,N_1957);
and U2452 (N_2452,N_1668,N_1794);
nor U2453 (N_2453,N_1532,N_1855);
xor U2454 (N_2454,N_1521,N_1828);
and U2455 (N_2455,N_1938,N_1996);
and U2456 (N_2456,N_1738,N_1560);
or U2457 (N_2457,N_1566,N_1895);
or U2458 (N_2458,N_1594,N_1894);
or U2459 (N_2459,N_1968,N_1744);
or U2460 (N_2460,N_1700,N_1914);
or U2461 (N_2461,N_1725,N_1733);
and U2462 (N_2462,N_1748,N_1843);
nand U2463 (N_2463,N_1744,N_1682);
nand U2464 (N_2464,N_1991,N_1966);
nand U2465 (N_2465,N_1826,N_1928);
nand U2466 (N_2466,N_1532,N_1990);
xnor U2467 (N_2467,N_1963,N_1753);
nor U2468 (N_2468,N_1716,N_1573);
nand U2469 (N_2469,N_1529,N_1915);
or U2470 (N_2470,N_1800,N_1875);
xnor U2471 (N_2471,N_1799,N_1965);
nor U2472 (N_2472,N_1823,N_1584);
or U2473 (N_2473,N_1763,N_1793);
nand U2474 (N_2474,N_1587,N_1957);
nor U2475 (N_2475,N_1782,N_1883);
and U2476 (N_2476,N_1977,N_1922);
nand U2477 (N_2477,N_1793,N_1613);
nor U2478 (N_2478,N_1570,N_1622);
nand U2479 (N_2479,N_1582,N_1676);
and U2480 (N_2480,N_1785,N_1734);
and U2481 (N_2481,N_1818,N_1507);
or U2482 (N_2482,N_1574,N_1875);
nand U2483 (N_2483,N_1844,N_1772);
xor U2484 (N_2484,N_1753,N_1965);
nor U2485 (N_2485,N_1763,N_1676);
or U2486 (N_2486,N_1831,N_1932);
and U2487 (N_2487,N_1833,N_1910);
nor U2488 (N_2488,N_1590,N_1914);
nor U2489 (N_2489,N_1912,N_1928);
nor U2490 (N_2490,N_1813,N_1871);
xnor U2491 (N_2491,N_1549,N_1895);
and U2492 (N_2492,N_1975,N_1856);
nand U2493 (N_2493,N_1752,N_1704);
nor U2494 (N_2494,N_1983,N_1644);
and U2495 (N_2495,N_1909,N_1820);
and U2496 (N_2496,N_1922,N_1852);
nor U2497 (N_2497,N_1789,N_1834);
or U2498 (N_2498,N_1669,N_1932);
nand U2499 (N_2499,N_1973,N_1551);
xnor U2500 (N_2500,N_2034,N_2232);
and U2501 (N_2501,N_2166,N_2271);
nand U2502 (N_2502,N_2195,N_2421);
or U2503 (N_2503,N_2458,N_2165);
and U2504 (N_2504,N_2192,N_2248);
nor U2505 (N_2505,N_2100,N_2368);
nand U2506 (N_2506,N_2099,N_2460);
or U2507 (N_2507,N_2146,N_2325);
nand U2508 (N_2508,N_2225,N_2019);
xnor U2509 (N_2509,N_2080,N_2183);
nand U2510 (N_2510,N_2212,N_2436);
nand U2511 (N_2511,N_2360,N_2109);
nor U2512 (N_2512,N_2367,N_2001);
and U2513 (N_2513,N_2017,N_2151);
and U2514 (N_2514,N_2011,N_2237);
nand U2515 (N_2515,N_2187,N_2293);
nor U2516 (N_2516,N_2224,N_2209);
or U2517 (N_2517,N_2089,N_2364);
nand U2518 (N_2518,N_2023,N_2198);
xnor U2519 (N_2519,N_2074,N_2136);
or U2520 (N_2520,N_2217,N_2082);
and U2521 (N_2521,N_2318,N_2277);
nor U2522 (N_2522,N_2407,N_2204);
and U2523 (N_2523,N_2384,N_2363);
nor U2524 (N_2524,N_2193,N_2276);
or U2525 (N_2525,N_2130,N_2266);
nor U2526 (N_2526,N_2274,N_2490);
nand U2527 (N_2527,N_2475,N_2438);
nor U2528 (N_2528,N_2372,N_2067);
or U2529 (N_2529,N_2284,N_2437);
nand U2530 (N_2530,N_2261,N_2115);
nand U2531 (N_2531,N_2466,N_2079);
nand U2532 (N_2532,N_2083,N_2194);
or U2533 (N_2533,N_2441,N_2341);
nor U2534 (N_2534,N_2162,N_2457);
nand U2535 (N_2535,N_2219,N_2215);
nor U2536 (N_2536,N_2308,N_2072);
nand U2537 (N_2537,N_2478,N_2331);
nor U2538 (N_2538,N_2294,N_2223);
or U2539 (N_2539,N_2035,N_2472);
or U2540 (N_2540,N_2141,N_2288);
or U2541 (N_2541,N_2428,N_2290);
and U2542 (N_2542,N_2137,N_2477);
xor U2543 (N_2543,N_2059,N_2275);
nor U2544 (N_2544,N_2126,N_2062);
xnor U2545 (N_2545,N_2312,N_2401);
or U2546 (N_2546,N_2201,N_2482);
xor U2547 (N_2547,N_2174,N_2152);
and U2548 (N_2548,N_2203,N_2040);
nand U2549 (N_2549,N_2353,N_2221);
nor U2550 (N_2550,N_2255,N_2425);
nor U2551 (N_2551,N_2296,N_2028);
nor U2552 (N_2552,N_2333,N_2461);
and U2553 (N_2553,N_2426,N_2159);
nor U2554 (N_2554,N_2263,N_2265);
and U2555 (N_2555,N_2379,N_2326);
and U2556 (N_2556,N_2065,N_2156);
nand U2557 (N_2557,N_2309,N_2434);
nor U2558 (N_2558,N_2007,N_2344);
nor U2559 (N_2559,N_2200,N_2279);
and U2560 (N_2560,N_2205,N_2238);
and U2561 (N_2561,N_2359,N_2234);
nand U2562 (N_2562,N_2345,N_2061);
nor U2563 (N_2563,N_2492,N_2487);
nand U2564 (N_2564,N_2108,N_2066);
nor U2565 (N_2565,N_2252,N_2375);
nor U2566 (N_2566,N_2105,N_2085);
or U2567 (N_2567,N_2496,N_2448);
xor U2568 (N_2568,N_2262,N_2471);
nand U2569 (N_2569,N_2175,N_2180);
xnor U2570 (N_2570,N_2332,N_2420);
or U2571 (N_2571,N_2354,N_2171);
nand U2572 (N_2572,N_2486,N_2469);
xnor U2573 (N_2573,N_2021,N_2050);
or U2574 (N_2574,N_2036,N_2418);
xnor U2575 (N_2575,N_2039,N_2207);
nor U2576 (N_2576,N_2150,N_2387);
nand U2577 (N_2577,N_2087,N_2303);
or U2578 (N_2578,N_2244,N_2411);
and U2579 (N_2579,N_2058,N_2348);
and U2580 (N_2580,N_2154,N_2101);
nand U2581 (N_2581,N_2328,N_2315);
and U2582 (N_2582,N_2313,N_2031);
and U2583 (N_2583,N_2049,N_2003);
or U2584 (N_2584,N_2107,N_2385);
or U2585 (N_2585,N_2015,N_2163);
or U2586 (N_2586,N_2455,N_2446);
or U2587 (N_2587,N_2149,N_2467);
nand U2588 (N_2588,N_2169,N_2301);
nor U2589 (N_2589,N_2230,N_2435);
or U2590 (N_2590,N_2063,N_2396);
nand U2591 (N_2591,N_2226,N_2386);
xnor U2592 (N_2592,N_2153,N_2071);
and U2593 (N_2593,N_2374,N_2316);
nand U2594 (N_2594,N_2051,N_2132);
nor U2595 (N_2595,N_2135,N_2433);
xor U2596 (N_2596,N_2283,N_2016);
nand U2597 (N_2597,N_2336,N_2213);
nand U2598 (N_2598,N_2114,N_2369);
nand U2599 (N_2599,N_2306,N_2362);
nor U2600 (N_2600,N_2009,N_2351);
or U2601 (N_2601,N_2260,N_2432);
nor U2602 (N_2602,N_2291,N_2229);
or U2603 (N_2603,N_2033,N_2392);
nand U2604 (N_2604,N_2366,N_2139);
and U2605 (N_2605,N_2349,N_2431);
nor U2606 (N_2606,N_2267,N_2117);
and U2607 (N_2607,N_2177,N_2417);
or U2608 (N_2608,N_2086,N_2214);
nor U2609 (N_2609,N_2254,N_2498);
and U2610 (N_2610,N_2479,N_2299);
nand U2611 (N_2611,N_2454,N_2416);
and U2612 (N_2612,N_2297,N_2305);
and U2613 (N_2613,N_2451,N_2122);
nand U2614 (N_2614,N_2464,N_2184);
and U2615 (N_2615,N_2389,N_2352);
nor U2616 (N_2616,N_2269,N_2022);
nor U2617 (N_2617,N_2282,N_2358);
or U2618 (N_2618,N_2295,N_2145);
xor U2619 (N_2619,N_2096,N_2335);
nand U2620 (N_2620,N_2347,N_2327);
nor U2621 (N_2621,N_2320,N_2340);
xnor U2622 (N_2622,N_2032,N_2323);
nor U2623 (N_2623,N_2125,N_2140);
or U2624 (N_2624,N_2172,N_2468);
or U2625 (N_2625,N_2413,N_2168);
and U2626 (N_2626,N_2285,N_2024);
and U2627 (N_2627,N_2245,N_2047);
or U2628 (N_2628,N_2013,N_2185);
and U2629 (N_2629,N_2106,N_2118);
nor U2630 (N_2630,N_2410,N_2112);
xor U2631 (N_2631,N_2134,N_2403);
or U2632 (N_2632,N_2429,N_2148);
nand U2633 (N_2633,N_2251,N_2493);
or U2634 (N_2634,N_2330,N_2317);
xnor U2635 (N_2635,N_2488,N_2197);
nor U2636 (N_2636,N_2361,N_2060);
nand U2637 (N_2637,N_2445,N_2414);
nor U2638 (N_2638,N_2300,N_2239);
xor U2639 (N_2639,N_2038,N_2246);
or U2640 (N_2640,N_2220,N_2444);
and U2641 (N_2641,N_2129,N_2030);
nand U2642 (N_2642,N_2131,N_2005);
nand U2643 (N_2643,N_2116,N_2055);
nor U2644 (N_2644,N_2018,N_2439);
and U2645 (N_2645,N_2324,N_2409);
xor U2646 (N_2646,N_2173,N_2481);
and U2647 (N_2647,N_2391,N_2376);
nand U2648 (N_2648,N_2272,N_2415);
nand U2649 (N_2649,N_2287,N_2462);
nand U2650 (N_2650,N_2405,N_2102);
nor U2651 (N_2651,N_2259,N_2243);
or U2652 (N_2652,N_2233,N_2449);
nor U2653 (N_2653,N_2042,N_2302);
or U2654 (N_2654,N_2247,N_2227);
and U2655 (N_2655,N_2064,N_2075);
nand U2656 (N_2656,N_2371,N_2278);
nor U2657 (N_2657,N_2499,N_2393);
or U2658 (N_2658,N_2158,N_2133);
and U2659 (N_2659,N_2043,N_2273);
and U2660 (N_2660,N_2378,N_2390);
or U2661 (N_2661,N_2179,N_2286);
nor U2662 (N_2662,N_2104,N_2406);
nand U2663 (N_2663,N_2440,N_2073);
and U2664 (N_2664,N_2298,N_2176);
and U2665 (N_2665,N_2138,N_2191);
nand U2666 (N_2666,N_2497,N_2000);
nor U2667 (N_2667,N_2381,N_2394);
and U2668 (N_2668,N_2143,N_2164);
nor U2669 (N_2669,N_2268,N_2076);
and U2670 (N_2670,N_2399,N_2370);
nand U2671 (N_2671,N_2250,N_2356);
and U2672 (N_2672,N_2070,N_2014);
and U2673 (N_2673,N_2447,N_2029);
nand U2674 (N_2674,N_2483,N_2020);
or U2675 (N_2675,N_2474,N_2357);
or U2676 (N_2676,N_2170,N_2218);
nand U2677 (N_2677,N_2453,N_2480);
nor U2678 (N_2678,N_2397,N_2144);
xor U2679 (N_2679,N_2319,N_2402);
nor U2680 (N_2680,N_2321,N_2121);
nor U2681 (N_2681,N_2157,N_2311);
nor U2682 (N_2682,N_2228,N_2006);
or U2683 (N_2683,N_2377,N_2068);
or U2684 (N_2684,N_2098,N_2091);
or U2685 (N_2685,N_2264,N_2240);
and U2686 (N_2686,N_2056,N_2078);
nor U2687 (N_2687,N_2452,N_2186);
nand U2688 (N_2688,N_2182,N_2343);
nand U2689 (N_2689,N_2476,N_2419);
nand U2690 (N_2690,N_2037,N_2189);
or U2691 (N_2691,N_2494,N_2155);
or U2692 (N_2692,N_2092,N_2337);
nor U2693 (N_2693,N_2142,N_2124);
or U2694 (N_2694,N_2491,N_2242);
xnor U2695 (N_2695,N_2008,N_2206);
or U2696 (N_2696,N_2280,N_2463);
or U2697 (N_2697,N_2094,N_2258);
nor U2698 (N_2698,N_2342,N_2211);
nor U2699 (N_2699,N_2196,N_2188);
or U2700 (N_2700,N_2012,N_2160);
nand U2701 (N_2701,N_2257,N_2057);
xnor U2702 (N_2702,N_2365,N_2256);
or U2703 (N_2703,N_2495,N_2382);
nand U2704 (N_2704,N_2281,N_2178);
nor U2705 (N_2705,N_2427,N_2222);
nand U2706 (N_2706,N_2010,N_2161);
and U2707 (N_2707,N_2235,N_2270);
xnor U2708 (N_2708,N_2470,N_2090);
xor U2709 (N_2709,N_2190,N_2123);
or U2710 (N_2710,N_2373,N_2334);
nand U2711 (N_2711,N_2119,N_2304);
nand U2712 (N_2712,N_2048,N_2484);
or U2713 (N_2713,N_2045,N_2128);
nand U2714 (N_2714,N_2400,N_2430);
or U2715 (N_2715,N_2465,N_2081);
nor U2716 (N_2716,N_2111,N_2292);
nor U2717 (N_2717,N_2167,N_2088);
and U2718 (N_2718,N_2054,N_2077);
nand U2719 (N_2719,N_2026,N_2307);
or U2720 (N_2720,N_2025,N_2355);
nand U2721 (N_2721,N_2241,N_2113);
and U2722 (N_2722,N_2084,N_2044);
nor U2723 (N_2723,N_2422,N_2346);
nor U2724 (N_2724,N_2052,N_2404);
nand U2725 (N_2725,N_2459,N_2450);
or U2726 (N_2726,N_2046,N_2199);
nand U2727 (N_2727,N_2069,N_2395);
nand U2728 (N_2728,N_2443,N_2380);
nand U2729 (N_2729,N_2103,N_2095);
nor U2730 (N_2730,N_2208,N_2423);
xnor U2731 (N_2731,N_2210,N_2489);
nor U2732 (N_2732,N_2339,N_2202);
xnor U2733 (N_2733,N_2097,N_2442);
and U2734 (N_2734,N_2424,N_2485);
and U2735 (N_2735,N_2002,N_2249);
or U2736 (N_2736,N_2093,N_2027);
or U2737 (N_2737,N_2289,N_2398);
or U2738 (N_2738,N_2127,N_2053);
nand U2739 (N_2739,N_2147,N_2216);
nor U2740 (N_2740,N_2473,N_2412);
and U2741 (N_2741,N_2329,N_2383);
and U2742 (N_2742,N_2041,N_2408);
nor U2743 (N_2743,N_2350,N_2236);
or U2744 (N_2744,N_2456,N_2004);
nand U2745 (N_2745,N_2314,N_2181);
nor U2746 (N_2746,N_2322,N_2231);
and U2747 (N_2747,N_2388,N_2253);
nand U2748 (N_2748,N_2338,N_2110);
and U2749 (N_2749,N_2120,N_2310);
nand U2750 (N_2750,N_2480,N_2289);
nand U2751 (N_2751,N_2452,N_2243);
nand U2752 (N_2752,N_2398,N_2331);
or U2753 (N_2753,N_2327,N_2093);
nor U2754 (N_2754,N_2440,N_2003);
xnor U2755 (N_2755,N_2353,N_2443);
nor U2756 (N_2756,N_2030,N_2465);
and U2757 (N_2757,N_2247,N_2162);
nor U2758 (N_2758,N_2061,N_2350);
nor U2759 (N_2759,N_2153,N_2303);
xor U2760 (N_2760,N_2306,N_2357);
xor U2761 (N_2761,N_2262,N_2378);
or U2762 (N_2762,N_2201,N_2044);
nor U2763 (N_2763,N_2285,N_2484);
nand U2764 (N_2764,N_2237,N_2017);
or U2765 (N_2765,N_2489,N_2461);
nand U2766 (N_2766,N_2051,N_2034);
nand U2767 (N_2767,N_2285,N_2183);
and U2768 (N_2768,N_2012,N_2180);
xnor U2769 (N_2769,N_2326,N_2189);
or U2770 (N_2770,N_2374,N_2278);
xnor U2771 (N_2771,N_2084,N_2241);
or U2772 (N_2772,N_2058,N_2264);
nor U2773 (N_2773,N_2249,N_2243);
or U2774 (N_2774,N_2476,N_2215);
nand U2775 (N_2775,N_2377,N_2217);
xor U2776 (N_2776,N_2440,N_2306);
or U2777 (N_2777,N_2157,N_2371);
nor U2778 (N_2778,N_2077,N_2397);
nor U2779 (N_2779,N_2428,N_2397);
and U2780 (N_2780,N_2024,N_2286);
nand U2781 (N_2781,N_2004,N_2269);
xnor U2782 (N_2782,N_2414,N_2449);
and U2783 (N_2783,N_2402,N_2222);
nor U2784 (N_2784,N_2095,N_2489);
nor U2785 (N_2785,N_2458,N_2393);
nor U2786 (N_2786,N_2303,N_2026);
or U2787 (N_2787,N_2496,N_2341);
nor U2788 (N_2788,N_2443,N_2338);
xnor U2789 (N_2789,N_2374,N_2275);
or U2790 (N_2790,N_2391,N_2392);
xor U2791 (N_2791,N_2354,N_2046);
and U2792 (N_2792,N_2394,N_2226);
xnor U2793 (N_2793,N_2108,N_2329);
nand U2794 (N_2794,N_2275,N_2437);
nand U2795 (N_2795,N_2374,N_2416);
or U2796 (N_2796,N_2372,N_2306);
and U2797 (N_2797,N_2158,N_2482);
nor U2798 (N_2798,N_2095,N_2055);
nand U2799 (N_2799,N_2025,N_2041);
nand U2800 (N_2800,N_2287,N_2110);
and U2801 (N_2801,N_2244,N_2269);
xor U2802 (N_2802,N_2331,N_2477);
nand U2803 (N_2803,N_2367,N_2226);
and U2804 (N_2804,N_2379,N_2139);
and U2805 (N_2805,N_2382,N_2246);
nor U2806 (N_2806,N_2350,N_2396);
nand U2807 (N_2807,N_2267,N_2426);
xor U2808 (N_2808,N_2486,N_2051);
and U2809 (N_2809,N_2245,N_2324);
nand U2810 (N_2810,N_2482,N_2105);
nor U2811 (N_2811,N_2014,N_2265);
nor U2812 (N_2812,N_2320,N_2295);
or U2813 (N_2813,N_2379,N_2468);
and U2814 (N_2814,N_2453,N_2012);
xor U2815 (N_2815,N_2160,N_2125);
nand U2816 (N_2816,N_2007,N_2090);
nand U2817 (N_2817,N_2460,N_2356);
xor U2818 (N_2818,N_2245,N_2381);
or U2819 (N_2819,N_2351,N_2418);
nor U2820 (N_2820,N_2088,N_2128);
xor U2821 (N_2821,N_2299,N_2347);
or U2822 (N_2822,N_2296,N_2026);
nor U2823 (N_2823,N_2185,N_2287);
or U2824 (N_2824,N_2063,N_2202);
nand U2825 (N_2825,N_2142,N_2092);
nor U2826 (N_2826,N_2036,N_2483);
or U2827 (N_2827,N_2485,N_2284);
nand U2828 (N_2828,N_2464,N_2102);
and U2829 (N_2829,N_2175,N_2416);
or U2830 (N_2830,N_2181,N_2308);
or U2831 (N_2831,N_2480,N_2096);
and U2832 (N_2832,N_2306,N_2054);
and U2833 (N_2833,N_2190,N_2061);
or U2834 (N_2834,N_2227,N_2281);
and U2835 (N_2835,N_2326,N_2378);
nor U2836 (N_2836,N_2157,N_2403);
nand U2837 (N_2837,N_2451,N_2372);
xnor U2838 (N_2838,N_2153,N_2083);
nor U2839 (N_2839,N_2124,N_2090);
nor U2840 (N_2840,N_2333,N_2004);
or U2841 (N_2841,N_2165,N_2386);
and U2842 (N_2842,N_2010,N_2486);
nand U2843 (N_2843,N_2389,N_2147);
and U2844 (N_2844,N_2038,N_2070);
and U2845 (N_2845,N_2412,N_2439);
xor U2846 (N_2846,N_2232,N_2191);
nand U2847 (N_2847,N_2308,N_2289);
nand U2848 (N_2848,N_2414,N_2366);
nor U2849 (N_2849,N_2417,N_2181);
nor U2850 (N_2850,N_2470,N_2223);
or U2851 (N_2851,N_2126,N_2450);
and U2852 (N_2852,N_2370,N_2014);
nor U2853 (N_2853,N_2091,N_2415);
nand U2854 (N_2854,N_2316,N_2157);
nor U2855 (N_2855,N_2179,N_2307);
nand U2856 (N_2856,N_2119,N_2000);
or U2857 (N_2857,N_2061,N_2197);
or U2858 (N_2858,N_2152,N_2185);
or U2859 (N_2859,N_2253,N_2042);
nand U2860 (N_2860,N_2273,N_2395);
and U2861 (N_2861,N_2361,N_2049);
nor U2862 (N_2862,N_2202,N_2494);
nand U2863 (N_2863,N_2167,N_2268);
nand U2864 (N_2864,N_2135,N_2322);
and U2865 (N_2865,N_2492,N_2141);
nand U2866 (N_2866,N_2402,N_2412);
and U2867 (N_2867,N_2413,N_2077);
nor U2868 (N_2868,N_2398,N_2199);
nand U2869 (N_2869,N_2141,N_2189);
or U2870 (N_2870,N_2165,N_2472);
and U2871 (N_2871,N_2000,N_2462);
xor U2872 (N_2872,N_2057,N_2141);
nand U2873 (N_2873,N_2185,N_2327);
and U2874 (N_2874,N_2003,N_2225);
nor U2875 (N_2875,N_2035,N_2401);
nor U2876 (N_2876,N_2308,N_2237);
and U2877 (N_2877,N_2346,N_2106);
nor U2878 (N_2878,N_2126,N_2433);
or U2879 (N_2879,N_2306,N_2197);
and U2880 (N_2880,N_2266,N_2489);
nand U2881 (N_2881,N_2096,N_2240);
nor U2882 (N_2882,N_2474,N_2488);
nor U2883 (N_2883,N_2179,N_2041);
and U2884 (N_2884,N_2058,N_2295);
or U2885 (N_2885,N_2139,N_2034);
or U2886 (N_2886,N_2380,N_2363);
or U2887 (N_2887,N_2160,N_2327);
nand U2888 (N_2888,N_2115,N_2450);
or U2889 (N_2889,N_2174,N_2269);
nand U2890 (N_2890,N_2020,N_2361);
and U2891 (N_2891,N_2272,N_2269);
nor U2892 (N_2892,N_2442,N_2420);
xor U2893 (N_2893,N_2176,N_2303);
nand U2894 (N_2894,N_2184,N_2097);
xnor U2895 (N_2895,N_2189,N_2099);
nand U2896 (N_2896,N_2116,N_2403);
and U2897 (N_2897,N_2233,N_2140);
and U2898 (N_2898,N_2117,N_2063);
xor U2899 (N_2899,N_2084,N_2081);
nor U2900 (N_2900,N_2309,N_2414);
or U2901 (N_2901,N_2451,N_2103);
nor U2902 (N_2902,N_2209,N_2260);
and U2903 (N_2903,N_2223,N_2457);
and U2904 (N_2904,N_2304,N_2408);
nand U2905 (N_2905,N_2174,N_2162);
nor U2906 (N_2906,N_2162,N_2001);
xor U2907 (N_2907,N_2233,N_2184);
or U2908 (N_2908,N_2216,N_2432);
xnor U2909 (N_2909,N_2222,N_2175);
and U2910 (N_2910,N_2303,N_2369);
or U2911 (N_2911,N_2470,N_2251);
nand U2912 (N_2912,N_2477,N_2114);
and U2913 (N_2913,N_2235,N_2352);
or U2914 (N_2914,N_2087,N_2467);
or U2915 (N_2915,N_2280,N_2299);
nand U2916 (N_2916,N_2075,N_2346);
nor U2917 (N_2917,N_2077,N_2151);
nand U2918 (N_2918,N_2201,N_2115);
and U2919 (N_2919,N_2381,N_2413);
or U2920 (N_2920,N_2112,N_2052);
or U2921 (N_2921,N_2304,N_2151);
nor U2922 (N_2922,N_2434,N_2326);
xor U2923 (N_2923,N_2078,N_2117);
or U2924 (N_2924,N_2038,N_2391);
and U2925 (N_2925,N_2492,N_2058);
and U2926 (N_2926,N_2481,N_2084);
or U2927 (N_2927,N_2009,N_2195);
nor U2928 (N_2928,N_2490,N_2180);
and U2929 (N_2929,N_2490,N_2382);
nand U2930 (N_2930,N_2041,N_2069);
or U2931 (N_2931,N_2287,N_2359);
or U2932 (N_2932,N_2402,N_2218);
nand U2933 (N_2933,N_2343,N_2107);
nand U2934 (N_2934,N_2273,N_2369);
or U2935 (N_2935,N_2393,N_2467);
nand U2936 (N_2936,N_2207,N_2186);
and U2937 (N_2937,N_2123,N_2168);
and U2938 (N_2938,N_2266,N_2128);
or U2939 (N_2939,N_2471,N_2096);
or U2940 (N_2940,N_2486,N_2156);
xor U2941 (N_2941,N_2266,N_2458);
xor U2942 (N_2942,N_2243,N_2109);
or U2943 (N_2943,N_2029,N_2426);
xnor U2944 (N_2944,N_2039,N_2019);
and U2945 (N_2945,N_2243,N_2307);
or U2946 (N_2946,N_2430,N_2217);
nand U2947 (N_2947,N_2225,N_2480);
xor U2948 (N_2948,N_2108,N_2128);
nor U2949 (N_2949,N_2487,N_2368);
or U2950 (N_2950,N_2144,N_2056);
nand U2951 (N_2951,N_2419,N_2349);
or U2952 (N_2952,N_2079,N_2248);
nor U2953 (N_2953,N_2347,N_2328);
or U2954 (N_2954,N_2449,N_2138);
nor U2955 (N_2955,N_2302,N_2287);
and U2956 (N_2956,N_2378,N_2138);
or U2957 (N_2957,N_2102,N_2371);
or U2958 (N_2958,N_2354,N_2349);
nand U2959 (N_2959,N_2100,N_2403);
and U2960 (N_2960,N_2252,N_2171);
and U2961 (N_2961,N_2316,N_2458);
and U2962 (N_2962,N_2097,N_2075);
or U2963 (N_2963,N_2065,N_2123);
or U2964 (N_2964,N_2000,N_2300);
or U2965 (N_2965,N_2413,N_2289);
or U2966 (N_2966,N_2469,N_2329);
or U2967 (N_2967,N_2442,N_2177);
nand U2968 (N_2968,N_2040,N_2469);
or U2969 (N_2969,N_2335,N_2146);
nand U2970 (N_2970,N_2434,N_2497);
nor U2971 (N_2971,N_2486,N_2069);
or U2972 (N_2972,N_2266,N_2272);
and U2973 (N_2973,N_2047,N_2213);
and U2974 (N_2974,N_2236,N_2123);
nor U2975 (N_2975,N_2118,N_2122);
nand U2976 (N_2976,N_2387,N_2456);
and U2977 (N_2977,N_2434,N_2355);
and U2978 (N_2978,N_2164,N_2367);
nand U2979 (N_2979,N_2083,N_2053);
nand U2980 (N_2980,N_2372,N_2001);
nor U2981 (N_2981,N_2367,N_2393);
or U2982 (N_2982,N_2318,N_2061);
or U2983 (N_2983,N_2131,N_2464);
nor U2984 (N_2984,N_2239,N_2011);
or U2985 (N_2985,N_2347,N_2318);
xnor U2986 (N_2986,N_2069,N_2407);
nand U2987 (N_2987,N_2401,N_2174);
nor U2988 (N_2988,N_2289,N_2474);
nand U2989 (N_2989,N_2472,N_2293);
nand U2990 (N_2990,N_2212,N_2007);
nand U2991 (N_2991,N_2440,N_2240);
or U2992 (N_2992,N_2334,N_2031);
nor U2993 (N_2993,N_2192,N_2113);
and U2994 (N_2994,N_2279,N_2238);
and U2995 (N_2995,N_2371,N_2208);
nor U2996 (N_2996,N_2454,N_2373);
or U2997 (N_2997,N_2497,N_2157);
xnor U2998 (N_2998,N_2110,N_2346);
or U2999 (N_2999,N_2119,N_2056);
nand U3000 (N_3000,N_2534,N_2781);
nand U3001 (N_3001,N_2521,N_2869);
xor U3002 (N_3002,N_2526,N_2801);
and U3003 (N_3003,N_2907,N_2537);
and U3004 (N_3004,N_2666,N_2562);
and U3005 (N_3005,N_2798,N_2807);
nor U3006 (N_3006,N_2620,N_2552);
or U3007 (N_3007,N_2993,N_2613);
and U3008 (N_3008,N_2771,N_2850);
nor U3009 (N_3009,N_2951,N_2877);
and U3010 (N_3010,N_2621,N_2797);
or U3011 (N_3011,N_2864,N_2954);
nor U3012 (N_3012,N_2512,N_2586);
or U3013 (N_3013,N_2751,N_2911);
nor U3014 (N_3014,N_2971,N_2626);
nand U3015 (N_3015,N_2873,N_2674);
xnor U3016 (N_3016,N_2592,N_2769);
nor U3017 (N_3017,N_2766,N_2573);
or U3018 (N_3018,N_2790,N_2646);
nor U3019 (N_3019,N_2729,N_2680);
and U3020 (N_3020,N_2833,N_2632);
nor U3021 (N_3021,N_2655,N_2831);
or U3022 (N_3022,N_2861,N_2882);
nor U3023 (N_3023,N_2890,N_2578);
nor U3024 (N_3024,N_2749,N_2881);
or U3025 (N_3025,N_2679,N_2788);
xor U3026 (N_3026,N_2709,N_2920);
nand U3027 (N_3027,N_2828,N_2683);
nor U3028 (N_3028,N_2803,N_2744);
nor U3029 (N_3029,N_2654,N_2970);
nor U3030 (N_3030,N_2530,N_2857);
nand U3031 (N_3031,N_2913,N_2564);
or U3032 (N_3032,N_2633,N_2746);
nand U3033 (N_3033,N_2956,N_2593);
xor U3034 (N_3034,N_2606,N_2952);
or U3035 (N_3035,N_2664,N_2967);
nand U3036 (N_3036,N_2717,N_2554);
and U3037 (N_3037,N_2539,N_2722);
or U3038 (N_3038,N_2663,N_2625);
or U3039 (N_3039,N_2533,N_2577);
nand U3040 (N_3040,N_2827,N_2763);
and U3041 (N_3041,N_2728,N_2906);
nor U3042 (N_3042,N_2692,N_2727);
or U3043 (N_3043,N_2768,N_2535);
and U3044 (N_3044,N_2600,N_2891);
or U3045 (N_3045,N_2931,N_2575);
xnor U3046 (N_3046,N_2884,N_2839);
or U3047 (N_3047,N_2942,N_2770);
xnor U3048 (N_3048,N_2567,N_2885);
nand U3049 (N_3049,N_2871,N_2550);
and U3050 (N_3050,N_2667,N_2838);
and U3051 (N_3051,N_2658,N_2962);
or U3052 (N_3052,N_2948,N_2914);
nand U3053 (N_3053,N_2514,N_2897);
nand U3054 (N_3054,N_2542,N_2583);
nor U3055 (N_3055,N_2739,N_2579);
or U3056 (N_3056,N_2826,N_2818);
or U3057 (N_3057,N_2947,N_2640);
nor U3058 (N_3058,N_2995,N_2983);
nor U3059 (N_3059,N_2689,N_2602);
or U3060 (N_3060,N_2693,N_2619);
nor U3061 (N_3061,N_2893,N_2662);
xor U3062 (N_3062,N_2509,N_2603);
and U3063 (N_3063,N_2946,N_2635);
nor U3064 (N_3064,N_2638,N_2915);
and U3065 (N_3065,N_2648,N_2989);
nand U3066 (N_3066,N_2782,N_2723);
and U3067 (N_3067,N_2794,N_2901);
or U3068 (N_3068,N_2713,N_2687);
nand U3069 (N_3069,N_2900,N_2529);
or U3070 (N_3070,N_2585,N_2960);
nor U3071 (N_3071,N_2531,N_2981);
nand U3072 (N_3072,N_2525,N_2651);
nor U3073 (N_3073,N_2936,N_2944);
nand U3074 (N_3074,N_2572,N_2966);
and U3075 (N_3075,N_2515,N_2580);
or U3076 (N_3076,N_2830,N_2725);
or U3077 (N_3077,N_2773,N_2842);
nand U3078 (N_3078,N_2819,N_2975);
and U3079 (N_3079,N_2916,N_2784);
nor U3080 (N_3080,N_2558,N_2817);
and U3081 (N_3081,N_2859,N_2779);
nor U3082 (N_3082,N_2671,N_2716);
or U3083 (N_3083,N_2935,N_2511);
nor U3084 (N_3084,N_2775,N_2776);
or U3085 (N_3085,N_2548,N_2595);
nand U3086 (N_3086,N_2591,N_2887);
nand U3087 (N_3087,N_2563,N_2841);
nand U3088 (N_3088,N_2642,N_2851);
nor U3089 (N_3089,N_2607,N_2933);
or U3090 (N_3090,N_2987,N_2661);
and U3091 (N_3091,N_2957,N_2825);
and U3092 (N_3092,N_2938,N_2734);
or U3093 (N_3093,N_2783,N_2964);
nor U3094 (N_3094,N_2852,N_2811);
nor U3095 (N_3095,N_2865,N_2502);
and U3096 (N_3096,N_2756,N_2866);
or U3097 (N_3097,N_2888,N_2574);
and U3098 (N_3098,N_2840,N_2556);
nand U3099 (N_3099,N_2611,N_2576);
or U3100 (N_3100,N_2919,N_2737);
and U3101 (N_3101,N_2999,N_2808);
xnor U3102 (N_3102,N_2774,N_2973);
or U3103 (N_3103,N_2868,N_2984);
or U3104 (N_3104,N_2681,N_2760);
and U3105 (N_3105,N_2872,N_2555);
or U3106 (N_3106,N_2753,N_2874);
xor U3107 (N_3107,N_2848,N_2581);
nor U3108 (N_3108,N_2924,N_2668);
nand U3109 (N_3109,N_2627,N_2615);
or U3110 (N_3110,N_2553,N_2714);
or U3111 (N_3111,N_2697,N_2785);
or U3112 (N_3112,N_2810,N_2707);
nand U3113 (N_3113,N_2650,N_2736);
nand U3114 (N_3114,N_2695,N_2812);
nand U3115 (N_3115,N_2718,N_2791);
or U3116 (N_3116,N_2898,N_2758);
or U3117 (N_3117,N_2623,N_2815);
and U3118 (N_3118,N_2880,N_2806);
and U3119 (N_3119,N_2832,N_2996);
or U3120 (N_3120,N_2904,N_2747);
nor U3121 (N_3121,N_2853,N_2943);
or U3122 (N_3122,N_2501,N_2672);
xor U3123 (N_3123,N_2802,N_2805);
or U3124 (N_3124,N_2703,N_2748);
nand U3125 (N_3125,N_2849,N_2657);
and U3126 (N_3126,N_2977,N_2767);
nand U3127 (N_3127,N_2757,N_2561);
or U3128 (N_3128,N_2738,N_2923);
nor U3129 (N_3129,N_2598,N_2641);
nand U3130 (N_3130,N_2837,N_2559);
nor U3131 (N_3131,N_2560,N_2653);
nor U3132 (N_3132,N_2990,N_2634);
and U3133 (N_3133,N_2959,N_2796);
nor U3134 (N_3134,N_2929,N_2862);
and U3135 (N_3135,N_2875,N_2659);
and U3136 (N_3136,N_2814,N_2590);
or U3137 (N_3137,N_2520,N_2597);
and U3138 (N_3138,N_2945,N_2712);
nor U3139 (N_3139,N_2986,N_2543);
and U3140 (N_3140,N_2675,N_2976);
nand U3141 (N_3141,N_2605,N_2587);
nor U3142 (N_3142,N_2510,N_2569);
nand U3143 (N_3143,N_2513,N_2961);
or U3144 (N_3144,N_2647,N_2980);
xnor U3145 (N_3145,N_2876,N_2541);
and U3146 (N_3146,N_2896,N_2596);
and U3147 (N_3147,N_2752,N_2545);
and U3148 (N_3148,N_2834,N_2557);
nor U3149 (N_3149,N_2816,N_2750);
and U3150 (N_3150,N_2799,N_2660);
and U3151 (N_3151,N_2649,N_2926);
nor U3152 (N_3152,N_2764,N_2604);
and U3153 (N_3153,N_2503,N_2965);
nand U3154 (N_3154,N_2892,N_2856);
nand U3155 (N_3155,N_2630,N_2677);
xor U3156 (N_3156,N_2844,N_2886);
and U3157 (N_3157,N_2795,N_2652);
nor U3158 (N_3158,N_2686,N_2691);
nor U3159 (N_3159,N_2594,N_2584);
or U3160 (N_3160,N_2628,N_2742);
nand U3161 (N_3161,N_2732,N_2883);
nand U3162 (N_3162,N_2889,N_2544);
nor U3163 (N_3163,N_2682,N_2870);
nor U3164 (N_3164,N_2616,N_2522);
and U3165 (N_3165,N_2762,N_2998);
nand U3166 (N_3166,N_2639,N_2684);
nand U3167 (N_3167,N_2822,N_2745);
or U3168 (N_3168,N_2787,N_2715);
and U3169 (N_3169,N_2972,N_2540);
nand U3170 (N_3170,N_2720,N_2932);
or U3171 (N_3171,N_2968,N_2710);
or U3172 (N_3172,N_2705,N_2608);
nor U3173 (N_3173,N_2676,N_2740);
xor U3174 (N_3174,N_2765,N_2517);
nand U3175 (N_3175,N_2800,N_2617);
nand U3176 (N_3176,N_2536,N_2912);
and U3177 (N_3177,N_2506,N_2867);
nand U3178 (N_3178,N_2702,N_2733);
nand U3179 (N_3179,N_2969,N_2994);
nor U3180 (N_3180,N_2988,N_2845);
nand U3181 (N_3181,N_2958,N_2527);
nor U3182 (N_3182,N_2982,N_2629);
and U3183 (N_3183,N_2846,N_2566);
and U3184 (N_3184,N_2631,N_2704);
nor U3185 (N_3185,N_2637,N_2588);
nand U3186 (N_3186,N_2847,N_2928);
nor U3187 (N_3187,N_2879,N_2902);
or U3188 (N_3188,N_2601,N_2645);
or U3189 (N_3189,N_2711,N_2665);
and U3190 (N_3190,N_2829,N_2524);
nor U3191 (N_3191,N_2698,N_2789);
and U3192 (N_3192,N_2792,N_2532);
or U3193 (N_3193,N_2690,N_2612);
nand U3194 (N_3194,N_2644,N_2974);
and U3195 (N_3195,N_2979,N_2685);
xor U3196 (N_3196,N_2528,N_2978);
xnor U3197 (N_3197,N_2854,N_2772);
nand U3198 (N_3198,N_2599,N_2820);
and U3199 (N_3199,N_2937,N_2678);
nand U3200 (N_3200,N_2699,N_2908);
xnor U3201 (N_3201,N_2508,N_2985);
nor U3202 (N_3202,N_2934,N_2696);
or U3203 (N_3203,N_2701,N_2836);
and U3204 (N_3204,N_2719,N_2504);
or U3205 (N_3205,N_2721,N_2878);
and U3206 (N_3206,N_2917,N_2571);
nand U3207 (N_3207,N_2963,N_2622);
nor U3208 (N_3208,N_2547,N_2505);
xnor U3209 (N_3209,N_2903,N_2918);
nand U3210 (N_3210,N_2700,N_2761);
and U3211 (N_3211,N_2743,N_2835);
or U3212 (N_3212,N_2921,N_2941);
and U3213 (N_3213,N_2804,N_2708);
nor U3214 (N_3214,N_2855,N_2565);
or U3215 (N_3215,N_2538,N_2939);
xnor U3216 (N_3216,N_2777,N_2930);
nor U3217 (N_3217,N_2636,N_2895);
nor U3218 (N_3218,N_2824,N_2991);
nand U3219 (N_3219,N_2910,N_2570);
nor U3220 (N_3220,N_2731,N_2780);
and U3221 (N_3221,N_2860,N_2656);
xor U3222 (N_3222,N_2519,N_2518);
nor U3223 (N_3223,N_2551,N_2741);
xnor U3224 (N_3224,N_2786,N_2992);
nand U3225 (N_3225,N_2670,N_2754);
nand U3226 (N_3226,N_2809,N_2500);
or U3227 (N_3227,N_2927,N_2955);
nand U3228 (N_3228,N_2823,N_2523);
nor U3229 (N_3229,N_2568,N_2759);
and U3230 (N_3230,N_2793,N_2863);
nor U3231 (N_3231,N_2858,N_2589);
and U3232 (N_3232,N_2894,N_2899);
nand U3233 (N_3233,N_2922,N_2516);
and U3234 (N_3234,N_2610,N_2673);
and U3235 (N_3235,N_2609,N_2813);
nand U3236 (N_3236,N_2706,N_2546);
or U3237 (N_3237,N_2950,N_2997);
or U3238 (N_3238,N_2755,N_2949);
or U3239 (N_3239,N_2724,N_2614);
and U3240 (N_3240,N_2735,N_2507);
and U3241 (N_3241,N_2730,N_2905);
or U3242 (N_3242,N_2688,N_2778);
and U3243 (N_3243,N_2726,N_2925);
or U3244 (N_3244,N_2618,N_2669);
and U3245 (N_3245,N_2643,N_2909);
nor U3246 (N_3246,N_2821,N_2549);
xor U3247 (N_3247,N_2694,N_2940);
nand U3248 (N_3248,N_2843,N_2953);
nor U3249 (N_3249,N_2582,N_2624);
nor U3250 (N_3250,N_2693,N_2962);
nand U3251 (N_3251,N_2500,N_2693);
xnor U3252 (N_3252,N_2795,N_2822);
xor U3253 (N_3253,N_2647,N_2843);
xnor U3254 (N_3254,N_2643,N_2622);
or U3255 (N_3255,N_2579,N_2559);
and U3256 (N_3256,N_2670,N_2820);
nand U3257 (N_3257,N_2829,N_2532);
or U3258 (N_3258,N_2537,N_2985);
nor U3259 (N_3259,N_2856,N_2631);
or U3260 (N_3260,N_2534,N_2724);
and U3261 (N_3261,N_2780,N_2619);
nor U3262 (N_3262,N_2659,N_2537);
xnor U3263 (N_3263,N_2533,N_2769);
nor U3264 (N_3264,N_2733,N_2599);
nand U3265 (N_3265,N_2616,N_2565);
or U3266 (N_3266,N_2992,N_2728);
and U3267 (N_3267,N_2738,N_2642);
nor U3268 (N_3268,N_2728,N_2816);
and U3269 (N_3269,N_2519,N_2671);
or U3270 (N_3270,N_2513,N_2909);
nand U3271 (N_3271,N_2790,N_2871);
nand U3272 (N_3272,N_2682,N_2787);
or U3273 (N_3273,N_2511,N_2701);
xnor U3274 (N_3274,N_2654,N_2743);
nand U3275 (N_3275,N_2905,N_2500);
or U3276 (N_3276,N_2851,N_2676);
and U3277 (N_3277,N_2946,N_2542);
or U3278 (N_3278,N_2855,N_2558);
or U3279 (N_3279,N_2916,N_2953);
and U3280 (N_3280,N_2834,N_2508);
or U3281 (N_3281,N_2916,N_2949);
xor U3282 (N_3282,N_2753,N_2904);
nor U3283 (N_3283,N_2869,N_2730);
xor U3284 (N_3284,N_2655,N_2925);
nand U3285 (N_3285,N_2943,N_2946);
and U3286 (N_3286,N_2671,N_2947);
or U3287 (N_3287,N_2548,N_2514);
or U3288 (N_3288,N_2514,N_2771);
and U3289 (N_3289,N_2744,N_2762);
nor U3290 (N_3290,N_2982,N_2700);
nand U3291 (N_3291,N_2600,N_2792);
nand U3292 (N_3292,N_2500,N_2977);
nor U3293 (N_3293,N_2916,N_2904);
nor U3294 (N_3294,N_2702,N_2567);
nand U3295 (N_3295,N_2933,N_2536);
and U3296 (N_3296,N_2593,N_2923);
or U3297 (N_3297,N_2963,N_2914);
nor U3298 (N_3298,N_2517,N_2534);
or U3299 (N_3299,N_2750,N_2587);
and U3300 (N_3300,N_2975,N_2996);
or U3301 (N_3301,N_2752,N_2556);
and U3302 (N_3302,N_2774,N_2849);
nand U3303 (N_3303,N_2820,N_2832);
nor U3304 (N_3304,N_2547,N_2934);
and U3305 (N_3305,N_2638,N_2897);
or U3306 (N_3306,N_2771,N_2994);
or U3307 (N_3307,N_2645,N_2878);
nor U3308 (N_3308,N_2885,N_2891);
or U3309 (N_3309,N_2699,N_2579);
or U3310 (N_3310,N_2817,N_2620);
and U3311 (N_3311,N_2749,N_2947);
nor U3312 (N_3312,N_2973,N_2914);
nor U3313 (N_3313,N_2788,N_2875);
and U3314 (N_3314,N_2633,N_2898);
and U3315 (N_3315,N_2881,N_2589);
nand U3316 (N_3316,N_2578,N_2777);
nand U3317 (N_3317,N_2933,N_2888);
xor U3318 (N_3318,N_2575,N_2760);
nand U3319 (N_3319,N_2741,N_2951);
and U3320 (N_3320,N_2513,N_2933);
nand U3321 (N_3321,N_2818,N_2516);
nand U3322 (N_3322,N_2913,N_2581);
xnor U3323 (N_3323,N_2848,N_2655);
nand U3324 (N_3324,N_2765,N_2885);
or U3325 (N_3325,N_2992,N_2538);
nand U3326 (N_3326,N_2682,N_2800);
nor U3327 (N_3327,N_2959,N_2929);
and U3328 (N_3328,N_2968,N_2793);
and U3329 (N_3329,N_2967,N_2524);
and U3330 (N_3330,N_2576,N_2532);
or U3331 (N_3331,N_2864,N_2600);
nor U3332 (N_3332,N_2582,N_2971);
nor U3333 (N_3333,N_2907,N_2611);
nand U3334 (N_3334,N_2949,N_2887);
xnor U3335 (N_3335,N_2647,N_2914);
nor U3336 (N_3336,N_2763,N_2754);
and U3337 (N_3337,N_2673,N_2722);
xor U3338 (N_3338,N_2534,N_2869);
nor U3339 (N_3339,N_2668,N_2821);
or U3340 (N_3340,N_2808,N_2610);
nand U3341 (N_3341,N_2524,N_2535);
nand U3342 (N_3342,N_2982,N_2719);
nor U3343 (N_3343,N_2615,N_2963);
nor U3344 (N_3344,N_2681,N_2556);
and U3345 (N_3345,N_2972,N_2747);
nor U3346 (N_3346,N_2805,N_2765);
or U3347 (N_3347,N_2863,N_2929);
or U3348 (N_3348,N_2559,N_2509);
nor U3349 (N_3349,N_2928,N_2632);
xnor U3350 (N_3350,N_2578,N_2645);
or U3351 (N_3351,N_2672,N_2744);
nor U3352 (N_3352,N_2687,N_2501);
nor U3353 (N_3353,N_2514,N_2658);
or U3354 (N_3354,N_2783,N_2871);
or U3355 (N_3355,N_2788,N_2865);
or U3356 (N_3356,N_2511,N_2589);
or U3357 (N_3357,N_2560,N_2621);
and U3358 (N_3358,N_2520,N_2882);
nand U3359 (N_3359,N_2798,N_2552);
or U3360 (N_3360,N_2716,N_2678);
or U3361 (N_3361,N_2740,N_2572);
nor U3362 (N_3362,N_2561,N_2957);
xor U3363 (N_3363,N_2876,N_2675);
nor U3364 (N_3364,N_2703,N_2648);
or U3365 (N_3365,N_2664,N_2830);
or U3366 (N_3366,N_2926,N_2734);
or U3367 (N_3367,N_2874,N_2935);
or U3368 (N_3368,N_2889,N_2766);
xnor U3369 (N_3369,N_2534,N_2982);
nand U3370 (N_3370,N_2792,N_2838);
nand U3371 (N_3371,N_2978,N_2881);
or U3372 (N_3372,N_2970,N_2989);
and U3373 (N_3373,N_2885,N_2868);
and U3374 (N_3374,N_2907,N_2945);
nand U3375 (N_3375,N_2567,N_2665);
xnor U3376 (N_3376,N_2549,N_2670);
or U3377 (N_3377,N_2617,N_2706);
xnor U3378 (N_3378,N_2597,N_2852);
nor U3379 (N_3379,N_2729,N_2979);
nand U3380 (N_3380,N_2544,N_2542);
nor U3381 (N_3381,N_2831,N_2792);
or U3382 (N_3382,N_2501,N_2505);
or U3383 (N_3383,N_2799,N_2702);
nand U3384 (N_3384,N_2615,N_2868);
and U3385 (N_3385,N_2883,N_2669);
xor U3386 (N_3386,N_2501,N_2697);
and U3387 (N_3387,N_2997,N_2779);
and U3388 (N_3388,N_2588,N_2537);
nor U3389 (N_3389,N_2632,N_2655);
nand U3390 (N_3390,N_2615,N_2772);
and U3391 (N_3391,N_2605,N_2880);
and U3392 (N_3392,N_2630,N_2682);
nand U3393 (N_3393,N_2630,N_2587);
xnor U3394 (N_3394,N_2709,N_2645);
nand U3395 (N_3395,N_2714,N_2835);
nand U3396 (N_3396,N_2537,N_2711);
nor U3397 (N_3397,N_2823,N_2837);
nor U3398 (N_3398,N_2737,N_2944);
and U3399 (N_3399,N_2722,N_2552);
nand U3400 (N_3400,N_2642,N_2527);
nand U3401 (N_3401,N_2701,N_2980);
nand U3402 (N_3402,N_2649,N_2989);
nor U3403 (N_3403,N_2651,N_2951);
nand U3404 (N_3404,N_2745,N_2904);
or U3405 (N_3405,N_2982,N_2554);
or U3406 (N_3406,N_2760,N_2875);
or U3407 (N_3407,N_2840,N_2733);
or U3408 (N_3408,N_2732,N_2594);
nor U3409 (N_3409,N_2769,N_2694);
or U3410 (N_3410,N_2886,N_2983);
nor U3411 (N_3411,N_2548,N_2852);
nand U3412 (N_3412,N_2611,N_2647);
nor U3413 (N_3413,N_2685,N_2957);
nand U3414 (N_3414,N_2988,N_2918);
nand U3415 (N_3415,N_2886,N_2911);
xor U3416 (N_3416,N_2944,N_2545);
or U3417 (N_3417,N_2811,N_2515);
or U3418 (N_3418,N_2804,N_2754);
and U3419 (N_3419,N_2644,N_2695);
nor U3420 (N_3420,N_2989,N_2566);
nand U3421 (N_3421,N_2505,N_2996);
xnor U3422 (N_3422,N_2973,N_2565);
and U3423 (N_3423,N_2785,N_2992);
nor U3424 (N_3424,N_2590,N_2606);
nand U3425 (N_3425,N_2611,N_2749);
nand U3426 (N_3426,N_2898,N_2650);
or U3427 (N_3427,N_2919,N_2674);
or U3428 (N_3428,N_2624,N_2570);
nor U3429 (N_3429,N_2881,N_2639);
or U3430 (N_3430,N_2734,N_2739);
or U3431 (N_3431,N_2525,N_2830);
nor U3432 (N_3432,N_2562,N_2701);
nor U3433 (N_3433,N_2590,N_2545);
nor U3434 (N_3434,N_2805,N_2524);
xnor U3435 (N_3435,N_2910,N_2926);
xor U3436 (N_3436,N_2982,N_2800);
and U3437 (N_3437,N_2501,N_2973);
xor U3438 (N_3438,N_2745,N_2972);
or U3439 (N_3439,N_2848,N_2790);
nor U3440 (N_3440,N_2781,N_2665);
and U3441 (N_3441,N_2591,N_2820);
nand U3442 (N_3442,N_2562,N_2708);
nand U3443 (N_3443,N_2784,N_2525);
nor U3444 (N_3444,N_2849,N_2626);
or U3445 (N_3445,N_2551,N_2966);
and U3446 (N_3446,N_2808,N_2920);
xnor U3447 (N_3447,N_2567,N_2716);
nand U3448 (N_3448,N_2809,N_2904);
xnor U3449 (N_3449,N_2656,N_2831);
nand U3450 (N_3450,N_2865,N_2612);
and U3451 (N_3451,N_2971,N_2853);
nor U3452 (N_3452,N_2944,N_2897);
or U3453 (N_3453,N_2700,N_2651);
nor U3454 (N_3454,N_2735,N_2847);
nor U3455 (N_3455,N_2526,N_2846);
nand U3456 (N_3456,N_2585,N_2946);
nand U3457 (N_3457,N_2781,N_2847);
or U3458 (N_3458,N_2766,N_2560);
and U3459 (N_3459,N_2917,N_2739);
nand U3460 (N_3460,N_2936,N_2874);
xor U3461 (N_3461,N_2825,N_2962);
xor U3462 (N_3462,N_2723,N_2951);
or U3463 (N_3463,N_2675,N_2575);
and U3464 (N_3464,N_2568,N_2776);
nor U3465 (N_3465,N_2750,N_2814);
nand U3466 (N_3466,N_2859,N_2799);
nor U3467 (N_3467,N_2658,N_2823);
nand U3468 (N_3468,N_2997,N_2811);
or U3469 (N_3469,N_2546,N_2916);
and U3470 (N_3470,N_2566,N_2929);
or U3471 (N_3471,N_2737,N_2631);
and U3472 (N_3472,N_2862,N_2623);
or U3473 (N_3473,N_2507,N_2891);
xor U3474 (N_3474,N_2624,N_2851);
or U3475 (N_3475,N_2648,N_2858);
nor U3476 (N_3476,N_2638,N_2560);
nor U3477 (N_3477,N_2632,N_2686);
nand U3478 (N_3478,N_2992,N_2818);
nand U3479 (N_3479,N_2501,N_2764);
or U3480 (N_3480,N_2664,N_2605);
nor U3481 (N_3481,N_2949,N_2839);
xnor U3482 (N_3482,N_2672,N_2736);
or U3483 (N_3483,N_2511,N_2866);
and U3484 (N_3484,N_2762,N_2706);
nor U3485 (N_3485,N_2628,N_2816);
nor U3486 (N_3486,N_2856,N_2726);
and U3487 (N_3487,N_2544,N_2593);
nor U3488 (N_3488,N_2788,N_2529);
nor U3489 (N_3489,N_2744,N_2958);
or U3490 (N_3490,N_2530,N_2611);
and U3491 (N_3491,N_2980,N_2800);
and U3492 (N_3492,N_2776,N_2904);
or U3493 (N_3493,N_2698,N_2737);
or U3494 (N_3494,N_2827,N_2667);
or U3495 (N_3495,N_2857,N_2609);
nand U3496 (N_3496,N_2736,N_2968);
or U3497 (N_3497,N_2962,N_2779);
or U3498 (N_3498,N_2628,N_2637);
nand U3499 (N_3499,N_2885,N_2860);
nor U3500 (N_3500,N_3111,N_3356);
or U3501 (N_3501,N_3087,N_3128);
and U3502 (N_3502,N_3306,N_3251);
and U3503 (N_3503,N_3149,N_3463);
nor U3504 (N_3504,N_3475,N_3345);
nor U3505 (N_3505,N_3190,N_3252);
and U3506 (N_3506,N_3127,N_3227);
or U3507 (N_3507,N_3214,N_3407);
nor U3508 (N_3508,N_3109,N_3362);
nand U3509 (N_3509,N_3402,N_3084);
nand U3510 (N_3510,N_3361,N_3279);
and U3511 (N_3511,N_3060,N_3488);
and U3512 (N_3512,N_3468,N_3273);
nand U3513 (N_3513,N_3492,N_3004);
xnor U3514 (N_3514,N_3496,N_3184);
and U3515 (N_3515,N_3470,N_3116);
xor U3516 (N_3516,N_3079,N_3048);
or U3517 (N_3517,N_3151,N_3082);
or U3518 (N_3518,N_3017,N_3158);
and U3519 (N_3519,N_3283,N_3040);
nor U3520 (N_3520,N_3423,N_3276);
nor U3521 (N_3521,N_3363,N_3066);
or U3522 (N_3522,N_3051,N_3445);
and U3523 (N_3523,N_3118,N_3350);
or U3524 (N_3524,N_3406,N_3333);
and U3525 (N_3525,N_3249,N_3254);
nor U3526 (N_3526,N_3392,N_3412);
nand U3527 (N_3527,N_3153,N_3452);
xor U3528 (N_3528,N_3381,N_3141);
nor U3529 (N_3529,N_3059,N_3437);
or U3530 (N_3530,N_3255,N_3372);
nand U3531 (N_3531,N_3162,N_3358);
or U3532 (N_3532,N_3387,N_3253);
and U3533 (N_3533,N_3164,N_3005);
and U3534 (N_3534,N_3009,N_3172);
nor U3535 (N_3535,N_3404,N_3025);
and U3536 (N_3536,N_3043,N_3115);
or U3537 (N_3537,N_3335,N_3261);
or U3538 (N_3538,N_3069,N_3444);
xor U3539 (N_3539,N_3319,N_3143);
or U3540 (N_3540,N_3070,N_3435);
nor U3541 (N_3541,N_3110,N_3411);
or U3542 (N_3542,N_3352,N_3077);
or U3543 (N_3543,N_3310,N_3133);
or U3544 (N_3544,N_3303,N_3467);
nor U3545 (N_3545,N_3036,N_3289);
and U3546 (N_3546,N_3293,N_3349);
or U3547 (N_3547,N_3135,N_3486);
or U3548 (N_3548,N_3003,N_3055);
nor U3549 (N_3549,N_3046,N_3420);
nand U3550 (N_3550,N_3068,N_3298);
or U3551 (N_3551,N_3365,N_3232);
nand U3552 (N_3552,N_3426,N_3160);
and U3553 (N_3553,N_3478,N_3413);
nand U3554 (N_3554,N_3489,N_3086);
and U3555 (N_3555,N_3176,N_3091);
and U3556 (N_3556,N_3099,N_3250);
nand U3557 (N_3557,N_3330,N_3321);
or U3558 (N_3558,N_3130,N_3433);
nand U3559 (N_3559,N_3331,N_3481);
or U3560 (N_3560,N_3295,N_3037);
and U3561 (N_3561,N_3226,N_3285);
nor U3562 (N_3562,N_3028,N_3113);
nor U3563 (N_3563,N_3181,N_3014);
and U3564 (N_3564,N_3373,N_3117);
or U3565 (N_3565,N_3067,N_3241);
nor U3566 (N_3566,N_3390,N_3104);
and U3567 (N_3567,N_3459,N_3403);
nand U3568 (N_3568,N_3409,N_3171);
nand U3569 (N_3569,N_3204,N_3443);
or U3570 (N_3570,N_3428,N_3073);
or U3571 (N_3571,N_3148,N_3192);
nor U3572 (N_3572,N_3446,N_3047);
nand U3573 (N_3573,N_3175,N_3200);
nand U3574 (N_3574,N_3439,N_3379);
xor U3575 (N_3575,N_3262,N_3026);
nand U3576 (N_3576,N_3215,N_3399);
or U3577 (N_3577,N_3105,N_3274);
and U3578 (N_3578,N_3264,N_3022);
and U3579 (N_3579,N_3245,N_3377);
nor U3580 (N_3580,N_3023,N_3010);
or U3581 (N_3581,N_3041,N_3346);
or U3582 (N_3582,N_3202,N_3242);
nor U3583 (N_3583,N_3355,N_3485);
nor U3584 (N_3584,N_3370,N_3369);
nand U3585 (N_3585,N_3178,N_3267);
xnor U3586 (N_3586,N_3271,N_3498);
nor U3587 (N_3587,N_3353,N_3326);
or U3588 (N_3588,N_3366,N_3432);
nand U3589 (N_3589,N_3132,N_3357);
or U3590 (N_3590,N_3400,N_3367);
and U3591 (N_3591,N_3035,N_3278);
nor U3592 (N_3592,N_3454,N_3228);
and U3593 (N_3593,N_3324,N_3163);
or U3594 (N_3594,N_3287,N_3016);
nand U3595 (N_3595,N_3179,N_3134);
nand U3596 (N_3596,N_3462,N_3374);
and U3597 (N_3597,N_3000,N_3029);
nor U3598 (N_3598,N_3408,N_3418);
nand U3599 (N_3599,N_3425,N_3229);
and U3600 (N_3600,N_3081,N_3263);
or U3601 (N_3601,N_3123,N_3144);
nor U3602 (N_3602,N_3429,N_3477);
and U3603 (N_3603,N_3193,N_3182);
nand U3604 (N_3604,N_3211,N_3024);
nor U3605 (N_3605,N_3210,N_3302);
nand U3606 (N_3606,N_3157,N_3385);
and U3607 (N_3607,N_3329,N_3054);
nor U3608 (N_3608,N_3398,N_3347);
nand U3609 (N_3609,N_3368,N_3327);
xnor U3610 (N_3610,N_3339,N_3001);
nor U3611 (N_3611,N_3042,N_3436);
xnor U3612 (N_3612,N_3240,N_3033);
or U3613 (N_3613,N_3480,N_3378);
or U3614 (N_3614,N_3225,N_3032);
nor U3615 (N_3615,N_3038,N_3216);
xor U3616 (N_3616,N_3447,N_3108);
nand U3617 (N_3617,N_3019,N_3057);
nor U3618 (N_3618,N_3020,N_3266);
nor U3619 (N_3619,N_3300,N_3259);
nand U3620 (N_3620,N_3102,N_3138);
nand U3621 (N_3621,N_3119,N_3464);
nand U3622 (N_3622,N_3056,N_3191);
nor U3623 (N_3623,N_3395,N_3169);
xor U3624 (N_3624,N_3247,N_3383);
or U3625 (N_3625,N_3305,N_3196);
nor U3626 (N_3626,N_3317,N_3071);
and U3627 (N_3627,N_3074,N_3294);
and U3628 (N_3628,N_3313,N_3297);
and U3629 (N_3629,N_3183,N_3018);
and U3630 (N_3630,N_3301,N_3320);
or U3631 (N_3631,N_3382,N_3461);
nor U3632 (N_3632,N_3323,N_3061);
nand U3633 (N_3633,N_3002,N_3277);
and U3634 (N_3634,N_3417,N_3465);
xnor U3635 (N_3635,N_3364,N_3044);
nor U3636 (N_3636,N_3248,N_3224);
or U3637 (N_3637,N_3188,N_3282);
nand U3638 (N_3638,N_3236,N_3474);
nor U3639 (N_3639,N_3159,N_3337);
and U3640 (N_3640,N_3451,N_3058);
nor U3641 (N_3641,N_3471,N_3286);
xnor U3642 (N_3642,N_3490,N_3371);
nand U3643 (N_3643,N_3410,N_3456);
xnor U3644 (N_3644,N_3007,N_3063);
nor U3645 (N_3645,N_3415,N_3360);
and U3646 (N_3646,N_3075,N_3209);
nor U3647 (N_3647,N_3220,N_3006);
or U3648 (N_3648,N_3348,N_3422);
and U3649 (N_3649,N_3483,N_3013);
nand U3650 (N_3650,N_3299,N_3218);
nand U3651 (N_3651,N_3328,N_3389);
nor U3652 (N_3652,N_3342,N_3097);
nand U3653 (N_3653,N_3343,N_3140);
nor U3654 (N_3654,N_3185,N_3269);
or U3655 (N_3655,N_3080,N_3137);
and U3656 (N_3656,N_3212,N_3491);
nand U3657 (N_3657,N_3206,N_3290);
nor U3658 (N_3658,N_3431,N_3053);
nor U3659 (N_3659,N_3416,N_3309);
nand U3660 (N_3660,N_3325,N_3499);
or U3661 (N_3661,N_3136,N_3351);
nor U3662 (N_3662,N_3145,N_3114);
or U3663 (N_3663,N_3161,N_3093);
nand U3664 (N_3664,N_3275,N_3238);
nand U3665 (N_3665,N_3394,N_3405);
xnor U3666 (N_3666,N_3072,N_3450);
nand U3667 (N_3667,N_3334,N_3341);
and U3668 (N_3668,N_3376,N_3095);
and U3669 (N_3669,N_3222,N_3121);
nand U3670 (N_3670,N_3235,N_3270);
nor U3671 (N_3671,N_3106,N_3064);
xor U3672 (N_3672,N_3280,N_3272);
and U3673 (N_3673,N_3170,N_3479);
or U3674 (N_3674,N_3312,N_3089);
nand U3675 (N_3675,N_3388,N_3112);
nor U3676 (N_3676,N_3015,N_3090);
or U3677 (N_3677,N_3239,N_3186);
nor U3678 (N_3678,N_3472,N_3180);
or U3679 (N_3679,N_3421,N_3484);
or U3680 (N_3680,N_3344,N_3078);
and U3681 (N_3681,N_3187,N_3438);
nor U3682 (N_3682,N_3125,N_3354);
nand U3683 (N_3683,N_3195,N_3156);
or U3684 (N_3684,N_3213,N_3049);
nor U3685 (N_3685,N_3359,N_3223);
nand U3686 (N_3686,N_3167,N_3307);
and U3687 (N_3687,N_3434,N_3011);
and U3688 (N_3688,N_3268,N_3197);
and U3689 (N_3689,N_3101,N_3281);
or U3690 (N_3690,N_3174,N_3457);
and U3691 (N_3691,N_3386,N_3460);
or U3692 (N_3692,N_3065,N_3031);
nand U3693 (N_3693,N_3414,N_3221);
and U3694 (N_3694,N_3311,N_3316);
nand U3695 (N_3695,N_3401,N_3217);
nor U3696 (N_3696,N_3194,N_3233);
nor U3697 (N_3697,N_3008,N_3393);
nor U3698 (N_3698,N_3256,N_3494);
nand U3699 (N_3699,N_3139,N_3050);
and U3700 (N_3700,N_3476,N_3304);
nor U3701 (N_3701,N_3427,N_3384);
nor U3702 (N_3702,N_3497,N_3288);
nand U3703 (N_3703,N_3315,N_3201);
xor U3704 (N_3704,N_3482,N_3495);
and U3705 (N_3705,N_3487,N_3203);
or U3706 (N_3706,N_3430,N_3338);
nor U3707 (N_3707,N_3088,N_3098);
and U3708 (N_3708,N_3292,N_3375);
and U3709 (N_3709,N_3096,N_3230);
or U3710 (N_3710,N_3092,N_3314);
nand U3711 (N_3711,N_3308,N_3246);
nand U3712 (N_3712,N_3126,N_3473);
or U3713 (N_3713,N_3419,N_3142);
nor U3714 (N_3714,N_3244,N_3103);
and U3715 (N_3715,N_3257,N_3094);
and U3716 (N_3716,N_3397,N_3030);
xor U3717 (N_3717,N_3458,N_3340);
and U3718 (N_3718,N_3318,N_3012);
and U3719 (N_3719,N_3155,N_3243);
nor U3720 (N_3720,N_3493,N_3062);
nand U3721 (N_3721,N_3219,N_3083);
nor U3722 (N_3722,N_3168,N_3469);
xor U3723 (N_3723,N_3189,N_3147);
and U3724 (N_3724,N_3296,N_3124);
xor U3725 (N_3725,N_3258,N_3039);
nand U3726 (N_3726,N_3284,N_3122);
or U3727 (N_3727,N_3332,N_3231);
xnor U3728 (N_3728,N_3146,N_3199);
or U3729 (N_3729,N_3260,N_3455);
nand U3730 (N_3730,N_3391,N_3205);
nand U3731 (N_3731,N_3322,N_3234);
xor U3732 (N_3732,N_3152,N_3449);
nor U3733 (N_3733,N_3208,N_3336);
nor U3734 (N_3734,N_3396,N_3165);
nor U3735 (N_3735,N_3027,N_3265);
nor U3736 (N_3736,N_3466,N_3150);
nor U3737 (N_3737,N_3052,N_3424);
nand U3738 (N_3738,N_3166,N_3173);
and U3739 (N_3739,N_3100,N_3380);
or U3740 (N_3740,N_3237,N_3076);
and U3741 (N_3741,N_3045,N_3291);
and U3742 (N_3742,N_3085,N_3442);
and U3743 (N_3743,N_3198,N_3448);
and U3744 (N_3744,N_3453,N_3207);
nand U3745 (N_3745,N_3154,N_3441);
xnor U3746 (N_3746,N_3120,N_3129);
nand U3747 (N_3747,N_3440,N_3034);
xnor U3748 (N_3748,N_3021,N_3107);
and U3749 (N_3749,N_3177,N_3131);
and U3750 (N_3750,N_3213,N_3333);
nand U3751 (N_3751,N_3057,N_3422);
nor U3752 (N_3752,N_3251,N_3490);
or U3753 (N_3753,N_3168,N_3106);
xor U3754 (N_3754,N_3124,N_3279);
nor U3755 (N_3755,N_3300,N_3349);
nor U3756 (N_3756,N_3301,N_3447);
nand U3757 (N_3757,N_3352,N_3280);
and U3758 (N_3758,N_3491,N_3107);
or U3759 (N_3759,N_3456,N_3176);
or U3760 (N_3760,N_3124,N_3302);
nand U3761 (N_3761,N_3126,N_3133);
nor U3762 (N_3762,N_3436,N_3010);
xnor U3763 (N_3763,N_3371,N_3416);
and U3764 (N_3764,N_3214,N_3223);
and U3765 (N_3765,N_3383,N_3326);
nand U3766 (N_3766,N_3228,N_3262);
nor U3767 (N_3767,N_3048,N_3465);
or U3768 (N_3768,N_3478,N_3415);
or U3769 (N_3769,N_3108,N_3023);
xnor U3770 (N_3770,N_3280,N_3285);
and U3771 (N_3771,N_3004,N_3170);
nor U3772 (N_3772,N_3322,N_3461);
xnor U3773 (N_3773,N_3171,N_3035);
nor U3774 (N_3774,N_3159,N_3275);
xor U3775 (N_3775,N_3150,N_3400);
or U3776 (N_3776,N_3420,N_3306);
nor U3777 (N_3777,N_3167,N_3432);
nand U3778 (N_3778,N_3070,N_3062);
and U3779 (N_3779,N_3124,N_3301);
or U3780 (N_3780,N_3483,N_3023);
nor U3781 (N_3781,N_3154,N_3194);
or U3782 (N_3782,N_3348,N_3098);
and U3783 (N_3783,N_3347,N_3154);
nor U3784 (N_3784,N_3322,N_3326);
nand U3785 (N_3785,N_3453,N_3222);
nand U3786 (N_3786,N_3489,N_3267);
nor U3787 (N_3787,N_3227,N_3263);
nand U3788 (N_3788,N_3082,N_3044);
and U3789 (N_3789,N_3386,N_3354);
or U3790 (N_3790,N_3419,N_3041);
and U3791 (N_3791,N_3096,N_3249);
or U3792 (N_3792,N_3216,N_3199);
xor U3793 (N_3793,N_3390,N_3132);
and U3794 (N_3794,N_3245,N_3209);
nand U3795 (N_3795,N_3115,N_3145);
nand U3796 (N_3796,N_3445,N_3334);
nand U3797 (N_3797,N_3113,N_3309);
nor U3798 (N_3798,N_3223,N_3405);
xnor U3799 (N_3799,N_3362,N_3170);
nand U3800 (N_3800,N_3489,N_3288);
or U3801 (N_3801,N_3362,N_3452);
nor U3802 (N_3802,N_3344,N_3002);
xnor U3803 (N_3803,N_3156,N_3094);
nor U3804 (N_3804,N_3348,N_3424);
and U3805 (N_3805,N_3370,N_3130);
nand U3806 (N_3806,N_3417,N_3082);
and U3807 (N_3807,N_3126,N_3391);
or U3808 (N_3808,N_3163,N_3229);
and U3809 (N_3809,N_3262,N_3055);
or U3810 (N_3810,N_3204,N_3138);
or U3811 (N_3811,N_3220,N_3089);
nand U3812 (N_3812,N_3260,N_3200);
nor U3813 (N_3813,N_3001,N_3109);
nand U3814 (N_3814,N_3267,N_3191);
and U3815 (N_3815,N_3440,N_3156);
nand U3816 (N_3816,N_3229,N_3170);
or U3817 (N_3817,N_3134,N_3315);
xor U3818 (N_3818,N_3179,N_3383);
nor U3819 (N_3819,N_3128,N_3313);
nand U3820 (N_3820,N_3237,N_3252);
nor U3821 (N_3821,N_3406,N_3079);
and U3822 (N_3822,N_3229,N_3349);
nand U3823 (N_3823,N_3037,N_3370);
nor U3824 (N_3824,N_3451,N_3230);
and U3825 (N_3825,N_3488,N_3256);
and U3826 (N_3826,N_3284,N_3400);
nand U3827 (N_3827,N_3371,N_3193);
nand U3828 (N_3828,N_3078,N_3197);
nor U3829 (N_3829,N_3305,N_3473);
or U3830 (N_3830,N_3038,N_3067);
and U3831 (N_3831,N_3183,N_3055);
nand U3832 (N_3832,N_3450,N_3319);
nor U3833 (N_3833,N_3209,N_3298);
nand U3834 (N_3834,N_3126,N_3100);
and U3835 (N_3835,N_3384,N_3232);
and U3836 (N_3836,N_3205,N_3021);
xnor U3837 (N_3837,N_3421,N_3473);
nand U3838 (N_3838,N_3000,N_3094);
nor U3839 (N_3839,N_3138,N_3164);
nor U3840 (N_3840,N_3439,N_3214);
xor U3841 (N_3841,N_3196,N_3415);
or U3842 (N_3842,N_3348,N_3272);
nand U3843 (N_3843,N_3446,N_3172);
nor U3844 (N_3844,N_3391,N_3079);
nor U3845 (N_3845,N_3204,N_3221);
nand U3846 (N_3846,N_3365,N_3192);
and U3847 (N_3847,N_3008,N_3048);
or U3848 (N_3848,N_3176,N_3432);
and U3849 (N_3849,N_3198,N_3256);
and U3850 (N_3850,N_3341,N_3076);
or U3851 (N_3851,N_3448,N_3271);
and U3852 (N_3852,N_3411,N_3492);
nand U3853 (N_3853,N_3051,N_3208);
and U3854 (N_3854,N_3331,N_3171);
and U3855 (N_3855,N_3141,N_3397);
or U3856 (N_3856,N_3472,N_3247);
and U3857 (N_3857,N_3138,N_3016);
and U3858 (N_3858,N_3475,N_3224);
nor U3859 (N_3859,N_3413,N_3260);
or U3860 (N_3860,N_3460,N_3378);
and U3861 (N_3861,N_3403,N_3179);
nand U3862 (N_3862,N_3410,N_3050);
and U3863 (N_3863,N_3413,N_3447);
nor U3864 (N_3864,N_3155,N_3249);
xor U3865 (N_3865,N_3451,N_3357);
nand U3866 (N_3866,N_3403,N_3251);
nand U3867 (N_3867,N_3407,N_3196);
or U3868 (N_3868,N_3260,N_3188);
xnor U3869 (N_3869,N_3192,N_3106);
nor U3870 (N_3870,N_3046,N_3066);
nor U3871 (N_3871,N_3008,N_3481);
and U3872 (N_3872,N_3285,N_3033);
or U3873 (N_3873,N_3099,N_3123);
nor U3874 (N_3874,N_3402,N_3028);
xnor U3875 (N_3875,N_3199,N_3247);
and U3876 (N_3876,N_3475,N_3283);
nor U3877 (N_3877,N_3154,N_3111);
or U3878 (N_3878,N_3135,N_3441);
nor U3879 (N_3879,N_3369,N_3423);
nand U3880 (N_3880,N_3247,N_3208);
xor U3881 (N_3881,N_3089,N_3131);
or U3882 (N_3882,N_3113,N_3234);
nor U3883 (N_3883,N_3073,N_3446);
and U3884 (N_3884,N_3307,N_3422);
and U3885 (N_3885,N_3169,N_3083);
nor U3886 (N_3886,N_3325,N_3223);
and U3887 (N_3887,N_3247,N_3481);
and U3888 (N_3888,N_3207,N_3337);
or U3889 (N_3889,N_3369,N_3032);
xor U3890 (N_3890,N_3484,N_3156);
nor U3891 (N_3891,N_3015,N_3138);
nor U3892 (N_3892,N_3442,N_3099);
nor U3893 (N_3893,N_3181,N_3190);
nor U3894 (N_3894,N_3139,N_3200);
xor U3895 (N_3895,N_3193,N_3221);
or U3896 (N_3896,N_3439,N_3384);
and U3897 (N_3897,N_3097,N_3323);
nor U3898 (N_3898,N_3391,N_3359);
nand U3899 (N_3899,N_3182,N_3090);
nor U3900 (N_3900,N_3434,N_3393);
nand U3901 (N_3901,N_3395,N_3195);
nor U3902 (N_3902,N_3170,N_3038);
or U3903 (N_3903,N_3395,N_3025);
nand U3904 (N_3904,N_3119,N_3218);
xor U3905 (N_3905,N_3338,N_3040);
xor U3906 (N_3906,N_3146,N_3071);
nor U3907 (N_3907,N_3187,N_3321);
nor U3908 (N_3908,N_3301,N_3250);
or U3909 (N_3909,N_3219,N_3265);
or U3910 (N_3910,N_3011,N_3273);
and U3911 (N_3911,N_3214,N_3321);
nand U3912 (N_3912,N_3011,N_3237);
nor U3913 (N_3913,N_3005,N_3077);
and U3914 (N_3914,N_3005,N_3325);
and U3915 (N_3915,N_3463,N_3168);
and U3916 (N_3916,N_3222,N_3473);
nor U3917 (N_3917,N_3013,N_3352);
or U3918 (N_3918,N_3188,N_3003);
nor U3919 (N_3919,N_3336,N_3039);
or U3920 (N_3920,N_3428,N_3450);
and U3921 (N_3921,N_3012,N_3404);
nand U3922 (N_3922,N_3232,N_3233);
or U3923 (N_3923,N_3402,N_3409);
xnor U3924 (N_3924,N_3099,N_3487);
and U3925 (N_3925,N_3061,N_3395);
or U3926 (N_3926,N_3030,N_3292);
nand U3927 (N_3927,N_3059,N_3228);
nor U3928 (N_3928,N_3062,N_3144);
or U3929 (N_3929,N_3186,N_3281);
or U3930 (N_3930,N_3090,N_3173);
nor U3931 (N_3931,N_3019,N_3481);
nand U3932 (N_3932,N_3111,N_3296);
or U3933 (N_3933,N_3090,N_3097);
nor U3934 (N_3934,N_3248,N_3210);
nor U3935 (N_3935,N_3222,N_3366);
and U3936 (N_3936,N_3253,N_3279);
and U3937 (N_3937,N_3031,N_3168);
or U3938 (N_3938,N_3229,N_3458);
xor U3939 (N_3939,N_3389,N_3441);
nand U3940 (N_3940,N_3377,N_3215);
nand U3941 (N_3941,N_3489,N_3468);
nand U3942 (N_3942,N_3260,N_3010);
or U3943 (N_3943,N_3397,N_3127);
or U3944 (N_3944,N_3427,N_3235);
or U3945 (N_3945,N_3457,N_3144);
nor U3946 (N_3946,N_3390,N_3090);
or U3947 (N_3947,N_3043,N_3063);
nand U3948 (N_3948,N_3117,N_3279);
nand U3949 (N_3949,N_3473,N_3175);
and U3950 (N_3950,N_3265,N_3482);
or U3951 (N_3951,N_3263,N_3495);
nand U3952 (N_3952,N_3226,N_3412);
nand U3953 (N_3953,N_3478,N_3410);
nand U3954 (N_3954,N_3496,N_3403);
xnor U3955 (N_3955,N_3002,N_3252);
nor U3956 (N_3956,N_3360,N_3333);
and U3957 (N_3957,N_3301,N_3309);
nor U3958 (N_3958,N_3017,N_3422);
nor U3959 (N_3959,N_3475,N_3472);
nor U3960 (N_3960,N_3212,N_3338);
and U3961 (N_3961,N_3094,N_3192);
nand U3962 (N_3962,N_3168,N_3468);
nor U3963 (N_3963,N_3397,N_3472);
nand U3964 (N_3964,N_3151,N_3052);
and U3965 (N_3965,N_3130,N_3188);
or U3966 (N_3966,N_3012,N_3067);
nor U3967 (N_3967,N_3076,N_3425);
or U3968 (N_3968,N_3311,N_3457);
or U3969 (N_3969,N_3427,N_3480);
nand U3970 (N_3970,N_3276,N_3151);
nand U3971 (N_3971,N_3411,N_3142);
or U3972 (N_3972,N_3264,N_3054);
nand U3973 (N_3973,N_3074,N_3336);
nor U3974 (N_3974,N_3316,N_3324);
or U3975 (N_3975,N_3368,N_3261);
xor U3976 (N_3976,N_3194,N_3048);
xnor U3977 (N_3977,N_3134,N_3252);
and U3978 (N_3978,N_3208,N_3390);
or U3979 (N_3979,N_3113,N_3066);
and U3980 (N_3980,N_3474,N_3190);
nand U3981 (N_3981,N_3295,N_3221);
xor U3982 (N_3982,N_3391,N_3265);
nor U3983 (N_3983,N_3323,N_3297);
and U3984 (N_3984,N_3266,N_3381);
xor U3985 (N_3985,N_3434,N_3051);
nand U3986 (N_3986,N_3457,N_3473);
nand U3987 (N_3987,N_3233,N_3442);
and U3988 (N_3988,N_3143,N_3069);
nand U3989 (N_3989,N_3305,N_3470);
nor U3990 (N_3990,N_3381,N_3038);
or U3991 (N_3991,N_3016,N_3279);
xor U3992 (N_3992,N_3410,N_3093);
nand U3993 (N_3993,N_3244,N_3350);
nor U3994 (N_3994,N_3470,N_3079);
nand U3995 (N_3995,N_3023,N_3172);
nand U3996 (N_3996,N_3431,N_3350);
nand U3997 (N_3997,N_3054,N_3363);
nor U3998 (N_3998,N_3048,N_3021);
or U3999 (N_3999,N_3070,N_3016);
xnor U4000 (N_4000,N_3949,N_3876);
or U4001 (N_4001,N_3581,N_3982);
nor U4002 (N_4002,N_3873,N_3723);
xor U4003 (N_4003,N_3843,N_3735);
nor U4004 (N_4004,N_3730,N_3734);
or U4005 (N_4005,N_3702,N_3961);
nand U4006 (N_4006,N_3912,N_3851);
or U4007 (N_4007,N_3819,N_3528);
and U4008 (N_4008,N_3775,N_3955);
and U4009 (N_4009,N_3750,N_3956);
nor U4010 (N_4010,N_3720,N_3579);
xor U4011 (N_4011,N_3512,N_3518);
nand U4012 (N_4012,N_3928,N_3918);
or U4013 (N_4013,N_3599,N_3810);
and U4014 (N_4014,N_3525,N_3764);
or U4015 (N_4015,N_3825,N_3954);
nor U4016 (N_4016,N_3564,N_3538);
nor U4017 (N_4017,N_3762,N_3548);
nand U4018 (N_4018,N_3753,N_3585);
or U4019 (N_4019,N_3900,N_3740);
or U4020 (N_4020,N_3914,N_3866);
xnor U4021 (N_4021,N_3526,N_3827);
nor U4022 (N_4022,N_3598,N_3771);
and U4023 (N_4023,N_3593,N_3559);
nand U4024 (N_4024,N_3539,N_3924);
nand U4025 (N_4025,N_3591,N_3976);
or U4026 (N_4026,N_3828,N_3536);
or U4027 (N_4027,N_3665,N_3765);
nand U4028 (N_4028,N_3658,N_3844);
or U4029 (N_4029,N_3670,N_3607);
or U4030 (N_4030,N_3703,N_3733);
nor U4031 (N_4031,N_3952,N_3556);
and U4032 (N_4032,N_3829,N_3576);
nor U4033 (N_4033,N_3929,N_3645);
and U4034 (N_4034,N_3690,N_3573);
nand U4035 (N_4035,N_3563,N_3784);
nor U4036 (N_4036,N_3738,N_3790);
nand U4037 (N_4037,N_3571,N_3853);
or U4038 (N_4038,N_3621,N_3562);
nor U4039 (N_4039,N_3916,N_3553);
and U4040 (N_4040,N_3502,N_3779);
and U4041 (N_4041,N_3551,N_3800);
nor U4042 (N_4042,N_3813,N_3572);
or U4043 (N_4043,N_3989,N_3904);
and U4044 (N_4044,N_3906,N_3774);
or U4045 (N_4045,N_3676,N_3991);
and U4046 (N_4046,N_3913,N_3922);
or U4047 (N_4047,N_3597,N_3641);
or U4048 (N_4048,N_3835,N_3809);
or U4049 (N_4049,N_3500,N_3729);
nor U4050 (N_4050,N_3660,N_3504);
nand U4051 (N_4051,N_3664,N_3520);
nand U4052 (N_4052,N_3944,N_3541);
nand U4053 (N_4053,N_3693,N_3637);
nor U4054 (N_4054,N_3647,N_3711);
nor U4055 (N_4055,N_3938,N_3847);
xor U4056 (N_4056,N_3725,N_3999);
or U4057 (N_4057,N_3569,N_3721);
nand U4058 (N_4058,N_3758,N_3974);
or U4059 (N_4059,N_3544,N_3656);
and U4060 (N_4060,N_3683,N_3542);
nor U4061 (N_4061,N_3950,N_3933);
nand U4062 (N_4062,N_3875,N_3507);
or U4063 (N_4063,N_3931,N_3651);
or U4064 (N_4064,N_3561,N_3659);
or U4065 (N_4065,N_3970,N_3527);
nand U4066 (N_4066,N_3503,N_3768);
and U4067 (N_4067,N_3627,N_3877);
and U4068 (N_4068,N_3617,N_3588);
and U4069 (N_4069,N_3718,N_3760);
nand U4070 (N_4070,N_3653,N_3675);
nor U4071 (N_4071,N_3977,N_3988);
and U4072 (N_4072,N_3555,N_3772);
nand U4073 (N_4073,N_3532,N_3523);
nor U4074 (N_4074,N_3602,N_3657);
or U4075 (N_4075,N_3787,N_3558);
nand U4076 (N_4076,N_3727,N_3707);
and U4077 (N_4077,N_3592,N_3742);
and U4078 (N_4078,N_3521,N_3574);
xnor U4079 (N_4079,N_3766,N_3975);
xnor U4080 (N_4080,N_3948,N_3782);
nor U4081 (N_4081,N_3698,N_3649);
or U4082 (N_4082,N_3880,N_3942);
nor U4083 (N_4083,N_3547,N_3600);
nor U4084 (N_4084,N_3717,N_3820);
nand U4085 (N_4085,N_3927,N_3613);
and U4086 (N_4086,N_3769,N_3537);
and U4087 (N_4087,N_3963,N_3508);
nor U4088 (N_4088,N_3966,N_3886);
or U4089 (N_4089,N_3728,N_3625);
nand U4090 (N_4090,N_3793,N_3618);
nand U4091 (N_4091,N_3823,N_3688);
and U4092 (N_4092,N_3752,N_3586);
and U4093 (N_4093,N_3953,N_3560);
or U4094 (N_4094,N_3650,N_3557);
or U4095 (N_4095,N_3919,N_3864);
nor U4096 (N_4096,N_3680,N_3798);
and U4097 (N_4097,N_3885,N_3980);
nand U4098 (N_4098,N_3812,N_3788);
nand U4099 (N_4099,N_3674,N_3601);
xor U4100 (N_4100,N_3856,N_3619);
or U4101 (N_4101,N_3673,N_3511);
or U4102 (N_4102,N_3892,N_3781);
or U4103 (N_4103,N_3540,N_3616);
xnor U4104 (N_4104,N_3614,N_3748);
nor U4105 (N_4105,N_3639,N_3965);
nand U4106 (N_4106,N_3794,N_3842);
and U4107 (N_4107,N_3958,N_3722);
or U4108 (N_4108,N_3979,N_3759);
nand U4109 (N_4109,N_3789,N_3524);
or U4110 (N_4110,N_3832,N_3552);
xor U4111 (N_4111,N_3749,N_3755);
nor U4112 (N_4112,N_3669,N_3509);
xor U4113 (N_4113,N_3663,N_3643);
nand U4114 (N_4114,N_3978,N_3802);
nor U4115 (N_4115,N_3939,N_3751);
nand U4116 (N_4116,N_3731,N_3681);
nor U4117 (N_4117,N_3898,N_3964);
nand U4118 (N_4118,N_3883,N_3830);
nand U4119 (N_4119,N_3887,N_3908);
nand U4120 (N_4120,N_3689,N_3902);
nor U4121 (N_4121,N_3865,N_3692);
nand U4122 (N_4122,N_3971,N_3773);
or U4123 (N_4123,N_3661,N_3807);
nand U4124 (N_4124,N_3850,N_3761);
nor U4125 (N_4125,N_3867,N_3513);
and U4126 (N_4126,N_3715,N_3917);
xor U4127 (N_4127,N_3724,N_3737);
or U4128 (N_4128,N_3567,N_3629);
and U4129 (N_4129,N_3841,N_3746);
and U4130 (N_4130,N_3947,N_3894);
and U4131 (N_4131,N_3668,N_3710);
nand U4132 (N_4132,N_3655,N_3854);
and U4133 (N_4133,N_3869,N_3652);
and U4134 (N_4134,N_3805,N_3684);
nor U4135 (N_4135,N_3691,N_3973);
and U4136 (N_4136,N_3714,N_3796);
nor U4137 (N_4137,N_3816,N_3967);
and U4138 (N_4138,N_3505,N_3905);
and U4139 (N_4139,N_3726,N_3943);
nand U4140 (N_4140,N_3682,N_3654);
and U4141 (N_4141,N_3550,N_3899);
or U4142 (N_4142,N_3837,N_3719);
nand U4143 (N_4143,N_3754,N_3662);
nor U4144 (N_4144,N_3833,N_3893);
nand U4145 (N_4145,N_3566,N_3868);
nand U4146 (N_4146,N_3695,N_3895);
xor U4147 (N_4147,N_3909,N_3612);
nor U4148 (N_4148,N_3584,N_3941);
nor U4149 (N_4149,N_3945,N_3763);
or U4150 (N_4150,N_3580,N_3845);
nor U4151 (N_4151,N_3852,N_3549);
or U4152 (N_4152,N_3926,N_3882);
or U4153 (N_4153,N_3708,N_3839);
or U4154 (N_4154,N_3596,N_3831);
or U4155 (N_4155,N_3861,N_3620);
or U4156 (N_4156,N_3879,N_3799);
xnor U4157 (N_4157,N_3777,N_3516);
nand U4158 (N_4158,N_3640,N_3935);
nand U4159 (N_4159,N_3628,N_3603);
nand U4160 (N_4160,N_3946,N_3545);
nand U4161 (N_4161,N_3756,N_3959);
and U4162 (N_4162,N_3747,N_3623);
or U4163 (N_4163,N_3815,N_3646);
or U4164 (N_4164,N_3694,N_3533);
nor U4165 (N_4165,N_3570,N_3510);
or U4166 (N_4166,N_3615,N_3677);
nor U4167 (N_4167,N_3604,N_3859);
nor U4168 (N_4168,N_3577,N_3804);
and U4169 (N_4169,N_3930,N_3817);
nand U4170 (N_4170,N_3834,N_3608);
and U4171 (N_4171,N_3872,N_3824);
nand U4172 (N_4172,N_3821,N_3811);
nand U4173 (N_4173,N_3531,N_3530);
xor U4174 (N_4174,N_3770,N_3814);
and U4175 (N_4175,N_3801,N_3934);
nand U4176 (N_4176,N_3910,N_3590);
or U4177 (N_4177,N_3960,N_3535);
nand U4178 (N_4178,N_3846,N_3757);
and U4179 (N_4179,N_3888,N_3701);
nor U4180 (N_4180,N_3632,N_3529);
or U4181 (N_4181,N_3803,N_3638);
and U4182 (N_4182,N_3672,N_3678);
and U4183 (N_4183,N_3870,N_3744);
nor U4184 (N_4184,N_3522,N_3685);
nand U4185 (N_4185,N_3626,N_3589);
xnor U4186 (N_4186,N_3915,N_3546);
and U4187 (N_4187,N_3595,N_3501);
nand U4188 (N_4188,N_3822,N_3648);
xor U4189 (N_4189,N_3587,N_3716);
nand U4190 (N_4190,N_3783,N_3786);
and U4191 (N_4191,N_3863,N_3611);
or U4192 (N_4192,N_3667,N_3514);
nor U4193 (N_4193,N_3849,N_3911);
or U4194 (N_4194,N_3986,N_3996);
or U4195 (N_4195,N_3709,N_3969);
or U4196 (N_4196,N_3679,N_3871);
and U4197 (N_4197,N_3713,N_3968);
and U4198 (N_4198,N_3994,N_3699);
and U4199 (N_4199,N_3897,N_3745);
nor U4200 (N_4200,N_3633,N_3998);
or U4201 (N_4201,N_3890,N_3700);
nand U4202 (N_4202,N_3818,N_3687);
nand U4203 (N_4203,N_3840,N_3605);
and U4204 (N_4204,N_3951,N_3889);
nor U4205 (N_4205,N_3862,N_3534);
or U4206 (N_4206,N_3568,N_3644);
nor U4207 (N_4207,N_3884,N_3920);
nand U4208 (N_4208,N_3797,N_3901);
or U4209 (N_4209,N_3878,N_3517);
and U4210 (N_4210,N_3778,N_3704);
nor U4211 (N_4211,N_3606,N_3666);
and U4212 (N_4212,N_3972,N_3506);
nor U4213 (N_4213,N_3519,N_3696);
nor U4214 (N_4214,N_3990,N_3848);
and U4215 (N_4215,N_3582,N_3780);
and U4216 (N_4216,N_3925,N_3836);
and U4217 (N_4217,N_3686,N_3860);
or U4218 (N_4218,N_3636,N_3962);
nand U4219 (N_4219,N_3808,N_3806);
nor U4220 (N_4220,N_3565,N_3543);
xnor U4221 (N_4221,N_3635,N_3515);
nor U4222 (N_4222,N_3712,N_3575);
and U4223 (N_4223,N_3743,N_3697);
nor U4224 (N_4224,N_3739,N_3983);
nor U4225 (N_4225,N_3921,N_3855);
and U4226 (N_4226,N_3630,N_3940);
or U4227 (N_4227,N_3984,N_3583);
or U4228 (N_4228,N_3671,N_3741);
nand U4229 (N_4229,N_3985,N_3858);
or U4230 (N_4230,N_3993,N_3795);
nor U4231 (N_4231,N_3874,N_3857);
or U4232 (N_4232,N_3732,N_3554);
nand U4233 (N_4233,N_3896,N_3622);
xnor U4234 (N_4234,N_3785,N_3838);
and U4235 (N_4235,N_3907,N_3776);
nor U4236 (N_4236,N_3937,N_3736);
or U4237 (N_4237,N_3903,N_3642);
nor U4238 (N_4238,N_3936,N_3624);
nand U4239 (N_4239,N_3997,N_3992);
or U4240 (N_4240,N_3705,N_3578);
and U4241 (N_4241,N_3881,N_3767);
xnor U4242 (N_4242,N_3981,N_3891);
and U4243 (N_4243,N_3957,N_3609);
xor U4244 (N_4244,N_3791,N_3610);
xnor U4245 (N_4245,N_3634,N_3594);
or U4246 (N_4246,N_3932,N_3631);
xor U4247 (N_4247,N_3923,N_3995);
nand U4248 (N_4248,N_3987,N_3706);
or U4249 (N_4249,N_3826,N_3792);
nor U4250 (N_4250,N_3731,N_3814);
nor U4251 (N_4251,N_3997,N_3553);
nand U4252 (N_4252,N_3593,N_3713);
nor U4253 (N_4253,N_3586,N_3628);
nor U4254 (N_4254,N_3743,N_3504);
or U4255 (N_4255,N_3948,N_3556);
nor U4256 (N_4256,N_3661,N_3858);
nor U4257 (N_4257,N_3659,N_3856);
or U4258 (N_4258,N_3702,N_3623);
or U4259 (N_4259,N_3976,N_3831);
and U4260 (N_4260,N_3795,N_3716);
and U4261 (N_4261,N_3571,N_3649);
and U4262 (N_4262,N_3624,N_3615);
nand U4263 (N_4263,N_3947,N_3605);
and U4264 (N_4264,N_3600,N_3818);
nand U4265 (N_4265,N_3584,N_3869);
or U4266 (N_4266,N_3543,N_3709);
and U4267 (N_4267,N_3887,N_3731);
nand U4268 (N_4268,N_3914,N_3537);
and U4269 (N_4269,N_3829,N_3676);
nand U4270 (N_4270,N_3701,N_3937);
or U4271 (N_4271,N_3767,N_3957);
nor U4272 (N_4272,N_3942,N_3790);
and U4273 (N_4273,N_3828,N_3629);
or U4274 (N_4274,N_3958,N_3577);
xnor U4275 (N_4275,N_3879,N_3536);
nor U4276 (N_4276,N_3956,N_3840);
and U4277 (N_4277,N_3873,N_3963);
nand U4278 (N_4278,N_3837,N_3911);
nand U4279 (N_4279,N_3664,N_3847);
nand U4280 (N_4280,N_3828,N_3803);
and U4281 (N_4281,N_3866,N_3634);
and U4282 (N_4282,N_3844,N_3857);
and U4283 (N_4283,N_3788,N_3830);
nor U4284 (N_4284,N_3620,N_3966);
xor U4285 (N_4285,N_3902,N_3969);
and U4286 (N_4286,N_3918,N_3516);
or U4287 (N_4287,N_3513,N_3573);
and U4288 (N_4288,N_3832,N_3757);
and U4289 (N_4289,N_3727,N_3734);
or U4290 (N_4290,N_3968,N_3707);
nand U4291 (N_4291,N_3741,N_3704);
xor U4292 (N_4292,N_3543,N_3712);
and U4293 (N_4293,N_3511,N_3655);
nor U4294 (N_4294,N_3577,N_3979);
nand U4295 (N_4295,N_3696,N_3749);
or U4296 (N_4296,N_3957,N_3763);
or U4297 (N_4297,N_3681,N_3851);
nor U4298 (N_4298,N_3945,N_3652);
nand U4299 (N_4299,N_3575,N_3871);
xnor U4300 (N_4300,N_3758,N_3943);
nor U4301 (N_4301,N_3925,N_3969);
or U4302 (N_4302,N_3999,N_3853);
or U4303 (N_4303,N_3726,N_3850);
xnor U4304 (N_4304,N_3776,N_3823);
and U4305 (N_4305,N_3720,N_3620);
nand U4306 (N_4306,N_3975,N_3620);
and U4307 (N_4307,N_3562,N_3524);
nor U4308 (N_4308,N_3777,N_3866);
and U4309 (N_4309,N_3571,N_3766);
nor U4310 (N_4310,N_3505,N_3709);
nand U4311 (N_4311,N_3981,N_3843);
xor U4312 (N_4312,N_3873,N_3913);
or U4313 (N_4313,N_3880,N_3927);
nand U4314 (N_4314,N_3574,N_3656);
and U4315 (N_4315,N_3699,N_3924);
or U4316 (N_4316,N_3635,N_3795);
or U4317 (N_4317,N_3912,N_3637);
and U4318 (N_4318,N_3677,N_3603);
nand U4319 (N_4319,N_3614,N_3540);
xor U4320 (N_4320,N_3985,N_3783);
or U4321 (N_4321,N_3589,N_3716);
nor U4322 (N_4322,N_3521,N_3502);
or U4323 (N_4323,N_3553,N_3979);
nand U4324 (N_4324,N_3802,N_3694);
and U4325 (N_4325,N_3886,N_3909);
nand U4326 (N_4326,N_3787,N_3960);
nand U4327 (N_4327,N_3561,N_3634);
and U4328 (N_4328,N_3893,N_3979);
nand U4329 (N_4329,N_3529,N_3676);
or U4330 (N_4330,N_3519,N_3661);
and U4331 (N_4331,N_3697,N_3662);
xor U4332 (N_4332,N_3694,N_3918);
and U4333 (N_4333,N_3750,N_3539);
nor U4334 (N_4334,N_3957,N_3704);
nand U4335 (N_4335,N_3550,N_3520);
and U4336 (N_4336,N_3938,N_3927);
and U4337 (N_4337,N_3854,N_3500);
and U4338 (N_4338,N_3857,N_3892);
and U4339 (N_4339,N_3951,N_3629);
xor U4340 (N_4340,N_3748,N_3827);
or U4341 (N_4341,N_3693,N_3628);
nor U4342 (N_4342,N_3883,N_3864);
nand U4343 (N_4343,N_3962,N_3550);
and U4344 (N_4344,N_3858,N_3892);
and U4345 (N_4345,N_3795,N_3695);
nor U4346 (N_4346,N_3689,N_3832);
and U4347 (N_4347,N_3564,N_3553);
nand U4348 (N_4348,N_3713,N_3909);
or U4349 (N_4349,N_3652,N_3679);
nor U4350 (N_4350,N_3849,N_3989);
nand U4351 (N_4351,N_3627,N_3921);
xor U4352 (N_4352,N_3574,N_3818);
xnor U4353 (N_4353,N_3981,N_3531);
xnor U4354 (N_4354,N_3595,N_3976);
or U4355 (N_4355,N_3501,N_3920);
nor U4356 (N_4356,N_3682,N_3975);
or U4357 (N_4357,N_3990,N_3630);
nand U4358 (N_4358,N_3916,N_3890);
nor U4359 (N_4359,N_3863,N_3528);
or U4360 (N_4360,N_3619,N_3789);
nor U4361 (N_4361,N_3847,N_3683);
and U4362 (N_4362,N_3613,N_3592);
nor U4363 (N_4363,N_3863,N_3837);
nand U4364 (N_4364,N_3744,N_3717);
and U4365 (N_4365,N_3980,N_3643);
and U4366 (N_4366,N_3724,N_3999);
or U4367 (N_4367,N_3647,N_3960);
nand U4368 (N_4368,N_3697,N_3972);
and U4369 (N_4369,N_3800,N_3602);
and U4370 (N_4370,N_3672,N_3901);
or U4371 (N_4371,N_3584,N_3523);
and U4372 (N_4372,N_3651,N_3851);
and U4373 (N_4373,N_3774,N_3969);
nand U4374 (N_4374,N_3800,N_3903);
xnor U4375 (N_4375,N_3874,N_3583);
nor U4376 (N_4376,N_3660,N_3537);
xnor U4377 (N_4377,N_3596,N_3542);
nor U4378 (N_4378,N_3710,N_3503);
and U4379 (N_4379,N_3591,N_3810);
nand U4380 (N_4380,N_3629,N_3738);
xnor U4381 (N_4381,N_3504,N_3693);
nor U4382 (N_4382,N_3618,N_3524);
nor U4383 (N_4383,N_3921,N_3546);
and U4384 (N_4384,N_3694,N_3705);
xor U4385 (N_4385,N_3619,N_3714);
nor U4386 (N_4386,N_3935,N_3898);
xnor U4387 (N_4387,N_3554,N_3503);
and U4388 (N_4388,N_3800,N_3645);
and U4389 (N_4389,N_3930,N_3707);
and U4390 (N_4390,N_3724,N_3826);
or U4391 (N_4391,N_3832,N_3968);
and U4392 (N_4392,N_3827,N_3714);
nor U4393 (N_4393,N_3855,N_3734);
nor U4394 (N_4394,N_3639,N_3946);
nand U4395 (N_4395,N_3673,N_3656);
nor U4396 (N_4396,N_3982,N_3702);
xnor U4397 (N_4397,N_3976,N_3966);
or U4398 (N_4398,N_3565,N_3966);
nor U4399 (N_4399,N_3967,N_3681);
nor U4400 (N_4400,N_3830,N_3695);
or U4401 (N_4401,N_3968,N_3791);
nor U4402 (N_4402,N_3672,N_3840);
or U4403 (N_4403,N_3669,N_3513);
nor U4404 (N_4404,N_3847,N_3755);
nor U4405 (N_4405,N_3895,N_3869);
nor U4406 (N_4406,N_3572,N_3545);
or U4407 (N_4407,N_3913,N_3802);
and U4408 (N_4408,N_3819,N_3798);
and U4409 (N_4409,N_3853,N_3918);
and U4410 (N_4410,N_3958,N_3798);
nand U4411 (N_4411,N_3987,N_3940);
nor U4412 (N_4412,N_3997,N_3959);
or U4413 (N_4413,N_3763,N_3703);
nand U4414 (N_4414,N_3829,N_3546);
nor U4415 (N_4415,N_3814,N_3771);
and U4416 (N_4416,N_3501,N_3580);
and U4417 (N_4417,N_3659,N_3858);
nor U4418 (N_4418,N_3693,N_3929);
xor U4419 (N_4419,N_3678,N_3922);
xor U4420 (N_4420,N_3811,N_3624);
and U4421 (N_4421,N_3531,N_3958);
nand U4422 (N_4422,N_3892,N_3567);
nor U4423 (N_4423,N_3761,N_3621);
nor U4424 (N_4424,N_3804,N_3870);
and U4425 (N_4425,N_3903,N_3574);
xnor U4426 (N_4426,N_3818,N_3810);
nand U4427 (N_4427,N_3973,N_3574);
nor U4428 (N_4428,N_3887,N_3813);
nand U4429 (N_4429,N_3868,N_3607);
or U4430 (N_4430,N_3649,N_3870);
and U4431 (N_4431,N_3680,N_3809);
nand U4432 (N_4432,N_3805,N_3902);
and U4433 (N_4433,N_3779,N_3660);
nand U4434 (N_4434,N_3923,N_3518);
nor U4435 (N_4435,N_3956,N_3953);
nand U4436 (N_4436,N_3867,N_3947);
nor U4437 (N_4437,N_3569,N_3981);
and U4438 (N_4438,N_3773,N_3749);
xnor U4439 (N_4439,N_3671,N_3725);
or U4440 (N_4440,N_3506,N_3773);
nor U4441 (N_4441,N_3689,N_3956);
and U4442 (N_4442,N_3581,N_3597);
xor U4443 (N_4443,N_3605,N_3892);
xnor U4444 (N_4444,N_3669,N_3666);
and U4445 (N_4445,N_3604,N_3916);
nand U4446 (N_4446,N_3616,N_3995);
and U4447 (N_4447,N_3961,N_3894);
nor U4448 (N_4448,N_3958,N_3746);
or U4449 (N_4449,N_3830,N_3661);
nand U4450 (N_4450,N_3523,N_3905);
nand U4451 (N_4451,N_3500,N_3987);
nor U4452 (N_4452,N_3972,N_3839);
nand U4453 (N_4453,N_3821,N_3664);
and U4454 (N_4454,N_3846,N_3817);
or U4455 (N_4455,N_3512,N_3781);
or U4456 (N_4456,N_3518,N_3716);
nand U4457 (N_4457,N_3841,N_3999);
nand U4458 (N_4458,N_3620,N_3876);
xnor U4459 (N_4459,N_3920,N_3825);
nand U4460 (N_4460,N_3592,N_3576);
nand U4461 (N_4461,N_3516,N_3906);
xor U4462 (N_4462,N_3680,N_3684);
or U4463 (N_4463,N_3770,N_3595);
or U4464 (N_4464,N_3854,N_3582);
and U4465 (N_4465,N_3505,N_3964);
nand U4466 (N_4466,N_3804,N_3930);
nor U4467 (N_4467,N_3613,N_3738);
xnor U4468 (N_4468,N_3590,N_3689);
nor U4469 (N_4469,N_3854,N_3748);
and U4470 (N_4470,N_3581,N_3940);
nor U4471 (N_4471,N_3989,N_3960);
nor U4472 (N_4472,N_3579,N_3765);
and U4473 (N_4473,N_3589,N_3692);
nor U4474 (N_4474,N_3535,N_3676);
nand U4475 (N_4475,N_3908,N_3819);
or U4476 (N_4476,N_3849,N_3999);
or U4477 (N_4477,N_3762,N_3935);
or U4478 (N_4478,N_3507,N_3697);
nor U4479 (N_4479,N_3874,N_3562);
nor U4480 (N_4480,N_3912,N_3804);
nand U4481 (N_4481,N_3811,N_3666);
or U4482 (N_4482,N_3504,N_3826);
nand U4483 (N_4483,N_3794,N_3658);
or U4484 (N_4484,N_3745,N_3622);
nand U4485 (N_4485,N_3578,N_3756);
or U4486 (N_4486,N_3818,N_3656);
and U4487 (N_4487,N_3813,N_3695);
and U4488 (N_4488,N_3727,N_3739);
or U4489 (N_4489,N_3883,N_3924);
nor U4490 (N_4490,N_3624,N_3507);
nor U4491 (N_4491,N_3920,N_3647);
nand U4492 (N_4492,N_3834,N_3515);
nand U4493 (N_4493,N_3947,N_3566);
xnor U4494 (N_4494,N_3606,N_3765);
nor U4495 (N_4495,N_3505,N_3824);
nor U4496 (N_4496,N_3795,N_3785);
nand U4497 (N_4497,N_3767,N_3907);
or U4498 (N_4498,N_3802,N_3918);
or U4499 (N_4499,N_3585,N_3710);
and U4500 (N_4500,N_4241,N_4066);
nor U4501 (N_4501,N_4094,N_4437);
xnor U4502 (N_4502,N_4170,N_4496);
or U4503 (N_4503,N_4065,N_4205);
xnor U4504 (N_4504,N_4275,N_4166);
nand U4505 (N_4505,N_4246,N_4089);
nand U4506 (N_4506,N_4353,N_4109);
nor U4507 (N_4507,N_4443,N_4338);
nor U4508 (N_4508,N_4261,N_4245);
nand U4509 (N_4509,N_4361,N_4177);
xnor U4510 (N_4510,N_4267,N_4175);
nand U4511 (N_4511,N_4279,N_4076);
and U4512 (N_4512,N_4337,N_4217);
or U4513 (N_4513,N_4373,N_4367);
nand U4514 (N_4514,N_4084,N_4440);
nand U4515 (N_4515,N_4482,N_4137);
and U4516 (N_4516,N_4017,N_4403);
and U4517 (N_4517,N_4271,N_4263);
and U4518 (N_4518,N_4215,N_4442);
and U4519 (N_4519,N_4023,N_4291);
and U4520 (N_4520,N_4332,N_4113);
nand U4521 (N_4521,N_4451,N_4457);
or U4522 (N_4522,N_4424,N_4420);
nor U4523 (N_4523,N_4476,N_4311);
or U4524 (N_4524,N_4499,N_4120);
nand U4525 (N_4525,N_4046,N_4003);
nor U4526 (N_4526,N_4301,N_4340);
nand U4527 (N_4527,N_4247,N_4320);
and U4528 (N_4528,N_4075,N_4011);
or U4529 (N_4529,N_4293,N_4185);
nor U4530 (N_4530,N_4411,N_4106);
nand U4531 (N_4531,N_4256,N_4386);
or U4532 (N_4532,N_4484,N_4232);
or U4533 (N_4533,N_4225,N_4234);
or U4534 (N_4534,N_4132,N_4221);
or U4535 (N_4535,N_4207,N_4134);
and U4536 (N_4536,N_4149,N_4196);
and U4537 (N_4537,N_4224,N_4313);
nor U4538 (N_4538,N_4264,N_4034);
and U4539 (N_4539,N_4053,N_4478);
nand U4540 (N_4540,N_4319,N_4074);
nand U4541 (N_4541,N_4335,N_4363);
or U4542 (N_4542,N_4125,N_4243);
nand U4543 (N_4543,N_4212,N_4200);
or U4544 (N_4544,N_4030,N_4356);
and U4545 (N_4545,N_4342,N_4376);
nor U4546 (N_4546,N_4325,N_4299);
nor U4547 (N_4547,N_4439,N_4460);
nor U4548 (N_4548,N_4024,N_4088);
nor U4549 (N_4549,N_4404,N_4131);
and U4550 (N_4550,N_4025,N_4292);
nor U4551 (N_4551,N_4485,N_4422);
and U4552 (N_4552,N_4248,N_4229);
nand U4553 (N_4553,N_4102,N_4123);
and U4554 (N_4554,N_4395,N_4298);
nand U4555 (N_4555,N_4050,N_4117);
and U4556 (N_4556,N_4461,N_4154);
xor U4557 (N_4557,N_4359,N_4231);
or U4558 (N_4558,N_4303,N_4242);
nor U4559 (N_4559,N_4161,N_4321);
and U4560 (N_4560,N_4103,N_4100);
xor U4561 (N_4561,N_4172,N_4198);
or U4562 (N_4562,N_4378,N_4474);
nand U4563 (N_4563,N_4312,N_4020);
xnor U4564 (N_4564,N_4428,N_4083);
nor U4565 (N_4565,N_4009,N_4111);
or U4566 (N_4566,N_4431,N_4368);
nand U4567 (N_4567,N_4223,N_4163);
nor U4568 (N_4568,N_4153,N_4080);
xor U4569 (N_4569,N_4458,N_4390);
nand U4570 (N_4570,N_4201,N_4369);
nor U4571 (N_4571,N_4262,N_4236);
or U4572 (N_4572,N_4018,N_4493);
nor U4573 (N_4573,N_4416,N_4189);
and U4574 (N_4574,N_4456,N_4060);
or U4575 (N_4575,N_4069,N_4391);
xnor U4576 (N_4576,N_4228,N_4194);
and U4577 (N_4577,N_4334,N_4494);
or U4578 (N_4578,N_4001,N_4021);
nand U4579 (N_4579,N_4164,N_4160);
nor U4580 (N_4580,N_4048,N_4341);
nand U4581 (N_4581,N_4295,N_4276);
nor U4582 (N_4582,N_4294,N_4097);
nand U4583 (N_4583,N_4366,N_4141);
nand U4584 (N_4584,N_4498,N_4202);
nor U4585 (N_4585,N_4426,N_4392);
nor U4586 (N_4586,N_4396,N_4107);
nor U4587 (N_4587,N_4054,N_4110);
nand U4588 (N_4588,N_4430,N_4441);
or U4589 (N_4589,N_4273,N_4220);
nand U4590 (N_4590,N_4027,N_4122);
or U4591 (N_4591,N_4381,N_4380);
and U4592 (N_4592,N_4272,N_4346);
and U4593 (N_4593,N_4310,N_4357);
nand U4594 (N_4594,N_4423,N_4049);
nor U4595 (N_4595,N_4007,N_4186);
or U4596 (N_4596,N_4324,N_4182);
and U4597 (N_4597,N_4281,N_4497);
or U4598 (N_4598,N_4093,N_4022);
and U4599 (N_4599,N_4147,N_4427);
and U4600 (N_4600,N_4173,N_4126);
and U4601 (N_4601,N_4284,N_4285);
or U4602 (N_4602,N_4429,N_4410);
xor U4603 (N_4603,N_4061,N_4377);
xnor U4604 (N_4604,N_4370,N_4056);
nand U4605 (N_4605,N_4387,N_4218);
nor U4606 (N_4606,N_4266,N_4032);
nor U4607 (N_4607,N_4468,N_4059);
and U4608 (N_4608,N_4128,N_4449);
or U4609 (N_4609,N_4283,N_4492);
and U4610 (N_4610,N_4150,N_4090);
xor U4611 (N_4611,N_4270,N_4286);
or U4612 (N_4612,N_4121,N_4167);
and U4613 (N_4613,N_4063,N_4214);
nor U4614 (N_4614,N_4033,N_4447);
and U4615 (N_4615,N_4406,N_4129);
and U4616 (N_4616,N_4462,N_4336);
or U4617 (N_4617,N_4136,N_4274);
and U4618 (N_4618,N_4133,N_4067);
nor U4619 (N_4619,N_4038,N_4290);
or U4620 (N_4620,N_4251,N_4385);
nand U4621 (N_4621,N_4178,N_4124);
nor U4622 (N_4622,N_4327,N_4148);
nor U4623 (N_4623,N_4306,N_4183);
nor U4624 (N_4624,N_4491,N_4344);
or U4625 (N_4625,N_4328,N_4415);
and U4626 (N_4626,N_4412,N_4058);
nor U4627 (N_4627,N_4176,N_4152);
and U4628 (N_4628,N_4169,N_4008);
nor U4629 (N_4629,N_4157,N_4216);
or U4630 (N_4630,N_4265,N_4471);
nand U4631 (N_4631,N_4179,N_4316);
xnor U4632 (N_4632,N_4425,N_4364);
xor U4633 (N_4633,N_4227,N_4195);
xnor U4634 (N_4634,N_4250,N_4397);
and U4635 (N_4635,N_4233,N_4401);
and U4636 (N_4636,N_4278,N_4486);
nor U4637 (N_4637,N_4039,N_4331);
xor U4638 (N_4638,N_4101,N_4091);
and U4639 (N_4639,N_4318,N_4288);
or U4640 (N_4640,N_4019,N_4255);
nor U4641 (N_4641,N_4098,N_4193);
nand U4642 (N_4642,N_4191,N_4105);
nand U4643 (N_4643,N_4143,N_4012);
or U4644 (N_4644,N_4052,N_4068);
nor U4645 (N_4645,N_4302,N_4419);
and U4646 (N_4646,N_4490,N_4211);
or U4647 (N_4647,N_4322,N_4037);
nor U4648 (N_4648,N_4145,N_4259);
nor U4649 (N_4649,N_4280,N_4174);
and U4650 (N_4650,N_4055,N_4465);
or U4651 (N_4651,N_4287,N_4297);
nand U4652 (N_4652,N_4467,N_4162);
nor U4653 (N_4653,N_4151,N_4488);
or U4654 (N_4654,N_4330,N_4454);
nand U4655 (N_4655,N_4070,N_4452);
nand U4656 (N_4656,N_4130,N_4345);
and U4657 (N_4657,N_4142,N_4146);
or U4658 (N_4658,N_4408,N_4190);
and U4659 (N_4659,N_4326,N_4495);
and U4660 (N_4660,N_4043,N_4282);
nand U4661 (N_4661,N_4477,N_4237);
nand U4662 (N_4662,N_4015,N_4144);
and U4663 (N_4663,N_4464,N_4343);
or U4664 (N_4664,N_4314,N_4064);
and U4665 (N_4665,N_4192,N_4339);
nand U4666 (N_4666,N_4184,N_4487);
or U4667 (N_4667,N_4383,N_4042);
or U4668 (N_4668,N_4206,N_4257);
or U4669 (N_4669,N_4300,N_4135);
nand U4670 (N_4670,N_4333,N_4140);
or U4671 (N_4671,N_4085,N_4252);
nand U4672 (N_4672,N_4036,N_4349);
or U4673 (N_4673,N_4219,N_4375);
xor U4674 (N_4674,N_4026,N_4139);
xnor U4675 (N_4675,N_4350,N_4400);
nand U4676 (N_4676,N_4099,N_4358);
nand U4677 (N_4677,N_4062,N_4365);
or U4678 (N_4678,N_4296,N_4096);
or U4679 (N_4679,N_4158,N_4388);
and U4680 (N_4680,N_4047,N_4181);
or U4681 (N_4681,N_4414,N_4116);
xnor U4682 (N_4682,N_4044,N_4014);
xnor U4683 (N_4683,N_4000,N_4006);
and U4684 (N_4684,N_4077,N_4435);
or U4685 (N_4685,N_4029,N_4384);
nand U4686 (N_4686,N_4071,N_4389);
or U4687 (N_4687,N_4244,N_4171);
nand U4688 (N_4688,N_4393,N_4118);
nor U4689 (N_4689,N_4348,N_4459);
or U4690 (N_4690,N_4114,N_4394);
xnor U4691 (N_4691,N_4479,N_4269);
and U4692 (N_4692,N_4455,N_4045);
nand U4693 (N_4693,N_4086,N_4226);
nor U4694 (N_4694,N_4413,N_4309);
or U4695 (N_4695,N_4204,N_4438);
xor U4696 (N_4696,N_4355,N_4407);
nor U4697 (N_4697,N_4238,N_4323);
nor U4698 (N_4698,N_4254,N_4127);
nor U4699 (N_4699,N_4010,N_4258);
or U4700 (N_4700,N_4445,N_4433);
nor U4701 (N_4701,N_4188,N_4379);
and U4702 (N_4702,N_4016,N_4031);
nand U4703 (N_4703,N_4304,N_4317);
nor U4704 (N_4704,N_4235,N_4253);
nand U4705 (N_4705,N_4277,N_4473);
nand U4706 (N_4706,N_4108,N_4448);
xnor U4707 (N_4707,N_4004,N_4453);
nand U4708 (N_4708,N_4035,N_4351);
nand U4709 (N_4709,N_4203,N_4450);
nand U4710 (N_4710,N_4308,N_4180);
nand U4711 (N_4711,N_4028,N_4472);
and U4712 (N_4712,N_4399,N_4230);
nor U4713 (N_4713,N_4347,N_4260);
or U4714 (N_4714,N_4409,N_4480);
xnor U4715 (N_4715,N_4095,N_4104);
and U4716 (N_4716,N_4268,N_4417);
or U4717 (N_4717,N_4371,N_4418);
and U4718 (N_4718,N_4240,N_4078);
and U4719 (N_4719,N_4168,N_4187);
xnor U4720 (N_4720,N_4469,N_4197);
xnor U4721 (N_4721,N_4115,N_4222);
or U4722 (N_4722,N_4307,N_4112);
and U4723 (N_4723,N_4041,N_4289);
xor U4724 (N_4724,N_4002,N_4398);
nor U4725 (N_4725,N_4329,N_4040);
and U4726 (N_4726,N_4057,N_4209);
or U4727 (N_4727,N_4072,N_4434);
xor U4728 (N_4728,N_4436,N_4082);
nand U4729 (N_4729,N_4483,N_4405);
nor U4730 (N_4730,N_4446,N_4315);
nand U4731 (N_4731,N_4374,N_4360);
and U4732 (N_4732,N_4092,N_4402);
and U4733 (N_4733,N_4073,N_4444);
and U4734 (N_4734,N_4470,N_4432);
nor U4735 (N_4735,N_4305,N_4466);
or U4736 (N_4736,N_4087,N_4489);
and U4737 (N_4737,N_4079,N_4249);
xnor U4738 (N_4738,N_4138,N_4155);
or U4739 (N_4739,N_4013,N_4199);
or U4740 (N_4740,N_4081,N_4051);
or U4741 (N_4741,N_4481,N_4165);
nand U4742 (N_4742,N_4005,N_4213);
nand U4743 (N_4743,N_4475,N_4119);
nand U4744 (N_4744,N_4156,N_4382);
or U4745 (N_4745,N_4239,N_4354);
nand U4746 (N_4746,N_4210,N_4372);
and U4747 (N_4747,N_4421,N_4352);
nand U4748 (N_4748,N_4208,N_4463);
nand U4749 (N_4749,N_4362,N_4159);
or U4750 (N_4750,N_4317,N_4145);
nand U4751 (N_4751,N_4449,N_4412);
nor U4752 (N_4752,N_4274,N_4271);
and U4753 (N_4753,N_4090,N_4399);
and U4754 (N_4754,N_4306,N_4339);
nor U4755 (N_4755,N_4467,N_4447);
nor U4756 (N_4756,N_4139,N_4296);
and U4757 (N_4757,N_4051,N_4097);
and U4758 (N_4758,N_4235,N_4217);
and U4759 (N_4759,N_4151,N_4017);
and U4760 (N_4760,N_4459,N_4358);
nor U4761 (N_4761,N_4361,N_4371);
or U4762 (N_4762,N_4290,N_4370);
and U4763 (N_4763,N_4426,N_4298);
nand U4764 (N_4764,N_4477,N_4423);
xor U4765 (N_4765,N_4074,N_4138);
or U4766 (N_4766,N_4175,N_4187);
or U4767 (N_4767,N_4003,N_4140);
or U4768 (N_4768,N_4277,N_4072);
nand U4769 (N_4769,N_4482,N_4090);
xnor U4770 (N_4770,N_4488,N_4387);
or U4771 (N_4771,N_4292,N_4329);
nand U4772 (N_4772,N_4304,N_4343);
or U4773 (N_4773,N_4263,N_4395);
nor U4774 (N_4774,N_4150,N_4104);
or U4775 (N_4775,N_4114,N_4473);
nor U4776 (N_4776,N_4483,N_4130);
nor U4777 (N_4777,N_4074,N_4429);
or U4778 (N_4778,N_4039,N_4373);
nand U4779 (N_4779,N_4196,N_4427);
nor U4780 (N_4780,N_4349,N_4060);
nand U4781 (N_4781,N_4016,N_4264);
nor U4782 (N_4782,N_4162,N_4034);
nand U4783 (N_4783,N_4413,N_4437);
nor U4784 (N_4784,N_4118,N_4264);
nand U4785 (N_4785,N_4119,N_4063);
and U4786 (N_4786,N_4419,N_4428);
and U4787 (N_4787,N_4324,N_4204);
and U4788 (N_4788,N_4180,N_4234);
nand U4789 (N_4789,N_4164,N_4125);
nand U4790 (N_4790,N_4425,N_4450);
nand U4791 (N_4791,N_4435,N_4316);
nand U4792 (N_4792,N_4492,N_4009);
or U4793 (N_4793,N_4256,N_4470);
and U4794 (N_4794,N_4317,N_4072);
xor U4795 (N_4795,N_4182,N_4293);
or U4796 (N_4796,N_4164,N_4366);
and U4797 (N_4797,N_4464,N_4089);
xor U4798 (N_4798,N_4126,N_4392);
nand U4799 (N_4799,N_4287,N_4213);
or U4800 (N_4800,N_4198,N_4415);
nor U4801 (N_4801,N_4212,N_4322);
nand U4802 (N_4802,N_4182,N_4049);
and U4803 (N_4803,N_4266,N_4022);
or U4804 (N_4804,N_4220,N_4310);
nand U4805 (N_4805,N_4018,N_4498);
nand U4806 (N_4806,N_4393,N_4056);
nand U4807 (N_4807,N_4166,N_4155);
or U4808 (N_4808,N_4041,N_4304);
nor U4809 (N_4809,N_4108,N_4455);
nor U4810 (N_4810,N_4239,N_4487);
and U4811 (N_4811,N_4050,N_4407);
and U4812 (N_4812,N_4302,N_4293);
or U4813 (N_4813,N_4342,N_4117);
and U4814 (N_4814,N_4139,N_4265);
or U4815 (N_4815,N_4231,N_4058);
nor U4816 (N_4816,N_4416,N_4200);
nand U4817 (N_4817,N_4171,N_4235);
or U4818 (N_4818,N_4341,N_4388);
or U4819 (N_4819,N_4106,N_4039);
nand U4820 (N_4820,N_4214,N_4273);
nand U4821 (N_4821,N_4247,N_4297);
nand U4822 (N_4822,N_4146,N_4085);
nor U4823 (N_4823,N_4383,N_4487);
nor U4824 (N_4824,N_4005,N_4148);
nand U4825 (N_4825,N_4445,N_4115);
nor U4826 (N_4826,N_4037,N_4248);
or U4827 (N_4827,N_4450,N_4300);
and U4828 (N_4828,N_4402,N_4070);
nand U4829 (N_4829,N_4449,N_4420);
nor U4830 (N_4830,N_4394,N_4049);
xor U4831 (N_4831,N_4411,N_4427);
nand U4832 (N_4832,N_4405,N_4263);
and U4833 (N_4833,N_4481,N_4230);
nand U4834 (N_4834,N_4055,N_4249);
nand U4835 (N_4835,N_4019,N_4444);
nor U4836 (N_4836,N_4132,N_4406);
or U4837 (N_4837,N_4242,N_4380);
and U4838 (N_4838,N_4285,N_4187);
and U4839 (N_4839,N_4076,N_4289);
nand U4840 (N_4840,N_4302,N_4499);
nor U4841 (N_4841,N_4415,N_4063);
nand U4842 (N_4842,N_4188,N_4361);
nor U4843 (N_4843,N_4060,N_4359);
xnor U4844 (N_4844,N_4444,N_4471);
or U4845 (N_4845,N_4240,N_4155);
or U4846 (N_4846,N_4261,N_4381);
or U4847 (N_4847,N_4226,N_4189);
nor U4848 (N_4848,N_4291,N_4224);
nor U4849 (N_4849,N_4382,N_4153);
and U4850 (N_4850,N_4044,N_4368);
xnor U4851 (N_4851,N_4116,N_4086);
and U4852 (N_4852,N_4376,N_4076);
xnor U4853 (N_4853,N_4254,N_4184);
nand U4854 (N_4854,N_4118,N_4107);
nor U4855 (N_4855,N_4023,N_4020);
nor U4856 (N_4856,N_4005,N_4076);
and U4857 (N_4857,N_4029,N_4387);
nor U4858 (N_4858,N_4034,N_4120);
nor U4859 (N_4859,N_4351,N_4189);
or U4860 (N_4860,N_4220,N_4227);
and U4861 (N_4861,N_4358,N_4463);
and U4862 (N_4862,N_4497,N_4327);
nand U4863 (N_4863,N_4180,N_4032);
or U4864 (N_4864,N_4226,N_4180);
and U4865 (N_4865,N_4026,N_4394);
xnor U4866 (N_4866,N_4123,N_4146);
and U4867 (N_4867,N_4413,N_4052);
and U4868 (N_4868,N_4218,N_4221);
xor U4869 (N_4869,N_4169,N_4009);
and U4870 (N_4870,N_4137,N_4391);
or U4871 (N_4871,N_4486,N_4377);
or U4872 (N_4872,N_4215,N_4032);
nor U4873 (N_4873,N_4490,N_4322);
nand U4874 (N_4874,N_4129,N_4027);
nor U4875 (N_4875,N_4185,N_4393);
nor U4876 (N_4876,N_4352,N_4077);
or U4877 (N_4877,N_4291,N_4064);
and U4878 (N_4878,N_4066,N_4408);
nor U4879 (N_4879,N_4250,N_4418);
nand U4880 (N_4880,N_4218,N_4070);
nand U4881 (N_4881,N_4126,N_4093);
or U4882 (N_4882,N_4451,N_4462);
or U4883 (N_4883,N_4060,N_4463);
nor U4884 (N_4884,N_4046,N_4437);
nor U4885 (N_4885,N_4497,N_4310);
and U4886 (N_4886,N_4140,N_4463);
or U4887 (N_4887,N_4074,N_4154);
and U4888 (N_4888,N_4054,N_4459);
nor U4889 (N_4889,N_4101,N_4471);
and U4890 (N_4890,N_4293,N_4047);
nand U4891 (N_4891,N_4439,N_4048);
nor U4892 (N_4892,N_4045,N_4268);
or U4893 (N_4893,N_4115,N_4473);
and U4894 (N_4894,N_4066,N_4007);
nand U4895 (N_4895,N_4275,N_4176);
or U4896 (N_4896,N_4101,N_4386);
nor U4897 (N_4897,N_4479,N_4276);
nor U4898 (N_4898,N_4307,N_4233);
or U4899 (N_4899,N_4120,N_4029);
and U4900 (N_4900,N_4111,N_4047);
nand U4901 (N_4901,N_4375,N_4252);
nor U4902 (N_4902,N_4449,N_4291);
or U4903 (N_4903,N_4065,N_4115);
or U4904 (N_4904,N_4104,N_4278);
nand U4905 (N_4905,N_4022,N_4468);
or U4906 (N_4906,N_4177,N_4388);
and U4907 (N_4907,N_4058,N_4128);
nor U4908 (N_4908,N_4397,N_4068);
xor U4909 (N_4909,N_4102,N_4116);
nor U4910 (N_4910,N_4308,N_4254);
or U4911 (N_4911,N_4312,N_4105);
or U4912 (N_4912,N_4490,N_4237);
xor U4913 (N_4913,N_4096,N_4421);
nand U4914 (N_4914,N_4341,N_4161);
or U4915 (N_4915,N_4006,N_4308);
nand U4916 (N_4916,N_4054,N_4463);
nor U4917 (N_4917,N_4082,N_4249);
xor U4918 (N_4918,N_4075,N_4067);
nand U4919 (N_4919,N_4355,N_4058);
and U4920 (N_4920,N_4272,N_4496);
nand U4921 (N_4921,N_4081,N_4281);
nand U4922 (N_4922,N_4139,N_4040);
and U4923 (N_4923,N_4273,N_4228);
nand U4924 (N_4924,N_4166,N_4262);
nand U4925 (N_4925,N_4144,N_4104);
nor U4926 (N_4926,N_4294,N_4193);
or U4927 (N_4927,N_4425,N_4068);
and U4928 (N_4928,N_4163,N_4170);
xnor U4929 (N_4929,N_4044,N_4038);
nand U4930 (N_4930,N_4019,N_4224);
and U4931 (N_4931,N_4353,N_4280);
xor U4932 (N_4932,N_4043,N_4019);
nand U4933 (N_4933,N_4488,N_4355);
nor U4934 (N_4934,N_4145,N_4013);
and U4935 (N_4935,N_4314,N_4336);
or U4936 (N_4936,N_4019,N_4212);
xnor U4937 (N_4937,N_4222,N_4276);
or U4938 (N_4938,N_4150,N_4093);
nor U4939 (N_4939,N_4106,N_4194);
and U4940 (N_4940,N_4493,N_4246);
or U4941 (N_4941,N_4253,N_4175);
xor U4942 (N_4942,N_4498,N_4401);
nor U4943 (N_4943,N_4442,N_4433);
nor U4944 (N_4944,N_4060,N_4384);
or U4945 (N_4945,N_4119,N_4025);
and U4946 (N_4946,N_4088,N_4412);
or U4947 (N_4947,N_4107,N_4161);
xnor U4948 (N_4948,N_4307,N_4353);
nor U4949 (N_4949,N_4418,N_4242);
nand U4950 (N_4950,N_4255,N_4191);
nor U4951 (N_4951,N_4372,N_4059);
and U4952 (N_4952,N_4255,N_4199);
nor U4953 (N_4953,N_4166,N_4296);
and U4954 (N_4954,N_4284,N_4346);
nor U4955 (N_4955,N_4212,N_4083);
nand U4956 (N_4956,N_4189,N_4404);
or U4957 (N_4957,N_4481,N_4483);
and U4958 (N_4958,N_4014,N_4104);
nand U4959 (N_4959,N_4307,N_4415);
or U4960 (N_4960,N_4100,N_4227);
nor U4961 (N_4961,N_4367,N_4294);
or U4962 (N_4962,N_4402,N_4459);
nand U4963 (N_4963,N_4426,N_4080);
nand U4964 (N_4964,N_4224,N_4288);
and U4965 (N_4965,N_4317,N_4253);
nor U4966 (N_4966,N_4084,N_4181);
and U4967 (N_4967,N_4063,N_4199);
or U4968 (N_4968,N_4176,N_4398);
nor U4969 (N_4969,N_4162,N_4201);
xor U4970 (N_4970,N_4190,N_4130);
nand U4971 (N_4971,N_4484,N_4169);
or U4972 (N_4972,N_4314,N_4176);
nor U4973 (N_4973,N_4427,N_4223);
or U4974 (N_4974,N_4082,N_4077);
nor U4975 (N_4975,N_4455,N_4459);
and U4976 (N_4976,N_4263,N_4472);
or U4977 (N_4977,N_4403,N_4263);
nand U4978 (N_4978,N_4187,N_4104);
nor U4979 (N_4979,N_4066,N_4154);
nand U4980 (N_4980,N_4083,N_4417);
or U4981 (N_4981,N_4318,N_4432);
nand U4982 (N_4982,N_4421,N_4006);
and U4983 (N_4983,N_4148,N_4224);
and U4984 (N_4984,N_4157,N_4425);
nand U4985 (N_4985,N_4258,N_4321);
nor U4986 (N_4986,N_4492,N_4226);
and U4987 (N_4987,N_4461,N_4460);
or U4988 (N_4988,N_4285,N_4112);
nor U4989 (N_4989,N_4336,N_4298);
xnor U4990 (N_4990,N_4143,N_4149);
and U4991 (N_4991,N_4143,N_4375);
and U4992 (N_4992,N_4273,N_4195);
xor U4993 (N_4993,N_4371,N_4012);
or U4994 (N_4994,N_4371,N_4289);
nand U4995 (N_4995,N_4001,N_4457);
nor U4996 (N_4996,N_4346,N_4356);
nand U4997 (N_4997,N_4158,N_4003);
nand U4998 (N_4998,N_4000,N_4470);
or U4999 (N_4999,N_4182,N_4349);
or U5000 (N_5000,N_4626,N_4500);
nand U5001 (N_5001,N_4980,N_4870);
and U5002 (N_5002,N_4922,N_4800);
or U5003 (N_5003,N_4576,N_4816);
nor U5004 (N_5004,N_4811,N_4911);
nor U5005 (N_5005,N_4621,N_4603);
or U5006 (N_5006,N_4827,N_4961);
xor U5007 (N_5007,N_4732,N_4503);
or U5008 (N_5008,N_4643,N_4650);
nor U5009 (N_5009,N_4677,N_4613);
or U5010 (N_5010,N_4652,N_4883);
nor U5011 (N_5011,N_4695,N_4644);
nor U5012 (N_5012,N_4558,N_4531);
xor U5013 (N_5013,N_4794,N_4769);
or U5014 (N_5014,N_4987,N_4688);
or U5015 (N_5015,N_4657,N_4886);
or U5016 (N_5016,N_4612,N_4895);
or U5017 (N_5017,N_4791,N_4519);
nor U5018 (N_5018,N_4983,N_4540);
and U5019 (N_5019,N_4855,N_4908);
nor U5020 (N_5020,N_4708,N_4590);
and U5021 (N_5021,N_4945,N_4937);
nor U5022 (N_5022,N_4593,N_4918);
nand U5023 (N_5023,N_4954,N_4507);
or U5024 (N_5024,N_4705,N_4990);
or U5025 (N_5025,N_4551,N_4736);
or U5026 (N_5026,N_4774,N_4524);
or U5027 (N_5027,N_4675,N_4521);
nor U5028 (N_5028,N_4926,N_4923);
xnor U5029 (N_5029,N_4698,N_4817);
or U5030 (N_5030,N_4998,N_4629);
nor U5031 (N_5031,N_4527,N_4869);
nor U5032 (N_5032,N_4599,N_4873);
xnor U5033 (N_5033,N_4820,N_4985);
and U5034 (N_5034,N_4938,N_4528);
nor U5035 (N_5035,N_4806,N_4824);
and U5036 (N_5036,N_4701,N_4501);
or U5037 (N_5037,N_4667,N_4766);
and U5038 (N_5038,N_4971,N_4569);
nand U5039 (N_5039,N_4964,N_4788);
nand U5040 (N_5040,N_4660,N_4738);
nor U5041 (N_5041,N_4856,N_4866);
or U5042 (N_5042,N_4796,N_4628);
nor U5043 (N_5043,N_4703,N_4608);
nor U5044 (N_5044,N_4779,N_4616);
and U5045 (N_5045,N_4823,N_4729);
nand U5046 (N_5046,N_4597,N_4720);
xnor U5047 (N_5047,N_4755,N_4741);
and U5048 (N_5048,N_4844,N_4826);
nor U5049 (N_5049,N_4759,N_4799);
and U5050 (N_5050,N_4902,N_4974);
xor U5051 (N_5051,N_4694,N_4790);
or U5052 (N_5052,N_4615,N_4950);
nand U5053 (N_5053,N_4589,N_4997);
nand U5054 (N_5054,N_4932,N_4511);
or U5055 (N_5055,N_4887,N_4994);
or U5056 (N_5056,N_4840,N_4762);
or U5057 (N_5057,N_4939,N_4696);
and U5058 (N_5058,N_4903,N_4999);
nor U5059 (N_5059,N_4967,N_4775);
and U5060 (N_5060,N_4525,N_4739);
or U5061 (N_5061,N_4929,N_4522);
xor U5062 (N_5062,N_4556,N_4976);
nor U5063 (N_5063,N_4829,N_4842);
nand U5064 (N_5064,N_4959,N_4965);
or U5065 (N_5065,N_4624,N_4515);
nor U5066 (N_5066,N_4570,N_4655);
or U5067 (N_5067,N_4575,N_4512);
xnor U5068 (N_5068,N_4681,N_4649);
and U5069 (N_5069,N_4863,N_4936);
nand U5070 (N_5070,N_4931,N_4854);
nand U5071 (N_5071,N_4952,N_4822);
and U5072 (N_5072,N_4735,N_4859);
nand U5073 (N_5073,N_4819,N_4927);
and U5074 (N_5074,N_4878,N_4901);
nand U5075 (N_5075,N_4921,N_4666);
or U5076 (N_5076,N_4579,N_4640);
and U5077 (N_5077,N_4723,N_4546);
or U5078 (N_5078,N_4710,N_4530);
or U5079 (N_5079,N_4958,N_4635);
or U5080 (N_5080,N_4913,N_4697);
or U5081 (N_5081,N_4646,N_4583);
nand U5082 (N_5082,N_4702,N_4880);
and U5083 (N_5083,N_4555,N_4768);
or U5084 (N_5084,N_4784,N_4719);
and U5085 (N_5085,N_4747,N_4944);
and U5086 (N_5086,N_4962,N_4773);
or U5087 (N_5087,N_4605,N_4673);
or U5088 (N_5088,N_4905,N_4686);
xor U5089 (N_5089,N_4843,N_4838);
nor U5090 (N_5090,N_4948,N_4641);
and U5091 (N_5091,N_4668,N_4510);
xor U5092 (N_5092,N_4912,N_4591);
and U5093 (N_5093,N_4632,N_4804);
nor U5094 (N_5094,N_4953,N_4991);
nor U5095 (N_5095,N_4572,N_4849);
nor U5096 (N_5096,N_4907,N_4864);
xnor U5097 (N_5097,N_4581,N_4969);
xnor U5098 (N_5098,N_4814,N_4627);
nor U5099 (N_5099,N_4853,N_4563);
and U5100 (N_5100,N_4847,N_4728);
nand U5101 (N_5101,N_4573,N_4834);
nand U5102 (N_5102,N_4692,N_4638);
nand U5103 (N_5103,N_4973,N_4665);
and U5104 (N_5104,N_4727,N_4809);
and U5105 (N_5105,N_4516,N_4781);
or U5106 (N_5106,N_4951,N_4956);
or U5107 (N_5107,N_4725,N_4566);
nand U5108 (N_5108,N_4633,N_4707);
and U5109 (N_5109,N_4808,N_4792);
and U5110 (N_5110,N_4682,N_4631);
nand U5111 (N_5111,N_4574,N_4656);
and U5112 (N_5112,N_4868,N_4831);
and U5113 (N_5113,N_4896,N_4722);
or U5114 (N_5114,N_4984,N_4772);
or U5115 (N_5115,N_4683,N_4639);
and U5116 (N_5116,N_4562,N_4552);
and U5117 (N_5117,N_4748,N_4687);
nand U5118 (N_5118,N_4770,N_4571);
or U5119 (N_5119,N_4716,N_4506);
or U5120 (N_5120,N_4882,N_4812);
and U5121 (N_5121,N_4715,N_4509);
nand U5122 (N_5122,N_4963,N_4798);
or U5123 (N_5123,N_4598,N_4737);
and U5124 (N_5124,N_4934,N_4744);
nand U5125 (N_5125,N_4915,N_4756);
nor U5126 (N_5126,N_4982,N_4925);
nor U5127 (N_5127,N_4596,N_4778);
and U5128 (N_5128,N_4928,N_4807);
and U5129 (N_5129,N_4797,N_4933);
nor U5130 (N_5130,N_4517,N_4542);
and U5131 (N_5131,N_4508,N_4718);
nand U5132 (N_5132,N_4502,N_4802);
nand U5133 (N_5133,N_4582,N_4654);
nor U5134 (N_5134,N_4536,N_4989);
and U5135 (N_5135,N_4610,N_4712);
nand U5136 (N_5136,N_4679,N_4753);
and U5137 (N_5137,N_4648,N_4529);
nand U5138 (N_5138,N_4609,N_4541);
nand U5139 (N_5139,N_4765,N_4543);
nand U5140 (N_5140,N_4520,N_4538);
nand U5141 (N_5141,N_4904,N_4504);
or U5142 (N_5142,N_4988,N_4604);
nor U5143 (N_5143,N_4978,N_4785);
or U5144 (N_5144,N_4601,N_4889);
nor U5145 (N_5145,N_4691,N_4595);
or U5146 (N_5146,N_4514,N_4890);
and U5147 (N_5147,N_4943,N_4949);
and U5148 (N_5148,N_4548,N_4783);
xnor U5149 (N_5149,N_4534,N_4565);
and U5150 (N_5150,N_4587,N_4545);
and U5151 (N_5151,N_4940,N_4602);
or U5152 (N_5152,N_4793,N_4600);
or U5153 (N_5153,N_4845,N_4841);
and U5154 (N_5154,N_4674,N_4975);
xnor U5155 (N_5155,N_4586,N_4625);
or U5156 (N_5156,N_4846,N_4771);
or U5157 (N_5157,N_4689,N_4815);
nand U5158 (N_5158,N_4761,N_4678);
nand U5159 (N_5159,N_4561,N_4850);
nor U5160 (N_5160,N_4557,N_4550);
nor U5161 (N_5161,N_4818,N_4726);
and U5162 (N_5162,N_4752,N_4981);
and U5163 (N_5163,N_4664,N_4754);
nor U5164 (N_5164,N_4955,N_4941);
or U5165 (N_5165,N_4700,N_4786);
or U5166 (N_5166,N_4881,N_4693);
and U5167 (N_5167,N_4833,N_4636);
nand U5168 (N_5168,N_4897,N_4659);
nand U5169 (N_5169,N_4885,N_4776);
and U5170 (N_5170,N_4651,N_4992);
and U5171 (N_5171,N_4935,N_4618);
or U5172 (N_5172,N_4709,N_4622);
and U5173 (N_5173,N_4544,N_4930);
nand U5174 (N_5174,N_4871,N_4505);
nor U5175 (N_5175,N_4642,N_4900);
xor U5176 (N_5176,N_4518,N_4730);
or U5177 (N_5177,N_4763,N_4825);
nand U5178 (N_5178,N_4924,N_4832);
nor U5179 (N_5179,N_4858,N_4690);
nor U5180 (N_5180,N_4917,N_4714);
nand U5181 (N_5181,N_4594,N_4749);
or U5182 (N_5182,N_4942,N_4580);
and U5183 (N_5183,N_4837,N_4611);
nand U5184 (N_5184,N_4526,N_4782);
and U5185 (N_5185,N_4828,N_4789);
nand U5186 (N_5186,N_4606,N_4877);
and U5187 (N_5187,N_4564,N_4711);
nand U5188 (N_5188,N_4879,N_4630);
and U5189 (N_5189,N_4746,N_4539);
nor U5190 (N_5190,N_4717,N_4685);
or U5191 (N_5191,N_4970,N_4872);
nor U5192 (N_5192,N_4852,N_4891);
xnor U5193 (N_5193,N_4875,N_4721);
nor U5194 (N_5194,N_4892,N_4742);
or U5195 (N_5195,N_4658,N_4745);
nand U5196 (N_5196,N_4713,N_4986);
nand U5197 (N_5197,N_4734,N_4906);
and U5198 (N_5198,N_4568,N_4767);
nor U5199 (N_5199,N_4513,N_4957);
nand U5200 (N_5200,N_4860,N_4647);
or U5201 (N_5201,N_4758,N_4966);
nand U5202 (N_5202,N_4920,N_4620);
nor U5203 (N_5203,N_4733,N_4909);
or U5204 (N_5204,N_4787,N_4740);
nand U5205 (N_5205,N_4663,N_4743);
or U5206 (N_5206,N_4995,N_4547);
or U5207 (N_5207,N_4862,N_4724);
or U5208 (N_5208,N_4757,N_4645);
or U5209 (N_5209,N_4588,N_4919);
nand U5210 (N_5210,N_4671,N_4795);
nor U5211 (N_5211,N_4848,N_4549);
xnor U5212 (N_5212,N_4780,N_4653);
or U5213 (N_5213,N_4607,N_4813);
nand U5214 (N_5214,N_4578,N_4968);
or U5215 (N_5215,N_4567,N_4554);
nor U5216 (N_5216,N_4876,N_4532);
xor U5217 (N_5217,N_4884,N_4836);
or U5218 (N_5218,N_4672,N_4592);
nand U5219 (N_5219,N_4559,N_4865);
nand U5220 (N_5220,N_4898,N_4947);
and U5221 (N_5221,N_4972,N_4751);
nor U5222 (N_5222,N_4979,N_4867);
xnor U5223 (N_5223,N_4704,N_4623);
and U5224 (N_5224,N_4993,N_4577);
nand U5225 (N_5225,N_4888,N_4894);
and U5226 (N_5226,N_4537,N_4670);
or U5227 (N_5227,N_4977,N_4662);
or U5228 (N_5228,N_4893,N_4560);
nand U5229 (N_5229,N_4760,N_4861);
or U5230 (N_5230,N_4821,N_4617);
xnor U5231 (N_5231,N_4637,N_4835);
nor U5232 (N_5232,N_4699,N_4533);
or U5233 (N_5233,N_4874,N_4553);
and U5234 (N_5234,N_4535,N_4669);
nor U5235 (N_5235,N_4839,N_4614);
nand U5236 (N_5236,N_4706,N_4661);
nand U5237 (N_5237,N_4810,N_4996);
and U5238 (N_5238,N_4634,N_4946);
and U5239 (N_5239,N_4960,N_4830);
and U5240 (N_5240,N_4916,N_4910);
and U5241 (N_5241,N_4619,N_4585);
nor U5242 (N_5242,N_4764,N_4851);
or U5243 (N_5243,N_4731,N_4899);
nor U5244 (N_5244,N_4750,N_4801);
nand U5245 (N_5245,N_4805,N_4803);
nand U5246 (N_5246,N_4857,N_4680);
or U5247 (N_5247,N_4676,N_4914);
or U5248 (N_5248,N_4684,N_4777);
and U5249 (N_5249,N_4523,N_4584);
nand U5250 (N_5250,N_4748,N_4601);
nor U5251 (N_5251,N_4959,N_4717);
nor U5252 (N_5252,N_4722,N_4639);
xor U5253 (N_5253,N_4954,N_4673);
nand U5254 (N_5254,N_4898,N_4651);
nand U5255 (N_5255,N_4810,N_4732);
nor U5256 (N_5256,N_4603,N_4665);
xnor U5257 (N_5257,N_4925,N_4850);
and U5258 (N_5258,N_4799,N_4967);
or U5259 (N_5259,N_4861,N_4611);
and U5260 (N_5260,N_4634,N_4971);
and U5261 (N_5261,N_4968,N_4832);
xor U5262 (N_5262,N_4910,N_4980);
nor U5263 (N_5263,N_4702,N_4600);
nor U5264 (N_5264,N_4678,N_4733);
nor U5265 (N_5265,N_4986,N_4602);
nand U5266 (N_5266,N_4845,N_4518);
or U5267 (N_5267,N_4735,N_4712);
and U5268 (N_5268,N_4566,N_4685);
nor U5269 (N_5269,N_4933,N_4905);
or U5270 (N_5270,N_4634,N_4998);
nor U5271 (N_5271,N_4843,N_4935);
xnor U5272 (N_5272,N_4914,N_4971);
xor U5273 (N_5273,N_4819,N_4693);
and U5274 (N_5274,N_4860,N_4535);
nor U5275 (N_5275,N_4806,N_4510);
nand U5276 (N_5276,N_4647,N_4729);
xnor U5277 (N_5277,N_4738,N_4965);
nor U5278 (N_5278,N_4567,N_4542);
nand U5279 (N_5279,N_4732,N_4870);
and U5280 (N_5280,N_4525,N_4906);
and U5281 (N_5281,N_4666,N_4860);
nand U5282 (N_5282,N_4956,N_4566);
and U5283 (N_5283,N_4809,N_4633);
or U5284 (N_5284,N_4758,N_4972);
nor U5285 (N_5285,N_4966,N_4595);
nor U5286 (N_5286,N_4585,N_4736);
and U5287 (N_5287,N_4554,N_4821);
and U5288 (N_5288,N_4890,N_4710);
and U5289 (N_5289,N_4765,N_4517);
or U5290 (N_5290,N_4976,N_4799);
or U5291 (N_5291,N_4916,N_4520);
nand U5292 (N_5292,N_4509,N_4561);
nand U5293 (N_5293,N_4745,N_4717);
and U5294 (N_5294,N_4688,N_4785);
and U5295 (N_5295,N_4825,N_4626);
or U5296 (N_5296,N_4667,N_4804);
and U5297 (N_5297,N_4761,N_4821);
and U5298 (N_5298,N_4900,N_4913);
and U5299 (N_5299,N_4505,N_4979);
nor U5300 (N_5300,N_4868,N_4726);
xnor U5301 (N_5301,N_4694,N_4678);
and U5302 (N_5302,N_4843,N_4544);
or U5303 (N_5303,N_4686,N_4868);
and U5304 (N_5304,N_4708,N_4786);
or U5305 (N_5305,N_4794,N_4979);
nor U5306 (N_5306,N_4576,N_4867);
nor U5307 (N_5307,N_4841,N_4972);
and U5308 (N_5308,N_4819,N_4716);
and U5309 (N_5309,N_4536,N_4921);
or U5310 (N_5310,N_4523,N_4723);
or U5311 (N_5311,N_4589,N_4787);
and U5312 (N_5312,N_4601,N_4679);
nor U5313 (N_5313,N_4527,N_4589);
xor U5314 (N_5314,N_4793,N_4881);
nor U5315 (N_5315,N_4917,N_4833);
nand U5316 (N_5316,N_4880,N_4969);
nand U5317 (N_5317,N_4864,N_4818);
nand U5318 (N_5318,N_4897,N_4613);
or U5319 (N_5319,N_4982,N_4929);
nand U5320 (N_5320,N_4601,N_4557);
nor U5321 (N_5321,N_4987,N_4824);
or U5322 (N_5322,N_4554,N_4764);
and U5323 (N_5323,N_4625,N_4554);
nand U5324 (N_5324,N_4618,N_4800);
nand U5325 (N_5325,N_4681,N_4720);
nor U5326 (N_5326,N_4645,N_4663);
nor U5327 (N_5327,N_4680,N_4756);
nand U5328 (N_5328,N_4749,N_4983);
and U5329 (N_5329,N_4980,N_4591);
nand U5330 (N_5330,N_4890,N_4931);
or U5331 (N_5331,N_4756,N_4551);
nand U5332 (N_5332,N_4558,N_4736);
nor U5333 (N_5333,N_4522,N_4524);
nor U5334 (N_5334,N_4971,N_4928);
and U5335 (N_5335,N_4712,N_4557);
or U5336 (N_5336,N_4746,N_4686);
nor U5337 (N_5337,N_4924,N_4610);
or U5338 (N_5338,N_4670,N_4591);
nor U5339 (N_5339,N_4747,N_4802);
or U5340 (N_5340,N_4904,N_4865);
and U5341 (N_5341,N_4880,N_4961);
or U5342 (N_5342,N_4660,N_4999);
nand U5343 (N_5343,N_4977,N_4691);
nand U5344 (N_5344,N_4596,N_4733);
nor U5345 (N_5345,N_4986,N_4941);
or U5346 (N_5346,N_4638,N_4602);
or U5347 (N_5347,N_4555,N_4661);
and U5348 (N_5348,N_4578,N_4519);
or U5349 (N_5349,N_4531,N_4925);
or U5350 (N_5350,N_4839,N_4753);
or U5351 (N_5351,N_4593,N_4666);
and U5352 (N_5352,N_4674,N_4528);
nor U5353 (N_5353,N_4532,N_4803);
or U5354 (N_5354,N_4584,N_4975);
nand U5355 (N_5355,N_4942,N_4565);
nor U5356 (N_5356,N_4653,N_4661);
nand U5357 (N_5357,N_4523,N_4830);
xnor U5358 (N_5358,N_4845,N_4649);
or U5359 (N_5359,N_4744,N_4964);
nor U5360 (N_5360,N_4585,N_4739);
nand U5361 (N_5361,N_4530,N_4612);
and U5362 (N_5362,N_4985,N_4578);
nand U5363 (N_5363,N_4573,N_4829);
nor U5364 (N_5364,N_4828,N_4695);
or U5365 (N_5365,N_4684,N_4946);
xor U5366 (N_5366,N_4749,N_4730);
and U5367 (N_5367,N_4704,N_4660);
nand U5368 (N_5368,N_4513,N_4542);
or U5369 (N_5369,N_4732,N_4505);
nor U5370 (N_5370,N_4599,N_4981);
nor U5371 (N_5371,N_4652,N_4721);
nand U5372 (N_5372,N_4860,N_4688);
or U5373 (N_5373,N_4666,N_4832);
nor U5374 (N_5374,N_4840,N_4831);
nand U5375 (N_5375,N_4580,N_4860);
and U5376 (N_5376,N_4543,N_4552);
nand U5377 (N_5377,N_4702,N_4555);
or U5378 (N_5378,N_4875,N_4707);
nor U5379 (N_5379,N_4591,N_4815);
nor U5380 (N_5380,N_4998,N_4718);
or U5381 (N_5381,N_4844,N_4993);
and U5382 (N_5382,N_4763,N_4565);
and U5383 (N_5383,N_4726,N_4675);
or U5384 (N_5384,N_4968,N_4882);
nor U5385 (N_5385,N_4974,N_4767);
or U5386 (N_5386,N_4828,N_4884);
or U5387 (N_5387,N_4818,N_4902);
nor U5388 (N_5388,N_4709,N_4623);
or U5389 (N_5389,N_4878,N_4592);
and U5390 (N_5390,N_4795,N_4833);
nor U5391 (N_5391,N_4771,N_4703);
or U5392 (N_5392,N_4912,N_4930);
nor U5393 (N_5393,N_4955,N_4542);
and U5394 (N_5394,N_4579,N_4861);
nand U5395 (N_5395,N_4660,N_4934);
or U5396 (N_5396,N_4572,N_4686);
nor U5397 (N_5397,N_4584,N_4621);
nand U5398 (N_5398,N_4593,N_4678);
nand U5399 (N_5399,N_4502,N_4571);
nor U5400 (N_5400,N_4536,N_4918);
xor U5401 (N_5401,N_4910,N_4659);
nand U5402 (N_5402,N_4881,N_4556);
or U5403 (N_5403,N_4651,N_4529);
or U5404 (N_5404,N_4845,N_4643);
nand U5405 (N_5405,N_4507,N_4790);
nor U5406 (N_5406,N_4643,N_4621);
nand U5407 (N_5407,N_4834,N_4969);
nand U5408 (N_5408,N_4913,N_4608);
or U5409 (N_5409,N_4706,N_4948);
or U5410 (N_5410,N_4817,N_4552);
nor U5411 (N_5411,N_4642,N_4858);
and U5412 (N_5412,N_4747,N_4698);
or U5413 (N_5413,N_4706,N_4934);
nor U5414 (N_5414,N_4826,N_4745);
xnor U5415 (N_5415,N_4529,N_4588);
nor U5416 (N_5416,N_4624,N_4541);
and U5417 (N_5417,N_4942,N_4730);
and U5418 (N_5418,N_4879,N_4858);
nor U5419 (N_5419,N_4913,N_4821);
nor U5420 (N_5420,N_4810,N_4806);
nor U5421 (N_5421,N_4916,N_4669);
nor U5422 (N_5422,N_4554,N_4575);
nand U5423 (N_5423,N_4914,N_4651);
and U5424 (N_5424,N_4932,N_4606);
nand U5425 (N_5425,N_4701,N_4968);
nand U5426 (N_5426,N_4934,N_4923);
nand U5427 (N_5427,N_4966,N_4897);
nand U5428 (N_5428,N_4681,N_4503);
nor U5429 (N_5429,N_4836,N_4799);
xor U5430 (N_5430,N_4833,N_4930);
nor U5431 (N_5431,N_4713,N_4593);
nand U5432 (N_5432,N_4593,N_4957);
or U5433 (N_5433,N_4589,N_4883);
nand U5434 (N_5434,N_4560,N_4679);
or U5435 (N_5435,N_4977,N_4811);
and U5436 (N_5436,N_4974,N_4512);
and U5437 (N_5437,N_4891,N_4934);
nor U5438 (N_5438,N_4779,N_4821);
nor U5439 (N_5439,N_4848,N_4906);
or U5440 (N_5440,N_4707,N_4823);
or U5441 (N_5441,N_4951,N_4976);
nor U5442 (N_5442,N_4959,N_4611);
nand U5443 (N_5443,N_4906,N_4791);
nor U5444 (N_5444,N_4540,N_4530);
nor U5445 (N_5445,N_4623,N_4659);
and U5446 (N_5446,N_4859,N_4895);
and U5447 (N_5447,N_4784,N_4772);
and U5448 (N_5448,N_4751,N_4788);
xnor U5449 (N_5449,N_4876,N_4730);
xor U5450 (N_5450,N_4877,N_4934);
nor U5451 (N_5451,N_4592,N_4797);
or U5452 (N_5452,N_4863,N_4833);
or U5453 (N_5453,N_4658,N_4600);
and U5454 (N_5454,N_4943,N_4628);
nand U5455 (N_5455,N_4876,N_4954);
nor U5456 (N_5456,N_4789,N_4514);
nor U5457 (N_5457,N_4814,N_4790);
or U5458 (N_5458,N_4552,N_4848);
and U5459 (N_5459,N_4959,N_4771);
and U5460 (N_5460,N_4523,N_4809);
and U5461 (N_5461,N_4735,N_4568);
or U5462 (N_5462,N_4578,N_4662);
or U5463 (N_5463,N_4646,N_4892);
or U5464 (N_5464,N_4804,N_4774);
xor U5465 (N_5465,N_4809,N_4685);
or U5466 (N_5466,N_4829,N_4844);
nand U5467 (N_5467,N_4707,N_4706);
nor U5468 (N_5468,N_4670,N_4586);
nor U5469 (N_5469,N_4526,N_4573);
nand U5470 (N_5470,N_4862,N_4566);
nor U5471 (N_5471,N_4812,N_4597);
nor U5472 (N_5472,N_4737,N_4929);
or U5473 (N_5473,N_4795,N_4955);
nor U5474 (N_5474,N_4524,N_4677);
or U5475 (N_5475,N_4926,N_4666);
nor U5476 (N_5476,N_4863,N_4949);
nor U5477 (N_5477,N_4602,N_4585);
nor U5478 (N_5478,N_4902,N_4574);
nor U5479 (N_5479,N_4612,N_4795);
and U5480 (N_5480,N_4996,N_4957);
and U5481 (N_5481,N_4540,N_4678);
and U5482 (N_5482,N_4955,N_4978);
and U5483 (N_5483,N_4573,N_4521);
or U5484 (N_5484,N_4530,N_4625);
and U5485 (N_5485,N_4687,N_4659);
or U5486 (N_5486,N_4783,N_4863);
nand U5487 (N_5487,N_4622,N_4568);
nand U5488 (N_5488,N_4858,N_4807);
or U5489 (N_5489,N_4653,N_4701);
and U5490 (N_5490,N_4716,N_4561);
xnor U5491 (N_5491,N_4804,N_4897);
nand U5492 (N_5492,N_4858,N_4848);
or U5493 (N_5493,N_4986,N_4623);
or U5494 (N_5494,N_4607,N_4941);
nor U5495 (N_5495,N_4520,N_4584);
xnor U5496 (N_5496,N_4682,N_4604);
or U5497 (N_5497,N_4728,N_4540);
or U5498 (N_5498,N_4605,N_4756);
or U5499 (N_5499,N_4769,N_4766);
or U5500 (N_5500,N_5471,N_5313);
and U5501 (N_5501,N_5261,N_5133);
nand U5502 (N_5502,N_5086,N_5426);
nand U5503 (N_5503,N_5135,N_5185);
or U5504 (N_5504,N_5168,N_5117);
nor U5505 (N_5505,N_5154,N_5397);
nor U5506 (N_5506,N_5083,N_5055);
nand U5507 (N_5507,N_5481,N_5267);
or U5508 (N_5508,N_5277,N_5102);
nand U5509 (N_5509,N_5349,N_5292);
or U5510 (N_5510,N_5177,N_5044);
nor U5511 (N_5511,N_5392,N_5434);
nand U5512 (N_5512,N_5061,N_5189);
nand U5513 (N_5513,N_5423,N_5028);
or U5514 (N_5514,N_5024,N_5370);
and U5515 (N_5515,N_5243,N_5458);
nor U5516 (N_5516,N_5163,N_5380);
and U5517 (N_5517,N_5118,N_5359);
and U5518 (N_5518,N_5202,N_5404);
or U5519 (N_5519,N_5220,N_5323);
or U5520 (N_5520,N_5057,N_5014);
or U5521 (N_5521,N_5005,N_5301);
nor U5522 (N_5522,N_5119,N_5222);
and U5523 (N_5523,N_5111,N_5475);
nor U5524 (N_5524,N_5469,N_5141);
nor U5525 (N_5525,N_5484,N_5258);
nand U5526 (N_5526,N_5023,N_5247);
xnor U5527 (N_5527,N_5081,N_5059);
nand U5528 (N_5528,N_5226,N_5113);
xor U5529 (N_5529,N_5476,N_5249);
nand U5530 (N_5530,N_5428,N_5071);
nor U5531 (N_5531,N_5215,N_5421);
nor U5532 (N_5532,N_5116,N_5329);
nand U5533 (N_5533,N_5418,N_5282);
nor U5534 (N_5534,N_5401,N_5008);
or U5535 (N_5535,N_5079,N_5333);
and U5536 (N_5536,N_5422,N_5228);
nand U5537 (N_5537,N_5097,N_5459);
and U5538 (N_5538,N_5046,N_5159);
nor U5539 (N_5539,N_5026,N_5120);
or U5540 (N_5540,N_5191,N_5307);
or U5541 (N_5541,N_5439,N_5407);
xnor U5542 (N_5542,N_5085,N_5472);
and U5543 (N_5543,N_5410,N_5477);
nor U5544 (N_5544,N_5390,N_5101);
nand U5545 (N_5545,N_5293,N_5264);
or U5546 (N_5546,N_5236,N_5321);
nand U5547 (N_5547,N_5088,N_5033);
and U5548 (N_5548,N_5002,N_5021);
nor U5549 (N_5549,N_5200,N_5164);
and U5550 (N_5550,N_5027,N_5308);
and U5551 (N_5551,N_5263,N_5336);
xor U5552 (N_5552,N_5140,N_5447);
nor U5553 (N_5553,N_5208,N_5373);
xnor U5554 (N_5554,N_5232,N_5411);
nand U5555 (N_5555,N_5365,N_5035);
nand U5556 (N_5556,N_5181,N_5147);
or U5557 (N_5557,N_5468,N_5358);
nand U5558 (N_5558,N_5280,N_5291);
or U5559 (N_5559,N_5092,N_5248);
and U5560 (N_5560,N_5417,N_5340);
nor U5561 (N_5561,N_5317,N_5433);
nor U5562 (N_5562,N_5091,N_5063);
and U5563 (N_5563,N_5151,N_5099);
nor U5564 (N_5564,N_5188,N_5309);
and U5565 (N_5565,N_5138,N_5001);
or U5566 (N_5566,N_5462,N_5209);
nor U5567 (N_5567,N_5204,N_5074);
xor U5568 (N_5568,N_5363,N_5003);
xnor U5569 (N_5569,N_5430,N_5213);
nand U5570 (N_5570,N_5326,N_5461);
nand U5571 (N_5571,N_5338,N_5446);
xnor U5572 (N_5572,N_5406,N_5227);
nor U5573 (N_5573,N_5094,N_5371);
nand U5574 (N_5574,N_5318,N_5056);
nor U5575 (N_5575,N_5274,N_5327);
nor U5576 (N_5576,N_5155,N_5105);
nand U5577 (N_5577,N_5123,N_5219);
nand U5578 (N_5578,N_5252,N_5286);
and U5579 (N_5579,N_5230,N_5429);
nor U5580 (N_5580,N_5069,N_5302);
or U5581 (N_5581,N_5259,N_5078);
nand U5582 (N_5582,N_5018,N_5443);
or U5583 (N_5583,N_5491,N_5171);
or U5584 (N_5584,N_5000,N_5130);
nand U5585 (N_5585,N_5045,N_5495);
nand U5586 (N_5586,N_5343,N_5207);
and U5587 (N_5587,N_5284,N_5285);
or U5588 (N_5588,N_5173,N_5149);
and U5589 (N_5589,N_5438,N_5346);
nor U5590 (N_5590,N_5187,N_5211);
nor U5591 (N_5591,N_5038,N_5129);
nand U5592 (N_5592,N_5052,N_5474);
or U5593 (N_5593,N_5250,N_5420);
nand U5594 (N_5594,N_5290,N_5360);
nand U5595 (N_5595,N_5466,N_5150);
or U5596 (N_5596,N_5139,N_5229);
xnor U5597 (N_5597,N_5016,N_5455);
nand U5598 (N_5598,N_5391,N_5270);
nor U5599 (N_5599,N_5496,N_5375);
nor U5600 (N_5600,N_5499,N_5331);
nor U5601 (N_5601,N_5362,N_5294);
or U5602 (N_5602,N_5271,N_5453);
xor U5603 (N_5603,N_5178,N_5409);
nor U5604 (N_5604,N_5257,N_5497);
and U5605 (N_5605,N_5265,N_5479);
nand U5606 (N_5606,N_5276,N_5457);
nand U5607 (N_5607,N_5167,N_5442);
or U5608 (N_5608,N_5166,N_5186);
nand U5609 (N_5609,N_5009,N_5395);
nand U5610 (N_5610,N_5075,N_5169);
nand U5611 (N_5611,N_5233,N_5393);
nor U5612 (N_5612,N_5482,N_5337);
or U5613 (N_5613,N_5054,N_5494);
and U5614 (N_5614,N_5451,N_5214);
nor U5615 (N_5615,N_5488,N_5047);
nand U5616 (N_5616,N_5049,N_5379);
xor U5617 (N_5617,N_5398,N_5234);
or U5618 (N_5618,N_5153,N_5165);
and U5619 (N_5619,N_5156,N_5152);
and U5620 (N_5620,N_5432,N_5192);
or U5621 (N_5621,N_5203,N_5256);
nor U5622 (N_5622,N_5062,N_5416);
nand U5623 (N_5623,N_5053,N_5449);
or U5624 (N_5624,N_5126,N_5316);
nor U5625 (N_5625,N_5435,N_5060);
and U5626 (N_5626,N_5223,N_5311);
or U5627 (N_5627,N_5090,N_5067);
or U5628 (N_5628,N_5383,N_5394);
nor U5629 (N_5629,N_5448,N_5431);
nand U5630 (N_5630,N_5465,N_5082);
or U5631 (N_5631,N_5369,N_5115);
nor U5632 (N_5632,N_5201,N_5224);
nor U5633 (N_5633,N_5344,N_5172);
nor U5634 (N_5634,N_5436,N_5158);
xor U5635 (N_5635,N_5254,N_5255);
or U5636 (N_5636,N_5412,N_5070);
and U5637 (N_5637,N_5405,N_5251);
nand U5638 (N_5638,N_5402,N_5330);
nor U5639 (N_5639,N_5460,N_5351);
xnor U5640 (N_5640,N_5015,N_5098);
xnor U5641 (N_5641,N_5493,N_5235);
nand U5642 (N_5642,N_5040,N_5095);
and U5643 (N_5643,N_5419,N_5287);
nand U5644 (N_5644,N_5314,N_5399);
nand U5645 (N_5645,N_5174,N_5332);
or U5646 (N_5646,N_5288,N_5361);
nand U5647 (N_5647,N_5010,N_5176);
xor U5648 (N_5648,N_5478,N_5198);
xnor U5649 (N_5649,N_5354,N_5162);
nor U5650 (N_5650,N_5041,N_5144);
or U5651 (N_5651,N_5073,N_5048);
nand U5652 (N_5652,N_5065,N_5304);
nand U5653 (N_5653,N_5456,N_5022);
xor U5654 (N_5654,N_5142,N_5483);
or U5655 (N_5655,N_5029,N_5058);
nand U5656 (N_5656,N_5128,N_5414);
xnor U5657 (N_5657,N_5148,N_5100);
or U5658 (N_5658,N_5020,N_5143);
or U5659 (N_5659,N_5110,N_5145);
nor U5660 (N_5660,N_5011,N_5076);
or U5661 (N_5661,N_5160,N_5295);
nand U5662 (N_5662,N_5444,N_5357);
or U5663 (N_5663,N_5352,N_5413);
and U5664 (N_5664,N_5454,N_5384);
nor U5665 (N_5665,N_5103,N_5463);
and U5666 (N_5666,N_5096,N_5134);
and U5667 (N_5667,N_5347,N_5108);
nand U5668 (N_5668,N_5231,N_5467);
or U5669 (N_5669,N_5218,N_5328);
xor U5670 (N_5670,N_5199,N_5266);
nor U5671 (N_5671,N_5272,N_5210);
nor U5672 (N_5672,N_5368,N_5170);
and U5673 (N_5673,N_5425,N_5107);
or U5674 (N_5674,N_5132,N_5437);
and U5675 (N_5675,N_5193,N_5385);
and U5676 (N_5676,N_5281,N_5335);
nor U5677 (N_5677,N_5137,N_5279);
or U5678 (N_5678,N_5216,N_5424);
nand U5679 (N_5679,N_5364,N_5068);
xnor U5680 (N_5680,N_5205,N_5486);
and U5681 (N_5681,N_5030,N_5310);
or U5682 (N_5682,N_5339,N_5382);
and U5683 (N_5683,N_5260,N_5366);
and U5684 (N_5684,N_5031,N_5253);
nor U5685 (N_5685,N_5037,N_5353);
nand U5686 (N_5686,N_5025,N_5464);
nor U5687 (N_5687,N_5066,N_5374);
xnor U5688 (N_5688,N_5355,N_5064);
nand U5689 (N_5689,N_5470,N_5007);
nand U5690 (N_5690,N_5125,N_5182);
and U5691 (N_5691,N_5445,N_5093);
nand U5692 (N_5692,N_5017,N_5403);
nand U5693 (N_5693,N_5322,N_5190);
or U5694 (N_5694,N_5032,N_5378);
nor U5695 (N_5695,N_5320,N_5319);
xnor U5696 (N_5696,N_5376,N_5237);
and U5697 (N_5697,N_5034,N_5341);
nand U5698 (N_5698,N_5089,N_5273);
xnor U5699 (N_5699,N_5489,N_5342);
nor U5700 (N_5700,N_5124,N_5131);
and U5701 (N_5701,N_5473,N_5206);
nand U5702 (N_5702,N_5408,N_5427);
nor U5703 (N_5703,N_5112,N_5241);
or U5704 (N_5704,N_5487,N_5240);
nand U5705 (N_5705,N_5051,N_5400);
or U5706 (N_5706,N_5183,N_5136);
nor U5707 (N_5707,N_5104,N_5396);
nor U5708 (N_5708,N_5345,N_5013);
or U5709 (N_5709,N_5036,N_5109);
xnor U5710 (N_5710,N_5221,N_5283);
or U5711 (N_5711,N_5324,N_5387);
nand U5712 (N_5712,N_5268,N_5196);
nor U5713 (N_5713,N_5122,N_5498);
nand U5714 (N_5714,N_5441,N_5386);
and U5715 (N_5715,N_5072,N_5296);
nor U5716 (N_5716,N_5305,N_5043);
nand U5717 (N_5717,N_5480,N_5452);
or U5718 (N_5718,N_5179,N_5275);
or U5719 (N_5719,N_5157,N_5300);
or U5720 (N_5720,N_5242,N_5348);
or U5721 (N_5721,N_5303,N_5377);
nor U5722 (N_5722,N_5175,N_5244);
nand U5723 (N_5723,N_5440,N_5197);
nand U5724 (N_5724,N_5004,N_5356);
or U5725 (N_5725,N_5325,N_5050);
nor U5726 (N_5726,N_5012,N_5299);
or U5727 (N_5727,N_5087,N_5084);
nand U5728 (N_5728,N_5127,N_5121);
nand U5729 (N_5729,N_5312,N_5306);
nor U5730 (N_5730,N_5350,N_5315);
and U5731 (N_5731,N_5217,N_5246);
nor U5732 (N_5732,N_5238,N_5006);
or U5733 (N_5733,N_5042,N_5184);
and U5734 (N_5734,N_5114,N_5080);
and U5735 (N_5735,N_5225,N_5146);
or U5736 (N_5736,N_5297,N_5077);
nand U5737 (N_5737,N_5490,N_5239);
nand U5738 (N_5738,N_5289,N_5372);
or U5739 (N_5739,N_5278,N_5388);
xor U5740 (N_5740,N_5106,N_5019);
or U5741 (N_5741,N_5194,N_5161);
or U5742 (N_5742,N_5381,N_5450);
nor U5743 (N_5743,N_5334,N_5367);
or U5744 (N_5744,N_5485,N_5269);
and U5745 (N_5745,N_5039,N_5415);
nand U5746 (N_5746,N_5195,N_5212);
nor U5747 (N_5747,N_5245,N_5492);
xnor U5748 (N_5748,N_5180,N_5298);
and U5749 (N_5749,N_5262,N_5389);
and U5750 (N_5750,N_5196,N_5286);
or U5751 (N_5751,N_5134,N_5058);
nand U5752 (N_5752,N_5203,N_5387);
nor U5753 (N_5753,N_5039,N_5133);
nor U5754 (N_5754,N_5285,N_5311);
nor U5755 (N_5755,N_5141,N_5042);
or U5756 (N_5756,N_5225,N_5283);
or U5757 (N_5757,N_5435,N_5059);
xnor U5758 (N_5758,N_5423,N_5072);
nor U5759 (N_5759,N_5006,N_5333);
nor U5760 (N_5760,N_5106,N_5256);
nand U5761 (N_5761,N_5075,N_5298);
and U5762 (N_5762,N_5161,N_5136);
nand U5763 (N_5763,N_5010,N_5073);
or U5764 (N_5764,N_5273,N_5040);
and U5765 (N_5765,N_5300,N_5081);
and U5766 (N_5766,N_5212,N_5457);
and U5767 (N_5767,N_5380,N_5111);
or U5768 (N_5768,N_5315,N_5401);
nor U5769 (N_5769,N_5451,N_5424);
nand U5770 (N_5770,N_5423,N_5382);
nand U5771 (N_5771,N_5255,N_5234);
or U5772 (N_5772,N_5080,N_5243);
nor U5773 (N_5773,N_5431,N_5338);
or U5774 (N_5774,N_5405,N_5141);
nor U5775 (N_5775,N_5048,N_5388);
nor U5776 (N_5776,N_5257,N_5170);
or U5777 (N_5777,N_5143,N_5436);
nand U5778 (N_5778,N_5363,N_5128);
nand U5779 (N_5779,N_5015,N_5287);
nor U5780 (N_5780,N_5311,N_5195);
nand U5781 (N_5781,N_5377,N_5457);
nor U5782 (N_5782,N_5446,N_5229);
or U5783 (N_5783,N_5398,N_5030);
nor U5784 (N_5784,N_5057,N_5100);
and U5785 (N_5785,N_5017,N_5067);
xnor U5786 (N_5786,N_5169,N_5209);
nand U5787 (N_5787,N_5294,N_5093);
or U5788 (N_5788,N_5434,N_5195);
xor U5789 (N_5789,N_5063,N_5343);
nor U5790 (N_5790,N_5465,N_5036);
or U5791 (N_5791,N_5267,N_5373);
or U5792 (N_5792,N_5180,N_5142);
xor U5793 (N_5793,N_5264,N_5396);
nor U5794 (N_5794,N_5331,N_5246);
or U5795 (N_5795,N_5178,N_5487);
and U5796 (N_5796,N_5478,N_5494);
nor U5797 (N_5797,N_5149,N_5486);
or U5798 (N_5798,N_5020,N_5376);
or U5799 (N_5799,N_5347,N_5006);
and U5800 (N_5800,N_5394,N_5376);
nor U5801 (N_5801,N_5365,N_5445);
nand U5802 (N_5802,N_5102,N_5183);
nand U5803 (N_5803,N_5452,N_5158);
or U5804 (N_5804,N_5313,N_5213);
or U5805 (N_5805,N_5135,N_5281);
or U5806 (N_5806,N_5064,N_5053);
and U5807 (N_5807,N_5230,N_5409);
or U5808 (N_5808,N_5341,N_5356);
and U5809 (N_5809,N_5076,N_5356);
nor U5810 (N_5810,N_5409,N_5281);
nand U5811 (N_5811,N_5330,N_5001);
or U5812 (N_5812,N_5481,N_5499);
nor U5813 (N_5813,N_5414,N_5231);
nor U5814 (N_5814,N_5029,N_5199);
nand U5815 (N_5815,N_5346,N_5453);
and U5816 (N_5816,N_5283,N_5415);
xor U5817 (N_5817,N_5149,N_5125);
and U5818 (N_5818,N_5209,N_5217);
nor U5819 (N_5819,N_5273,N_5177);
nor U5820 (N_5820,N_5411,N_5240);
xor U5821 (N_5821,N_5483,N_5205);
nand U5822 (N_5822,N_5283,N_5220);
nor U5823 (N_5823,N_5154,N_5421);
nor U5824 (N_5824,N_5283,N_5310);
nor U5825 (N_5825,N_5293,N_5087);
nand U5826 (N_5826,N_5035,N_5354);
nor U5827 (N_5827,N_5328,N_5272);
or U5828 (N_5828,N_5149,N_5226);
nor U5829 (N_5829,N_5429,N_5327);
nand U5830 (N_5830,N_5338,N_5334);
nor U5831 (N_5831,N_5227,N_5476);
nor U5832 (N_5832,N_5469,N_5045);
or U5833 (N_5833,N_5482,N_5292);
nand U5834 (N_5834,N_5471,N_5144);
or U5835 (N_5835,N_5302,N_5136);
nand U5836 (N_5836,N_5217,N_5052);
xor U5837 (N_5837,N_5236,N_5170);
xnor U5838 (N_5838,N_5068,N_5267);
or U5839 (N_5839,N_5423,N_5207);
and U5840 (N_5840,N_5334,N_5163);
or U5841 (N_5841,N_5354,N_5427);
xnor U5842 (N_5842,N_5045,N_5109);
nor U5843 (N_5843,N_5168,N_5489);
or U5844 (N_5844,N_5486,N_5188);
and U5845 (N_5845,N_5480,N_5155);
nand U5846 (N_5846,N_5276,N_5362);
and U5847 (N_5847,N_5335,N_5290);
nand U5848 (N_5848,N_5079,N_5167);
nand U5849 (N_5849,N_5055,N_5360);
nand U5850 (N_5850,N_5028,N_5133);
xnor U5851 (N_5851,N_5135,N_5410);
nor U5852 (N_5852,N_5290,N_5143);
and U5853 (N_5853,N_5285,N_5324);
or U5854 (N_5854,N_5258,N_5365);
xor U5855 (N_5855,N_5427,N_5404);
or U5856 (N_5856,N_5001,N_5300);
nand U5857 (N_5857,N_5376,N_5171);
nand U5858 (N_5858,N_5442,N_5260);
or U5859 (N_5859,N_5175,N_5015);
xnor U5860 (N_5860,N_5207,N_5183);
nor U5861 (N_5861,N_5291,N_5307);
and U5862 (N_5862,N_5169,N_5314);
or U5863 (N_5863,N_5233,N_5477);
or U5864 (N_5864,N_5459,N_5146);
nand U5865 (N_5865,N_5040,N_5461);
nand U5866 (N_5866,N_5025,N_5098);
or U5867 (N_5867,N_5104,N_5395);
or U5868 (N_5868,N_5148,N_5166);
xor U5869 (N_5869,N_5044,N_5383);
nand U5870 (N_5870,N_5452,N_5342);
xor U5871 (N_5871,N_5418,N_5013);
and U5872 (N_5872,N_5449,N_5005);
and U5873 (N_5873,N_5042,N_5316);
or U5874 (N_5874,N_5051,N_5093);
nor U5875 (N_5875,N_5371,N_5364);
nor U5876 (N_5876,N_5454,N_5069);
or U5877 (N_5877,N_5006,N_5044);
or U5878 (N_5878,N_5307,N_5240);
or U5879 (N_5879,N_5469,N_5117);
or U5880 (N_5880,N_5164,N_5363);
xnor U5881 (N_5881,N_5333,N_5059);
or U5882 (N_5882,N_5306,N_5361);
nor U5883 (N_5883,N_5145,N_5026);
nand U5884 (N_5884,N_5161,N_5476);
nand U5885 (N_5885,N_5498,N_5000);
nand U5886 (N_5886,N_5437,N_5199);
and U5887 (N_5887,N_5469,N_5331);
nor U5888 (N_5888,N_5385,N_5148);
nor U5889 (N_5889,N_5382,N_5324);
and U5890 (N_5890,N_5157,N_5211);
xnor U5891 (N_5891,N_5486,N_5329);
nor U5892 (N_5892,N_5415,N_5238);
nor U5893 (N_5893,N_5314,N_5197);
and U5894 (N_5894,N_5387,N_5148);
nand U5895 (N_5895,N_5347,N_5329);
nor U5896 (N_5896,N_5274,N_5013);
nand U5897 (N_5897,N_5228,N_5039);
nand U5898 (N_5898,N_5131,N_5112);
nand U5899 (N_5899,N_5358,N_5433);
nor U5900 (N_5900,N_5374,N_5499);
nand U5901 (N_5901,N_5394,N_5283);
or U5902 (N_5902,N_5467,N_5109);
nand U5903 (N_5903,N_5464,N_5287);
nor U5904 (N_5904,N_5060,N_5392);
nor U5905 (N_5905,N_5366,N_5006);
nand U5906 (N_5906,N_5165,N_5362);
or U5907 (N_5907,N_5439,N_5078);
and U5908 (N_5908,N_5461,N_5310);
nor U5909 (N_5909,N_5003,N_5405);
and U5910 (N_5910,N_5033,N_5237);
or U5911 (N_5911,N_5023,N_5326);
nor U5912 (N_5912,N_5161,N_5441);
or U5913 (N_5913,N_5281,N_5305);
nor U5914 (N_5914,N_5079,N_5027);
nand U5915 (N_5915,N_5122,N_5108);
nand U5916 (N_5916,N_5198,N_5237);
nand U5917 (N_5917,N_5149,N_5143);
and U5918 (N_5918,N_5234,N_5465);
nand U5919 (N_5919,N_5059,N_5296);
nor U5920 (N_5920,N_5334,N_5063);
or U5921 (N_5921,N_5255,N_5271);
nor U5922 (N_5922,N_5093,N_5057);
nand U5923 (N_5923,N_5029,N_5178);
or U5924 (N_5924,N_5269,N_5341);
nand U5925 (N_5925,N_5417,N_5056);
and U5926 (N_5926,N_5054,N_5419);
nor U5927 (N_5927,N_5157,N_5030);
nor U5928 (N_5928,N_5161,N_5331);
or U5929 (N_5929,N_5088,N_5282);
xor U5930 (N_5930,N_5449,N_5155);
nor U5931 (N_5931,N_5387,N_5394);
and U5932 (N_5932,N_5101,N_5301);
or U5933 (N_5933,N_5112,N_5163);
xor U5934 (N_5934,N_5259,N_5032);
nand U5935 (N_5935,N_5420,N_5252);
and U5936 (N_5936,N_5381,N_5118);
nor U5937 (N_5937,N_5380,N_5090);
or U5938 (N_5938,N_5012,N_5001);
nor U5939 (N_5939,N_5465,N_5351);
and U5940 (N_5940,N_5467,N_5074);
nand U5941 (N_5941,N_5045,N_5471);
xor U5942 (N_5942,N_5249,N_5363);
nand U5943 (N_5943,N_5143,N_5014);
and U5944 (N_5944,N_5242,N_5394);
nand U5945 (N_5945,N_5031,N_5402);
and U5946 (N_5946,N_5367,N_5050);
or U5947 (N_5947,N_5359,N_5122);
and U5948 (N_5948,N_5410,N_5096);
or U5949 (N_5949,N_5018,N_5340);
xnor U5950 (N_5950,N_5039,N_5197);
or U5951 (N_5951,N_5011,N_5136);
nor U5952 (N_5952,N_5365,N_5312);
xor U5953 (N_5953,N_5335,N_5025);
nand U5954 (N_5954,N_5368,N_5291);
nor U5955 (N_5955,N_5301,N_5209);
nor U5956 (N_5956,N_5196,N_5078);
or U5957 (N_5957,N_5464,N_5042);
nand U5958 (N_5958,N_5396,N_5175);
nand U5959 (N_5959,N_5379,N_5155);
nor U5960 (N_5960,N_5353,N_5494);
or U5961 (N_5961,N_5320,N_5436);
and U5962 (N_5962,N_5018,N_5254);
or U5963 (N_5963,N_5262,N_5336);
nor U5964 (N_5964,N_5267,N_5302);
xnor U5965 (N_5965,N_5162,N_5380);
nor U5966 (N_5966,N_5035,N_5352);
or U5967 (N_5967,N_5080,N_5255);
or U5968 (N_5968,N_5047,N_5439);
and U5969 (N_5969,N_5110,N_5313);
nor U5970 (N_5970,N_5433,N_5212);
or U5971 (N_5971,N_5129,N_5101);
nor U5972 (N_5972,N_5379,N_5380);
nand U5973 (N_5973,N_5115,N_5456);
nand U5974 (N_5974,N_5096,N_5442);
nor U5975 (N_5975,N_5210,N_5434);
nor U5976 (N_5976,N_5187,N_5283);
or U5977 (N_5977,N_5203,N_5289);
nor U5978 (N_5978,N_5220,N_5231);
nor U5979 (N_5979,N_5258,N_5438);
and U5980 (N_5980,N_5384,N_5292);
and U5981 (N_5981,N_5341,N_5066);
nor U5982 (N_5982,N_5144,N_5125);
or U5983 (N_5983,N_5180,N_5090);
or U5984 (N_5984,N_5499,N_5326);
nor U5985 (N_5985,N_5498,N_5302);
xnor U5986 (N_5986,N_5485,N_5096);
nor U5987 (N_5987,N_5216,N_5255);
and U5988 (N_5988,N_5251,N_5100);
and U5989 (N_5989,N_5023,N_5441);
nor U5990 (N_5990,N_5155,N_5222);
and U5991 (N_5991,N_5322,N_5367);
nor U5992 (N_5992,N_5092,N_5478);
and U5993 (N_5993,N_5360,N_5449);
xor U5994 (N_5994,N_5341,N_5076);
nand U5995 (N_5995,N_5417,N_5467);
or U5996 (N_5996,N_5222,N_5446);
nand U5997 (N_5997,N_5492,N_5175);
or U5998 (N_5998,N_5494,N_5154);
nor U5999 (N_5999,N_5364,N_5338);
and U6000 (N_6000,N_5653,N_5805);
or U6001 (N_6001,N_5713,N_5665);
nand U6002 (N_6002,N_5877,N_5558);
or U6003 (N_6003,N_5998,N_5857);
nor U6004 (N_6004,N_5548,N_5594);
xnor U6005 (N_6005,N_5528,N_5911);
xor U6006 (N_6006,N_5979,N_5975);
or U6007 (N_6007,N_5677,N_5702);
and U6008 (N_6008,N_5917,N_5918);
xnor U6009 (N_6009,N_5899,N_5790);
nand U6010 (N_6010,N_5572,N_5988);
xnor U6011 (N_6011,N_5934,N_5871);
nor U6012 (N_6012,N_5815,N_5648);
and U6013 (N_6013,N_5534,N_5681);
nor U6014 (N_6014,N_5808,N_5818);
xnor U6015 (N_6015,N_5506,N_5848);
nor U6016 (N_6016,N_5726,N_5944);
and U6017 (N_6017,N_5872,N_5601);
and U6018 (N_6018,N_5524,N_5959);
nand U6019 (N_6019,N_5755,N_5650);
nor U6020 (N_6020,N_5887,N_5651);
or U6021 (N_6021,N_5974,N_5616);
or U6022 (N_6022,N_5747,N_5763);
xnor U6023 (N_6023,N_5622,N_5728);
or U6024 (N_6024,N_5860,N_5811);
and U6025 (N_6025,N_5845,N_5893);
and U6026 (N_6026,N_5641,N_5654);
xor U6027 (N_6027,N_5715,N_5853);
and U6028 (N_6028,N_5706,N_5787);
nand U6029 (N_6029,N_5664,N_5637);
nand U6030 (N_6030,N_5926,N_5510);
nand U6031 (N_6031,N_5519,N_5813);
or U6032 (N_6032,N_5631,N_5780);
nand U6033 (N_6033,N_5957,N_5769);
nand U6034 (N_6034,N_5810,N_5609);
nand U6035 (N_6035,N_5547,N_5846);
nand U6036 (N_6036,N_5670,N_5858);
and U6037 (N_6037,N_5717,N_5646);
and U6038 (N_6038,N_5723,N_5643);
and U6039 (N_6039,N_5603,N_5590);
xnor U6040 (N_6040,N_5898,N_5718);
nand U6041 (N_6041,N_5844,N_5593);
or U6042 (N_6042,N_5686,N_5995);
nand U6043 (N_6043,N_5512,N_5869);
nor U6044 (N_6044,N_5972,N_5910);
nand U6045 (N_6045,N_5854,N_5950);
or U6046 (N_6046,N_5970,N_5765);
and U6047 (N_6047,N_5913,N_5921);
or U6048 (N_6048,N_5838,N_5938);
xor U6049 (N_6049,N_5701,N_5573);
or U6050 (N_6050,N_5612,N_5965);
or U6051 (N_6051,N_5835,N_5564);
nand U6052 (N_6052,N_5630,N_5855);
nand U6053 (N_6053,N_5733,N_5731);
and U6054 (N_6054,N_5884,N_5748);
or U6055 (N_6055,N_5782,N_5909);
nor U6056 (N_6056,N_5864,N_5736);
xnor U6057 (N_6057,N_5929,N_5674);
or U6058 (N_6058,N_5649,N_5513);
or U6059 (N_6059,N_5978,N_5508);
or U6060 (N_6060,N_5742,N_5840);
nor U6061 (N_6061,N_5746,N_5941);
and U6062 (N_6062,N_5891,N_5894);
or U6063 (N_6063,N_5886,N_5541);
and U6064 (N_6064,N_5740,N_5791);
and U6065 (N_6065,N_5623,N_5669);
or U6066 (N_6066,N_5737,N_5596);
and U6067 (N_6067,N_5850,N_5682);
nor U6068 (N_6068,N_5885,N_5947);
or U6069 (N_6069,N_5517,N_5831);
or U6070 (N_6070,N_5936,N_5614);
nand U6071 (N_6071,N_5552,N_5916);
and U6072 (N_6072,N_5764,N_5667);
nor U6073 (N_6073,N_5565,N_5536);
nor U6074 (N_6074,N_5684,N_5874);
nand U6075 (N_6075,N_5833,N_5961);
and U6076 (N_6076,N_5793,N_5656);
or U6077 (N_6077,N_5559,N_5621);
and U6078 (N_6078,N_5561,N_5505);
nand U6079 (N_6079,N_5930,N_5977);
and U6080 (N_6080,N_5618,N_5819);
or U6081 (N_6081,N_5696,N_5515);
or U6082 (N_6082,N_5583,N_5673);
xnor U6083 (N_6083,N_5504,N_5946);
or U6084 (N_6084,N_5925,N_5849);
nor U6085 (N_6085,N_5535,N_5927);
nor U6086 (N_6086,N_5794,N_5514);
nor U6087 (N_6087,N_5908,N_5915);
nor U6088 (N_6088,N_5557,N_5923);
or U6089 (N_6089,N_5716,N_5830);
nand U6090 (N_6090,N_5628,N_5645);
and U6091 (N_6091,N_5705,N_5574);
nand U6092 (N_6092,N_5738,N_5700);
nand U6093 (N_6093,N_5903,N_5962);
nor U6094 (N_6094,N_5620,N_5779);
and U6095 (N_6095,N_5757,N_5642);
or U6096 (N_6096,N_5671,N_5803);
and U6097 (N_6097,N_5533,N_5553);
and U6098 (N_6098,N_5735,N_5501);
and U6099 (N_6099,N_5841,N_5963);
nand U6100 (N_6100,N_5598,N_5729);
nor U6101 (N_6101,N_5525,N_5602);
nor U6102 (N_6102,N_5710,N_5861);
and U6103 (N_6103,N_5798,N_5543);
and U6104 (N_6104,N_5683,N_5968);
nor U6105 (N_6105,N_5532,N_5586);
and U6106 (N_6106,N_5719,N_5741);
nor U6107 (N_6107,N_5568,N_5924);
nor U6108 (N_6108,N_5881,N_5912);
or U6109 (N_6109,N_5580,N_5599);
and U6110 (N_6110,N_5851,N_5986);
xnor U6111 (N_6111,N_5588,N_5821);
or U6112 (N_6112,N_5743,N_5807);
nor U6113 (N_6113,N_5822,N_5999);
nand U6114 (N_6114,N_5906,N_5942);
nand U6115 (N_6115,N_5816,N_5868);
nand U6116 (N_6116,N_5870,N_5775);
nand U6117 (N_6117,N_5672,N_5966);
nor U6118 (N_6118,N_5953,N_5576);
and U6119 (N_6119,N_5920,N_5949);
xor U6120 (N_6120,N_5866,N_5889);
and U6121 (N_6121,N_5617,N_5919);
xor U6122 (N_6122,N_5652,N_5638);
nand U6123 (N_6123,N_5882,N_5973);
nor U6124 (N_6124,N_5875,N_5661);
nand U6125 (N_6125,N_5933,N_5626);
xor U6126 (N_6126,N_5992,N_5577);
or U6127 (N_6127,N_5571,N_5823);
and U6128 (N_6128,N_5876,N_5595);
nand U6129 (N_6129,N_5592,N_5507);
and U6130 (N_6130,N_5640,N_5502);
xor U6131 (N_6131,N_5636,N_5827);
or U6132 (N_6132,N_5660,N_5619);
and U6133 (N_6133,N_5680,N_5605);
nand U6134 (N_6134,N_5967,N_5629);
and U6135 (N_6135,N_5768,N_5767);
and U6136 (N_6136,N_5549,N_5806);
nor U6137 (N_6137,N_5801,N_5523);
nor U6138 (N_6138,N_5996,N_5878);
nor U6139 (N_6139,N_5985,N_5778);
and U6140 (N_6140,N_5714,N_5948);
or U6141 (N_6141,N_5809,N_5792);
nor U6142 (N_6142,N_5896,N_5865);
nand U6143 (N_6143,N_5550,N_5624);
and U6144 (N_6144,N_5759,N_5607);
or U6145 (N_6145,N_5703,N_5522);
nand U6146 (N_6146,N_5707,N_5608);
xnor U6147 (N_6147,N_5538,N_5509);
and U6148 (N_6148,N_5783,N_5597);
nand U6149 (N_6149,N_5632,N_5964);
nand U6150 (N_6150,N_5732,N_5969);
nor U6151 (N_6151,N_5774,N_5812);
or U6152 (N_6152,N_5863,N_5951);
and U6153 (N_6153,N_5799,N_5862);
or U6154 (N_6154,N_5545,N_5982);
and U6155 (N_6155,N_5721,N_5634);
nand U6156 (N_6156,N_5540,N_5688);
or U6157 (N_6157,N_5633,N_5575);
or U6158 (N_6158,N_5606,N_5754);
nor U6159 (N_6159,N_5907,N_5697);
and U6160 (N_6160,N_5687,N_5668);
and U6161 (N_6161,N_5569,N_5613);
nand U6162 (N_6162,N_5730,N_5960);
nor U6163 (N_6163,N_5635,N_5584);
or U6164 (N_6164,N_5530,N_5750);
nand U6165 (N_6165,N_5901,N_5773);
xnor U6166 (N_6166,N_5712,N_5727);
nor U6167 (N_6167,N_5954,N_5711);
and U6168 (N_6168,N_5647,N_5662);
nor U6169 (N_6169,N_5983,N_5679);
or U6170 (N_6170,N_5837,N_5879);
nand U6171 (N_6171,N_5663,N_5758);
nor U6172 (N_6172,N_5981,N_5788);
and U6173 (N_6173,N_5658,N_5867);
and U6174 (N_6174,N_5826,N_5690);
or U6175 (N_6175,N_5900,N_5824);
nand U6176 (N_6176,N_5776,N_5888);
nand U6177 (N_6177,N_5698,N_5956);
and U6178 (N_6178,N_5675,N_5852);
and U6179 (N_6179,N_5520,N_5814);
or U6180 (N_6180,N_5937,N_5739);
xnor U6181 (N_6181,N_5709,N_5760);
nand U6182 (N_6182,N_5828,N_5989);
or U6183 (N_6183,N_5804,N_5579);
and U6184 (N_6184,N_5753,N_5581);
and U6185 (N_6185,N_5611,N_5516);
nor U6186 (N_6186,N_5722,N_5699);
and U6187 (N_6187,N_5980,N_5749);
xnor U6188 (N_6188,N_5562,N_5859);
or U6189 (N_6189,N_5566,N_5537);
nand U6190 (N_6190,N_5685,N_5997);
nor U6191 (N_6191,N_5990,N_5786);
xnor U6192 (N_6192,N_5570,N_5745);
and U6193 (N_6193,N_5762,N_5615);
xor U6194 (N_6194,N_5527,N_5834);
and U6195 (N_6195,N_5785,N_5800);
or U6196 (N_6196,N_5836,N_5657);
nand U6197 (N_6197,N_5905,N_5708);
nand U6198 (N_6198,N_5526,N_5902);
and U6199 (N_6199,N_5610,N_5625);
nor U6200 (N_6200,N_5639,N_5529);
or U6201 (N_6201,N_5692,N_5503);
xnor U6202 (N_6202,N_5689,N_5802);
and U6203 (N_6203,N_5531,N_5724);
nand U6204 (N_6204,N_5817,N_5932);
nand U6205 (N_6205,N_5914,N_5839);
nor U6206 (N_6206,N_5772,N_5587);
nor U6207 (N_6207,N_5544,N_5627);
nand U6208 (N_6208,N_5756,N_5781);
and U6209 (N_6209,N_5589,N_5695);
or U6210 (N_6210,N_5744,N_5600);
and U6211 (N_6211,N_5659,N_5770);
nor U6212 (N_6212,N_5825,N_5940);
and U6213 (N_6213,N_5987,N_5766);
nand U6214 (N_6214,N_5939,N_5897);
or U6215 (N_6215,N_5945,N_5518);
nor U6216 (N_6216,N_5551,N_5751);
nor U6217 (N_6217,N_5556,N_5795);
nand U6218 (N_6218,N_5704,N_5761);
or U6219 (N_6219,N_5943,N_5971);
nor U6220 (N_6220,N_5734,N_5797);
and U6221 (N_6221,N_5931,N_5991);
nand U6222 (N_6222,N_5976,N_5993);
or U6223 (N_6223,N_5771,N_5691);
nor U6224 (N_6224,N_5676,N_5694);
nor U6225 (N_6225,N_5560,N_5500);
nor U6226 (N_6226,N_5856,N_5892);
nor U6227 (N_6227,N_5511,N_5820);
nor U6228 (N_6228,N_5666,N_5952);
nand U6229 (N_6229,N_5555,N_5678);
and U6230 (N_6230,N_5984,N_5958);
or U6231 (N_6231,N_5644,N_5955);
nand U6232 (N_6232,N_5655,N_5777);
xnor U6233 (N_6233,N_5585,N_5578);
or U6234 (N_6234,N_5784,N_5829);
nor U6235 (N_6235,N_5539,N_5546);
nand U6236 (N_6236,N_5582,N_5752);
nor U6237 (N_6237,N_5883,N_5563);
nand U6238 (N_6238,N_5842,N_5725);
nand U6239 (N_6239,N_5847,N_5922);
xnor U6240 (N_6240,N_5928,N_5843);
nand U6241 (N_6241,N_5604,N_5796);
nand U6242 (N_6242,N_5693,N_5895);
nand U6243 (N_6243,N_5873,N_5591);
and U6244 (N_6244,N_5890,N_5789);
or U6245 (N_6245,N_5880,N_5521);
nand U6246 (N_6246,N_5904,N_5994);
nand U6247 (N_6247,N_5935,N_5542);
or U6248 (N_6248,N_5832,N_5554);
xnor U6249 (N_6249,N_5567,N_5720);
nand U6250 (N_6250,N_5517,N_5842);
or U6251 (N_6251,N_5902,N_5659);
or U6252 (N_6252,N_5515,N_5657);
nand U6253 (N_6253,N_5888,N_5619);
nor U6254 (N_6254,N_5809,N_5938);
nor U6255 (N_6255,N_5521,N_5723);
or U6256 (N_6256,N_5527,N_5761);
nor U6257 (N_6257,N_5654,N_5716);
nor U6258 (N_6258,N_5708,N_5955);
and U6259 (N_6259,N_5985,N_5741);
and U6260 (N_6260,N_5975,N_5895);
nor U6261 (N_6261,N_5794,N_5702);
xnor U6262 (N_6262,N_5718,N_5635);
nor U6263 (N_6263,N_5943,N_5912);
or U6264 (N_6264,N_5610,N_5878);
nand U6265 (N_6265,N_5995,N_5690);
and U6266 (N_6266,N_5970,N_5990);
xor U6267 (N_6267,N_5999,N_5798);
nor U6268 (N_6268,N_5547,N_5700);
xor U6269 (N_6269,N_5597,N_5840);
nor U6270 (N_6270,N_5924,N_5901);
or U6271 (N_6271,N_5673,N_5856);
xor U6272 (N_6272,N_5950,N_5543);
and U6273 (N_6273,N_5844,N_5548);
nand U6274 (N_6274,N_5596,N_5587);
nor U6275 (N_6275,N_5644,N_5566);
or U6276 (N_6276,N_5514,N_5904);
xnor U6277 (N_6277,N_5685,N_5963);
nand U6278 (N_6278,N_5673,N_5894);
nor U6279 (N_6279,N_5780,N_5613);
xor U6280 (N_6280,N_5844,N_5761);
and U6281 (N_6281,N_5776,N_5990);
nor U6282 (N_6282,N_5712,N_5829);
and U6283 (N_6283,N_5882,N_5892);
nand U6284 (N_6284,N_5587,N_5690);
nor U6285 (N_6285,N_5609,N_5757);
or U6286 (N_6286,N_5824,N_5643);
nor U6287 (N_6287,N_5598,N_5543);
nor U6288 (N_6288,N_5723,N_5778);
and U6289 (N_6289,N_5898,N_5624);
or U6290 (N_6290,N_5739,N_5992);
nor U6291 (N_6291,N_5533,N_5775);
and U6292 (N_6292,N_5941,N_5949);
nand U6293 (N_6293,N_5650,N_5756);
nor U6294 (N_6294,N_5676,N_5506);
nand U6295 (N_6295,N_5816,N_5761);
nand U6296 (N_6296,N_5551,N_5747);
nor U6297 (N_6297,N_5773,N_5910);
or U6298 (N_6298,N_5609,N_5893);
and U6299 (N_6299,N_5889,N_5612);
xor U6300 (N_6300,N_5888,N_5740);
nor U6301 (N_6301,N_5688,N_5873);
and U6302 (N_6302,N_5532,N_5695);
xor U6303 (N_6303,N_5978,N_5690);
or U6304 (N_6304,N_5523,N_5623);
and U6305 (N_6305,N_5601,N_5642);
or U6306 (N_6306,N_5765,N_5593);
or U6307 (N_6307,N_5970,N_5822);
xnor U6308 (N_6308,N_5733,N_5865);
or U6309 (N_6309,N_5947,N_5992);
xor U6310 (N_6310,N_5744,N_5949);
nor U6311 (N_6311,N_5944,N_5861);
nor U6312 (N_6312,N_5527,N_5539);
nand U6313 (N_6313,N_5751,N_5944);
or U6314 (N_6314,N_5837,N_5919);
or U6315 (N_6315,N_5857,N_5701);
and U6316 (N_6316,N_5846,N_5552);
nand U6317 (N_6317,N_5579,N_5688);
nor U6318 (N_6318,N_5696,N_5785);
or U6319 (N_6319,N_5940,N_5856);
nand U6320 (N_6320,N_5500,N_5691);
nor U6321 (N_6321,N_5841,N_5734);
nor U6322 (N_6322,N_5564,N_5819);
and U6323 (N_6323,N_5641,N_5956);
or U6324 (N_6324,N_5949,N_5501);
nand U6325 (N_6325,N_5987,N_5801);
nand U6326 (N_6326,N_5801,N_5812);
xnor U6327 (N_6327,N_5653,N_5768);
and U6328 (N_6328,N_5878,N_5600);
or U6329 (N_6329,N_5516,N_5691);
nand U6330 (N_6330,N_5945,N_5501);
xor U6331 (N_6331,N_5714,N_5511);
nor U6332 (N_6332,N_5790,N_5687);
nand U6333 (N_6333,N_5894,N_5867);
and U6334 (N_6334,N_5689,N_5652);
xor U6335 (N_6335,N_5744,N_5775);
nor U6336 (N_6336,N_5521,N_5829);
and U6337 (N_6337,N_5904,N_5871);
nor U6338 (N_6338,N_5839,N_5595);
or U6339 (N_6339,N_5649,N_5924);
nor U6340 (N_6340,N_5539,N_5842);
and U6341 (N_6341,N_5731,N_5551);
nor U6342 (N_6342,N_5779,N_5508);
nand U6343 (N_6343,N_5780,N_5753);
or U6344 (N_6344,N_5712,N_5651);
nand U6345 (N_6345,N_5968,N_5992);
xor U6346 (N_6346,N_5818,N_5686);
or U6347 (N_6347,N_5982,N_5907);
or U6348 (N_6348,N_5623,N_5512);
xor U6349 (N_6349,N_5505,N_5676);
and U6350 (N_6350,N_5534,N_5670);
and U6351 (N_6351,N_5640,N_5875);
or U6352 (N_6352,N_5960,N_5742);
xor U6353 (N_6353,N_5771,N_5688);
or U6354 (N_6354,N_5749,N_5772);
xnor U6355 (N_6355,N_5976,N_5693);
nor U6356 (N_6356,N_5577,N_5799);
nor U6357 (N_6357,N_5661,N_5710);
nor U6358 (N_6358,N_5747,N_5816);
xnor U6359 (N_6359,N_5938,N_5803);
xor U6360 (N_6360,N_5902,N_5549);
or U6361 (N_6361,N_5861,N_5530);
nand U6362 (N_6362,N_5771,N_5827);
nor U6363 (N_6363,N_5813,N_5517);
or U6364 (N_6364,N_5554,N_5544);
and U6365 (N_6365,N_5550,N_5793);
xnor U6366 (N_6366,N_5845,N_5832);
and U6367 (N_6367,N_5954,N_5724);
and U6368 (N_6368,N_5591,N_5781);
and U6369 (N_6369,N_5635,N_5784);
or U6370 (N_6370,N_5640,N_5877);
nand U6371 (N_6371,N_5543,N_5680);
nor U6372 (N_6372,N_5923,N_5636);
or U6373 (N_6373,N_5602,N_5929);
nand U6374 (N_6374,N_5842,N_5994);
or U6375 (N_6375,N_5784,N_5935);
nor U6376 (N_6376,N_5556,N_5939);
and U6377 (N_6377,N_5736,N_5637);
nand U6378 (N_6378,N_5588,N_5733);
nand U6379 (N_6379,N_5817,N_5828);
and U6380 (N_6380,N_5642,N_5813);
nand U6381 (N_6381,N_5924,N_5959);
and U6382 (N_6382,N_5902,N_5539);
nor U6383 (N_6383,N_5726,N_5681);
nor U6384 (N_6384,N_5584,N_5825);
nor U6385 (N_6385,N_5690,N_5964);
nand U6386 (N_6386,N_5861,N_5735);
and U6387 (N_6387,N_5847,N_5899);
nand U6388 (N_6388,N_5812,N_5875);
and U6389 (N_6389,N_5846,N_5704);
nand U6390 (N_6390,N_5629,N_5593);
and U6391 (N_6391,N_5955,N_5747);
xnor U6392 (N_6392,N_5695,N_5772);
nor U6393 (N_6393,N_5660,N_5589);
or U6394 (N_6394,N_5885,N_5623);
and U6395 (N_6395,N_5509,N_5506);
xor U6396 (N_6396,N_5821,N_5663);
xor U6397 (N_6397,N_5637,N_5593);
and U6398 (N_6398,N_5519,N_5889);
or U6399 (N_6399,N_5697,N_5572);
nand U6400 (N_6400,N_5773,N_5941);
nand U6401 (N_6401,N_5811,N_5638);
nor U6402 (N_6402,N_5699,N_5550);
and U6403 (N_6403,N_5990,N_5561);
nor U6404 (N_6404,N_5749,N_5612);
and U6405 (N_6405,N_5599,N_5957);
or U6406 (N_6406,N_5965,N_5844);
nand U6407 (N_6407,N_5549,N_5986);
or U6408 (N_6408,N_5879,N_5577);
and U6409 (N_6409,N_5742,N_5780);
nor U6410 (N_6410,N_5675,N_5515);
xnor U6411 (N_6411,N_5541,N_5534);
nand U6412 (N_6412,N_5918,N_5856);
and U6413 (N_6413,N_5803,N_5696);
nand U6414 (N_6414,N_5864,N_5973);
nand U6415 (N_6415,N_5997,N_5894);
and U6416 (N_6416,N_5529,N_5695);
nand U6417 (N_6417,N_5551,N_5532);
and U6418 (N_6418,N_5771,N_5730);
nand U6419 (N_6419,N_5963,N_5717);
nand U6420 (N_6420,N_5853,N_5909);
nor U6421 (N_6421,N_5618,N_5601);
xnor U6422 (N_6422,N_5773,N_5520);
xor U6423 (N_6423,N_5712,N_5611);
nand U6424 (N_6424,N_5961,N_5706);
and U6425 (N_6425,N_5759,N_5960);
nand U6426 (N_6426,N_5906,N_5819);
or U6427 (N_6427,N_5657,N_5756);
xor U6428 (N_6428,N_5514,N_5600);
nand U6429 (N_6429,N_5598,N_5980);
xnor U6430 (N_6430,N_5546,N_5988);
nor U6431 (N_6431,N_5935,N_5559);
xnor U6432 (N_6432,N_5854,N_5836);
nand U6433 (N_6433,N_5977,N_5990);
nand U6434 (N_6434,N_5846,N_5578);
nand U6435 (N_6435,N_5526,N_5840);
nor U6436 (N_6436,N_5715,N_5963);
or U6437 (N_6437,N_5605,N_5721);
and U6438 (N_6438,N_5633,N_5923);
and U6439 (N_6439,N_5728,N_5922);
nand U6440 (N_6440,N_5791,N_5812);
nand U6441 (N_6441,N_5816,N_5677);
or U6442 (N_6442,N_5992,N_5662);
nand U6443 (N_6443,N_5773,N_5665);
and U6444 (N_6444,N_5512,N_5561);
nor U6445 (N_6445,N_5674,N_5786);
nand U6446 (N_6446,N_5674,N_5829);
nor U6447 (N_6447,N_5933,N_5890);
or U6448 (N_6448,N_5598,N_5739);
or U6449 (N_6449,N_5648,N_5963);
and U6450 (N_6450,N_5803,N_5975);
xor U6451 (N_6451,N_5598,N_5849);
or U6452 (N_6452,N_5937,N_5773);
and U6453 (N_6453,N_5878,N_5875);
nand U6454 (N_6454,N_5548,N_5654);
nor U6455 (N_6455,N_5943,N_5824);
or U6456 (N_6456,N_5592,N_5716);
and U6457 (N_6457,N_5547,N_5545);
or U6458 (N_6458,N_5938,N_5875);
or U6459 (N_6459,N_5613,N_5647);
nor U6460 (N_6460,N_5650,N_5559);
and U6461 (N_6461,N_5876,N_5555);
xor U6462 (N_6462,N_5893,N_5859);
or U6463 (N_6463,N_5906,N_5588);
xor U6464 (N_6464,N_5890,N_5833);
xnor U6465 (N_6465,N_5564,N_5701);
xor U6466 (N_6466,N_5666,N_5593);
nor U6467 (N_6467,N_5754,N_5781);
nand U6468 (N_6468,N_5685,N_5560);
xnor U6469 (N_6469,N_5535,N_5579);
nand U6470 (N_6470,N_5889,N_5548);
xnor U6471 (N_6471,N_5977,N_5738);
or U6472 (N_6472,N_5728,N_5524);
and U6473 (N_6473,N_5641,N_5769);
xor U6474 (N_6474,N_5738,N_5662);
nor U6475 (N_6475,N_5652,N_5656);
xnor U6476 (N_6476,N_5953,N_5546);
or U6477 (N_6477,N_5575,N_5785);
xnor U6478 (N_6478,N_5860,N_5832);
xnor U6479 (N_6479,N_5913,N_5537);
nand U6480 (N_6480,N_5505,N_5559);
nor U6481 (N_6481,N_5929,N_5650);
nand U6482 (N_6482,N_5615,N_5986);
or U6483 (N_6483,N_5858,N_5582);
or U6484 (N_6484,N_5769,N_5884);
nor U6485 (N_6485,N_5573,N_5782);
nand U6486 (N_6486,N_5564,N_5887);
or U6487 (N_6487,N_5986,N_5934);
and U6488 (N_6488,N_5582,N_5933);
and U6489 (N_6489,N_5932,N_5562);
nor U6490 (N_6490,N_5766,N_5654);
nor U6491 (N_6491,N_5739,N_5991);
or U6492 (N_6492,N_5567,N_5577);
nand U6493 (N_6493,N_5535,N_5501);
nand U6494 (N_6494,N_5894,N_5825);
nor U6495 (N_6495,N_5710,N_5949);
nand U6496 (N_6496,N_5957,N_5708);
or U6497 (N_6497,N_5589,N_5763);
and U6498 (N_6498,N_5786,N_5612);
and U6499 (N_6499,N_5675,N_5559);
nand U6500 (N_6500,N_6087,N_6090);
nand U6501 (N_6501,N_6135,N_6138);
nor U6502 (N_6502,N_6312,N_6273);
nor U6503 (N_6503,N_6427,N_6349);
and U6504 (N_6504,N_6451,N_6156);
nor U6505 (N_6505,N_6259,N_6444);
and U6506 (N_6506,N_6472,N_6228);
and U6507 (N_6507,N_6084,N_6030);
xor U6508 (N_6508,N_6343,N_6042);
and U6509 (N_6509,N_6152,N_6418);
nand U6510 (N_6510,N_6112,N_6245);
and U6511 (N_6511,N_6464,N_6484);
nand U6512 (N_6512,N_6403,N_6426);
nand U6513 (N_6513,N_6244,N_6026);
or U6514 (N_6514,N_6424,N_6260);
nor U6515 (N_6515,N_6121,N_6256);
nand U6516 (N_6516,N_6191,N_6449);
nor U6517 (N_6517,N_6198,N_6368);
nor U6518 (N_6518,N_6194,N_6345);
nor U6519 (N_6519,N_6351,N_6226);
and U6520 (N_6520,N_6432,N_6077);
and U6521 (N_6521,N_6328,N_6159);
and U6522 (N_6522,N_6045,N_6028);
nand U6523 (N_6523,N_6267,N_6285);
nor U6524 (N_6524,N_6443,N_6387);
and U6525 (N_6525,N_6329,N_6347);
or U6526 (N_6526,N_6208,N_6115);
or U6527 (N_6527,N_6106,N_6411);
nand U6528 (N_6528,N_6335,N_6086);
nor U6529 (N_6529,N_6496,N_6127);
and U6530 (N_6530,N_6441,N_6033);
and U6531 (N_6531,N_6295,N_6122);
xor U6532 (N_6532,N_6342,N_6110);
xnor U6533 (N_6533,N_6108,N_6300);
or U6534 (N_6534,N_6423,N_6410);
and U6535 (N_6535,N_6275,N_6271);
or U6536 (N_6536,N_6249,N_6333);
nand U6537 (N_6537,N_6209,N_6177);
nand U6538 (N_6538,N_6397,N_6440);
nor U6539 (N_6539,N_6014,N_6361);
nor U6540 (N_6540,N_6337,N_6216);
and U6541 (N_6541,N_6400,N_6499);
nor U6542 (N_6542,N_6034,N_6105);
or U6543 (N_6543,N_6079,N_6057);
or U6544 (N_6544,N_6120,N_6479);
or U6545 (N_6545,N_6100,N_6221);
nand U6546 (N_6546,N_6303,N_6085);
and U6547 (N_6547,N_6016,N_6011);
nor U6548 (N_6548,N_6032,N_6224);
or U6549 (N_6549,N_6294,N_6075);
or U6550 (N_6550,N_6438,N_6185);
nor U6551 (N_6551,N_6453,N_6407);
nor U6552 (N_6552,N_6282,N_6281);
nand U6553 (N_6553,N_6182,N_6466);
nand U6554 (N_6554,N_6165,N_6018);
or U6555 (N_6555,N_6459,N_6416);
nand U6556 (N_6556,N_6072,N_6098);
nor U6557 (N_6557,N_6048,N_6131);
or U6558 (N_6558,N_6354,N_6067);
nor U6559 (N_6559,N_6492,N_6398);
or U6560 (N_6560,N_6157,N_6266);
and U6561 (N_6561,N_6477,N_6377);
or U6562 (N_6562,N_6279,N_6174);
and U6563 (N_6563,N_6237,N_6413);
and U6564 (N_6564,N_6362,N_6483);
nor U6565 (N_6565,N_6463,N_6024);
and U6566 (N_6566,N_6020,N_6471);
xnor U6567 (N_6567,N_6289,N_6164);
or U6568 (N_6568,N_6036,N_6031);
nor U6569 (N_6569,N_6378,N_6417);
and U6570 (N_6570,N_6145,N_6091);
nor U6571 (N_6571,N_6405,N_6428);
or U6572 (N_6572,N_6231,N_6118);
and U6573 (N_6573,N_6317,N_6313);
nor U6574 (N_6574,N_6461,N_6311);
or U6575 (N_6575,N_6205,N_6066);
nor U6576 (N_6576,N_6211,N_6324);
nand U6577 (N_6577,N_6462,N_6161);
xnor U6578 (N_6578,N_6059,N_6227);
or U6579 (N_6579,N_6327,N_6478);
or U6580 (N_6580,N_6450,N_6035);
nand U6581 (N_6581,N_6151,N_6366);
nand U6582 (N_6582,N_6125,N_6095);
and U6583 (N_6583,N_6040,N_6242);
xnor U6584 (N_6584,N_6265,N_6027);
nor U6585 (N_6585,N_6334,N_6186);
xnor U6586 (N_6586,N_6207,N_6263);
and U6587 (N_6587,N_6485,N_6482);
or U6588 (N_6588,N_6234,N_6204);
and U6589 (N_6589,N_6447,N_6247);
nor U6590 (N_6590,N_6232,N_6310);
and U6591 (N_6591,N_6128,N_6065);
or U6592 (N_6592,N_6049,N_6308);
nor U6593 (N_6593,N_6376,N_6465);
or U6594 (N_6594,N_6195,N_6150);
nor U6595 (N_6595,N_6214,N_6364);
nand U6596 (N_6596,N_6332,N_6350);
nand U6597 (N_6597,N_6352,N_6458);
and U6598 (N_6598,N_6415,N_6010);
and U6599 (N_6599,N_6373,N_6215);
or U6600 (N_6600,N_6060,N_6488);
or U6601 (N_6601,N_6047,N_6253);
or U6602 (N_6602,N_6183,N_6004);
and U6603 (N_6603,N_6448,N_6494);
nand U6604 (N_6604,N_6046,N_6068);
nand U6605 (N_6605,N_6480,N_6358);
nand U6606 (N_6606,N_6469,N_6139);
and U6607 (N_6607,N_6379,N_6076);
or U6608 (N_6608,N_6476,N_6369);
nor U6609 (N_6609,N_6434,N_6320);
and U6610 (N_6610,N_6339,N_6061);
nor U6611 (N_6611,N_6173,N_6326);
nor U6612 (N_6612,N_6201,N_6495);
and U6613 (N_6613,N_6390,N_6467);
and U6614 (N_6614,N_6154,N_6168);
nand U6615 (N_6615,N_6013,N_6055);
and U6616 (N_6616,N_6305,N_6435);
nor U6617 (N_6617,N_6223,N_6250);
nor U6618 (N_6618,N_6491,N_6180);
or U6619 (N_6619,N_6497,N_6370);
xor U6620 (N_6620,N_6070,N_6129);
and U6621 (N_6621,N_6371,N_6425);
and U6622 (N_6622,N_6096,N_6431);
or U6623 (N_6623,N_6330,N_6318);
and U6624 (N_6624,N_6325,N_6296);
or U6625 (N_6625,N_6130,N_6074);
nor U6626 (N_6626,N_6172,N_6419);
nor U6627 (N_6627,N_6290,N_6019);
nor U6628 (N_6628,N_6468,N_6422);
nand U6629 (N_6629,N_6230,N_6007);
and U6630 (N_6630,N_6261,N_6162);
nor U6631 (N_6631,N_6147,N_6489);
nor U6632 (N_6632,N_6141,N_6103);
or U6633 (N_6633,N_6252,N_6420);
nor U6634 (N_6634,N_6301,N_6088);
and U6635 (N_6635,N_6190,N_6299);
and U6636 (N_6636,N_6365,N_6283);
nor U6637 (N_6637,N_6023,N_6430);
nor U6638 (N_6638,N_6386,N_6192);
nand U6639 (N_6639,N_6175,N_6439);
nor U6640 (N_6640,N_6291,N_6081);
nand U6641 (N_6641,N_6189,N_6113);
nor U6642 (N_6642,N_6184,N_6187);
or U6643 (N_6643,N_6382,N_6298);
and U6644 (N_6644,N_6243,N_6063);
nor U6645 (N_6645,N_6475,N_6302);
nand U6646 (N_6646,N_6064,N_6481);
or U6647 (N_6647,N_6384,N_6414);
nand U6648 (N_6648,N_6277,N_6452);
nor U6649 (N_6649,N_6314,N_6153);
nand U6650 (N_6650,N_6341,N_6225);
and U6651 (N_6651,N_6235,N_6136);
xnor U6652 (N_6652,N_6241,N_6394);
and U6653 (N_6653,N_6071,N_6197);
or U6654 (N_6654,N_6169,N_6356);
or U6655 (N_6655,N_6078,N_6179);
nand U6656 (N_6656,N_6321,N_6372);
and U6657 (N_6657,N_6490,N_6089);
xor U6658 (N_6658,N_6137,N_6114);
xnor U6659 (N_6659,N_6437,N_6346);
and U6660 (N_6660,N_6486,N_6493);
nand U6661 (N_6661,N_6170,N_6022);
and U6662 (N_6662,N_6017,N_6163);
and U6663 (N_6663,N_6158,N_6116);
nand U6664 (N_6664,N_6240,N_6012);
and U6665 (N_6665,N_6248,N_6206);
nand U6666 (N_6666,N_6276,N_6003);
or U6667 (N_6667,N_6412,N_6393);
or U6668 (N_6668,N_6119,N_6353);
or U6669 (N_6669,N_6094,N_6280);
nand U6670 (N_6670,N_6188,N_6196);
nand U6671 (N_6671,N_6293,N_6268);
nor U6672 (N_6672,N_6322,N_6093);
nand U6673 (N_6673,N_6203,N_6257);
or U6674 (N_6674,N_6446,N_6166);
and U6675 (N_6675,N_6238,N_6274);
nor U6676 (N_6676,N_6001,N_6392);
or U6677 (N_6677,N_6178,N_6388);
nor U6678 (N_6678,N_6021,N_6292);
nor U6679 (N_6679,N_6236,N_6142);
nand U6680 (N_6680,N_6404,N_6455);
and U6681 (N_6681,N_6336,N_6391);
nand U6682 (N_6682,N_6133,N_6286);
xnor U6683 (N_6683,N_6155,N_6383);
nor U6684 (N_6684,N_6340,N_6357);
nand U6685 (N_6685,N_6050,N_6304);
and U6686 (N_6686,N_6210,N_6367);
or U6687 (N_6687,N_6399,N_6044);
or U6688 (N_6688,N_6134,N_6073);
nor U6689 (N_6689,N_6009,N_6456);
nor U6690 (N_6690,N_6396,N_6262);
or U6691 (N_6691,N_6360,N_6316);
or U6692 (N_6692,N_6385,N_6278);
nor U6693 (N_6693,N_6000,N_6309);
nor U6694 (N_6694,N_6251,N_6212);
and U6695 (N_6695,N_6052,N_6144);
nor U6696 (N_6696,N_6421,N_6083);
nor U6697 (N_6697,N_6233,N_6069);
and U6698 (N_6698,N_6111,N_6143);
nor U6699 (N_6699,N_6053,N_6005);
nor U6700 (N_6700,N_6474,N_6389);
nor U6701 (N_6701,N_6470,N_6307);
nor U6702 (N_6702,N_6123,N_6355);
nand U6703 (N_6703,N_6109,N_6270);
or U6704 (N_6704,N_6460,N_6315);
nor U6705 (N_6705,N_6222,N_6015);
nand U6706 (N_6706,N_6038,N_6176);
xor U6707 (N_6707,N_6097,N_6445);
nor U6708 (N_6708,N_6008,N_6104);
nand U6709 (N_6709,N_6338,N_6043);
and U6710 (N_6710,N_6487,N_6433);
and U6711 (N_6711,N_6126,N_6062);
xnor U6712 (N_6712,N_6148,N_6099);
nor U6713 (N_6713,N_6348,N_6284);
and U6714 (N_6714,N_6442,N_6374);
nand U6715 (N_6715,N_6058,N_6375);
or U6716 (N_6716,N_6082,N_6102);
nand U6717 (N_6717,N_6101,N_6297);
or U6718 (N_6718,N_6331,N_6002);
and U6719 (N_6719,N_6402,N_6473);
and U6720 (N_6720,N_6429,N_6344);
nand U6721 (N_6721,N_6037,N_6039);
nor U6722 (N_6722,N_6269,N_6199);
nor U6723 (N_6723,N_6160,N_6006);
nand U6724 (N_6724,N_6246,N_6051);
and U6725 (N_6725,N_6239,N_6395);
and U6726 (N_6726,N_6149,N_6167);
or U6727 (N_6727,N_6381,N_6219);
and U6728 (N_6728,N_6408,N_6146);
nand U6729 (N_6729,N_6254,N_6132);
nor U6730 (N_6730,N_6080,N_6171);
xnor U6731 (N_6731,N_6056,N_6200);
nand U6732 (N_6732,N_6218,N_6054);
nor U6733 (N_6733,N_6140,N_6306);
or U6734 (N_6734,N_6220,N_6229);
and U6735 (N_6735,N_6272,N_6107);
or U6736 (N_6736,N_6287,N_6202);
nand U6737 (N_6737,N_6401,N_6193);
or U6738 (N_6738,N_6323,N_6436);
nor U6739 (N_6739,N_6457,N_6498);
nand U6740 (N_6740,N_6217,N_6406);
and U6741 (N_6741,N_6029,N_6255);
or U6742 (N_6742,N_6213,N_6025);
or U6743 (N_6743,N_6319,N_6454);
or U6744 (N_6744,N_6409,N_6258);
xnor U6745 (N_6745,N_6124,N_6264);
or U6746 (N_6746,N_6359,N_6181);
or U6747 (N_6747,N_6363,N_6288);
or U6748 (N_6748,N_6117,N_6092);
nand U6749 (N_6749,N_6380,N_6041);
and U6750 (N_6750,N_6102,N_6294);
or U6751 (N_6751,N_6342,N_6031);
nand U6752 (N_6752,N_6250,N_6305);
nand U6753 (N_6753,N_6071,N_6140);
and U6754 (N_6754,N_6006,N_6278);
and U6755 (N_6755,N_6263,N_6479);
or U6756 (N_6756,N_6419,N_6427);
nand U6757 (N_6757,N_6399,N_6458);
and U6758 (N_6758,N_6054,N_6222);
nor U6759 (N_6759,N_6300,N_6464);
nor U6760 (N_6760,N_6417,N_6200);
nand U6761 (N_6761,N_6043,N_6319);
xnor U6762 (N_6762,N_6066,N_6053);
nand U6763 (N_6763,N_6167,N_6195);
and U6764 (N_6764,N_6289,N_6131);
and U6765 (N_6765,N_6410,N_6401);
or U6766 (N_6766,N_6090,N_6239);
xnor U6767 (N_6767,N_6020,N_6056);
and U6768 (N_6768,N_6299,N_6077);
and U6769 (N_6769,N_6182,N_6252);
and U6770 (N_6770,N_6415,N_6208);
and U6771 (N_6771,N_6132,N_6314);
or U6772 (N_6772,N_6378,N_6136);
nor U6773 (N_6773,N_6138,N_6296);
or U6774 (N_6774,N_6395,N_6197);
nand U6775 (N_6775,N_6454,N_6337);
and U6776 (N_6776,N_6257,N_6188);
or U6777 (N_6777,N_6405,N_6145);
nor U6778 (N_6778,N_6163,N_6218);
nor U6779 (N_6779,N_6425,N_6195);
or U6780 (N_6780,N_6372,N_6170);
nand U6781 (N_6781,N_6388,N_6275);
nand U6782 (N_6782,N_6293,N_6247);
xor U6783 (N_6783,N_6378,N_6493);
or U6784 (N_6784,N_6485,N_6428);
nand U6785 (N_6785,N_6056,N_6296);
nor U6786 (N_6786,N_6410,N_6326);
or U6787 (N_6787,N_6483,N_6077);
nor U6788 (N_6788,N_6275,N_6097);
or U6789 (N_6789,N_6368,N_6404);
nor U6790 (N_6790,N_6111,N_6318);
nand U6791 (N_6791,N_6247,N_6367);
or U6792 (N_6792,N_6161,N_6204);
nor U6793 (N_6793,N_6398,N_6200);
nand U6794 (N_6794,N_6426,N_6111);
and U6795 (N_6795,N_6050,N_6204);
nand U6796 (N_6796,N_6023,N_6148);
nor U6797 (N_6797,N_6337,N_6174);
nor U6798 (N_6798,N_6366,N_6303);
nand U6799 (N_6799,N_6277,N_6145);
and U6800 (N_6800,N_6140,N_6176);
nand U6801 (N_6801,N_6240,N_6414);
nor U6802 (N_6802,N_6185,N_6133);
or U6803 (N_6803,N_6035,N_6080);
nand U6804 (N_6804,N_6097,N_6180);
and U6805 (N_6805,N_6296,N_6239);
nor U6806 (N_6806,N_6021,N_6087);
xor U6807 (N_6807,N_6284,N_6398);
or U6808 (N_6808,N_6361,N_6081);
nor U6809 (N_6809,N_6137,N_6194);
nand U6810 (N_6810,N_6307,N_6474);
nand U6811 (N_6811,N_6021,N_6390);
nand U6812 (N_6812,N_6135,N_6198);
or U6813 (N_6813,N_6468,N_6113);
nand U6814 (N_6814,N_6021,N_6409);
nand U6815 (N_6815,N_6265,N_6195);
and U6816 (N_6816,N_6151,N_6434);
nand U6817 (N_6817,N_6419,N_6047);
nand U6818 (N_6818,N_6177,N_6418);
and U6819 (N_6819,N_6191,N_6053);
nor U6820 (N_6820,N_6102,N_6190);
xnor U6821 (N_6821,N_6020,N_6301);
xnor U6822 (N_6822,N_6214,N_6394);
nor U6823 (N_6823,N_6058,N_6345);
or U6824 (N_6824,N_6082,N_6455);
nand U6825 (N_6825,N_6150,N_6443);
or U6826 (N_6826,N_6398,N_6394);
or U6827 (N_6827,N_6206,N_6418);
nand U6828 (N_6828,N_6491,N_6160);
or U6829 (N_6829,N_6073,N_6111);
nand U6830 (N_6830,N_6449,N_6335);
nand U6831 (N_6831,N_6465,N_6256);
nor U6832 (N_6832,N_6016,N_6131);
and U6833 (N_6833,N_6330,N_6231);
nor U6834 (N_6834,N_6415,N_6385);
and U6835 (N_6835,N_6323,N_6097);
xor U6836 (N_6836,N_6097,N_6492);
or U6837 (N_6837,N_6454,N_6023);
nand U6838 (N_6838,N_6161,N_6108);
nand U6839 (N_6839,N_6317,N_6396);
or U6840 (N_6840,N_6386,N_6180);
and U6841 (N_6841,N_6372,N_6129);
or U6842 (N_6842,N_6368,N_6362);
and U6843 (N_6843,N_6083,N_6369);
or U6844 (N_6844,N_6262,N_6395);
nor U6845 (N_6845,N_6081,N_6383);
nor U6846 (N_6846,N_6224,N_6043);
and U6847 (N_6847,N_6302,N_6084);
nand U6848 (N_6848,N_6406,N_6389);
or U6849 (N_6849,N_6243,N_6357);
or U6850 (N_6850,N_6357,N_6224);
and U6851 (N_6851,N_6361,N_6326);
and U6852 (N_6852,N_6023,N_6245);
nand U6853 (N_6853,N_6295,N_6285);
nand U6854 (N_6854,N_6369,N_6275);
and U6855 (N_6855,N_6308,N_6001);
xor U6856 (N_6856,N_6328,N_6103);
or U6857 (N_6857,N_6255,N_6411);
or U6858 (N_6858,N_6184,N_6219);
nor U6859 (N_6859,N_6115,N_6085);
or U6860 (N_6860,N_6106,N_6100);
and U6861 (N_6861,N_6461,N_6268);
nand U6862 (N_6862,N_6034,N_6139);
nor U6863 (N_6863,N_6117,N_6486);
or U6864 (N_6864,N_6420,N_6164);
or U6865 (N_6865,N_6341,N_6409);
nor U6866 (N_6866,N_6442,N_6134);
nor U6867 (N_6867,N_6298,N_6164);
nand U6868 (N_6868,N_6130,N_6100);
and U6869 (N_6869,N_6286,N_6095);
and U6870 (N_6870,N_6227,N_6461);
xnor U6871 (N_6871,N_6232,N_6189);
xnor U6872 (N_6872,N_6092,N_6423);
and U6873 (N_6873,N_6152,N_6334);
and U6874 (N_6874,N_6181,N_6012);
xor U6875 (N_6875,N_6254,N_6476);
and U6876 (N_6876,N_6087,N_6245);
nor U6877 (N_6877,N_6190,N_6372);
and U6878 (N_6878,N_6377,N_6146);
or U6879 (N_6879,N_6291,N_6012);
nor U6880 (N_6880,N_6264,N_6069);
xor U6881 (N_6881,N_6286,N_6160);
nor U6882 (N_6882,N_6223,N_6316);
nand U6883 (N_6883,N_6202,N_6164);
and U6884 (N_6884,N_6433,N_6148);
nand U6885 (N_6885,N_6409,N_6370);
xor U6886 (N_6886,N_6445,N_6273);
nand U6887 (N_6887,N_6343,N_6319);
and U6888 (N_6888,N_6372,N_6187);
and U6889 (N_6889,N_6387,N_6310);
or U6890 (N_6890,N_6109,N_6063);
nor U6891 (N_6891,N_6424,N_6038);
and U6892 (N_6892,N_6371,N_6121);
and U6893 (N_6893,N_6192,N_6080);
and U6894 (N_6894,N_6236,N_6004);
nor U6895 (N_6895,N_6278,N_6362);
or U6896 (N_6896,N_6355,N_6474);
and U6897 (N_6897,N_6372,N_6310);
xnor U6898 (N_6898,N_6036,N_6062);
xor U6899 (N_6899,N_6444,N_6215);
nand U6900 (N_6900,N_6179,N_6177);
and U6901 (N_6901,N_6491,N_6298);
and U6902 (N_6902,N_6072,N_6104);
or U6903 (N_6903,N_6491,N_6280);
and U6904 (N_6904,N_6056,N_6216);
and U6905 (N_6905,N_6028,N_6292);
or U6906 (N_6906,N_6134,N_6182);
nor U6907 (N_6907,N_6187,N_6377);
nor U6908 (N_6908,N_6437,N_6391);
nor U6909 (N_6909,N_6343,N_6278);
and U6910 (N_6910,N_6145,N_6391);
or U6911 (N_6911,N_6131,N_6069);
and U6912 (N_6912,N_6351,N_6234);
nand U6913 (N_6913,N_6410,N_6350);
nand U6914 (N_6914,N_6249,N_6394);
or U6915 (N_6915,N_6020,N_6436);
and U6916 (N_6916,N_6288,N_6255);
or U6917 (N_6917,N_6375,N_6362);
nand U6918 (N_6918,N_6025,N_6138);
nor U6919 (N_6919,N_6440,N_6066);
and U6920 (N_6920,N_6010,N_6089);
nand U6921 (N_6921,N_6221,N_6261);
or U6922 (N_6922,N_6054,N_6156);
nand U6923 (N_6923,N_6425,N_6064);
and U6924 (N_6924,N_6277,N_6475);
nor U6925 (N_6925,N_6351,N_6252);
and U6926 (N_6926,N_6211,N_6421);
or U6927 (N_6927,N_6293,N_6313);
and U6928 (N_6928,N_6181,N_6062);
and U6929 (N_6929,N_6109,N_6036);
nand U6930 (N_6930,N_6078,N_6269);
nand U6931 (N_6931,N_6449,N_6454);
nand U6932 (N_6932,N_6086,N_6156);
or U6933 (N_6933,N_6377,N_6314);
nand U6934 (N_6934,N_6191,N_6181);
nand U6935 (N_6935,N_6288,N_6239);
and U6936 (N_6936,N_6380,N_6420);
and U6937 (N_6937,N_6409,N_6162);
nor U6938 (N_6938,N_6201,N_6414);
nand U6939 (N_6939,N_6249,N_6425);
nand U6940 (N_6940,N_6421,N_6189);
nor U6941 (N_6941,N_6166,N_6383);
nand U6942 (N_6942,N_6078,N_6173);
nor U6943 (N_6943,N_6309,N_6345);
nor U6944 (N_6944,N_6245,N_6473);
or U6945 (N_6945,N_6394,N_6361);
nor U6946 (N_6946,N_6051,N_6095);
nor U6947 (N_6947,N_6090,N_6102);
xnor U6948 (N_6948,N_6014,N_6028);
nor U6949 (N_6949,N_6022,N_6029);
nor U6950 (N_6950,N_6143,N_6467);
or U6951 (N_6951,N_6008,N_6466);
nand U6952 (N_6952,N_6416,N_6031);
nor U6953 (N_6953,N_6486,N_6133);
or U6954 (N_6954,N_6288,N_6180);
and U6955 (N_6955,N_6106,N_6317);
and U6956 (N_6956,N_6427,N_6361);
nand U6957 (N_6957,N_6115,N_6224);
and U6958 (N_6958,N_6240,N_6379);
and U6959 (N_6959,N_6352,N_6077);
nand U6960 (N_6960,N_6108,N_6094);
or U6961 (N_6961,N_6238,N_6130);
nand U6962 (N_6962,N_6057,N_6226);
and U6963 (N_6963,N_6305,N_6312);
nor U6964 (N_6964,N_6384,N_6354);
nand U6965 (N_6965,N_6085,N_6495);
nor U6966 (N_6966,N_6038,N_6136);
nand U6967 (N_6967,N_6200,N_6469);
nand U6968 (N_6968,N_6054,N_6347);
nor U6969 (N_6969,N_6321,N_6026);
xnor U6970 (N_6970,N_6433,N_6010);
or U6971 (N_6971,N_6307,N_6294);
xnor U6972 (N_6972,N_6219,N_6450);
xnor U6973 (N_6973,N_6244,N_6059);
and U6974 (N_6974,N_6330,N_6058);
and U6975 (N_6975,N_6353,N_6448);
nand U6976 (N_6976,N_6326,N_6177);
or U6977 (N_6977,N_6170,N_6478);
nand U6978 (N_6978,N_6128,N_6244);
and U6979 (N_6979,N_6133,N_6449);
nor U6980 (N_6980,N_6477,N_6284);
nand U6981 (N_6981,N_6312,N_6143);
nor U6982 (N_6982,N_6291,N_6403);
nand U6983 (N_6983,N_6251,N_6455);
or U6984 (N_6984,N_6247,N_6084);
and U6985 (N_6985,N_6443,N_6036);
xor U6986 (N_6986,N_6480,N_6450);
xnor U6987 (N_6987,N_6447,N_6361);
nor U6988 (N_6988,N_6213,N_6261);
and U6989 (N_6989,N_6008,N_6431);
nor U6990 (N_6990,N_6153,N_6315);
xnor U6991 (N_6991,N_6210,N_6078);
nor U6992 (N_6992,N_6021,N_6007);
xnor U6993 (N_6993,N_6142,N_6404);
and U6994 (N_6994,N_6443,N_6496);
nand U6995 (N_6995,N_6090,N_6391);
nor U6996 (N_6996,N_6312,N_6005);
nor U6997 (N_6997,N_6342,N_6442);
nor U6998 (N_6998,N_6167,N_6179);
xnor U6999 (N_6999,N_6139,N_6093);
nand U7000 (N_7000,N_6606,N_6886);
nor U7001 (N_7001,N_6749,N_6548);
and U7002 (N_7002,N_6636,N_6754);
or U7003 (N_7003,N_6511,N_6753);
and U7004 (N_7004,N_6744,N_6848);
or U7005 (N_7005,N_6619,N_6656);
nor U7006 (N_7006,N_6766,N_6569);
and U7007 (N_7007,N_6964,N_6947);
or U7008 (N_7008,N_6705,N_6893);
nand U7009 (N_7009,N_6602,N_6661);
nand U7010 (N_7010,N_6919,N_6629);
or U7011 (N_7011,N_6706,N_6934);
nand U7012 (N_7012,N_6707,N_6741);
xnor U7013 (N_7013,N_6570,N_6853);
nor U7014 (N_7014,N_6679,N_6609);
nand U7015 (N_7015,N_6946,N_6502);
nor U7016 (N_7016,N_6750,N_6697);
xnor U7017 (N_7017,N_6740,N_6614);
nor U7018 (N_7018,N_6748,N_6880);
nand U7019 (N_7019,N_6824,N_6850);
or U7020 (N_7020,N_6993,N_6516);
nor U7021 (N_7021,N_6896,N_6581);
and U7022 (N_7022,N_6857,N_6696);
and U7023 (N_7023,N_6774,N_6873);
and U7024 (N_7024,N_6508,N_6959);
or U7025 (N_7025,N_6898,N_6835);
or U7026 (N_7026,N_6802,N_6621);
nor U7027 (N_7027,N_6586,N_6555);
nand U7028 (N_7028,N_6522,N_6683);
nor U7029 (N_7029,N_6885,N_6541);
xnor U7030 (N_7030,N_6889,N_6550);
and U7031 (N_7031,N_6940,N_6876);
nand U7032 (N_7032,N_6540,N_6616);
or U7033 (N_7033,N_6657,N_6643);
nand U7034 (N_7034,N_6858,N_6836);
and U7035 (N_7035,N_6899,N_6622);
xor U7036 (N_7036,N_6952,N_6674);
and U7037 (N_7037,N_6930,N_6973);
nor U7038 (N_7038,N_6726,N_6637);
xor U7039 (N_7039,N_6936,N_6743);
or U7040 (N_7040,N_6554,N_6784);
or U7041 (N_7041,N_6829,N_6735);
nor U7042 (N_7042,N_6755,N_6975);
and U7043 (N_7043,N_6813,N_6684);
xnor U7044 (N_7044,N_6982,N_6931);
nand U7045 (N_7045,N_6807,N_6709);
and U7046 (N_7046,N_6939,N_6579);
nor U7047 (N_7047,N_6590,N_6632);
nor U7048 (N_7048,N_6781,N_6715);
nand U7049 (N_7049,N_6641,N_6830);
nand U7050 (N_7050,N_6504,N_6675);
or U7051 (N_7051,N_6926,N_6794);
nor U7052 (N_7052,N_6659,N_6509);
and U7053 (N_7053,N_6694,N_6681);
nor U7054 (N_7054,N_6861,N_6686);
nor U7055 (N_7055,N_6669,N_6551);
nor U7056 (N_7056,N_6994,N_6860);
and U7057 (N_7057,N_6957,N_6595);
and U7058 (N_7058,N_6881,N_6981);
and U7059 (N_7059,N_6950,N_6534);
xor U7060 (N_7060,N_6729,N_6601);
and U7061 (N_7061,N_6834,N_6600);
or U7062 (N_7062,N_6867,N_6650);
nor U7063 (N_7063,N_6677,N_6800);
or U7064 (N_7064,N_6965,N_6539);
nand U7065 (N_7065,N_6587,N_6529);
nor U7066 (N_7066,N_6877,N_6756);
nor U7067 (N_7067,N_6764,N_6521);
or U7068 (N_7068,N_6627,N_6501);
nor U7069 (N_7069,N_6838,N_6678);
and U7070 (N_7070,N_6514,N_6699);
and U7071 (N_7071,N_6820,N_6623);
and U7072 (N_7072,N_6597,N_6953);
or U7073 (N_7073,N_6640,N_6798);
nor U7074 (N_7074,N_6634,N_6689);
nand U7075 (N_7075,N_6728,N_6865);
nand U7076 (N_7076,N_6943,N_6868);
nand U7077 (N_7077,N_6759,N_6917);
nor U7078 (N_7078,N_6546,N_6701);
nand U7079 (N_7079,N_6664,N_6773);
or U7080 (N_7080,N_6969,N_6900);
or U7081 (N_7081,N_6929,N_6779);
xnor U7082 (N_7082,N_6823,N_6770);
or U7083 (N_7083,N_6882,N_6788);
nor U7084 (N_7084,N_6870,N_6879);
or U7085 (N_7085,N_6908,N_6512);
and U7086 (N_7086,N_6513,N_6812);
nor U7087 (N_7087,N_6518,N_6523);
nor U7088 (N_7088,N_6817,N_6665);
and U7089 (N_7089,N_6777,N_6765);
or U7090 (N_7090,N_6574,N_6789);
xor U7091 (N_7091,N_6702,N_6792);
and U7092 (N_7092,N_6951,N_6670);
nand U7093 (N_7093,N_6575,N_6978);
nor U7094 (N_7094,N_6577,N_6713);
xnor U7095 (N_7095,N_6795,N_6814);
nand U7096 (N_7096,N_6971,N_6724);
nor U7097 (N_7097,N_6653,N_6685);
nand U7098 (N_7098,N_6588,N_6598);
nor U7099 (N_7099,N_6954,N_6872);
nor U7100 (N_7100,N_6688,N_6822);
nor U7101 (N_7101,N_6758,N_6974);
and U7102 (N_7102,N_6630,N_6763);
and U7103 (N_7103,N_6801,N_6921);
and U7104 (N_7104,N_6966,N_6985);
nand U7105 (N_7105,N_6720,N_6768);
or U7106 (N_7106,N_6840,N_6628);
nor U7107 (N_7107,N_6576,N_6785);
nand U7108 (N_7108,N_6552,N_6827);
and U7109 (N_7109,N_6625,N_6998);
or U7110 (N_7110,N_6646,N_6658);
or U7111 (N_7111,N_6914,N_6560);
and U7112 (N_7112,N_6949,N_6986);
and U7113 (N_7113,N_6567,N_6673);
nor U7114 (N_7114,N_6797,N_6533);
nand U7115 (N_7115,N_6517,N_6837);
nor U7116 (N_7116,N_6922,N_6693);
nor U7117 (N_7117,N_6531,N_6895);
or U7118 (N_7118,N_6948,N_6935);
nor U7119 (N_7119,N_6642,N_6912);
nor U7120 (N_7120,N_6866,N_6730);
nand U7121 (N_7121,N_6941,N_6903);
nand U7122 (N_7122,N_6825,N_6704);
nand U7123 (N_7123,N_6992,N_6762);
nor U7124 (N_7124,N_6584,N_6938);
and U7125 (N_7125,N_6894,N_6663);
and U7126 (N_7126,N_6796,N_6736);
and U7127 (N_7127,N_6902,N_6901);
nand U7128 (N_7128,N_6828,N_6725);
and U7129 (N_7129,N_6542,N_6582);
and U7130 (N_7130,N_6972,N_6937);
or U7131 (N_7131,N_6718,N_6568);
nor U7132 (N_7132,N_6624,N_6589);
nand U7133 (N_7133,N_6869,N_6769);
or U7134 (N_7134,N_6671,N_6710);
or U7135 (N_7135,N_6703,N_6803);
nor U7136 (N_7136,N_6549,N_6532);
nand U7137 (N_7137,N_6591,N_6594);
or U7138 (N_7138,N_6578,N_6841);
nor U7139 (N_7139,N_6553,N_6995);
xnor U7140 (N_7140,N_6644,N_6832);
and U7141 (N_7141,N_6721,N_6698);
and U7142 (N_7142,N_6535,N_6660);
nand U7143 (N_7143,N_6847,N_6500);
or U7144 (N_7144,N_6599,N_6536);
nand U7145 (N_7145,N_6846,N_6558);
nand U7146 (N_7146,N_6617,N_6910);
nor U7147 (N_7147,N_6719,N_6733);
or U7148 (N_7148,N_6888,N_6810);
nor U7149 (N_7149,N_6708,N_6615);
or U7150 (N_7150,N_6571,N_6566);
or U7151 (N_7151,N_6647,N_6676);
nand U7152 (N_7152,N_6690,N_6804);
xnor U7153 (N_7153,N_6849,N_6855);
and U7154 (N_7154,N_6808,N_6700);
and U7155 (N_7155,N_6916,N_6924);
nor U7156 (N_7156,N_6731,N_6976);
or U7157 (N_7157,N_6906,N_6528);
or U7158 (N_7158,N_6933,N_6815);
nor U7159 (N_7159,N_6852,N_6944);
and U7160 (N_7160,N_6526,N_6716);
nand U7161 (N_7161,N_6883,N_6775);
or U7162 (N_7162,N_6778,N_6672);
or U7163 (N_7163,N_6923,N_6510);
and U7164 (N_7164,N_6562,N_6955);
or U7165 (N_7165,N_6932,N_6737);
or U7166 (N_7166,N_6648,N_6863);
nor U7167 (N_7167,N_6787,N_6727);
xnor U7168 (N_7168,N_6816,N_6907);
and U7169 (N_7169,N_6842,N_6874);
nand U7170 (N_7170,N_6927,N_6610);
or U7171 (N_7171,N_6572,N_6742);
nor U7172 (N_7172,N_6620,N_6618);
nor U7173 (N_7173,N_6603,N_6891);
or U7174 (N_7174,N_6682,N_6958);
nand U7175 (N_7175,N_6585,N_6605);
nor U7176 (N_7176,N_6593,N_6864);
or U7177 (N_7177,N_6772,N_6738);
nor U7178 (N_7178,N_6984,N_6928);
and U7179 (N_7179,N_6913,N_6780);
and U7180 (N_7180,N_6524,N_6996);
or U7181 (N_7181,N_6732,N_6988);
nand U7182 (N_7182,N_6854,N_6680);
or U7183 (N_7183,N_6503,N_6687);
nand U7184 (N_7184,N_6544,N_6547);
nor U7185 (N_7185,N_6989,N_6545);
or U7186 (N_7186,N_6862,N_6638);
nor U7187 (N_7187,N_6890,N_6525);
or U7188 (N_7188,N_6875,N_6915);
nor U7189 (N_7189,N_6734,N_6563);
or U7190 (N_7190,N_6592,N_6811);
and U7191 (N_7191,N_6979,N_6859);
and U7192 (N_7192,N_6608,N_6945);
nand U7193 (N_7193,N_6564,N_6892);
nor U7194 (N_7194,N_6918,N_6538);
xor U7195 (N_7195,N_6712,N_6826);
or U7196 (N_7196,N_6666,N_6667);
and U7197 (N_7197,N_6845,N_6782);
or U7198 (N_7198,N_6505,N_6987);
nor U7199 (N_7199,N_6723,N_6767);
nand U7200 (N_7200,N_6839,N_6583);
nand U7201 (N_7201,N_6999,N_6960);
and U7202 (N_7202,N_6956,N_6980);
and U7203 (N_7203,N_6559,N_6695);
and U7204 (N_7204,N_6543,N_6771);
or U7205 (N_7205,N_6920,N_6821);
nand U7206 (N_7206,N_6851,N_6612);
nand U7207 (N_7207,N_6613,N_6604);
xor U7208 (N_7208,N_6904,N_6909);
nand U7209 (N_7209,N_6805,N_6791);
and U7210 (N_7210,N_6990,N_6833);
nor U7211 (N_7211,N_6911,N_6652);
xor U7212 (N_7212,N_6760,N_6668);
nor U7213 (N_7213,N_6651,N_6633);
and U7214 (N_7214,N_6515,N_6962);
nor U7215 (N_7215,N_6596,N_6506);
nor U7216 (N_7216,N_6925,N_6635);
or U7217 (N_7217,N_6739,N_6809);
and U7218 (N_7218,N_6799,N_6897);
and U7219 (N_7219,N_6557,N_6968);
xnor U7220 (N_7220,N_6819,N_6818);
nand U7221 (N_7221,N_6806,N_6580);
nand U7222 (N_7222,N_6757,N_6507);
and U7223 (N_7223,N_6711,N_6843);
and U7224 (N_7224,N_6717,N_6991);
or U7225 (N_7225,N_6963,N_6783);
xnor U7226 (N_7226,N_6747,N_6977);
nand U7227 (N_7227,N_6573,N_6752);
and U7228 (N_7228,N_6790,N_6970);
and U7229 (N_7229,N_6983,N_6691);
xor U7230 (N_7230,N_6856,N_6631);
and U7231 (N_7231,N_6520,N_6692);
and U7232 (N_7232,N_6565,N_6662);
nand U7233 (N_7233,N_6626,N_6745);
xor U7234 (N_7234,N_6649,N_6611);
or U7235 (N_7235,N_6831,N_6967);
or U7236 (N_7236,N_6639,N_6878);
or U7237 (N_7237,N_6654,N_6530);
or U7238 (N_7238,N_6961,N_6884);
nand U7239 (N_7239,N_6905,N_6607);
nor U7240 (N_7240,N_6942,N_6722);
xnor U7241 (N_7241,N_6655,N_6844);
xor U7242 (N_7242,N_6997,N_6776);
nor U7243 (N_7243,N_6561,N_6871);
xor U7244 (N_7244,N_6645,N_6887);
or U7245 (N_7245,N_6751,N_6556);
nand U7246 (N_7246,N_6786,N_6537);
nor U7247 (N_7247,N_6793,N_6714);
or U7248 (N_7248,N_6527,N_6761);
or U7249 (N_7249,N_6519,N_6746);
and U7250 (N_7250,N_6850,N_6532);
and U7251 (N_7251,N_6829,N_6813);
and U7252 (N_7252,N_6828,N_6942);
or U7253 (N_7253,N_6599,N_6668);
nor U7254 (N_7254,N_6950,N_6706);
nand U7255 (N_7255,N_6976,N_6825);
and U7256 (N_7256,N_6823,N_6614);
nor U7257 (N_7257,N_6804,N_6541);
xnor U7258 (N_7258,N_6975,N_6960);
nor U7259 (N_7259,N_6574,N_6686);
nor U7260 (N_7260,N_6668,N_6986);
nand U7261 (N_7261,N_6993,N_6749);
and U7262 (N_7262,N_6667,N_6765);
nor U7263 (N_7263,N_6913,N_6563);
or U7264 (N_7264,N_6972,N_6759);
nor U7265 (N_7265,N_6960,N_6605);
or U7266 (N_7266,N_6750,N_6860);
and U7267 (N_7267,N_6831,N_6878);
nand U7268 (N_7268,N_6583,N_6905);
or U7269 (N_7269,N_6960,N_6568);
and U7270 (N_7270,N_6848,N_6940);
and U7271 (N_7271,N_6958,N_6812);
and U7272 (N_7272,N_6686,N_6611);
and U7273 (N_7273,N_6816,N_6765);
and U7274 (N_7274,N_6964,N_6597);
nand U7275 (N_7275,N_6796,N_6829);
xnor U7276 (N_7276,N_6693,N_6956);
nand U7277 (N_7277,N_6782,N_6825);
and U7278 (N_7278,N_6983,N_6578);
nor U7279 (N_7279,N_6559,N_6752);
nor U7280 (N_7280,N_6765,N_6687);
or U7281 (N_7281,N_6772,N_6996);
xnor U7282 (N_7282,N_6822,N_6739);
and U7283 (N_7283,N_6693,N_6963);
nor U7284 (N_7284,N_6716,N_6770);
and U7285 (N_7285,N_6641,N_6905);
or U7286 (N_7286,N_6728,N_6924);
and U7287 (N_7287,N_6633,N_6635);
xnor U7288 (N_7288,N_6999,N_6660);
nand U7289 (N_7289,N_6855,N_6942);
or U7290 (N_7290,N_6595,N_6505);
nor U7291 (N_7291,N_6784,N_6659);
nor U7292 (N_7292,N_6734,N_6570);
nor U7293 (N_7293,N_6881,N_6897);
and U7294 (N_7294,N_6751,N_6508);
nor U7295 (N_7295,N_6708,N_6752);
xnor U7296 (N_7296,N_6836,N_6545);
or U7297 (N_7297,N_6688,N_6825);
xnor U7298 (N_7298,N_6727,N_6595);
nand U7299 (N_7299,N_6985,N_6764);
nor U7300 (N_7300,N_6955,N_6793);
or U7301 (N_7301,N_6767,N_6837);
and U7302 (N_7302,N_6854,N_6907);
or U7303 (N_7303,N_6676,N_6906);
and U7304 (N_7304,N_6797,N_6706);
or U7305 (N_7305,N_6785,N_6767);
or U7306 (N_7306,N_6757,N_6815);
xor U7307 (N_7307,N_6745,N_6784);
nand U7308 (N_7308,N_6614,N_6732);
and U7309 (N_7309,N_6919,N_6538);
or U7310 (N_7310,N_6851,N_6534);
xor U7311 (N_7311,N_6801,N_6600);
nand U7312 (N_7312,N_6642,N_6765);
xnor U7313 (N_7313,N_6866,N_6775);
nor U7314 (N_7314,N_6652,N_6820);
nor U7315 (N_7315,N_6895,N_6928);
or U7316 (N_7316,N_6872,N_6554);
and U7317 (N_7317,N_6717,N_6633);
nand U7318 (N_7318,N_6852,N_6816);
or U7319 (N_7319,N_6723,N_6819);
xnor U7320 (N_7320,N_6915,N_6596);
or U7321 (N_7321,N_6802,N_6735);
or U7322 (N_7322,N_6645,N_6987);
and U7323 (N_7323,N_6702,N_6802);
nor U7324 (N_7324,N_6563,N_6905);
or U7325 (N_7325,N_6692,N_6529);
nand U7326 (N_7326,N_6907,N_6736);
xor U7327 (N_7327,N_6785,N_6723);
and U7328 (N_7328,N_6994,N_6990);
and U7329 (N_7329,N_6574,N_6980);
nand U7330 (N_7330,N_6724,N_6764);
and U7331 (N_7331,N_6817,N_6608);
nor U7332 (N_7332,N_6980,N_6511);
and U7333 (N_7333,N_6797,N_6843);
nor U7334 (N_7334,N_6528,N_6694);
or U7335 (N_7335,N_6884,N_6798);
nand U7336 (N_7336,N_6732,N_6809);
xor U7337 (N_7337,N_6585,N_6844);
xor U7338 (N_7338,N_6552,N_6958);
nand U7339 (N_7339,N_6823,N_6581);
or U7340 (N_7340,N_6641,N_6668);
and U7341 (N_7341,N_6566,N_6903);
and U7342 (N_7342,N_6754,N_6553);
xnor U7343 (N_7343,N_6919,N_6735);
nand U7344 (N_7344,N_6971,N_6678);
xnor U7345 (N_7345,N_6878,N_6706);
nor U7346 (N_7346,N_6679,N_6795);
nand U7347 (N_7347,N_6643,N_6992);
or U7348 (N_7348,N_6693,N_6528);
xor U7349 (N_7349,N_6529,N_6761);
xnor U7350 (N_7350,N_6595,N_6713);
nand U7351 (N_7351,N_6599,N_6706);
nand U7352 (N_7352,N_6573,N_6853);
nor U7353 (N_7353,N_6968,N_6667);
xor U7354 (N_7354,N_6547,N_6698);
nand U7355 (N_7355,N_6656,N_6827);
or U7356 (N_7356,N_6563,N_6595);
and U7357 (N_7357,N_6559,N_6519);
and U7358 (N_7358,N_6992,N_6659);
nand U7359 (N_7359,N_6966,N_6851);
xor U7360 (N_7360,N_6632,N_6549);
nor U7361 (N_7361,N_6728,N_6516);
and U7362 (N_7362,N_6669,N_6873);
and U7363 (N_7363,N_6525,N_6748);
nor U7364 (N_7364,N_6543,N_6999);
and U7365 (N_7365,N_6980,N_6925);
nand U7366 (N_7366,N_6895,N_6610);
and U7367 (N_7367,N_6971,N_6671);
nor U7368 (N_7368,N_6641,N_6566);
xnor U7369 (N_7369,N_6928,N_6595);
and U7370 (N_7370,N_6749,N_6873);
nor U7371 (N_7371,N_6676,N_6823);
xnor U7372 (N_7372,N_6545,N_6711);
nand U7373 (N_7373,N_6779,N_6519);
nand U7374 (N_7374,N_6519,N_6724);
or U7375 (N_7375,N_6956,N_6676);
nand U7376 (N_7376,N_6965,N_6671);
and U7377 (N_7377,N_6664,N_6525);
and U7378 (N_7378,N_6764,N_6911);
and U7379 (N_7379,N_6854,N_6710);
or U7380 (N_7380,N_6784,N_6632);
xnor U7381 (N_7381,N_6806,N_6990);
nand U7382 (N_7382,N_6860,N_6591);
or U7383 (N_7383,N_6707,N_6601);
and U7384 (N_7384,N_6637,N_6819);
xnor U7385 (N_7385,N_6772,N_6720);
xor U7386 (N_7386,N_6811,N_6606);
nor U7387 (N_7387,N_6714,N_6874);
nand U7388 (N_7388,N_6512,N_6519);
and U7389 (N_7389,N_6512,N_6749);
nand U7390 (N_7390,N_6923,N_6961);
and U7391 (N_7391,N_6774,N_6912);
nand U7392 (N_7392,N_6898,N_6737);
nand U7393 (N_7393,N_6609,N_6824);
nor U7394 (N_7394,N_6888,N_6599);
or U7395 (N_7395,N_6642,N_6517);
or U7396 (N_7396,N_6829,N_6668);
nand U7397 (N_7397,N_6690,N_6600);
nor U7398 (N_7398,N_6791,N_6971);
and U7399 (N_7399,N_6722,N_6840);
and U7400 (N_7400,N_6884,N_6969);
nor U7401 (N_7401,N_6725,N_6665);
and U7402 (N_7402,N_6722,N_6600);
nand U7403 (N_7403,N_6764,N_6609);
or U7404 (N_7404,N_6932,N_6696);
or U7405 (N_7405,N_6731,N_6512);
nor U7406 (N_7406,N_6528,N_6705);
xor U7407 (N_7407,N_6609,N_6886);
nor U7408 (N_7408,N_6774,N_6968);
nand U7409 (N_7409,N_6996,N_6677);
nor U7410 (N_7410,N_6929,N_6685);
xnor U7411 (N_7411,N_6768,N_6895);
nand U7412 (N_7412,N_6525,N_6677);
nand U7413 (N_7413,N_6861,N_6875);
nand U7414 (N_7414,N_6867,N_6875);
nand U7415 (N_7415,N_6725,N_6527);
xor U7416 (N_7416,N_6995,N_6566);
nor U7417 (N_7417,N_6920,N_6640);
nor U7418 (N_7418,N_6637,N_6601);
nand U7419 (N_7419,N_6923,N_6980);
or U7420 (N_7420,N_6780,N_6873);
and U7421 (N_7421,N_6790,N_6686);
nand U7422 (N_7422,N_6613,N_6850);
and U7423 (N_7423,N_6760,N_6649);
nor U7424 (N_7424,N_6679,N_6812);
and U7425 (N_7425,N_6917,N_6615);
nor U7426 (N_7426,N_6961,N_6913);
nor U7427 (N_7427,N_6737,N_6775);
nand U7428 (N_7428,N_6811,N_6934);
or U7429 (N_7429,N_6759,N_6862);
nor U7430 (N_7430,N_6750,N_6695);
nand U7431 (N_7431,N_6963,N_6913);
or U7432 (N_7432,N_6929,N_6528);
xnor U7433 (N_7433,N_6758,N_6820);
nand U7434 (N_7434,N_6809,N_6706);
xnor U7435 (N_7435,N_6928,N_6926);
or U7436 (N_7436,N_6561,N_6788);
nor U7437 (N_7437,N_6500,N_6904);
and U7438 (N_7438,N_6832,N_6564);
or U7439 (N_7439,N_6780,N_6729);
and U7440 (N_7440,N_6570,N_6908);
and U7441 (N_7441,N_6755,N_6700);
nor U7442 (N_7442,N_6787,N_6966);
and U7443 (N_7443,N_6877,N_6762);
xor U7444 (N_7444,N_6868,N_6966);
nand U7445 (N_7445,N_6796,N_6848);
nand U7446 (N_7446,N_6905,N_6577);
or U7447 (N_7447,N_6748,N_6800);
nor U7448 (N_7448,N_6731,N_6669);
nand U7449 (N_7449,N_6731,N_6690);
nor U7450 (N_7450,N_6566,N_6841);
nor U7451 (N_7451,N_6949,N_6599);
or U7452 (N_7452,N_6997,N_6876);
and U7453 (N_7453,N_6779,N_6699);
and U7454 (N_7454,N_6780,N_6604);
and U7455 (N_7455,N_6596,N_6844);
or U7456 (N_7456,N_6939,N_6890);
nor U7457 (N_7457,N_6584,N_6664);
or U7458 (N_7458,N_6703,N_6720);
nand U7459 (N_7459,N_6929,N_6784);
nor U7460 (N_7460,N_6774,N_6637);
nand U7461 (N_7461,N_6773,N_6698);
nand U7462 (N_7462,N_6832,N_6982);
and U7463 (N_7463,N_6543,N_6597);
nor U7464 (N_7464,N_6778,N_6929);
xor U7465 (N_7465,N_6936,N_6782);
nor U7466 (N_7466,N_6903,N_6780);
or U7467 (N_7467,N_6835,N_6896);
nor U7468 (N_7468,N_6848,N_6699);
xor U7469 (N_7469,N_6556,N_6525);
nor U7470 (N_7470,N_6857,N_6513);
nand U7471 (N_7471,N_6878,N_6994);
and U7472 (N_7472,N_6854,N_6762);
or U7473 (N_7473,N_6570,N_6666);
and U7474 (N_7474,N_6787,N_6535);
and U7475 (N_7475,N_6619,N_6638);
nor U7476 (N_7476,N_6751,N_6510);
or U7477 (N_7477,N_6943,N_6537);
nor U7478 (N_7478,N_6633,N_6694);
nand U7479 (N_7479,N_6706,N_6866);
and U7480 (N_7480,N_6824,N_6547);
nor U7481 (N_7481,N_6817,N_6774);
nand U7482 (N_7482,N_6643,N_6965);
nand U7483 (N_7483,N_6645,N_6852);
nand U7484 (N_7484,N_6553,N_6552);
and U7485 (N_7485,N_6506,N_6587);
or U7486 (N_7486,N_6627,N_6743);
nand U7487 (N_7487,N_6905,N_6982);
nand U7488 (N_7488,N_6951,N_6723);
nor U7489 (N_7489,N_6587,N_6827);
and U7490 (N_7490,N_6892,N_6950);
nand U7491 (N_7491,N_6920,N_6778);
nor U7492 (N_7492,N_6768,N_6966);
or U7493 (N_7493,N_6975,N_6820);
nand U7494 (N_7494,N_6809,N_6787);
nand U7495 (N_7495,N_6940,N_6955);
nand U7496 (N_7496,N_6804,N_6768);
or U7497 (N_7497,N_6869,N_6738);
nor U7498 (N_7498,N_6699,N_6747);
and U7499 (N_7499,N_6920,N_6600);
nand U7500 (N_7500,N_7067,N_7435);
or U7501 (N_7501,N_7429,N_7446);
or U7502 (N_7502,N_7102,N_7253);
xnor U7503 (N_7503,N_7337,N_7191);
and U7504 (N_7504,N_7027,N_7257);
nand U7505 (N_7505,N_7388,N_7270);
nor U7506 (N_7506,N_7148,N_7371);
xor U7507 (N_7507,N_7251,N_7195);
nand U7508 (N_7508,N_7013,N_7322);
or U7509 (N_7509,N_7202,N_7350);
or U7510 (N_7510,N_7121,N_7294);
and U7511 (N_7511,N_7053,N_7050);
nand U7512 (N_7512,N_7291,N_7106);
nand U7513 (N_7513,N_7184,N_7468);
and U7514 (N_7514,N_7002,N_7494);
and U7515 (N_7515,N_7036,N_7323);
and U7516 (N_7516,N_7464,N_7223);
and U7517 (N_7517,N_7096,N_7345);
nor U7518 (N_7518,N_7135,N_7165);
nor U7519 (N_7519,N_7153,N_7230);
or U7520 (N_7520,N_7144,N_7343);
xor U7521 (N_7521,N_7437,N_7283);
and U7522 (N_7522,N_7387,N_7383);
xnor U7523 (N_7523,N_7489,N_7240);
or U7524 (N_7524,N_7373,N_7031);
and U7525 (N_7525,N_7344,N_7335);
or U7526 (N_7526,N_7288,N_7427);
or U7527 (N_7527,N_7124,N_7378);
and U7528 (N_7528,N_7136,N_7442);
nand U7529 (N_7529,N_7439,N_7089);
nand U7530 (N_7530,N_7358,N_7363);
or U7531 (N_7531,N_7414,N_7222);
nand U7532 (N_7532,N_7411,N_7483);
nand U7533 (N_7533,N_7110,N_7271);
or U7534 (N_7534,N_7095,N_7274);
nor U7535 (N_7535,N_7267,N_7317);
nand U7536 (N_7536,N_7187,N_7478);
or U7537 (N_7537,N_7289,N_7134);
nand U7538 (N_7538,N_7086,N_7261);
nor U7539 (N_7539,N_7269,N_7349);
or U7540 (N_7540,N_7171,N_7119);
xor U7541 (N_7541,N_7475,N_7448);
and U7542 (N_7542,N_7168,N_7318);
and U7543 (N_7543,N_7145,N_7149);
nor U7544 (N_7544,N_7329,N_7122);
or U7545 (N_7545,N_7452,N_7120);
nand U7546 (N_7546,N_7417,N_7028);
and U7547 (N_7547,N_7212,N_7425);
and U7548 (N_7548,N_7381,N_7405);
or U7549 (N_7549,N_7104,N_7037);
nand U7550 (N_7550,N_7156,N_7476);
nand U7551 (N_7551,N_7473,N_7313);
nand U7552 (N_7552,N_7008,N_7142);
nand U7553 (N_7553,N_7484,N_7377);
nand U7554 (N_7554,N_7308,N_7192);
and U7555 (N_7555,N_7232,N_7210);
or U7556 (N_7556,N_7055,N_7157);
nor U7557 (N_7557,N_7266,N_7118);
xnor U7558 (N_7558,N_7433,N_7457);
nor U7559 (N_7559,N_7301,N_7091);
nor U7560 (N_7560,N_7175,N_7268);
nor U7561 (N_7561,N_7022,N_7430);
xor U7562 (N_7562,N_7169,N_7461);
nor U7563 (N_7563,N_7048,N_7341);
nand U7564 (N_7564,N_7088,N_7237);
and U7565 (N_7565,N_7131,N_7493);
nand U7566 (N_7566,N_7176,N_7282);
and U7567 (N_7567,N_7005,N_7458);
nand U7568 (N_7568,N_7426,N_7316);
or U7569 (N_7569,N_7077,N_7178);
nor U7570 (N_7570,N_7382,N_7044);
nor U7571 (N_7571,N_7141,N_7256);
nand U7572 (N_7572,N_7233,N_7200);
xor U7573 (N_7573,N_7273,N_7026);
and U7574 (N_7574,N_7278,N_7471);
or U7575 (N_7575,N_7391,N_7432);
nand U7576 (N_7576,N_7115,N_7482);
nand U7577 (N_7577,N_7113,N_7047);
nand U7578 (N_7578,N_7172,N_7163);
or U7579 (N_7579,N_7132,N_7205);
nand U7580 (N_7580,N_7087,N_7216);
nand U7581 (N_7581,N_7190,N_7114);
and U7582 (N_7582,N_7249,N_7389);
nand U7583 (N_7583,N_7443,N_7182);
and U7584 (N_7584,N_7444,N_7059);
or U7585 (N_7585,N_7219,N_7060);
nand U7586 (N_7586,N_7162,N_7263);
nand U7587 (N_7587,N_7133,N_7260);
or U7588 (N_7588,N_7398,N_7465);
or U7589 (N_7589,N_7409,N_7150);
and U7590 (N_7590,N_7072,N_7220);
and U7591 (N_7591,N_7231,N_7364);
nand U7592 (N_7592,N_7147,N_7459);
nand U7593 (N_7593,N_7116,N_7472);
or U7594 (N_7594,N_7392,N_7319);
nor U7595 (N_7595,N_7075,N_7183);
nor U7596 (N_7596,N_7185,N_7057);
and U7597 (N_7597,N_7030,N_7339);
nand U7598 (N_7598,N_7495,N_7040);
xor U7599 (N_7599,N_7234,N_7338);
xnor U7600 (N_7600,N_7159,N_7491);
nand U7601 (N_7601,N_7453,N_7369);
and U7602 (N_7602,N_7440,N_7245);
or U7603 (N_7603,N_7211,N_7297);
nand U7604 (N_7604,N_7361,N_7360);
nor U7605 (N_7605,N_7431,N_7352);
nor U7606 (N_7606,N_7395,N_7239);
nor U7607 (N_7607,N_7138,N_7177);
or U7608 (N_7608,N_7385,N_7023);
nand U7609 (N_7609,N_7259,N_7347);
nor U7610 (N_7610,N_7334,N_7073);
xor U7611 (N_7611,N_7038,N_7451);
or U7612 (N_7612,N_7214,N_7324);
or U7613 (N_7613,N_7128,N_7217);
nand U7614 (N_7614,N_7406,N_7054);
nand U7615 (N_7615,N_7342,N_7137);
and U7616 (N_7616,N_7112,N_7094);
xnor U7617 (N_7617,N_7080,N_7359);
or U7618 (N_7618,N_7330,N_7085);
nand U7619 (N_7619,N_7079,N_7011);
nor U7620 (N_7620,N_7333,N_7332);
nor U7621 (N_7621,N_7170,N_7227);
nor U7622 (N_7622,N_7328,N_7246);
nand U7623 (N_7623,N_7151,N_7296);
nand U7624 (N_7624,N_7140,N_7481);
nor U7625 (N_7625,N_7479,N_7236);
or U7626 (N_7626,N_7033,N_7196);
nand U7627 (N_7627,N_7413,N_7092);
nand U7628 (N_7628,N_7445,N_7416);
nand U7629 (N_7629,N_7423,N_7203);
nand U7630 (N_7630,N_7139,N_7229);
xnor U7631 (N_7631,N_7181,N_7407);
or U7632 (N_7632,N_7298,N_7194);
and U7633 (N_7633,N_7064,N_7455);
or U7634 (N_7634,N_7415,N_7056);
or U7635 (N_7635,N_7404,N_7068);
xnor U7636 (N_7636,N_7017,N_7370);
nor U7637 (N_7637,N_7126,N_7403);
nand U7638 (N_7638,N_7093,N_7254);
and U7639 (N_7639,N_7412,N_7469);
or U7640 (N_7640,N_7486,N_7143);
nor U7641 (N_7641,N_7300,N_7252);
or U7642 (N_7642,N_7366,N_7420);
and U7643 (N_7643,N_7204,N_7146);
and U7644 (N_7644,N_7496,N_7419);
and U7645 (N_7645,N_7326,N_7111);
or U7646 (N_7646,N_7401,N_7250);
nor U7647 (N_7647,N_7394,N_7109);
nor U7648 (N_7648,N_7123,N_7428);
or U7649 (N_7649,N_7365,N_7315);
nor U7650 (N_7650,N_7228,N_7006);
and U7651 (N_7651,N_7155,N_7167);
nor U7652 (N_7652,N_7255,N_7390);
and U7653 (N_7653,N_7325,N_7215);
nor U7654 (N_7654,N_7348,N_7065);
xnor U7655 (N_7655,N_7293,N_7490);
nand U7656 (N_7656,N_7393,N_7025);
nand U7657 (N_7657,N_7016,N_7275);
nand U7658 (N_7658,N_7499,N_7010);
nor U7659 (N_7659,N_7331,N_7374);
nor U7660 (N_7660,N_7083,N_7173);
and U7661 (N_7661,N_7043,N_7336);
nand U7662 (N_7662,N_7277,N_7280);
nor U7663 (N_7663,N_7052,N_7058);
nor U7664 (N_7664,N_7379,N_7105);
nand U7665 (N_7665,N_7353,N_7243);
and U7666 (N_7666,N_7356,N_7117);
nor U7667 (N_7667,N_7265,N_7049);
or U7668 (N_7668,N_7004,N_7450);
xor U7669 (N_7669,N_7281,N_7474);
nor U7670 (N_7670,N_7497,N_7480);
nor U7671 (N_7671,N_7303,N_7076);
nor U7672 (N_7672,N_7470,N_7287);
and U7673 (N_7673,N_7090,N_7161);
nand U7674 (N_7674,N_7351,N_7197);
or U7675 (N_7675,N_7380,N_7107);
or U7676 (N_7676,N_7295,N_7041);
xnor U7677 (N_7677,N_7180,N_7456);
nor U7678 (N_7678,N_7018,N_7305);
nor U7679 (N_7679,N_7154,N_7264);
nand U7680 (N_7680,N_7462,N_7032);
or U7681 (N_7681,N_7447,N_7129);
nand U7682 (N_7682,N_7368,N_7396);
nand U7683 (N_7683,N_7258,N_7436);
or U7684 (N_7684,N_7001,N_7320);
or U7685 (N_7685,N_7046,N_7063);
nand U7686 (N_7686,N_7125,N_7158);
nand U7687 (N_7687,N_7312,N_7221);
nor U7688 (N_7688,N_7224,N_7367);
nand U7689 (N_7689,N_7101,N_7164);
and U7690 (N_7690,N_7186,N_7492);
nand U7691 (N_7691,N_7286,N_7012);
nor U7692 (N_7692,N_7242,N_7020);
and U7693 (N_7693,N_7103,N_7069);
or U7694 (N_7694,N_7238,N_7130);
and U7695 (N_7695,N_7386,N_7188);
or U7696 (N_7696,N_7007,N_7201);
nand U7697 (N_7697,N_7179,N_7304);
nor U7698 (N_7698,N_7071,N_7310);
and U7699 (N_7699,N_7424,N_7397);
and U7700 (N_7700,N_7463,N_7421);
nand U7701 (N_7701,N_7015,N_7160);
or U7702 (N_7702,N_7019,N_7021);
xor U7703 (N_7703,N_7285,N_7003);
nand U7704 (N_7704,N_7070,N_7066);
nand U7705 (N_7705,N_7247,N_7399);
nand U7706 (N_7706,N_7354,N_7262);
nand U7707 (N_7707,N_7039,N_7209);
or U7708 (N_7708,N_7108,N_7248);
nor U7709 (N_7709,N_7174,N_7078);
and U7710 (N_7710,N_7098,N_7000);
or U7711 (N_7711,N_7485,N_7309);
nand U7712 (N_7712,N_7290,N_7488);
or U7713 (N_7713,N_7084,N_7081);
nand U7714 (N_7714,N_7498,N_7376);
and U7715 (N_7715,N_7042,N_7438);
xnor U7716 (N_7716,N_7166,N_7082);
and U7717 (N_7717,N_7357,N_7099);
and U7718 (N_7718,N_7127,N_7418);
xor U7719 (N_7719,N_7311,N_7226);
nor U7720 (N_7720,N_7218,N_7284);
and U7721 (N_7721,N_7074,N_7346);
or U7722 (N_7722,N_7400,N_7410);
nand U7723 (N_7723,N_7279,N_7307);
or U7724 (N_7724,N_7340,N_7276);
nor U7725 (N_7725,N_7235,N_7207);
xnor U7726 (N_7726,N_7299,N_7208);
and U7727 (N_7727,N_7213,N_7024);
or U7728 (N_7728,N_7062,N_7355);
xnor U7729 (N_7729,N_7384,N_7292);
and U7730 (N_7730,N_7051,N_7206);
or U7731 (N_7731,N_7408,N_7375);
nand U7732 (N_7732,N_7422,N_7272);
nor U7733 (N_7733,N_7402,N_7045);
or U7734 (N_7734,N_7314,N_7189);
and U7735 (N_7735,N_7014,N_7034);
nor U7736 (N_7736,N_7372,N_7302);
or U7737 (N_7737,N_7454,N_7306);
nor U7738 (N_7738,N_7244,N_7362);
or U7739 (N_7739,N_7241,N_7152);
and U7740 (N_7740,N_7434,N_7199);
nor U7741 (N_7741,N_7061,N_7097);
and U7742 (N_7742,N_7009,N_7449);
nor U7743 (N_7743,N_7441,N_7327);
nor U7744 (N_7744,N_7467,N_7487);
nor U7745 (N_7745,N_7321,N_7460);
or U7746 (N_7746,N_7225,N_7477);
nor U7747 (N_7747,N_7100,N_7035);
and U7748 (N_7748,N_7193,N_7466);
nor U7749 (N_7749,N_7198,N_7029);
nand U7750 (N_7750,N_7216,N_7057);
nand U7751 (N_7751,N_7083,N_7373);
nand U7752 (N_7752,N_7253,N_7266);
or U7753 (N_7753,N_7293,N_7150);
xor U7754 (N_7754,N_7455,N_7437);
nand U7755 (N_7755,N_7235,N_7282);
nand U7756 (N_7756,N_7140,N_7453);
and U7757 (N_7757,N_7199,N_7222);
nand U7758 (N_7758,N_7374,N_7307);
and U7759 (N_7759,N_7235,N_7279);
and U7760 (N_7760,N_7498,N_7145);
xor U7761 (N_7761,N_7073,N_7306);
nand U7762 (N_7762,N_7150,N_7424);
xnor U7763 (N_7763,N_7068,N_7217);
nand U7764 (N_7764,N_7257,N_7018);
nor U7765 (N_7765,N_7277,N_7234);
nand U7766 (N_7766,N_7437,N_7499);
and U7767 (N_7767,N_7396,N_7160);
or U7768 (N_7768,N_7371,N_7008);
or U7769 (N_7769,N_7445,N_7085);
and U7770 (N_7770,N_7250,N_7424);
or U7771 (N_7771,N_7392,N_7024);
nor U7772 (N_7772,N_7404,N_7354);
and U7773 (N_7773,N_7388,N_7047);
nor U7774 (N_7774,N_7133,N_7248);
xnor U7775 (N_7775,N_7264,N_7463);
xor U7776 (N_7776,N_7056,N_7256);
nand U7777 (N_7777,N_7124,N_7346);
xnor U7778 (N_7778,N_7341,N_7454);
nand U7779 (N_7779,N_7317,N_7245);
or U7780 (N_7780,N_7057,N_7103);
nand U7781 (N_7781,N_7460,N_7191);
nand U7782 (N_7782,N_7345,N_7491);
or U7783 (N_7783,N_7406,N_7124);
nand U7784 (N_7784,N_7008,N_7109);
nor U7785 (N_7785,N_7415,N_7253);
nor U7786 (N_7786,N_7436,N_7260);
or U7787 (N_7787,N_7009,N_7092);
nand U7788 (N_7788,N_7028,N_7101);
nor U7789 (N_7789,N_7284,N_7439);
nand U7790 (N_7790,N_7011,N_7114);
nor U7791 (N_7791,N_7400,N_7373);
nor U7792 (N_7792,N_7315,N_7012);
and U7793 (N_7793,N_7159,N_7137);
nor U7794 (N_7794,N_7354,N_7021);
nand U7795 (N_7795,N_7250,N_7209);
or U7796 (N_7796,N_7370,N_7072);
nor U7797 (N_7797,N_7067,N_7203);
nor U7798 (N_7798,N_7148,N_7127);
nor U7799 (N_7799,N_7210,N_7265);
and U7800 (N_7800,N_7352,N_7087);
and U7801 (N_7801,N_7402,N_7428);
and U7802 (N_7802,N_7238,N_7302);
nor U7803 (N_7803,N_7237,N_7087);
or U7804 (N_7804,N_7412,N_7117);
nor U7805 (N_7805,N_7479,N_7086);
and U7806 (N_7806,N_7279,N_7238);
and U7807 (N_7807,N_7183,N_7290);
or U7808 (N_7808,N_7104,N_7040);
and U7809 (N_7809,N_7491,N_7121);
nand U7810 (N_7810,N_7364,N_7037);
and U7811 (N_7811,N_7062,N_7085);
xor U7812 (N_7812,N_7370,N_7381);
nor U7813 (N_7813,N_7295,N_7221);
nor U7814 (N_7814,N_7328,N_7322);
xor U7815 (N_7815,N_7402,N_7060);
nor U7816 (N_7816,N_7469,N_7368);
nand U7817 (N_7817,N_7395,N_7119);
or U7818 (N_7818,N_7349,N_7376);
nor U7819 (N_7819,N_7214,N_7134);
nand U7820 (N_7820,N_7141,N_7453);
and U7821 (N_7821,N_7247,N_7384);
nand U7822 (N_7822,N_7270,N_7150);
nor U7823 (N_7823,N_7353,N_7444);
xnor U7824 (N_7824,N_7433,N_7424);
nor U7825 (N_7825,N_7483,N_7418);
nor U7826 (N_7826,N_7162,N_7234);
nand U7827 (N_7827,N_7394,N_7040);
or U7828 (N_7828,N_7429,N_7142);
nor U7829 (N_7829,N_7404,N_7169);
xnor U7830 (N_7830,N_7360,N_7144);
or U7831 (N_7831,N_7403,N_7281);
xor U7832 (N_7832,N_7245,N_7367);
or U7833 (N_7833,N_7246,N_7191);
nor U7834 (N_7834,N_7056,N_7419);
nand U7835 (N_7835,N_7382,N_7142);
or U7836 (N_7836,N_7435,N_7367);
nand U7837 (N_7837,N_7375,N_7052);
nor U7838 (N_7838,N_7461,N_7261);
or U7839 (N_7839,N_7016,N_7181);
nand U7840 (N_7840,N_7030,N_7483);
or U7841 (N_7841,N_7096,N_7326);
nand U7842 (N_7842,N_7179,N_7281);
or U7843 (N_7843,N_7287,N_7313);
nand U7844 (N_7844,N_7155,N_7074);
or U7845 (N_7845,N_7361,N_7183);
nand U7846 (N_7846,N_7343,N_7239);
xor U7847 (N_7847,N_7455,N_7024);
nor U7848 (N_7848,N_7205,N_7126);
nand U7849 (N_7849,N_7223,N_7118);
and U7850 (N_7850,N_7222,N_7268);
or U7851 (N_7851,N_7492,N_7278);
and U7852 (N_7852,N_7019,N_7155);
xor U7853 (N_7853,N_7176,N_7232);
or U7854 (N_7854,N_7121,N_7215);
nand U7855 (N_7855,N_7064,N_7458);
nand U7856 (N_7856,N_7139,N_7178);
or U7857 (N_7857,N_7401,N_7265);
and U7858 (N_7858,N_7496,N_7262);
nand U7859 (N_7859,N_7386,N_7165);
xor U7860 (N_7860,N_7034,N_7318);
xor U7861 (N_7861,N_7239,N_7170);
nor U7862 (N_7862,N_7013,N_7167);
nand U7863 (N_7863,N_7371,N_7363);
or U7864 (N_7864,N_7418,N_7342);
nand U7865 (N_7865,N_7479,N_7316);
nor U7866 (N_7866,N_7335,N_7231);
xnor U7867 (N_7867,N_7130,N_7439);
nor U7868 (N_7868,N_7484,N_7160);
and U7869 (N_7869,N_7142,N_7243);
and U7870 (N_7870,N_7456,N_7306);
nor U7871 (N_7871,N_7428,N_7027);
or U7872 (N_7872,N_7243,N_7471);
xor U7873 (N_7873,N_7411,N_7449);
or U7874 (N_7874,N_7423,N_7493);
nand U7875 (N_7875,N_7225,N_7172);
nand U7876 (N_7876,N_7347,N_7492);
nor U7877 (N_7877,N_7330,N_7141);
or U7878 (N_7878,N_7134,N_7171);
or U7879 (N_7879,N_7048,N_7025);
nor U7880 (N_7880,N_7070,N_7376);
or U7881 (N_7881,N_7071,N_7147);
and U7882 (N_7882,N_7248,N_7065);
xor U7883 (N_7883,N_7326,N_7478);
and U7884 (N_7884,N_7004,N_7292);
xor U7885 (N_7885,N_7068,N_7408);
or U7886 (N_7886,N_7207,N_7438);
or U7887 (N_7887,N_7127,N_7419);
nor U7888 (N_7888,N_7009,N_7305);
or U7889 (N_7889,N_7105,N_7258);
and U7890 (N_7890,N_7183,N_7161);
nand U7891 (N_7891,N_7233,N_7093);
nor U7892 (N_7892,N_7413,N_7385);
and U7893 (N_7893,N_7012,N_7138);
nor U7894 (N_7894,N_7334,N_7155);
nand U7895 (N_7895,N_7122,N_7393);
and U7896 (N_7896,N_7456,N_7163);
or U7897 (N_7897,N_7358,N_7197);
xnor U7898 (N_7898,N_7217,N_7239);
nand U7899 (N_7899,N_7069,N_7327);
nand U7900 (N_7900,N_7238,N_7158);
nor U7901 (N_7901,N_7288,N_7175);
or U7902 (N_7902,N_7139,N_7079);
nor U7903 (N_7903,N_7439,N_7461);
nand U7904 (N_7904,N_7223,N_7150);
or U7905 (N_7905,N_7154,N_7432);
xnor U7906 (N_7906,N_7310,N_7123);
or U7907 (N_7907,N_7187,N_7005);
nor U7908 (N_7908,N_7164,N_7040);
and U7909 (N_7909,N_7370,N_7380);
xnor U7910 (N_7910,N_7070,N_7199);
and U7911 (N_7911,N_7164,N_7123);
or U7912 (N_7912,N_7323,N_7498);
or U7913 (N_7913,N_7211,N_7373);
or U7914 (N_7914,N_7216,N_7005);
and U7915 (N_7915,N_7472,N_7145);
nand U7916 (N_7916,N_7377,N_7353);
and U7917 (N_7917,N_7200,N_7335);
nor U7918 (N_7918,N_7453,N_7262);
nand U7919 (N_7919,N_7213,N_7306);
nand U7920 (N_7920,N_7299,N_7058);
or U7921 (N_7921,N_7074,N_7313);
nand U7922 (N_7922,N_7073,N_7186);
nor U7923 (N_7923,N_7102,N_7143);
nand U7924 (N_7924,N_7355,N_7296);
and U7925 (N_7925,N_7218,N_7212);
and U7926 (N_7926,N_7420,N_7028);
nand U7927 (N_7927,N_7395,N_7289);
and U7928 (N_7928,N_7079,N_7337);
and U7929 (N_7929,N_7187,N_7314);
nand U7930 (N_7930,N_7292,N_7298);
nand U7931 (N_7931,N_7401,N_7026);
nand U7932 (N_7932,N_7456,N_7336);
nand U7933 (N_7933,N_7225,N_7170);
nand U7934 (N_7934,N_7010,N_7122);
or U7935 (N_7935,N_7227,N_7242);
xor U7936 (N_7936,N_7148,N_7472);
xnor U7937 (N_7937,N_7084,N_7029);
and U7938 (N_7938,N_7486,N_7331);
and U7939 (N_7939,N_7278,N_7191);
and U7940 (N_7940,N_7297,N_7480);
and U7941 (N_7941,N_7485,N_7240);
nor U7942 (N_7942,N_7202,N_7487);
nor U7943 (N_7943,N_7068,N_7055);
and U7944 (N_7944,N_7150,N_7137);
and U7945 (N_7945,N_7444,N_7295);
and U7946 (N_7946,N_7419,N_7389);
nor U7947 (N_7947,N_7143,N_7289);
and U7948 (N_7948,N_7046,N_7187);
xnor U7949 (N_7949,N_7146,N_7337);
nor U7950 (N_7950,N_7183,N_7104);
or U7951 (N_7951,N_7459,N_7338);
and U7952 (N_7952,N_7498,N_7228);
nand U7953 (N_7953,N_7145,N_7353);
nor U7954 (N_7954,N_7430,N_7299);
nor U7955 (N_7955,N_7341,N_7103);
or U7956 (N_7956,N_7163,N_7156);
or U7957 (N_7957,N_7214,N_7123);
and U7958 (N_7958,N_7318,N_7499);
or U7959 (N_7959,N_7393,N_7453);
or U7960 (N_7960,N_7216,N_7224);
nor U7961 (N_7961,N_7304,N_7302);
and U7962 (N_7962,N_7026,N_7463);
nand U7963 (N_7963,N_7040,N_7093);
and U7964 (N_7964,N_7288,N_7095);
nand U7965 (N_7965,N_7425,N_7123);
or U7966 (N_7966,N_7469,N_7170);
nor U7967 (N_7967,N_7231,N_7460);
xor U7968 (N_7968,N_7235,N_7015);
xnor U7969 (N_7969,N_7123,N_7035);
or U7970 (N_7970,N_7134,N_7343);
nand U7971 (N_7971,N_7481,N_7082);
or U7972 (N_7972,N_7217,N_7269);
and U7973 (N_7973,N_7319,N_7227);
xor U7974 (N_7974,N_7357,N_7472);
xor U7975 (N_7975,N_7114,N_7431);
nand U7976 (N_7976,N_7185,N_7086);
or U7977 (N_7977,N_7285,N_7376);
nand U7978 (N_7978,N_7029,N_7256);
xor U7979 (N_7979,N_7429,N_7416);
nor U7980 (N_7980,N_7182,N_7437);
nand U7981 (N_7981,N_7000,N_7392);
xnor U7982 (N_7982,N_7335,N_7384);
nor U7983 (N_7983,N_7440,N_7317);
xor U7984 (N_7984,N_7124,N_7070);
nor U7985 (N_7985,N_7247,N_7099);
nor U7986 (N_7986,N_7338,N_7341);
and U7987 (N_7987,N_7363,N_7246);
nand U7988 (N_7988,N_7201,N_7309);
nand U7989 (N_7989,N_7328,N_7389);
and U7990 (N_7990,N_7194,N_7339);
xnor U7991 (N_7991,N_7326,N_7392);
xnor U7992 (N_7992,N_7013,N_7395);
xnor U7993 (N_7993,N_7426,N_7186);
nand U7994 (N_7994,N_7364,N_7071);
xnor U7995 (N_7995,N_7388,N_7368);
nor U7996 (N_7996,N_7394,N_7042);
nand U7997 (N_7997,N_7076,N_7213);
nor U7998 (N_7998,N_7057,N_7226);
and U7999 (N_7999,N_7189,N_7390);
and U8000 (N_8000,N_7994,N_7986);
and U8001 (N_8001,N_7639,N_7656);
or U8002 (N_8002,N_7873,N_7874);
or U8003 (N_8003,N_7970,N_7562);
nor U8004 (N_8004,N_7515,N_7935);
or U8005 (N_8005,N_7502,N_7847);
nand U8006 (N_8006,N_7889,N_7551);
and U8007 (N_8007,N_7514,N_7649);
nand U8008 (N_8008,N_7575,N_7932);
nand U8009 (N_8009,N_7964,N_7794);
nand U8010 (N_8010,N_7771,N_7851);
and U8011 (N_8011,N_7927,N_7952);
or U8012 (N_8012,N_7734,N_7721);
nor U8013 (N_8013,N_7720,N_7988);
nor U8014 (N_8014,N_7733,N_7744);
nor U8015 (N_8015,N_7888,N_7629);
nand U8016 (N_8016,N_7563,N_7680);
and U8017 (N_8017,N_7858,N_7921);
or U8018 (N_8018,N_7728,N_7710);
nor U8019 (N_8019,N_7613,N_7813);
nor U8020 (N_8020,N_7907,N_7810);
nand U8021 (N_8021,N_7602,N_7600);
or U8022 (N_8022,N_7931,N_7506);
and U8023 (N_8023,N_7642,N_7749);
nor U8024 (N_8024,N_7962,N_7700);
nand U8025 (N_8025,N_7553,N_7542);
or U8026 (N_8026,N_7683,N_7902);
nor U8027 (N_8027,N_7606,N_7916);
or U8028 (N_8028,N_7691,N_7740);
xor U8029 (N_8029,N_7996,N_7567);
nand U8030 (N_8030,N_7912,N_7779);
or U8031 (N_8031,N_7516,N_7584);
and U8032 (N_8032,N_7971,N_7676);
nor U8033 (N_8033,N_7636,N_7992);
xor U8034 (N_8034,N_7974,N_7845);
nor U8035 (N_8035,N_7635,N_7622);
nand U8036 (N_8036,N_7752,N_7886);
nand U8037 (N_8037,N_7539,N_7903);
nor U8038 (N_8038,N_7648,N_7624);
or U8039 (N_8039,N_7596,N_7780);
nor U8040 (N_8040,N_7755,N_7781);
or U8041 (N_8041,N_7538,N_7709);
nand U8042 (N_8042,N_7601,N_7999);
and U8043 (N_8043,N_7520,N_7808);
xnor U8044 (N_8044,N_7532,N_7793);
or U8045 (N_8045,N_7603,N_7647);
or U8046 (N_8046,N_7876,N_7993);
nand U8047 (N_8047,N_7640,N_7938);
and U8048 (N_8048,N_7678,N_7564);
and U8049 (N_8049,N_7594,N_7791);
and U8050 (N_8050,N_7894,N_7669);
or U8051 (N_8051,N_7548,N_7834);
or U8052 (N_8052,N_7616,N_7763);
or U8053 (N_8053,N_7544,N_7821);
and U8054 (N_8054,N_7929,N_7574);
and U8055 (N_8055,N_7809,N_7995);
and U8056 (N_8056,N_7849,N_7658);
nor U8057 (N_8057,N_7754,N_7933);
xnor U8058 (N_8058,N_7922,N_7920);
and U8059 (N_8059,N_7893,N_7586);
xor U8060 (N_8060,N_7925,N_7628);
xor U8061 (N_8061,N_7765,N_7558);
and U8062 (N_8062,N_7766,N_7513);
or U8063 (N_8063,N_7688,N_7707);
nor U8064 (N_8064,N_7919,N_7812);
nand U8065 (N_8065,N_7891,N_7589);
xor U8066 (N_8066,N_7565,N_7623);
and U8067 (N_8067,N_7802,N_7725);
or U8068 (N_8068,N_7985,N_7905);
and U8069 (N_8069,N_7738,N_7896);
or U8070 (N_8070,N_7778,N_7850);
and U8071 (N_8071,N_7987,N_7819);
nand U8072 (N_8072,N_7915,N_7528);
nand U8073 (N_8073,N_7832,N_7543);
nor U8074 (N_8074,N_7698,N_7942);
or U8075 (N_8075,N_7652,N_7829);
or U8076 (N_8076,N_7972,N_7718);
and U8077 (N_8077,N_7941,N_7981);
nand U8078 (N_8078,N_7662,N_7879);
xnor U8079 (N_8079,N_7913,N_7897);
nor U8080 (N_8080,N_7536,N_7732);
nor U8081 (N_8081,N_7965,N_7863);
nand U8082 (N_8082,N_7541,N_7782);
nand U8083 (N_8083,N_7670,N_7830);
nand U8084 (N_8084,N_7762,N_7671);
and U8085 (N_8085,N_7654,N_7751);
and U8086 (N_8086,N_7880,N_7895);
and U8087 (N_8087,N_7547,N_7523);
xnor U8088 (N_8088,N_7769,N_7645);
nand U8089 (N_8089,N_7610,N_7742);
nand U8090 (N_8090,N_7522,N_7588);
nor U8091 (N_8091,N_7869,N_7590);
and U8092 (N_8092,N_7504,N_7665);
xnor U8093 (N_8093,N_7815,N_7825);
or U8094 (N_8094,N_7783,N_7572);
nand U8095 (N_8095,N_7776,N_7803);
nor U8096 (N_8096,N_7509,N_7862);
xnor U8097 (N_8097,N_7577,N_7911);
or U8098 (N_8098,N_7702,N_7521);
or U8099 (N_8099,N_7615,N_7978);
or U8100 (N_8100,N_7704,N_7500);
and U8101 (N_8101,N_7653,N_7634);
and U8102 (N_8102,N_7580,N_7861);
nor U8103 (N_8103,N_7945,N_7944);
and U8104 (N_8104,N_7597,N_7887);
nor U8105 (N_8105,N_7806,N_7787);
nand U8106 (N_8106,N_7626,N_7904);
or U8107 (N_8107,N_7956,N_7646);
or U8108 (N_8108,N_7609,N_7729);
nand U8109 (N_8109,N_7814,N_7570);
xnor U8110 (N_8110,N_7818,N_7883);
nor U8111 (N_8111,N_7591,N_7901);
nor U8112 (N_8112,N_7881,N_7675);
nor U8113 (N_8113,N_7790,N_7836);
nor U8114 (N_8114,N_7756,N_7655);
nand U8115 (N_8115,N_7966,N_7875);
nand U8116 (N_8116,N_7661,N_7840);
nor U8117 (N_8117,N_7923,N_7573);
nand U8118 (N_8118,N_7864,N_7918);
and U8119 (N_8119,N_7554,N_7726);
nand U8120 (N_8120,N_7585,N_7617);
nor U8121 (N_8121,N_7526,N_7795);
and U8122 (N_8122,N_7768,N_7770);
and U8123 (N_8123,N_7946,N_7885);
nand U8124 (N_8124,N_7550,N_7519);
nor U8125 (N_8125,N_7871,N_7736);
and U8126 (N_8126,N_7943,N_7898);
and U8127 (N_8127,N_7882,N_7837);
and U8128 (N_8128,N_7637,N_7761);
nor U8129 (N_8129,N_7699,N_7805);
and U8130 (N_8130,N_7578,N_7870);
nand U8131 (N_8131,N_7684,N_7960);
nand U8132 (N_8132,N_7817,N_7644);
nor U8133 (N_8133,N_7797,N_7682);
nor U8134 (N_8134,N_7576,N_7583);
xor U8135 (N_8135,N_7690,N_7745);
and U8136 (N_8136,N_7844,N_7841);
nor U8137 (N_8137,N_7846,N_7663);
nor U8138 (N_8138,N_7731,N_7786);
and U8139 (N_8139,N_7712,N_7664);
or U8140 (N_8140,N_7529,N_7743);
nand U8141 (N_8141,N_7711,N_7959);
nand U8142 (N_8142,N_7801,N_7552);
nand U8143 (N_8143,N_7884,N_7593);
xor U8144 (N_8144,N_7854,N_7505);
nand U8145 (N_8145,N_7827,N_7679);
nand U8146 (N_8146,N_7828,N_7632);
nand U8147 (N_8147,N_7820,N_7650);
nand U8148 (N_8148,N_7503,N_7757);
nand U8149 (N_8149,N_7612,N_7724);
nand U8150 (N_8150,N_7872,N_7822);
nand U8151 (N_8151,N_7982,N_7701);
or U8152 (N_8152,N_7799,N_7706);
xor U8153 (N_8153,N_7792,N_7848);
and U8154 (N_8154,N_7937,N_7659);
and U8155 (N_8155,N_7716,N_7674);
nand U8156 (N_8156,N_7967,N_7950);
nor U8157 (N_8157,N_7619,N_7697);
nor U8158 (N_8158,N_7865,N_7605);
nand U8159 (N_8159,N_7714,N_7686);
or U8160 (N_8160,N_7530,N_7677);
or U8161 (N_8161,N_7668,N_7512);
nor U8162 (N_8162,N_7607,N_7940);
or U8163 (N_8163,N_7730,N_7816);
and U8164 (N_8164,N_7977,N_7741);
or U8165 (N_8165,N_7804,N_7673);
nand U8166 (N_8166,N_7775,N_7651);
nand U8167 (N_8167,N_7777,N_7908);
nor U8168 (N_8168,N_7860,N_7560);
and U8169 (N_8169,N_7826,N_7511);
nor U8170 (N_8170,N_7934,N_7517);
or U8171 (N_8171,N_7693,N_7930);
and U8172 (N_8172,N_7900,N_7703);
and U8173 (N_8173,N_7501,N_7708);
nand U8174 (N_8174,N_7899,N_7980);
nor U8175 (N_8175,N_7638,N_7853);
nor U8176 (N_8176,N_7625,N_7961);
or U8177 (N_8177,N_7997,N_7975);
and U8178 (N_8178,N_7569,N_7559);
or U8179 (N_8179,N_7811,N_7525);
nor U8180 (N_8180,N_7568,N_7954);
nand U8181 (N_8181,N_7852,N_7892);
nand U8182 (N_8182,N_7633,N_7877);
or U8183 (N_8183,N_7592,N_7758);
and U8184 (N_8184,N_7890,N_7687);
nand U8185 (N_8185,N_7695,N_7753);
or U8186 (N_8186,N_7608,N_7604);
nor U8187 (N_8187,N_7939,N_7936);
nor U8188 (N_8188,N_7917,N_7722);
or U8189 (N_8189,N_7540,N_7856);
and U8190 (N_8190,N_7735,N_7681);
or U8191 (N_8191,N_7556,N_7969);
nor U8192 (N_8192,N_7507,N_7582);
nor U8193 (N_8193,N_7859,N_7527);
or U8194 (N_8194,N_7773,N_7842);
or U8195 (N_8195,N_7598,N_7785);
nand U8196 (N_8196,N_7914,N_7833);
or U8197 (N_8197,N_7566,N_7549);
nor U8198 (N_8198,N_7823,N_7947);
or U8199 (N_8199,N_7689,N_7831);
nor U8200 (N_8200,N_7747,N_7909);
xor U8201 (N_8201,N_7599,N_7581);
nand U8202 (N_8202,N_7705,N_7561);
and U8203 (N_8203,N_7926,N_7571);
and U8204 (N_8204,N_7928,N_7533);
nand U8205 (N_8205,N_7643,N_7534);
nor U8206 (N_8206,N_7685,N_7948);
nand U8207 (N_8207,N_7723,N_7746);
or U8208 (N_8208,N_7727,N_7667);
nor U8209 (N_8209,N_7984,N_7772);
or U8210 (N_8210,N_7717,N_7910);
nand U8211 (N_8211,N_7672,N_7990);
xor U8212 (N_8212,N_7949,N_7748);
xor U8213 (N_8213,N_7991,N_7621);
nand U8214 (N_8214,N_7979,N_7759);
and U8215 (N_8215,N_7555,N_7968);
or U8216 (N_8216,N_7508,N_7838);
or U8217 (N_8217,N_7694,N_7951);
nand U8218 (N_8218,N_7953,N_7535);
xnor U8219 (N_8219,N_7955,N_7867);
and U8220 (N_8220,N_7510,N_7537);
or U8221 (N_8221,N_7798,N_7627);
xor U8222 (N_8222,N_7579,N_7857);
nand U8223 (N_8223,N_7587,N_7767);
or U8224 (N_8224,N_7618,N_7878);
nand U8225 (N_8225,N_7713,N_7524);
nor U8226 (N_8226,N_7750,N_7692);
nor U8227 (N_8227,N_7518,N_7739);
and U8228 (N_8228,N_7839,N_7715);
and U8229 (N_8229,N_7719,N_7788);
or U8230 (N_8230,N_7546,N_7760);
and U8231 (N_8231,N_7835,N_7855);
or U8232 (N_8232,N_7631,N_7657);
and U8233 (N_8233,N_7963,N_7630);
xnor U8234 (N_8234,N_7824,N_7660);
nand U8235 (N_8235,N_7868,N_7800);
or U8236 (N_8236,N_7957,N_7998);
and U8237 (N_8237,N_7958,N_7924);
nand U8238 (N_8238,N_7620,N_7737);
or U8239 (N_8239,N_7789,N_7807);
nand U8240 (N_8240,N_7866,N_7774);
or U8241 (N_8241,N_7614,N_7983);
nor U8242 (N_8242,N_7989,N_7784);
nand U8243 (N_8243,N_7843,N_7976);
nor U8244 (N_8244,N_7696,N_7611);
or U8245 (N_8245,N_7973,N_7906);
nand U8246 (N_8246,N_7666,N_7545);
or U8247 (N_8247,N_7595,N_7641);
and U8248 (N_8248,N_7531,N_7557);
and U8249 (N_8249,N_7764,N_7796);
nand U8250 (N_8250,N_7956,N_7894);
xnor U8251 (N_8251,N_7932,N_7744);
nor U8252 (N_8252,N_7749,N_7713);
nand U8253 (N_8253,N_7544,N_7827);
nor U8254 (N_8254,N_7864,N_7949);
or U8255 (N_8255,N_7603,N_7879);
nor U8256 (N_8256,N_7708,N_7821);
nand U8257 (N_8257,N_7546,N_7920);
and U8258 (N_8258,N_7886,N_7978);
nand U8259 (N_8259,N_7722,N_7678);
or U8260 (N_8260,N_7965,N_7671);
nor U8261 (N_8261,N_7780,N_7524);
and U8262 (N_8262,N_7928,N_7905);
and U8263 (N_8263,N_7985,N_7895);
and U8264 (N_8264,N_7728,N_7616);
nand U8265 (N_8265,N_7807,N_7898);
nor U8266 (N_8266,N_7803,N_7804);
and U8267 (N_8267,N_7923,N_7971);
nand U8268 (N_8268,N_7697,N_7896);
xor U8269 (N_8269,N_7619,N_7758);
and U8270 (N_8270,N_7516,N_7718);
nand U8271 (N_8271,N_7838,N_7959);
and U8272 (N_8272,N_7961,N_7631);
nor U8273 (N_8273,N_7833,N_7987);
or U8274 (N_8274,N_7998,N_7902);
xor U8275 (N_8275,N_7504,N_7734);
and U8276 (N_8276,N_7801,N_7555);
nor U8277 (N_8277,N_7570,N_7539);
nand U8278 (N_8278,N_7545,N_7714);
and U8279 (N_8279,N_7742,N_7752);
or U8280 (N_8280,N_7677,N_7821);
or U8281 (N_8281,N_7970,N_7538);
nor U8282 (N_8282,N_7878,N_7868);
nor U8283 (N_8283,N_7991,N_7539);
nand U8284 (N_8284,N_7775,N_7666);
xnor U8285 (N_8285,N_7920,N_7625);
or U8286 (N_8286,N_7883,N_7639);
nor U8287 (N_8287,N_7710,N_7721);
or U8288 (N_8288,N_7922,N_7503);
or U8289 (N_8289,N_7647,N_7652);
and U8290 (N_8290,N_7749,N_7547);
or U8291 (N_8291,N_7784,N_7985);
nand U8292 (N_8292,N_7592,N_7547);
or U8293 (N_8293,N_7851,N_7917);
xor U8294 (N_8294,N_7547,N_7520);
nand U8295 (N_8295,N_7639,N_7716);
xor U8296 (N_8296,N_7835,N_7876);
xnor U8297 (N_8297,N_7975,N_7961);
and U8298 (N_8298,N_7783,N_7698);
or U8299 (N_8299,N_7637,N_7915);
and U8300 (N_8300,N_7600,N_7903);
xor U8301 (N_8301,N_7655,N_7711);
nand U8302 (N_8302,N_7636,N_7766);
nor U8303 (N_8303,N_7582,N_7785);
xnor U8304 (N_8304,N_7988,N_7770);
or U8305 (N_8305,N_7565,N_7838);
or U8306 (N_8306,N_7877,N_7651);
xnor U8307 (N_8307,N_7948,N_7564);
and U8308 (N_8308,N_7966,N_7954);
and U8309 (N_8309,N_7729,N_7834);
and U8310 (N_8310,N_7721,N_7665);
nor U8311 (N_8311,N_7527,N_7999);
xor U8312 (N_8312,N_7804,N_7596);
nand U8313 (N_8313,N_7548,N_7597);
and U8314 (N_8314,N_7562,N_7501);
xor U8315 (N_8315,N_7561,N_7922);
nand U8316 (N_8316,N_7595,N_7876);
nand U8317 (N_8317,N_7602,N_7808);
or U8318 (N_8318,N_7949,N_7845);
or U8319 (N_8319,N_7721,N_7521);
xnor U8320 (N_8320,N_7973,N_7725);
nor U8321 (N_8321,N_7984,N_7600);
and U8322 (N_8322,N_7513,N_7733);
nor U8323 (N_8323,N_7968,N_7891);
nor U8324 (N_8324,N_7533,N_7513);
or U8325 (N_8325,N_7586,N_7684);
or U8326 (N_8326,N_7569,N_7991);
nor U8327 (N_8327,N_7744,N_7568);
xnor U8328 (N_8328,N_7597,N_7595);
or U8329 (N_8329,N_7934,N_7738);
nand U8330 (N_8330,N_7698,N_7869);
and U8331 (N_8331,N_7536,N_7540);
or U8332 (N_8332,N_7920,N_7693);
or U8333 (N_8333,N_7965,N_7822);
nand U8334 (N_8334,N_7574,N_7946);
xor U8335 (N_8335,N_7673,N_7741);
nor U8336 (N_8336,N_7701,N_7606);
xnor U8337 (N_8337,N_7927,N_7968);
nand U8338 (N_8338,N_7600,N_7762);
and U8339 (N_8339,N_7949,N_7540);
and U8340 (N_8340,N_7510,N_7769);
and U8341 (N_8341,N_7961,N_7667);
and U8342 (N_8342,N_7695,N_7869);
nor U8343 (N_8343,N_7813,N_7632);
or U8344 (N_8344,N_7728,N_7767);
or U8345 (N_8345,N_7740,N_7778);
nand U8346 (N_8346,N_7669,N_7504);
nand U8347 (N_8347,N_7766,N_7891);
nand U8348 (N_8348,N_7823,N_7708);
and U8349 (N_8349,N_7955,N_7856);
xor U8350 (N_8350,N_7901,N_7863);
nand U8351 (N_8351,N_7815,N_7751);
or U8352 (N_8352,N_7631,N_7682);
nand U8353 (N_8353,N_7807,N_7870);
and U8354 (N_8354,N_7949,N_7896);
nor U8355 (N_8355,N_7573,N_7862);
nand U8356 (N_8356,N_7672,N_7634);
nand U8357 (N_8357,N_7938,N_7632);
nand U8358 (N_8358,N_7830,N_7815);
or U8359 (N_8359,N_7644,N_7639);
and U8360 (N_8360,N_7819,N_7887);
nand U8361 (N_8361,N_7944,N_7954);
or U8362 (N_8362,N_7629,N_7667);
or U8363 (N_8363,N_7721,N_7849);
xor U8364 (N_8364,N_7984,N_7927);
nor U8365 (N_8365,N_7891,N_7952);
or U8366 (N_8366,N_7838,N_7786);
nand U8367 (N_8367,N_7936,N_7970);
and U8368 (N_8368,N_7967,N_7589);
nand U8369 (N_8369,N_7712,N_7950);
xnor U8370 (N_8370,N_7534,N_7829);
nand U8371 (N_8371,N_7773,N_7806);
and U8372 (N_8372,N_7502,N_7588);
nand U8373 (N_8373,N_7517,N_7850);
or U8374 (N_8374,N_7889,N_7721);
or U8375 (N_8375,N_7841,N_7759);
and U8376 (N_8376,N_7630,N_7937);
and U8377 (N_8377,N_7819,N_7685);
nand U8378 (N_8378,N_7641,N_7707);
nor U8379 (N_8379,N_7641,N_7874);
nor U8380 (N_8380,N_7712,N_7922);
nor U8381 (N_8381,N_7684,N_7562);
xor U8382 (N_8382,N_7513,N_7788);
and U8383 (N_8383,N_7819,N_7521);
and U8384 (N_8384,N_7571,N_7881);
and U8385 (N_8385,N_7683,N_7901);
nand U8386 (N_8386,N_7637,N_7853);
and U8387 (N_8387,N_7855,N_7653);
nand U8388 (N_8388,N_7861,N_7734);
nand U8389 (N_8389,N_7738,N_7736);
nand U8390 (N_8390,N_7896,N_7779);
and U8391 (N_8391,N_7630,N_7964);
nor U8392 (N_8392,N_7664,N_7505);
or U8393 (N_8393,N_7662,N_7925);
or U8394 (N_8394,N_7796,N_7686);
nand U8395 (N_8395,N_7891,N_7759);
nor U8396 (N_8396,N_7593,N_7962);
nor U8397 (N_8397,N_7903,N_7570);
nor U8398 (N_8398,N_7756,N_7638);
nor U8399 (N_8399,N_7955,N_7673);
and U8400 (N_8400,N_7846,N_7682);
nor U8401 (N_8401,N_7840,N_7781);
nand U8402 (N_8402,N_7948,N_7758);
nand U8403 (N_8403,N_7984,N_7855);
nor U8404 (N_8404,N_7837,N_7900);
nor U8405 (N_8405,N_7510,N_7970);
nor U8406 (N_8406,N_7991,N_7981);
and U8407 (N_8407,N_7920,N_7527);
or U8408 (N_8408,N_7809,N_7657);
or U8409 (N_8409,N_7776,N_7663);
xor U8410 (N_8410,N_7993,N_7853);
and U8411 (N_8411,N_7698,N_7638);
nand U8412 (N_8412,N_7853,N_7963);
and U8413 (N_8413,N_7702,N_7546);
and U8414 (N_8414,N_7830,N_7916);
nor U8415 (N_8415,N_7843,N_7556);
nand U8416 (N_8416,N_7697,N_7635);
or U8417 (N_8417,N_7574,N_7956);
and U8418 (N_8418,N_7743,N_7606);
nand U8419 (N_8419,N_7606,N_7737);
xnor U8420 (N_8420,N_7838,N_7800);
and U8421 (N_8421,N_7639,N_7881);
and U8422 (N_8422,N_7872,N_7944);
nor U8423 (N_8423,N_7813,N_7673);
xnor U8424 (N_8424,N_7779,N_7721);
nor U8425 (N_8425,N_7991,N_7743);
nand U8426 (N_8426,N_7881,N_7744);
and U8427 (N_8427,N_7635,N_7886);
xnor U8428 (N_8428,N_7652,N_7910);
nand U8429 (N_8429,N_7670,N_7937);
nand U8430 (N_8430,N_7951,N_7860);
nand U8431 (N_8431,N_7530,N_7935);
or U8432 (N_8432,N_7564,N_7877);
nor U8433 (N_8433,N_7548,N_7974);
or U8434 (N_8434,N_7821,N_7882);
or U8435 (N_8435,N_7863,N_7510);
xnor U8436 (N_8436,N_7628,N_7746);
nor U8437 (N_8437,N_7566,N_7944);
or U8438 (N_8438,N_7576,N_7998);
nor U8439 (N_8439,N_7877,N_7568);
nand U8440 (N_8440,N_7796,N_7769);
or U8441 (N_8441,N_7935,N_7786);
nand U8442 (N_8442,N_7558,N_7700);
nand U8443 (N_8443,N_7995,N_7562);
nor U8444 (N_8444,N_7770,N_7827);
xnor U8445 (N_8445,N_7860,N_7845);
nor U8446 (N_8446,N_7833,N_7529);
or U8447 (N_8447,N_7536,N_7645);
xnor U8448 (N_8448,N_7550,N_7879);
nor U8449 (N_8449,N_7729,N_7524);
nor U8450 (N_8450,N_7834,N_7762);
nor U8451 (N_8451,N_7637,N_7919);
and U8452 (N_8452,N_7772,N_7535);
nand U8453 (N_8453,N_7595,N_7713);
nor U8454 (N_8454,N_7705,N_7944);
or U8455 (N_8455,N_7974,N_7704);
nand U8456 (N_8456,N_7520,N_7657);
nor U8457 (N_8457,N_7752,N_7583);
nor U8458 (N_8458,N_7974,N_7601);
xor U8459 (N_8459,N_7876,N_7501);
nand U8460 (N_8460,N_7829,N_7564);
xnor U8461 (N_8461,N_7612,N_7864);
or U8462 (N_8462,N_7953,N_7935);
nand U8463 (N_8463,N_7805,N_7638);
nand U8464 (N_8464,N_7947,N_7745);
nand U8465 (N_8465,N_7938,N_7741);
xor U8466 (N_8466,N_7716,N_7798);
nor U8467 (N_8467,N_7696,N_7910);
and U8468 (N_8468,N_7748,N_7581);
and U8469 (N_8469,N_7717,N_7698);
xnor U8470 (N_8470,N_7806,N_7728);
nand U8471 (N_8471,N_7852,N_7606);
or U8472 (N_8472,N_7913,N_7584);
and U8473 (N_8473,N_7502,N_7748);
or U8474 (N_8474,N_7652,N_7786);
and U8475 (N_8475,N_7977,N_7982);
and U8476 (N_8476,N_7761,N_7629);
or U8477 (N_8477,N_7587,N_7690);
nand U8478 (N_8478,N_7557,N_7971);
nor U8479 (N_8479,N_7990,N_7952);
nand U8480 (N_8480,N_7938,N_7847);
and U8481 (N_8481,N_7913,N_7861);
nor U8482 (N_8482,N_7765,N_7791);
nand U8483 (N_8483,N_7925,N_7547);
and U8484 (N_8484,N_7521,N_7511);
nand U8485 (N_8485,N_7674,N_7597);
nand U8486 (N_8486,N_7640,N_7555);
or U8487 (N_8487,N_7982,N_7878);
and U8488 (N_8488,N_7871,N_7763);
or U8489 (N_8489,N_7815,N_7534);
nand U8490 (N_8490,N_7618,N_7715);
nor U8491 (N_8491,N_7656,N_7795);
or U8492 (N_8492,N_7691,N_7690);
nand U8493 (N_8493,N_7831,N_7774);
xnor U8494 (N_8494,N_7776,N_7652);
nand U8495 (N_8495,N_7732,N_7982);
nand U8496 (N_8496,N_7537,N_7944);
nand U8497 (N_8497,N_7893,N_7997);
nand U8498 (N_8498,N_7818,N_7716);
nor U8499 (N_8499,N_7746,N_7511);
and U8500 (N_8500,N_8213,N_8413);
and U8501 (N_8501,N_8072,N_8462);
nand U8502 (N_8502,N_8007,N_8266);
or U8503 (N_8503,N_8202,N_8187);
nor U8504 (N_8504,N_8281,N_8456);
nand U8505 (N_8505,N_8130,N_8285);
nand U8506 (N_8506,N_8359,N_8217);
nor U8507 (N_8507,N_8200,N_8077);
xor U8508 (N_8508,N_8050,N_8319);
and U8509 (N_8509,N_8051,N_8028);
nand U8510 (N_8510,N_8149,N_8396);
or U8511 (N_8511,N_8435,N_8243);
xnor U8512 (N_8512,N_8086,N_8001);
and U8513 (N_8513,N_8487,N_8417);
nor U8514 (N_8514,N_8412,N_8401);
xor U8515 (N_8515,N_8238,N_8268);
and U8516 (N_8516,N_8191,N_8037);
nand U8517 (N_8517,N_8152,N_8458);
and U8518 (N_8518,N_8492,N_8208);
xnor U8519 (N_8519,N_8354,N_8450);
xnor U8520 (N_8520,N_8375,N_8157);
nand U8521 (N_8521,N_8372,N_8170);
nor U8522 (N_8522,N_8443,N_8475);
or U8523 (N_8523,N_8025,N_8033);
nand U8524 (N_8524,N_8128,N_8315);
nand U8525 (N_8525,N_8175,N_8111);
nor U8526 (N_8526,N_8383,N_8089);
nand U8527 (N_8527,N_8437,N_8044);
nand U8528 (N_8528,N_8054,N_8369);
and U8529 (N_8529,N_8222,N_8153);
nor U8530 (N_8530,N_8184,N_8063);
nor U8531 (N_8531,N_8296,N_8498);
nor U8532 (N_8532,N_8232,N_8134);
nand U8533 (N_8533,N_8465,N_8382);
nor U8534 (N_8534,N_8259,N_8103);
nor U8535 (N_8535,N_8303,N_8236);
nor U8536 (N_8536,N_8003,N_8047);
nand U8537 (N_8537,N_8404,N_8022);
and U8538 (N_8538,N_8101,N_8166);
or U8539 (N_8539,N_8224,N_8280);
nand U8540 (N_8540,N_8029,N_8004);
nand U8541 (N_8541,N_8373,N_8317);
xor U8542 (N_8542,N_8242,N_8485);
and U8543 (N_8543,N_8334,N_8239);
nor U8544 (N_8544,N_8035,N_8364);
or U8545 (N_8545,N_8381,N_8488);
nand U8546 (N_8546,N_8362,N_8415);
and U8547 (N_8547,N_8418,N_8489);
or U8548 (N_8548,N_8341,N_8034);
or U8549 (N_8549,N_8366,N_8091);
or U8550 (N_8550,N_8146,N_8444);
nand U8551 (N_8551,N_8172,N_8246);
and U8552 (N_8552,N_8350,N_8019);
or U8553 (N_8553,N_8347,N_8137);
nor U8554 (N_8554,N_8141,N_8289);
xor U8555 (N_8555,N_8446,N_8041);
nand U8556 (N_8556,N_8258,N_8231);
nor U8557 (N_8557,N_8247,N_8066);
nand U8558 (N_8558,N_8169,N_8371);
xor U8559 (N_8559,N_8235,N_8457);
or U8560 (N_8560,N_8297,N_8438);
nor U8561 (N_8561,N_8422,N_8240);
nand U8562 (N_8562,N_8429,N_8336);
nand U8563 (N_8563,N_8244,N_8448);
nor U8564 (N_8564,N_8271,N_8349);
nor U8565 (N_8565,N_8279,N_8305);
and U8566 (N_8566,N_8110,N_8274);
nor U8567 (N_8567,N_8299,N_8138);
and U8568 (N_8568,N_8181,N_8178);
or U8569 (N_8569,N_8070,N_8132);
nor U8570 (N_8570,N_8008,N_8218);
nand U8571 (N_8571,N_8339,N_8405);
nor U8572 (N_8572,N_8333,N_8447);
or U8573 (N_8573,N_8201,N_8384);
nor U8574 (N_8574,N_8049,N_8420);
nand U8575 (N_8575,N_8156,N_8433);
nand U8576 (N_8576,N_8131,N_8300);
or U8577 (N_8577,N_8451,N_8469);
and U8578 (N_8578,N_8223,N_8030);
or U8579 (N_8579,N_8490,N_8264);
nand U8580 (N_8580,N_8343,N_8379);
and U8581 (N_8581,N_8411,N_8024);
nor U8582 (N_8582,N_8278,N_8093);
and U8583 (N_8583,N_8416,N_8251);
or U8584 (N_8584,N_8291,N_8171);
and U8585 (N_8585,N_8430,N_8073);
xor U8586 (N_8586,N_8257,N_8102);
nor U8587 (N_8587,N_8174,N_8160);
and U8588 (N_8588,N_8021,N_8309);
nand U8589 (N_8589,N_8229,N_8112);
xor U8590 (N_8590,N_8183,N_8253);
or U8591 (N_8591,N_8467,N_8431);
nand U8592 (N_8592,N_8476,N_8150);
xor U8593 (N_8593,N_8064,N_8026);
and U8594 (N_8594,N_8220,N_8290);
nor U8595 (N_8595,N_8387,N_8454);
nand U8596 (N_8596,N_8075,N_8313);
or U8597 (N_8597,N_8393,N_8331);
or U8598 (N_8598,N_8298,N_8212);
and U8599 (N_8599,N_8227,N_8079);
or U8600 (N_8600,N_8085,N_8464);
xor U8601 (N_8601,N_8479,N_8321);
nand U8602 (N_8602,N_8302,N_8282);
and U8603 (N_8603,N_8460,N_8482);
nand U8604 (N_8604,N_8159,N_8392);
or U8605 (N_8605,N_8256,N_8306);
and U8606 (N_8606,N_8409,N_8012);
and U8607 (N_8607,N_8328,N_8228);
or U8608 (N_8608,N_8318,N_8142);
nor U8609 (N_8609,N_8121,N_8173);
nor U8610 (N_8610,N_8324,N_8310);
nand U8611 (N_8611,N_8252,N_8267);
nor U8612 (N_8612,N_8126,N_8378);
xor U8613 (N_8613,N_8164,N_8006);
nor U8614 (N_8614,N_8403,N_8076);
nand U8615 (N_8615,N_8081,N_8145);
nand U8616 (N_8616,N_8090,N_8052);
nor U8617 (N_8617,N_8261,N_8494);
and U8618 (N_8618,N_8391,N_8071);
or U8619 (N_8619,N_8365,N_8196);
and U8620 (N_8620,N_8214,N_8406);
nand U8621 (N_8621,N_8165,N_8046);
xor U8622 (N_8622,N_8162,N_8277);
nand U8623 (N_8623,N_8136,N_8345);
xnor U8624 (N_8624,N_8135,N_8140);
or U8625 (N_8625,N_8179,N_8120);
or U8626 (N_8626,N_8427,N_8316);
nand U8627 (N_8627,N_8002,N_8441);
and U8628 (N_8628,N_8186,N_8499);
xor U8629 (N_8629,N_8481,N_8432);
and U8630 (N_8630,N_8275,N_8468);
and U8631 (N_8631,N_8395,N_8105);
nand U8632 (N_8632,N_8107,N_8419);
nand U8633 (N_8633,N_8389,N_8158);
nor U8634 (N_8634,N_8342,N_8118);
nand U8635 (N_8635,N_8211,N_8470);
nor U8636 (N_8636,N_8304,N_8486);
nand U8637 (N_8637,N_8058,N_8491);
or U8638 (N_8638,N_8016,N_8466);
and U8639 (N_8639,N_8320,N_8209);
xnor U8640 (N_8640,N_8151,N_8356);
and U8641 (N_8641,N_8119,N_8276);
or U8642 (N_8642,N_8097,N_8043);
nor U8643 (N_8643,N_8327,N_8376);
and U8644 (N_8644,N_8332,N_8445);
nor U8645 (N_8645,N_8286,N_8358);
and U8646 (N_8646,N_8036,N_8326);
nor U8647 (N_8647,N_8067,N_8199);
nor U8648 (N_8648,N_8361,N_8380);
nor U8649 (N_8649,N_8233,N_8061);
or U8650 (N_8650,N_8100,N_8497);
or U8651 (N_8651,N_8283,N_8250);
nand U8652 (N_8652,N_8189,N_8322);
or U8653 (N_8653,N_8000,N_8292);
nor U8654 (N_8654,N_8254,N_8068);
and U8655 (N_8655,N_8032,N_8198);
nand U8656 (N_8656,N_8014,N_8386);
nor U8657 (N_8657,N_8206,N_8125);
nor U8658 (N_8658,N_8203,N_8057);
nand U8659 (N_8659,N_8474,N_8426);
or U8660 (N_8660,N_8461,N_8069);
xor U8661 (N_8661,N_8225,N_8344);
xor U8662 (N_8662,N_8330,N_8098);
nand U8663 (N_8663,N_8104,N_8230);
or U8664 (N_8664,N_8095,N_8010);
nor U8665 (N_8665,N_8018,N_8295);
xor U8666 (N_8666,N_8452,N_8092);
nand U8667 (N_8667,N_8477,N_8493);
xor U8668 (N_8668,N_8219,N_8205);
or U8669 (N_8669,N_8117,N_8195);
or U8670 (N_8670,N_8423,N_8325);
nor U8671 (N_8671,N_8323,N_8115);
or U8672 (N_8672,N_8301,N_8442);
nand U8673 (N_8673,N_8062,N_8352);
or U8674 (N_8674,N_8221,N_8122);
and U8675 (N_8675,N_8059,N_8048);
or U8676 (N_8676,N_8155,N_8367);
and U8677 (N_8677,N_8394,N_8484);
or U8678 (N_8678,N_8353,N_8408);
and U8679 (N_8679,N_8038,N_8216);
nand U8680 (N_8680,N_8397,N_8180);
nor U8681 (N_8681,N_8124,N_8197);
or U8682 (N_8682,N_8357,N_8449);
nor U8683 (N_8683,N_8255,N_8428);
or U8684 (N_8684,N_8414,N_8440);
nand U8685 (N_8685,N_8154,N_8288);
nor U8686 (N_8686,N_8472,N_8060);
nand U8687 (N_8687,N_8087,N_8190);
and U8688 (N_8688,N_8215,N_8177);
nor U8689 (N_8689,N_8390,N_8065);
nor U8690 (N_8690,N_8015,N_8193);
nor U8691 (N_8691,N_8312,N_8346);
nand U8692 (N_8692,N_8096,N_8351);
nand U8693 (N_8693,N_8053,N_8192);
and U8694 (N_8694,N_8400,N_8455);
nor U8695 (N_8695,N_8385,N_8168);
and U8696 (N_8696,N_8039,N_8473);
or U8697 (N_8697,N_8148,N_8308);
or U8698 (N_8698,N_8338,N_8082);
nand U8699 (N_8699,N_8377,N_8495);
nand U8700 (N_8700,N_8471,N_8139);
nor U8701 (N_8701,N_8410,N_8020);
and U8702 (N_8702,N_8088,N_8094);
nor U8703 (N_8703,N_8270,N_8311);
nand U8704 (N_8704,N_8335,N_8355);
nand U8705 (N_8705,N_8055,N_8116);
or U8706 (N_8706,N_8241,N_8388);
or U8707 (N_8707,N_8269,N_8307);
nand U8708 (N_8708,N_8478,N_8237);
or U8709 (N_8709,N_8084,N_8496);
nand U8710 (N_8710,N_8340,N_8127);
and U8711 (N_8711,N_8374,N_8109);
nor U8712 (N_8712,N_8287,N_8245);
nor U8713 (N_8713,N_8045,N_8176);
and U8714 (N_8714,N_8398,N_8161);
nand U8715 (N_8715,N_8078,N_8234);
nand U8716 (N_8716,N_8249,N_8133);
nand U8717 (N_8717,N_8348,N_8263);
nor U8718 (N_8718,N_8248,N_8011);
or U8719 (N_8719,N_8106,N_8027);
xor U8720 (N_8720,N_8017,N_8260);
and U8721 (N_8721,N_8273,N_8337);
and U8722 (N_8722,N_8009,N_8013);
nor U8723 (N_8723,N_8483,N_8363);
nand U8724 (N_8724,N_8329,N_8163);
and U8725 (N_8725,N_8129,N_8421);
nand U8726 (N_8726,N_8042,N_8123);
or U8727 (N_8727,N_8144,N_8294);
nand U8728 (N_8728,N_8143,N_8424);
nor U8729 (N_8729,N_8083,N_8182);
nor U8730 (N_8730,N_8188,N_8099);
and U8731 (N_8731,N_8425,N_8114);
nor U8732 (N_8732,N_8207,N_8204);
nand U8733 (N_8733,N_8399,N_8113);
nor U8734 (N_8734,N_8368,N_8265);
nor U8735 (N_8735,N_8262,N_8272);
nand U8736 (N_8736,N_8108,N_8459);
xnor U8737 (N_8737,N_8210,N_8436);
nand U8738 (N_8738,N_8185,N_8434);
nand U8739 (N_8739,N_8453,N_8463);
nor U8740 (N_8740,N_8040,N_8005);
and U8741 (N_8741,N_8480,N_8194);
or U8742 (N_8742,N_8056,N_8293);
xnor U8743 (N_8743,N_8370,N_8407);
or U8744 (N_8744,N_8226,N_8167);
and U8745 (N_8745,N_8031,N_8080);
or U8746 (N_8746,N_8360,N_8147);
or U8747 (N_8747,N_8439,N_8314);
nand U8748 (N_8748,N_8402,N_8284);
nand U8749 (N_8749,N_8023,N_8074);
nor U8750 (N_8750,N_8402,N_8060);
or U8751 (N_8751,N_8353,N_8210);
xor U8752 (N_8752,N_8488,N_8103);
nor U8753 (N_8753,N_8027,N_8001);
nor U8754 (N_8754,N_8349,N_8129);
nor U8755 (N_8755,N_8490,N_8355);
nand U8756 (N_8756,N_8214,N_8235);
nor U8757 (N_8757,N_8249,N_8090);
nand U8758 (N_8758,N_8273,N_8137);
nor U8759 (N_8759,N_8410,N_8292);
or U8760 (N_8760,N_8100,N_8287);
nand U8761 (N_8761,N_8368,N_8141);
nor U8762 (N_8762,N_8415,N_8490);
nor U8763 (N_8763,N_8028,N_8036);
or U8764 (N_8764,N_8134,N_8218);
nor U8765 (N_8765,N_8026,N_8415);
nor U8766 (N_8766,N_8439,N_8436);
nor U8767 (N_8767,N_8330,N_8453);
and U8768 (N_8768,N_8322,N_8245);
or U8769 (N_8769,N_8125,N_8242);
nand U8770 (N_8770,N_8008,N_8448);
or U8771 (N_8771,N_8323,N_8081);
and U8772 (N_8772,N_8499,N_8047);
or U8773 (N_8773,N_8365,N_8465);
nor U8774 (N_8774,N_8399,N_8171);
nor U8775 (N_8775,N_8388,N_8358);
or U8776 (N_8776,N_8141,N_8257);
xor U8777 (N_8777,N_8096,N_8287);
or U8778 (N_8778,N_8225,N_8496);
nand U8779 (N_8779,N_8163,N_8174);
nand U8780 (N_8780,N_8393,N_8228);
or U8781 (N_8781,N_8311,N_8015);
and U8782 (N_8782,N_8309,N_8038);
or U8783 (N_8783,N_8089,N_8200);
nand U8784 (N_8784,N_8441,N_8058);
or U8785 (N_8785,N_8476,N_8134);
nand U8786 (N_8786,N_8476,N_8211);
nand U8787 (N_8787,N_8289,N_8319);
and U8788 (N_8788,N_8433,N_8179);
and U8789 (N_8789,N_8475,N_8066);
and U8790 (N_8790,N_8074,N_8392);
nand U8791 (N_8791,N_8160,N_8311);
or U8792 (N_8792,N_8222,N_8486);
nand U8793 (N_8793,N_8157,N_8303);
nor U8794 (N_8794,N_8179,N_8223);
nand U8795 (N_8795,N_8339,N_8242);
or U8796 (N_8796,N_8109,N_8200);
or U8797 (N_8797,N_8455,N_8350);
and U8798 (N_8798,N_8252,N_8239);
xor U8799 (N_8799,N_8029,N_8118);
nor U8800 (N_8800,N_8262,N_8482);
xnor U8801 (N_8801,N_8145,N_8489);
nor U8802 (N_8802,N_8260,N_8423);
and U8803 (N_8803,N_8152,N_8314);
nor U8804 (N_8804,N_8127,N_8273);
or U8805 (N_8805,N_8323,N_8238);
or U8806 (N_8806,N_8411,N_8129);
nor U8807 (N_8807,N_8141,N_8251);
nand U8808 (N_8808,N_8101,N_8232);
and U8809 (N_8809,N_8301,N_8499);
nand U8810 (N_8810,N_8343,N_8154);
or U8811 (N_8811,N_8498,N_8427);
nor U8812 (N_8812,N_8157,N_8158);
or U8813 (N_8813,N_8057,N_8286);
nor U8814 (N_8814,N_8160,N_8080);
and U8815 (N_8815,N_8164,N_8270);
nand U8816 (N_8816,N_8075,N_8479);
nor U8817 (N_8817,N_8154,N_8080);
or U8818 (N_8818,N_8264,N_8323);
nor U8819 (N_8819,N_8132,N_8281);
and U8820 (N_8820,N_8211,N_8374);
nor U8821 (N_8821,N_8201,N_8013);
or U8822 (N_8822,N_8372,N_8289);
or U8823 (N_8823,N_8418,N_8414);
and U8824 (N_8824,N_8480,N_8182);
and U8825 (N_8825,N_8458,N_8100);
nor U8826 (N_8826,N_8476,N_8457);
or U8827 (N_8827,N_8076,N_8382);
or U8828 (N_8828,N_8160,N_8222);
or U8829 (N_8829,N_8101,N_8416);
nand U8830 (N_8830,N_8026,N_8079);
nor U8831 (N_8831,N_8289,N_8373);
or U8832 (N_8832,N_8221,N_8184);
or U8833 (N_8833,N_8210,N_8181);
and U8834 (N_8834,N_8214,N_8022);
nor U8835 (N_8835,N_8333,N_8232);
and U8836 (N_8836,N_8450,N_8064);
or U8837 (N_8837,N_8067,N_8002);
or U8838 (N_8838,N_8061,N_8119);
xnor U8839 (N_8839,N_8232,N_8156);
and U8840 (N_8840,N_8262,N_8389);
or U8841 (N_8841,N_8480,N_8018);
or U8842 (N_8842,N_8325,N_8322);
nor U8843 (N_8843,N_8083,N_8101);
and U8844 (N_8844,N_8014,N_8225);
nand U8845 (N_8845,N_8239,N_8261);
nand U8846 (N_8846,N_8067,N_8423);
xnor U8847 (N_8847,N_8281,N_8328);
nor U8848 (N_8848,N_8317,N_8405);
nand U8849 (N_8849,N_8216,N_8360);
and U8850 (N_8850,N_8209,N_8256);
nor U8851 (N_8851,N_8129,N_8146);
nand U8852 (N_8852,N_8386,N_8476);
or U8853 (N_8853,N_8394,N_8423);
nand U8854 (N_8854,N_8161,N_8099);
and U8855 (N_8855,N_8162,N_8226);
nor U8856 (N_8856,N_8317,N_8350);
xor U8857 (N_8857,N_8162,N_8203);
or U8858 (N_8858,N_8390,N_8384);
and U8859 (N_8859,N_8013,N_8422);
nand U8860 (N_8860,N_8162,N_8329);
nand U8861 (N_8861,N_8493,N_8129);
nor U8862 (N_8862,N_8482,N_8058);
and U8863 (N_8863,N_8063,N_8415);
and U8864 (N_8864,N_8294,N_8050);
or U8865 (N_8865,N_8397,N_8156);
nand U8866 (N_8866,N_8076,N_8270);
or U8867 (N_8867,N_8450,N_8499);
and U8868 (N_8868,N_8306,N_8359);
and U8869 (N_8869,N_8418,N_8460);
and U8870 (N_8870,N_8205,N_8143);
and U8871 (N_8871,N_8153,N_8445);
nor U8872 (N_8872,N_8286,N_8039);
nand U8873 (N_8873,N_8206,N_8436);
nand U8874 (N_8874,N_8120,N_8454);
nand U8875 (N_8875,N_8102,N_8042);
nand U8876 (N_8876,N_8415,N_8496);
or U8877 (N_8877,N_8156,N_8162);
nand U8878 (N_8878,N_8200,N_8481);
xor U8879 (N_8879,N_8062,N_8042);
or U8880 (N_8880,N_8428,N_8026);
nor U8881 (N_8881,N_8311,N_8221);
or U8882 (N_8882,N_8174,N_8486);
or U8883 (N_8883,N_8252,N_8345);
and U8884 (N_8884,N_8140,N_8139);
or U8885 (N_8885,N_8421,N_8105);
nor U8886 (N_8886,N_8422,N_8304);
and U8887 (N_8887,N_8311,N_8182);
and U8888 (N_8888,N_8361,N_8252);
xor U8889 (N_8889,N_8305,N_8361);
and U8890 (N_8890,N_8232,N_8256);
or U8891 (N_8891,N_8000,N_8330);
nand U8892 (N_8892,N_8340,N_8215);
or U8893 (N_8893,N_8273,N_8209);
nor U8894 (N_8894,N_8450,N_8284);
or U8895 (N_8895,N_8333,N_8024);
or U8896 (N_8896,N_8406,N_8371);
nand U8897 (N_8897,N_8484,N_8204);
nor U8898 (N_8898,N_8459,N_8389);
and U8899 (N_8899,N_8263,N_8022);
xor U8900 (N_8900,N_8099,N_8088);
and U8901 (N_8901,N_8274,N_8138);
nand U8902 (N_8902,N_8352,N_8003);
and U8903 (N_8903,N_8059,N_8345);
nor U8904 (N_8904,N_8444,N_8065);
xor U8905 (N_8905,N_8053,N_8393);
or U8906 (N_8906,N_8170,N_8214);
nand U8907 (N_8907,N_8286,N_8494);
nand U8908 (N_8908,N_8270,N_8033);
nor U8909 (N_8909,N_8376,N_8449);
nor U8910 (N_8910,N_8218,N_8143);
or U8911 (N_8911,N_8313,N_8484);
nand U8912 (N_8912,N_8136,N_8054);
and U8913 (N_8913,N_8179,N_8157);
and U8914 (N_8914,N_8089,N_8228);
nor U8915 (N_8915,N_8343,N_8395);
and U8916 (N_8916,N_8432,N_8115);
and U8917 (N_8917,N_8156,N_8353);
xor U8918 (N_8918,N_8138,N_8108);
nor U8919 (N_8919,N_8322,N_8108);
or U8920 (N_8920,N_8120,N_8447);
and U8921 (N_8921,N_8100,N_8129);
nand U8922 (N_8922,N_8389,N_8041);
and U8923 (N_8923,N_8030,N_8156);
nor U8924 (N_8924,N_8498,N_8060);
or U8925 (N_8925,N_8032,N_8337);
and U8926 (N_8926,N_8038,N_8467);
and U8927 (N_8927,N_8104,N_8174);
nor U8928 (N_8928,N_8278,N_8018);
and U8929 (N_8929,N_8163,N_8382);
nand U8930 (N_8930,N_8381,N_8329);
or U8931 (N_8931,N_8076,N_8242);
or U8932 (N_8932,N_8258,N_8288);
or U8933 (N_8933,N_8472,N_8049);
nand U8934 (N_8934,N_8473,N_8113);
or U8935 (N_8935,N_8288,N_8101);
xor U8936 (N_8936,N_8486,N_8149);
nand U8937 (N_8937,N_8475,N_8005);
nor U8938 (N_8938,N_8007,N_8282);
nand U8939 (N_8939,N_8411,N_8073);
or U8940 (N_8940,N_8039,N_8431);
nand U8941 (N_8941,N_8467,N_8082);
and U8942 (N_8942,N_8204,N_8223);
and U8943 (N_8943,N_8130,N_8194);
and U8944 (N_8944,N_8403,N_8390);
nand U8945 (N_8945,N_8319,N_8447);
xnor U8946 (N_8946,N_8393,N_8032);
nand U8947 (N_8947,N_8285,N_8388);
or U8948 (N_8948,N_8403,N_8361);
and U8949 (N_8949,N_8460,N_8189);
or U8950 (N_8950,N_8311,N_8238);
xor U8951 (N_8951,N_8265,N_8031);
or U8952 (N_8952,N_8042,N_8414);
or U8953 (N_8953,N_8420,N_8397);
nor U8954 (N_8954,N_8438,N_8489);
or U8955 (N_8955,N_8193,N_8255);
and U8956 (N_8956,N_8442,N_8051);
or U8957 (N_8957,N_8358,N_8319);
and U8958 (N_8958,N_8327,N_8043);
and U8959 (N_8959,N_8089,N_8334);
or U8960 (N_8960,N_8271,N_8298);
nand U8961 (N_8961,N_8153,N_8481);
nor U8962 (N_8962,N_8019,N_8205);
or U8963 (N_8963,N_8331,N_8291);
and U8964 (N_8964,N_8458,N_8206);
nor U8965 (N_8965,N_8208,N_8322);
or U8966 (N_8966,N_8160,N_8067);
nor U8967 (N_8967,N_8246,N_8383);
nor U8968 (N_8968,N_8124,N_8344);
and U8969 (N_8969,N_8030,N_8141);
and U8970 (N_8970,N_8316,N_8228);
or U8971 (N_8971,N_8203,N_8146);
or U8972 (N_8972,N_8110,N_8395);
and U8973 (N_8973,N_8157,N_8371);
nand U8974 (N_8974,N_8191,N_8440);
nor U8975 (N_8975,N_8172,N_8282);
xor U8976 (N_8976,N_8465,N_8346);
nand U8977 (N_8977,N_8235,N_8138);
and U8978 (N_8978,N_8382,N_8430);
or U8979 (N_8979,N_8216,N_8437);
and U8980 (N_8980,N_8441,N_8434);
and U8981 (N_8981,N_8160,N_8354);
nor U8982 (N_8982,N_8312,N_8140);
nor U8983 (N_8983,N_8196,N_8232);
nor U8984 (N_8984,N_8134,N_8164);
or U8985 (N_8985,N_8194,N_8449);
xnor U8986 (N_8986,N_8294,N_8306);
nor U8987 (N_8987,N_8096,N_8148);
nor U8988 (N_8988,N_8242,N_8350);
xor U8989 (N_8989,N_8237,N_8481);
or U8990 (N_8990,N_8335,N_8025);
and U8991 (N_8991,N_8480,N_8015);
nand U8992 (N_8992,N_8294,N_8005);
nand U8993 (N_8993,N_8183,N_8265);
or U8994 (N_8994,N_8244,N_8440);
xor U8995 (N_8995,N_8266,N_8014);
or U8996 (N_8996,N_8069,N_8027);
or U8997 (N_8997,N_8007,N_8094);
nand U8998 (N_8998,N_8322,N_8072);
nand U8999 (N_8999,N_8370,N_8042);
xnor U9000 (N_9000,N_8589,N_8966);
nand U9001 (N_9001,N_8780,N_8871);
and U9002 (N_9002,N_8773,N_8869);
and U9003 (N_9003,N_8691,N_8853);
nor U9004 (N_9004,N_8860,N_8760);
nor U9005 (N_9005,N_8502,N_8587);
and U9006 (N_9006,N_8920,N_8891);
nor U9007 (N_9007,N_8796,N_8875);
and U9008 (N_9008,N_8671,N_8595);
xnor U9009 (N_9009,N_8872,N_8880);
nand U9010 (N_9010,N_8904,N_8665);
nand U9011 (N_9011,N_8682,N_8890);
nor U9012 (N_9012,N_8503,N_8652);
nand U9013 (N_9013,N_8613,N_8805);
nand U9014 (N_9014,N_8969,N_8584);
or U9015 (N_9015,N_8590,N_8634);
nand U9016 (N_9016,N_8812,N_8896);
or U9017 (N_9017,N_8789,N_8585);
or U9018 (N_9018,N_8995,N_8688);
nand U9019 (N_9019,N_8928,N_8670);
or U9020 (N_9020,N_8628,N_8675);
xor U9021 (N_9021,N_8599,N_8787);
and U9022 (N_9022,N_8956,N_8882);
nor U9023 (N_9023,N_8817,N_8727);
and U9024 (N_9024,N_8603,N_8678);
and U9025 (N_9025,N_8621,N_8862);
or U9026 (N_9026,N_8982,N_8709);
nand U9027 (N_9027,N_8838,N_8627);
nor U9028 (N_9028,N_8633,N_8537);
nand U9029 (N_9029,N_8522,N_8570);
nand U9030 (N_9030,N_8563,N_8915);
or U9031 (N_9031,N_8663,N_8979);
or U9032 (N_9032,N_8819,N_8782);
and U9033 (N_9033,N_8724,N_8818);
or U9034 (N_9034,N_8978,N_8643);
nor U9035 (N_9035,N_8770,N_8746);
and U9036 (N_9036,N_8935,N_8861);
nand U9037 (N_9037,N_8857,N_8751);
xnor U9038 (N_9038,N_8834,N_8912);
and U9039 (N_9039,N_8926,N_8743);
nor U9040 (N_9040,N_8656,N_8514);
nor U9041 (N_9041,N_8703,N_8747);
nand U9042 (N_9042,N_8850,N_8874);
and U9043 (N_9043,N_8843,N_8661);
or U9044 (N_9044,N_8863,N_8500);
nand U9045 (N_9045,N_8555,N_8545);
nor U9046 (N_9046,N_8944,N_8901);
and U9047 (N_9047,N_8933,N_8638);
and U9048 (N_9048,N_8837,N_8740);
or U9049 (N_9049,N_8771,N_8617);
or U9050 (N_9050,N_8594,N_8681);
or U9051 (N_9051,N_8521,N_8799);
and U9052 (N_9052,N_8801,N_8717);
nand U9053 (N_9053,N_8741,N_8677);
nand U9054 (N_9054,N_8794,N_8898);
nor U9055 (N_9055,N_8826,N_8878);
nand U9056 (N_9056,N_8839,N_8856);
or U9057 (N_9057,N_8811,N_8532);
nor U9058 (N_9058,N_8632,N_8757);
nor U9059 (N_9059,N_8824,N_8636);
nor U9060 (N_9060,N_8650,N_8725);
nand U9061 (N_9061,N_8997,N_8547);
nor U9062 (N_9062,N_8985,N_8629);
nor U9063 (N_9063,N_8511,N_8753);
nand U9064 (N_9064,N_8833,N_8961);
or U9065 (N_9065,N_8533,N_8560);
nor U9066 (N_9066,N_8695,N_8778);
and U9067 (N_9067,N_8802,N_8637);
nand U9068 (N_9068,N_8921,N_8945);
or U9069 (N_9069,N_8752,N_8842);
and U9070 (N_9070,N_8685,N_8649);
or U9071 (N_9071,N_8994,N_8932);
nor U9072 (N_9072,N_8948,N_8776);
nand U9073 (N_9073,N_8607,N_8750);
nand U9074 (N_9074,N_8957,N_8561);
or U9075 (N_9075,N_8669,N_8586);
nor U9076 (N_9076,N_8601,N_8855);
xnor U9077 (N_9077,N_8798,N_8544);
nand U9078 (N_9078,N_8734,N_8516);
nor U9079 (N_9079,N_8943,N_8934);
nand U9080 (N_9080,N_8914,N_8714);
and U9081 (N_9081,N_8726,N_8907);
xor U9082 (N_9082,N_8910,N_8523);
or U9083 (N_9083,N_8729,N_8791);
xnor U9084 (N_9084,N_8518,N_8885);
nor U9085 (N_9085,N_8832,N_8936);
or U9086 (N_9086,N_8785,N_8639);
or U9087 (N_9087,N_8686,N_8528);
nand U9088 (N_9088,N_8998,N_8930);
nor U9089 (N_9089,N_8551,N_8951);
and U9090 (N_9090,N_8755,N_8536);
and U9091 (N_9091,N_8761,N_8909);
or U9092 (N_9092,N_8575,N_8504);
nand U9093 (N_9093,N_8783,N_8911);
nor U9094 (N_9094,N_8611,N_8772);
nand U9095 (N_9095,N_8831,N_8823);
and U9096 (N_9096,N_8604,N_8836);
nand U9097 (N_9097,N_8800,N_8655);
nand U9098 (N_9098,N_8572,N_8540);
nand U9099 (N_9099,N_8647,N_8756);
or U9100 (N_9100,N_8806,N_8923);
nand U9101 (N_9101,N_8881,N_8640);
nand U9102 (N_9102,N_8793,N_8868);
xor U9103 (N_9103,N_8707,N_8705);
nor U9104 (N_9104,N_8674,N_8990);
nor U9105 (N_9105,N_8645,N_8596);
nand U9106 (N_9106,N_8929,N_8615);
nand U9107 (N_9107,N_8538,N_8716);
nor U9108 (N_9108,N_8680,N_8892);
and U9109 (N_9109,N_8947,N_8973);
or U9110 (N_9110,N_8720,N_8989);
nand U9111 (N_9111,N_8942,N_8676);
and U9112 (N_9112,N_8507,N_8769);
nand U9113 (N_9113,N_8513,N_8664);
nand U9114 (N_9114,N_8510,N_8712);
nand U9115 (N_9115,N_8758,N_8512);
and U9116 (N_9116,N_8991,N_8775);
or U9117 (N_9117,N_8918,N_8554);
nor U9118 (N_9118,N_8900,N_8583);
or U9119 (N_9119,N_8981,N_8902);
nor U9120 (N_9120,N_8524,N_8795);
xor U9121 (N_9121,N_8964,N_8591);
or U9122 (N_9122,N_8672,N_8975);
nand U9123 (N_9123,N_8535,N_8745);
xor U9124 (N_9124,N_8807,N_8899);
and U9125 (N_9125,N_8764,N_8949);
and U9126 (N_9126,N_8866,N_8515);
and U9127 (N_9127,N_8840,N_8849);
nand U9128 (N_9128,N_8765,N_8820);
nand U9129 (N_9129,N_8955,N_8865);
nor U9130 (N_9130,N_8684,N_8623);
or U9131 (N_9131,N_8530,N_8895);
nand U9132 (N_9132,N_8959,N_8905);
xor U9133 (N_9133,N_8694,N_8592);
or U9134 (N_9134,N_8704,N_8574);
xnor U9135 (N_9135,N_8786,N_8618);
and U9136 (N_9136,N_8852,N_8630);
nor U9137 (N_9137,N_8814,N_8550);
and U9138 (N_9138,N_8673,N_8619);
or U9139 (N_9139,N_8542,N_8602);
xnor U9140 (N_9140,N_8922,N_8917);
and U9141 (N_9141,N_8557,N_8767);
nand U9142 (N_9142,N_8830,N_8988);
or U9143 (N_9143,N_8809,N_8897);
or U9144 (N_9144,N_8748,N_8658);
nand U9145 (N_9145,N_8626,N_8841);
and U9146 (N_9146,N_8701,N_8567);
nor U9147 (N_9147,N_8854,N_8762);
nor U9148 (N_9148,N_8744,N_8559);
or U9149 (N_9149,N_8941,N_8562);
or U9150 (N_9150,N_8582,N_8713);
nand U9151 (N_9151,N_8822,N_8960);
nand U9152 (N_9152,N_8784,N_8827);
xnor U9153 (N_9153,N_8710,N_8699);
nand U9154 (N_9154,N_8763,N_8702);
and U9155 (N_9155,N_8527,N_8730);
nand U9156 (N_9156,N_8877,N_8999);
nand U9157 (N_9157,N_8723,N_8579);
and U9158 (N_9158,N_8883,N_8828);
and U9159 (N_9159,N_8573,N_8858);
nor U9160 (N_9160,N_8846,N_8690);
xor U9161 (N_9161,N_8644,N_8668);
nor U9162 (N_9162,N_8593,N_8870);
nand U9163 (N_9163,N_8946,N_8777);
or U9164 (N_9164,N_8987,N_8976);
nand U9165 (N_9165,N_8908,N_8864);
nor U9166 (N_9166,N_8708,N_8706);
nor U9167 (N_9167,N_8736,N_8968);
nand U9168 (N_9168,N_8816,N_8641);
or U9169 (N_9169,N_8893,N_8938);
and U9170 (N_9170,N_8894,N_8971);
nor U9171 (N_9171,N_8581,N_8625);
or U9172 (N_9172,N_8738,N_8648);
nor U9173 (N_9173,N_8851,N_8867);
nand U9174 (N_9174,N_8580,N_8697);
xor U9175 (N_9175,N_8578,N_8693);
nor U9176 (N_9176,N_8733,N_8835);
nand U9177 (N_9177,N_8808,N_8813);
nand U9178 (N_9178,N_8829,N_8937);
and U9179 (N_9179,N_8597,N_8768);
nor U9180 (N_9180,N_8919,N_8543);
and U9181 (N_9181,N_8631,N_8552);
nor U9182 (N_9182,N_8667,N_8963);
and U9183 (N_9183,N_8577,N_8742);
xnor U9184 (N_9184,N_8931,N_8588);
or U9185 (N_9185,N_8689,N_8803);
and U9186 (N_9186,N_8598,N_8501);
and U9187 (N_9187,N_8698,N_8605);
and U9188 (N_9188,N_8531,N_8654);
or U9189 (N_9189,N_8821,N_8749);
nor U9190 (N_9190,N_8692,N_8952);
xnor U9191 (N_9191,N_8759,N_8984);
xor U9192 (N_9192,N_8506,N_8983);
and U9193 (N_9193,N_8566,N_8666);
nand U9194 (N_9194,N_8642,N_8549);
and U9195 (N_9195,N_8810,N_8711);
nor U9196 (N_9196,N_8620,N_8509);
nand U9197 (N_9197,N_8953,N_8600);
and U9198 (N_9198,N_8887,N_8974);
or U9199 (N_9199,N_8790,N_8614);
nand U9200 (N_9200,N_8848,N_8906);
nand U9201 (N_9201,N_8722,N_8739);
nand U9202 (N_9202,N_8565,N_8608);
nand U9203 (N_9203,N_8967,N_8815);
and U9204 (N_9204,N_8992,N_8525);
nor U9205 (N_9205,N_8859,N_8616);
xnor U9206 (N_9206,N_8541,N_8606);
nor U9207 (N_9207,N_8996,N_8927);
nor U9208 (N_9208,N_8986,N_8735);
or U9209 (N_9209,N_8825,N_8779);
nand U9210 (N_9210,N_8657,N_8888);
xor U9211 (N_9211,N_8972,N_8646);
nor U9212 (N_9212,N_8965,N_8553);
xnor U9213 (N_9213,N_8556,N_8766);
nand U9214 (N_9214,N_8774,N_8970);
nand U9215 (N_9215,N_8925,N_8876);
xnor U9216 (N_9216,N_8653,N_8879);
nand U9217 (N_9217,N_8719,N_8505);
nand U9218 (N_9218,N_8700,N_8950);
xor U9219 (N_9219,N_8508,N_8954);
or U9220 (N_9220,N_8886,N_8715);
nand U9221 (N_9221,N_8526,N_8977);
xor U9222 (N_9222,N_8564,N_8958);
or U9223 (N_9223,N_8718,N_8939);
or U9224 (N_9224,N_8962,N_8610);
nor U9225 (N_9225,N_8683,N_8844);
or U9226 (N_9226,N_8781,N_8662);
or U9227 (N_9227,N_8696,N_8558);
nand U9228 (N_9228,N_8635,N_8847);
or U9229 (N_9229,N_8940,N_8721);
or U9230 (N_9230,N_8609,N_8884);
nand U9231 (N_9231,N_8804,N_8916);
or U9232 (N_9232,N_8576,N_8754);
nor U9233 (N_9233,N_8659,N_8548);
nor U9234 (N_9234,N_8569,N_8529);
and U9235 (N_9235,N_8519,N_8980);
nor U9236 (N_9236,N_8792,N_8913);
or U9237 (N_9237,N_8546,N_8889);
xnor U9238 (N_9238,N_8520,N_8534);
nor U9239 (N_9239,N_8788,N_8651);
nor U9240 (N_9240,N_8612,N_8624);
nand U9241 (N_9241,N_8731,N_8728);
nor U9242 (N_9242,N_8903,N_8687);
or U9243 (N_9243,N_8517,N_8660);
and U9244 (N_9244,N_8679,N_8797);
xnor U9245 (N_9245,N_8845,N_8539);
nor U9246 (N_9246,N_8622,N_8568);
or U9247 (N_9247,N_8732,N_8993);
nand U9248 (N_9248,N_8737,N_8873);
or U9249 (N_9249,N_8571,N_8924);
and U9250 (N_9250,N_8971,N_8781);
nor U9251 (N_9251,N_8869,N_8674);
nor U9252 (N_9252,N_8500,N_8852);
nor U9253 (N_9253,N_8820,N_8721);
xnor U9254 (N_9254,N_8743,N_8551);
nor U9255 (N_9255,N_8588,N_8669);
or U9256 (N_9256,N_8760,N_8866);
and U9257 (N_9257,N_8907,N_8879);
nor U9258 (N_9258,N_8651,N_8557);
nor U9259 (N_9259,N_8914,N_8814);
nor U9260 (N_9260,N_8684,N_8643);
and U9261 (N_9261,N_8657,N_8794);
or U9262 (N_9262,N_8869,N_8789);
or U9263 (N_9263,N_8953,N_8745);
nor U9264 (N_9264,N_8812,N_8986);
nor U9265 (N_9265,N_8522,N_8938);
nand U9266 (N_9266,N_8623,N_8931);
nor U9267 (N_9267,N_8600,N_8745);
nor U9268 (N_9268,N_8708,N_8772);
nand U9269 (N_9269,N_8560,N_8845);
nor U9270 (N_9270,N_8732,N_8935);
nand U9271 (N_9271,N_8560,N_8890);
nor U9272 (N_9272,N_8628,N_8742);
or U9273 (N_9273,N_8692,N_8879);
nand U9274 (N_9274,N_8908,N_8640);
nor U9275 (N_9275,N_8784,N_8592);
xnor U9276 (N_9276,N_8885,N_8810);
xnor U9277 (N_9277,N_8542,N_8977);
and U9278 (N_9278,N_8923,N_8605);
or U9279 (N_9279,N_8913,N_8832);
and U9280 (N_9280,N_8595,N_8704);
and U9281 (N_9281,N_8756,N_8925);
or U9282 (N_9282,N_8568,N_8781);
and U9283 (N_9283,N_8572,N_8569);
nor U9284 (N_9284,N_8593,N_8722);
xnor U9285 (N_9285,N_8642,N_8877);
or U9286 (N_9286,N_8873,N_8976);
nor U9287 (N_9287,N_8591,N_8873);
and U9288 (N_9288,N_8586,N_8576);
xor U9289 (N_9289,N_8849,N_8545);
or U9290 (N_9290,N_8545,N_8719);
and U9291 (N_9291,N_8783,N_8519);
nand U9292 (N_9292,N_8964,N_8563);
or U9293 (N_9293,N_8637,N_8699);
or U9294 (N_9294,N_8624,N_8895);
or U9295 (N_9295,N_8727,N_8764);
xor U9296 (N_9296,N_8660,N_8688);
nor U9297 (N_9297,N_8919,N_8874);
and U9298 (N_9298,N_8595,N_8964);
or U9299 (N_9299,N_8741,N_8959);
nand U9300 (N_9300,N_8764,N_8587);
or U9301 (N_9301,N_8770,N_8905);
and U9302 (N_9302,N_8664,N_8859);
or U9303 (N_9303,N_8799,N_8543);
nor U9304 (N_9304,N_8680,N_8818);
xnor U9305 (N_9305,N_8554,N_8576);
or U9306 (N_9306,N_8725,N_8727);
nand U9307 (N_9307,N_8578,N_8990);
xor U9308 (N_9308,N_8703,N_8608);
nand U9309 (N_9309,N_8547,N_8965);
xor U9310 (N_9310,N_8968,N_8657);
xnor U9311 (N_9311,N_8613,N_8960);
or U9312 (N_9312,N_8869,N_8858);
or U9313 (N_9313,N_8918,N_8843);
nand U9314 (N_9314,N_8548,N_8838);
nor U9315 (N_9315,N_8558,N_8622);
nor U9316 (N_9316,N_8655,N_8552);
and U9317 (N_9317,N_8529,N_8604);
and U9318 (N_9318,N_8690,N_8743);
and U9319 (N_9319,N_8991,N_8540);
and U9320 (N_9320,N_8544,N_8503);
and U9321 (N_9321,N_8625,N_8915);
or U9322 (N_9322,N_8584,N_8888);
xnor U9323 (N_9323,N_8583,N_8802);
or U9324 (N_9324,N_8611,N_8705);
nand U9325 (N_9325,N_8853,N_8832);
and U9326 (N_9326,N_8824,N_8996);
xor U9327 (N_9327,N_8776,N_8605);
nand U9328 (N_9328,N_8525,N_8603);
and U9329 (N_9329,N_8615,N_8743);
xor U9330 (N_9330,N_8762,N_8654);
nor U9331 (N_9331,N_8757,N_8864);
and U9332 (N_9332,N_8677,N_8869);
or U9333 (N_9333,N_8910,N_8822);
and U9334 (N_9334,N_8733,N_8833);
xnor U9335 (N_9335,N_8999,N_8766);
nor U9336 (N_9336,N_8522,N_8516);
and U9337 (N_9337,N_8995,N_8996);
nand U9338 (N_9338,N_8942,N_8893);
nand U9339 (N_9339,N_8687,N_8577);
nor U9340 (N_9340,N_8999,N_8714);
nand U9341 (N_9341,N_8931,N_8506);
nand U9342 (N_9342,N_8745,N_8766);
nor U9343 (N_9343,N_8837,N_8624);
and U9344 (N_9344,N_8998,N_8581);
and U9345 (N_9345,N_8912,N_8907);
or U9346 (N_9346,N_8757,N_8669);
and U9347 (N_9347,N_8587,N_8965);
and U9348 (N_9348,N_8565,N_8629);
nor U9349 (N_9349,N_8590,N_8575);
xnor U9350 (N_9350,N_8659,N_8621);
nand U9351 (N_9351,N_8855,N_8534);
nor U9352 (N_9352,N_8608,N_8645);
and U9353 (N_9353,N_8844,N_8576);
and U9354 (N_9354,N_8859,N_8924);
and U9355 (N_9355,N_8932,N_8737);
or U9356 (N_9356,N_8899,N_8992);
and U9357 (N_9357,N_8644,N_8897);
and U9358 (N_9358,N_8560,N_8684);
nand U9359 (N_9359,N_8883,N_8955);
nor U9360 (N_9360,N_8719,N_8905);
or U9361 (N_9361,N_8939,N_8541);
or U9362 (N_9362,N_8551,N_8977);
nor U9363 (N_9363,N_8903,N_8583);
or U9364 (N_9364,N_8977,N_8831);
and U9365 (N_9365,N_8977,N_8556);
and U9366 (N_9366,N_8664,N_8675);
nor U9367 (N_9367,N_8982,N_8838);
and U9368 (N_9368,N_8854,N_8611);
nor U9369 (N_9369,N_8760,N_8953);
and U9370 (N_9370,N_8893,N_8678);
nand U9371 (N_9371,N_8651,N_8947);
nor U9372 (N_9372,N_8640,N_8693);
nand U9373 (N_9373,N_8554,N_8795);
or U9374 (N_9374,N_8526,N_8514);
or U9375 (N_9375,N_8771,N_8650);
nand U9376 (N_9376,N_8854,N_8639);
nor U9377 (N_9377,N_8936,N_8625);
nand U9378 (N_9378,N_8644,N_8972);
nor U9379 (N_9379,N_8976,N_8707);
nor U9380 (N_9380,N_8522,N_8978);
and U9381 (N_9381,N_8571,N_8663);
xor U9382 (N_9382,N_8754,N_8765);
and U9383 (N_9383,N_8993,N_8668);
and U9384 (N_9384,N_8787,N_8752);
nor U9385 (N_9385,N_8672,N_8654);
xor U9386 (N_9386,N_8888,N_8634);
or U9387 (N_9387,N_8922,N_8510);
nor U9388 (N_9388,N_8955,N_8810);
and U9389 (N_9389,N_8788,N_8728);
and U9390 (N_9390,N_8735,N_8985);
xnor U9391 (N_9391,N_8947,N_8946);
nor U9392 (N_9392,N_8977,N_8686);
and U9393 (N_9393,N_8777,N_8589);
or U9394 (N_9394,N_8573,N_8527);
nand U9395 (N_9395,N_8978,N_8766);
xor U9396 (N_9396,N_8560,N_8521);
or U9397 (N_9397,N_8733,N_8888);
nand U9398 (N_9398,N_8875,N_8663);
nand U9399 (N_9399,N_8544,N_8678);
and U9400 (N_9400,N_8655,N_8885);
nor U9401 (N_9401,N_8622,N_8870);
and U9402 (N_9402,N_8772,N_8985);
and U9403 (N_9403,N_8573,N_8678);
nand U9404 (N_9404,N_8943,N_8595);
or U9405 (N_9405,N_8766,N_8674);
and U9406 (N_9406,N_8783,N_8805);
and U9407 (N_9407,N_8648,N_8562);
or U9408 (N_9408,N_8700,N_8666);
nor U9409 (N_9409,N_8879,N_8698);
or U9410 (N_9410,N_8905,N_8844);
xor U9411 (N_9411,N_8621,N_8840);
or U9412 (N_9412,N_8993,N_8891);
nand U9413 (N_9413,N_8905,N_8780);
nor U9414 (N_9414,N_8739,N_8547);
and U9415 (N_9415,N_8906,N_8574);
xor U9416 (N_9416,N_8965,N_8790);
xor U9417 (N_9417,N_8636,N_8534);
or U9418 (N_9418,N_8637,N_8868);
or U9419 (N_9419,N_8892,N_8670);
and U9420 (N_9420,N_8620,N_8852);
nand U9421 (N_9421,N_8726,N_8656);
nor U9422 (N_9422,N_8748,N_8790);
nand U9423 (N_9423,N_8572,N_8831);
or U9424 (N_9424,N_8646,N_8631);
and U9425 (N_9425,N_8611,N_8590);
nor U9426 (N_9426,N_8899,N_8834);
and U9427 (N_9427,N_8727,N_8572);
and U9428 (N_9428,N_8681,N_8535);
and U9429 (N_9429,N_8539,N_8725);
or U9430 (N_9430,N_8528,N_8898);
and U9431 (N_9431,N_8831,N_8773);
or U9432 (N_9432,N_8793,N_8525);
or U9433 (N_9433,N_8993,N_8924);
nand U9434 (N_9434,N_8597,N_8516);
xor U9435 (N_9435,N_8760,N_8755);
and U9436 (N_9436,N_8886,N_8698);
nor U9437 (N_9437,N_8789,N_8726);
nand U9438 (N_9438,N_8728,N_8598);
nand U9439 (N_9439,N_8676,N_8975);
nand U9440 (N_9440,N_8883,N_8503);
nand U9441 (N_9441,N_8785,N_8545);
nand U9442 (N_9442,N_8704,N_8815);
nand U9443 (N_9443,N_8803,N_8556);
and U9444 (N_9444,N_8994,N_8676);
xor U9445 (N_9445,N_8717,N_8568);
xnor U9446 (N_9446,N_8746,N_8925);
nand U9447 (N_9447,N_8945,N_8553);
or U9448 (N_9448,N_8844,N_8635);
and U9449 (N_9449,N_8806,N_8818);
and U9450 (N_9450,N_8561,N_8502);
or U9451 (N_9451,N_8595,N_8903);
and U9452 (N_9452,N_8803,N_8540);
nor U9453 (N_9453,N_8830,N_8736);
xnor U9454 (N_9454,N_8787,N_8523);
and U9455 (N_9455,N_8513,N_8556);
nand U9456 (N_9456,N_8987,N_8741);
and U9457 (N_9457,N_8869,N_8855);
and U9458 (N_9458,N_8852,N_8936);
nor U9459 (N_9459,N_8659,N_8535);
xor U9460 (N_9460,N_8649,N_8515);
nand U9461 (N_9461,N_8832,N_8701);
or U9462 (N_9462,N_8808,N_8848);
nor U9463 (N_9463,N_8967,N_8589);
nor U9464 (N_9464,N_8979,N_8710);
and U9465 (N_9465,N_8885,N_8658);
and U9466 (N_9466,N_8625,N_8839);
xnor U9467 (N_9467,N_8703,N_8872);
and U9468 (N_9468,N_8611,N_8574);
nor U9469 (N_9469,N_8891,N_8504);
and U9470 (N_9470,N_8517,N_8635);
or U9471 (N_9471,N_8618,N_8798);
or U9472 (N_9472,N_8959,N_8667);
nand U9473 (N_9473,N_8802,N_8696);
nand U9474 (N_9474,N_8540,N_8855);
or U9475 (N_9475,N_8804,N_8722);
nand U9476 (N_9476,N_8529,N_8626);
nand U9477 (N_9477,N_8678,N_8752);
nor U9478 (N_9478,N_8775,N_8641);
or U9479 (N_9479,N_8903,N_8695);
nor U9480 (N_9480,N_8581,N_8993);
nand U9481 (N_9481,N_8668,N_8699);
or U9482 (N_9482,N_8633,N_8779);
xnor U9483 (N_9483,N_8881,N_8776);
and U9484 (N_9484,N_8680,N_8839);
and U9485 (N_9485,N_8538,N_8809);
nand U9486 (N_9486,N_8533,N_8640);
xnor U9487 (N_9487,N_8816,N_8737);
and U9488 (N_9488,N_8546,N_8867);
or U9489 (N_9489,N_8712,N_8578);
or U9490 (N_9490,N_8524,N_8762);
and U9491 (N_9491,N_8888,N_8923);
nor U9492 (N_9492,N_8664,N_8623);
or U9493 (N_9493,N_8762,N_8764);
nor U9494 (N_9494,N_8899,N_8728);
or U9495 (N_9495,N_8561,N_8733);
nand U9496 (N_9496,N_8948,N_8922);
or U9497 (N_9497,N_8543,N_8539);
and U9498 (N_9498,N_8635,N_8838);
nor U9499 (N_9499,N_8791,N_8903);
nand U9500 (N_9500,N_9218,N_9342);
xnor U9501 (N_9501,N_9232,N_9375);
and U9502 (N_9502,N_9301,N_9182);
and U9503 (N_9503,N_9118,N_9429);
and U9504 (N_9504,N_9496,N_9236);
and U9505 (N_9505,N_9312,N_9169);
or U9506 (N_9506,N_9122,N_9027);
nand U9507 (N_9507,N_9059,N_9066);
nand U9508 (N_9508,N_9190,N_9069);
nor U9509 (N_9509,N_9061,N_9436);
or U9510 (N_9510,N_9444,N_9425);
nand U9511 (N_9511,N_9217,N_9263);
nand U9512 (N_9512,N_9349,N_9255);
or U9513 (N_9513,N_9078,N_9421);
nand U9514 (N_9514,N_9120,N_9102);
nor U9515 (N_9515,N_9195,N_9030);
nor U9516 (N_9516,N_9464,N_9274);
nand U9517 (N_9517,N_9399,N_9362);
nor U9518 (N_9518,N_9402,N_9155);
nor U9519 (N_9519,N_9447,N_9446);
and U9520 (N_9520,N_9434,N_9032);
nor U9521 (N_9521,N_9415,N_9337);
and U9522 (N_9522,N_9035,N_9076);
nor U9523 (N_9523,N_9260,N_9098);
nand U9524 (N_9524,N_9373,N_9156);
nand U9525 (N_9525,N_9177,N_9314);
xnor U9526 (N_9526,N_9105,N_9485);
nor U9527 (N_9527,N_9132,N_9227);
and U9528 (N_9528,N_9298,N_9046);
and U9529 (N_9529,N_9081,N_9219);
or U9530 (N_9530,N_9367,N_9345);
nor U9531 (N_9531,N_9222,N_9137);
or U9532 (N_9532,N_9273,N_9110);
and U9533 (N_9533,N_9271,N_9099);
or U9534 (N_9534,N_9481,N_9103);
nand U9535 (N_9535,N_9168,N_9051);
xor U9536 (N_9536,N_9248,N_9378);
nand U9537 (N_9537,N_9489,N_9357);
or U9538 (N_9538,N_9256,N_9004);
xnor U9539 (N_9539,N_9318,N_9072);
nor U9540 (N_9540,N_9281,N_9224);
and U9541 (N_9541,N_9463,N_9238);
nor U9542 (N_9542,N_9055,N_9426);
and U9543 (N_9543,N_9029,N_9131);
nand U9544 (N_9544,N_9171,N_9358);
nand U9545 (N_9545,N_9243,N_9453);
xnor U9546 (N_9546,N_9012,N_9418);
nor U9547 (N_9547,N_9254,N_9094);
and U9548 (N_9548,N_9139,N_9422);
xnor U9549 (N_9549,N_9466,N_9336);
xnor U9550 (N_9550,N_9075,N_9441);
nor U9551 (N_9551,N_9006,N_9036);
xor U9552 (N_9552,N_9235,N_9244);
nand U9553 (N_9553,N_9183,N_9034);
nor U9554 (N_9554,N_9424,N_9465);
nor U9555 (N_9555,N_9347,N_9293);
nor U9556 (N_9556,N_9354,N_9319);
nor U9557 (N_9557,N_9024,N_9449);
xor U9558 (N_9558,N_9133,N_9262);
and U9559 (N_9559,N_9161,N_9246);
or U9560 (N_9560,N_9049,N_9136);
nor U9561 (N_9561,N_9234,N_9428);
and U9562 (N_9562,N_9292,N_9186);
or U9563 (N_9563,N_9355,N_9296);
and U9564 (N_9564,N_9162,N_9390);
nand U9565 (N_9565,N_9229,N_9269);
and U9566 (N_9566,N_9460,N_9491);
or U9567 (N_9567,N_9450,N_9164);
nand U9568 (N_9568,N_9093,N_9279);
xnor U9569 (N_9569,N_9041,N_9458);
nand U9570 (N_9570,N_9062,N_9052);
and U9571 (N_9571,N_9070,N_9258);
and U9572 (N_9572,N_9230,N_9208);
nor U9573 (N_9573,N_9050,N_9384);
or U9574 (N_9574,N_9083,N_9172);
or U9575 (N_9575,N_9495,N_9247);
nor U9576 (N_9576,N_9225,N_9060);
nor U9577 (N_9577,N_9149,N_9025);
nand U9578 (N_9578,N_9226,N_9023);
nand U9579 (N_9579,N_9391,N_9115);
nand U9580 (N_9580,N_9474,N_9303);
nand U9581 (N_9581,N_9278,N_9090);
nand U9582 (N_9582,N_9284,N_9443);
nand U9583 (N_9583,N_9416,N_9205);
nor U9584 (N_9584,N_9328,N_9175);
and U9585 (N_9585,N_9045,N_9397);
and U9586 (N_9586,N_9321,N_9287);
and U9587 (N_9587,N_9191,N_9251);
or U9588 (N_9588,N_9154,N_9374);
nor U9589 (N_9589,N_9356,N_9343);
nand U9590 (N_9590,N_9000,N_9308);
nor U9591 (N_9591,N_9112,N_9237);
and U9592 (N_9592,N_9400,N_9233);
nand U9593 (N_9593,N_9488,N_9280);
nand U9594 (N_9594,N_9445,N_9272);
nor U9595 (N_9595,N_9268,N_9001);
nand U9596 (N_9596,N_9092,N_9123);
nand U9597 (N_9597,N_9077,N_9184);
and U9598 (N_9598,N_9145,N_9157);
and U9599 (N_9599,N_9207,N_9146);
or U9600 (N_9600,N_9338,N_9439);
and U9601 (N_9601,N_9325,N_9039);
and U9602 (N_9602,N_9265,N_9142);
nand U9603 (N_9603,N_9043,N_9388);
xnor U9604 (N_9604,N_9433,N_9499);
nand U9605 (N_9605,N_9108,N_9179);
or U9606 (N_9606,N_9277,N_9192);
and U9607 (N_9607,N_9461,N_9085);
nand U9608 (N_9608,N_9117,N_9320);
or U9609 (N_9609,N_9166,N_9158);
nand U9610 (N_9610,N_9151,N_9040);
nor U9611 (N_9611,N_9215,N_9437);
and U9612 (N_9612,N_9057,N_9221);
nand U9613 (N_9613,N_9138,N_9253);
nor U9614 (N_9614,N_9140,N_9387);
nand U9615 (N_9615,N_9359,N_9194);
nand U9616 (N_9616,N_9369,N_9323);
xor U9617 (N_9617,N_9412,N_9189);
nor U9618 (N_9618,N_9200,N_9071);
and U9619 (N_9619,N_9020,N_9417);
xor U9620 (N_9620,N_9411,N_9483);
nand U9621 (N_9621,N_9405,N_9173);
nor U9622 (N_9622,N_9315,N_9261);
nand U9623 (N_9623,N_9327,N_9361);
and U9624 (N_9624,N_9409,N_9352);
nor U9625 (N_9625,N_9324,N_9129);
or U9626 (N_9626,N_9119,N_9017);
nand U9627 (N_9627,N_9366,N_9407);
nand U9628 (N_9628,N_9259,N_9150);
or U9629 (N_9629,N_9322,N_9198);
and U9630 (N_9630,N_9372,N_9467);
nand U9631 (N_9631,N_9159,N_9404);
nand U9632 (N_9632,N_9294,N_9365);
xnor U9633 (N_9633,N_9240,N_9199);
nor U9634 (N_9634,N_9126,N_9360);
and U9635 (N_9635,N_9087,N_9497);
nand U9636 (N_9636,N_9239,N_9209);
xor U9637 (N_9637,N_9231,N_9044);
or U9638 (N_9638,N_9165,N_9371);
and U9639 (N_9639,N_9455,N_9220);
and U9640 (N_9640,N_9080,N_9019);
or U9641 (N_9641,N_9468,N_9054);
nand U9642 (N_9642,N_9479,N_9480);
xor U9643 (N_9643,N_9185,N_9282);
nor U9644 (N_9644,N_9064,N_9249);
nor U9645 (N_9645,N_9210,N_9267);
nand U9646 (N_9646,N_9414,N_9038);
nor U9647 (N_9647,N_9058,N_9302);
nand U9648 (N_9648,N_9266,N_9063);
or U9649 (N_9649,N_9478,N_9285);
nor U9650 (N_9650,N_9305,N_9241);
or U9651 (N_9651,N_9385,N_9187);
and U9652 (N_9652,N_9309,N_9289);
and U9653 (N_9653,N_9016,N_9329);
and U9654 (N_9654,N_9068,N_9393);
and U9655 (N_9655,N_9427,N_9291);
nand U9656 (N_9656,N_9176,N_9121);
or U9657 (N_9657,N_9297,N_9410);
and U9658 (N_9658,N_9452,N_9348);
or U9659 (N_9659,N_9128,N_9167);
nor U9660 (N_9660,N_9276,N_9022);
nor U9661 (N_9661,N_9073,N_9015);
xnor U9662 (N_9662,N_9430,N_9379);
nand U9663 (N_9663,N_9475,N_9257);
nand U9664 (N_9664,N_9088,N_9332);
nand U9665 (N_9665,N_9471,N_9037);
nor U9666 (N_9666,N_9107,N_9100);
nor U9667 (N_9667,N_9482,N_9334);
or U9668 (N_9668,N_9440,N_9275);
nand U9669 (N_9669,N_9392,N_9326);
nand U9670 (N_9670,N_9188,N_9346);
and U9671 (N_9671,N_9310,N_9286);
nand U9672 (N_9672,N_9005,N_9330);
or U9673 (N_9673,N_9065,N_9214);
or U9674 (N_9674,N_9096,N_9377);
or U9675 (N_9675,N_9473,N_9290);
xor U9676 (N_9676,N_9484,N_9113);
nand U9677 (N_9677,N_9304,N_9228);
nand U9678 (N_9678,N_9053,N_9344);
or U9679 (N_9679,N_9487,N_9353);
or U9680 (N_9680,N_9370,N_9490);
xor U9681 (N_9681,N_9013,N_9086);
or U9682 (N_9682,N_9106,N_9316);
or U9683 (N_9683,N_9163,N_9389);
nor U9684 (N_9684,N_9420,N_9295);
or U9685 (N_9685,N_9135,N_9395);
or U9686 (N_9686,N_9213,N_9394);
and U9687 (N_9687,N_9147,N_9026);
and U9688 (N_9688,N_9451,N_9494);
and U9689 (N_9689,N_9007,N_9382);
or U9690 (N_9690,N_9242,N_9014);
and U9691 (N_9691,N_9091,N_9144);
xor U9692 (N_9692,N_9398,N_9335);
or U9693 (N_9693,N_9380,N_9386);
xnor U9694 (N_9694,N_9498,N_9376);
or U9695 (N_9695,N_9114,N_9074);
or U9696 (N_9696,N_9442,N_9250);
and U9697 (N_9697,N_9413,N_9307);
nand U9698 (N_9698,N_9454,N_9245);
and U9699 (N_9699,N_9493,N_9300);
nor U9700 (N_9700,N_9435,N_9492);
and U9701 (N_9701,N_9095,N_9201);
and U9702 (N_9702,N_9104,N_9470);
nand U9703 (N_9703,N_9031,N_9202);
nand U9704 (N_9704,N_9010,N_9306);
and U9705 (N_9705,N_9124,N_9042);
and U9706 (N_9706,N_9383,N_9148);
nor U9707 (N_9707,N_9178,N_9180);
nand U9708 (N_9708,N_9211,N_9082);
or U9709 (N_9709,N_9152,N_9403);
or U9710 (N_9710,N_9351,N_9438);
or U9711 (N_9711,N_9127,N_9341);
nand U9712 (N_9712,N_9197,N_9448);
nor U9713 (N_9713,N_9270,N_9456);
or U9714 (N_9714,N_9047,N_9313);
nand U9715 (N_9715,N_9141,N_9028);
and U9716 (N_9716,N_9067,N_9364);
xor U9717 (N_9717,N_9472,N_9339);
xor U9718 (N_9718,N_9048,N_9432);
and U9719 (N_9719,N_9381,N_9196);
and U9720 (N_9720,N_9401,N_9396);
or U9721 (N_9721,N_9143,N_9419);
or U9722 (N_9722,N_9079,N_9476);
or U9723 (N_9723,N_9317,N_9363);
nor U9724 (N_9724,N_9193,N_9011);
nor U9725 (N_9725,N_9340,N_9459);
or U9726 (N_9726,N_9264,N_9408);
xor U9727 (N_9727,N_9223,N_9486);
and U9728 (N_9728,N_9204,N_9368);
nor U9729 (N_9729,N_9252,N_9283);
or U9730 (N_9730,N_9153,N_9206);
or U9731 (N_9731,N_9056,N_9033);
and U9732 (N_9732,N_9212,N_9311);
nor U9733 (N_9733,N_9457,N_9203);
and U9734 (N_9734,N_9021,N_9288);
nor U9735 (N_9735,N_9431,N_9462);
or U9736 (N_9736,N_9125,N_9002);
or U9737 (N_9737,N_9477,N_9130);
and U9738 (N_9738,N_9134,N_9181);
xor U9739 (N_9739,N_9009,N_9097);
nor U9740 (N_9740,N_9469,N_9333);
and U9741 (N_9741,N_9160,N_9018);
nand U9742 (N_9742,N_9109,N_9216);
xor U9743 (N_9743,N_9299,N_9111);
nand U9744 (N_9744,N_9101,N_9008);
and U9745 (N_9745,N_9116,N_9174);
and U9746 (N_9746,N_9084,N_9406);
or U9747 (N_9747,N_9423,N_9331);
xor U9748 (N_9748,N_9003,N_9350);
nand U9749 (N_9749,N_9170,N_9089);
and U9750 (N_9750,N_9368,N_9322);
or U9751 (N_9751,N_9010,N_9442);
or U9752 (N_9752,N_9221,N_9032);
nand U9753 (N_9753,N_9495,N_9300);
and U9754 (N_9754,N_9212,N_9468);
or U9755 (N_9755,N_9133,N_9338);
nor U9756 (N_9756,N_9419,N_9040);
and U9757 (N_9757,N_9247,N_9078);
and U9758 (N_9758,N_9110,N_9297);
nand U9759 (N_9759,N_9451,N_9080);
nand U9760 (N_9760,N_9077,N_9406);
and U9761 (N_9761,N_9005,N_9343);
nor U9762 (N_9762,N_9106,N_9259);
nand U9763 (N_9763,N_9420,N_9247);
and U9764 (N_9764,N_9422,N_9050);
nor U9765 (N_9765,N_9143,N_9184);
and U9766 (N_9766,N_9371,N_9015);
and U9767 (N_9767,N_9378,N_9190);
nand U9768 (N_9768,N_9272,N_9010);
or U9769 (N_9769,N_9321,N_9217);
or U9770 (N_9770,N_9421,N_9154);
and U9771 (N_9771,N_9435,N_9373);
xnor U9772 (N_9772,N_9175,N_9156);
and U9773 (N_9773,N_9361,N_9269);
xnor U9774 (N_9774,N_9318,N_9340);
nand U9775 (N_9775,N_9247,N_9015);
xnor U9776 (N_9776,N_9427,N_9359);
nor U9777 (N_9777,N_9173,N_9133);
or U9778 (N_9778,N_9245,N_9203);
or U9779 (N_9779,N_9399,N_9044);
or U9780 (N_9780,N_9140,N_9336);
and U9781 (N_9781,N_9042,N_9149);
nand U9782 (N_9782,N_9271,N_9320);
nor U9783 (N_9783,N_9128,N_9063);
or U9784 (N_9784,N_9341,N_9486);
nand U9785 (N_9785,N_9133,N_9469);
nand U9786 (N_9786,N_9183,N_9118);
nand U9787 (N_9787,N_9224,N_9163);
nand U9788 (N_9788,N_9374,N_9076);
nand U9789 (N_9789,N_9314,N_9456);
nor U9790 (N_9790,N_9305,N_9353);
nor U9791 (N_9791,N_9050,N_9036);
nor U9792 (N_9792,N_9297,N_9309);
and U9793 (N_9793,N_9301,N_9053);
nor U9794 (N_9794,N_9288,N_9263);
or U9795 (N_9795,N_9259,N_9336);
nor U9796 (N_9796,N_9356,N_9272);
and U9797 (N_9797,N_9001,N_9338);
or U9798 (N_9798,N_9426,N_9304);
and U9799 (N_9799,N_9113,N_9327);
nand U9800 (N_9800,N_9022,N_9207);
nor U9801 (N_9801,N_9024,N_9399);
xnor U9802 (N_9802,N_9212,N_9241);
nor U9803 (N_9803,N_9259,N_9062);
nor U9804 (N_9804,N_9085,N_9046);
or U9805 (N_9805,N_9080,N_9204);
nand U9806 (N_9806,N_9404,N_9342);
nand U9807 (N_9807,N_9282,N_9217);
nor U9808 (N_9808,N_9407,N_9210);
xnor U9809 (N_9809,N_9477,N_9118);
nor U9810 (N_9810,N_9414,N_9451);
nand U9811 (N_9811,N_9471,N_9332);
or U9812 (N_9812,N_9111,N_9118);
and U9813 (N_9813,N_9214,N_9484);
nor U9814 (N_9814,N_9307,N_9373);
nor U9815 (N_9815,N_9255,N_9081);
and U9816 (N_9816,N_9296,N_9237);
and U9817 (N_9817,N_9494,N_9189);
nor U9818 (N_9818,N_9016,N_9380);
nor U9819 (N_9819,N_9401,N_9406);
nor U9820 (N_9820,N_9471,N_9433);
nor U9821 (N_9821,N_9413,N_9189);
and U9822 (N_9822,N_9456,N_9126);
and U9823 (N_9823,N_9071,N_9373);
nand U9824 (N_9824,N_9164,N_9429);
or U9825 (N_9825,N_9160,N_9357);
nor U9826 (N_9826,N_9052,N_9092);
and U9827 (N_9827,N_9460,N_9414);
nor U9828 (N_9828,N_9035,N_9317);
or U9829 (N_9829,N_9470,N_9244);
nand U9830 (N_9830,N_9067,N_9038);
nor U9831 (N_9831,N_9244,N_9284);
nand U9832 (N_9832,N_9238,N_9447);
and U9833 (N_9833,N_9474,N_9003);
and U9834 (N_9834,N_9063,N_9332);
nand U9835 (N_9835,N_9373,N_9481);
nor U9836 (N_9836,N_9343,N_9032);
and U9837 (N_9837,N_9340,N_9363);
nor U9838 (N_9838,N_9412,N_9026);
and U9839 (N_9839,N_9281,N_9122);
or U9840 (N_9840,N_9152,N_9134);
nor U9841 (N_9841,N_9242,N_9203);
and U9842 (N_9842,N_9451,N_9474);
or U9843 (N_9843,N_9136,N_9091);
or U9844 (N_9844,N_9056,N_9240);
nand U9845 (N_9845,N_9377,N_9399);
and U9846 (N_9846,N_9007,N_9373);
nor U9847 (N_9847,N_9194,N_9418);
nor U9848 (N_9848,N_9029,N_9255);
nand U9849 (N_9849,N_9160,N_9097);
or U9850 (N_9850,N_9124,N_9248);
and U9851 (N_9851,N_9009,N_9316);
nor U9852 (N_9852,N_9256,N_9015);
xor U9853 (N_9853,N_9315,N_9487);
nor U9854 (N_9854,N_9220,N_9472);
xor U9855 (N_9855,N_9286,N_9306);
nand U9856 (N_9856,N_9388,N_9038);
or U9857 (N_9857,N_9029,N_9081);
nor U9858 (N_9858,N_9181,N_9205);
nor U9859 (N_9859,N_9297,N_9462);
and U9860 (N_9860,N_9205,N_9422);
xnor U9861 (N_9861,N_9260,N_9054);
and U9862 (N_9862,N_9090,N_9003);
xor U9863 (N_9863,N_9099,N_9257);
or U9864 (N_9864,N_9460,N_9489);
nor U9865 (N_9865,N_9024,N_9117);
or U9866 (N_9866,N_9144,N_9269);
xor U9867 (N_9867,N_9112,N_9333);
xnor U9868 (N_9868,N_9486,N_9111);
nand U9869 (N_9869,N_9492,N_9001);
nand U9870 (N_9870,N_9065,N_9260);
or U9871 (N_9871,N_9275,N_9274);
or U9872 (N_9872,N_9476,N_9173);
nand U9873 (N_9873,N_9021,N_9199);
nand U9874 (N_9874,N_9229,N_9149);
xor U9875 (N_9875,N_9204,N_9006);
and U9876 (N_9876,N_9146,N_9449);
and U9877 (N_9877,N_9141,N_9100);
nand U9878 (N_9878,N_9385,N_9096);
and U9879 (N_9879,N_9345,N_9099);
nor U9880 (N_9880,N_9360,N_9422);
or U9881 (N_9881,N_9424,N_9055);
nor U9882 (N_9882,N_9154,N_9241);
xor U9883 (N_9883,N_9305,N_9043);
xor U9884 (N_9884,N_9406,N_9454);
xor U9885 (N_9885,N_9238,N_9180);
nor U9886 (N_9886,N_9335,N_9154);
nor U9887 (N_9887,N_9032,N_9404);
nand U9888 (N_9888,N_9132,N_9386);
nand U9889 (N_9889,N_9424,N_9328);
nand U9890 (N_9890,N_9291,N_9140);
and U9891 (N_9891,N_9117,N_9161);
or U9892 (N_9892,N_9382,N_9461);
xnor U9893 (N_9893,N_9008,N_9396);
nand U9894 (N_9894,N_9164,N_9410);
nor U9895 (N_9895,N_9385,N_9244);
and U9896 (N_9896,N_9181,N_9196);
or U9897 (N_9897,N_9282,N_9000);
nor U9898 (N_9898,N_9474,N_9389);
nand U9899 (N_9899,N_9024,N_9394);
nor U9900 (N_9900,N_9034,N_9434);
nand U9901 (N_9901,N_9038,N_9136);
xnor U9902 (N_9902,N_9413,N_9169);
nor U9903 (N_9903,N_9033,N_9499);
xnor U9904 (N_9904,N_9454,N_9404);
xor U9905 (N_9905,N_9082,N_9160);
and U9906 (N_9906,N_9229,N_9186);
and U9907 (N_9907,N_9336,N_9238);
or U9908 (N_9908,N_9179,N_9147);
or U9909 (N_9909,N_9260,N_9392);
and U9910 (N_9910,N_9042,N_9041);
nand U9911 (N_9911,N_9271,N_9304);
xnor U9912 (N_9912,N_9475,N_9024);
nor U9913 (N_9913,N_9201,N_9394);
nor U9914 (N_9914,N_9068,N_9316);
or U9915 (N_9915,N_9139,N_9480);
and U9916 (N_9916,N_9427,N_9203);
or U9917 (N_9917,N_9337,N_9076);
and U9918 (N_9918,N_9232,N_9170);
nor U9919 (N_9919,N_9188,N_9458);
and U9920 (N_9920,N_9046,N_9032);
nor U9921 (N_9921,N_9262,N_9291);
nand U9922 (N_9922,N_9392,N_9082);
nand U9923 (N_9923,N_9061,N_9397);
nand U9924 (N_9924,N_9289,N_9193);
or U9925 (N_9925,N_9103,N_9342);
nor U9926 (N_9926,N_9287,N_9040);
and U9927 (N_9927,N_9106,N_9357);
and U9928 (N_9928,N_9219,N_9303);
and U9929 (N_9929,N_9035,N_9490);
nand U9930 (N_9930,N_9413,N_9339);
nor U9931 (N_9931,N_9364,N_9421);
nor U9932 (N_9932,N_9386,N_9052);
xor U9933 (N_9933,N_9310,N_9180);
or U9934 (N_9934,N_9195,N_9088);
and U9935 (N_9935,N_9475,N_9274);
nand U9936 (N_9936,N_9256,N_9316);
xnor U9937 (N_9937,N_9006,N_9057);
and U9938 (N_9938,N_9395,N_9317);
nor U9939 (N_9939,N_9021,N_9354);
and U9940 (N_9940,N_9352,N_9182);
nand U9941 (N_9941,N_9144,N_9167);
and U9942 (N_9942,N_9317,N_9377);
nand U9943 (N_9943,N_9429,N_9190);
xor U9944 (N_9944,N_9389,N_9394);
nor U9945 (N_9945,N_9375,N_9480);
nor U9946 (N_9946,N_9286,N_9395);
or U9947 (N_9947,N_9175,N_9050);
nor U9948 (N_9948,N_9041,N_9437);
nand U9949 (N_9949,N_9498,N_9178);
or U9950 (N_9950,N_9235,N_9420);
nand U9951 (N_9951,N_9415,N_9305);
and U9952 (N_9952,N_9256,N_9057);
nor U9953 (N_9953,N_9415,N_9172);
or U9954 (N_9954,N_9213,N_9015);
and U9955 (N_9955,N_9049,N_9371);
nor U9956 (N_9956,N_9137,N_9301);
xnor U9957 (N_9957,N_9096,N_9136);
nand U9958 (N_9958,N_9357,N_9337);
and U9959 (N_9959,N_9459,N_9488);
or U9960 (N_9960,N_9091,N_9478);
nor U9961 (N_9961,N_9212,N_9488);
or U9962 (N_9962,N_9293,N_9182);
nand U9963 (N_9963,N_9377,N_9463);
and U9964 (N_9964,N_9179,N_9237);
nor U9965 (N_9965,N_9346,N_9474);
or U9966 (N_9966,N_9043,N_9192);
nor U9967 (N_9967,N_9086,N_9236);
nand U9968 (N_9968,N_9119,N_9295);
or U9969 (N_9969,N_9232,N_9045);
and U9970 (N_9970,N_9281,N_9222);
and U9971 (N_9971,N_9443,N_9430);
or U9972 (N_9972,N_9266,N_9168);
or U9973 (N_9973,N_9238,N_9452);
nor U9974 (N_9974,N_9027,N_9120);
or U9975 (N_9975,N_9347,N_9428);
and U9976 (N_9976,N_9453,N_9006);
and U9977 (N_9977,N_9297,N_9050);
nand U9978 (N_9978,N_9115,N_9078);
nand U9979 (N_9979,N_9294,N_9073);
or U9980 (N_9980,N_9425,N_9272);
nor U9981 (N_9981,N_9456,N_9200);
nand U9982 (N_9982,N_9191,N_9305);
and U9983 (N_9983,N_9366,N_9426);
or U9984 (N_9984,N_9326,N_9183);
nand U9985 (N_9985,N_9156,N_9497);
and U9986 (N_9986,N_9194,N_9337);
nand U9987 (N_9987,N_9229,N_9347);
xnor U9988 (N_9988,N_9024,N_9000);
or U9989 (N_9989,N_9359,N_9432);
nand U9990 (N_9990,N_9439,N_9269);
nor U9991 (N_9991,N_9257,N_9448);
nor U9992 (N_9992,N_9382,N_9488);
nand U9993 (N_9993,N_9439,N_9180);
nor U9994 (N_9994,N_9105,N_9223);
nand U9995 (N_9995,N_9346,N_9023);
nor U9996 (N_9996,N_9177,N_9321);
xnor U9997 (N_9997,N_9094,N_9262);
and U9998 (N_9998,N_9088,N_9129);
and U9999 (N_9999,N_9213,N_9459);
and UO_0 (O_0,N_9854,N_9811);
nand UO_1 (O_1,N_9529,N_9765);
xor UO_2 (O_2,N_9527,N_9972);
nor UO_3 (O_3,N_9718,N_9986);
and UO_4 (O_4,N_9513,N_9514);
nor UO_5 (O_5,N_9767,N_9993);
and UO_6 (O_6,N_9917,N_9611);
or UO_7 (O_7,N_9868,N_9659);
or UO_8 (O_8,N_9915,N_9542);
nand UO_9 (O_9,N_9627,N_9769);
nand UO_10 (O_10,N_9825,N_9980);
nor UO_11 (O_11,N_9601,N_9537);
xnor UO_12 (O_12,N_9755,N_9961);
or UO_13 (O_13,N_9969,N_9760);
nand UO_14 (O_14,N_9728,N_9736);
or UO_15 (O_15,N_9598,N_9776);
nor UO_16 (O_16,N_9931,N_9691);
or UO_17 (O_17,N_9948,N_9852);
nor UO_18 (O_18,N_9684,N_9914);
nor UO_19 (O_19,N_9748,N_9875);
xnor UO_20 (O_20,N_9906,N_9511);
and UO_21 (O_21,N_9833,N_9701);
nand UO_22 (O_22,N_9730,N_9562);
nand UO_23 (O_23,N_9928,N_9884);
or UO_24 (O_24,N_9871,N_9580);
and UO_25 (O_25,N_9773,N_9757);
nor UO_26 (O_26,N_9965,N_9665);
or UO_27 (O_27,N_9662,N_9711);
nor UO_28 (O_28,N_9652,N_9922);
xor UO_29 (O_29,N_9716,N_9680);
xnor UO_30 (O_30,N_9509,N_9717);
nor UO_31 (O_31,N_9644,N_9824);
nor UO_32 (O_32,N_9524,N_9878);
nor UO_33 (O_33,N_9747,N_9621);
xnor UO_34 (O_34,N_9532,N_9837);
xnor UO_35 (O_35,N_9912,N_9698);
nand UO_36 (O_36,N_9819,N_9975);
nor UO_37 (O_37,N_9528,N_9626);
and UO_38 (O_38,N_9913,N_9813);
and UO_39 (O_39,N_9639,N_9669);
nand UO_40 (O_40,N_9733,N_9779);
or UO_41 (O_41,N_9602,N_9821);
and UO_42 (O_42,N_9688,N_9617);
or UO_43 (O_43,N_9749,N_9789);
nand UO_44 (O_44,N_9849,N_9800);
xnor UO_45 (O_45,N_9879,N_9804);
xnor UO_46 (O_46,N_9681,N_9941);
and UO_47 (O_47,N_9771,N_9904);
nand UO_48 (O_48,N_9561,N_9866);
nand UO_49 (O_49,N_9628,N_9766);
and UO_50 (O_50,N_9835,N_9959);
nand UO_51 (O_51,N_9907,N_9918);
or UO_52 (O_52,N_9889,N_9794);
nand UO_53 (O_53,N_9859,N_9775);
nand UO_54 (O_54,N_9533,N_9584);
and UO_55 (O_55,N_9505,N_9786);
nand UO_56 (O_56,N_9905,N_9982);
nor UO_57 (O_57,N_9520,N_9696);
nor UO_58 (O_58,N_9805,N_9809);
and UO_59 (O_59,N_9739,N_9838);
xnor UO_60 (O_60,N_9929,N_9890);
or UO_61 (O_61,N_9792,N_9512);
nand UO_62 (O_62,N_9892,N_9839);
or UO_63 (O_63,N_9958,N_9936);
nor UO_64 (O_64,N_9842,N_9585);
xnor UO_65 (O_65,N_9802,N_9785);
nor UO_66 (O_66,N_9899,N_9850);
and UO_67 (O_67,N_9615,N_9977);
and UO_68 (O_68,N_9950,N_9731);
or UO_69 (O_69,N_9783,N_9501);
xnor UO_70 (O_70,N_9937,N_9604);
nand UO_71 (O_71,N_9575,N_9699);
nor UO_72 (O_72,N_9844,N_9920);
and UO_73 (O_73,N_9857,N_9847);
or UO_74 (O_74,N_9654,N_9940);
nor UO_75 (O_75,N_9843,N_9964);
nor UO_76 (O_76,N_9740,N_9943);
or UO_77 (O_77,N_9548,N_9553);
xnor UO_78 (O_78,N_9591,N_9634);
or UO_79 (O_79,N_9933,N_9953);
nor UO_80 (O_80,N_9797,N_9796);
and UO_81 (O_81,N_9582,N_9834);
nand UO_82 (O_82,N_9620,N_9944);
nor UO_83 (O_83,N_9810,N_9795);
or UO_84 (O_84,N_9687,N_9721);
nor UO_85 (O_85,N_9791,N_9600);
and UO_86 (O_86,N_9506,N_9567);
and UO_87 (O_87,N_9947,N_9761);
or UO_88 (O_88,N_9738,N_9778);
xnor UO_89 (O_89,N_9873,N_9863);
nor UO_90 (O_90,N_9571,N_9517);
or UO_91 (O_91,N_9596,N_9777);
nor UO_92 (O_92,N_9876,N_9710);
and UO_93 (O_93,N_9935,N_9645);
and UO_94 (O_94,N_9559,N_9581);
and UO_95 (O_95,N_9881,N_9885);
nor UO_96 (O_96,N_9586,N_9994);
nand UO_97 (O_97,N_9543,N_9675);
or UO_98 (O_98,N_9784,N_9754);
nor UO_99 (O_99,N_9660,N_9702);
nand UO_100 (O_100,N_9763,N_9525);
or UO_101 (O_101,N_9573,N_9829);
xor UO_102 (O_102,N_9606,N_9832);
xnor UO_103 (O_103,N_9820,N_9744);
nand UO_104 (O_104,N_9891,N_9633);
or UO_105 (O_105,N_9724,N_9945);
xnor UO_106 (O_106,N_9607,N_9894);
nor UO_107 (O_107,N_9672,N_9510);
nor UO_108 (O_108,N_9707,N_9949);
nor UO_109 (O_109,N_9787,N_9996);
nor UO_110 (O_110,N_9897,N_9973);
nor UO_111 (O_111,N_9729,N_9605);
xnor UO_112 (O_112,N_9822,N_9998);
or UO_113 (O_113,N_9921,N_9690);
nor UO_114 (O_114,N_9614,N_9540);
and UO_115 (O_115,N_9869,N_9807);
and UO_116 (O_116,N_9656,N_9901);
or UO_117 (O_117,N_9706,N_9723);
or UO_118 (O_118,N_9874,N_9910);
nand UO_119 (O_119,N_9923,N_9756);
or UO_120 (O_120,N_9530,N_9911);
nor UO_121 (O_121,N_9693,N_9828);
or UO_122 (O_122,N_9741,N_9700);
nand UO_123 (O_123,N_9768,N_9909);
and UO_124 (O_124,N_9815,N_9742);
nand UO_125 (O_125,N_9546,N_9694);
and UO_126 (O_126,N_9570,N_9704);
nor UO_127 (O_127,N_9919,N_9841);
and UO_128 (O_128,N_9732,N_9535);
nand UO_129 (O_129,N_9872,N_9951);
or UO_130 (O_130,N_9599,N_9563);
or UO_131 (O_131,N_9708,N_9623);
or UO_132 (O_132,N_9870,N_9595);
or UO_133 (O_133,N_9927,N_9709);
nor UO_134 (O_134,N_9984,N_9649);
or UO_135 (O_135,N_9974,N_9774);
nor UO_136 (O_136,N_9727,N_9853);
nor UO_137 (O_137,N_9764,N_9893);
or UO_138 (O_138,N_9719,N_9572);
nand UO_139 (O_139,N_9564,N_9858);
and UO_140 (O_140,N_9619,N_9737);
nand UO_141 (O_141,N_9641,N_9930);
or UO_142 (O_142,N_9577,N_9938);
nor UO_143 (O_143,N_9753,N_9968);
or UO_144 (O_144,N_9677,N_9772);
nand UO_145 (O_145,N_9806,N_9569);
or UO_146 (O_146,N_9855,N_9579);
or UO_147 (O_147,N_9657,N_9647);
nand UO_148 (O_148,N_9550,N_9713);
nor UO_149 (O_149,N_9799,N_9743);
or UO_150 (O_150,N_9593,N_9712);
and UO_151 (O_151,N_9664,N_9552);
xor UO_152 (O_152,N_9685,N_9587);
and UO_153 (O_153,N_9538,N_9515);
or UO_154 (O_154,N_9612,N_9782);
nand UO_155 (O_155,N_9545,N_9608);
nand UO_156 (O_156,N_9999,N_9566);
nand UO_157 (O_157,N_9865,N_9589);
nand UO_158 (O_158,N_9817,N_9518);
nand UO_159 (O_159,N_9750,N_9848);
nand UO_160 (O_160,N_9745,N_9934);
xnor UO_161 (O_161,N_9955,N_9597);
nor UO_162 (O_162,N_9500,N_9836);
and UO_163 (O_163,N_9565,N_9823);
or UO_164 (O_164,N_9642,N_9674);
nand UO_165 (O_165,N_9671,N_9678);
xnor UO_166 (O_166,N_9703,N_9502);
xnor UO_167 (O_167,N_9908,N_9650);
or UO_168 (O_168,N_9618,N_9803);
and UO_169 (O_169,N_9661,N_9578);
nor UO_170 (O_170,N_9722,N_9970);
nand UO_171 (O_171,N_9705,N_9646);
nor UO_172 (O_172,N_9735,N_9673);
and UO_173 (O_173,N_9840,N_9900);
and UO_174 (O_174,N_9963,N_9523);
nand UO_175 (O_175,N_9883,N_9668);
nor UO_176 (O_176,N_9504,N_9946);
nor UO_177 (O_177,N_9638,N_9983);
xor UO_178 (O_178,N_9594,N_9629);
nand UO_179 (O_179,N_9846,N_9603);
nor UO_180 (O_180,N_9534,N_9882);
or UO_181 (O_181,N_9676,N_9588);
nor UO_182 (O_182,N_9536,N_9898);
and UO_183 (O_183,N_9568,N_9845);
nor UO_184 (O_184,N_9616,N_9888);
nor UO_185 (O_185,N_9544,N_9679);
nor UO_186 (O_186,N_9516,N_9507);
nor UO_187 (O_187,N_9653,N_9555);
nor UO_188 (O_188,N_9924,N_9957);
and UO_189 (O_189,N_9814,N_9793);
or UO_190 (O_190,N_9610,N_9720);
nand UO_191 (O_191,N_9895,N_9864);
nor UO_192 (O_192,N_9631,N_9503);
nor UO_193 (O_193,N_9670,N_9549);
nor UO_194 (O_194,N_9637,N_9609);
or UO_195 (O_195,N_9560,N_9658);
and UO_196 (O_196,N_9808,N_9997);
nand UO_197 (O_197,N_9992,N_9902);
nand UO_198 (O_198,N_9925,N_9655);
or UO_199 (O_199,N_9683,N_9886);
xor UO_200 (O_200,N_9861,N_9667);
nand UO_201 (O_201,N_9826,N_9976);
nor UO_202 (O_202,N_9812,N_9887);
or UO_203 (O_203,N_9867,N_9989);
and UO_204 (O_204,N_9695,N_9962);
or UO_205 (O_205,N_9522,N_9583);
xnor UO_206 (O_206,N_9877,N_9971);
and UO_207 (O_207,N_9926,N_9827);
nor UO_208 (O_208,N_9952,N_9551);
xnor UO_209 (O_209,N_9860,N_9954);
nor UO_210 (O_210,N_9798,N_9625);
nand UO_211 (O_211,N_9526,N_9682);
nor UO_212 (O_212,N_9635,N_9942);
and UO_213 (O_213,N_9995,N_9788);
and UO_214 (O_214,N_9666,N_9818);
nand UO_215 (O_215,N_9547,N_9541);
nor UO_216 (O_216,N_9896,N_9960);
nand UO_217 (O_217,N_9851,N_9903);
and UO_218 (O_218,N_9770,N_9715);
nor UO_219 (O_219,N_9640,N_9758);
nand UO_220 (O_220,N_9988,N_9880);
and UO_221 (O_221,N_9558,N_9726);
or UO_222 (O_222,N_9987,N_9990);
nand UO_223 (O_223,N_9801,N_9816);
nand UO_224 (O_224,N_9966,N_9734);
nand UO_225 (O_225,N_9648,N_9556);
nand UO_226 (O_226,N_9978,N_9697);
or UO_227 (O_227,N_9636,N_9630);
nor UO_228 (O_228,N_9686,N_9780);
or UO_229 (O_229,N_9508,N_9956);
nor UO_230 (O_230,N_9651,N_9916);
xnor UO_231 (O_231,N_9531,N_9762);
or UO_232 (O_232,N_9554,N_9752);
or UO_233 (O_233,N_9692,N_9939);
nand UO_234 (O_234,N_9751,N_9521);
and UO_235 (O_235,N_9624,N_9725);
nor UO_236 (O_236,N_9622,N_9985);
xor UO_237 (O_237,N_9539,N_9663);
and UO_238 (O_238,N_9576,N_9714);
xnor UO_239 (O_239,N_9981,N_9979);
or UO_240 (O_240,N_9519,N_9831);
and UO_241 (O_241,N_9759,N_9932);
nor UO_242 (O_242,N_9790,N_9613);
nand UO_243 (O_243,N_9746,N_9574);
or UO_244 (O_244,N_9689,N_9592);
nand UO_245 (O_245,N_9830,N_9632);
nor UO_246 (O_246,N_9862,N_9967);
nor UO_247 (O_247,N_9781,N_9643);
nand UO_248 (O_248,N_9557,N_9856);
and UO_249 (O_249,N_9590,N_9991);
and UO_250 (O_250,N_9872,N_9843);
nor UO_251 (O_251,N_9786,N_9845);
and UO_252 (O_252,N_9917,N_9584);
nand UO_253 (O_253,N_9581,N_9509);
or UO_254 (O_254,N_9513,N_9534);
or UO_255 (O_255,N_9761,N_9603);
nand UO_256 (O_256,N_9676,N_9544);
or UO_257 (O_257,N_9565,N_9637);
or UO_258 (O_258,N_9805,N_9734);
nor UO_259 (O_259,N_9906,N_9686);
nand UO_260 (O_260,N_9739,N_9598);
nor UO_261 (O_261,N_9781,N_9548);
xnor UO_262 (O_262,N_9649,N_9547);
nor UO_263 (O_263,N_9583,N_9638);
xor UO_264 (O_264,N_9542,N_9619);
nor UO_265 (O_265,N_9935,N_9523);
nand UO_266 (O_266,N_9735,N_9881);
nor UO_267 (O_267,N_9971,N_9777);
and UO_268 (O_268,N_9969,N_9521);
nor UO_269 (O_269,N_9795,N_9674);
xnor UO_270 (O_270,N_9514,N_9918);
nor UO_271 (O_271,N_9962,N_9936);
nand UO_272 (O_272,N_9935,N_9679);
and UO_273 (O_273,N_9801,N_9877);
or UO_274 (O_274,N_9872,N_9966);
and UO_275 (O_275,N_9866,N_9974);
or UO_276 (O_276,N_9726,N_9683);
nand UO_277 (O_277,N_9962,N_9980);
nor UO_278 (O_278,N_9894,N_9846);
or UO_279 (O_279,N_9983,N_9596);
xor UO_280 (O_280,N_9665,N_9597);
and UO_281 (O_281,N_9762,N_9577);
or UO_282 (O_282,N_9542,N_9830);
nand UO_283 (O_283,N_9821,N_9500);
nand UO_284 (O_284,N_9508,N_9942);
and UO_285 (O_285,N_9969,N_9954);
or UO_286 (O_286,N_9861,N_9755);
or UO_287 (O_287,N_9789,N_9760);
nand UO_288 (O_288,N_9562,N_9847);
xor UO_289 (O_289,N_9684,N_9582);
nor UO_290 (O_290,N_9768,N_9523);
and UO_291 (O_291,N_9773,N_9917);
or UO_292 (O_292,N_9506,N_9825);
xnor UO_293 (O_293,N_9874,N_9517);
nor UO_294 (O_294,N_9685,N_9769);
nand UO_295 (O_295,N_9918,N_9603);
nand UO_296 (O_296,N_9727,N_9550);
nand UO_297 (O_297,N_9846,N_9670);
nand UO_298 (O_298,N_9939,N_9569);
nand UO_299 (O_299,N_9608,N_9942);
nor UO_300 (O_300,N_9990,N_9528);
or UO_301 (O_301,N_9544,N_9828);
or UO_302 (O_302,N_9803,N_9802);
and UO_303 (O_303,N_9796,N_9598);
xnor UO_304 (O_304,N_9686,N_9764);
nand UO_305 (O_305,N_9711,N_9822);
nand UO_306 (O_306,N_9647,N_9723);
and UO_307 (O_307,N_9782,N_9711);
or UO_308 (O_308,N_9521,N_9813);
nor UO_309 (O_309,N_9797,N_9533);
xnor UO_310 (O_310,N_9688,N_9891);
and UO_311 (O_311,N_9841,N_9685);
nor UO_312 (O_312,N_9984,N_9715);
or UO_313 (O_313,N_9531,N_9765);
and UO_314 (O_314,N_9800,N_9770);
nand UO_315 (O_315,N_9857,N_9900);
nor UO_316 (O_316,N_9563,N_9607);
and UO_317 (O_317,N_9873,N_9835);
nor UO_318 (O_318,N_9999,N_9835);
nor UO_319 (O_319,N_9956,N_9812);
nand UO_320 (O_320,N_9837,N_9738);
and UO_321 (O_321,N_9572,N_9838);
nand UO_322 (O_322,N_9820,N_9748);
or UO_323 (O_323,N_9974,N_9837);
nor UO_324 (O_324,N_9521,N_9914);
or UO_325 (O_325,N_9715,N_9917);
or UO_326 (O_326,N_9930,N_9823);
and UO_327 (O_327,N_9729,N_9698);
nand UO_328 (O_328,N_9898,N_9776);
nand UO_329 (O_329,N_9936,N_9808);
xnor UO_330 (O_330,N_9828,N_9636);
and UO_331 (O_331,N_9909,N_9567);
or UO_332 (O_332,N_9539,N_9612);
nor UO_333 (O_333,N_9990,N_9543);
nand UO_334 (O_334,N_9722,N_9797);
nand UO_335 (O_335,N_9914,N_9908);
nor UO_336 (O_336,N_9671,N_9593);
and UO_337 (O_337,N_9963,N_9611);
or UO_338 (O_338,N_9547,N_9977);
or UO_339 (O_339,N_9741,N_9691);
and UO_340 (O_340,N_9743,N_9787);
or UO_341 (O_341,N_9703,N_9713);
nor UO_342 (O_342,N_9659,N_9514);
and UO_343 (O_343,N_9723,N_9915);
nand UO_344 (O_344,N_9768,N_9839);
nor UO_345 (O_345,N_9729,N_9897);
or UO_346 (O_346,N_9937,N_9984);
xor UO_347 (O_347,N_9651,N_9548);
nand UO_348 (O_348,N_9727,N_9611);
or UO_349 (O_349,N_9914,N_9714);
nor UO_350 (O_350,N_9627,N_9539);
nor UO_351 (O_351,N_9937,N_9753);
or UO_352 (O_352,N_9594,N_9563);
or UO_353 (O_353,N_9985,N_9884);
or UO_354 (O_354,N_9536,N_9623);
and UO_355 (O_355,N_9651,N_9928);
nand UO_356 (O_356,N_9906,N_9702);
or UO_357 (O_357,N_9812,N_9896);
nor UO_358 (O_358,N_9651,N_9924);
and UO_359 (O_359,N_9542,N_9812);
or UO_360 (O_360,N_9772,N_9703);
nor UO_361 (O_361,N_9895,N_9962);
or UO_362 (O_362,N_9928,N_9712);
xor UO_363 (O_363,N_9588,N_9852);
nand UO_364 (O_364,N_9716,N_9727);
nor UO_365 (O_365,N_9615,N_9590);
nand UO_366 (O_366,N_9715,N_9987);
nand UO_367 (O_367,N_9861,N_9876);
and UO_368 (O_368,N_9820,N_9758);
xor UO_369 (O_369,N_9567,N_9711);
nor UO_370 (O_370,N_9911,N_9512);
nor UO_371 (O_371,N_9734,N_9842);
xnor UO_372 (O_372,N_9509,N_9512);
nor UO_373 (O_373,N_9643,N_9921);
and UO_374 (O_374,N_9839,N_9646);
or UO_375 (O_375,N_9743,N_9981);
or UO_376 (O_376,N_9629,N_9595);
nand UO_377 (O_377,N_9893,N_9580);
nand UO_378 (O_378,N_9870,N_9881);
and UO_379 (O_379,N_9990,N_9680);
or UO_380 (O_380,N_9612,N_9538);
or UO_381 (O_381,N_9646,N_9735);
and UO_382 (O_382,N_9637,N_9589);
or UO_383 (O_383,N_9844,N_9753);
nand UO_384 (O_384,N_9523,N_9649);
nand UO_385 (O_385,N_9879,N_9848);
nor UO_386 (O_386,N_9881,N_9971);
nand UO_387 (O_387,N_9913,N_9602);
and UO_388 (O_388,N_9621,N_9983);
and UO_389 (O_389,N_9672,N_9830);
nand UO_390 (O_390,N_9706,N_9898);
and UO_391 (O_391,N_9984,N_9979);
nand UO_392 (O_392,N_9672,N_9667);
or UO_393 (O_393,N_9610,N_9911);
and UO_394 (O_394,N_9729,N_9730);
xor UO_395 (O_395,N_9566,N_9604);
or UO_396 (O_396,N_9897,N_9824);
and UO_397 (O_397,N_9617,N_9785);
or UO_398 (O_398,N_9675,N_9604);
and UO_399 (O_399,N_9668,N_9764);
nor UO_400 (O_400,N_9691,N_9730);
nor UO_401 (O_401,N_9839,N_9696);
nand UO_402 (O_402,N_9753,N_9729);
or UO_403 (O_403,N_9925,N_9540);
nand UO_404 (O_404,N_9527,N_9963);
or UO_405 (O_405,N_9768,N_9781);
or UO_406 (O_406,N_9767,N_9722);
nor UO_407 (O_407,N_9866,N_9548);
or UO_408 (O_408,N_9909,N_9791);
nor UO_409 (O_409,N_9601,N_9904);
nand UO_410 (O_410,N_9520,N_9651);
nand UO_411 (O_411,N_9985,N_9692);
nor UO_412 (O_412,N_9540,N_9558);
and UO_413 (O_413,N_9835,N_9920);
or UO_414 (O_414,N_9557,N_9560);
nand UO_415 (O_415,N_9965,N_9964);
nor UO_416 (O_416,N_9580,N_9761);
xnor UO_417 (O_417,N_9583,N_9575);
nor UO_418 (O_418,N_9708,N_9874);
nand UO_419 (O_419,N_9767,N_9966);
nor UO_420 (O_420,N_9635,N_9569);
nor UO_421 (O_421,N_9825,N_9860);
nor UO_422 (O_422,N_9934,N_9685);
and UO_423 (O_423,N_9651,N_9799);
nor UO_424 (O_424,N_9628,N_9824);
xor UO_425 (O_425,N_9606,N_9644);
and UO_426 (O_426,N_9904,N_9909);
or UO_427 (O_427,N_9780,N_9931);
nand UO_428 (O_428,N_9766,N_9526);
nand UO_429 (O_429,N_9544,N_9682);
nand UO_430 (O_430,N_9902,N_9834);
nor UO_431 (O_431,N_9876,N_9647);
and UO_432 (O_432,N_9953,N_9536);
nor UO_433 (O_433,N_9512,N_9717);
nor UO_434 (O_434,N_9984,N_9952);
nor UO_435 (O_435,N_9885,N_9988);
nand UO_436 (O_436,N_9799,N_9899);
nor UO_437 (O_437,N_9556,N_9702);
and UO_438 (O_438,N_9870,N_9761);
or UO_439 (O_439,N_9634,N_9560);
nor UO_440 (O_440,N_9709,N_9801);
nand UO_441 (O_441,N_9876,N_9911);
and UO_442 (O_442,N_9929,N_9685);
nor UO_443 (O_443,N_9833,N_9915);
or UO_444 (O_444,N_9850,N_9517);
nor UO_445 (O_445,N_9846,N_9659);
and UO_446 (O_446,N_9777,N_9802);
nor UO_447 (O_447,N_9987,N_9797);
nand UO_448 (O_448,N_9554,N_9687);
or UO_449 (O_449,N_9940,N_9794);
or UO_450 (O_450,N_9550,N_9641);
and UO_451 (O_451,N_9816,N_9706);
nand UO_452 (O_452,N_9983,N_9922);
nor UO_453 (O_453,N_9874,N_9516);
or UO_454 (O_454,N_9719,N_9981);
xor UO_455 (O_455,N_9542,N_9864);
or UO_456 (O_456,N_9750,N_9516);
and UO_457 (O_457,N_9703,N_9807);
nor UO_458 (O_458,N_9639,N_9757);
and UO_459 (O_459,N_9911,N_9537);
and UO_460 (O_460,N_9617,N_9552);
xnor UO_461 (O_461,N_9977,N_9855);
or UO_462 (O_462,N_9742,N_9611);
and UO_463 (O_463,N_9618,N_9890);
or UO_464 (O_464,N_9757,N_9874);
nand UO_465 (O_465,N_9542,N_9687);
or UO_466 (O_466,N_9930,N_9776);
and UO_467 (O_467,N_9684,N_9740);
and UO_468 (O_468,N_9950,N_9849);
nor UO_469 (O_469,N_9712,N_9843);
nand UO_470 (O_470,N_9957,N_9962);
or UO_471 (O_471,N_9805,N_9991);
or UO_472 (O_472,N_9992,N_9551);
nor UO_473 (O_473,N_9808,N_9801);
or UO_474 (O_474,N_9634,N_9703);
nor UO_475 (O_475,N_9602,N_9723);
nor UO_476 (O_476,N_9952,N_9808);
xor UO_477 (O_477,N_9559,N_9675);
and UO_478 (O_478,N_9744,N_9784);
and UO_479 (O_479,N_9821,N_9805);
nor UO_480 (O_480,N_9568,N_9933);
nand UO_481 (O_481,N_9506,N_9822);
xor UO_482 (O_482,N_9901,N_9924);
xor UO_483 (O_483,N_9593,N_9937);
or UO_484 (O_484,N_9876,N_9624);
and UO_485 (O_485,N_9924,N_9577);
nor UO_486 (O_486,N_9634,N_9743);
xor UO_487 (O_487,N_9597,N_9849);
nand UO_488 (O_488,N_9588,N_9656);
xor UO_489 (O_489,N_9797,N_9827);
nor UO_490 (O_490,N_9650,N_9881);
nand UO_491 (O_491,N_9922,N_9821);
nand UO_492 (O_492,N_9846,N_9868);
nor UO_493 (O_493,N_9768,N_9899);
nand UO_494 (O_494,N_9762,N_9570);
and UO_495 (O_495,N_9647,N_9945);
nand UO_496 (O_496,N_9546,N_9659);
or UO_497 (O_497,N_9635,N_9768);
xor UO_498 (O_498,N_9535,N_9658);
nand UO_499 (O_499,N_9929,N_9719);
and UO_500 (O_500,N_9634,N_9981);
or UO_501 (O_501,N_9757,N_9977);
or UO_502 (O_502,N_9733,N_9739);
and UO_503 (O_503,N_9784,N_9730);
xnor UO_504 (O_504,N_9507,N_9759);
nand UO_505 (O_505,N_9677,N_9798);
nand UO_506 (O_506,N_9885,N_9992);
and UO_507 (O_507,N_9785,N_9912);
xnor UO_508 (O_508,N_9748,N_9539);
or UO_509 (O_509,N_9650,N_9598);
nand UO_510 (O_510,N_9766,N_9943);
nor UO_511 (O_511,N_9579,N_9558);
nor UO_512 (O_512,N_9597,N_9667);
nand UO_513 (O_513,N_9556,N_9809);
nand UO_514 (O_514,N_9891,N_9715);
nand UO_515 (O_515,N_9710,N_9530);
and UO_516 (O_516,N_9887,N_9633);
and UO_517 (O_517,N_9957,N_9665);
or UO_518 (O_518,N_9777,N_9922);
xor UO_519 (O_519,N_9606,N_9699);
and UO_520 (O_520,N_9705,N_9547);
or UO_521 (O_521,N_9806,N_9666);
nor UO_522 (O_522,N_9570,N_9562);
xor UO_523 (O_523,N_9923,N_9857);
or UO_524 (O_524,N_9564,N_9713);
or UO_525 (O_525,N_9692,N_9781);
nand UO_526 (O_526,N_9551,N_9927);
nand UO_527 (O_527,N_9964,N_9818);
nand UO_528 (O_528,N_9965,N_9704);
or UO_529 (O_529,N_9895,N_9989);
or UO_530 (O_530,N_9567,N_9991);
nand UO_531 (O_531,N_9989,N_9939);
nor UO_532 (O_532,N_9932,N_9746);
and UO_533 (O_533,N_9821,N_9702);
nor UO_534 (O_534,N_9658,N_9525);
or UO_535 (O_535,N_9904,N_9608);
nand UO_536 (O_536,N_9903,N_9718);
or UO_537 (O_537,N_9811,N_9756);
nor UO_538 (O_538,N_9796,N_9503);
and UO_539 (O_539,N_9883,N_9617);
and UO_540 (O_540,N_9588,N_9936);
nand UO_541 (O_541,N_9800,N_9960);
and UO_542 (O_542,N_9647,N_9673);
nand UO_543 (O_543,N_9525,N_9904);
nand UO_544 (O_544,N_9515,N_9742);
nand UO_545 (O_545,N_9906,N_9606);
and UO_546 (O_546,N_9777,N_9973);
nand UO_547 (O_547,N_9525,N_9771);
nand UO_548 (O_548,N_9880,N_9783);
xor UO_549 (O_549,N_9947,N_9543);
xnor UO_550 (O_550,N_9904,N_9760);
or UO_551 (O_551,N_9881,N_9872);
nor UO_552 (O_552,N_9792,N_9606);
nand UO_553 (O_553,N_9688,N_9938);
or UO_554 (O_554,N_9772,N_9879);
or UO_555 (O_555,N_9956,N_9832);
nor UO_556 (O_556,N_9947,N_9918);
and UO_557 (O_557,N_9904,N_9690);
or UO_558 (O_558,N_9728,N_9910);
xor UO_559 (O_559,N_9851,N_9622);
and UO_560 (O_560,N_9921,N_9682);
and UO_561 (O_561,N_9571,N_9958);
or UO_562 (O_562,N_9719,N_9973);
nor UO_563 (O_563,N_9586,N_9802);
nor UO_564 (O_564,N_9798,N_9678);
nand UO_565 (O_565,N_9839,N_9562);
xor UO_566 (O_566,N_9978,N_9806);
and UO_567 (O_567,N_9648,N_9789);
or UO_568 (O_568,N_9504,N_9630);
or UO_569 (O_569,N_9753,N_9727);
or UO_570 (O_570,N_9866,N_9579);
nor UO_571 (O_571,N_9951,N_9717);
or UO_572 (O_572,N_9653,N_9800);
nand UO_573 (O_573,N_9656,N_9613);
and UO_574 (O_574,N_9998,N_9729);
nor UO_575 (O_575,N_9899,N_9789);
nand UO_576 (O_576,N_9965,N_9678);
nor UO_577 (O_577,N_9951,N_9531);
or UO_578 (O_578,N_9514,N_9700);
and UO_579 (O_579,N_9638,N_9565);
nor UO_580 (O_580,N_9822,N_9763);
and UO_581 (O_581,N_9887,N_9874);
nand UO_582 (O_582,N_9622,N_9912);
or UO_583 (O_583,N_9889,N_9888);
nand UO_584 (O_584,N_9615,N_9992);
and UO_585 (O_585,N_9794,N_9865);
or UO_586 (O_586,N_9807,N_9720);
nor UO_587 (O_587,N_9730,N_9896);
or UO_588 (O_588,N_9972,N_9743);
and UO_589 (O_589,N_9761,N_9514);
nor UO_590 (O_590,N_9598,N_9667);
nor UO_591 (O_591,N_9583,N_9953);
nor UO_592 (O_592,N_9527,N_9962);
and UO_593 (O_593,N_9762,N_9978);
nor UO_594 (O_594,N_9544,N_9681);
nor UO_595 (O_595,N_9712,N_9560);
or UO_596 (O_596,N_9960,N_9888);
or UO_597 (O_597,N_9934,N_9870);
nand UO_598 (O_598,N_9724,N_9851);
nor UO_599 (O_599,N_9947,N_9931);
nand UO_600 (O_600,N_9702,N_9916);
xor UO_601 (O_601,N_9885,N_9756);
nor UO_602 (O_602,N_9719,N_9891);
nand UO_603 (O_603,N_9543,N_9693);
nor UO_604 (O_604,N_9737,N_9952);
nand UO_605 (O_605,N_9732,N_9793);
or UO_606 (O_606,N_9778,N_9849);
xnor UO_607 (O_607,N_9757,N_9641);
or UO_608 (O_608,N_9520,N_9582);
nor UO_609 (O_609,N_9736,N_9793);
and UO_610 (O_610,N_9650,N_9668);
nor UO_611 (O_611,N_9880,N_9708);
nand UO_612 (O_612,N_9728,N_9902);
and UO_613 (O_613,N_9887,N_9822);
or UO_614 (O_614,N_9913,N_9903);
xor UO_615 (O_615,N_9940,N_9605);
and UO_616 (O_616,N_9555,N_9796);
nand UO_617 (O_617,N_9871,N_9724);
xor UO_618 (O_618,N_9580,N_9921);
or UO_619 (O_619,N_9590,N_9729);
nor UO_620 (O_620,N_9577,N_9878);
nand UO_621 (O_621,N_9626,N_9682);
or UO_622 (O_622,N_9860,N_9885);
and UO_623 (O_623,N_9791,N_9843);
and UO_624 (O_624,N_9508,N_9633);
nand UO_625 (O_625,N_9648,N_9700);
and UO_626 (O_626,N_9871,N_9817);
and UO_627 (O_627,N_9764,N_9895);
nand UO_628 (O_628,N_9865,N_9995);
or UO_629 (O_629,N_9700,N_9956);
or UO_630 (O_630,N_9877,N_9681);
xor UO_631 (O_631,N_9826,N_9640);
nor UO_632 (O_632,N_9926,N_9740);
and UO_633 (O_633,N_9557,N_9840);
nand UO_634 (O_634,N_9994,N_9602);
and UO_635 (O_635,N_9997,N_9604);
or UO_636 (O_636,N_9595,N_9914);
or UO_637 (O_637,N_9911,N_9894);
xnor UO_638 (O_638,N_9992,N_9820);
and UO_639 (O_639,N_9859,N_9684);
nand UO_640 (O_640,N_9863,N_9847);
xor UO_641 (O_641,N_9881,N_9565);
or UO_642 (O_642,N_9500,N_9992);
nand UO_643 (O_643,N_9644,N_9568);
nor UO_644 (O_644,N_9945,N_9605);
or UO_645 (O_645,N_9571,N_9581);
nand UO_646 (O_646,N_9998,N_9936);
nand UO_647 (O_647,N_9855,N_9908);
nor UO_648 (O_648,N_9530,N_9712);
or UO_649 (O_649,N_9948,N_9512);
and UO_650 (O_650,N_9696,N_9903);
xnor UO_651 (O_651,N_9879,N_9617);
xor UO_652 (O_652,N_9683,N_9617);
nor UO_653 (O_653,N_9525,N_9612);
nor UO_654 (O_654,N_9976,N_9951);
nor UO_655 (O_655,N_9517,N_9524);
nor UO_656 (O_656,N_9528,N_9835);
and UO_657 (O_657,N_9612,N_9887);
or UO_658 (O_658,N_9911,N_9908);
or UO_659 (O_659,N_9595,N_9657);
or UO_660 (O_660,N_9601,N_9554);
and UO_661 (O_661,N_9907,N_9597);
xor UO_662 (O_662,N_9915,N_9864);
nand UO_663 (O_663,N_9919,N_9604);
and UO_664 (O_664,N_9642,N_9713);
nor UO_665 (O_665,N_9680,N_9603);
xor UO_666 (O_666,N_9576,N_9504);
and UO_667 (O_667,N_9548,N_9813);
and UO_668 (O_668,N_9505,N_9567);
nor UO_669 (O_669,N_9817,N_9851);
and UO_670 (O_670,N_9697,N_9914);
nor UO_671 (O_671,N_9806,N_9544);
or UO_672 (O_672,N_9857,N_9611);
and UO_673 (O_673,N_9648,N_9615);
xnor UO_674 (O_674,N_9734,N_9840);
nand UO_675 (O_675,N_9917,N_9890);
or UO_676 (O_676,N_9855,N_9966);
nor UO_677 (O_677,N_9655,N_9507);
and UO_678 (O_678,N_9868,N_9546);
xor UO_679 (O_679,N_9688,N_9998);
or UO_680 (O_680,N_9832,N_9734);
and UO_681 (O_681,N_9979,N_9923);
nor UO_682 (O_682,N_9605,N_9863);
xor UO_683 (O_683,N_9735,N_9966);
xnor UO_684 (O_684,N_9786,N_9538);
nand UO_685 (O_685,N_9593,N_9889);
and UO_686 (O_686,N_9676,N_9646);
nor UO_687 (O_687,N_9815,N_9598);
xor UO_688 (O_688,N_9926,N_9578);
or UO_689 (O_689,N_9767,N_9606);
and UO_690 (O_690,N_9516,N_9959);
and UO_691 (O_691,N_9766,N_9532);
or UO_692 (O_692,N_9961,N_9847);
nor UO_693 (O_693,N_9707,N_9859);
nor UO_694 (O_694,N_9591,N_9610);
or UO_695 (O_695,N_9519,N_9816);
xor UO_696 (O_696,N_9963,N_9672);
nor UO_697 (O_697,N_9625,N_9570);
nand UO_698 (O_698,N_9558,N_9718);
nor UO_699 (O_699,N_9686,N_9579);
or UO_700 (O_700,N_9733,N_9845);
or UO_701 (O_701,N_9749,N_9771);
and UO_702 (O_702,N_9546,N_9735);
or UO_703 (O_703,N_9950,N_9683);
and UO_704 (O_704,N_9644,N_9551);
or UO_705 (O_705,N_9876,N_9890);
and UO_706 (O_706,N_9917,N_9694);
xnor UO_707 (O_707,N_9963,N_9514);
or UO_708 (O_708,N_9836,N_9977);
nand UO_709 (O_709,N_9557,N_9938);
or UO_710 (O_710,N_9878,N_9757);
nand UO_711 (O_711,N_9944,N_9772);
and UO_712 (O_712,N_9979,N_9849);
and UO_713 (O_713,N_9764,N_9542);
nor UO_714 (O_714,N_9530,N_9874);
or UO_715 (O_715,N_9760,N_9647);
nand UO_716 (O_716,N_9862,N_9988);
and UO_717 (O_717,N_9556,N_9567);
and UO_718 (O_718,N_9854,N_9550);
or UO_719 (O_719,N_9834,N_9777);
nor UO_720 (O_720,N_9994,N_9639);
or UO_721 (O_721,N_9693,N_9585);
nor UO_722 (O_722,N_9568,N_9922);
or UO_723 (O_723,N_9855,N_9988);
or UO_724 (O_724,N_9597,N_9970);
and UO_725 (O_725,N_9880,N_9678);
nand UO_726 (O_726,N_9934,N_9640);
nand UO_727 (O_727,N_9774,N_9650);
or UO_728 (O_728,N_9959,N_9751);
nor UO_729 (O_729,N_9512,N_9878);
xor UO_730 (O_730,N_9859,N_9955);
nand UO_731 (O_731,N_9837,N_9590);
nor UO_732 (O_732,N_9995,N_9561);
nor UO_733 (O_733,N_9978,N_9942);
nor UO_734 (O_734,N_9649,N_9514);
nand UO_735 (O_735,N_9767,N_9975);
nor UO_736 (O_736,N_9586,N_9819);
or UO_737 (O_737,N_9989,N_9778);
or UO_738 (O_738,N_9649,N_9797);
nand UO_739 (O_739,N_9694,N_9994);
and UO_740 (O_740,N_9529,N_9719);
nor UO_741 (O_741,N_9635,N_9698);
or UO_742 (O_742,N_9922,N_9909);
and UO_743 (O_743,N_9684,N_9827);
nand UO_744 (O_744,N_9613,N_9927);
and UO_745 (O_745,N_9818,N_9924);
nor UO_746 (O_746,N_9899,N_9839);
or UO_747 (O_747,N_9946,N_9943);
and UO_748 (O_748,N_9508,N_9784);
nand UO_749 (O_749,N_9711,N_9867);
xnor UO_750 (O_750,N_9863,N_9884);
nand UO_751 (O_751,N_9731,N_9593);
nand UO_752 (O_752,N_9898,N_9925);
or UO_753 (O_753,N_9534,N_9832);
or UO_754 (O_754,N_9753,N_9888);
nor UO_755 (O_755,N_9579,N_9764);
or UO_756 (O_756,N_9580,N_9518);
nand UO_757 (O_757,N_9856,N_9517);
nor UO_758 (O_758,N_9534,N_9921);
and UO_759 (O_759,N_9688,N_9531);
and UO_760 (O_760,N_9617,N_9897);
nand UO_761 (O_761,N_9610,N_9842);
or UO_762 (O_762,N_9572,N_9785);
and UO_763 (O_763,N_9984,N_9739);
and UO_764 (O_764,N_9950,N_9666);
and UO_765 (O_765,N_9574,N_9559);
nand UO_766 (O_766,N_9653,N_9772);
nand UO_767 (O_767,N_9917,N_9956);
and UO_768 (O_768,N_9521,N_9534);
and UO_769 (O_769,N_9841,N_9550);
and UO_770 (O_770,N_9529,N_9743);
and UO_771 (O_771,N_9957,N_9571);
or UO_772 (O_772,N_9544,N_9948);
xor UO_773 (O_773,N_9540,N_9781);
nor UO_774 (O_774,N_9575,N_9660);
nand UO_775 (O_775,N_9702,N_9558);
and UO_776 (O_776,N_9775,N_9886);
and UO_777 (O_777,N_9674,N_9986);
nand UO_778 (O_778,N_9609,N_9679);
nor UO_779 (O_779,N_9604,N_9865);
xor UO_780 (O_780,N_9811,N_9750);
xnor UO_781 (O_781,N_9552,N_9906);
or UO_782 (O_782,N_9553,N_9564);
nor UO_783 (O_783,N_9874,N_9889);
nand UO_784 (O_784,N_9941,N_9894);
or UO_785 (O_785,N_9924,N_9873);
nand UO_786 (O_786,N_9876,N_9695);
and UO_787 (O_787,N_9696,N_9999);
nand UO_788 (O_788,N_9796,N_9802);
or UO_789 (O_789,N_9918,N_9932);
nand UO_790 (O_790,N_9811,N_9661);
nand UO_791 (O_791,N_9973,N_9513);
and UO_792 (O_792,N_9835,N_9855);
and UO_793 (O_793,N_9513,N_9595);
or UO_794 (O_794,N_9559,N_9938);
and UO_795 (O_795,N_9554,N_9809);
or UO_796 (O_796,N_9890,N_9728);
nor UO_797 (O_797,N_9662,N_9733);
or UO_798 (O_798,N_9705,N_9876);
nor UO_799 (O_799,N_9694,N_9861);
and UO_800 (O_800,N_9905,N_9679);
nand UO_801 (O_801,N_9541,N_9698);
nor UO_802 (O_802,N_9987,N_9771);
nor UO_803 (O_803,N_9526,N_9959);
and UO_804 (O_804,N_9683,N_9941);
and UO_805 (O_805,N_9904,N_9544);
and UO_806 (O_806,N_9671,N_9772);
nor UO_807 (O_807,N_9771,N_9891);
and UO_808 (O_808,N_9554,N_9935);
xor UO_809 (O_809,N_9514,N_9973);
nand UO_810 (O_810,N_9822,N_9900);
and UO_811 (O_811,N_9790,N_9547);
xnor UO_812 (O_812,N_9600,N_9586);
nand UO_813 (O_813,N_9555,N_9894);
and UO_814 (O_814,N_9888,N_9759);
nand UO_815 (O_815,N_9768,N_9963);
nor UO_816 (O_816,N_9782,N_9643);
and UO_817 (O_817,N_9897,N_9579);
or UO_818 (O_818,N_9576,N_9749);
nor UO_819 (O_819,N_9542,N_9658);
xor UO_820 (O_820,N_9530,N_9995);
nor UO_821 (O_821,N_9703,N_9652);
or UO_822 (O_822,N_9564,N_9709);
or UO_823 (O_823,N_9652,N_9620);
and UO_824 (O_824,N_9880,N_9990);
nand UO_825 (O_825,N_9562,N_9824);
nand UO_826 (O_826,N_9597,N_9946);
or UO_827 (O_827,N_9531,N_9881);
and UO_828 (O_828,N_9565,N_9628);
or UO_829 (O_829,N_9911,N_9783);
nand UO_830 (O_830,N_9539,N_9933);
nand UO_831 (O_831,N_9514,N_9579);
or UO_832 (O_832,N_9692,N_9833);
or UO_833 (O_833,N_9898,N_9705);
and UO_834 (O_834,N_9566,N_9764);
and UO_835 (O_835,N_9571,N_9955);
or UO_836 (O_836,N_9886,N_9721);
nand UO_837 (O_837,N_9981,N_9686);
nor UO_838 (O_838,N_9903,N_9952);
or UO_839 (O_839,N_9582,N_9968);
nand UO_840 (O_840,N_9557,N_9532);
nor UO_841 (O_841,N_9761,N_9583);
and UO_842 (O_842,N_9956,N_9674);
nand UO_843 (O_843,N_9960,N_9661);
xor UO_844 (O_844,N_9613,N_9617);
or UO_845 (O_845,N_9786,N_9529);
or UO_846 (O_846,N_9861,N_9638);
xnor UO_847 (O_847,N_9667,N_9626);
xor UO_848 (O_848,N_9853,N_9846);
and UO_849 (O_849,N_9536,N_9699);
or UO_850 (O_850,N_9829,N_9761);
xnor UO_851 (O_851,N_9800,N_9903);
nor UO_852 (O_852,N_9889,N_9769);
and UO_853 (O_853,N_9974,N_9758);
xnor UO_854 (O_854,N_9579,N_9649);
nor UO_855 (O_855,N_9869,N_9565);
or UO_856 (O_856,N_9581,N_9619);
xnor UO_857 (O_857,N_9908,N_9574);
nand UO_858 (O_858,N_9724,N_9934);
nand UO_859 (O_859,N_9872,N_9545);
nor UO_860 (O_860,N_9621,N_9890);
nand UO_861 (O_861,N_9737,N_9577);
nor UO_862 (O_862,N_9954,N_9613);
and UO_863 (O_863,N_9503,N_9985);
nand UO_864 (O_864,N_9970,N_9900);
nand UO_865 (O_865,N_9906,N_9938);
and UO_866 (O_866,N_9733,N_9690);
or UO_867 (O_867,N_9689,N_9848);
nor UO_868 (O_868,N_9691,N_9998);
nand UO_869 (O_869,N_9884,N_9951);
and UO_870 (O_870,N_9826,N_9744);
xor UO_871 (O_871,N_9522,N_9982);
nand UO_872 (O_872,N_9642,N_9667);
nand UO_873 (O_873,N_9542,N_9803);
nand UO_874 (O_874,N_9902,N_9841);
nand UO_875 (O_875,N_9579,N_9904);
nand UO_876 (O_876,N_9761,N_9522);
nand UO_877 (O_877,N_9860,N_9571);
nor UO_878 (O_878,N_9978,N_9706);
or UO_879 (O_879,N_9903,N_9975);
nand UO_880 (O_880,N_9682,N_9970);
nor UO_881 (O_881,N_9928,N_9780);
or UO_882 (O_882,N_9719,N_9641);
or UO_883 (O_883,N_9867,N_9629);
xor UO_884 (O_884,N_9613,N_9583);
or UO_885 (O_885,N_9502,N_9667);
or UO_886 (O_886,N_9706,N_9734);
nor UO_887 (O_887,N_9821,N_9616);
or UO_888 (O_888,N_9720,N_9723);
nor UO_889 (O_889,N_9610,N_9555);
nand UO_890 (O_890,N_9525,N_9778);
nor UO_891 (O_891,N_9651,N_9679);
nor UO_892 (O_892,N_9947,N_9610);
nand UO_893 (O_893,N_9991,N_9815);
nand UO_894 (O_894,N_9557,N_9639);
or UO_895 (O_895,N_9746,N_9827);
nor UO_896 (O_896,N_9831,N_9962);
or UO_897 (O_897,N_9745,N_9962);
nor UO_898 (O_898,N_9751,N_9634);
nor UO_899 (O_899,N_9999,N_9763);
and UO_900 (O_900,N_9681,N_9811);
or UO_901 (O_901,N_9925,N_9728);
nor UO_902 (O_902,N_9691,N_9879);
nand UO_903 (O_903,N_9958,N_9643);
nor UO_904 (O_904,N_9603,N_9919);
nand UO_905 (O_905,N_9591,N_9611);
and UO_906 (O_906,N_9971,N_9927);
nor UO_907 (O_907,N_9734,N_9874);
nand UO_908 (O_908,N_9560,N_9567);
nand UO_909 (O_909,N_9572,N_9854);
and UO_910 (O_910,N_9638,N_9712);
or UO_911 (O_911,N_9809,N_9803);
and UO_912 (O_912,N_9652,N_9906);
nand UO_913 (O_913,N_9936,N_9914);
or UO_914 (O_914,N_9782,N_9736);
nor UO_915 (O_915,N_9805,N_9625);
nor UO_916 (O_916,N_9580,N_9830);
and UO_917 (O_917,N_9805,N_9717);
nor UO_918 (O_918,N_9928,N_9544);
nand UO_919 (O_919,N_9738,N_9612);
and UO_920 (O_920,N_9897,N_9892);
nor UO_921 (O_921,N_9548,N_9857);
nand UO_922 (O_922,N_9945,N_9626);
or UO_923 (O_923,N_9806,N_9677);
and UO_924 (O_924,N_9694,N_9668);
nand UO_925 (O_925,N_9689,N_9981);
nor UO_926 (O_926,N_9599,N_9826);
nor UO_927 (O_927,N_9883,N_9513);
nor UO_928 (O_928,N_9700,N_9520);
or UO_929 (O_929,N_9540,N_9949);
or UO_930 (O_930,N_9685,N_9993);
or UO_931 (O_931,N_9590,N_9783);
and UO_932 (O_932,N_9756,N_9915);
nand UO_933 (O_933,N_9549,N_9928);
and UO_934 (O_934,N_9808,N_9873);
nand UO_935 (O_935,N_9966,N_9809);
xnor UO_936 (O_936,N_9772,N_9779);
nor UO_937 (O_937,N_9572,N_9694);
and UO_938 (O_938,N_9717,N_9942);
nand UO_939 (O_939,N_9508,N_9893);
nand UO_940 (O_940,N_9700,N_9616);
nand UO_941 (O_941,N_9676,N_9917);
nor UO_942 (O_942,N_9704,N_9743);
xor UO_943 (O_943,N_9970,N_9923);
or UO_944 (O_944,N_9541,N_9525);
xnor UO_945 (O_945,N_9745,N_9773);
xor UO_946 (O_946,N_9533,N_9933);
or UO_947 (O_947,N_9909,N_9700);
nor UO_948 (O_948,N_9800,N_9614);
nand UO_949 (O_949,N_9593,N_9788);
and UO_950 (O_950,N_9859,N_9716);
and UO_951 (O_951,N_9670,N_9532);
and UO_952 (O_952,N_9570,N_9981);
xor UO_953 (O_953,N_9670,N_9891);
nor UO_954 (O_954,N_9732,N_9960);
xor UO_955 (O_955,N_9830,N_9581);
or UO_956 (O_956,N_9935,N_9977);
nand UO_957 (O_957,N_9596,N_9544);
nor UO_958 (O_958,N_9813,N_9896);
nand UO_959 (O_959,N_9736,N_9942);
and UO_960 (O_960,N_9596,N_9581);
nand UO_961 (O_961,N_9764,N_9720);
or UO_962 (O_962,N_9842,N_9618);
xor UO_963 (O_963,N_9853,N_9833);
nor UO_964 (O_964,N_9592,N_9909);
or UO_965 (O_965,N_9569,N_9879);
nand UO_966 (O_966,N_9829,N_9929);
and UO_967 (O_967,N_9546,N_9542);
xnor UO_968 (O_968,N_9677,N_9977);
or UO_969 (O_969,N_9788,N_9987);
and UO_970 (O_970,N_9707,N_9613);
or UO_971 (O_971,N_9587,N_9677);
nor UO_972 (O_972,N_9505,N_9593);
nor UO_973 (O_973,N_9845,N_9538);
nor UO_974 (O_974,N_9797,N_9672);
nor UO_975 (O_975,N_9566,N_9639);
xnor UO_976 (O_976,N_9924,N_9717);
and UO_977 (O_977,N_9801,N_9611);
nand UO_978 (O_978,N_9863,N_9993);
nor UO_979 (O_979,N_9898,N_9916);
nand UO_980 (O_980,N_9680,N_9598);
and UO_981 (O_981,N_9521,N_9770);
xor UO_982 (O_982,N_9520,N_9572);
and UO_983 (O_983,N_9980,N_9509);
xnor UO_984 (O_984,N_9861,N_9829);
nor UO_985 (O_985,N_9953,N_9935);
xnor UO_986 (O_986,N_9950,N_9827);
and UO_987 (O_987,N_9706,N_9710);
xor UO_988 (O_988,N_9756,N_9927);
or UO_989 (O_989,N_9514,N_9919);
nand UO_990 (O_990,N_9758,N_9736);
and UO_991 (O_991,N_9928,N_9605);
nor UO_992 (O_992,N_9902,N_9743);
and UO_993 (O_993,N_9734,N_9515);
xnor UO_994 (O_994,N_9931,N_9594);
and UO_995 (O_995,N_9876,N_9849);
nor UO_996 (O_996,N_9830,N_9877);
or UO_997 (O_997,N_9934,N_9554);
or UO_998 (O_998,N_9899,N_9852);
nand UO_999 (O_999,N_9874,N_9585);
or UO_1000 (O_1000,N_9692,N_9804);
nor UO_1001 (O_1001,N_9673,N_9692);
and UO_1002 (O_1002,N_9981,N_9748);
nand UO_1003 (O_1003,N_9624,N_9679);
xor UO_1004 (O_1004,N_9532,N_9588);
nor UO_1005 (O_1005,N_9956,N_9535);
and UO_1006 (O_1006,N_9556,N_9598);
or UO_1007 (O_1007,N_9585,N_9898);
nor UO_1008 (O_1008,N_9955,N_9689);
or UO_1009 (O_1009,N_9798,N_9987);
xor UO_1010 (O_1010,N_9512,N_9660);
and UO_1011 (O_1011,N_9884,N_9829);
or UO_1012 (O_1012,N_9769,N_9556);
xnor UO_1013 (O_1013,N_9962,N_9984);
nand UO_1014 (O_1014,N_9728,N_9595);
nor UO_1015 (O_1015,N_9982,N_9714);
nand UO_1016 (O_1016,N_9840,N_9623);
nor UO_1017 (O_1017,N_9800,N_9863);
nand UO_1018 (O_1018,N_9838,N_9579);
and UO_1019 (O_1019,N_9585,N_9958);
and UO_1020 (O_1020,N_9890,N_9794);
nor UO_1021 (O_1021,N_9763,N_9865);
or UO_1022 (O_1022,N_9902,N_9994);
nand UO_1023 (O_1023,N_9785,N_9987);
or UO_1024 (O_1024,N_9801,N_9837);
and UO_1025 (O_1025,N_9667,N_9770);
or UO_1026 (O_1026,N_9901,N_9532);
and UO_1027 (O_1027,N_9928,N_9608);
or UO_1028 (O_1028,N_9932,N_9693);
nor UO_1029 (O_1029,N_9844,N_9577);
or UO_1030 (O_1030,N_9906,N_9619);
nor UO_1031 (O_1031,N_9806,N_9536);
nor UO_1032 (O_1032,N_9908,N_9507);
nor UO_1033 (O_1033,N_9543,N_9718);
nor UO_1034 (O_1034,N_9927,N_9521);
nor UO_1035 (O_1035,N_9702,N_9773);
or UO_1036 (O_1036,N_9791,N_9522);
nand UO_1037 (O_1037,N_9640,N_9734);
and UO_1038 (O_1038,N_9925,N_9928);
and UO_1039 (O_1039,N_9516,N_9925);
or UO_1040 (O_1040,N_9735,N_9832);
or UO_1041 (O_1041,N_9800,N_9822);
and UO_1042 (O_1042,N_9931,N_9612);
nand UO_1043 (O_1043,N_9999,N_9679);
nor UO_1044 (O_1044,N_9892,N_9917);
or UO_1045 (O_1045,N_9707,N_9774);
or UO_1046 (O_1046,N_9732,N_9809);
and UO_1047 (O_1047,N_9691,N_9682);
nand UO_1048 (O_1048,N_9866,N_9518);
and UO_1049 (O_1049,N_9965,N_9520);
and UO_1050 (O_1050,N_9910,N_9928);
nor UO_1051 (O_1051,N_9836,N_9625);
or UO_1052 (O_1052,N_9634,N_9955);
and UO_1053 (O_1053,N_9654,N_9741);
or UO_1054 (O_1054,N_9806,N_9559);
or UO_1055 (O_1055,N_9652,N_9956);
and UO_1056 (O_1056,N_9506,N_9654);
and UO_1057 (O_1057,N_9942,N_9840);
nand UO_1058 (O_1058,N_9778,N_9693);
or UO_1059 (O_1059,N_9930,N_9621);
or UO_1060 (O_1060,N_9914,N_9642);
xnor UO_1061 (O_1061,N_9562,N_9935);
nand UO_1062 (O_1062,N_9637,N_9857);
nand UO_1063 (O_1063,N_9617,N_9668);
nor UO_1064 (O_1064,N_9985,N_9616);
nor UO_1065 (O_1065,N_9677,N_9747);
nor UO_1066 (O_1066,N_9648,N_9559);
or UO_1067 (O_1067,N_9967,N_9998);
nand UO_1068 (O_1068,N_9677,N_9745);
or UO_1069 (O_1069,N_9938,N_9927);
and UO_1070 (O_1070,N_9660,N_9658);
xnor UO_1071 (O_1071,N_9752,N_9745);
and UO_1072 (O_1072,N_9537,N_9686);
nand UO_1073 (O_1073,N_9741,N_9870);
xnor UO_1074 (O_1074,N_9797,N_9614);
xor UO_1075 (O_1075,N_9755,N_9719);
nand UO_1076 (O_1076,N_9661,N_9823);
or UO_1077 (O_1077,N_9557,N_9512);
and UO_1078 (O_1078,N_9800,N_9906);
nand UO_1079 (O_1079,N_9952,N_9719);
nor UO_1080 (O_1080,N_9507,N_9751);
nand UO_1081 (O_1081,N_9834,N_9503);
nor UO_1082 (O_1082,N_9563,N_9959);
nand UO_1083 (O_1083,N_9510,N_9800);
or UO_1084 (O_1084,N_9698,N_9625);
nand UO_1085 (O_1085,N_9646,N_9909);
nand UO_1086 (O_1086,N_9845,N_9750);
nand UO_1087 (O_1087,N_9821,N_9655);
nor UO_1088 (O_1088,N_9761,N_9924);
and UO_1089 (O_1089,N_9765,N_9771);
or UO_1090 (O_1090,N_9903,N_9598);
or UO_1091 (O_1091,N_9734,N_9771);
nor UO_1092 (O_1092,N_9613,N_9844);
xor UO_1093 (O_1093,N_9698,N_9630);
nand UO_1094 (O_1094,N_9572,N_9984);
nor UO_1095 (O_1095,N_9948,N_9622);
nor UO_1096 (O_1096,N_9701,N_9569);
xnor UO_1097 (O_1097,N_9809,N_9574);
xor UO_1098 (O_1098,N_9686,N_9795);
or UO_1099 (O_1099,N_9673,N_9967);
nand UO_1100 (O_1100,N_9834,N_9511);
nand UO_1101 (O_1101,N_9701,N_9978);
and UO_1102 (O_1102,N_9798,N_9730);
xnor UO_1103 (O_1103,N_9983,N_9723);
nand UO_1104 (O_1104,N_9722,N_9929);
nand UO_1105 (O_1105,N_9594,N_9847);
and UO_1106 (O_1106,N_9693,N_9689);
nor UO_1107 (O_1107,N_9933,N_9844);
or UO_1108 (O_1108,N_9571,N_9660);
xor UO_1109 (O_1109,N_9792,N_9705);
and UO_1110 (O_1110,N_9983,N_9960);
and UO_1111 (O_1111,N_9704,N_9717);
nor UO_1112 (O_1112,N_9781,N_9848);
xnor UO_1113 (O_1113,N_9791,N_9945);
nor UO_1114 (O_1114,N_9837,N_9641);
nor UO_1115 (O_1115,N_9727,N_9907);
xnor UO_1116 (O_1116,N_9892,N_9602);
nor UO_1117 (O_1117,N_9781,N_9711);
or UO_1118 (O_1118,N_9737,N_9584);
nor UO_1119 (O_1119,N_9898,N_9604);
and UO_1120 (O_1120,N_9942,N_9526);
nand UO_1121 (O_1121,N_9762,N_9648);
nand UO_1122 (O_1122,N_9784,N_9617);
nor UO_1123 (O_1123,N_9525,N_9655);
or UO_1124 (O_1124,N_9716,N_9711);
or UO_1125 (O_1125,N_9557,N_9591);
or UO_1126 (O_1126,N_9829,N_9907);
or UO_1127 (O_1127,N_9641,N_9987);
nor UO_1128 (O_1128,N_9565,N_9654);
and UO_1129 (O_1129,N_9794,N_9982);
nand UO_1130 (O_1130,N_9643,N_9530);
xor UO_1131 (O_1131,N_9591,N_9972);
or UO_1132 (O_1132,N_9633,N_9944);
or UO_1133 (O_1133,N_9698,N_9845);
or UO_1134 (O_1134,N_9817,N_9573);
nand UO_1135 (O_1135,N_9549,N_9911);
and UO_1136 (O_1136,N_9992,N_9867);
and UO_1137 (O_1137,N_9727,N_9617);
xnor UO_1138 (O_1138,N_9688,N_9581);
nand UO_1139 (O_1139,N_9886,N_9560);
nand UO_1140 (O_1140,N_9645,N_9658);
or UO_1141 (O_1141,N_9636,N_9551);
nor UO_1142 (O_1142,N_9520,N_9818);
and UO_1143 (O_1143,N_9787,N_9629);
and UO_1144 (O_1144,N_9540,N_9759);
or UO_1145 (O_1145,N_9636,N_9545);
nor UO_1146 (O_1146,N_9698,N_9822);
or UO_1147 (O_1147,N_9986,N_9561);
nand UO_1148 (O_1148,N_9700,N_9821);
and UO_1149 (O_1149,N_9768,N_9802);
nor UO_1150 (O_1150,N_9762,N_9584);
and UO_1151 (O_1151,N_9547,N_9704);
xnor UO_1152 (O_1152,N_9767,N_9542);
xnor UO_1153 (O_1153,N_9911,N_9977);
and UO_1154 (O_1154,N_9655,N_9880);
or UO_1155 (O_1155,N_9581,N_9977);
nor UO_1156 (O_1156,N_9862,N_9740);
or UO_1157 (O_1157,N_9949,N_9773);
and UO_1158 (O_1158,N_9563,N_9586);
nor UO_1159 (O_1159,N_9952,N_9842);
nand UO_1160 (O_1160,N_9996,N_9879);
nor UO_1161 (O_1161,N_9634,N_9787);
nand UO_1162 (O_1162,N_9901,N_9839);
nor UO_1163 (O_1163,N_9832,N_9977);
nand UO_1164 (O_1164,N_9846,N_9773);
nor UO_1165 (O_1165,N_9982,N_9891);
and UO_1166 (O_1166,N_9655,N_9817);
nor UO_1167 (O_1167,N_9790,N_9753);
or UO_1168 (O_1168,N_9678,N_9680);
or UO_1169 (O_1169,N_9885,N_9594);
or UO_1170 (O_1170,N_9868,N_9858);
and UO_1171 (O_1171,N_9506,N_9821);
nor UO_1172 (O_1172,N_9598,N_9937);
or UO_1173 (O_1173,N_9824,N_9699);
or UO_1174 (O_1174,N_9738,N_9517);
nor UO_1175 (O_1175,N_9793,N_9887);
nor UO_1176 (O_1176,N_9900,N_9624);
or UO_1177 (O_1177,N_9658,N_9720);
and UO_1178 (O_1178,N_9517,N_9682);
nor UO_1179 (O_1179,N_9536,N_9755);
or UO_1180 (O_1180,N_9615,N_9717);
and UO_1181 (O_1181,N_9580,N_9583);
and UO_1182 (O_1182,N_9913,N_9555);
nand UO_1183 (O_1183,N_9765,N_9564);
or UO_1184 (O_1184,N_9702,N_9960);
nor UO_1185 (O_1185,N_9963,N_9538);
nand UO_1186 (O_1186,N_9570,N_9655);
or UO_1187 (O_1187,N_9562,N_9893);
nand UO_1188 (O_1188,N_9856,N_9745);
and UO_1189 (O_1189,N_9975,N_9526);
xnor UO_1190 (O_1190,N_9958,N_9538);
or UO_1191 (O_1191,N_9809,N_9842);
nand UO_1192 (O_1192,N_9561,N_9577);
or UO_1193 (O_1193,N_9500,N_9842);
nand UO_1194 (O_1194,N_9799,N_9914);
nand UO_1195 (O_1195,N_9790,N_9718);
and UO_1196 (O_1196,N_9834,N_9557);
xnor UO_1197 (O_1197,N_9974,N_9633);
xor UO_1198 (O_1198,N_9806,N_9638);
nor UO_1199 (O_1199,N_9500,N_9771);
nand UO_1200 (O_1200,N_9575,N_9539);
xnor UO_1201 (O_1201,N_9923,N_9941);
nor UO_1202 (O_1202,N_9767,N_9520);
nor UO_1203 (O_1203,N_9546,N_9574);
or UO_1204 (O_1204,N_9707,N_9531);
and UO_1205 (O_1205,N_9614,N_9763);
nor UO_1206 (O_1206,N_9745,N_9876);
and UO_1207 (O_1207,N_9839,N_9759);
nor UO_1208 (O_1208,N_9965,N_9550);
xor UO_1209 (O_1209,N_9530,N_9621);
nand UO_1210 (O_1210,N_9673,N_9521);
and UO_1211 (O_1211,N_9929,N_9535);
nor UO_1212 (O_1212,N_9657,N_9975);
or UO_1213 (O_1213,N_9537,N_9690);
or UO_1214 (O_1214,N_9742,N_9935);
or UO_1215 (O_1215,N_9618,N_9505);
or UO_1216 (O_1216,N_9527,N_9664);
and UO_1217 (O_1217,N_9528,N_9665);
xnor UO_1218 (O_1218,N_9745,N_9711);
nand UO_1219 (O_1219,N_9585,N_9904);
nor UO_1220 (O_1220,N_9941,N_9664);
nor UO_1221 (O_1221,N_9503,N_9937);
and UO_1222 (O_1222,N_9923,N_9797);
nand UO_1223 (O_1223,N_9729,N_9869);
nor UO_1224 (O_1224,N_9996,N_9926);
or UO_1225 (O_1225,N_9702,N_9891);
or UO_1226 (O_1226,N_9507,N_9978);
or UO_1227 (O_1227,N_9962,N_9806);
or UO_1228 (O_1228,N_9712,N_9705);
nor UO_1229 (O_1229,N_9568,N_9778);
xnor UO_1230 (O_1230,N_9629,N_9634);
nor UO_1231 (O_1231,N_9604,N_9958);
nor UO_1232 (O_1232,N_9841,N_9687);
or UO_1233 (O_1233,N_9952,N_9649);
and UO_1234 (O_1234,N_9522,N_9777);
and UO_1235 (O_1235,N_9930,N_9754);
or UO_1236 (O_1236,N_9947,N_9937);
nand UO_1237 (O_1237,N_9573,N_9937);
xnor UO_1238 (O_1238,N_9569,N_9868);
nand UO_1239 (O_1239,N_9952,N_9523);
or UO_1240 (O_1240,N_9841,N_9662);
nand UO_1241 (O_1241,N_9864,N_9782);
nor UO_1242 (O_1242,N_9538,N_9998);
nand UO_1243 (O_1243,N_9818,N_9753);
nor UO_1244 (O_1244,N_9838,N_9515);
and UO_1245 (O_1245,N_9840,N_9673);
nor UO_1246 (O_1246,N_9946,N_9757);
nor UO_1247 (O_1247,N_9702,N_9749);
nand UO_1248 (O_1248,N_9765,N_9659);
or UO_1249 (O_1249,N_9503,N_9950);
xnor UO_1250 (O_1250,N_9775,N_9560);
nor UO_1251 (O_1251,N_9503,N_9916);
or UO_1252 (O_1252,N_9924,N_9539);
or UO_1253 (O_1253,N_9654,N_9668);
nor UO_1254 (O_1254,N_9594,N_9822);
nor UO_1255 (O_1255,N_9626,N_9660);
nand UO_1256 (O_1256,N_9848,N_9943);
and UO_1257 (O_1257,N_9624,N_9924);
nand UO_1258 (O_1258,N_9872,N_9935);
and UO_1259 (O_1259,N_9578,N_9723);
nor UO_1260 (O_1260,N_9845,N_9770);
or UO_1261 (O_1261,N_9814,N_9638);
and UO_1262 (O_1262,N_9856,N_9622);
nand UO_1263 (O_1263,N_9520,N_9690);
xor UO_1264 (O_1264,N_9574,N_9530);
nor UO_1265 (O_1265,N_9545,N_9731);
or UO_1266 (O_1266,N_9828,N_9713);
nand UO_1267 (O_1267,N_9786,N_9561);
and UO_1268 (O_1268,N_9853,N_9564);
and UO_1269 (O_1269,N_9886,N_9587);
or UO_1270 (O_1270,N_9890,N_9922);
nand UO_1271 (O_1271,N_9752,N_9527);
and UO_1272 (O_1272,N_9578,N_9857);
and UO_1273 (O_1273,N_9727,N_9529);
nor UO_1274 (O_1274,N_9585,N_9543);
and UO_1275 (O_1275,N_9638,N_9739);
nand UO_1276 (O_1276,N_9532,N_9844);
nor UO_1277 (O_1277,N_9765,N_9882);
or UO_1278 (O_1278,N_9923,N_9642);
or UO_1279 (O_1279,N_9925,N_9720);
and UO_1280 (O_1280,N_9799,N_9771);
nand UO_1281 (O_1281,N_9534,N_9686);
and UO_1282 (O_1282,N_9848,N_9912);
and UO_1283 (O_1283,N_9862,N_9621);
or UO_1284 (O_1284,N_9730,N_9821);
or UO_1285 (O_1285,N_9927,N_9590);
nor UO_1286 (O_1286,N_9585,N_9924);
or UO_1287 (O_1287,N_9990,N_9916);
or UO_1288 (O_1288,N_9505,N_9827);
xnor UO_1289 (O_1289,N_9996,N_9708);
or UO_1290 (O_1290,N_9644,N_9654);
xor UO_1291 (O_1291,N_9592,N_9676);
nor UO_1292 (O_1292,N_9789,N_9624);
and UO_1293 (O_1293,N_9699,N_9675);
nor UO_1294 (O_1294,N_9697,N_9837);
and UO_1295 (O_1295,N_9657,N_9720);
and UO_1296 (O_1296,N_9702,N_9580);
xor UO_1297 (O_1297,N_9586,N_9809);
nand UO_1298 (O_1298,N_9962,N_9561);
nor UO_1299 (O_1299,N_9681,N_9905);
nand UO_1300 (O_1300,N_9936,N_9957);
xor UO_1301 (O_1301,N_9644,N_9891);
or UO_1302 (O_1302,N_9576,N_9642);
or UO_1303 (O_1303,N_9835,N_9720);
and UO_1304 (O_1304,N_9696,N_9974);
nor UO_1305 (O_1305,N_9860,N_9778);
xnor UO_1306 (O_1306,N_9722,N_9944);
nor UO_1307 (O_1307,N_9563,N_9725);
or UO_1308 (O_1308,N_9925,N_9844);
or UO_1309 (O_1309,N_9511,N_9930);
or UO_1310 (O_1310,N_9783,N_9534);
and UO_1311 (O_1311,N_9558,N_9624);
nand UO_1312 (O_1312,N_9858,N_9532);
or UO_1313 (O_1313,N_9522,N_9703);
nor UO_1314 (O_1314,N_9500,N_9812);
and UO_1315 (O_1315,N_9612,N_9866);
and UO_1316 (O_1316,N_9925,N_9526);
xnor UO_1317 (O_1317,N_9799,N_9783);
nor UO_1318 (O_1318,N_9738,N_9679);
and UO_1319 (O_1319,N_9676,N_9858);
or UO_1320 (O_1320,N_9573,N_9959);
xor UO_1321 (O_1321,N_9886,N_9995);
nand UO_1322 (O_1322,N_9626,N_9860);
and UO_1323 (O_1323,N_9861,N_9990);
xnor UO_1324 (O_1324,N_9935,N_9806);
or UO_1325 (O_1325,N_9503,N_9624);
and UO_1326 (O_1326,N_9596,N_9656);
nor UO_1327 (O_1327,N_9573,N_9998);
and UO_1328 (O_1328,N_9507,N_9802);
nand UO_1329 (O_1329,N_9630,N_9839);
or UO_1330 (O_1330,N_9966,N_9723);
nand UO_1331 (O_1331,N_9799,N_9669);
nand UO_1332 (O_1332,N_9613,N_9861);
or UO_1333 (O_1333,N_9971,N_9932);
nand UO_1334 (O_1334,N_9579,N_9710);
nor UO_1335 (O_1335,N_9599,N_9676);
and UO_1336 (O_1336,N_9911,N_9718);
nor UO_1337 (O_1337,N_9695,N_9557);
nor UO_1338 (O_1338,N_9814,N_9894);
nand UO_1339 (O_1339,N_9619,N_9847);
nor UO_1340 (O_1340,N_9645,N_9868);
or UO_1341 (O_1341,N_9716,N_9634);
or UO_1342 (O_1342,N_9936,N_9831);
nor UO_1343 (O_1343,N_9852,N_9629);
and UO_1344 (O_1344,N_9854,N_9528);
or UO_1345 (O_1345,N_9743,N_9804);
or UO_1346 (O_1346,N_9725,N_9540);
and UO_1347 (O_1347,N_9985,N_9770);
nand UO_1348 (O_1348,N_9982,N_9835);
and UO_1349 (O_1349,N_9943,N_9879);
nor UO_1350 (O_1350,N_9567,N_9713);
nand UO_1351 (O_1351,N_9558,N_9836);
nand UO_1352 (O_1352,N_9504,N_9745);
nand UO_1353 (O_1353,N_9745,N_9751);
and UO_1354 (O_1354,N_9599,N_9991);
nor UO_1355 (O_1355,N_9705,N_9914);
nand UO_1356 (O_1356,N_9656,N_9982);
nor UO_1357 (O_1357,N_9749,N_9570);
and UO_1358 (O_1358,N_9739,N_9537);
or UO_1359 (O_1359,N_9882,N_9629);
nand UO_1360 (O_1360,N_9992,N_9552);
and UO_1361 (O_1361,N_9837,N_9831);
xor UO_1362 (O_1362,N_9937,N_9815);
and UO_1363 (O_1363,N_9771,N_9951);
or UO_1364 (O_1364,N_9534,N_9763);
or UO_1365 (O_1365,N_9733,N_9889);
or UO_1366 (O_1366,N_9635,N_9619);
or UO_1367 (O_1367,N_9833,N_9884);
nor UO_1368 (O_1368,N_9518,N_9986);
xor UO_1369 (O_1369,N_9770,N_9901);
nor UO_1370 (O_1370,N_9695,N_9660);
or UO_1371 (O_1371,N_9539,N_9720);
and UO_1372 (O_1372,N_9708,N_9699);
nor UO_1373 (O_1373,N_9930,N_9898);
nor UO_1374 (O_1374,N_9697,N_9502);
nand UO_1375 (O_1375,N_9643,N_9911);
and UO_1376 (O_1376,N_9622,N_9895);
nor UO_1377 (O_1377,N_9819,N_9954);
nand UO_1378 (O_1378,N_9890,N_9508);
or UO_1379 (O_1379,N_9874,N_9710);
or UO_1380 (O_1380,N_9686,N_9613);
nor UO_1381 (O_1381,N_9583,N_9699);
nor UO_1382 (O_1382,N_9641,N_9569);
nor UO_1383 (O_1383,N_9646,N_9984);
nor UO_1384 (O_1384,N_9547,N_9861);
nor UO_1385 (O_1385,N_9564,N_9611);
nand UO_1386 (O_1386,N_9981,N_9530);
and UO_1387 (O_1387,N_9623,N_9743);
nor UO_1388 (O_1388,N_9889,N_9576);
nand UO_1389 (O_1389,N_9975,N_9727);
nor UO_1390 (O_1390,N_9798,N_9675);
and UO_1391 (O_1391,N_9977,N_9678);
or UO_1392 (O_1392,N_9784,N_9876);
nor UO_1393 (O_1393,N_9711,N_9687);
and UO_1394 (O_1394,N_9866,N_9820);
nand UO_1395 (O_1395,N_9740,N_9686);
or UO_1396 (O_1396,N_9955,N_9784);
nor UO_1397 (O_1397,N_9817,N_9631);
nand UO_1398 (O_1398,N_9906,N_9612);
nor UO_1399 (O_1399,N_9722,N_9917);
nor UO_1400 (O_1400,N_9581,N_9911);
and UO_1401 (O_1401,N_9912,N_9745);
and UO_1402 (O_1402,N_9877,N_9938);
and UO_1403 (O_1403,N_9713,N_9937);
nand UO_1404 (O_1404,N_9799,N_9723);
and UO_1405 (O_1405,N_9632,N_9645);
and UO_1406 (O_1406,N_9565,N_9642);
and UO_1407 (O_1407,N_9622,N_9966);
nand UO_1408 (O_1408,N_9998,N_9947);
nand UO_1409 (O_1409,N_9531,N_9577);
nand UO_1410 (O_1410,N_9574,N_9937);
nor UO_1411 (O_1411,N_9536,N_9741);
nand UO_1412 (O_1412,N_9586,N_9989);
xor UO_1413 (O_1413,N_9960,N_9989);
nand UO_1414 (O_1414,N_9633,N_9789);
nor UO_1415 (O_1415,N_9512,N_9935);
or UO_1416 (O_1416,N_9819,N_9683);
nand UO_1417 (O_1417,N_9866,N_9928);
or UO_1418 (O_1418,N_9917,N_9844);
or UO_1419 (O_1419,N_9894,N_9657);
xnor UO_1420 (O_1420,N_9674,N_9988);
and UO_1421 (O_1421,N_9962,N_9570);
nand UO_1422 (O_1422,N_9875,N_9878);
or UO_1423 (O_1423,N_9930,N_9743);
and UO_1424 (O_1424,N_9588,N_9680);
nor UO_1425 (O_1425,N_9981,N_9708);
and UO_1426 (O_1426,N_9981,N_9903);
nor UO_1427 (O_1427,N_9536,N_9529);
nor UO_1428 (O_1428,N_9989,N_9671);
nor UO_1429 (O_1429,N_9920,N_9918);
or UO_1430 (O_1430,N_9532,N_9566);
or UO_1431 (O_1431,N_9633,N_9833);
or UO_1432 (O_1432,N_9696,N_9733);
and UO_1433 (O_1433,N_9734,N_9716);
or UO_1434 (O_1434,N_9989,N_9757);
nand UO_1435 (O_1435,N_9855,N_9780);
or UO_1436 (O_1436,N_9810,N_9622);
or UO_1437 (O_1437,N_9858,N_9541);
nor UO_1438 (O_1438,N_9732,N_9773);
or UO_1439 (O_1439,N_9514,N_9926);
nand UO_1440 (O_1440,N_9913,N_9835);
or UO_1441 (O_1441,N_9595,N_9761);
nand UO_1442 (O_1442,N_9664,N_9915);
and UO_1443 (O_1443,N_9784,N_9877);
and UO_1444 (O_1444,N_9809,N_9872);
and UO_1445 (O_1445,N_9727,N_9507);
xnor UO_1446 (O_1446,N_9995,N_9884);
nand UO_1447 (O_1447,N_9784,N_9778);
and UO_1448 (O_1448,N_9584,N_9851);
nor UO_1449 (O_1449,N_9762,N_9880);
nor UO_1450 (O_1450,N_9795,N_9584);
and UO_1451 (O_1451,N_9904,N_9849);
nand UO_1452 (O_1452,N_9681,N_9772);
and UO_1453 (O_1453,N_9598,N_9581);
nor UO_1454 (O_1454,N_9774,N_9861);
or UO_1455 (O_1455,N_9606,N_9877);
or UO_1456 (O_1456,N_9993,N_9922);
nand UO_1457 (O_1457,N_9893,N_9728);
nor UO_1458 (O_1458,N_9527,N_9938);
or UO_1459 (O_1459,N_9837,N_9995);
nor UO_1460 (O_1460,N_9675,N_9868);
nand UO_1461 (O_1461,N_9710,N_9635);
and UO_1462 (O_1462,N_9503,N_9640);
or UO_1463 (O_1463,N_9720,N_9619);
xor UO_1464 (O_1464,N_9768,N_9573);
and UO_1465 (O_1465,N_9822,N_9829);
nor UO_1466 (O_1466,N_9535,N_9742);
and UO_1467 (O_1467,N_9532,N_9680);
and UO_1468 (O_1468,N_9638,N_9598);
or UO_1469 (O_1469,N_9631,N_9513);
and UO_1470 (O_1470,N_9723,N_9623);
nand UO_1471 (O_1471,N_9548,N_9533);
nor UO_1472 (O_1472,N_9854,N_9843);
xnor UO_1473 (O_1473,N_9824,N_9973);
nor UO_1474 (O_1474,N_9538,N_9832);
nor UO_1475 (O_1475,N_9544,N_9816);
nand UO_1476 (O_1476,N_9528,N_9677);
and UO_1477 (O_1477,N_9939,N_9673);
nand UO_1478 (O_1478,N_9617,N_9753);
nand UO_1479 (O_1479,N_9531,N_9914);
and UO_1480 (O_1480,N_9878,N_9929);
xnor UO_1481 (O_1481,N_9734,N_9662);
or UO_1482 (O_1482,N_9962,N_9889);
and UO_1483 (O_1483,N_9599,N_9588);
xor UO_1484 (O_1484,N_9902,N_9622);
nor UO_1485 (O_1485,N_9929,N_9784);
nand UO_1486 (O_1486,N_9619,N_9618);
nand UO_1487 (O_1487,N_9874,N_9538);
or UO_1488 (O_1488,N_9856,N_9992);
nor UO_1489 (O_1489,N_9551,N_9863);
and UO_1490 (O_1490,N_9886,N_9555);
and UO_1491 (O_1491,N_9547,N_9662);
and UO_1492 (O_1492,N_9985,N_9859);
xor UO_1493 (O_1493,N_9691,N_9722);
nor UO_1494 (O_1494,N_9789,N_9718);
and UO_1495 (O_1495,N_9672,N_9996);
nand UO_1496 (O_1496,N_9629,N_9775);
and UO_1497 (O_1497,N_9748,N_9649);
and UO_1498 (O_1498,N_9735,N_9517);
nand UO_1499 (O_1499,N_9692,N_9551);
endmodule