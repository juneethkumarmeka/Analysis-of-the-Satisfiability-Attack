module basic_2000_20000_2500_10_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
xor U0 (N_0,In_356,In_261);
or U1 (N_1,In_957,In_1030);
or U2 (N_2,In_1325,In_1168);
nor U3 (N_3,In_1853,In_1666);
nand U4 (N_4,In_1899,In_1454);
nor U5 (N_5,In_1073,In_414);
or U6 (N_6,In_701,In_65);
or U7 (N_7,In_1163,In_1694);
or U8 (N_8,In_1814,In_447);
nand U9 (N_9,In_1486,In_1581);
nor U10 (N_10,In_1265,In_245);
nor U11 (N_11,In_933,In_1852);
nand U12 (N_12,In_321,In_1643);
or U13 (N_13,In_15,In_379);
xor U14 (N_14,In_1287,In_1092);
or U15 (N_15,In_1578,In_1941);
nor U16 (N_16,In_738,In_365);
or U17 (N_17,In_1065,In_707);
nand U18 (N_18,In_1904,In_1742);
xor U19 (N_19,In_75,In_1562);
and U20 (N_20,In_1056,In_1902);
nand U21 (N_21,In_1681,In_1826);
nor U22 (N_22,In_1245,In_1131);
nand U23 (N_23,In_146,In_1232);
or U24 (N_24,In_1790,In_887);
xnor U25 (N_25,In_1502,In_1665);
xnor U26 (N_26,In_541,In_680);
and U27 (N_27,In_1521,In_740);
and U28 (N_28,In_1858,In_499);
and U29 (N_29,In_1690,In_1607);
or U30 (N_30,In_880,In_684);
xor U31 (N_31,In_478,In_861);
or U32 (N_32,In_1201,In_609);
xor U33 (N_33,In_1239,In_1836);
or U34 (N_34,In_1250,In_1039);
nand U35 (N_35,In_1376,In_813);
and U36 (N_36,In_1133,In_1429);
and U37 (N_37,In_605,In_612);
and U38 (N_38,In_1362,In_1075);
and U39 (N_39,In_885,In_1687);
or U40 (N_40,In_1512,In_675);
xor U41 (N_41,In_1328,In_1886);
xor U42 (N_42,In_1017,In_390);
nand U43 (N_43,In_194,In_1966);
xnor U44 (N_44,In_656,In_1164);
or U45 (N_45,In_1008,In_399);
and U46 (N_46,In_1156,In_1262);
xor U47 (N_47,In_662,In_1276);
and U48 (N_48,In_255,In_1183);
or U49 (N_49,In_529,In_1530);
nor U50 (N_50,In_1942,In_1612);
xnor U51 (N_51,In_1700,In_1460);
nand U52 (N_52,In_1476,In_1193);
xor U53 (N_53,In_905,In_1069);
xnor U54 (N_54,In_1820,In_98);
nand U55 (N_55,In_442,In_988);
nand U56 (N_56,In_1273,In_185);
nand U57 (N_57,In_1304,In_1206);
nand U58 (N_58,In_372,In_79);
nand U59 (N_59,In_1103,In_1513);
and U60 (N_60,In_275,In_1055);
nand U61 (N_61,In_470,In_1586);
xnor U62 (N_62,In_1060,In_1143);
nand U63 (N_63,In_1237,In_1182);
nand U64 (N_64,In_491,In_1811);
nand U65 (N_65,In_20,In_1072);
and U66 (N_66,In_434,In_1360);
nor U67 (N_67,In_1741,In_117);
or U68 (N_68,In_103,In_1518);
nand U69 (N_69,In_1257,In_980);
or U70 (N_70,In_133,In_1298);
nor U71 (N_71,In_1652,In_1441);
nand U72 (N_72,In_697,In_949);
nand U73 (N_73,In_235,In_52);
nand U74 (N_74,In_500,In_1846);
nor U75 (N_75,In_741,In_349);
and U76 (N_76,In_1228,In_1863);
nand U77 (N_77,In_918,In_213);
nand U78 (N_78,In_281,In_420);
nor U79 (N_79,In_144,In_1340);
nor U80 (N_80,In_1988,In_1765);
nand U81 (N_81,In_1301,In_833);
nor U82 (N_82,In_712,In_1939);
or U83 (N_83,In_1066,In_579);
nor U84 (N_84,In_1884,In_1189);
nor U85 (N_85,In_200,In_790);
nand U86 (N_86,In_318,In_1745);
and U87 (N_87,In_1599,In_222);
nor U88 (N_88,In_114,In_1480);
nand U89 (N_89,In_1209,In_815);
and U90 (N_90,In_601,In_538);
and U91 (N_91,In_550,In_1874);
nor U92 (N_92,In_1554,In_882);
xor U93 (N_93,In_1491,In_1101);
xor U94 (N_94,In_1013,In_630);
or U95 (N_95,In_1217,In_11);
or U96 (N_96,In_839,In_273);
and U97 (N_97,In_182,In_92);
nor U98 (N_98,In_651,In_331);
nand U99 (N_99,In_1947,In_821);
and U100 (N_100,In_5,In_1061);
nor U101 (N_101,In_565,In_1969);
nand U102 (N_102,In_46,In_1769);
xnor U103 (N_103,In_115,In_1608);
and U104 (N_104,In_1383,In_1087);
nand U105 (N_105,In_1719,In_644);
xor U106 (N_106,In_181,In_867);
and U107 (N_107,In_421,In_663);
and U108 (N_108,In_1354,In_418);
or U109 (N_109,In_1344,In_483);
or U110 (N_110,In_568,In_1597);
and U111 (N_111,In_472,In_971);
nor U112 (N_112,In_551,In_1861);
or U113 (N_113,In_505,In_1181);
xor U114 (N_114,In_919,In_1375);
or U115 (N_115,In_481,In_105);
or U116 (N_116,In_1960,In_485);
and U117 (N_117,In_567,In_804);
and U118 (N_118,In_1248,In_1161);
or U119 (N_119,In_1099,In_308);
nor U120 (N_120,In_1869,In_307);
xor U121 (N_121,In_888,In_299);
nand U122 (N_122,In_409,In_1705);
nand U123 (N_123,In_860,In_960);
nand U124 (N_124,In_1366,In_454);
xnor U125 (N_125,In_566,In_1457);
or U126 (N_126,In_891,In_25);
and U127 (N_127,In_1272,In_1726);
nand U128 (N_128,In_31,In_315);
xor U129 (N_129,In_337,In_934);
nor U130 (N_130,In_1179,In_1762);
nor U131 (N_131,In_1370,In_973);
nor U132 (N_132,In_1444,In_294);
and U133 (N_133,In_141,In_456);
xnor U134 (N_134,In_1016,In_224);
xnor U135 (N_135,In_1924,In_527);
or U136 (N_136,In_1724,In_1355);
and U137 (N_137,In_822,In_1033);
or U138 (N_138,In_1675,In_234);
xor U139 (N_139,In_608,In_1054);
or U140 (N_140,In_1159,In_1630);
xnor U141 (N_141,In_1199,In_1832);
xor U142 (N_142,In_1496,In_652);
or U143 (N_143,In_1645,In_367);
xnor U144 (N_144,In_649,In_1835);
nand U145 (N_145,In_1777,In_1499);
or U146 (N_146,In_1656,In_589);
and U147 (N_147,In_86,In_1542);
xnor U148 (N_148,In_1729,In_1443);
nor U149 (N_149,In_1644,In_1312);
or U150 (N_150,In_266,In_441);
and U151 (N_151,In_1459,In_1322);
or U152 (N_152,In_1368,In_354);
xnor U153 (N_153,In_686,In_532);
and U154 (N_154,In_1242,In_1012);
and U155 (N_155,In_1549,In_993);
xor U156 (N_156,In_295,In_1091);
or U157 (N_157,In_1019,In_1658);
nor U158 (N_158,In_1109,In_215);
nand U159 (N_159,In_1816,In_335);
nor U160 (N_160,In_625,In_1600);
nand U161 (N_161,In_89,In_1428);
nor U162 (N_162,In_1978,In_467);
and U163 (N_163,In_348,In_1905);
or U164 (N_164,In_484,In_1489);
nor U165 (N_165,In_1912,In_476);
nand U166 (N_166,In_1748,In_1083);
or U167 (N_167,In_1105,In_921);
xnor U168 (N_168,In_1359,In_143);
xnor U169 (N_169,In_387,In_926);
xor U170 (N_170,In_1350,In_850);
nor U171 (N_171,In_1919,In_800);
and U172 (N_172,In_645,In_638);
nor U173 (N_173,In_1509,In_1559);
nor U174 (N_174,In_946,In_1169);
and U175 (N_175,In_1048,In_139);
and U176 (N_176,In_1649,In_1653);
nor U177 (N_177,In_1771,In_1634);
nor U178 (N_178,In_121,In_70);
nor U179 (N_179,In_1632,In_1246);
or U180 (N_180,In_203,In_575);
nand U181 (N_181,In_474,In_1856);
xnor U182 (N_182,In_1841,In_570);
nand U183 (N_183,In_257,In_986);
xor U184 (N_184,In_1531,In_344);
or U185 (N_185,In_410,In_95);
nand U186 (N_186,In_157,In_293);
nor U187 (N_187,In_48,In_935);
xor U188 (N_188,In_947,In_429);
and U189 (N_189,In_1041,In_866);
nand U190 (N_190,In_554,In_809);
nor U191 (N_191,In_1333,In_1439);
or U192 (N_192,In_1381,In_985);
nor U193 (N_193,In_746,In_1330);
and U194 (N_194,In_108,In_910);
nand U195 (N_195,In_526,In_1519);
nor U196 (N_196,In_966,In_1845);
xnor U197 (N_197,In_1598,In_1445);
nor U198 (N_198,In_1281,In_469);
or U199 (N_199,In_1674,In_1959);
nand U200 (N_200,In_832,In_1946);
and U201 (N_201,In_1077,In_975);
and U202 (N_202,In_1763,In_238);
xor U203 (N_203,In_1002,In_1976);
and U204 (N_204,In_324,In_1187);
or U205 (N_205,In_149,In_1948);
and U206 (N_206,In_1575,In_10);
nor U207 (N_207,In_1725,In_1815);
or U208 (N_208,In_1931,In_844);
or U209 (N_209,In_1172,In_1200);
and U210 (N_210,In_480,In_104);
or U211 (N_211,In_584,In_1515);
xnor U212 (N_212,In_976,In_607);
and U213 (N_213,In_719,In_646);
xor U214 (N_214,In_1926,In_1498);
nor U215 (N_215,In_784,In_1718);
nor U216 (N_216,In_1753,In_1430);
nor U217 (N_217,In_1446,In_1523);
nand U218 (N_218,In_1470,In_1024);
xnor U219 (N_219,In_248,In_1233);
and U220 (N_220,In_902,In_1174);
nand U221 (N_221,In_1136,In_460);
or U222 (N_222,In_655,In_131);
or U223 (N_223,In_342,In_53);
and U224 (N_224,In_823,In_537);
nand U225 (N_225,In_209,In_1928);
xnor U226 (N_226,In_1141,In_1098);
nor U227 (N_227,In_404,In_892);
nand U228 (N_228,In_1282,In_1838);
and U229 (N_229,In_217,In_962);
and U230 (N_230,In_19,In_1416);
nor U231 (N_231,In_936,In_1638);
xor U232 (N_232,In_1842,In_895);
and U233 (N_233,In_1721,In_97);
xor U234 (N_234,In_1032,In_1728);
nor U235 (N_235,In_1167,In_1999);
or U236 (N_236,In_464,In_969);
xor U237 (N_237,In_759,In_1637);
nand U238 (N_238,In_1794,In_1197);
xnor U239 (N_239,In_101,In_1025);
xor U240 (N_240,In_300,In_1567);
nor U241 (N_241,In_1119,In_325);
nor U242 (N_242,In_289,In_1920);
nand U243 (N_243,In_193,In_818);
nor U244 (N_244,In_610,In_1146);
nand U245 (N_245,In_285,In_1749);
or U246 (N_246,In_0,In_1615);
xnor U247 (N_247,In_1400,In_1042);
or U248 (N_248,In_1731,In_1453);
and U249 (N_249,In_578,In_1613);
and U250 (N_250,In_828,In_159);
xnor U251 (N_251,In_924,In_794);
nor U252 (N_252,In_1035,In_243);
nand U253 (N_253,In_1448,In_1142);
or U254 (N_254,In_1260,In_1932);
or U255 (N_255,In_1536,In_1252);
nand U256 (N_256,In_373,In_620);
or U257 (N_257,In_35,In_1129);
and U258 (N_258,In_368,In_1064);
and U259 (N_259,In_1538,In_750);
nand U260 (N_260,In_657,In_1641);
and U261 (N_261,In_1831,In_582);
nor U262 (N_262,In_436,In_1647);
nand U263 (N_263,In_893,In_1433);
xor U264 (N_264,In_1456,In_282);
and U265 (N_265,In_580,In_1053);
nor U266 (N_266,In_1402,In_717);
and U267 (N_267,In_1507,In_1399);
xor U268 (N_268,In_703,In_1766);
and U269 (N_269,In_774,In_1238);
or U270 (N_270,In_397,In_183);
and U271 (N_271,In_1481,In_1894);
nand U272 (N_272,In_298,In_1697);
nand U273 (N_273,In_1198,In_17);
nand U274 (N_274,In_78,In_636);
or U275 (N_275,In_359,In_639);
nor U276 (N_276,In_425,In_381);
nor U277 (N_277,In_504,In_953);
or U278 (N_278,In_1903,In_1533);
nor U279 (N_279,In_870,In_1361);
nand U280 (N_280,In_1052,In_59);
nor U281 (N_281,In_1236,In_653);
nor U282 (N_282,In_1933,In_1524);
xor U283 (N_283,In_956,In_1093);
or U284 (N_284,In_278,In_863);
or U285 (N_285,In_147,In_1138);
xnor U286 (N_286,In_455,In_1195);
xor U287 (N_287,In_1396,In_477);
nand U288 (N_288,In_1648,In_1689);
nand U289 (N_289,In_1810,In_1930);
nand U290 (N_290,In_847,In_1422);
xnor U291 (N_291,In_498,In_1935);
xnor U292 (N_292,In_350,In_1365);
nor U293 (N_293,In_585,In_268);
xor U294 (N_294,In_173,In_333);
nand U295 (N_295,In_112,In_1264);
xnor U296 (N_296,In_68,In_1547);
xor U297 (N_297,In_279,In_594);
nand U298 (N_298,In_711,In_450);
nor U299 (N_299,In_1225,In_357);
nor U300 (N_300,In_1971,In_1337);
xnor U301 (N_301,In_246,In_1384);
xnor U302 (N_302,In_1631,In_1230);
and U303 (N_303,In_916,In_1390);
and U304 (N_304,In_1377,In_1995);
and U305 (N_305,In_1194,In_24);
nor U306 (N_306,In_14,In_58);
xor U307 (N_307,In_1254,In_958);
nand U308 (N_308,In_812,In_1078);
or U309 (N_309,In_1898,In_286);
or U310 (N_310,In_328,In_72);
nand U311 (N_311,In_1879,In_792);
or U312 (N_312,In_922,In_525);
nand U313 (N_313,In_44,In_127);
xnor U314 (N_314,In_1274,In_1692);
and U315 (N_315,In_782,In_1759);
xor U316 (N_316,In_1944,In_1235);
nor U317 (N_317,In_1984,In_1349);
or U318 (N_318,In_1124,In_1802);
or U319 (N_319,In_319,In_71);
and U320 (N_320,In_290,In_1351);
xnor U321 (N_321,In_1412,In_1510);
or U322 (N_322,In_136,In_1503);
or U323 (N_323,In_1385,In_1202);
nand U324 (N_324,In_1405,In_1309);
xnor U325 (N_325,In_1571,In_1781);
nand U326 (N_326,In_842,In_1011);
or U327 (N_327,In_959,In_6);
nand U328 (N_328,In_1038,In_1699);
or U329 (N_329,In_1302,In_1543);
xor U330 (N_330,In_1353,In_1626);
and U331 (N_331,In_1421,In_827);
nor U332 (N_332,In_1261,In_1711);
or U333 (N_333,In_1911,In_881);
and U334 (N_334,In_494,In_292);
and U335 (N_335,In_145,In_374);
or U336 (N_336,In_1537,In_346);
xnor U337 (N_337,In_1642,In_770);
nand U338 (N_338,In_1867,In_621);
xnor U339 (N_339,In_631,In_789);
nor U340 (N_340,In_40,In_230);
xnor U341 (N_341,In_1226,In_1121);
or U342 (N_342,In_1015,In_1830);
nor U343 (N_343,In_523,In_1602);
or U344 (N_344,In_1266,In_852);
or U345 (N_345,In_214,In_1321);
and U346 (N_346,In_187,In_1208);
or U347 (N_347,In_1625,In_1676);
or U348 (N_348,In_617,In_1149);
and U349 (N_349,In_1994,In_803);
nor U350 (N_350,In_647,In_1378);
or U351 (N_351,In_1715,In_2);
and U352 (N_352,In_3,In_1908);
nand U353 (N_353,In_760,In_1916);
or U354 (N_354,In_559,In_119);
xnor U355 (N_355,In_1918,In_1082);
nand U356 (N_356,In_130,In_1278);
or U357 (N_357,In_1892,In_937);
and U358 (N_358,In_761,In_534);
xnor U359 (N_359,In_679,In_1750);
nor U360 (N_360,In_326,In_87);
nor U361 (N_361,In_763,In_125);
and U362 (N_362,In_13,In_398);
or U363 (N_363,In_694,In_501);
nor U364 (N_364,In_1822,In_1722);
and U365 (N_365,In_1983,In_1680);
xor U366 (N_366,In_443,In_1154);
or U367 (N_367,In_514,In_1849);
nor U368 (N_368,In_1318,In_1629);
nand U369 (N_369,In_689,In_854);
or U370 (N_370,In_994,In_1686);
nor U371 (N_371,In_1992,In_74);
or U372 (N_372,In_876,In_1868);
or U373 (N_373,In_757,In_744);
nand U374 (N_374,In_170,In_1097);
nand U375 (N_375,In_1371,In_383);
xor U376 (N_376,In_1606,In_1859);
xor U377 (N_377,In_999,In_29);
nand U378 (N_378,In_195,In_941);
or U379 (N_379,In_948,In_507);
nor U380 (N_380,In_63,In_1807);
or U381 (N_381,In_831,In_1591);
xnor U382 (N_382,In_1224,In_403);
nand U383 (N_383,In_1432,In_1819);
xnor U384 (N_384,In_1323,In_1331);
and U385 (N_385,In_1847,In_1655);
xor U386 (N_386,In_1601,In_1031);
nand U387 (N_387,In_561,In_982);
nand U388 (N_388,In_1391,In_496);
and U389 (N_389,In_666,In_297);
or U390 (N_390,In_465,In_685);
and U391 (N_391,In_1938,In_1335);
and U392 (N_392,In_1921,In_1808);
or U393 (N_393,In_204,In_683);
xor U394 (N_394,In_1395,In_493);
and U395 (N_395,In_416,In_156);
or U396 (N_396,In_1477,In_424);
xnor U397 (N_397,In_164,In_597);
or U398 (N_398,In_1247,In_388);
and U399 (N_399,In_1043,In_1511);
xnor U400 (N_400,In_543,In_1345);
nor U401 (N_401,In_392,In_406);
nor U402 (N_402,In_380,In_152);
nand U403 (N_403,In_968,In_1425);
nor U404 (N_404,In_1411,In_524);
nand U405 (N_405,In_178,In_1279);
xnor U406 (N_406,In_431,In_1184);
and U407 (N_407,In_252,In_1770);
or U408 (N_408,In_558,In_1881);
xnor U409 (N_409,In_1691,In_1348);
xor U410 (N_410,In_1752,In_670);
and U411 (N_411,In_1463,In_1914);
nand U412 (N_412,In_1840,In_176);
nand U413 (N_413,In_509,In_731);
or U414 (N_414,In_944,In_1572);
nand U415 (N_415,In_1501,In_950);
and U416 (N_416,In_1394,In_423);
or U417 (N_417,In_210,In_1186);
xor U418 (N_418,In_641,In_49);
nand U419 (N_419,In_1541,In_1901);
nand U420 (N_420,In_624,In_244);
xor U421 (N_421,In_1305,In_1525);
nand U422 (N_422,In_899,In_884);
and U423 (N_423,In_1191,In_36);
and U424 (N_424,In_26,In_1222);
nor U425 (N_425,In_879,In_1640);
nor U426 (N_426,In_415,In_723);
and U427 (N_427,In_309,In_438);
or U428 (N_428,In_1442,In_629);
xor U429 (N_429,In_577,In_236);
xor U430 (N_430,In_1380,In_1267);
nand U431 (N_431,In_188,In_1427);
or U432 (N_432,In_227,In_1044);
nand U433 (N_433,In_1423,In_506);
nor U434 (N_434,In_385,In_1825);
and U435 (N_435,In_742,In_851);
nand U436 (N_436,In_1756,In_845);
and U437 (N_437,In_1660,In_91);
and U438 (N_438,In_1410,In_1864);
nand U439 (N_439,In_1404,In_726);
or U440 (N_440,In_829,In_312);
nand U441 (N_441,In_7,In_1673);
nand U442 (N_442,In_1165,In_231);
nand U443 (N_443,In_1047,In_665);
xnor U444 (N_444,In_1296,In_1307);
xor U445 (N_445,In_730,In_1871);
nand U446 (N_446,In_1990,In_9);
and U447 (N_447,In_274,In_857);
and U448 (N_448,In_1621,In_1954);
nor U449 (N_449,In_778,In_417);
or U450 (N_450,In_1215,In_47);
or U451 (N_451,In_1364,In_681);
and U452 (N_452,In_277,In_637);
or U453 (N_453,In_725,In_1732);
xnor U454 (N_454,In_1545,In_1004);
or U455 (N_455,In_1848,In_932);
nor U456 (N_456,In_284,In_613);
nor U457 (N_457,In_199,In_262);
xnor U458 (N_458,In_595,In_733);
xnor U459 (N_459,In_1500,In_1672);
nor U460 (N_460,In_1843,In_1688);
xor U461 (N_461,In_1299,In_1356);
and U462 (N_462,In_1270,In_184);
and U463 (N_463,In_1034,In_654);
and U464 (N_464,In_1603,In_978);
or U465 (N_465,In_1627,In_739);
nor U466 (N_466,In_1593,In_107);
xor U467 (N_467,In_732,In_444);
nand U468 (N_468,In_1426,In_702);
nor U469 (N_469,In_1455,In_1107);
nand U470 (N_470,In_30,In_1682);
nor U471 (N_471,In_1112,In_898);
xnor U472 (N_472,In_1341,In_386);
or U473 (N_473,In_618,In_1461);
and U474 (N_474,In_1982,In_1592);
and U475 (N_475,In_198,In_1160);
xnor U476 (N_476,In_106,In_797);
and U477 (N_477,In_1565,In_1839);
and U478 (N_478,In_352,In_1363);
and U479 (N_479,In_1397,In_1492);
and U480 (N_480,In_316,In_890);
nand U481 (N_481,In_1028,In_1624);
or U482 (N_482,In_642,In_773);
or U483 (N_483,In_1857,In_1720);
or U484 (N_484,In_1434,In_788);
and U485 (N_485,In_1409,In_1162);
nand U486 (N_486,In_313,In_755);
or U487 (N_487,In_520,In_370);
nor U488 (N_488,In_232,In_1114);
nand U489 (N_489,In_1214,In_1128);
nand U490 (N_490,In_564,In_206);
and U491 (N_491,In_1407,In_1618);
nand U492 (N_492,In_497,In_998);
nand U493 (N_493,In_327,In_1890);
xor U494 (N_494,In_627,In_775);
and U495 (N_495,In_834,In_1595);
or U496 (N_496,In_1285,In_1981);
xnor U497 (N_497,In_824,In_1824);
nor U498 (N_498,In_673,In_154);
nand U499 (N_499,In_1558,In_604);
or U500 (N_500,In_671,In_682);
nor U501 (N_501,In_545,In_1180);
or U502 (N_502,In_806,In_1227);
or U503 (N_503,In_780,In_22);
nand U504 (N_504,In_355,In_171);
nand U505 (N_505,In_615,In_1204);
nand U506 (N_506,In_43,In_877);
xor U507 (N_507,In_1229,In_271);
nand U508 (N_508,In_1910,In_1555);
nor U509 (N_509,In_1873,In_1374);
and U510 (N_510,In_1369,In_263);
and U511 (N_511,In_1520,In_706);
or U512 (N_512,In_1166,In_1084);
nand U513 (N_513,In_1922,In_1219);
nand U514 (N_514,In_695,In_883);
and U515 (N_515,In_1135,In_419);
xnor U516 (N_516,In_1367,In_785);
and U517 (N_517,In_1561,In_1315);
and U518 (N_518,In_407,In_533);
or U519 (N_519,In_1468,In_1100);
or U520 (N_520,In_389,In_855);
and U521 (N_521,In_1962,In_1244);
or U522 (N_522,In_362,In_155);
or U523 (N_523,In_488,In_1424);
or U524 (N_524,In_276,In_989);
xnor U525 (N_525,In_169,In_1817);
nor U526 (N_526,In_1104,In_713);
and U527 (N_527,In_459,In_915);
nor U528 (N_528,In_1927,In_303);
nand U529 (N_529,In_1122,In_375);
nand U530 (N_530,In_1818,In_179);
nand U531 (N_531,In_1584,In_503);
nor U532 (N_532,In_556,In_1277);
xnor U533 (N_533,In_1139,In_1268);
nor U534 (N_534,In_250,In_979);
nand U535 (N_535,In_635,In_1059);
nand U536 (N_536,In_1452,In_751);
nand U537 (N_537,In_1472,In_1014);
xor U538 (N_538,In_192,In_1196);
xnor U539 (N_539,In_648,In_886);
and U540 (N_540,In_1737,In_320);
xnor U541 (N_541,In_603,In_667);
nor U542 (N_542,In_1783,In_1440);
or U543 (N_543,In_1714,In_317);
xor U544 (N_544,In_1258,In_1259);
nor U545 (N_545,In_728,In_1635);
and U546 (N_546,In_1570,In_1804);
and U547 (N_547,In_1563,In_1577);
nand U548 (N_548,In_1482,In_555);
or U549 (N_549,In_253,In_1177);
and U550 (N_550,In_64,In_990);
nor U551 (N_551,In_825,In_1089);
or U552 (N_552,In_837,In_1450);
nand U553 (N_553,In_1823,In_1583);
nand U554 (N_554,In_592,In_1679);
nor U555 (N_555,In_952,In_1293);
xor U556 (N_556,In_267,In_1079);
and U557 (N_557,In_288,In_1828);
nand U558 (N_558,In_205,In_889);
and U559 (N_559,In_1211,In_1067);
and U560 (N_560,In_668,In_628);
xnor U561 (N_561,In_1552,In_168);
xor U562 (N_562,In_1698,In_1294);
nand U563 (N_563,In_1223,In_1548);
or U564 (N_564,In_1956,In_1062);
and U565 (N_565,In_826,In_599);
nor U566 (N_566,In_283,In_901);
or U567 (N_567,In_967,In_661);
nand U568 (N_568,In_264,In_475);
and U569 (N_569,In_931,In_1280);
nor U570 (N_570,In_913,In_1474);
or U571 (N_571,In_1579,In_846);
xnor U572 (N_572,In_1408,In_1891);
or U573 (N_573,In_1306,In_402);
xnor U574 (N_574,In_1018,In_1557);
or U575 (N_575,In_172,In_914);
or U576 (N_576,In_1701,In_1508);
and U577 (N_577,In_366,In_1271);
and U578 (N_578,In_1005,In_220);
xor U579 (N_579,In_16,In_446);
xor U580 (N_580,In_1088,In_987);
and U581 (N_581,In_771,In_1253);
and U582 (N_582,In_1393,In_1487);
nor U583 (N_583,In_1576,In_1338);
and U584 (N_584,In_428,In_858);
nor U585 (N_585,In_1068,In_80);
or U586 (N_586,In_1473,In_161);
xor U587 (N_587,In_329,In_376);
or U588 (N_588,In_838,In_489);
nor U589 (N_589,In_1049,In_593);
or U590 (N_590,In_1784,In_1144);
nor U591 (N_591,In_301,In_124);
and U592 (N_592,In_468,In_820);
xnor U593 (N_593,In_1684,In_531);
xor U594 (N_594,In_207,In_1466);
xnor U595 (N_595,In_1106,In_1494);
or U596 (N_596,In_96,In_451);
nand U597 (N_597,In_132,In_1505);
and U598 (N_598,In_1693,In_1739);
and U599 (N_599,In_259,In_1546);
nand U600 (N_600,In_581,In_1788);
or U601 (N_601,In_1834,In_1733);
nor U602 (N_602,In_1566,In_664);
nor U603 (N_603,In_569,In_1010);
nand U604 (N_604,In_906,In_783);
and U605 (N_605,In_1801,In_1115);
xor U606 (N_606,In_219,In_737);
xor U607 (N_607,In_1964,In_1708);
and U608 (N_608,In_1778,In_614);
nand U609 (N_609,In_1875,In_1774);
xnor U610 (N_610,In_51,In_109);
nand U611 (N_611,In_1185,In_1934);
nand U612 (N_612,In_1564,In_1171);
xnor U613 (N_613,In_1961,In_1006);
or U614 (N_614,In_807,In_395);
nand U615 (N_615,In_449,In_1528);
and U616 (N_616,In_1590,In_1556);
nor U617 (N_617,In_700,In_1650);
nand U618 (N_618,In_571,In_1300);
nor U619 (N_619,In_1153,In_241);
nand U620 (N_620,In_596,In_1495);
and U621 (N_621,In_1147,In_1622);
nor U622 (N_622,In_810,In_323);
nand U623 (N_623,In_942,In_1574);
and U624 (N_624,In_1667,In_539);
or U625 (N_625,In_983,In_1646);
and U626 (N_626,In_716,In_517);
and U627 (N_627,In_634,In_1102);
xnor U628 (N_628,In_66,In_1140);
xor U629 (N_629,In_88,In_912);
xor U630 (N_630,In_1516,In_1730);
nand U631 (N_631,In_433,In_709);
nor U632 (N_632,In_391,In_369);
xnor U633 (N_633,In_992,In_1437);
xnor U634 (N_634,In_27,In_1449);
nand U635 (N_635,In_736,In_767);
xnor U636 (N_636,In_1544,In_1465);
xor U637 (N_637,In_1469,In_995);
xor U638 (N_638,In_1560,In_81);
nor U639 (N_639,In_1118,In_1659);
nand U640 (N_640,In_50,In_466);
or U641 (N_641,In_688,In_1123);
nor U642 (N_642,In_439,In_1913);
nor U643 (N_643,In_1023,In_492);
and U644 (N_644,In_1915,In_69);
and U645 (N_645,In_587,In_1882);
nor U646 (N_646,In_1683,In_1540);
nand U647 (N_647,In_1289,In_1095);
and U648 (N_648,In_1851,In_1972);
and U649 (N_649,In_799,In_113);
and U650 (N_650,In_39,In_1387);
nand U651 (N_651,In_1878,In_1134);
nor U652 (N_652,In_90,In_1573);
xnor U653 (N_653,In_747,In_1373);
and U654 (N_654,In_457,In_904);
nor U655 (N_655,In_1799,In_1797);
nand U656 (N_656,In_1483,In_1094);
nor U657 (N_657,In_55,In_1485);
and U658 (N_658,In_868,In_1782);
xor U659 (N_659,In_1113,In_1313);
nand U660 (N_660,In_573,In_338);
or U661 (N_661,In_223,In_452);
xor U662 (N_662,In_1880,In_1295);
or U663 (N_663,In_1314,In_229);
or U664 (N_664,In_228,In_1532);
and U665 (N_665,In_1695,In_692);
xor U666 (N_666,In_1589,In_1490);
and U667 (N_667,In_77,In_1772);
nor U668 (N_668,In_1775,In_1677);
nor U669 (N_669,In_848,In_849);
xnor U670 (N_670,In_269,In_1803);
or U671 (N_671,In_1283,In_557);
nand U672 (N_672,In_122,In_482);
and U673 (N_673,In_486,In_343);
nand U674 (N_674,In_340,In_56);
or U675 (N_675,In_1255,In_781);
nor U676 (N_676,In_186,In_1923);
or U677 (N_677,In_1058,In_840);
nor U678 (N_678,In_118,In_221);
nand U679 (N_679,In_1288,In_1897);
or U680 (N_680,In_1716,In_353);
nor U681 (N_681,In_1967,In_927);
nand U682 (N_682,In_84,In_1761);
nor U683 (N_683,In_768,In_691);
xor U684 (N_684,In_260,In_1740);
nand U685 (N_685,In_769,In_1872);
nand U686 (N_686,In_1026,In_111);
or U687 (N_687,In_1241,In_371);
nor U688 (N_688,In_1401,In_1707);
or U689 (N_689,In_1096,In_721);
or U690 (N_690,In_41,In_552);
nor U691 (N_691,In_413,In_611);
and U692 (N_692,In_1334,In_1506);
nor U693 (N_693,In_1462,In_548);
nand U694 (N_694,In_110,In_129);
and U695 (N_695,In_1029,In_1310);
and U696 (N_696,In_1205,In_535);
and U697 (N_697,In_616,In_1998);
and U698 (N_698,In_1604,In_856);
xor U699 (N_699,In_1866,In_1654);
and U700 (N_700,In_530,In_165);
nand U701 (N_701,In_160,In_1076);
nand U702 (N_702,In_1175,In_254);
and U703 (N_703,In_588,In_1081);
or U704 (N_704,In_1917,In_1989);
and U705 (N_705,In_393,In_1623);
and U706 (N_706,In_518,In_1190);
xor U707 (N_707,In_1120,In_177);
or U708 (N_708,In_82,In_430);
nor U709 (N_709,In_1888,In_669);
or U710 (N_710,In_819,In_358);
nand U711 (N_711,In_1968,In_21);
nand U712 (N_712,In_676,In_776);
nand U713 (N_713,In_1158,In_1970);
or U714 (N_714,In_1940,In_1320);
nand U715 (N_715,In_1037,In_1787);
nor U716 (N_716,In_553,In_1806);
or U717 (N_717,In_678,In_1986);
or U718 (N_718,In_871,In_626);
nor U719 (N_719,In_754,In_1965);
nand U720 (N_720,In_1389,In_1001);
nor U721 (N_721,In_1757,In_1311);
or U722 (N_722,In_83,In_1020);
and U723 (N_723,In_1431,In_408);
nand U724 (N_724,In_458,In_777);
or U725 (N_725,In_1170,In_1231);
nor U726 (N_726,In_698,In_361);
nor U727 (N_727,In_1661,In_1414);
xor U728 (N_728,In_516,In_378);
nand U729 (N_729,In_1308,In_772);
nand U730 (N_730,In_749,In_1497);
or U731 (N_731,In_60,In_1885);
nand U732 (N_732,In_339,In_1398);
nand U733 (N_733,In_37,In_574);
and U734 (N_734,In_1286,In_562);
nor U735 (N_735,In_1319,In_1249);
and U736 (N_736,In_1529,In_1747);
xnor U737 (N_737,In_1827,In_1657);
or U738 (N_738,In_1275,In_1145);
xnor U739 (N_739,In_1789,In_528);
nor U740 (N_740,In_1779,In_1009);
xor U741 (N_741,In_23,In_1504);
nor U742 (N_742,In_1007,In_218);
nor U743 (N_743,In_1663,In_148);
and U744 (N_744,In_1793,In_1116);
nor U745 (N_745,In_1850,In_306);
nor U746 (N_746,In_965,In_512);
or U747 (N_747,In_1130,In_1985);
nor U748 (N_748,In_1022,In_128);
xor U749 (N_749,In_1447,In_1760);
or U750 (N_750,In_576,In_963);
nand U751 (N_751,In_964,In_1619);
nor U752 (N_752,In_1213,In_1668);
nor U753 (N_753,In_563,In_930);
or U754 (N_754,In_382,In_519);
or U755 (N_755,In_302,In_1837);
or U756 (N_756,In_1,In_163);
xnor U757 (N_757,In_1860,In_872);
nand U758 (N_758,In_38,In_705);
nor U759 (N_759,In_1150,In_1332);
and U760 (N_760,In_1417,In_153);
nor U761 (N_761,In_1773,In_99);
nand U762 (N_762,In_1829,In_1003);
and U763 (N_763,In_1324,In_411);
nand U764 (N_764,In_123,In_853);
or U765 (N_765,In_1620,In_1792);
and U766 (N_766,In_1436,In_334);
or U767 (N_767,In_1896,In_1786);
xor U768 (N_768,In_1352,In_1568);
nand U769 (N_769,In_1738,In_1585);
or U770 (N_770,In_714,In_1388);
and U771 (N_771,In_1220,In_1925);
xor U772 (N_772,In_1550,In_1876);
and U773 (N_773,In_1240,In_448);
xnor U774 (N_774,In_791,In_240);
xor U775 (N_775,In_180,In_1125);
and U776 (N_776,In_938,In_1734);
xnor U777 (N_777,In_623,In_1735);
nand U778 (N_778,In_212,In_727);
or U779 (N_779,In_1768,In_1063);
nor U780 (N_780,In_830,In_1243);
and U781 (N_781,In_798,In_590);
nand U782 (N_782,In_158,In_1471);
and U783 (N_783,In_364,In_510);
nand U784 (N_784,In_1269,In_1800);
nor U785 (N_785,In_805,In_900);
xor U786 (N_786,In_1833,In_1936);
or U787 (N_787,In_1937,In_1406);
and U788 (N_788,In_542,In_1303);
nor U789 (N_789,In_247,In_1751);
or U790 (N_790,In_196,In_137);
or U791 (N_791,In_802,In_1074);
or U792 (N_792,In_93,In_1251);
nor U793 (N_793,In_674,In_296);
nor U794 (N_794,In_508,In_622);
or U795 (N_795,In_640,In_18);
xor U796 (N_796,In_1517,In_1951);
xor U797 (N_797,In_1117,In_909);
nor U798 (N_798,In_748,In_190);
or U799 (N_799,In_151,In_1127);
and U800 (N_800,In_1111,In_76);
xnor U801 (N_801,In_841,In_743);
and U802 (N_802,In_1706,In_1435);
xor U803 (N_803,In_134,In_633);
or U804 (N_804,In_336,In_715);
nand U805 (N_805,In_835,In_1594);
nor U806 (N_806,In_981,In_1478);
and U807 (N_807,In_67,In_764);
xor U808 (N_808,In_1743,In_487);
and U809 (N_809,In_762,In_786);
nand U810 (N_810,In_1767,In_1991);
or U811 (N_811,In_911,In_45);
or U812 (N_812,In_710,In_1382);
or U813 (N_813,In_1796,In_1717);
nor U814 (N_814,In_1221,In_1475);
xor U815 (N_815,In_1346,In_843);
or U816 (N_816,In_1671,In_560);
xor U817 (N_817,In_445,In_57);
and U818 (N_818,In_598,In_1758);
xor U819 (N_819,In_606,In_1188);
and U820 (N_820,In_400,In_1974);
and U821 (N_821,In_955,In_859);
and U822 (N_822,In_1192,In_1479);
xor U823 (N_823,In_1297,In_1805);
nand U824 (N_824,In_1943,In_974);
nand U825 (N_825,In_1316,In_1929);
and U826 (N_826,In_256,In_704);
nand U827 (N_827,In_540,In_1958);
nor U828 (N_828,In_479,In_1534);
nand U829 (N_829,In_1336,In_875);
nor U830 (N_830,In_1080,In_1973);
nand U831 (N_831,In_1844,In_1949);
xnor U832 (N_832,In_515,In_536);
nor U833 (N_833,In_1764,In_1291);
xor U834 (N_834,In_765,In_216);
or U835 (N_835,In_1662,In_305);
nor U836 (N_836,In_140,In_304);
and U837 (N_837,In_1212,In_660);
nand U838 (N_838,In_1909,In_94);
nor U839 (N_839,In_322,In_461);
and U840 (N_840,In_191,In_1292);
or U841 (N_841,In_1535,In_473);
xnor U842 (N_842,In_341,In_756);
or U843 (N_843,In_142,In_619);
xor U844 (N_844,In_1609,In_1317);
nor U845 (N_845,In_34,In_795);
nor U846 (N_846,In_1854,In_1605);
nand U847 (N_847,In_412,In_522);
nor U848 (N_848,In_1617,In_1403);
and U849 (N_849,In_347,In_1610);
nor U850 (N_850,In_708,In_1132);
or U851 (N_851,In_211,In_1975);
and U852 (N_852,In_1290,In_591);
nor U853 (N_853,In_85,In_787);
nand U854 (N_854,In_1057,In_363);
nor U855 (N_855,In_817,In_1484);
nand U856 (N_856,In_1950,In_672);
xor U857 (N_857,In_1342,In_970);
or U858 (N_858,In_1870,In_793);
or U859 (N_859,In_440,In_766);
nor U860 (N_860,In_32,In_897);
xor U861 (N_861,In_33,In_360);
nor U862 (N_862,In_310,In_435);
xor U863 (N_863,In_925,In_996);
nand U864 (N_864,In_1046,In_42);
nor U865 (N_865,In_1438,In_437);
nor U866 (N_866,In_939,In_427);
and U867 (N_867,In_940,In_1000);
nor U868 (N_868,In_4,In_126);
and U869 (N_869,In_1108,In_1696);
and U870 (N_870,In_471,In_1178);
nand U871 (N_871,In_270,In_1553);
nor U872 (N_872,In_1703,In_720);
xnor U873 (N_873,In_314,In_249);
xnor U874 (N_874,In_758,In_801);
or U875 (N_875,In_1685,In_1284);
nor U876 (N_876,In_396,In_1580);
and U877 (N_877,In_1636,In_600);
xnor U878 (N_878,In_1027,In_954);
or U879 (N_879,In_917,In_1887);
nor U880 (N_880,In_864,In_1347);
nand U881 (N_881,In_135,In_779);
or U882 (N_882,In_265,In_862);
nor U883 (N_883,In_1263,In_1488);
and U884 (N_884,In_197,In_1900);
nand U885 (N_885,In_1085,In_1980);
and U886 (N_886,In_1813,In_873);
or U887 (N_887,In_1256,In_1358);
nand U888 (N_888,In_1493,In_1086);
nor U889 (N_889,In_929,In_908);
or U890 (N_890,In_1754,In_945);
xnor U891 (N_891,In_1218,In_1669);
nand U892 (N_892,In_632,In_920);
nor U893 (N_893,In_658,In_394);
nor U894 (N_894,In_690,In_1415);
xnor U895 (N_895,In_735,In_202);
and U896 (N_896,In_100,In_977);
xor U897 (N_897,In_878,In_1713);
and U898 (N_898,In_687,In_1736);
nor U899 (N_899,In_502,In_1327);
nor U900 (N_900,In_189,In_1582);
xor U901 (N_901,In_1791,In_1588);
xor U902 (N_902,In_495,In_1798);
or U903 (N_903,In_102,In_345);
and U904 (N_904,In_814,In_1670);
nor U905 (N_905,In_1996,In_1137);
or U906 (N_906,In_1616,In_650);
nor U907 (N_907,In_237,In_1746);
and U908 (N_908,In_1957,In_116);
or U909 (N_909,In_1210,In_311);
nand U910 (N_910,In_903,In_997);
or U911 (N_911,In_865,In_1467);
nand U912 (N_912,In_745,In_896);
nor U913 (N_913,In_677,In_138);
nand U914 (N_914,In_377,In_1392);
xnor U915 (N_915,In_718,In_511);
xor U916 (N_916,In_1216,In_696);
and U917 (N_917,In_724,In_432);
xnor U918 (N_918,In_928,In_1357);
nor U919 (N_919,In_1877,In_490);
nor U920 (N_920,In_242,In_811);
or U921 (N_921,In_583,In_287);
and U922 (N_922,In_1727,In_1379);
nor U923 (N_923,In_1865,In_1963);
and U924 (N_924,In_1596,In_521);
nand U925 (N_925,In_1587,In_453);
and U926 (N_926,In_1071,In_8);
or U927 (N_927,In_549,In_869);
xnor U928 (N_928,In_1776,In_462);
or U929 (N_929,In_1464,In_175);
nor U930 (N_930,In_1945,In_233);
nand U931 (N_931,In_1953,In_951);
nor U932 (N_932,In_426,In_1997);
xor U933 (N_933,In_174,In_1977);
or U934 (N_934,In_405,In_1539);
xnor U935 (N_935,In_1812,In_1173);
nor U936 (N_936,In_734,In_1329);
or U937 (N_937,In_1152,In_1372);
xor U938 (N_938,In_1785,In_1522);
or U939 (N_939,In_1710,In_1458);
nor U940 (N_940,In_1955,In_1326);
or U941 (N_941,In_1821,In_1451);
and U942 (N_942,In_1021,In_162);
nor U943 (N_943,In_166,In_1723);
or U944 (N_944,In_1889,In_1895);
nand U945 (N_945,In_602,In_61);
xnor U946 (N_946,In_1614,In_291);
or U947 (N_947,In_586,In_544);
or U948 (N_948,In_1993,In_1155);
xor U949 (N_949,In_332,In_722);
nand U950 (N_950,In_1611,In_258);
xnor U951 (N_951,In_1639,In_907);
xnor U952 (N_952,In_874,In_1126);
nand U953 (N_953,In_422,In_1855);
and U954 (N_954,In_752,In_1051);
xnor U955 (N_955,In_1664,In_1704);
and U956 (N_956,In_1090,In_1339);
or U957 (N_957,In_643,In_208);
nor U958 (N_958,In_1413,In_150);
xor U959 (N_959,In_1040,In_226);
or U960 (N_960,In_693,In_972);
and U961 (N_961,In_1110,In_280);
and U962 (N_962,In_1419,In_1893);
xor U963 (N_963,In_1987,In_12);
xor U964 (N_964,In_894,In_1386);
xor U965 (N_965,In_943,In_836);
nand U966 (N_966,In_753,In_1050);
nor U967 (N_967,In_659,In_1207);
nor U968 (N_968,In_1527,In_1551);
xnor U969 (N_969,In_28,In_546);
and U970 (N_970,In_1036,In_1234);
and U971 (N_971,In_923,In_1952);
or U972 (N_972,In_699,In_1651);
nor U973 (N_973,In_1418,In_1628);
and U974 (N_974,In_572,In_547);
nor U975 (N_975,In_167,In_120);
nor U976 (N_976,In_1979,In_73);
nand U977 (N_977,In_62,In_251);
nand U978 (N_978,In_816,In_463);
or U979 (N_979,In_984,In_991);
xor U980 (N_980,In_239,In_1678);
nand U981 (N_981,In_330,In_513);
nor U982 (N_982,In_1709,In_1569);
nand U983 (N_983,In_1526,In_54);
nand U984 (N_984,In_1203,In_1176);
nor U985 (N_985,In_1151,In_808);
and U986 (N_986,In_272,In_1070);
or U987 (N_987,In_201,In_351);
nand U988 (N_988,In_1883,In_384);
xor U989 (N_989,In_1712,In_1343);
and U990 (N_990,In_729,In_1809);
xor U991 (N_991,In_1906,In_1045);
or U992 (N_992,In_1862,In_401);
or U993 (N_993,In_1148,In_1633);
and U994 (N_994,In_961,In_1420);
nand U995 (N_995,In_1780,In_1744);
nor U996 (N_996,In_1795,In_1755);
nand U997 (N_997,In_225,In_796);
nor U998 (N_998,In_1157,In_1702);
nor U999 (N_999,In_1514,In_1907);
xor U1000 (N_1000,In_1807,In_1565);
nand U1001 (N_1001,In_324,In_1162);
nand U1002 (N_1002,In_616,In_58);
or U1003 (N_1003,In_1070,In_121);
nor U1004 (N_1004,In_890,In_1431);
nand U1005 (N_1005,In_671,In_668);
xnor U1006 (N_1006,In_473,In_197);
nor U1007 (N_1007,In_1260,In_1980);
and U1008 (N_1008,In_1793,In_755);
or U1009 (N_1009,In_768,In_1279);
nand U1010 (N_1010,In_950,In_51);
and U1011 (N_1011,In_1026,In_440);
xnor U1012 (N_1012,In_927,In_1138);
nor U1013 (N_1013,In_1918,In_271);
nor U1014 (N_1014,In_1939,In_864);
nor U1015 (N_1015,In_572,In_503);
and U1016 (N_1016,In_1121,In_1677);
and U1017 (N_1017,In_1016,In_1482);
and U1018 (N_1018,In_850,In_987);
or U1019 (N_1019,In_651,In_1862);
or U1020 (N_1020,In_844,In_1472);
xor U1021 (N_1021,In_511,In_1159);
nor U1022 (N_1022,In_923,In_613);
nand U1023 (N_1023,In_45,In_867);
nand U1024 (N_1024,In_99,In_1934);
xnor U1025 (N_1025,In_499,In_990);
and U1026 (N_1026,In_516,In_1349);
nor U1027 (N_1027,In_1588,In_688);
and U1028 (N_1028,In_477,In_1210);
or U1029 (N_1029,In_1035,In_150);
nand U1030 (N_1030,In_1442,In_178);
nand U1031 (N_1031,In_235,In_409);
xnor U1032 (N_1032,In_1296,In_1441);
nand U1033 (N_1033,In_1463,In_199);
and U1034 (N_1034,In_1001,In_1956);
xor U1035 (N_1035,In_1268,In_482);
and U1036 (N_1036,In_1440,In_363);
nand U1037 (N_1037,In_457,In_365);
nand U1038 (N_1038,In_491,In_1173);
nand U1039 (N_1039,In_1180,In_508);
nand U1040 (N_1040,In_1227,In_125);
or U1041 (N_1041,In_305,In_1669);
xnor U1042 (N_1042,In_253,In_1681);
nand U1043 (N_1043,In_41,In_250);
and U1044 (N_1044,In_149,In_548);
nand U1045 (N_1045,In_460,In_1729);
or U1046 (N_1046,In_1218,In_1633);
xor U1047 (N_1047,In_389,In_55);
nor U1048 (N_1048,In_1065,In_1606);
nand U1049 (N_1049,In_102,In_1378);
or U1050 (N_1050,In_1929,In_235);
and U1051 (N_1051,In_887,In_544);
xnor U1052 (N_1052,In_1018,In_35);
or U1053 (N_1053,In_144,In_1428);
nand U1054 (N_1054,In_726,In_692);
nand U1055 (N_1055,In_194,In_704);
nand U1056 (N_1056,In_918,In_897);
and U1057 (N_1057,In_756,In_1928);
and U1058 (N_1058,In_773,In_825);
xor U1059 (N_1059,In_1459,In_17);
and U1060 (N_1060,In_1326,In_1737);
xnor U1061 (N_1061,In_604,In_1220);
and U1062 (N_1062,In_448,In_1142);
nor U1063 (N_1063,In_1420,In_295);
xnor U1064 (N_1064,In_1412,In_860);
xnor U1065 (N_1065,In_1870,In_797);
xnor U1066 (N_1066,In_307,In_1011);
or U1067 (N_1067,In_796,In_489);
nor U1068 (N_1068,In_947,In_551);
xnor U1069 (N_1069,In_1002,In_1491);
and U1070 (N_1070,In_972,In_1765);
and U1071 (N_1071,In_1395,In_1016);
nor U1072 (N_1072,In_79,In_793);
or U1073 (N_1073,In_1367,In_237);
xor U1074 (N_1074,In_180,In_557);
xor U1075 (N_1075,In_2,In_1171);
nor U1076 (N_1076,In_223,In_381);
or U1077 (N_1077,In_1029,In_1488);
nor U1078 (N_1078,In_1749,In_1730);
xor U1079 (N_1079,In_1850,In_920);
nor U1080 (N_1080,In_1004,In_1241);
or U1081 (N_1081,In_1971,In_1692);
nor U1082 (N_1082,In_1406,In_1217);
or U1083 (N_1083,In_1221,In_759);
xnor U1084 (N_1084,In_317,In_575);
or U1085 (N_1085,In_90,In_1006);
or U1086 (N_1086,In_1392,In_658);
and U1087 (N_1087,In_105,In_1658);
nor U1088 (N_1088,In_1357,In_1287);
and U1089 (N_1089,In_1714,In_1894);
nor U1090 (N_1090,In_1829,In_902);
nand U1091 (N_1091,In_1168,In_1265);
and U1092 (N_1092,In_1159,In_1460);
xnor U1093 (N_1093,In_1950,In_1066);
nand U1094 (N_1094,In_235,In_1576);
nand U1095 (N_1095,In_735,In_1571);
nand U1096 (N_1096,In_1017,In_191);
or U1097 (N_1097,In_363,In_1468);
or U1098 (N_1098,In_36,In_592);
xor U1099 (N_1099,In_1636,In_924);
and U1100 (N_1100,In_1253,In_1859);
and U1101 (N_1101,In_1621,In_52);
nand U1102 (N_1102,In_400,In_362);
nor U1103 (N_1103,In_712,In_841);
or U1104 (N_1104,In_936,In_1235);
or U1105 (N_1105,In_1455,In_940);
or U1106 (N_1106,In_607,In_264);
nor U1107 (N_1107,In_781,In_73);
nand U1108 (N_1108,In_1466,In_609);
xor U1109 (N_1109,In_364,In_1456);
and U1110 (N_1110,In_221,In_481);
and U1111 (N_1111,In_1762,In_714);
nor U1112 (N_1112,In_324,In_336);
nor U1113 (N_1113,In_1544,In_909);
xor U1114 (N_1114,In_830,In_1012);
or U1115 (N_1115,In_40,In_1685);
or U1116 (N_1116,In_975,In_978);
nor U1117 (N_1117,In_1225,In_780);
xnor U1118 (N_1118,In_195,In_1715);
nor U1119 (N_1119,In_1280,In_898);
or U1120 (N_1120,In_730,In_889);
or U1121 (N_1121,In_2,In_320);
nand U1122 (N_1122,In_150,In_390);
and U1123 (N_1123,In_487,In_709);
and U1124 (N_1124,In_621,In_959);
xnor U1125 (N_1125,In_1614,In_1379);
nor U1126 (N_1126,In_352,In_1423);
or U1127 (N_1127,In_1652,In_1492);
or U1128 (N_1128,In_109,In_174);
or U1129 (N_1129,In_1069,In_795);
and U1130 (N_1130,In_448,In_14);
nand U1131 (N_1131,In_526,In_194);
nor U1132 (N_1132,In_520,In_1515);
nand U1133 (N_1133,In_524,In_594);
nor U1134 (N_1134,In_896,In_991);
xor U1135 (N_1135,In_631,In_1648);
nand U1136 (N_1136,In_1902,In_905);
and U1137 (N_1137,In_1741,In_92);
or U1138 (N_1138,In_1941,In_730);
or U1139 (N_1139,In_783,In_1686);
nand U1140 (N_1140,In_1364,In_253);
xor U1141 (N_1141,In_1467,In_515);
nor U1142 (N_1142,In_551,In_1655);
or U1143 (N_1143,In_1916,In_1256);
xnor U1144 (N_1144,In_168,In_820);
nand U1145 (N_1145,In_1645,In_5);
or U1146 (N_1146,In_782,In_1159);
or U1147 (N_1147,In_367,In_1566);
and U1148 (N_1148,In_138,In_364);
xor U1149 (N_1149,In_167,In_407);
or U1150 (N_1150,In_1091,In_1372);
and U1151 (N_1151,In_1508,In_632);
or U1152 (N_1152,In_196,In_87);
xor U1153 (N_1153,In_1952,In_812);
xnor U1154 (N_1154,In_926,In_1134);
nor U1155 (N_1155,In_231,In_621);
or U1156 (N_1156,In_1569,In_1320);
xor U1157 (N_1157,In_389,In_1444);
and U1158 (N_1158,In_164,In_641);
and U1159 (N_1159,In_61,In_106);
or U1160 (N_1160,In_1488,In_1972);
nor U1161 (N_1161,In_1261,In_1445);
nand U1162 (N_1162,In_1574,In_1796);
nand U1163 (N_1163,In_1030,In_540);
nand U1164 (N_1164,In_1460,In_55);
xor U1165 (N_1165,In_1690,In_89);
xnor U1166 (N_1166,In_1215,In_755);
xor U1167 (N_1167,In_1662,In_107);
and U1168 (N_1168,In_377,In_852);
nor U1169 (N_1169,In_182,In_798);
and U1170 (N_1170,In_19,In_1352);
or U1171 (N_1171,In_1242,In_215);
xnor U1172 (N_1172,In_1898,In_856);
nor U1173 (N_1173,In_165,In_26);
nor U1174 (N_1174,In_321,In_101);
or U1175 (N_1175,In_243,In_276);
nand U1176 (N_1176,In_1565,In_1343);
nand U1177 (N_1177,In_1244,In_1064);
or U1178 (N_1178,In_1950,In_82);
nor U1179 (N_1179,In_788,In_1718);
nand U1180 (N_1180,In_1233,In_375);
or U1181 (N_1181,In_1142,In_1859);
xor U1182 (N_1182,In_894,In_1044);
and U1183 (N_1183,In_401,In_921);
nand U1184 (N_1184,In_652,In_1902);
nor U1185 (N_1185,In_1244,In_171);
xor U1186 (N_1186,In_1027,In_1252);
or U1187 (N_1187,In_422,In_605);
nor U1188 (N_1188,In_1605,In_1717);
or U1189 (N_1189,In_173,In_1385);
nor U1190 (N_1190,In_97,In_1912);
nor U1191 (N_1191,In_1044,In_1040);
nand U1192 (N_1192,In_579,In_330);
nor U1193 (N_1193,In_517,In_1890);
nor U1194 (N_1194,In_1399,In_886);
and U1195 (N_1195,In_1360,In_1246);
and U1196 (N_1196,In_647,In_1763);
nor U1197 (N_1197,In_1125,In_108);
or U1198 (N_1198,In_1795,In_1740);
xor U1199 (N_1199,In_1060,In_711);
and U1200 (N_1200,In_1687,In_834);
nand U1201 (N_1201,In_431,In_195);
and U1202 (N_1202,In_1882,In_1546);
xor U1203 (N_1203,In_1860,In_69);
and U1204 (N_1204,In_1684,In_592);
and U1205 (N_1205,In_847,In_1931);
and U1206 (N_1206,In_92,In_352);
nor U1207 (N_1207,In_317,In_708);
and U1208 (N_1208,In_29,In_301);
nor U1209 (N_1209,In_1867,In_1030);
xor U1210 (N_1210,In_477,In_511);
and U1211 (N_1211,In_1001,In_737);
and U1212 (N_1212,In_204,In_1252);
or U1213 (N_1213,In_883,In_1353);
xnor U1214 (N_1214,In_1134,In_348);
and U1215 (N_1215,In_1702,In_1344);
nor U1216 (N_1216,In_1417,In_113);
xor U1217 (N_1217,In_287,In_1811);
nor U1218 (N_1218,In_1064,In_1467);
xnor U1219 (N_1219,In_209,In_1836);
nor U1220 (N_1220,In_1009,In_303);
nor U1221 (N_1221,In_282,In_607);
nand U1222 (N_1222,In_1550,In_791);
nor U1223 (N_1223,In_537,In_38);
or U1224 (N_1224,In_1632,In_331);
and U1225 (N_1225,In_816,In_1817);
xnor U1226 (N_1226,In_54,In_1366);
or U1227 (N_1227,In_378,In_1552);
xnor U1228 (N_1228,In_36,In_367);
or U1229 (N_1229,In_1502,In_397);
and U1230 (N_1230,In_1583,In_628);
or U1231 (N_1231,In_900,In_1627);
nand U1232 (N_1232,In_1265,In_69);
or U1233 (N_1233,In_265,In_930);
xnor U1234 (N_1234,In_1797,In_850);
nor U1235 (N_1235,In_62,In_664);
nor U1236 (N_1236,In_1557,In_379);
and U1237 (N_1237,In_18,In_578);
and U1238 (N_1238,In_1614,In_809);
nand U1239 (N_1239,In_1554,In_1884);
nand U1240 (N_1240,In_1091,In_1863);
or U1241 (N_1241,In_581,In_97);
or U1242 (N_1242,In_1797,In_162);
nor U1243 (N_1243,In_1779,In_1748);
or U1244 (N_1244,In_699,In_886);
xor U1245 (N_1245,In_1006,In_1413);
or U1246 (N_1246,In_809,In_1354);
xor U1247 (N_1247,In_1225,In_1223);
nand U1248 (N_1248,In_1740,In_1166);
xnor U1249 (N_1249,In_3,In_663);
nand U1250 (N_1250,In_131,In_1520);
and U1251 (N_1251,In_1388,In_36);
or U1252 (N_1252,In_236,In_310);
or U1253 (N_1253,In_1936,In_60);
or U1254 (N_1254,In_529,In_1149);
or U1255 (N_1255,In_1047,In_559);
and U1256 (N_1256,In_1025,In_1654);
and U1257 (N_1257,In_1686,In_130);
and U1258 (N_1258,In_793,In_1452);
or U1259 (N_1259,In_1694,In_1550);
nand U1260 (N_1260,In_70,In_838);
xnor U1261 (N_1261,In_1394,In_474);
xor U1262 (N_1262,In_303,In_180);
xor U1263 (N_1263,In_1797,In_1336);
or U1264 (N_1264,In_1240,In_1422);
xor U1265 (N_1265,In_125,In_1737);
and U1266 (N_1266,In_104,In_280);
nand U1267 (N_1267,In_1386,In_1914);
nor U1268 (N_1268,In_1393,In_1207);
nand U1269 (N_1269,In_779,In_654);
or U1270 (N_1270,In_1453,In_143);
nand U1271 (N_1271,In_799,In_31);
xor U1272 (N_1272,In_827,In_20);
and U1273 (N_1273,In_1333,In_238);
nor U1274 (N_1274,In_1054,In_792);
nand U1275 (N_1275,In_1471,In_1650);
nand U1276 (N_1276,In_1953,In_1794);
xor U1277 (N_1277,In_1989,In_670);
nand U1278 (N_1278,In_1288,In_1915);
xor U1279 (N_1279,In_390,In_1879);
nand U1280 (N_1280,In_1369,In_1414);
or U1281 (N_1281,In_1434,In_1760);
or U1282 (N_1282,In_1998,In_483);
nor U1283 (N_1283,In_1851,In_1621);
nor U1284 (N_1284,In_647,In_616);
and U1285 (N_1285,In_481,In_1708);
or U1286 (N_1286,In_1857,In_387);
nand U1287 (N_1287,In_701,In_1630);
or U1288 (N_1288,In_1372,In_936);
nor U1289 (N_1289,In_918,In_1975);
or U1290 (N_1290,In_1138,In_1855);
xnor U1291 (N_1291,In_1725,In_259);
xnor U1292 (N_1292,In_1887,In_702);
nor U1293 (N_1293,In_40,In_930);
nand U1294 (N_1294,In_884,In_1908);
and U1295 (N_1295,In_1224,In_872);
nor U1296 (N_1296,In_455,In_30);
xor U1297 (N_1297,In_647,In_223);
nand U1298 (N_1298,In_483,In_659);
and U1299 (N_1299,In_396,In_1323);
and U1300 (N_1300,In_1114,In_1253);
or U1301 (N_1301,In_1042,In_1789);
nand U1302 (N_1302,In_219,In_1432);
nand U1303 (N_1303,In_1799,In_85);
and U1304 (N_1304,In_1367,In_830);
xnor U1305 (N_1305,In_1949,In_1388);
or U1306 (N_1306,In_701,In_823);
xnor U1307 (N_1307,In_877,In_593);
xnor U1308 (N_1308,In_249,In_913);
nor U1309 (N_1309,In_260,In_712);
or U1310 (N_1310,In_1669,In_1563);
and U1311 (N_1311,In_515,In_565);
and U1312 (N_1312,In_1920,In_317);
nor U1313 (N_1313,In_822,In_832);
and U1314 (N_1314,In_620,In_453);
nand U1315 (N_1315,In_1288,In_1162);
xor U1316 (N_1316,In_1854,In_280);
or U1317 (N_1317,In_1769,In_1608);
and U1318 (N_1318,In_1531,In_1211);
nor U1319 (N_1319,In_939,In_155);
nand U1320 (N_1320,In_1739,In_1761);
nand U1321 (N_1321,In_513,In_1633);
nor U1322 (N_1322,In_492,In_1934);
or U1323 (N_1323,In_348,In_603);
nor U1324 (N_1324,In_678,In_900);
xor U1325 (N_1325,In_210,In_1205);
nor U1326 (N_1326,In_866,In_1624);
or U1327 (N_1327,In_352,In_1060);
and U1328 (N_1328,In_1608,In_279);
and U1329 (N_1329,In_979,In_180);
and U1330 (N_1330,In_925,In_358);
xnor U1331 (N_1331,In_35,In_165);
nand U1332 (N_1332,In_1173,In_1081);
xor U1333 (N_1333,In_1348,In_63);
nand U1334 (N_1334,In_1215,In_1399);
xor U1335 (N_1335,In_1605,In_300);
or U1336 (N_1336,In_651,In_1724);
nand U1337 (N_1337,In_1589,In_1485);
and U1338 (N_1338,In_346,In_212);
nand U1339 (N_1339,In_1928,In_434);
and U1340 (N_1340,In_973,In_638);
xor U1341 (N_1341,In_186,In_1622);
or U1342 (N_1342,In_54,In_475);
and U1343 (N_1343,In_1056,In_1429);
nor U1344 (N_1344,In_414,In_1801);
or U1345 (N_1345,In_575,In_762);
nand U1346 (N_1346,In_1097,In_976);
nand U1347 (N_1347,In_1325,In_1770);
xnor U1348 (N_1348,In_1068,In_131);
nor U1349 (N_1349,In_891,In_1427);
xor U1350 (N_1350,In_1091,In_355);
nand U1351 (N_1351,In_420,In_1241);
nor U1352 (N_1352,In_1131,In_1004);
and U1353 (N_1353,In_1960,In_1465);
nor U1354 (N_1354,In_1111,In_515);
nand U1355 (N_1355,In_779,In_1469);
or U1356 (N_1356,In_1528,In_1667);
or U1357 (N_1357,In_93,In_606);
nor U1358 (N_1358,In_96,In_1862);
xor U1359 (N_1359,In_330,In_1740);
and U1360 (N_1360,In_234,In_1668);
nand U1361 (N_1361,In_644,In_387);
or U1362 (N_1362,In_624,In_890);
nand U1363 (N_1363,In_523,In_1371);
nor U1364 (N_1364,In_603,In_442);
or U1365 (N_1365,In_1426,In_714);
nand U1366 (N_1366,In_1437,In_1137);
nand U1367 (N_1367,In_1991,In_1334);
nor U1368 (N_1368,In_454,In_1059);
or U1369 (N_1369,In_1819,In_814);
and U1370 (N_1370,In_622,In_1054);
nor U1371 (N_1371,In_366,In_401);
and U1372 (N_1372,In_1688,In_235);
nor U1373 (N_1373,In_661,In_1051);
and U1374 (N_1374,In_656,In_424);
or U1375 (N_1375,In_479,In_1840);
or U1376 (N_1376,In_1552,In_635);
nor U1377 (N_1377,In_773,In_1966);
xnor U1378 (N_1378,In_1968,In_941);
and U1379 (N_1379,In_537,In_41);
and U1380 (N_1380,In_1842,In_812);
nor U1381 (N_1381,In_384,In_430);
and U1382 (N_1382,In_670,In_1101);
and U1383 (N_1383,In_1590,In_767);
or U1384 (N_1384,In_1519,In_1252);
and U1385 (N_1385,In_19,In_681);
nor U1386 (N_1386,In_1170,In_739);
nor U1387 (N_1387,In_1197,In_840);
nand U1388 (N_1388,In_897,In_1558);
or U1389 (N_1389,In_1186,In_577);
or U1390 (N_1390,In_484,In_872);
xor U1391 (N_1391,In_1754,In_1919);
xnor U1392 (N_1392,In_423,In_1037);
nand U1393 (N_1393,In_1354,In_280);
nand U1394 (N_1394,In_1896,In_37);
nand U1395 (N_1395,In_496,In_1708);
xor U1396 (N_1396,In_422,In_1619);
or U1397 (N_1397,In_653,In_1858);
nand U1398 (N_1398,In_95,In_453);
or U1399 (N_1399,In_836,In_1970);
nor U1400 (N_1400,In_1747,In_1732);
nand U1401 (N_1401,In_1139,In_1541);
or U1402 (N_1402,In_1622,In_1415);
or U1403 (N_1403,In_573,In_386);
nand U1404 (N_1404,In_1901,In_1502);
nor U1405 (N_1405,In_1779,In_781);
xor U1406 (N_1406,In_1513,In_1975);
and U1407 (N_1407,In_1389,In_691);
and U1408 (N_1408,In_249,In_1528);
nor U1409 (N_1409,In_1997,In_674);
and U1410 (N_1410,In_1054,In_1509);
nand U1411 (N_1411,In_133,In_864);
or U1412 (N_1412,In_708,In_87);
nor U1413 (N_1413,In_747,In_1332);
xor U1414 (N_1414,In_1597,In_1351);
and U1415 (N_1415,In_407,In_1997);
and U1416 (N_1416,In_1998,In_137);
nand U1417 (N_1417,In_1455,In_1132);
and U1418 (N_1418,In_1930,In_227);
nand U1419 (N_1419,In_246,In_775);
xor U1420 (N_1420,In_741,In_1643);
xnor U1421 (N_1421,In_1368,In_792);
xnor U1422 (N_1422,In_1812,In_542);
and U1423 (N_1423,In_1905,In_444);
nor U1424 (N_1424,In_1287,In_120);
or U1425 (N_1425,In_417,In_1672);
nand U1426 (N_1426,In_574,In_1833);
nor U1427 (N_1427,In_399,In_1377);
nor U1428 (N_1428,In_819,In_1745);
nand U1429 (N_1429,In_665,In_1557);
nand U1430 (N_1430,In_1493,In_656);
or U1431 (N_1431,In_559,In_984);
nand U1432 (N_1432,In_700,In_1468);
or U1433 (N_1433,In_1714,In_1349);
or U1434 (N_1434,In_1218,In_1061);
xor U1435 (N_1435,In_1045,In_668);
nand U1436 (N_1436,In_255,In_403);
nor U1437 (N_1437,In_1634,In_825);
and U1438 (N_1438,In_978,In_1445);
xor U1439 (N_1439,In_880,In_1499);
nor U1440 (N_1440,In_799,In_46);
xnor U1441 (N_1441,In_1778,In_157);
and U1442 (N_1442,In_1414,In_132);
xnor U1443 (N_1443,In_82,In_1245);
xor U1444 (N_1444,In_743,In_922);
or U1445 (N_1445,In_1747,In_732);
and U1446 (N_1446,In_1692,In_491);
xor U1447 (N_1447,In_573,In_815);
xnor U1448 (N_1448,In_1357,In_1710);
or U1449 (N_1449,In_147,In_337);
and U1450 (N_1450,In_1406,In_89);
or U1451 (N_1451,In_1869,In_1228);
or U1452 (N_1452,In_1655,In_1313);
nor U1453 (N_1453,In_266,In_184);
or U1454 (N_1454,In_21,In_1037);
and U1455 (N_1455,In_134,In_1449);
nand U1456 (N_1456,In_68,In_43);
and U1457 (N_1457,In_1040,In_71);
or U1458 (N_1458,In_1822,In_1870);
and U1459 (N_1459,In_1926,In_680);
nand U1460 (N_1460,In_1574,In_1330);
xnor U1461 (N_1461,In_688,In_548);
nor U1462 (N_1462,In_1223,In_1246);
xor U1463 (N_1463,In_583,In_651);
nand U1464 (N_1464,In_1301,In_1221);
nand U1465 (N_1465,In_141,In_593);
or U1466 (N_1466,In_825,In_779);
or U1467 (N_1467,In_652,In_1497);
nand U1468 (N_1468,In_69,In_507);
xnor U1469 (N_1469,In_1536,In_656);
nor U1470 (N_1470,In_1321,In_812);
or U1471 (N_1471,In_1302,In_1553);
nor U1472 (N_1472,In_1488,In_1859);
or U1473 (N_1473,In_1596,In_991);
and U1474 (N_1474,In_1773,In_865);
nor U1475 (N_1475,In_1292,In_1668);
nand U1476 (N_1476,In_24,In_1187);
and U1477 (N_1477,In_911,In_1183);
or U1478 (N_1478,In_2,In_1642);
nand U1479 (N_1479,In_25,In_1081);
or U1480 (N_1480,In_743,In_1079);
xnor U1481 (N_1481,In_1648,In_919);
and U1482 (N_1482,In_1108,In_1725);
nand U1483 (N_1483,In_715,In_1516);
or U1484 (N_1484,In_614,In_1697);
and U1485 (N_1485,In_537,In_74);
or U1486 (N_1486,In_1767,In_188);
and U1487 (N_1487,In_1629,In_444);
and U1488 (N_1488,In_1630,In_633);
and U1489 (N_1489,In_809,In_1505);
and U1490 (N_1490,In_890,In_1735);
or U1491 (N_1491,In_49,In_1521);
or U1492 (N_1492,In_93,In_1072);
and U1493 (N_1493,In_1671,In_1064);
nor U1494 (N_1494,In_1479,In_1746);
xor U1495 (N_1495,In_760,In_705);
or U1496 (N_1496,In_1921,In_558);
nand U1497 (N_1497,In_678,In_155);
or U1498 (N_1498,In_1751,In_1772);
nand U1499 (N_1499,In_838,In_23);
xor U1500 (N_1500,In_915,In_1920);
nand U1501 (N_1501,In_954,In_1088);
or U1502 (N_1502,In_325,In_1946);
nand U1503 (N_1503,In_694,In_245);
xor U1504 (N_1504,In_320,In_810);
xnor U1505 (N_1505,In_1124,In_1767);
xor U1506 (N_1506,In_1586,In_401);
nand U1507 (N_1507,In_1604,In_1598);
nand U1508 (N_1508,In_1991,In_513);
or U1509 (N_1509,In_205,In_306);
xnor U1510 (N_1510,In_412,In_1770);
nand U1511 (N_1511,In_1983,In_788);
xnor U1512 (N_1512,In_1153,In_216);
and U1513 (N_1513,In_1838,In_1448);
or U1514 (N_1514,In_1712,In_773);
or U1515 (N_1515,In_374,In_1378);
xor U1516 (N_1516,In_460,In_213);
nand U1517 (N_1517,In_1858,In_522);
nand U1518 (N_1518,In_1838,In_1191);
and U1519 (N_1519,In_255,In_86);
or U1520 (N_1520,In_634,In_1202);
nand U1521 (N_1521,In_886,In_1900);
nor U1522 (N_1522,In_63,In_1589);
and U1523 (N_1523,In_1401,In_1960);
xnor U1524 (N_1524,In_271,In_1810);
xor U1525 (N_1525,In_763,In_1517);
nor U1526 (N_1526,In_763,In_1018);
and U1527 (N_1527,In_90,In_1060);
and U1528 (N_1528,In_692,In_1476);
xor U1529 (N_1529,In_928,In_1924);
or U1530 (N_1530,In_1619,In_1184);
nor U1531 (N_1531,In_639,In_949);
nand U1532 (N_1532,In_236,In_1317);
and U1533 (N_1533,In_1677,In_21);
nand U1534 (N_1534,In_421,In_1562);
nand U1535 (N_1535,In_18,In_591);
and U1536 (N_1536,In_1638,In_895);
and U1537 (N_1537,In_317,In_1214);
and U1538 (N_1538,In_211,In_577);
nor U1539 (N_1539,In_1478,In_1151);
nor U1540 (N_1540,In_1985,In_877);
nand U1541 (N_1541,In_654,In_523);
and U1542 (N_1542,In_175,In_635);
and U1543 (N_1543,In_1847,In_1669);
nor U1544 (N_1544,In_308,In_1783);
nor U1545 (N_1545,In_1766,In_1857);
nor U1546 (N_1546,In_1744,In_1418);
or U1547 (N_1547,In_1258,In_93);
nor U1548 (N_1548,In_1643,In_1183);
or U1549 (N_1549,In_664,In_1089);
xor U1550 (N_1550,In_1946,In_1087);
xnor U1551 (N_1551,In_1061,In_1968);
nor U1552 (N_1552,In_1740,In_589);
or U1553 (N_1553,In_1198,In_994);
nand U1554 (N_1554,In_1362,In_1184);
or U1555 (N_1555,In_1561,In_38);
xnor U1556 (N_1556,In_1829,In_779);
xor U1557 (N_1557,In_995,In_233);
and U1558 (N_1558,In_1054,In_1206);
xor U1559 (N_1559,In_1249,In_1746);
xor U1560 (N_1560,In_876,In_1851);
and U1561 (N_1561,In_639,In_1766);
nand U1562 (N_1562,In_293,In_1376);
xnor U1563 (N_1563,In_868,In_1173);
or U1564 (N_1564,In_259,In_966);
nand U1565 (N_1565,In_1556,In_1206);
xor U1566 (N_1566,In_986,In_1536);
nand U1567 (N_1567,In_858,In_176);
xnor U1568 (N_1568,In_709,In_1784);
or U1569 (N_1569,In_1387,In_662);
nand U1570 (N_1570,In_955,In_610);
and U1571 (N_1571,In_17,In_812);
or U1572 (N_1572,In_47,In_16);
xor U1573 (N_1573,In_1599,In_875);
xor U1574 (N_1574,In_836,In_622);
nand U1575 (N_1575,In_186,In_375);
or U1576 (N_1576,In_1772,In_472);
xnor U1577 (N_1577,In_1825,In_30);
xor U1578 (N_1578,In_838,In_882);
nand U1579 (N_1579,In_291,In_445);
and U1580 (N_1580,In_421,In_1829);
nor U1581 (N_1581,In_73,In_1357);
xnor U1582 (N_1582,In_1200,In_1827);
and U1583 (N_1583,In_95,In_269);
or U1584 (N_1584,In_1568,In_467);
nand U1585 (N_1585,In_330,In_736);
xor U1586 (N_1586,In_210,In_1207);
and U1587 (N_1587,In_1471,In_1230);
or U1588 (N_1588,In_870,In_1405);
or U1589 (N_1589,In_839,In_1545);
nand U1590 (N_1590,In_1164,In_22);
xor U1591 (N_1591,In_656,In_1660);
nor U1592 (N_1592,In_1124,In_1205);
nor U1593 (N_1593,In_1099,In_851);
or U1594 (N_1594,In_224,In_286);
nand U1595 (N_1595,In_597,In_846);
and U1596 (N_1596,In_905,In_220);
and U1597 (N_1597,In_1093,In_157);
and U1598 (N_1598,In_303,In_127);
nand U1599 (N_1599,In_1896,In_779);
nand U1600 (N_1600,In_1562,In_1513);
or U1601 (N_1601,In_1854,In_1979);
or U1602 (N_1602,In_1889,In_1622);
nand U1603 (N_1603,In_1568,In_1725);
and U1604 (N_1604,In_17,In_1064);
nand U1605 (N_1605,In_415,In_210);
or U1606 (N_1606,In_284,In_1044);
xnor U1607 (N_1607,In_775,In_1003);
nor U1608 (N_1608,In_887,In_95);
or U1609 (N_1609,In_575,In_1010);
xnor U1610 (N_1610,In_1045,In_1056);
or U1611 (N_1611,In_1567,In_255);
nor U1612 (N_1612,In_204,In_1107);
and U1613 (N_1613,In_1796,In_849);
nor U1614 (N_1614,In_1493,In_158);
nand U1615 (N_1615,In_444,In_450);
nor U1616 (N_1616,In_889,In_953);
xor U1617 (N_1617,In_1832,In_959);
or U1618 (N_1618,In_1342,In_740);
or U1619 (N_1619,In_502,In_546);
and U1620 (N_1620,In_697,In_568);
or U1621 (N_1621,In_1665,In_1029);
nor U1622 (N_1622,In_1910,In_1625);
xor U1623 (N_1623,In_1867,In_195);
or U1624 (N_1624,In_1015,In_1354);
nand U1625 (N_1625,In_981,In_1659);
or U1626 (N_1626,In_1813,In_1772);
nand U1627 (N_1627,In_1032,In_1607);
xnor U1628 (N_1628,In_0,In_398);
and U1629 (N_1629,In_781,In_1919);
nand U1630 (N_1630,In_1066,In_810);
and U1631 (N_1631,In_1016,In_619);
nand U1632 (N_1632,In_1955,In_1012);
nand U1633 (N_1633,In_1059,In_1796);
or U1634 (N_1634,In_1655,In_1682);
nand U1635 (N_1635,In_648,In_1935);
nand U1636 (N_1636,In_613,In_996);
or U1637 (N_1637,In_1763,In_208);
or U1638 (N_1638,In_1341,In_1060);
nor U1639 (N_1639,In_1766,In_1399);
and U1640 (N_1640,In_466,In_1783);
or U1641 (N_1641,In_1963,In_929);
xnor U1642 (N_1642,In_44,In_524);
xnor U1643 (N_1643,In_517,In_1436);
nor U1644 (N_1644,In_907,In_81);
and U1645 (N_1645,In_491,In_371);
or U1646 (N_1646,In_1041,In_83);
nor U1647 (N_1647,In_145,In_519);
and U1648 (N_1648,In_181,In_1315);
and U1649 (N_1649,In_608,In_620);
and U1650 (N_1650,In_509,In_26);
nand U1651 (N_1651,In_192,In_1410);
or U1652 (N_1652,In_1434,In_1438);
and U1653 (N_1653,In_1192,In_733);
and U1654 (N_1654,In_1569,In_226);
nand U1655 (N_1655,In_100,In_800);
and U1656 (N_1656,In_715,In_892);
xor U1657 (N_1657,In_800,In_1084);
xor U1658 (N_1658,In_469,In_1087);
nand U1659 (N_1659,In_1882,In_944);
nand U1660 (N_1660,In_125,In_1006);
xor U1661 (N_1661,In_148,In_1182);
nor U1662 (N_1662,In_1253,In_352);
nand U1663 (N_1663,In_1555,In_1163);
xor U1664 (N_1664,In_1204,In_777);
nor U1665 (N_1665,In_359,In_1291);
xnor U1666 (N_1666,In_485,In_1921);
xor U1667 (N_1667,In_1932,In_1922);
or U1668 (N_1668,In_1629,In_92);
or U1669 (N_1669,In_311,In_1672);
nand U1670 (N_1670,In_1662,In_1734);
xor U1671 (N_1671,In_53,In_263);
nand U1672 (N_1672,In_1326,In_1541);
or U1673 (N_1673,In_1339,In_1100);
nand U1674 (N_1674,In_1051,In_1455);
or U1675 (N_1675,In_0,In_1855);
nor U1676 (N_1676,In_1110,In_1774);
nand U1677 (N_1677,In_1821,In_1137);
or U1678 (N_1678,In_1040,In_939);
and U1679 (N_1679,In_1728,In_1838);
nand U1680 (N_1680,In_346,In_517);
nor U1681 (N_1681,In_12,In_1311);
nand U1682 (N_1682,In_1875,In_471);
or U1683 (N_1683,In_1735,In_1859);
xor U1684 (N_1684,In_311,In_1357);
and U1685 (N_1685,In_1390,In_923);
nand U1686 (N_1686,In_1624,In_1933);
xnor U1687 (N_1687,In_1792,In_1);
or U1688 (N_1688,In_1905,In_633);
and U1689 (N_1689,In_1702,In_162);
nand U1690 (N_1690,In_994,In_684);
nand U1691 (N_1691,In_985,In_161);
nor U1692 (N_1692,In_1930,In_1240);
or U1693 (N_1693,In_493,In_1387);
nand U1694 (N_1694,In_576,In_1847);
nor U1695 (N_1695,In_1317,In_1326);
and U1696 (N_1696,In_892,In_1253);
or U1697 (N_1697,In_1015,In_1765);
nand U1698 (N_1698,In_590,In_1282);
xnor U1699 (N_1699,In_951,In_1166);
nand U1700 (N_1700,In_521,In_1268);
or U1701 (N_1701,In_1598,In_378);
or U1702 (N_1702,In_1203,In_1046);
nor U1703 (N_1703,In_220,In_142);
xor U1704 (N_1704,In_1665,In_590);
and U1705 (N_1705,In_1092,In_538);
or U1706 (N_1706,In_1063,In_373);
nor U1707 (N_1707,In_360,In_1783);
nor U1708 (N_1708,In_771,In_539);
and U1709 (N_1709,In_371,In_1602);
xor U1710 (N_1710,In_851,In_1562);
and U1711 (N_1711,In_177,In_285);
nand U1712 (N_1712,In_1912,In_808);
and U1713 (N_1713,In_752,In_1343);
or U1714 (N_1714,In_22,In_672);
xnor U1715 (N_1715,In_753,In_1642);
or U1716 (N_1716,In_1256,In_294);
or U1717 (N_1717,In_799,In_1799);
and U1718 (N_1718,In_977,In_735);
nand U1719 (N_1719,In_23,In_1324);
and U1720 (N_1720,In_512,In_1289);
xnor U1721 (N_1721,In_1764,In_1834);
nor U1722 (N_1722,In_272,In_1428);
and U1723 (N_1723,In_1374,In_1901);
xor U1724 (N_1724,In_886,In_91);
nor U1725 (N_1725,In_1580,In_411);
nor U1726 (N_1726,In_1210,In_1987);
xnor U1727 (N_1727,In_25,In_377);
nor U1728 (N_1728,In_1340,In_1121);
xor U1729 (N_1729,In_250,In_1045);
and U1730 (N_1730,In_465,In_670);
nand U1731 (N_1731,In_136,In_719);
nand U1732 (N_1732,In_179,In_176);
nand U1733 (N_1733,In_1124,In_1309);
and U1734 (N_1734,In_481,In_265);
or U1735 (N_1735,In_265,In_1587);
nand U1736 (N_1736,In_486,In_1938);
nor U1737 (N_1737,In_84,In_227);
nor U1738 (N_1738,In_908,In_1280);
nand U1739 (N_1739,In_1745,In_331);
or U1740 (N_1740,In_1620,In_1679);
nand U1741 (N_1741,In_953,In_1641);
xnor U1742 (N_1742,In_1928,In_1687);
and U1743 (N_1743,In_1403,In_497);
or U1744 (N_1744,In_414,In_1269);
nor U1745 (N_1745,In_1485,In_1091);
nand U1746 (N_1746,In_1157,In_1759);
and U1747 (N_1747,In_638,In_643);
and U1748 (N_1748,In_1389,In_1922);
nand U1749 (N_1749,In_1764,In_26);
or U1750 (N_1750,In_1124,In_360);
nand U1751 (N_1751,In_411,In_1581);
or U1752 (N_1752,In_1257,In_506);
nor U1753 (N_1753,In_1578,In_671);
or U1754 (N_1754,In_1118,In_1133);
nand U1755 (N_1755,In_1852,In_1550);
and U1756 (N_1756,In_53,In_1180);
and U1757 (N_1757,In_383,In_370);
and U1758 (N_1758,In_625,In_1315);
nand U1759 (N_1759,In_1883,In_1721);
xor U1760 (N_1760,In_1045,In_620);
and U1761 (N_1761,In_342,In_1599);
and U1762 (N_1762,In_1453,In_1293);
xor U1763 (N_1763,In_1149,In_1139);
or U1764 (N_1764,In_1752,In_1621);
and U1765 (N_1765,In_739,In_553);
xnor U1766 (N_1766,In_594,In_1488);
nor U1767 (N_1767,In_1281,In_1745);
nor U1768 (N_1768,In_1262,In_1242);
and U1769 (N_1769,In_670,In_1148);
and U1770 (N_1770,In_547,In_1033);
nand U1771 (N_1771,In_1344,In_1393);
nand U1772 (N_1772,In_829,In_1000);
xnor U1773 (N_1773,In_637,In_129);
nor U1774 (N_1774,In_1266,In_49);
nand U1775 (N_1775,In_869,In_788);
and U1776 (N_1776,In_1956,In_137);
xor U1777 (N_1777,In_493,In_781);
and U1778 (N_1778,In_521,In_483);
nand U1779 (N_1779,In_1166,In_116);
or U1780 (N_1780,In_1724,In_579);
nor U1781 (N_1781,In_1191,In_889);
nand U1782 (N_1782,In_284,In_1590);
nor U1783 (N_1783,In_1574,In_647);
or U1784 (N_1784,In_1038,In_1550);
and U1785 (N_1785,In_1474,In_941);
and U1786 (N_1786,In_298,In_335);
xnor U1787 (N_1787,In_40,In_1000);
or U1788 (N_1788,In_1345,In_793);
nor U1789 (N_1789,In_960,In_1931);
nand U1790 (N_1790,In_717,In_1236);
or U1791 (N_1791,In_371,In_271);
and U1792 (N_1792,In_1457,In_237);
or U1793 (N_1793,In_34,In_1092);
and U1794 (N_1794,In_1035,In_1071);
nor U1795 (N_1795,In_823,In_926);
nand U1796 (N_1796,In_1464,In_666);
or U1797 (N_1797,In_737,In_1880);
or U1798 (N_1798,In_1988,In_1340);
and U1799 (N_1799,In_534,In_956);
xnor U1800 (N_1800,In_1705,In_1029);
nor U1801 (N_1801,In_216,In_1776);
nand U1802 (N_1802,In_1738,In_585);
nor U1803 (N_1803,In_1421,In_1371);
nand U1804 (N_1804,In_1920,In_1150);
nor U1805 (N_1805,In_1226,In_51);
xnor U1806 (N_1806,In_1032,In_582);
and U1807 (N_1807,In_646,In_1926);
nor U1808 (N_1808,In_887,In_529);
nand U1809 (N_1809,In_26,In_1007);
or U1810 (N_1810,In_1696,In_294);
or U1811 (N_1811,In_235,In_1973);
or U1812 (N_1812,In_466,In_1349);
or U1813 (N_1813,In_1450,In_1531);
nand U1814 (N_1814,In_1984,In_116);
and U1815 (N_1815,In_754,In_1119);
nor U1816 (N_1816,In_774,In_1679);
and U1817 (N_1817,In_83,In_870);
and U1818 (N_1818,In_1605,In_1780);
and U1819 (N_1819,In_1780,In_1869);
and U1820 (N_1820,In_1923,In_974);
nor U1821 (N_1821,In_43,In_1061);
nor U1822 (N_1822,In_1461,In_94);
and U1823 (N_1823,In_1944,In_178);
nor U1824 (N_1824,In_1808,In_969);
nor U1825 (N_1825,In_1487,In_1624);
or U1826 (N_1826,In_1721,In_1321);
and U1827 (N_1827,In_299,In_698);
nor U1828 (N_1828,In_511,In_663);
nor U1829 (N_1829,In_1152,In_1835);
or U1830 (N_1830,In_1738,In_571);
or U1831 (N_1831,In_1152,In_963);
or U1832 (N_1832,In_1815,In_142);
nand U1833 (N_1833,In_405,In_1631);
and U1834 (N_1834,In_1600,In_1175);
xnor U1835 (N_1835,In_1533,In_579);
nor U1836 (N_1836,In_1508,In_304);
nor U1837 (N_1837,In_1392,In_934);
and U1838 (N_1838,In_1696,In_1998);
nand U1839 (N_1839,In_364,In_134);
nor U1840 (N_1840,In_243,In_1645);
nor U1841 (N_1841,In_129,In_731);
or U1842 (N_1842,In_1987,In_1059);
xnor U1843 (N_1843,In_223,In_1804);
or U1844 (N_1844,In_1871,In_1990);
nand U1845 (N_1845,In_1770,In_1093);
nor U1846 (N_1846,In_544,In_1939);
nand U1847 (N_1847,In_1734,In_1394);
xnor U1848 (N_1848,In_186,In_837);
or U1849 (N_1849,In_1648,In_1164);
xnor U1850 (N_1850,In_503,In_878);
or U1851 (N_1851,In_992,In_994);
xor U1852 (N_1852,In_920,In_1502);
or U1853 (N_1853,In_572,In_1665);
nor U1854 (N_1854,In_315,In_84);
and U1855 (N_1855,In_105,In_712);
and U1856 (N_1856,In_176,In_456);
nor U1857 (N_1857,In_985,In_1494);
nor U1858 (N_1858,In_480,In_819);
nand U1859 (N_1859,In_206,In_798);
nor U1860 (N_1860,In_72,In_601);
and U1861 (N_1861,In_42,In_829);
nand U1862 (N_1862,In_1138,In_434);
or U1863 (N_1863,In_950,In_1050);
or U1864 (N_1864,In_722,In_716);
nor U1865 (N_1865,In_1996,In_1959);
nor U1866 (N_1866,In_764,In_1459);
nor U1867 (N_1867,In_1283,In_1574);
xor U1868 (N_1868,In_1366,In_860);
nand U1869 (N_1869,In_1505,In_1185);
xor U1870 (N_1870,In_796,In_1221);
nand U1871 (N_1871,In_1328,In_654);
xnor U1872 (N_1872,In_377,In_7);
or U1873 (N_1873,In_275,In_1307);
or U1874 (N_1874,In_409,In_1357);
and U1875 (N_1875,In_1424,In_1766);
nor U1876 (N_1876,In_828,In_1311);
or U1877 (N_1877,In_1119,In_1771);
or U1878 (N_1878,In_231,In_1028);
nor U1879 (N_1879,In_640,In_1101);
xnor U1880 (N_1880,In_1870,In_151);
nor U1881 (N_1881,In_358,In_394);
nand U1882 (N_1882,In_1193,In_558);
nand U1883 (N_1883,In_774,In_1139);
and U1884 (N_1884,In_596,In_1987);
nand U1885 (N_1885,In_1812,In_1117);
or U1886 (N_1886,In_624,In_155);
xor U1887 (N_1887,In_1625,In_1054);
or U1888 (N_1888,In_598,In_1412);
xor U1889 (N_1889,In_705,In_1269);
and U1890 (N_1890,In_1492,In_1335);
nand U1891 (N_1891,In_689,In_1019);
nor U1892 (N_1892,In_40,In_224);
or U1893 (N_1893,In_1567,In_1825);
nor U1894 (N_1894,In_857,In_1094);
nor U1895 (N_1895,In_626,In_1820);
or U1896 (N_1896,In_965,In_1004);
and U1897 (N_1897,In_277,In_1434);
nand U1898 (N_1898,In_634,In_471);
and U1899 (N_1899,In_337,In_91);
xnor U1900 (N_1900,In_93,In_315);
and U1901 (N_1901,In_1211,In_102);
nor U1902 (N_1902,In_868,In_679);
xor U1903 (N_1903,In_430,In_600);
and U1904 (N_1904,In_479,In_1120);
nor U1905 (N_1905,In_378,In_1983);
or U1906 (N_1906,In_580,In_259);
nor U1907 (N_1907,In_88,In_1566);
nor U1908 (N_1908,In_1881,In_807);
and U1909 (N_1909,In_1500,In_676);
nand U1910 (N_1910,In_734,In_1598);
nor U1911 (N_1911,In_1881,In_468);
or U1912 (N_1912,In_1239,In_780);
or U1913 (N_1913,In_1971,In_1341);
nor U1914 (N_1914,In_1533,In_1431);
and U1915 (N_1915,In_604,In_1048);
or U1916 (N_1916,In_1413,In_1469);
xnor U1917 (N_1917,In_590,In_81);
or U1918 (N_1918,In_1022,In_817);
and U1919 (N_1919,In_1609,In_1760);
and U1920 (N_1920,In_1075,In_766);
nand U1921 (N_1921,In_355,In_347);
or U1922 (N_1922,In_54,In_1500);
and U1923 (N_1923,In_1693,In_1969);
nand U1924 (N_1924,In_290,In_382);
nor U1925 (N_1925,In_1979,In_1414);
or U1926 (N_1926,In_1677,In_1013);
nor U1927 (N_1927,In_1523,In_1199);
and U1928 (N_1928,In_1570,In_88);
or U1929 (N_1929,In_1404,In_281);
or U1930 (N_1930,In_1015,In_235);
and U1931 (N_1931,In_1154,In_823);
nand U1932 (N_1932,In_1914,In_1014);
or U1933 (N_1933,In_798,In_682);
and U1934 (N_1934,In_1864,In_970);
nor U1935 (N_1935,In_381,In_1466);
nand U1936 (N_1936,In_1690,In_390);
xor U1937 (N_1937,In_1191,In_505);
xnor U1938 (N_1938,In_1571,In_1533);
xnor U1939 (N_1939,In_286,In_20);
nand U1940 (N_1940,In_1612,In_1547);
nor U1941 (N_1941,In_552,In_1472);
nand U1942 (N_1942,In_1250,In_1496);
xor U1943 (N_1943,In_1226,In_670);
xor U1944 (N_1944,In_1954,In_96);
nor U1945 (N_1945,In_1843,In_444);
nand U1946 (N_1946,In_1591,In_411);
xnor U1947 (N_1947,In_1992,In_1787);
nor U1948 (N_1948,In_1495,In_896);
or U1949 (N_1949,In_1175,In_387);
xor U1950 (N_1950,In_990,In_1141);
or U1951 (N_1951,In_1567,In_1873);
nand U1952 (N_1952,In_1747,In_364);
nand U1953 (N_1953,In_778,In_786);
and U1954 (N_1954,In_732,In_1920);
and U1955 (N_1955,In_1095,In_99);
or U1956 (N_1956,In_1391,In_41);
nor U1957 (N_1957,In_100,In_1644);
xor U1958 (N_1958,In_1548,In_895);
nor U1959 (N_1959,In_46,In_823);
nand U1960 (N_1960,In_1411,In_1321);
nand U1961 (N_1961,In_1143,In_656);
and U1962 (N_1962,In_255,In_1235);
and U1963 (N_1963,In_871,In_601);
or U1964 (N_1964,In_766,In_1090);
and U1965 (N_1965,In_438,In_1197);
nand U1966 (N_1966,In_118,In_654);
or U1967 (N_1967,In_779,In_1183);
or U1968 (N_1968,In_422,In_1726);
or U1969 (N_1969,In_1126,In_1522);
or U1970 (N_1970,In_917,In_635);
and U1971 (N_1971,In_610,In_1256);
xor U1972 (N_1972,In_333,In_646);
xor U1973 (N_1973,In_1612,In_1849);
nor U1974 (N_1974,In_151,In_1569);
xor U1975 (N_1975,In_52,In_1953);
and U1976 (N_1976,In_458,In_1349);
nor U1977 (N_1977,In_1061,In_1106);
or U1978 (N_1978,In_813,In_1709);
or U1979 (N_1979,In_1725,In_711);
or U1980 (N_1980,In_677,In_124);
and U1981 (N_1981,In_1570,In_1178);
nor U1982 (N_1982,In_23,In_43);
nand U1983 (N_1983,In_1310,In_525);
xnor U1984 (N_1984,In_1206,In_317);
or U1985 (N_1985,In_534,In_931);
nor U1986 (N_1986,In_1160,In_843);
xor U1987 (N_1987,In_1752,In_618);
and U1988 (N_1988,In_619,In_669);
xnor U1989 (N_1989,In_304,In_1561);
xor U1990 (N_1990,In_1228,In_396);
nand U1991 (N_1991,In_395,In_1748);
nand U1992 (N_1992,In_1753,In_1825);
nand U1993 (N_1993,In_814,In_1723);
nand U1994 (N_1994,In_136,In_1902);
xnor U1995 (N_1995,In_612,In_1630);
xor U1996 (N_1996,In_769,In_1192);
and U1997 (N_1997,In_483,In_279);
or U1998 (N_1998,In_1193,In_1522);
and U1999 (N_1999,In_753,In_1360);
and U2000 (N_2000,N_1187,N_1850);
and U2001 (N_2001,N_1009,N_1615);
or U2002 (N_2002,N_1713,N_1621);
nor U2003 (N_2003,N_236,N_1231);
and U2004 (N_2004,N_867,N_1354);
nor U2005 (N_2005,N_857,N_1948);
or U2006 (N_2006,N_541,N_1788);
and U2007 (N_2007,N_227,N_815);
and U2008 (N_2008,N_61,N_1498);
nand U2009 (N_2009,N_506,N_1366);
or U2010 (N_2010,N_1232,N_1329);
nor U2011 (N_2011,N_465,N_379);
and U2012 (N_2012,N_285,N_1571);
xnor U2013 (N_2013,N_10,N_1090);
or U2014 (N_2014,N_563,N_284);
or U2015 (N_2015,N_1899,N_1891);
and U2016 (N_2016,N_1198,N_1676);
and U2017 (N_2017,N_73,N_380);
or U2018 (N_2018,N_249,N_397);
nor U2019 (N_2019,N_1826,N_1039);
and U2020 (N_2020,N_1443,N_1549);
nand U2021 (N_2021,N_771,N_1776);
or U2022 (N_2022,N_915,N_840);
or U2023 (N_2023,N_1757,N_346);
nand U2024 (N_2024,N_1800,N_558);
and U2025 (N_2025,N_418,N_750);
nor U2026 (N_2026,N_338,N_896);
xor U2027 (N_2027,N_1897,N_138);
nand U2028 (N_2028,N_1646,N_315);
nor U2029 (N_2029,N_643,N_481);
xnor U2030 (N_2030,N_163,N_942);
or U2031 (N_2031,N_1092,N_1803);
nor U2032 (N_2032,N_1482,N_855);
and U2033 (N_2033,N_1520,N_1712);
or U2034 (N_2034,N_58,N_260);
and U2035 (N_2035,N_677,N_1315);
nand U2036 (N_2036,N_439,N_1977);
and U2037 (N_2037,N_407,N_116);
nor U2038 (N_2038,N_652,N_193);
nand U2039 (N_2039,N_1043,N_169);
nand U2040 (N_2040,N_924,N_542);
nor U2041 (N_2041,N_1679,N_1873);
and U2042 (N_2042,N_442,N_1408);
and U2043 (N_2043,N_882,N_641);
and U2044 (N_2044,N_1106,N_185);
xor U2045 (N_2045,N_1032,N_1410);
or U2046 (N_2046,N_160,N_588);
xor U2047 (N_2047,N_74,N_1244);
xnor U2048 (N_2048,N_436,N_330);
or U2049 (N_2049,N_533,N_1230);
nand U2050 (N_2050,N_953,N_837);
nor U2051 (N_2051,N_630,N_1490);
nor U2052 (N_2052,N_1184,N_134);
or U2053 (N_2053,N_1389,N_1840);
nand U2054 (N_2054,N_1377,N_871);
xor U2055 (N_2055,N_309,N_1169);
nor U2056 (N_2056,N_804,N_715);
nor U2057 (N_2057,N_1626,N_299);
xor U2058 (N_2058,N_1367,N_589);
nand U2059 (N_2059,N_1538,N_318);
and U2060 (N_2060,N_578,N_665);
nand U2061 (N_2061,N_1743,N_1220);
or U2062 (N_2062,N_1218,N_1682);
xor U2063 (N_2063,N_467,N_1732);
xor U2064 (N_2064,N_901,N_1185);
xnor U2065 (N_2065,N_1052,N_961);
nand U2066 (N_2066,N_1215,N_62);
nor U2067 (N_2067,N_707,N_1640);
and U2068 (N_2068,N_1174,N_660);
xor U2069 (N_2069,N_14,N_1099);
nor U2070 (N_2070,N_54,N_1990);
xnor U2071 (N_2071,N_673,N_1160);
xor U2072 (N_2072,N_635,N_1501);
nor U2073 (N_2073,N_229,N_1412);
nand U2074 (N_2074,N_415,N_388);
xnor U2075 (N_2075,N_1647,N_1924);
or U2076 (N_2076,N_1003,N_248);
or U2077 (N_2077,N_1260,N_605);
or U2078 (N_2078,N_949,N_1249);
nand U2079 (N_2079,N_852,N_1431);
nor U2080 (N_2080,N_1228,N_409);
nand U2081 (N_2081,N_1175,N_441);
nor U2082 (N_2082,N_1363,N_564);
and U2083 (N_2083,N_50,N_1736);
xor U2084 (N_2084,N_25,N_1478);
and U2085 (N_2085,N_631,N_1468);
nor U2086 (N_2086,N_1818,N_1305);
xnor U2087 (N_2087,N_1606,N_1950);
nand U2088 (N_2088,N_0,N_477);
nand U2089 (N_2089,N_1652,N_1123);
and U2090 (N_2090,N_1857,N_458);
xnor U2091 (N_2091,N_344,N_1296);
nor U2092 (N_2092,N_489,N_1060);
nand U2093 (N_2093,N_1759,N_352);
and U2094 (N_2094,N_734,N_28);
xnor U2095 (N_2095,N_684,N_1845);
xnor U2096 (N_2096,N_623,N_1282);
nand U2097 (N_2097,N_860,N_1864);
or U2098 (N_2098,N_1082,N_1325);
xnor U2099 (N_2099,N_1378,N_405);
nand U2100 (N_2100,N_56,N_1648);
xor U2101 (N_2101,N_547,N_688);
nor U2102 (N_2102,N_827,N_657);
or U2103 (N_2103,N_744,N_256);
nand U2104 (N_2104,N_1373,N_341);
and U2105 (N_2105,N_1726,N_647);
nand U2106 (N_2106,N_457,N_1956);
xor U2107 (N_2107,N_1669,N_199);
nor U2108 (N_2108,N_1855,N_1080);
and U2109 (N_2109,N_1239,N_1789);
nand U2110 (N_2110,N_1464,N_392);
or U2111 (N_2111,N_76,N_1341);
nand U2112 (N_2112,N_1774,N_246);
nand U2113 (N_2113,N_1405,N_1460);
nand U2114 (N_2114,N_1319,N_1739);
nand U2115 (N_2115,N_461,N_327);
nand U2116 (N_2116,N_1702,N_775);
nor U2117 (N_2117,N_1276,N_196);
nor U2118 (N_2118,N_1399,N_1946);
nand U2119 (N_2119,N_534,N_1890);
and U2120 (N_2120,N_1382,N_191);
and U2121 (N_2121,N_764,N_713);
nand U2122 (N_2122,N_30,N_1452);
xor U2123 (N_2123,N_1432,N_719);
nand U2124 (N_2124,N_1847,N_1439);
nor U2125 (N_2125,N_650,N_767);
nand U2126 (N_2126,N_1863,N_1653);
or U2127 (N_2127,N_222,N_1799);
xor U2128 (N_2128,N_640,N_1544);
and U2129 (N_2129,N_851,N_894);
and U2130 (N_2130,N_819,N_440);
xor U2131 (N_2131,N_44,N_1714);
and U2132 (N_2132,N_1256,N_1865);
nand U2133 (N_2133,N_1791,N_85);
nand U2134 (N_2134,N_1983,N_1271);
or U2135 (N_2135,N_128,N_1756);
or U2136 (N_2136,N_847,N_1278);
xor U2137 (N_2137,N_1938,N_991);
or U2138 (N_2138,N_381,N_216);
xnor U2139 (N_2139,N_472,N_1094);
nand U2140 (N_2140,N_41,N_1144);
and U2141 (N_2141,N_1006,N_416);
nor U2142 (N_2142,N_1115,N_1164);
nor U2143 (N_2143,N_549,N_1116);
and U2144 (N_2144,N_1595,N_1131);
xnor U2145 (N_2145,N_414,N_703);
nor U2146 (N_2146,N_520,N_270);
and U2147 (N_2147,N_1985,N_1825);
nand U2148 (N_2148,N_709,N_865);
and U2149 (N_2149,N_1364,N_878);
and U2150 (N_2150,N_297,N_1807);
nor U2151 (N_2151,N_1196,N_1212);
and U2152 (N_2152,N_447,N_220);
and U2153 (N_2153,N_1134,N_879);
or U2154 (N_2154,N_1969,N_658);
xnor U2155 (N_2155,N_1497,N_125);
or U2156 (N_2156,N_1604,N_1804);
xnor U2157 (N_2157,N_1635,N_551);
or U2158 (N_2158,N_259,N_853);
xor U2159 (N_2159,N_625,N_1479);
xor U2160 (N_2160,N_1475,N_36);
or U2161 (N_2161,N_1331,N_292);
or U2162 (N_2162,N_322,N_9);
xor U2163 (N_2163,N_121,N_1266);
xor U2164 (N_2164,N_1416,N_1775);
xnor U2165 (N_2165,N_947,N_8);
or U2166 (N_2166,N_258,N_96);
nor U2167 (N_2167,N_763,N_1058);
nor U2168 (N_2168,N_480,N_1254);
and U2169 (N_2169,N_1406,N_821);
nand U2170 (N_2170,N_733,N_1356);
xnor U2171 (N_2171,N_722,N_1274);
nor U2172 (N_2172,N_842,N_724);
nor U2173 (N_2173,N_1573,N_790);
and U2174 (N_2174,N_1022,N_1124);
nand U2175 (N_2175,N_1014,N_780);
nand U2176 (N_2176,N_88,N_752);
xnor U2177 (N_2177,N_264,N_65);
xor U2178 (N_2178,N_1978,N_221);
nor U2179 (N_2179,N_1411,N_336);
and U2180 (N_2180,N_1369,N_1081);
xor U2181 (N_2181,N_1062,N_1332);
or U2182 (N_2182,N_527,N_1659);
xnor U2183 (N_2183,N_437,N_130);
and U2184 (N_2184,N_1071,N_1495);
and U2185 (N_2185,N_612,N_1545);
xor U2186 (N_2186,N_404,N_376);
xnor U2187 (N_2187,N_693,N_1654);
xor U2188 (N_2188,N_124,N_1001);
nand U2189 (N_2189,N_602,N_1381);
xor U2190 (N_2190,N_166,N_353);
nand U2191 (N_2191,N_793,N_47);
nor U2192 (N_2192,N_769,N_1380);
xnor U2193 (N_2193,N_1010,N_1002);
xnor U2194 (N_2194,N_1979,N_1936);
nor U2195 (N_2195,N_1597,N_1217);
nor U2196 (N_2196,N_664,N_883);
nor U2197 (N_2197,N_1214,N_1425);
nand U2198 (N_2198,N_964,N_1592);
xor U2199 (N_2199,N_818,N_462);
or U2200 (N_2200,N_178,N_742);
and U2201 (N_2201,N_71,N_1324);
xnor U2202 (N_2202,N_1744,N_1967);
and U2203 (N_2203,N_508,N_267);
nor U2204 (N_2204,N_1657,N_543);
xor U2205 (N_2205,N_1289,N_1666);
or U2206 (N_2206,N_539,N_137);
xnor U2207 (N_2207,N_718,N_500);
and U2208 (N_2208,N_1110,N_1995);
nor U2209 (N_2209,N_1913,N_354);
xnor U2210 (N_2210,N_1072,N_203);
and U2211 (N_2211,N_1844,N_1686);
nor U2212 (N_2212,N_966,N_566);
nor U2213 (N_2213,N_432,N_908);
nand U2214 (N_2214,N_1579,N_591);
and U2215 (N_2215,N_784,N_369);
nand U2216 (N_2216,N_60,N_811);
nand U2217 (N_2217,N_778,N_911);
xor U2218 (N_2218,N_357,N_1236);
and U2219 (N_2219,N_1334,N_366);
and U2220 (N_2220,N_1581,N_826);
nand U2221 (N_2221,N_317,N_180);
or U2222 (N_2222,N_287,N_1910);
or U2223 (N_2223,N_1834,N_573);
and U2224 (N_2224,N_600,N_651);
nor U2225 (N_2225,N_708,N_799);
and U2226 (N_2226,N_1601,N_1546);
or U2227 (N_2227,N_1753,N_204);
and U2228 (N_2228,N_1028,N_721);
xnor U2229 (N_2229,N_1031,N_532);
and U2230 (N_2230,N_546,N_1991);
or U2231 (N_2231,N_998,N_1740);
or U2232 (N_2232,N_1209,N_3);
xor U2233 (N_2233,N_300,N_536);
or U2234 (N_2234,N_306,N_1513);
nor U2235 (N_2235,N_1610,N_1359);
nor U2236 (N_2236,N_1121,N_999);
or U2237 (N_2237,N_1414,N_922);
xor U2238 (N_2238,N_1782,N_38);
or U2239 (N_2239,N_522,N_1917);
xor U2240 (N_2240,N_1245,N_240);
or U2241 (N_2241,N_1643,N_1565);
or U2242 (N_2242,N_152,N_401);
nand U2243 (N_2243,N_599,N_776);
and U2244 (N_2244,N_893,N_1450);
nand U2245 (N_2245,N_1088,N_21);
nand U2246 (N_2246,N_704,N_412);
and U2247 (N_2247,N_1469,N_1277);
nand U2248 (N_2248,N_754,N_282);
and U2249 (N_2249,N_213,N_269);
nand U2250 (N_2250,N_1057,N_385);
or U2251 (N_2251,N_1663,N_1104);
and U2252 (N_2252,N_490,N_1383);
nand U2253 (N_2253,N_413,N_1190);
or U2254 (N_2254,N_1293,N_1777);
nor U2255 (N_2255,N_325,N_615);
and U2256 (N_2256,N_1178,N_601);
nand U2257 (N_2257,N_1859,N_459);
nor U2258 (N_2258,N_1824,N_792);
xnor U2259 (N_2259,N_604,N_1179);
and U2260 (N_2260,N_1896,N_503);
nand U2261 (N_2261,N_1612,N_1519);
and U2262 (N_2262,N_1150,N_984);
nor U2263 (N_2263,N_759,N_123);
xnor U2264 (N_2264,N_177,N_181);
nand U2265 (N_2265,N_271,N_934);
xor U2266 (N_2266,N_1133,N_1201);
nand U2267 (N_2267,N_1441,N_788);
nand U2268 (N_2268,N_1370,N_861);
nor U2269 (N_2269,N_841,N_510);
nor U2270 (N_2270,N_1697,N_1958);
or U2271 (N_2271,N_1151,N_1858);
nor U2272 (N_2272,N_712,N_476);
and U2273 (N_2273,N_1837,N_1079);
nand U2274 (N_2274,N_1024,N_1182);
nor U2275 (N_2275,N_424,N_1591);
xor U2276 (N_2276,N_498,N_1796);
nand U2277 (N_2277,N_1255,N_1516);
or U2278 (N_2278,N_349,N_1842);
nor U2279 (N_2279,N_1993,N_176);
nor U2280 (N_2280,N_823,N_323);
or U2281 (N_2281,N_1314,N_807);
xor U2282 (N_2282,N_1534,N_175);
or U2283 (N_2283,N_512,N_740);
or U2284 (N_2284,N_1132,N_1952);
xor U2285 (N_2285,N_830,N_1030);
or U2286 (N_2286,N_530,N_581);
nor U2287 (N_2287,N_1698,N_399);
nor U2288 (N_2288,N_988,N_279);
xor U2289 (N_2289,N_79,N_1149);
xor U2290 (N_2290,N_1407,N_1881);
nand U2291 (N_2291,N_24,N_1103);
or U2292 (N_2292,N_1651,N_1265);
and U2293 (N_2293,N_691,N_1922);
and U2294 (N_2294,N_828,N_1846);
xor U2295 (N_2295,N_219,N_314);
and U2296 (N_2296,N_1729,N_945);
or U2297 (N_2297,N_1795,N_1784);
nand U2298 (N_2298,N_1045,N_245);
and U2299 (N_2299,N_812,N_1869);
nor U2300 (N_2300,N_1529,N_1507);
or U2301 (N_2301,N_449,N_854);
and U2302 (N_2302,N_1980,N_1394);
nand U2303 (N_2303,N_629,N_1456);
or U2304 (N_2304,N_1303,N_1861);
and U2305 (N_2305,N_1954,N_1633);
xnor U2306 (N_2306,N_210,N_1477);
or U2307 (N_2307,N_482,N_1848);
nand U2308 (N_2308,N_694,N_406);
and U2309 (N_2309,N_1570,N_1792);
nor U2310 (N_2310,N_11,N_585);
or U2311 (N_2311,N_1975,N_1596);
nand U2312 (N_2312,N_1902,N_1476);
nand U2313 (N_2313,N_126,N_302);
nand U2314 (N_2314,N_1880,N_904);
xnor U2315 (N_2315,N_1594,N_295);
xor U2316 (N_2316,N_286,N_745);
nor U2317 (N_2317,N_1561,N_749);
or U2318 (N_2318,N_1639,N_897);
xnor U2319 (N_2319,N_39,N_777);
or U2320 (N_2320,N_311,N_1912);
nor U2321 (N_2321,N_1790,N_1283);
xnor U2322 (N_2322,N_948,N_202);
and U2323 (N_2323,N_900,N_732);
or U2324 (N_2324,N_1253,N_1100);
nand U2325 (N_2325,N_782,N_632);
or U2326 (N_2326,N_1553,N_1629);
nand U2327 (N_2327,N_570,N_189);
nand U2328 (N_2328,N_765,N_686);
nor U2329 (N_2329,N_1734,N_1981);
and U2330 (N_2330,N_918,N_16);
nor U2331 (N_2331,N_114,N_1462);
nor U2332 (N_2332,N_682,N_1420);
and U2333 (N_2333,N_577,N_976);
and U2334 (N_2334,N_1749,N_603);
or U2335 (N_2335,N_1430,N_1291);
nand U2336 (N_2336,N_119,N_1176);
or U2337 (N_2337,N_726,N_1101);
or U2338 (N_2338,N_212,N_339);
nand U2339 (N_2339,N_1091,N_610);
nor U2340 (N_2340,N_170,N_319);
or U2341 (N_2341,N_968,N_567);
or U2342 (N_2342,N_1424,N_1620);
nor U2343 (N_2343,N_1871,N_120);
xor U2344 (N_2344,N_201,N_312);
nand U2345 (N_2345,N_1158,N_1717);
xnor U2346 (N_2346,N_766,N_328);
and U2347 (N_2347,N_293,N_1488);
nor U2348 (N_2348,N_829,N_298);
xnor U2349 (N_2349,N_1445,N_89);
nor U2350 (N_2350,N_45,N_624);
nor U2351 (N_2351,N_1280,N_1210);
xor U2352 (N_2352,N_1645,N_1680);
nor U2353 (N_2353,N_102,N_875);
xor U2354 (N_2354,N_186,N_1168);
nand U2355 (N_2355,N_1016,N_1999);
xor U2356 (N_2356,N_411,N_932);
xnor U2357 (N_2357,N_1270,N_173);
xor U2358 (N_2358,N_758,N_1572);
nand U2359 (N_2359,N_1547,N_1427);
and U2360 (N_2360,N_1550,N_1055);
xnor U2361 (N_2361,N_1418,N_1578);
or U2362 (N_2362,N_198,N_1773);
nor U2363 (N_2363,N_485,N_1203);
and U2364 (N_2364,N_1018,N_335);
and U2365 (N_2365,N_1649,N_1066);
xor U2366 (N_2366,N_639,N_429);
xor U2367 (N_2367,N_946,N_1607);
nor U2368 (N_2368,N_468,N_977);
xor U2369 (N_2369,N_197,N_22);
and U2370 (N_2370,N_1668,N_504);
nand U2371 (N_2371,N_1141,N_142);
nor U2372 (N_2372,N_797,N_1021);
xnor U2373 (N_2373,N_408,N_1339);
and U2374 (N_2374,N_1047,N_1748);
xnor U2375 (N_2375,N_87,N_192);
or U2376 (N_2376,N_1357,N_19);
nor U2377 (N_2377,N_456,N_954);
and U2378 (N_2378,N_511,N_756);
nand U2379 (N_2379,N_348,N_4);
nand U2380 (N_2380,N_1755,N_957);
and U2381 (N_2381,N_1780,N_1987);
xnor U2382 (N_2382,N_12,N_731);
and U2383 (N_2383,N_31,N_736);
nor U2384 (N_2384,N_184,N_435);
nand U2385 (N_2385,N_813,N_98);
and U2386 (N_2386,N_1959,N_149);
xor U2387 (N_2387,N_1392,N_1556);
nor U2388 (N_2388,N_1049,N_1388);
and U2389 (N_2389,N_1148,N_1290);
nor U2390 (N_2390,N_1710,N_729);
nor U2391 (N_2391,N_1955,N_994);
nor U2392 (N_2392,N_1502,N_1306);
or U2393 (N_2393,N_1191,N_1583);
nand U2394 (N_2394,N_1754,N_1204);
nand U2395 (N_2395,N_428,N_1471);
nand U2396 (N_2396,N_1761,N_1361);
nor U2397 (N_2397,N_1437,N_773);
xor U2398 (N_2398,N_272,N_1461);
nor U2399 (N_2399,N_1984,N_23);
nand U2400 (N_2400,N_316,N_993);
nor U2401 (N_2401,N_1994,N_862);
and U2402 (N_2402,N_1200,N_1586);
nand U2403 (N_2403,N_1084,N_873);
and U2404 (N_2404,N_1321,N_289);
and U2405 (N_2405,N_1111,N_1269);
and U2406 (N_2406,N_890,N_1292);
nand U2407 (N_2407,N_1281,N_675);
and U2408 (N_2408,N_1409,N_1493);
xnor U2409 (N_2409,N_1707,N_383);
nor U2410 (N_2410,N_1608,N_460);
or U2411 (N_2411,N_556,N_1309);
nand U2412 (N_2412,N_86,N_291);
nand U2413 (N_2413,N_1605,N_1355);
xnor U2414 (N_2414,N_760,N_362);
nand U2415 (N_2415,N_1527,N_1500);
xor U2416 (N_2416,N_1262,N_872);
nor U2417 (N_2417,N_1568,N_810);
and U2418 (N_2418,N_214,N_334);
and U2419 (N_2419,N_1806,N_1772);
xor U2420 (N_2420,N_35,N_685);
or U2421 (N_2421,N_1767,N_448);
xnor U2422 (N_2422,N_1423,N_1900);
xnor U2423 (N_2423,N_478,N_1240);
or U2424 (N_2424,N_1536,N_1102);
nor U2425 (N_2425,N_746,N_1375);
nor U2426 (N_2426,N_1046,N_1085);
nor U2427 (N_2427,N_275,N_843);
nor U2428 (N_2428,N_583,N_1816);
nor U2429 (N_2429,N_1429,N_1944);
and U2430 (N_2430,N_1470,N_1294);
and U2431 (N_2431,N_244,N_1693);
xor U2432 (N_2432,N_1559,N_820);
nand U2433 (N_2433,N_347,N_653);
xor U2434 (N_2434,N_1075,N_1787);
xor U2435 (N_2435,N_1154,N_1171);
nor U2436 (N_2436,N_1827,N_1499);
nand U2437 (N_2437,N_678,N_223);
xor U2438 (N_2438,N_1876,N_1558);
or U2439 (N_2439,N_1867,N_1590);
nor U2440 (N_2440,N_1786,N_1718);
nand U2441 (N_2441,N_1831,N_238);
nor U2442 (N_2442,N_104,N_1333);
or U2443 (N_2443,N_1078,N_1636);
or U2444 (N_2444,N_737,N_326);
and U2445 (N_2445,N_105,N_1349);
xnor U2446 (N_2446,N_273,N_303);
xor U2447 (N_2447,N_1735,N_951);
and U2448 (N_2448,N_419,N_1634);
nor U2449 (N_2449,N_649,N_928);
or U2450 (N_2450,N_1918,N_1838);
and U2451 (N_2451,N_518,N_1968);
xor U2452 (N_2452,N_450,N_1797);
xnor U2453 (N_2453,N_1617,N_1962);
nand U2454 (N_2454,N_898,N_569);
xnor U2455 (N_2455,N_32,N_455);
nor U2456 (N_2456,N_739,N_1927);
nor U2457 (N_2457,N_638,N_288);
nand U2458 (N_2458,N_1223,N_1953);
and U2459 (N_2459,N_1036,N_1338);
xnor U2460 (N_2460,N_1130,N_153);
xnor U2461 (N_2461,N_1008,N_356);
or U2462 (N_2462,N_1487,N_43);
nand U2463 (N_2463,N_1798,N_91);
nor U2464 (N_2464,N_1575,N_27);
or U2465 (N_2465,N_1086,N_848);
and U2466 (N_2466,N_580,N_529);
nor U2467 (N_2467,N_1322,N_738);
or U2468 (N_2468,N_422,N_1692);
nand U2469 (N_2469,N_805,N_1644);
xnor U2470 (N_2470,N_1167,N_57);
and U2471 (N_2471,N_1785,N_1073);
xor U2472 (N_2472,N_107,N_1385);
and U2473 (N_2473,N_753,N_905);
nor U2474 (N_2474,N_1397,N_963);
nand U2475 (N_2475,N_1812,N_1225);
and U2476 (N_2476,N_705,N_1199);
nand U2477 (N_2477,N_1569,N_127);
and U2478 (N_2478,N_164,N_1989);
nand U2479 (N_2479,N_1161,N_935);
nand U2480 (N_2480,N_1793,N_195);
xnor U2481 (N_2481,N_1852,N_59);
nand U2482 (N_2482,N_1000,N_495);
and U2483 (N_2483,N_1543,N_690);
or U2484 (N_2484,N_239,N_1770);
xnor U2485 (N_2485,N_1898,N_962);
xnor U2486 (N_2486,N_243,N_836);
xor U2487 (N_2487,N_108,N_1893);
and U2488 (N_2488,N_1853,N_674);
xnor U2489 (N_2489,N_1901,N_755);
or U2490 (N_2490,N_1828,N_1390);
or U2491 (N_2491,N_1802,N_1737);
xnor U2492 (N_2492,N_1672,N_880);
and U2493 (N_2493,N_1308,N_553);
nor U2494 (N_2494,N_562,N_941);
nor U2495 (N_2495,N_394,N_117);
nand U2496 (N_2496,N_1760,N_717);
nand U2497 (N_2497,N_1973,N_1465);
nor U2498 (N_2498,N_524,N_711);
and U2499 (N_2499,N_1731,N_1384);
nand U2500 (N_2500,N_1165,N_990);
or U2501 (N_2501,N_475,N_725);
xnor U2502 (N_2502,N_1940,N_1267);
and U2503 (N_2503,N_1275,N_84);
and U2504 (N_2504,N_1170,N_1069);
or U2505 (N_2505,N_1971,N_1709);
and U2506 (N_2506,N_365,N_1525);
nand U2507 (N_2507,N_735,N_1263);
or U2508 (N_2508,N_617,N_1741);
or U2509 (N_2509,N_235,N_967);
and U2510 (N_2510,N_1642,N_774);
nand U2511 (N_2511,N_42,N_1413);
nand U2512 (N_2512,N_1667,N_78);
and U2513 (N_2513,N_226,N_157);
and U2514 (N_2514,N_785,N_892);
xnor U2515 (N_2515,N_262,N_1112);
and U2516 (N_2516,N_131,N_26);
nor U2517 (N_2517,N_743,N_1417);
or U2518 (N_2518,N_1751,N_1662);
and U2519 (N_2519,N_1746,N_1945);
and U2520 (N_2520,N_1699,N_208);
xnor U2521 (N_2521,N_1942,N_697);
or U2522 (N_2522,N_215,N_1350);
or U2523 (N_2523,N_1152,N_521);
and U2524 (N_2524,N_1421,N_613);
nand U2525 (N_2525,N_1474,N_595);
and U2526 (N_2526,N_676,N_1823);
xnor U2527 (N_2527,N_1555,N_519);
and U2528 (N_2528,N_382,N_1691);
or U2529 (N_2529,N_331,N_329);
and U2530 (N_2530,N_1162,N_135);
nor U2531 (N_2531,N_1630,N_492);
or U2532 (N_2532,N_225,N_474);
nor U2533 (N_2533,N_1140,N_155);
and U2534 (N_2534,N_1295,N_560);
xnor U2535 (N_2535,N_1221,N_1207);
nor U2536 (N_2536,N_1526,N_1195);
or U2537 (N_2537,N_1318,N_1126);
nor U2538 (N_2538,N_584,N_582);
and U2539 (N_2539,N_844,N_1554);
xor U2540 (N_2540,N_1467,N_156);
nand U2541 (N_2541,N_1401,N_863);
nand U2542 (N_2542,N_1933,N_1076);
nand U2543 (N_2543,N_1584,N_514);
xor U2544 (N_2544,N_592,N_1506);
xor U2545 (N_2545,N_310,N_806);
xor U2546 (N_2546,N_1234,N_516);
nand U2547 (N_2547,N_1451,N_1909);
xnor U2548 (N_2548,N_110,N_143);
xnor U2549 (N_2549,N_274,N_132);
nor U2550 (N_2550,N_913,N_1213);
or U2551 (N_2551,N_473,N_206);
nand U2552 (N_2552,N_1061,N_888);
nand U2553 (N_2553,N_200,N_1173);
nor U2554 (N_2554,N_634,N_1326);
nand U2555 (N_2555,N_970,N_895);
and U2556 (N_2556,N_261,N_118);
and U2557 (N_2557,N_1832,N_655);
and U2558 (N_2558,N_614,N_596);
and U2559 (N_2559,N_1386,N_748);
xor U2560 (N_2560,N_1532,N_1723);
nand U2561 (N_2561,N_49,N_1317);
and U2562 (N_2562,N_1434,N_1599);
or U2563 (N_2563,N_1906,N_876);
or U2564 (N_2564,N_608,N_681);
or U2565 (N_2565,N_1997,N_796);
or U2566 (N_2566,N_1611,N_723);
nor U2567 (N_2567,N_1929,N_611);
and U2568 (N_2568,N_80,N_1783);
or U2569 (N_2569,N_1587,N_525);
nor U2570 (N_2570,N_846,N_1539);
or U2571 (N_2571,N_554,N_190);
xnor U2572 (N_2572,N_1136,N_241);
xnor U2573 (N_2573,N_133,N_1779);
and U2574 (N_2574,N_1435,N_885);
xnor U2575 (N_2575,N_230,N_955);
or U2576 (N_2576,N_343,N_710);
xnor U2577 (N_2577,N_1172,N_1866);
xnor U2578 (N_2578,N_93,N_903);
nand U2579 (N_2579,N_1820,N_587);
and U2580 (N_2580,N_1518,N_1042);
and U2581 (N_2581,N_1851,N_1738);
or U2582 (N_2582,N_1700,N_1562);
nor U2583 (N_2583,N_907,N_1323);
xnor U2584 (N_2584,N_1026,N_1892);
nor U2585 (N_2585,N_277,N_1705);
and U2586 (N_2586,N_835,N_368);
nand U2587 (N_2587,N_1048,N_1352);
nor U2588 (N_2588,N_1229,N_607);
and U2589 (N_2589,N_1466,N_798);
xor U2590 (N_2590,N_1129,N_1004);
and U2591 (N_2591,N_598,N_433);
nand U2592 (N_2592,N_390,N_906);
or U2593 (N_2593,N_1730,N_670);
nand U2594 (N_2594,N_502,N_921);
and U2595 (N_2595,N_63,N_1135);
xnor U2596 (N_2596,N_444,N_66);
nand U2597 (N_2597,N_1678,N_1972);
or U2598 (N_2598,N_1733,N_1986);
xnor U2599 (N_2599,N_68,N_978);
or U2600 (N_2600,N_250,N_1879);
nor U2601 (N_2601,N_616,N_1480);
nor U2602 (N_2602,N_886,N_1618);
xor U2603 (N_2603,N_992,N_831);
nand U2604 (N_2604,N_1551,N_486);
xor U2605 (N_2605,N_1689,N_783);
or U2606 (N_2606,N_420,N_972);
and U2607 (N_2607,N_257,N_730);
or U2608 (N_2608,N_1877,N_1279);
or U2609 (N_2609,N_622,N_1521);
or U2610 (N_2610,N_1919,N_1932);
and U2611 (N_2611,N_351,N_1023);
xor U2612 (N_2612,N_989,N_1119);
nor U2613 (N_2613,N_927,N_1528);
nand U2614 (N_2614,N_692,N_874);
xnor U2615 (N_2615,N_923,N_816);
xor U2616 (N_2616,N_1183,N_1448);
nand U2617 (N_2617,N_801,N_1365);
and U2618 (N_2618,N_1083,N_430);
nand U2619 (N_2619,N_702,N_1624);
or U2620 (N_2620,N_1193,N_1044);
or U2621 (N_2621,N_454,N_561);
and U2622 (N_2622,N_1564,N_786);
nand U2623 (N_2623,N_1614,N_165);
nand U2624 (N_2624,N_680,N_618);
or U2625 (N_2625,N_1233,N_1928);
or U2626 (N_2626,N_207,N_1181);
xor U2627 (N_2627,N_13,N_1219);
xnor U2628 (N_2628,N_548,N_1345);
or U2629 (N_2629,N_1064,N_889);
or U2630 (N_2630,N_699,N_1655);
xor U2631 (N_2631,N_426,N_939);
or U2632 (N_2632,N_689,N_122);
xor U2633 (N_2633,N_389,N_802);
nand U2634 (N_2634,N_1298,N_1402);
nor U2635 (N_2635,N_662,N_1725);
and U2636 (N_2636,N_912,N_1348);
xor U2637 (N_2637,N_1288,N_1449);
and U2638 (N_2638,N_1301,N_590);
nor U2639 (N_2639,N_959,N_1878);
nand U2640 (N_2640,N_345,N_845);
xor U2641 (N_2641,N_400,N_825);
nand U2642 (N_2642,N_1387,N_1750);
and U2643 (N_2643,N_1671,N_695);
and U2644 (N_2644,N_20,N_263);
nor U2645 (N_2645,N_301,N_565);
or U2646 (N_2646,N_531,N_1914);
nand U2647 (N_2647,N_1284,N_1415);
nor U2648 (N_2648,N_1426,N_507);
nor U2649 (N_2649,N_147,N_150);
xor U2650 (N_2650,N_1379,N_211);
nor U2651 (N_2651,N_231,N_296);
or U2652 (N_2652,N_1576,N_1089);
and U2653 (N_2653,N_1593,N_1517);
nand U2654 (N_2654,N_1433,N_1704);
nor U2655 (N_2655,N_645,N_1603);
xor U2656 (N_2656,N_205,N_1988);
nand U2657 (N_2657,N_1481,N_82);
nor U2658 (N_2658,N_1904,N_513);
xnor U2659 (N_2659,N_517,N_283);
nand U2660 (N_2660,N_1656,N_1765);
and U2661 (N_2661,N_159,N_768);
nand U2662 (N_2662,N_1934,N_1809);
nand U2663 (N_2663,N_822,N_969);
xnor U2664 (N_2664,N_112,N_727);
or U2665 (N_2665,N_321,N_1304);
nor U2666 (N_2666,N_1247,N_1719);
xnor U2667 (N_2667,N_253,N_1063);
or U2668 (N_2668,N_1884,N_1778);
or U2669 (N_2669,N_1849,N_1907);
and U2670 (N_2670,N_716,N_1391);
or U2671 (N_2671,N_167,N_266);
and U2672 (N_2672,N_1540,N_1157);
and U2673 (N_2673,N_800,N_1665);
or U2674 (N_2674,N_859,N_1522);
or U2675 (N_2675,N_1664,N_973);
nand U2676 (N_2676,N_779,N_1163);
nor U2677 (N_2677,N_687,N_679);
or U2678 (N_2678,N_1715,N_1483);
nand U2679 (N_2679,N_1065,N_1272);
or U2680 (N_2680,N_1860,N_342);
or U2681 (N_2681,N_7,N_1567);
nand U2682 (N_2682,N_1485,N_669);
nor U2683 (N_2683,N_1582,N_1109);
nand U2684 (N_2684,N_1925,N_464);
nor U2685 (N_2685,N_637,N_1285);
nand U2686 (N_2686,N_609,N_1114);
nor U2687 (N_2687,N_866,N_1374);
xnor U2688 (N_2688,N_224,N_997);
xnor U2689 (N_2689,N_741,N_1155);
nand U2690 (N_2690,N_762,N_1473);
and U2691 (N_2691,N_706,N_1235);
and U2692 (N_2692,N_537,N_1224);
nor U2693 (N_2693,N_1312,N_359);
and U2694 (N_2694,N_1346,N_1589);
and U2695 (N_2695,N_1628,N_90);
or U2696 (N_2696,N_1616,N_242);
and U2697 (N_2697,N_656,N_1336);
xnor U2698 (N_2698,N_1895,N_926);
or U2699 (N_2699,N_1264,N_858);
nor U2700 (N_2700,N_986,N_597);
xor U2701 (N_2701,N_761,N_1251);
xnor U2702 (N_2702,N_971,N_1371);
xor U2703 (N_2703,N_268,N_1297);
xor U2704 (N_2704,N_666,N_183);
nor U2705 (N_2705,N_1137,N_1588);
nor U2706 (N_2706,N_1,N_501);
and U2707 (N_2707,N_1747,N_1996);
and U2708 (N_2708,N_367,N_899);
xnor U2709 (N_2709,N_576,N_552);
xnor U2710 (N_2710,N_75,N_1268);
or U2711 (N_2711,N_1964,N_427);
and U2712 (N_2712,N_1683,N_644);
nand U2713 (N_2713,N_1113,N_559);
nand U2714 (N_2714,N_1742,N_920);
xor U2715 (N_2715,N_499,N_1320);
and U2716 (N_2716,N_1769,N_1243);
and U2717 (N_2717,N_15,N_252);
and U2718 (N_2718,N_233,N_1147);
xor U2719 (N_2719,N_938,N_109);
xnor U2720 (N_2720,N_877,N_996);
or U2721 (N_2721,N_391,N_909);
nand U2722 (N_2722,N_1025,N_77);
nand U2723 (N_2723,N_887,N_371);
or U2724 (N_2724,N_1019,N_1856);
or U2725 (N_2725,N_1206,N_1396);
and U2726 (N_2726,N_55,N_1248);
xnor U2727 (N_2727,N_307,N_1923);
xor U2728 (N_2728,N_1781,N_833);
and U2729 (N_2729,N_95,N_696);
nor U2730 (N_2730,N_1108,N_1054);
and U2731 (N_2731,N_1530,N_870);
nand U2732 (N_2732,N_747,N_849);
or U2733 (N_2733,N_940,N_1600);
xnor U2734 (N_2734,N_1491,N_937);
or U2735 (N_2735,N_1970,N_1768);
or U2736 (N_2736,N_1237,N_1261);
nor U2737 (N_2737,N_659,N_1038);
xor U2738 (N_2738,N_103,N_40);
xnor U2739 (N_2739,N_1241,N_1340);
nand U2740 (N_2740,N_1728,N_396);
xor U2741 (N_2741,N_1650,N_1492);
nand U2742 (N_2742,N_1096,N_438);
nor U2743 (N_2743,N_1098,N_333);
nor U2744 (N_2744,N_1454,N_1903);
or U2745 (N_2745,N_1685,N_350);
xor U2746 (N_2746,N_914,N_1311);
and U2747 (N_2747,N_434,N_1360);
nand U2748 (N_2748,N_1040,N_1337);
nor U2749 (N_2749,N_1868,N_982);
and U2750 (N_2750,N_809,N_1523);
xor U2751 (N_2751,N_1419,N_671);
or U2752 (N_2752,N_278,N_540);
xor U2753 (N_2753,N_1560,N_575);
nand U2754 (N_2754,N_808,N_304);
nor U2755 (N_2755,N_965,N_1695);
and U2756 (N_2756,N_6,N_1186);
xor U2757 (N_2757,N_672,N_1694);
xor U2758 (N_2758,N_1194,N_1189);
nor U2759 (N_2759,N_728,N_1422);
nand U2760 (N_2760,N_148,N_1222);
and U2761 (N_2761,N_237,N_463);
and U2762 (N_2762,N_1541,N_1931);
nand U2763 (N_2763,N_1395,N_70);
and U2764 (N_2764,N_1463,N_1724);
and U2765 (N_2765,N_1146,N_1974);
xor U2766 (N_2766,N_360,N_1299);
or U2767 (N_2767,N_484,N_1808);
and U2768 (N_2768,N_384,N_1926);
xnor U2769 (N_2769,N_290,N_1960);
and U2770 (N_2770,N_526,N_1327);
nand U2771 (N_2771,N_1566,N_1436);
nor U2772 (N_2772,N_1514,N_1677);
nor U2773 (N_2773,N_789,N_917);
nor U2774 (N_2774,N_1242,N_101);
and U2775 (N_2775,N_1376,N_1505);
or U2776 (N_2776,N_1034,N_361);
or U2777 (N_2777,N_839,N_579);
nand U2778 (N_2778,N_1313,N_144);
nor U2779 (N_2779,N_308,N_29);
or U2780 (N_2780,N_1627,N_1882);
nand U2781 (N_2781,N_980,N_140);
or U2782 (N_2782,N_1625,N_324);
nand U2783 (N_2783,N_1508,N_557);
nand U2784 (N_2784,N_884,N_1690);
nand U2785 (N_2785,N_145,N_1344);
nor U2786 (N_2786,N_83,N_1455);
and U2787 (N_2787,N_1688,N_1829);
nor U2788 (N_2788,N_1216,N_373);
and U2789 (N_2789,N_1011,N_683);
xnor U2790 (N_2790,N_1074,N_1310);
and U2791 (N_2791,N_337,N_1939);
or U2792 (N_2792,N_431,N_46);
or U2793 (N_2793,N_1504,N_1670);
and U2794 (N_2794,N_494,N_952);
nand U2795 (N_2795,N_1638,N_1335);
nand U2796 (N_2796,N_1051,N_1708);
xor U2797 (N_2797,N_154,N_280);
nand U2798 (N_2798,N_228,N_1835);
or U2799 (N_2799,N_1428,N_1509);
nand U2800 (N_2800,N_313,N_981);
and U2801 (N_2801,N_1442,N_593);
and U2802 (N_2802,N_1097,N_1342);
nor U2803 (N_2803,N_1810,N_1328);
and U2804 (N_2804,N_1343,N_1815);
or U2805 (N_2805,N_1117,N_1453);
xor U2806 (N_2806,N_1957,N_1961);
and U2807 (N_2807,N_451,N_1585);
and U2808 (N_2808,N_1368,N_781);
nand U2809 (N_2809,N_34,N_642);
and U2810 (N_2810,N_574,N_1720);
nor U2811 (N_2811,N_1015,N_1794);
or U2812 (N_2812,N_139,N_281);
nand U2813 (N_2813,N_1300,N_386);
nand U2814 (N_2814,N_97,N_1180);
or U2815 (N_2815,N_834,N_1351);
nor U2816 (N_2816,N_1302,N_452);
nor U2817 (N_2817,N_523,N_1703);
nor U2818 (N_2818,N_1013,N_423);
or U2819 (N_2819,N_1515,N_1813);
and U2820 (N_2820,N_496,N_1673);
or U2821 (N_2821,N_417,N_1205);
nor U2822 (N_2822,N_1403,N_1949);
nand U2823 (N_2823,N_757,N_1841);
nor U2824 (N_2824,N_479,N_1675);
xor U2825 (N_2825,N_1602,N_1613);
or U2826 (N_2826,N_1118,N_232);
xor U2827 (N_2827,N_1801,N_33);
xnor U2828 (N_2828,N_1819,N_1142);
nand U2829 (N_2829,N_487,N_1524);
or U2830 (N_2830,N_443,N_466);
and U2831 (N_2831,N_358,N_1446);
xor U2832 (N_2832,N_1035,N_1935);
or U2833 (N_2833,N_902,N_387);
nand U2834 (N_2834,N_960,N_1510);
xor U2835 (N_2835,N_355,N_1353);
xnor U2836 (N_2836,N_1444,N_470);
or U2837 (N_2837,N_1020,N_1836);
or U2838 (N_2838,N_410,N_568);
nand U2839 (N_2839,N_838,N_987);
and U2840 (N_2840,N_218,N_81);
xnor U2841 (N_2841,N_1494,N_1400);
or U2842 (N_2842,N_1674,N_1992);
nand U2843 (N_2843,N_136,N_1125);
or U2844 (N_2844,N_958,N_483);
xor U2845 (N_2845,N_393,N_1887);
nor U2846 (N_2846,N_544,N_1658);
and U2847 (N_2847,N_469,N_1316);
nor U2848 (N_2848,N_1883,N_1862);
or U2849 (N_2849,N_1763,N_1166);
nand U2850 (N_2850,N_1438,N_1976);
nand U2851 (N_2851,N_620,N_814);
and U2852 (N_2852,N_48,N_2);
nand U2853 (N_2853,N_856,N_1752);
and U2854 (N_2854,N_1548,N_751);
nor U2855 (N_2855,N_1107,N_1889);
nand U2856 (N_2856,N_340,N_654);
xor U2857 (N_2857,N_5,N_129);
xor U2858 (N_2858,N_372,N_891);
and U2859 (N_2859,N_1029,N_1580);
and U2860 (N_2860,N_943,N_1053);
xnor U2861 (N_2861,N_1041,N_1998);
or U2862 (N_2862,N_1886,N_1503);
and U2863 (N_2863,N_636,N_1722);
nand U2864 (N_2864,N_332,N_1227);
or U2865 (N_2865,N_648,N_161);
xor U2866 (N_2866,N_172,N_1486);
or U2867 (N_2867,N_1854,N_374);
nand U2868 (N_2868,N_535,N_1764);
or U2869 (N_2869,N_265,N_661);
nand U2870 (N_2870,N_1758,N_1535);
xnor U2871 (N_2871,N_667,N_1921);
xor U2872 (N_2872,N_1458,N_398);
xor U2873 (N_2873,N_188,N_395);
and U2874 (N_2874,N_294,N_1684);
and U2875 (N_2875,N_493,N_1496);
or U2876 (N_2876,N_1138,N_1489);
or U2877 (N_2877,N_471,N_668);
or U2878 (N_2878,N_1095,N_179);
and U2879 (N_2879,N_1637,N_868);
xor U2880 (N_2880,N_1398,N_572);
xnor U2881 (N_2881,N_983,N_69);
or U2882 (N_2882,N_1372,N_1087);
or U2883 (N_2883,N_141,N_370);
or U2884 (N_2884,N_1622,N_1905);
and U2885 (N_2885,N_1457,N_106);
and U2886 (N_2886,N_1027,N_1156);
nand U2887 (N_2887,N_217,N_187);
or U2888 (N_2888,N_944,N_1727);
xor U2889 (N_2889,N_1177,N_1347);
nor U2890 (N_2890,N_1930,N_425);
or U2891 (N_2891,N_1093,N_453);
nand U2892 (N_2892,N_606,N_850);
xor U2893 (N_2893,N_113,N_497);
nand U2894 (N_2894,N_1552,N_1894);
or U2895 (N_2895,N_633,N_1598);
or U2896 (N_2896,N_505,N_1721);
or U2897 (N_2897,N_1056,N_528);
xor U2898 (N_2898,N_586,N_1077);
nor U2899 (N_2899,N_985,N_1745);
xor U2900 (N_2900,N_621,N_1911);
nand U2901 (N_2901,N_1259,N_627);
and U2902 (N_2902,N_1609,N_377);
nor U2903 (N_2903,N_255,N_720);
nor U2904 (N_2904,N_979,N_950);
and U2905 (N_2905,N_919,N_1821);
or U2906 (N_2906,N_1660,N_1145);
and U2907 (N_2907,N_1805,N_67);
and U2908 (N_2908,N_538,N_555);
or U2909 (N_2909,N_1153,N_1885);
and U2910 (N_2910,N_1632,N_700);
xor U2911 (N_2911,N_794,N_515);
or U2912 (N_2912,N_1830,N_663);
nor U2913 (N_2913,N_1512,N_1711);
or U2914 (N_2914,N_1404,N_305);
nand U2915 (N_2915,N_1537,N_910);
nand U2916 (N_2916,N_1982,N_1070);
nand U2917 (N_2917,N_646,N_1771);
or U2918 (N_2918,N_1943,N_824);
nand U2919 (N_2919,N_1542,N_1007);
or U2920 (N_2920,N_378,N_94);
nand U2921 (N_2921,N_491,N_37);
xnor U2922 (N_2922,N_364,N_1563);
nor U2923 (N_2923,N_1833,N_1706);
xnor U2924 (N_2924,N_1916,N_1017);
or U2925 (N_2925,N_701,N_1843);
and U2926 (N_2926,N_1128,N_772);
xnor U2927 (N_2927,N_1701,N_1822);
xor U2928 (N_2928,N_1966,N_162);
and U2929 (N_2929,N_171,N_916);
or U2930 (N_2930,N_375,N_1459);
nand U2931 (N_2931,N_1037,N_1941);
nand U2932 (N_2932,N_974,N_1287);
xnor U2933 (N_2933,N_18,N_1059);
nor U2934 (N_2934,N_403,N_936);
xor U2935 (N_2935,N_864,N_1362);
nand U2936 (N_2936,N_1920,N_168);
and U2937 (N_2937,N_1915,N_1811);
nand U2938 (N_2938,N_1226,N_1197);
and U2939 (N_2939,N_1286,N_53);
nand U2940 (N_2940,N_1951,N_1872);
or U2941 (N_2941,N_594,N_1358);
xnor U2942 (N_2942,N_1211,N_1252);
nor U2943 (N_2943,N_817,N_1696);
or U2944 (N_2944,N_930,N_1143);
nand U2945 (N_2945,N_182,N_363);
and U2946 (N_2946,N_209,N_1681);
nand U2947 (N_2947,N_1208,N_1005);
nor U2948 (N_2948,N_234,N_1947);
or U2949 (N_2949,N_795,N_1273);
and U2950 (N_2950,N_92,N_1557);
nor U2951 (N_2951,N_995,N_146);
and U2952 (N_2952,N_956,N_488);
xor U2953 (N_2953,N_17,N_1472);
nand U2954 (N_2954,N_1965,N_1393);
xnor U2955 (N_2955,N_1766,N_619);
and U2956 (N_2956,N_1870,N_1937);
or U2957 (N_2957,N_421,N_445);
nand U2958 (N_2958,N_1631,N_803);
nand U2959 (N_2959,N_1250,N_1068);
nor U2960 (N_2960,N_787,N_1814);
nand U2961 (N_2961,N_869,N_446);
nand U2962 (N_2962,N_72,N_64);
or U2963 (N_2963,N_925,N_1192);
or U2964 (N_2964,N_1531,N_51);
nand U2965 (N_2965,N_1238,N_52);
and U2966 (N_2966,N_1762,N_550);
and U2967 (N_2967,N_1050,N_1817);
and U2968 (N_2968,N_509,N_158);
nor U2969 (N_2969,N_1716,N_320);
or U2970 (N_2970,N_1246,N_1122);
nor U2971 (N_2971,N_571,N_1188);
or U2972 (N_2972,N_1511,N_714);
and U2973 (N_2973,N_1641,N_1330);
nand U2974 (N_2974,N_770,N_1875);
or U2975 (N_2975,N_1067,N_1574);
and U2976 (N_2976,N_1623,N_1120);
xnor U2977 (N_2977,N_174,N_1577);
nand U2978 (N_2978,N_115,N_151);
nand U2979 (N_2979,N_254,N_1307);
or U2980 (N_2980,N_1687,N_111);
and U2981 (N_2981,N_1159,N_933);
nand U2982 (N_2982,N_1533,N_402);
nor U2983 (N_2983,N_1202,N_1258);
nand U2984 (N_2984,N_1839,N_791);
and U2985 (N_2985,N_832,N_100);
nor U2986 (N_2986,N_1661,N_626);
or U2987 (N_2987,N_1139,N_1447);
or U2988 (N_2988,N_1484,N_1963);
nor U2989 (N_2989,N_247,N_1874);
nand U2990 (N_2990,N_975,N_251);
or U2991 (N_2991,N_1888,N_931);
xnor U2992 (N_2992,N_628,N_1257);
and U2993 (N_2993,N_1127,N_99);
and U2994 (N_2994,N_929,N_276);
nor U2995 (N_2995,N_194,N_1440);
and U2996 (N_2996,N_1908,N_545);
and U2997 (N_2997,N_1619,N_881);
nor U2998 (N_2998,N_1033,N_1012);
nand U2999 (N_2999,N_1105,N_698);
nor U3000 (N_3000,N_681,N_554);
xnor U3001 (N_3001,N_611,N_249);
and U3002 (N_3002,N_786,N_47);
nor U3003 (N_3003,N_1220,N_1629);
and U3004 (N_3004,N_735,N_555);
nor U3005 (N_3005,N_239,N_418);
nand U3006 (N_3006,N_1761,N_1826);
nand U3007 (N_3007,N_1227,N_562);
and U3008 (N_3008,N_1439,N_614);
nand U3009 (N_3009,N_1080,N_1691);
nor U3010 (N_3010,N_1191,N_1570);
nor U3011 (N_3011,N_895,N_925);
and U3012 (N_3012,N_922,N_501);
or U3013 (N_3013,N_1439,N_1168);
xor U3014 (N_3014,N_202,N_1253);
nor U3015 (N_3015,N_1057,N_158);
and U3016 (N_3016,N_751,N_1207);
nand U3017 (N_3017,N_1130,N_1873);
or U3018 (N_3018,N_1265,N_562);
and U3019 (N_3019,N_1429,N_683);
xor U3020 (N_3020,N_1170,N_1221);
or U3021 (N_3021,N_816,N_1095);
or U3022 (N_3022,N_201,N_1836);
or U3023 (N_3023,N_664,N_1033);
and U3024 (N_3024,N_1826,N_1164);
nand U3025 (N_3025,N_1255,N_611);
or U3026 (N_3026,N_617,N_1351);
xor U3027 (N_3027,N_1777,N_633);
nor U3028 (N_3028,N_1593,N_468);
and U3029 (N_3029,N_1403,N_1525);
xnor U3030 (N_3030,N_971,N_1277);
xnor U3031 (N_3031,N_62,N_815);
or U3032 (N_3032,N_1624,N_1110);
xor U3033 (N_3033,N_244,N_947);
xnor U3034 (N_3034,N_1662,N_1409);
nand U3035 (N_3035,N_1620,N_887);
nor U3036 (N_3036,N_355,N_366);
and U3037 (N_3037,N_865,N_1284);
and U3038 (N_3038,N_1826,N_1525);
and U3039 (N_3039,N_78,N_1622);
and U3040 (N_3040,N_1029,N_791);
and U3041 (N_3041,N_14,N_1471);
xnor U3042 (N_3042,N_1025,N_1112);
xnor U3043 (N_3043,N_878,N_1095);
nor U3044 (N_3044,N_1281,N_882);
or U3045 (N_3045,N_948,N_164);
or U3046 (N_3046,N_1702,N_586);
nand U3047 (N_3047,N_5,N_530);
xor U3048 (N_3048,N_354,N_320);
xnor U3049 (N_3049,N_1469,N_661);
xor U3050 (N_3050,N_1537,N_1938);
xnor U3051 (N_3051,N_898,N_773);
nor U3052 (N_3052,N_902,N_1362);
nor U3053 (N_3053,N_737,N_541);
nor U3054 (N_3054,N_1882,N_179);
or U3055 (N_3055,N_626,N_1164);
nand U3056 (N_3056,N_905,N_137);
and U3057 (N_3057,N_852,N_1985);
nand U3058 (N_3058,N_1942,N_1731);
nand U3059 (N_3059,N_128,N_1210);
nand U3060 (N_3060,N_996,N_129);
or U3061 (N_3061,N_691,N_140);
and U3062 (N_3062,N_1902,N_322);
nor U3063 (N_3063,N_749,N_1760);
and U3064 (N_3064,N_27,N_432);
and U3065 (N_3065,N_1534,N_1472);
and U3066 (N_3066,N_282,N_1877);
nor U3067 (N_3067,N_1738,N_1491);
nor U3068 (N_3068,N_1033,N_123);
nand U3069 (N_3069,N_182,N_1015);
xnor U3070 (N_3070,N_772,N_198);
xnor U3071 (N_3071,N_1077,N_464);
nor U3072 (N_3072,N_515,N_1487);
xnor U3073 (N_3073,N_110,N_1853);
or U3074 (N_3074,N_674,N_1283);
nor U3075 (N_3075,N_1761,N_614);
and U3076 (N_3076,N_1171,N_545);
nand U3077 (N_3077,N_1621,N_1780);
or U3078 (N_3078,N_635,N_176);
and U3079 (N_3079,N_485,N_739);
nand U3080 (N_3080,N_1223,N_1191);
or U3081 (N_3081,N_1861,N_324);
nor U3082 (N_3082,N_758,N_846);
xor U3083 (N_3083,N_1669,N_1800);
nor U3084 (N_3084,N_786,N_341);
and U3085 (N_3085,N_1554,N_1957);
nor U3086 (N_3086,N_149,N_990);
nand U3087 (N_3087,N_46,N_1826);
xnor U3088 (N_3088,N_1633,N_596);
and U3089 (N_3089,N_1625,N_406);
xnor U3090 (N_3090,N_1131,N_1153);
or U3091 (N_3091,N_289,N_1457);
and U3092 (N_3092,N_1053,N_95);
or U3093 (N_3093,N_1978,N_477);
nand U3094 (N_3094,N_1387,N_47);
nand U3095 (N_3095,N_1486,N_96);
or U3096 (N_3096,N_1545,N_116);
and U3097 (N_3097,N_177,N_687);
xnor U3098 (N_3098,N_309,N_1979);
or U3099 (N_3099,N_949,N_1655);
nand U3100 (N_3100,N_1839,N_1479);
nand U3101 (N_3101,N_1250,N_759);
nand U3102 (N_3102,N_1299,N_609);
nor U3103 (N_3103,N_1240,N_1698);
and U3104 (N_3104,N_1490,N_423);
nor U3105 (N_3105,N_57,N_640);
nor U3106 (N_3106,N_1027,N_1313);
nor U3107 (N_3107,N_552,N_45);
xnor U3108 (N_3108,N_1902,N_706);
nand U3109 (N_3109,N_561,N_380);
xor U3110 (N_3110,N_322,N_1047);
xor U3111 (N_3111,N_397,N_315);
and U3112 (N_3112,N_1449,N_966);
or U3113 (N_3113,N_230,N_163);
or U3114 (N_3114,N_1607,N_861);
and U3115 (N_3115,N_458,N_1510);
nand U3116 (N_3116,N_113,N_1044);
and U3117 (N_3117,N_253,N_1985);
and U3118 (N_3118,N_1345,N_255);
or U3119 (N_3119,N_1372,N_1808);
nor U3120 (N_3120,N_897,N_1874);
nor U3121 (N_3121,N_1960,N_1243);
xnor U3122 (N_3122,N_406,N_1466);
nor U3123 (N_3123,N_296,N_169);
xor U3124 (N_3124,N_628,N_1269);
xnor U3125 (N_3125,N_1663,N_623);
nor U3126 (N_3126,N_1731,N_1955);
or U3127 (N_3127,N_1734,N_1436);
xnor U3128 (N_3128,N_1791,N_1022);
or U3129 (N_3129,N_1974,N_497);
or U3130 (N_3130,N_1667,N_652);
xnor U3131 (N_3131,N_613,N_129);
nand U3132 (N_3132,N_289,N_1650);
xor U3133 (N_3133,N_760,N_1854);
xor U3134 (N_3134,N_763,N_1581);
nand U3135 (N_3135,N_1182,N_693);
or U3136 (N_3136,N_1314,N_1956);
or U3137 (N_3137,N_1201,N_517);
nand U3138 (N_3138,N_345,N_1866);
xor U3139 (N_3139,N_1845,N_143);
and U3140 (N_3140,N_1889,N_1850);
or U3141 (N_3141,N_1328,N_1565);
or U3142 (N_3142,N_206,N_1248);
nand U3143 (N_3143,N_567,N_495);
and U3144 (N_3144,N_121,N_1696);
xor U3145 (N_3145,N_1034,N_1680);
and U3146 (N_3146,N_565,N_1133);
nor U3147 (N_3147,N_80,N_1781);
xnor U3148 (N_3148,N_219,N_1796);
nor U3149 (N_3149,N_1789,N_1268);
xor U3150 (N_3150,N_319,N_743);
and U3151 (N_3151,N_1439,N_1029);
nand U3152 (N_3152,N_209,N_1635);
nor U3153 (N_3153,N_867,N_1192);
and U3154 (N_3154,N_1885,N_1839);
nor U3155 (N_3155,N_847,N_895);
xor U3156 (N_3156,N_1679,N_530);
nand U3157 (N_3157,N_1660,N_958);
and U3158 (N_3158,N_1074,N_388);
nand U3159 (N_3159,N_864,N_439);
xor U3160 (N_3160,N_378,N_985);
or U3161 (N_3161,N_1857,N_1011);
and U3162 (N_3162,N_1564,N_1107);
nand U3163 (N_3163,N_1238,N_1719);
nor U3164 (N_3164,N_705,N_1994);
nand U3165 (N_3165,N_1366,N_676);
and U3166 (N_3166,N_851,N_992);
nand U3167 (N_3167,N_940,N_865);
nand U3168 (N_3168,N_1400,N_970);
and U3169 (N_3169,N_114,N_192);
nand U3170 (N_3170,N_1532,N_1059);
xnor U3171 (N_3171,N_1706,N_876);
nor U3172 (N_3172,N_742,N_1731);
nor U3173 (N_3173,N_242,N_358);
or U3174 (N_3174,N_611,N_1661);
or U3175 (N_3175,N_642,N_122);
nor U3176 (N_3176,N_1918,N_1698);
and U3177 (N_3177,N_1381,N_1214);
nand U3178 (N_3178,N_429,N_1584);
nor U3179 (N_3179,N_1290,N_103);
xor U3180 (N_3180,N_354,N_434);
and U3181 (N_3181,N_1172,N_1365);
xnor U3182 (N_3182,N_180,N_1418);
and U3183 (N_3183,N_1222,N_46);
xor U3184 (N_3184,N_127,N_108);
nor U3185 (N_3185,N_234,N_74);
or U3186 (N_3186,N_884,N_602);
xnor U3187 (N_3187,N_484,N_84);
and U3188 (N_3188,N_1648,N_1580);
and U3189 (N_3189,N_1751,N_218);
nand U3190 (N_3190,N_159,N_267);
nand U3191 (N_3191,N_976,N_369);
nand U3192 (N_3192,N_394,N_37);
xor U3193 (N_3193,N_1409,N_342);
nand U3194 (N_3194,N_736,N_1389);
and U3195 (N_3195,N_1936,N_714);
and U3196 (N_3196,N_1377,N_878);
or U3197 (N_3197,N_1099,N_379);
nor U3198 (N_3198,N_963,N_874);
and U3199 (N_3199,N_1005,N_1649);
nor U3200 (N_3200,N_1211,N_1994);
nor U3201 (N_3201,N_1481,N_1012);
nor U3202 (N_3202,N_1621,N_1677);
and U3203 (N_3203,N_1756,N_967);
or U3204 (N_3204,N_554,N_829);
or U3205 (N_3205,N_1780,N_950);
or U3206 (N_3206,N_1304,N_232);
xor U3207 (N_3207,N_281,N_178);
nor U3208 (N_3208,N_1204,N_1835);
nor U3209 (N_3209,N_456,N_1863);
nand U3210 (N_3210,N_1391,N_1296);
or U3211 (N_3211,N_1704,N_1804);
or U3212 (N_3212,N_357,N_1884);
nor U3213 (N_3213,N_372,N_500);
xor U3214 (N_3214,N_872,N_662);
nand U3215 (N_3215,N_1330,N_1911);
xnor U3216 (N_3216,N_1445,N_1474);
and U3217 (N_3217,N_829,N_16);
xnor U3218 (N_3218,N_384,N_650);
or U3219 (N_3219,N_622,N_713);
or U3220 (N_3220,N_866,N_576);
nor U3221 (N_3221,N_662,N_1550);
or U3222 (N_3222,N_1010,N_1372);
nand U3223 (N_3223,N_1106,N_662);
xor U3224 (N_3224,N_724,N_1382);
or U3225 (N_3225,N_1447,N_1793);
xnor U3226 (N_3226,N_1616,N_566);
and U3227 (N_3227,N_1615,N_1213);
and U3228 (N_3228,N_365,N_1408);
nor U3229 (N_3229,N_786,N_750);
nand U3230 (N_3230,N_965,N_1518);
nor U3231 (N_3231,N_1648,N_889);
or U3232 (N_3232,N_1284,N_1536);
or U3233 (N_3233,N_1248,N_1905);
or U3234 (N_3234,N_133,N_1832);
or U3235 (N_3235,N_1073,N_115);
or U3236 (N_3236,N_1473,N_1500);
or U3237 (N_3237,N_1940,N_520);
nor U3238 (N_3238,N_593,N_785);
nor U3239 (N_3239,N_1376,N_933);
nand U3240 (N_3240,N_70,N_265);
xnor U3241 (N_3241,N_197,N_1068);
xor U3242 (N_3242,N_154,N_304);
nor U3243 (N_3243,N_467,N_614);
and U3244 (N_3244,N_291,N_131);
xnor U3245 (N_3245,N_897,N_1844);
nand U3246 (N_3246,N_1880,N_1737);
and U3247 (N_3247,N_640,N_833);
and U3248 (N_3248,N_877,N_964);
xnor U3249 (N_3249,N_292,N_198);
nand U3250 (N_3250,N_1721,N_1252);
or U3251 (N_3251,N_1919,N_1908);
nor U3252 (N_3252,N_409,N_1844);
and U3253 (N_3253,N_1341,N_1373);
xor U3254 (N_3254,N_623,N_384);
xnor U3255 (N_3255,N_1992,N_390);
or U3256 (N_3256,N_578,N_771);
and U3257 (N_3257,N_1045,N_813);
or U3258 (N_3258,N_1869,N_1132);
xor U3259 (N_3259,N_1536,N_735);
nor U3260 (N_3260,N_847,N_411);
nand U3261 (N_3261,N_588,N_310);
or U3262 (N_3262,N_234,N_1909);
nand U3263 (N_3263,N_1993,N_150);
xor U3264 (N_3264,N_573,N_556);
nand U3265 (N_3265,N_924,N_1632);
and U3266 (N_3266,N_1569,N_515);
or U3267 (N_3267,N_118,N_487);
xor U3268 (N_3268,N_648,N_79);
nor U3269 (N_3269,N_764,N_554);
or U3270 (N_3270,N_275,N_1903);
or U3271 (N_3271,N_93,N_1528);
and U3272 (N_3272,N_1085,N_1095);
xnor U3273 (N_3273,N_909,N_1086);
nand U3274 (N_3274,N_1014,N_1707);
or U3275 (N_3275,N_1158,N_1379);
or U3276 (N_3276,N_546,N_1483);
or U3277 (N_3277,N_1279,N_1116);
xnor U3278 (N_3278,N_923,N_1341);
nor U3279 (N_3279,N_668,N_1420);
and U3280 (N_3280,N_1134,N_1809);
nand U3281 (N_3281,N_1341,N_140);
and U3282 (N_3282,N_1389,N_110);
nor U3283 (N_3283,N_460,N_474);
nor U3284 (N_3284,N_821,N_461);
or U3285 (N_3285,N_1230,N_192);
and U3286 (N_3286,N_886,N_1858);
nand U3287 (N_3287,N_1471,N_1180);
or U3288 (N_3288,N_218,N_1285);
nand U3289 (N_3289,N_1418,N_162);
xor U3290 (N_3290,N_1910,N_1848);
or U3291 (N_3291,N_317,N_531);
xnor U3292 (N_3292,N_963,N_299);
nor U3293 (N_3293,N_297,N_961);
nor U3294 (N_3294,N_799,N_1900);
or U3295 (N_3295,N_1372,N_494);
xnor U3296 (N_3296,N_1444,N_474);
xnor U3297 (N_3297,N_37,N_1544);
xor U3298 (N_3298,N_741,N_1602);
and U3299 (N_3299,N_810,N_1059);
nor U3300 (N_3300,N_1750,N_685);
or U3301 (N_3301,N_1056,N_762);
and U3302 (N_3302,N_892,N_1153);
nand U3303 (N_3303,N_140,N_904);
nor U3304 (N_3304,N_1220,N_227);
nand U3305 (N_3305,N_1383,N_1284);
or U3306 (N_3306,N_1326,N_400);
or U3307 (N_3307,N_541,N_57);
or U3308 (N_3308,N_0,N_881);
xnor U3309 (N_3309,N_1425,N_559);
xnor U3310 (N_3310,N_1806,N_1263);
or U3311 (N_3311,N_198,N_1830);
or U3312 (N_3312,N_363,N_1270);
or U3313 (N_3313,N_1821,N_1942);
xor U3314 (N_3314,N_915,N_1008);
and U3315 (N_3315,N_773,N_1954);
xnor U3316 (N_3316,N_395,N_55);
nor U3317 (N_3317,N_1785,N_1253);
and U3318 (N_3318,N_962,N_1490);
and U3319 (N_3319,N_269,N_1892);
xor U3320 (N_3320,N_185,N_1227);
xnor U3321 (N_3321,N_1024,N_820);
nor U3322 (N_3322,N_89,N_1470);
xnor U3323 (N_3323,N_41,N_667);
nor U3324 (N_3324,N_1352,N_1626);
or U3325 (N_3325,N_812,N_600);
xnor U3326 (N_3326,N_718,N_1992);
nor U3327 (N_3327,N_1776,N_1020);
and U3328 (N_3328,N_1122,N_1386);
or U3329 (N_3329,N_369,N_931);
xnor U3330 (N_3330,N_1153,N_1700);
and U3331 (N_3331,N_1222,N_1595);
nor U3332 (N_3332,N_395,N_1031);
xnor U3333 (N_3333,N_1624,N_247);
xnor U3334 (N_3334,N_454,N_1061);
nand U3335 (N_3335,N_939,N_954);
nand U3336 (N_3336,N_1211,N_1631);
or U3337 (N_3337,N_598,N_1669);
xor U3338 (N_3338,N_836,N_1885);
nor U3339 (N_3339,N_807,N_1332);
xor U3340 (N_3340,N_1891,N_262);
nor U3341 (N_3341,N_1382,N_1094);
and U3342 (N_3342,N_1711,N_481);
xnor U3343 (N_3343,N_1133,N_1295);
nor U3344 (N_3344,N_1014,N_1567);
nand U3345 (N_3345,N_541,N_621);
nand U3346 (N_3346,N_1657,N_1949);
xor U3347 (N_3347,N_1490,N_899);
and U3348 (N_3348,N_956,N_163);
or U3349 (N_3349,N_1153,N_961);
nand U3350 (N_3350,N_752,N_1256);
nand U3351 (N_3351,N_1612,N_916);
nor U3352 (N_3352,N_1428,N_418);
or U3353 (N_3353,N_1686,N_402);
nor U3354 (N_3354,N_397,N_340);
nor U3355 (N_3355,N_1960,N_753);
or U3356 (N_3356,N_412,N_1526);
and U3357 (N_3357,N_295,N_1593);
nand U3358 (N_3358,N_219,N_1070);
nand U3359 (N_3359,N_1930,N_662);
and U3360 (N_3360,N_1133,N_1518);
nor U3361 (N_3361,N_1769,N_715);
nor U3362 (N_3362,N_1108,N_809);
xor U3363 (N_3363,N_1360,N_188);
nor U3364 (N_3364,N_777,N_1845);
xnor U3365 (N_3365,N_1159,N_1219);
xor U3366 (N_3366,N_1035,N_890);
xnor U3367 (N_3367,N_1723,N_1872);
nand U3368 (N_3368,N_1086,N_1042);
nor U3369 (N_3369,N_1410,N_395);
nand U3370 (N_3370,N_1570,N_1772);
xnor U3371 (N_3371,N_1687,N_1154);
or U3372 (N_3372,N_249,N_983);
or U3373 (N_3373,N_353,N_163);
nand U3374 (N_3374,N_663,N_605);
xnor U3375 (N_3375,N_1771,N_326);
or U3376 (N_3376,N_1353,N_1119);
and U3377 (N_3377,N_188,N_644);
and U3378 (N_3378,N_866,N_138);
nand U3379 (N_3379,N_1910,N_570);
or U3380 (N_3380,N_1492,N_1556);
xor U3381 (N_3381,N_1206,N_651);
or U3382 (N_3382,N_577,N_559);
nor U3383 (N_3383,N_323,N_1671);
and U3384 (N_3384,N_1242,N_409);
xor U3385 (N_3385,N_1925,N_250);
nand U3386 (N_3386,N_538,N_1916);
nor U3387 (N_3387,N_1201,N_210);
nor U3388 (N_3388,N_854,N_1899);
nor U3389 (N_3389,N_1064,N_304);
xnor U3390 (N_3390,N_1510,N_1964);
and U3391 (N_3391,N_5,N_1812);
nor U3392 (N_3392,N_741,N_1369);
nor U3393 (N_3393,N_512,N_451);
nor U3394 (N_3394,N_1852,N_486);
nor U3395 (N_3395,N_738,N_494);
nor U3396 (N_3396,N_432,N_344);
xor U3397 (N_3397,N_832,N_514);
and U3398 (N_3398,N_931,N_1396);
nor U3399 (N_3399,N_1189,N_903);
or U3400 (N_3400,N_1275,N_1473);
or U3401 (N_3401,N_1983,N_1796);
and U3402 (N_3402,N_579,N_272);
and U3403 (N_3403,N_436,N_471);
nand U3404 (N_3404,N_1840,N_278);
xor U3405 (N_3405,N_1291,N_835);
xnor U3406 (N_3406,N_1465,N_1207);
xnor U3407 (N_3407,N_1312,N_565);
or U3408 (N_3408,N_1713,N_972);
and U3409 (N_3409,N_536,N_1990);
and U3410 (N_3410,N_1488,N_1260);
or U3411 (N_3411,N_1085,N_151);
xnor U3412 (N_3412,N_1270,N_890);
and U3413 (N_3413,N_1422,N_338);
and U3414 (N_3414,N_1665,N_1483);
nor U3415 (N_3415,N_1780,N_71);
xnor U3416 (N_3416,N_526,N_1498);
nand U3417 (N_3417,N_1164,N_61);
and U3418 (N_3418,N_740,N_1219);
xor U3419 (N_3419,N_649,N_253);
nor U3420 (N_3420,N_541,N_510);
and U3421 (N_3421,N_1827,N_1977);
nand U3422 (N_3422,N_1262,N_1822);
nor U3423 (N_3423,N_1422,N_559);
nand U3424 (N_3424,N_1300,N_104);
or U3425 (N_3425,N_705,N_743);
nand U3426 (N_3426,N_1606,N_581);
and U3427 (N_3427,N_405,N_342);
xor U3428 (N_3428,N_157,N_80);
xor U3429 (N_3429,N_1938,N_748);
xor U3430 (N_3430,N_1607,N_822);
or U3431 (N_3431,N_1513,N_489);
nand U3432 (N_3432,N_312,N_1441);
nand U3433 (N_3433,N_33,N_55);
nor U3434 (N_3434,N_762,N_981);
nor U3435 (N_3435,N_1005,N_429);
nor U3436 (N_3436,N_1860,N_564);
nor U3437 (N_3437,N_1470,N_978);
xor U3438 (N_3438,N_1475,N_107);
and U3439 (N_3439,N_1234,N_1494);
nand U3440 (N_3440,N_643,N_1898);
xnor U3441 (N_3441,N_1072,N_30);
xor U3442 (N_3442,N_814,N_1856);
nor U3443 (N_3443,N_1662,N_1530);
or U3444 (N_3444,N_1241,N_987);
nor U3445 (N_3445,N_598,N_172);
or U3446 (N_3446,N_333,N_1874);
nand U3447 (N_3447,N_1503,N_219);
or U3448 (N_3448,N_119,N_365);
xor U3449 (N_3449,N_575,N_696);
or U3450 (N_3450,N_446,N_889);
or U3451 (N_3451,N_1545,N_1422);
nand U3452 (N_3452,N_248,N_1375);
and U3453 (N_3453,N_1405,N_439);
nand U3454 (N_3454,N_1932,N_743);
nand U3455 (N_3455,N_1699,N_1961);
nand U3456 (N_3456,N_1827,N_1151);
nor U3457 (N_3457,N_595,N_1704);
nor U3458 (N_3458,N_1615,N_904);
nor U3459 (N_3459,N_1021,N_435);
nor U3460 (N_3460,N_1702,N_53);
nand U3461 (N_3461,N_1947,N_294);
nand U3462 (N_3462,N_173,N_1867);
nand U3463 (N_3463,N_332,N_1990);
or U3464 (N_3464,N_144,N_1526);
or U3465 (N_3465,N_1004,N_993);
nand U3466 (N_3466,N_438,N_271);
and U3467 (N_3467,N_952,N_947);
nor U3468 (N_3468,N_502,N_422);
nor U3469 (N_3469,N_1035,N_966);
or U3470 (N_3470,N_1605,N_347);
nand U3471 (N_3471,N_87,N_385);
and U3472 (N_3472,N_1927,N_723);
and U3473 (N_3473,N_1747,N_1644);
or U3474 (N_3474,N_387,N_1495);
or U3475 (N_3475,N_1478,N_1658);
nor U3476 (N_3476,N_70,N_1724);
nor U3477 (N_3477,N_1971,N_1575);
xor U3478 (N_3478,N_1699,N_1167);
nor U3479 (N_3479,N_1598,N_1729);
nand U3480 (N_3480,N_1627,N_1932);
or U3481 (N_3481,N_359,N_964);
and U3482 (N_3482,N_1136,N_456);
nor U3483 (N_3483,N_358,N_236);
and U3484 (N_3484,N_519,N_452);
nor U3485 (N_3485,N_338,N_5);
nand U3486 (N_3486,N_416,N_1698);
and U3487 (N_3487,N_805,N_1453);
nor U3488 (N_3488,N_991,N_914);
xnor U3489 (N_3489,N_106,N_1663);
nor U3490 (N_3490,N_1064,N_1797);
xnor U3491 (N_3491,N_1229,N_1722);
or U3492 (N_3492,N_1538,N_272);
nor U3493 (N_3493,N_753,N_964);
or U3494 (N_3494,N_535,N_791);
nor U3495 (N_3495,N_813,N_379);
nor U3496 (N_3496,N_1531,N_972);
and U3497 (N_3497,N_437,N_1408);
xnor U3498 (N_3498,N_269,N_1122);
xor U3499 (N_3499,N_981,N_402);
and U3500 (N_3500,N_270,N_1971);
or U3501 (N_3501,N_1471,N_476);
and U3502 (N_3502,N_1220,N_578);
and U3503 (N_3503,N_1597,N_851);
nor U3504 (N_3504,N_1990,N_159);
nor U3505 (N_3505,N_6,N_296);
nor U3506 (N_3506,N_343,N_1324);
and U3507 (N_3507,N_1382,N_611);
xor U3508 (N_3508,N_888,N_1343);
xnor U3509 (N_3509,N_1537,N_1731);
xnor U3510 (N_3510,N_1362,N_1970);
or U3511 (N_3511,N_437,N_1460);
nor U3512 (N_3512,N_1679,N_1739);
nor U3513 (N_3513,N_1397,N_1491);
nor U3514 (N_3514,N_83,N_1033);
nor U3515 (N_3515,N_588,N_1814);
nor U3516 (N_3516,N_1236,N_1234);
and U3517 (N_3517,N_616,N_209);
or U3518 (N_3518,N_799,N_104);
and U3519 (N_3519,N_827,N_924);
or U3520 (N_3520,N_1928,N_1418);
and U3521 (N_3521,N_1297,N_1803);
xnor U3522 (N_3522,N_1578,N_1572);
xor U3523 (N_3523,N_9,N_1336);
nor U3524 (N_3524,N_853,N_1155);
nand U3525 (N_3525,N_1877,N_1193);
or U3526 (N_3526,N_442,N_123);
nor U3527 (N_3527,N_1872,N_201);
nand U3528 (N_3528,N_847,N_387);
or U3529 (N_3529,N_398,N_1369);
and U3530 (N_3530,N_151,N_259);
or U3531 (N_3531,N_366,N_1683);
nor U3532 (N_3532,N_1358,N_1555);
nor U3533 (N_3533,N_581,N_1943);
and U3534 (N_3534,N_1913,N_1881);
xnor U3535 (N_3535,N_1949,N_1936);
or U3536 (N_3536,N_1276,N_600);
or U3537 (N_3537,N_619,N_1244);
and U3538 (N_3538,N_1746,N_723);
nand U3539 (N_3539,N_573,N_422);
nor U3540 (N_3540,N_399,N_1781);
or U3541 (N_3541,N_968,N_1940);
and U3542 (N_3542,N_964,N_458);
and U3543 (N_3543,N_1632,N_158);
nor U3544 (N_3544,N_86,N_1891);
or U3545 (N_3545,N_1574,N_1296);
xor U3546 (N_3546,N_542,N_460);
nand U3547 (N_3547,N_523,N_1857);
nand U3548 (N_3548,N_772,N_1578);
xnor U3549 (N_3549,N_1080,N_1842);
nand U3550 (N_3550,N_233,N_1294);
nand U3551 (N_3551,N_1416,N_434);
nor U3552 (N_3552,N_257,N_1840);
xnor U3553 (N_3553,N_1473,N_1998);
or U3554 (N_3554,N_410,N_1916);
and U3555 (N_3555,N_1954,N_231);
and U3556 (N_3556,N_606,N_621);
xor U3557 (N_3557,N_447,N_281);
nand U3558 (N_3558,N_905,N_1122);
or U3559 (N_3559,N_66,N_62);
or U3560 (N_3560,N_1886,N_768);
nand U3561 (N_3561,N_1119,N_1420);
or U3562 (N_3562,N_739,N_1363);
nor U3563 (N_3563,N_208,N_1345);
and U3564 (N_3564,N_653,N_424);
or U3565 (N_3565,N_343,N_1770);
nand U3566 (N_3566,N_1711,N_1433);
and U3567 (N_3567,N_1241,N_1421);
nand U3568 (N_3568,N_1539,N_1870);
xor U3569 (N_3569,N_164,N_951);
nor U3570 (N_3570,N_1787,N_1124);
nand U3571 (N_3571,N_205,N_153);
nor U3572 (N_3572,N_240,N_409);
and U3573 (N_3573,N_84,N_1431);
or U3574 (N_3574,N_972,N_1082);
nor U3575 (N_3575,N_1665,N_942);
and U3576 (N_3576,N_1162,N_1834);
nand U3577 (N_3577,N_292,N_1515);
and U3578 (N_3578,N_1024,N_961);
or U3579 (N_3579,N_1417,N_909);
xor U3580 (N_3580,N_1469,N_288);
nand U3581 (N_3581,N_1107,N_428);
or U3582 (N_3582,N_1377,N_548);
or U3583 (N_3583,N_775,N_1289);
nor U3584 (N_3584,N_1037,N_1709);
nor U3585 (N_3585,N_539,N_628);
nand U3586 (N_3586,N_1811,N_64);
xor U3587 (N_3587,N_1517,N_1258);
nand U3588 (N_3588,N_830,N_1524);
and U3589 (N_3589,N_373,N_1900);
and U3590 (N_3590,N_461,N_1280);
and U3591 (N_3591,N_1924,N_427);
or U3592 (N_3592,N_1755,N_1848);
nand U3593 (N_3593,N_274,N_1827);
and U3594 (N_3594,N_619,N_1125);
nor U3595 (N_3595,N_1761,N_1804);
and U3596 (N_3596,N_10,N_32);
xor U3597 (N_3597,N_1305,N_251);
nor U3598 (N_3598,N_101,N_149);
or U3599 (N_3599,N_508,N_1905);
or U3600 (N_3600,N_418,N_930);
or U3601 (N_3601,N_1364,N_1176);
or U3602 (N_3602,N_1296,N_90);
or U3603 (N_3603,N_1117,N_188);
and U3604 (N_3604,N_1041,N_302);
or U3605 (N_3605,N_1187,N_24);
or U3606 (N_3606,N_626,N_204);
nor U3607 (N_3607,N_264,N_1607);
and U3608 (N_3608,N_543,N_1622);
or U3609 (N_3609,N_344,N_1242);
xnor U3610 (N_3610,N_576,N_705);
nor U3611 (N_3611,N_1271,N_387);
nor U3612 (N_3612,N_1060,N_220);
or U3613 (N_3613,N_1847,N_1305);
xnor U3614 (N_3614,N_1390,N_1553);
nand U3615 (N_3615,N_1609,N_1587);
or U3616 (N_3616,N_871,N_9);
and U3617 (N_3617,N_426,N_1674);
xor U3618 (N_3618,N_58,N_1899);
or U3619 (N_3619,N_560,N_964);
xor U3620 (N_3620,N_157,N_1339);
xor U3621 (N_3621,N_333,N_424);
or U3622 (N_3622,N_1248,N_664);
xor U3623 (N_3623,N_490,N_95);
or U3624 (N_3624,N_173,N_766);
nor U3625 (N_3625,N_436,N_1258);
nand U3626 (N_3626,N_748,N_1368);
or U3627 (N_3627,N_1818,N_118);
xnor U3628 (N_3628,N_650,N_1862);
nor U3629 (N_3629,N_1771,N_15);
and U3630 (N_3630,N_63,N_1020);
nand U3631 (N_3631,N_1076,N_271);
nor U3632 (N_3632,N_1969,N_70);
xor U3633 (N_3633,N_25,N_1593);
and U3634 (N_3634,N_577,N_913);
or U3635 (N_3635,N_720,N_655);
nand U3636 (N_3636,N_1944,N_243);
xor U3637 (N_3637,N_1037,N_168);
nand U3638 (N_3638,N_1644,N_401);
nand U3639 (N_3639,N_354,N_131);
xnor U3640 (N_3640,N_1913,N_1449);
or U3641 (N_3641,N_1698,N_1019);
xor U3642 (N_3642,N_584,N_1295);
or U3643 (N_3643,N_1879,N_1087);
or U3644 (N_3644,N_1564,N_286);
xnor U3645 (N_3645,N_315,N_1290);
xnor U3646 (N_3646,N_1806,N_1718);
nor U3647 (N_3647,N_1309,N_1001);
and U3648 (N_3648,N_478,N_566);
or U3649 (N_3649,N_303,N_353);
nor U3650 (N_3650,N_185,N_377);
or U3651 (N_3651,N_659,N_1567);
and U3652 (N_3652,N_11,N_1844);
xor U3653 (N_3653,N_1833,N_283);
nand U3654 (N_3654,N_220,N_1517);
nor U3655 (N_3655,N_1567,N_1641);
nor U3656 (N_3656,N_1514,N_1959);
nor U3657 (N_3657,N_1921,N_1482);
xor U3658 (N_3658,N_1229,N_1782);
xor U3659 (N_3659,N_328,N_704);
xnor U3660 (N_3660,N_1449,N_1548);
nor U3661 (N_3661,N_999,N_1366);
and U3662 (N_3662,N_246,N_452);
or U3663 (N_3663,N_1261,N_1157);
xnor U3664 (N_3664,N_987,N_865);
nor U3665 (N_3665,N_1796,N_1436);
xnor U3666 (N_3666,N_326,N_334);
xnor U3667 (N_3667,N_1967,N_115);
and U3668 (N_3668,N_1745,N_1660);
or U3669 (N_3669,N_547,N_1139);
nor U3670 (N_3670,N_1916,N_1282);
nand U3671 (N_3671,N_1300,N_1738);
nor U3672 (N_3672,N_312,N_960);
nor U3673 (N_3673,N_620,N_372);
or U3674 (N_3674,N_1966,N_1148);
nand U3675 (N_3675,N_1992,N_1595);
or U3676 (N_3676,N_1605,N_1159);
and U3677 (N_3677,N_640,N_1679);
and U3678 (N_3678,N_1964,N_1340);
and U3679 (N_3679,N_1369,N_1998);
xnor U3680 (N_3680,N_1879,N_631);
nor U3681 (N_3681,N_1160,N_744);
nand U3682 (N_3682,N_562,N_1488);
and U3683 (N_3683,N_210,N_1900);
and U3684 (N_3684,N_302,N_876);
xor U3685 (N_3685,N_1219,N_207);
or U3686 (N_3686,N_474,N_379);
and U3687 (N_3687,N_929,N_1813);
or U3688 (N_3688,N_178,N_428);
or U3689 (N_3689,N_1035,N_1160);
xnor U3690 (N_3690,N_169,N_1412);
nand U3691 (N_3691,N_1274,N_259);
or U3692 (N_3692,N_231,N_912);
or U3693 (N_3693,N_1106,N_1969);
nor U3694 (N_3694,N_1418,N_1832);
nand U3695 (N_3695,N_1214,N_524);
and U3696 (N_3696,N_1177,N_1972);
and U3697 (N_3697,N_1449,N_1815);
and U3698 (N_3698,N_1826,N_1801);
and U3699 (N_3699,N_435,N_950);
or U3700 (N_3700,N_439,N_1133);
or U3701 (N_3701,N_1424,N_917);
nand U3702 (N_3702,N_834,N_1154);
nor U3703 (N_3703,N_737,N_1993);
nand U3704 (N_3704,N_972,N_1322);
nand U3705 (N_3705,N_589,N_240);
and U3706 (N_3706,N_377,N_1418);
nand U3707 (N_3707,N_1356,N_991);
xor U3708 (N_3708,N_1347,N_247);
nand U3709 (N_3709,N_829,N_1286);
and U3710 (N_3710,N_1151,N_472);
xor U3711 (N_3711,N_1514,N_93);
xnor U3712 (N_3712,N_402,N_262);
and U3713 (N_3713,N_1758,N_1565);
or U3714 (N_3714,N_1684,N_1215);
nor U3715 (N_3715,N_1914,N_1677);
or U3716 (N_3716,N_724,N_320);
nor U3717 (N_3717,N_1203,N_371);
nor U3718 (N_3718,N_1277,N_1270);
xnor U3719 (N_3719,N_1160,N_1521);
and U3720 (N_3720,N_597,N_977);
xor U3721 (N_3721,N_1965,N_807);
or U3722 (N_3722,N_1814,N_1522);
xnor U3723 (N_3723,N_1718,N_1364);
and U3724 (N_3724,N_18,N_426);
and U3725 (N_3725,N_120,N_1493);
nand U3726 (N_3726,N_1199,N_848);
xor U3727 (N_3727,N_1352,N_1251);
nand U3728 (N_3728,N_1465,N_241);
and U3729 (N_3729,N_1831,N_1083);
or U3730 (N_3730,N_1847,N_1399);
nand U3731 (N_3731,N_1280,N_1452);
or U3732 (N_3732,N_825,N_1150);
nand U3733 (N_3733,N_1710,N_1093);
nand U3734 (N_3734,N_332,N_1119);
nor U3735 (N_3735,N_36,N_1810);
and U3736 (N_3736,N_1729,N_553);
nor U3737 (N_3737,N_182,N_915);
nor U3738 (N_3738,N_1194,N_1011);
and U3739 (N_3739,N_962,N_1910);
xnor U3740 (N_3740,N_1725,N_1569);
nor U3741 (N_3741,N_1832,N_1381);
nor U3742 (N_3742,N_1176,N_1174);
nor U3743 (N_3743,N_375,N_1081);
nand U3744 (N_3744,N_1807,N_628);
and U3745 (N_3745,N_825,N_143);
nor U3746 (N_3746,N_1039,N_581);
nor U3747 (N_3747,N_1895,N_154);
xnor U3748 (N_3748,N_1884,N_1737);
and U3749 (N_3749,N_1484,N_525);
and U3750 (N_3750,N_1133,N_209);
xor U3751 (N_3751,N_912,N_857);
or U3752 (N_3752,N_1993,N_1202);
or U3753 (N_3753,N_821,N_1163);
or U3754 (N_3754,N_1676,N_799);
or U3755 (N_3755,N_214,N_482);
or U3756 (N_3756,N_998,N_1603);
and U3757 (N_3757,N_1701,N_1595);
and U3758 (N_3758,N_263,N_1137);
nand U3759 (N_3759,N_162,N_193);
nor U3760 (N_3760,N_64,N_1469);
or U3761 (N_3761,N_479,N_182);
nor U3762 (N_3762,N_756,N_1635);
xnor U3763 (N_3763,N_1205,N_584);
or U3764 (N_3764,N_1836,N_1321);
and U3765 (N_3765,N_1257,N_303);
xnor U3766 (N_3766,N_564,N_1037);
nand U3767 (N_3767,N_1171,N_1858);
and U3768 (N_3768,N_988,N_87);
nor U3769 (N_3769,N_1735,N_597);
nand U3770 (N_3770,N_329,N_961);
and U3771 (N_3771,N_1594,N_631);
xnor U3772 (N_3772,N_71,N_192);
nor U3773 (N_3773,N_1343,N_554);
or U3774 (N_3774,N_579,N_1173);
and U3775 (N_3775,N_1116,N_803);
and U3776 (N_3776,N_1185,N_1258);
and U3777 (N_3777,N_92,N_465);
nand U3778 (N_3778,N_733,N_1096);
nand U3779 (N_3779,N_643,N_858);
nor U3780 (N_3780,N_108,N_291);
nor U3781 (N_3781,N_198,N_1597);
nor U3782 (N_3782,N_1499,N_574);
or U3783 (N_3783,N_283,N_1321);
or U3784 (N_3784,N_1934,N_1020);
xnor U3785 (N_3785,N_1811,N_199);
and U3786 (N_3786,N_1555,N_1294);
nand U3787 (N_3787,N_815,N_1181);
and U3788 (N_3788,N_856,N_1256);
nand U3789 (N_3789,N_1031,N_1939);
or U3790 (N_3790,N_892,N_1647);
and U3791 (N_3791,N_766,N_1666);
nor U3792 (N_3792,N_1798,N_667);
xnor U3793 (N_3793,N_35,N_1648);
nand U3794 (N_3794,N_173,N_1164);
nor U3795 (N_3795,N_934,N_244);
nor U3796 (N_3796,N_695,N_1726);
nor U3797 (N_3797,N_476,N_1574);
xnor U3798 (N_3798,N_1356,N_1146);
nand U3799 (N_3799,N_1160,N_1153);
and U3800 (N_3800,N_1453,N_1034);
or U3801 (N_3801,N_1581,N_320);
xor U3802 (N_3802,N_539,N_796);
nor U3803 (N_3803,N_848,N_1804);
xor U3804 (N_3804,N_40,N_1354);
nor U3805 (N_3805,N_1968,N_1052);
or U3806 (N_3806,N_1113,N_97);
nor U3807 (N_3807,N_1667,N_508);
nand U3808 (N_3808,N_1565,N_492);
or U3809 (N_3809,N_1994,N_1864);
nor U3810 (N_3810,N_999,N_313);
nand U3811 (N_3811,N_1341,N_334);
nor U3812 (N_3812,N_1693,N_1142);
and U3813 (N_3813,N_1955,N_1764);
xor U3814 (N_3814,N_819,N_1390);
nor U3815 (N_3815,N_1666,N_1860);
xor U3816 (N_3816,N_1396,N_102);
nor U3817 (N_3817,N_934,N_1038);
or U3818 (N_3818,N_359,N_821);
nor U3819 (N_3819,N_1944,N_1382);
or U3820 (N_3820,N_112,N_40);
nor U3821 (N_3821,N_1536,N_694);
nand U3822 (N_3822,N_1024,N_135);
nand U3823 (N_3823,N_566,N_1820);
and U3824 (N_3824,N_143,N_1539);
nor U3825 (N_3825,N_1627,N_1302);
xor U3826 (N_3826,N_1127,N_1331);
xor U3827 (N_3827,N_1893,N_1789);
nand U3828 (N_3828,N_36,N_1115);
nand U3829 (N_3829,N_131,N_1772);
nor U3830 (N_3830,N_1895,N_202);
xor U3831 (N_3831,N_1212,N_1213);
nand U3832 (N_3832,N_971,N_581);
nand U3833 (N_3833,N_1055,N_1327);
or U3834 (N_3834,N_322,N_685);
nand U3835 (N_3835,N_1349,N_1925);
nor U3836 (N_3836,N_1837,N_1742);
nand U3837 (N_3837,N_191,N_1028);
nand U3838 (N_3838,N_866,N_229);
nor U3839 (N_3839,N_1965,N_1414);
nand U3840 (N_3840,N_410,N_815);
nand U3841 (N_3841,N_1234,N_1532);
nor U3842 (N_3842,N_1146,N_651);
or U3843 (N_3843,N_994,N_446);
nor U3844 (N_3844,N_1103,N_1639);
or U3845 (N_3845,N_903,N_1461);
nor U3846 (N_3846,N_1583,N_555);
or U3847 (N_3847,N_101,N_389);
nor U3848 (N_3848,N_828,N_218);
nand U3849 (N_3849,N_579,N_697);
xor U3850 (N_3850,N_1764,N_1388);
or U3851 (N_3851,N_715,N_1315);
nor U3852 (N_3852,N_1467,N_1610);
and U3853 (N_3853,N_1845,N_469);
or U3854 (N_3854,N_1591,N_1919);
xor U3855 (N_3855,N_727,N_231);
or U3856 (N_3856,N_381,N_907);
or U3857 (N_3857,N_837,N_1338);
nand U3858 (N_3858,N_333,N_1448);
and U3859 (N_3859,N_1787,N_413);
nor U3860 (N_3860,N_849,N_1960);
or U3861 (N_3861,N_964,N_1365);
and U3862 (N_3862,N_1343,N_1771);
nor U3863 (N_3863,N_1684,N_1655);
nor U3864 (N_3864,N_565,N_1292);
xnor U3865 (N_3865,N_442,N_1084);
or U3866 (N_3866,N_1788,N_1588);
and U3867 (N_3867,N_490,N_77);
and U3868 (N_3868,N_1869,N_1926);
nand U3869 (N_3869,N_1339,N_599);
nand U3870 (N_3870,N_1002,N_116);
nor U3871 (N_3871,N_1888,N_615);
nor U3872 (N_3872,N_317,N_1077);
and U3873 (N_3873,N_1190,N_1631);
nand U3874 (N_3874,N_559,N_1849);
nor U3875 (N_3875,N_1609,N_699);
xor U3876 (N_3876,N_978,N_313);
xnor U3877 (N_3877,N_21,N_1121);
and U3878 (N_3878,N_681,N_560);
nand U3879 (N_3879,N_247,N_453);
nand U3880 (N_3880,N_838,N_371);
nor U3881 (N_3881,N_1246,N_1684);
or U3882 (N_3882,N_837,N_336);
or U3883 (N_3883,N_603,N_891);
or U3884 (N_3884,N_273,N_1223);
nor U3885 (N_3885,N_972,N_1820);
or U3886 (N_3886,N_113,N_1420);
xor U3887 (N_3887,N_1988,N_1760);
and U3888 (N_3888,N_457,N_1580);
nand U3889 (N_3889,N_367,N_28);
nor U3890 (N_3890,N_1071,N_571);
and U3891 (N_3891,N_478,N_858);
and U3892 (N_3892,N_951,N_408);
and U3893 (N_3893,N_1732,N_1091);
xor U3894 (N_3894,N_433,N_978);
or U3895 (N_3895,N_1715,N_432);
xnor U3896 (N_3896,N_509,N_436);
and U3897 (N_3897,N_609,N_134);
and U3898 (N_3898,N_853,N_1565);
nor U3899 (N_3899,N_1839,N_1762);
and U3900 (N_3900,N_1267,N_211);
nor U3901 (N_3901,N_1763,N_338);
xnor U3902 (N_3902,N_1594,N_205);
and U3903 (N_3903,N_538,N_1043);
xor U3904 (N_3904,N_947,N_1691);
nand U3905 (N_3905,N_1976,N_66);
nand U3906 (N_3906,N_667,N_1541);
or U3907 (N_3907,N_628,N_576);
nand U3908 (N_3908,N_1719,N_1877);
or U3909 (N_3909,N_1840,N_686);
xor U3910 (N_3910,N_381,N_1801);
or U3911 (N_3911,N_1803,N_1094);
nand U3912 (N_3912,N_350,N_898);
nor U3913 (N_3913,N_1345,N_671);
nor U3914 (N_3914,N_205,N_492);
xor U3915 (N_3915,N_1372,N_171);
xor U3916 (N_3916,N_1426,N_1001);
nor U3917 (N_3917,N_1644,N_1651);
nand U3918 (N_3918,N_425,N_1347);
or U3919 (N_3919,N_381,N_843);
nand U3920 (N_3920,N_565,N_1458);
or U3921 (N_3921,N_954,N_1387);
nor U3922 (N_3922,N_1726,N_604);
or U3923 (N_3923,N_1305,N_52);
xor U3924 (N_3924,N_327,N_900);
xnor U3925 (N_3925,N_1958,N_1295);
xnor U3926 (N_3926,N_994,N_1015);
nand U3927 (N_3927,N_104,N_1189);
nand U3928 (N_3928,N_62,N_823);
and U3929 (N_3929,N_341,N_60);
nor U3930 (N_3930,N_1831,N_1145);
or U3931 (N_3931,N_1458,N_591);
and U3932 (N_3932,N_872,N_1138);
or U3933 (N_3933,N_1335,N_1132);
nor U3934 (N_3934,N_393,N_375);
or U3935 (N_3935,N_239,N_1302);
and U3936 (N_3936,N_1824,N_694);
xnor U3937 (N_3937,N_281,N_1579);
or U3938 (N_3938,N_99,N_1968);
or U3939 (N_3939,N_1919,N_245);
xor U3940 (N_3940,N_1718,N_629);
xnor U3941 (N_3941,N_1606,N_475);
xnor U3942 (N_3942,N_1161,N_1277);
and U3943 (N_3943,N_1586,N_919);
and U3944 (N_3944,N_1025,N_339);
or U3945 (N_3945,N_265,N_1642);
or U3946 (N_3946,N_1775,N_1674);
and U3947 (N_3947,N_371,N_1681);
nand U3948 (N_3948,N_533,N_1112);
and U3949 (N_3949,N_703,N_1467);
or U3950 (N_3950,N_228,N_1964);
nor U3951 (N_3951,N_1733,N_593);
nand U3952 (N_3952,N_1310,N_1505);
nor U3953 (N_3953,N_1265,N_34);
nor U3954 (N_3954,N_1300,N_706);
xnor U3955 (N_3955,N_1427,N_1088);
nor U3956 (N_3956,N_307,N_1614);
nor U3957 (N_3957,N_1160,N_1864);
nand U3958 (N_3958,N_1199,N_1259);
or U3959 (N_3959,N_1603,N_1992);
xnor U3960 (N_3960,N_1372,N_25);
nor U3961 (N_3961,N_992,N_1072);
nand U3962 (N_3962,N_962,N_1735);
xnor U3963 (N_3963,N_208,N_1536);
or U3964 (N_3964,N_1926,N_1410);
or U3965 (N_3965,N_1556,N_1215);
nor U3966 (N_3966,N_454,N_1941);
or U3967 (N_3967,N_1560,N_853);
or U3968 (N_3968,N_1935,N_1110);
nand U3969 (N_3969,N_186,N_408);
or U3970 (N_3970,N_1965,N_1935);
nor U3971 (N_3971,N_542,N_420);
nor U3972 (N_3972,N_1018,N_160);
and U3973 (N_3973,N_975,N_751);
nand U3974 (N_3974,N_477,N_1808);
nor U3975 (N_3975,N_1517,N_1546);
and U3976 (N_3976,N_270,N_535);
or U3977 (N_3977,N_1936,N_1471);
nor U3978 (N_3978,N_1747,N_93);
or U3979 (N_3979,N_1125,N_445);
nand U3980 (N_3980,N_1450,N_260);
nor U3981 (N_3981,N_967,N_1832);
xor U3982 (N_3982,N_880,N_373);
nor U3983 (N_3983,N_772,N_268);
or U3984 (N_3984,N_175,N_406);
or U3985 (N_3985,N_1348,N_1639);
nand U3986 (N_3986,N_1306,N_1388);
and U3987 (N_3987,N_1412,N_990);
xnor U3988 (N_3988,N_1893,N_212);
nand U3989 (N_3989,N_1318,N_108);
and U3990 (N_3990,N_1119,N_1551);
xor U3991 (N_3991,N_1310,N_1687);
or U3992 (N_3992,N_1810,N_873);
nand U3993 (N_3993,N_569,N_110);
or U3994 (N_3994,N_264,N_650);
or U3995 (N_3995,N_404,N_414);
and U3996 (N_3996,N_515,N_453);
xnor U3997 (N_3997,N_644,N_1241);
nand U3998 (N_3998,N_1409,N_993);
xnor U3999 (N_3999,N_1058,N_1124);
or U4000 (N_4000,N_3541,N_3514);
xor U4001 (N_4001,N_2700,N_2507);
nand U4002 (N_4002,N_2305,N_3678);
xor U4003 (N_4003,N_2698,N_3240);
xor U4004 (N_4004,N_2918,N_2039);
or U4005 (N_4005,N_2397,N_3712);
xor U4006 (N_4006,N_2536,N_3256);
xnor U4007 (N_4007,N_2870,N_3647);
or U4008 (N_4008,N_3774,N_3233);
nand U4009 (N_4009,N_2036,N_3727);
or U4010 (N_4010,N_2586,N_2907);
xor U4011 (N_4011,N_3065,N_3892);
or U4012 (N_4012,N_2773,N_2845);
xnor U4013 (N_4013,N_3023,N_2974);
or U4014 (N_4014,N_3329,N_2243);
and U4015 (N_4015,N_2483,N_2994);
nor U4016 (N_4016,N_3166,N_2263);
or U4017 (N_4017,N_3399,N_3562);
or U4018 (N_4018,N_2349,N_2929);
nor U4019 (N_4019,N_3553,N_3605);
xor U4020 (N_4020,N_2205,N_3001);
xnor U4021 (N_4021,N_3397,N_2290);
nor U4022 (N_4022,N_3633,N_2407);
nor U4023 (N_4023,N_2748,N_2682);
nand U4024 (N_4024,N_3851,N_2135);
nor U4025 (N_4025,N_2514,N_3013);
xor U4026 (N_4026,N_3243,N_2401);
nor U4027 (N_4027,N_3050,N_3803);
nor U4028 (N_4028,N_2474,N_2011);
xor U4029 (N_4029,N_2687,N_3281);
or U4030 (N_4030,N_3832,N_2498);
nor U4031 (N_4031,N_2123,N_2463);
or U4032 (N_4032,N_3759,N_3003);
and U4033 (N_4033,N_2440,N_3781);
nor U4034 (N_4034,N_2647,N_2598);
and U4035 (N_4035,N_3254,N_2165);
or U4036 (N_4036,N_2889,N_2551);
or U4037 (N_4037,N_3952,N_2371);
or U4038 (N_4038,N_3807,N_3419);
and U4039 (N_4039,N_2340,N_3905);
nand U4040 (N_4040,N_3915,N_3356);
nor U4041 (N_4041,N_3932,N_3371);
nor U4042 (N_4042,N_2983,N_3015);
and U4043 (N_4043,N_3696,N_3485);
nor U4044 (N_4044,N_2755,N_2074);
xnor U4045 (N_4045,N_2325,N_3768);
and U4046 (N_4046,N_3685,N_2527);
xor U4047 (N_4047,N_2726,N_3101);
xnor U4048 (N_4048,N_3285,N_2570);
nor U4049 (N_4049,N_2057,N_3303);
nor U4050 (N_4050,N_3720,N_2688);
or U4051 (N_4051,N_2099,N_3394);
nand U4052 (N_4052,N_3388,N_3436);
nor U4053 (N_4053,N_3891,N_2991);
xnor U4054 (N_4054,N_3816,N_2424);
or U4055 (N_4055,N_2716,N_2920);
nor U4056 (N_4056,N_3095,N_3366);
nor U4057 (N_4057,N_2620,N_3653);
and U4058 (N_4058,N_3513,N_2078);
or U4059 (N_4059,N_2177,N_3483);
or U4060 (N_4060,N_3568,N_3118);
or U4061 (N_4061,N_3955,N_3214);
nor U4062 (N_4062,N_3462,N_2254);
nand U4063 (N_4063,N_3636,N_2959);
xor U4064 (N_4064,N_3471,N_3822);
or U4065 (N_4065,N_2164,N_3149);
nand U4066 (N_4066,N_2942,N_3081);
or U4067 (N_4067,N_3334,N_3472);
or U4068 (N_4068,N_3398,N_3326);
or U4069 (N_4069,N_3802,N_3474);
or U4070 (N_4070,N_3617,N_2249);
nor U4071 (N_4071,N_2840,N_2893);
or U4072 (N_4072,N_2010,N_3710);
or U4073 (N_4073,N_3817,N_2533);
nand U4074 (N_4074,N_3224,N_3193);
and U4075 (N_4075,N_2579,N_3921);
nand U4076 (N_4076,N_3523,N_2188);
xor U4077 (N_4077,N_3194,N_3931);
nand U4078 (N_4078,N_2418,N_3898);
nand U4079 (N_4079,N_3092,N_3411);
or U4080 (N_4080,N_2382,N_3086);
xnor U4081 (N_4081,N_2098,N_2990);
nor U4082 (N_4082,N_3190,N_3819);
nor U4083 (N_4083,N_2442,N_2226);
and U4084 (N_4084,N_2882,N_3229);
nand U4085 (N_4085,N_2832,N_3967);
nor U4086 (N_4086,N_3631,N_2623);
or U4087 (N_4087,N_2545,N_2992);
or U4088 (N_4088,N_2152,N_3746);
nor U4089 (N_4089,N_2842,N_3940);
or U4090 (N_4090,N_3694,N_2691);
nor U4091 (N_4091,N_3055,N_3794);
nor U4092 (N_4092,N_3219,N_3524);
xnor U4093 (N_4093,N_3521,N_3943);
or U4094 (N_4094,N_2492,N_3908);
nand U4095 (N_4095,N_2095,N_3255);
and U4096 (N_4096,N_2602,N_3151);
nand U4097 (N_4097,N_3742,N_2689);
xor U4098 (N_4098,N_2847,N_2330);
or U4099 (N_4099,N_2635,N_2471);
and U4100 (N_4100,N_3016,N_3335);
nor U4101 (N_4101,N_3903,N_3032);
xnor U4102 (N_4102,N_2791,N_2276);
or U4103 (N_4103,N_3800,N_3043);
nor U4104 (N_4104,N_2601,N_3215);
xor U4105 (N_4105,N_3555,N_2625);
nor U4106 (N_4106,N_3522,N_2841);
xnor U4107 (N_4107,N_3161,N_3295);
nor U4108 (N_4108,N_3619,N_3960);
or U4109 (N_4109,N_2106,N_3992);
nand U4110 (N_4110,N_2192,N_2119);
and U4111 (N_4111,N_2684,N_3236);
and U4112 (N_4112,N_2334,N_2000);
xnor U4113 (N_4113,N_2049,N_2589);
or U4114 (N_4114,N_2599,N_2658);
nor U4115 (N_4115,N_2491,N_2828);
and U4116 (N_4116,N_3845,N_2420);
nand U4117 (N_4117,N_3939,N_2278);
nor U4118 (N_4118,N_2757,N_3038);
or U4119 (N_4119,N_2391,N_3478);
or U4120 (N_4120,N_3597,N_2664);
or U4121 (N_4121,N_2643,N_2131);
nand U4122 (N_4122,N_3789,N_3866);
nor U4123 (N_4123,N_2052,N_3876);
xnor U4124 (N_4124,N_2260,N_2202);
xor U4125 (N_4125,N_3075,N_3705);
or U4126 (N_4126,N_2796,N_3094);
nor U4127 (N_4127,N_2298,N_3646);
nand U4128 (N_4128,N_3682,N_2677);
or U4129 (N_4129,N_2028,N_2128);
and U4130 (N_4130,N_2056,N_3917);
and U4131 (N_4131,N_2680,N_3466);
and U4132 (N_4132,N_3404,N_2523);
xor U4133 (N_4133,N_3582,N_3993);
and U4134 (N_4134,N_2862,N_3676);
and U4135 (N_4135,N_2425,N_2718);
and U4136 (N_4136,N_2332,N_3155);
nand U4137 (N_4137,N_2631,N_2987);
and U4138 (N_4138,N_2692,N_3362);
or U4139 (N_4139,N_3307,N_3990);
nor U4140 (N_4140,N_2110,N_3089);
and U4141 (N_4141,N_2590,N_3687);
and U4142 (N_4142,N_2565,N_2952);
xnor U4143 (N_4143,N_3811,N_3278);
or U4144 (N_4144,N_2734,N_3706);
or U4145 (N_4145,N_3480,N_3137);
and U4146 (N_4146,N_2389,N_2253);
nor U4147 (N_4147,N_3998,N_3359);
and U4148 (N_4148,N_2093,N_2609);
xnor U4149 (N_4149,N_3709,N_3099);
xnor U4150 (N_4150,N_3263,N_3573);
xnor U4151 (N_4151,N_3292,N_2279);
nand U4152 (N_4152,N_3721,N_2663);
and U4153 (N_4153,N_3907,N_3028);
and U4154 (N_4154,N_3925,N_3130);
or U4155 (N_4155,N_2416,N_3987);
nor U4156 (N_4156,N_2070,N_3426);
or U4157 (N_4157,N_3743,N_3077);
nand U4158 (N_4158,N_3838,N_2393);
nand U4159 (N_4159,N_3225,N_3490);
xnor U4160 (N_4160,N_2233,N_3873);
nand U4161 (N_4161,N_2848,N_3324);
xor U4162 (N_4162,N_2676,N_3806);
and U4163 (N_4163,N_3723,N_2489);
and U4164 (N_4164,N_3574,N_2096);
nand U4165 (N_4165,N_2229,N_3121);
or U4166 (N_4166,N_3422,N_2813);
and U4167 (N_4167,N_2013,N_3588);
or U4168 (N_4168,N_2464,N_3639);
nand U4169 (N_4169,N_3184,N_2752);
xnor U4170 (N_4170,N_3280,N_2354);
xnor U4171 (N_4171,N_2733,N_3584);
xnor U4172 (N_4172,N_2512,N_2931);
or U4173 (N_4173,N_3073,N_3569);
xor U4174 (N_4174,N_3748,N_2670);
nand U4175 (N_4175,N_3831,N_2534);
or U4176 (N_4176,N_2854,N_2809);
and U4177 (N_4177,N_3519,N_3577);
nand U4178 (N_4178,N_3464,N_2975);
nor U4179 (N_4179,N_2380,N_3064);
xnor U4180 (N_4180,N_2295,N_3616);
and U4181 (N_4181,N_3009,N_3545);
nand U4182 (N_4182,N_2029,N_3100);
nor U4183 (N_4183,N_2896,N_2517);
nand U4184 (N_4184,N_2657,N_3542);
and U4185 (N_4185,N_2368,N_2493);
xnor U4186 (N_4186,N_2331,N_2034);
xor U4187 (N_4187,N_2549,N_3276);
and U4188 (N_4188,N_2083,N_3056);
nand U4189 (N_4189,N_2428,N_2894);
and U4190 (N_4190,N_2981,N_3841);
nand U4191 (N_4191,N_2802,N_2091);
xnor U4192 (N_4192,N_2877,N_3782);
nor U4193 (N_4193,N_3048,N_3097);
and U4194 (N_4194,N_2208,N_3156);
or U4195 (N_4195,N_3024,N_2482);
and U4196 (N_4196,N_3707,N_3487);
and U4197 (N_4197,N_3864,N_2007);
and U4198 (N_4198,N_3409,N_2210);
nand U4199 (N_4199,N_3714,N_2729);
xor U4200 (N_4200,N_3400,N_2139);
xor U4201 (N_4201,N_3871,N_3423);
or U4202 (N_4202,N_3951,N_3425);
nor U4203 (N_4203,N_3935,N_3637);
nand U4204 (N_4204,N_2741,N_2652);
and U4205 (N_4205,N_3332,N_3237);
or U4206 (N_4206,N_2329,N_3345);
and U4207 (N_4207,N_3516,N_3752);
xnor U4208 (N_4208,N_3235,N_3679);
nor U4209 (N_4209,N_2120,N_2137);
nor U4210 (N_4210,N_3614,N_3405);
or U4211 (N_4211,N_2426,N_2221);
nand U4212 (N_4212,N_3284,N_3327);
nor U4213 (N_4213,N_3942,N_2820);
nor U4214 (N_4214,N_2540,N_2234);
nand U4215 (N_4215,N_2318,N_2417);
nand U4216 (N_4216,N_2793,N_2708);
xor U4217 (N_4217,N_3729,N_2481);
nor U4218 (N_4218,N_3451,N_3188);
nor U4219 (N_4219,N_3078,N_2798);
nor U4220 (N_4220,N_3854,N_2694);
nor U4221 (N_4221,N_3306,N_3842);
and U4222 (N_4222,N_2005,N_2858);
and U4223 (N_4223,N_3860,N_3098);
xnor U4224 (N_4224,N_2693,N_3799);
nor U4225 (N_4225,N_2812,N_3146);
nand U4226 (N_4226,N_3889,N_3596);
and U4227 (N_4227,N_2112,N_2107);
xnor U4228 (N_4228,N_2488,N_3719);
xor U4229 (N_4229,N_2563,N_2525);
xor U4230 (N_4230,N_3196,N_3527);
xnor U4231 (N_4231,N_2582,N_2788);
nand U4232 (N_4232,N_2966,N_2584);
or U4233 (N_4233,N_3595,N_3390);
and U4234 (N_4234,N_2421,N_3493);
nand U4235 (N_4235,N_3543,N_2588);
or U4236 (N_4236,N_2683,N_3063);
nor U4237 (N_4237,N_2486,N_2556);
nor U4238 (N_4238,N_3642,N_3693);
xnor U4239 (N_4239,N_2129,N_3695);
and U4240 (N_4240,N_2115,N_2903);
nor U4241 (N_4241,N_3823,N_2315);
nor U4242 (N_4242,N_3777,N_3771);
xnor U4243 (N_4243,N_2374,N_3894);
and U4244 (N_4244,N_2508,N_3176);
nand U4245 (N_4245,N_2504,N_3269);
or U4246 (N_4246,N_3628,N_2906);
or U4247 (N_4247,N_3966,N_3997);
nor U4248 (N_4248,N_2972,N_3000);
nand U4249 (N_4249,N_3376,N_3883);
nand U4250 (N_4250,N_2134,N_3242);
or U4251 (N_4251,N_3593,N_2580);
or U4252 (N_4252,N_3826,N_3949);
nand U4253 (N_4253,N_3780,N_3648);
xor U4254 (N_4254,N_2344,N_3395);
nor U4255 (N_4255,N_2366,N_3208);
nor U4256 (N_4256,N_3618,N_2785);
and U4257 (N_4257,N_2406,N_2963);
and U4258 (N_4258,N_3052,N_2561);
or U4259 (N_4259,N_3266,N_2101);
or U4260 (N_4260,N_2160,N_2247);
or U4261 (N_4261,N_2776,N_2568);
nor U4262 (N_4262,N_3191,N_2833);
nand U4263 (N_4263,N_3333,N_3624);
or U4264 (N_4264,N_3994,N_3981);
or U4265 (N_4265,N_2255,N_2228);
nor U4266 (N_4266,N_2238,N_3034);
or U4267 (N_4267,N_3289,N_3258);
nand U4268 (N_4268,N_2869,N_2242);
nand U4269 (N_4269,N_3890,N_2521);
and U4270 (N_4270,N_2660,N_2470);
and U4271 (N_4271,N_3260,N_3491);
xor U4272 (N_4272,N_2714,N_2654);
and U4273 (N_4273,N_3173,N_2302);
nand U4274 (N_4274,N_3297,N_3933);
and U4275 (N_4275,N_3186,N_2182);
or U4276 (N_4276,N_3415,N_3004);
xnor U4277 (N_4277,N_3205,N_2412);
xnor U4278 (N_4278,N_2913,N_3899);
xnor U4279 (N_4279,N_3231,N_2600);
nor U4280 (N_4280,N_3878,N_2023);
nand U4281 (N_4281,N_3259,N_2411);
or U4282 (N_4282,N_3911,N_3136);
and U4283 (N_4283,N_3557,N_2665);
xnor U4284 (N_4284,N_2114,N_2460);
or U4285 (N_4285,N_2312,N_2581);
and U4286 (N_4286,N_2447,N_2308);
nand U4287 (N_4287,N_3470,N_2054);
xnor U4288 (N_4288,N_2853,N_2985);
nand U4289 (N_4289,N_3182,N_3717);
xor U4290 (N_4290,N_2476,N_3054);
nor U4291 (N_4291,N_3529,N_2433);
or U4292 (N_4292,N_3393,N_3020);
nand U4293 (N_4293,N_3066,N_2430);
nor U4294 (N_4294,N_3670,N_2267);
nor U4295 (N_4295,N_3758,N_3881);
and U4296 (N_4296,N_3677,N_2899);
nor U4297 (N_4297,N_2431,N_3251);
nor U4298 (N_4298,N_3927,N_2797);
nor U4299 (N_4299,N_3872,N_3575);
nand U4300 (N_4300,N_2436,N_2458);
or U4301 (N_4301,N_3314,N_3041);
nand U4302 (N_4302,N_3657,N_3414);
and U4303 (N_4303,N_2587,N_2520);
nor U4304 (N_4304,N_2980,N_2209);
or U4305 (N_4305,N_2022,N_2358);
nor U4306 (N_4306,N_3510,N_3726);
nor U4307 (N_4307,N_3632,N_2863);
nor U4308 (N_4308,N_3133,N_2457);
and U4309 (N_4309,N_3681,N_2145);
nor U4310 (N_4310,N_2956,N_2954);
xnor U4311 (N_4311,N_2810,N_3152);
xor U4312 (N_4312,N_2958,N_2178);
or U4313 (N_4313,N_2880,N_2567);
nand U4314 (N_4314,N_2050,N_2136);
nand U4315 (N_4315,N_3974,N_3621);
nand U4316 (N_4316,N_2257,N_2180);
nand U4317 (N_4317,N_3120,N_2181);
or U4318 (N_4318,N_2675,N_2284);
xor U4319 (N_4319,N_3587,N_2686);
xor U4320 (N_4320,N_2744,N_2821);
or U4321 (N_4321,N_2021,N_2914);
and U4322 (N_4322,N_3355,N_3879);
nor U4323 (N_4323,N_2807,N_3068);
nand U4324 (N_4324,N_2085,N_2794);
nand U4325 (N_4325,N_2876,N_3548);
nand U4326 (N_4326,N_3975,N_3641);
or U4327 (N_4327,N_3740,N_2736);
nor U4328 (N_4328,N_3164,N_3241);
xor U4329 (N_4329,N_2968,N_2575);
xnor U4330 (N_4330,N_3459,N_3906);
or U4331 (N_4331,N_2891,N_2189);
and U4332 (N_4332,N_2272,N_3420);
nor U4333 (N_4333,N_2113,N_2452);
and U4334 (N_4334,N_2496,N_3924);
nor U4335 (N_4335,N_3517,N_2065);
xor U4336 (N_4336,N_2775,N_2381);
or U4337 (N_4337,N_2611,N_3358);
xor U4338 (N_4338,N_3686,N_3223);
xnor U4339 (N_4339,N_3107,N_3724);
nand U4340 (N_4340,N_3311,N_3102);
or U4341 (N_4341,N_3279,N_3572);
xor U4342 (N_4342,N_2289,N_3535);
or U4343 (N_4343,N_2341,N_2976);
and U4344 (N_4344,N_3812,N_3814);
or U4345 (N_4345,N_2232,N_2634);
and U4346 (N_4346,N_2058,N_2090);
and U4347 (N_4347,N_2740,N_2307);
or U4348 (N_4348,N_2199,N_2695);
nand U4349 (N_4349,N_3827,N_3318);
and U4350 (N_4350,N_2337,N_3167);
or U4351 (N_4351,N_3185,N_3886);
and U4352 (N_4352,N_3112,N_3505);
xnor U4353 (N_4353,N_2617,N_3021);
nand U4354 (N_4354,N_3407,N_2604);
nand U4355 (N_4355,N_2443,N_2500);
and U4356 (N_4356,N_3689,N_2328);
nor U4357 (N_4357,N_2583,N_2917);
or U4358 (N_4358,N_3045,N_2273);
nand U4359 (N_4359,N_3109,N_2150);
and U4360 (N_4360,N_2200,N_3901);
nand U4361 (N_4361,N_3058,N_2978);
and U4362 (N_4362,N_2535,N_3843);
xnor U4363 (N_4363,N_3210,N_2553);
and U4364 (N_4364,N_2361,N_2047);
xnor U4365 (N_4365,N_2154,N_3716);
xor U4366 (N_4366,N_3923,N_2701);
and U4367 (N_4367,N_2495,N_3382);
nor U4368 (N_4368,N_3357,N_3808);
nand U4369 (N_4369,N_3127,N_3410);
xnor U4370 (N_4370,N_2747,N_2395);
xor U4371 (N_4371,N_2613,N_3790);
nor U4372 (N_4372,N_2211,N_2649);
nand U4373 (N_4373,N_3005,N_3928);
and U4374 (N_4374,N_3732,N_2979);
or U4375 (N_4375,N_3668,N_3062);
or U4376 (N_4376,N_3140,N_2014);
nor U4377 (N_4377,N_2759,N_2127);
xnor U4378 (N_4378,N_2105,N_3507);
nor U4379 (N_4379,N_3406,N_3738);
xnor U4380 (N_4380,N_2711,N_2285);
or U4381 (N_4381,N_3262,N_2288);
nand U4382 (N_4382,N_2944,N_2518);
and U4383 (N_4383,N_3046,N_3948);
nor U4384 (N_4384,N_3785,N_3837);
or U4385 (N_4385,N_2002,N_2666);
nand U4386 (N_4386,N_3500,N_2133);
xor U4387 (N_4387,N_3551,N_2097);
xnor U4388 (N_4388,N_2286,N_2887);
and U4389 (N_4389,N_3010,N_2051);
xnor U4390 (N_4390,N_3435,N_3481);
nand U4391 (N_4391,N_2179,N_2450);
nor U4392 (N_4392,N_3143,N_3914);
nor U4393 (N_4393,N_3468,N_3683);
nand U4394 (N_4394,N_2453,N_2789);
nand U4395 (N_4395,N_2819,N_2277);
xor U4396 (N_4396,N_2597,N_3565);
or U4397 (N_4397,N_2161,N_3469);
xor U4398 (N_4398,N_3135,N_3502);
nor U4399 (N_4399,N_3116,N_2557);
xor U4400 (N_4400,N_3867,N_3440);
and U4401 (N_4401,N_3042,N_2859);
xnor U4402 (N_4402,N_2373,N_3110);
xnor U4403 (N_4403,N_2068,N_3764);
and U4404 (N_4404,N_2938,N_2851);
and U4405 (N_4405,N_2158,N_2902);
or U4406 (N_4406,N_2445,N_3762);
nor U4407 (N_4407,N_3498,N_2792);
nand U4408 (N_4408,N_3609,N_2356);
xor U4409 (N_4409,N_2313,N_2142);
and U4410 (N_4410,N_3037,N_2259);
xor U4411 (N_4411,N_3375,N_2048);
xnor U4412 (N_4412,N_3373,N_3141);
nand U4413 (N_4413,N_2351,N_3700);
xor U4414 (N_4414,N_3608,N_3713);
nor U4415 (N_4415,N_2388,N_2915);
and U4416 (N_4416,N_2219,N_3044);
nand U4417 (N_4417,N_2637,N_2001);
nor U4418 (N_4418,N_3880,N_2075);
or U4419 (N_4419,N_3014,N_3699);
nor U4420 (N_4420,N_2564,N_3634);
xnor U4421 (N_4421,N_3735,N_3512);
and U4422 (N_4422,N_3850,N_3348);
and U4423 (N_4423,N_3217,N_2619);
or U4424 (N_4424,N_2799,N_3627);
or U4425 (N_4425,N_3200,N_3970);
nor U4426 (N_4426,N_3783,N_3980);
nor U4427 (N_4427,N_2172,N_2645);
nand U4428 (N_4428,N_3766,N_3652);
and U4429 (N_4429,N_2861,N_3600);
or U4430 (N_4430,N_3660,N_2541);
xor U4431 (N_4431,N_2667,N_2860);
and U4432 (N_4432,N_3773,N_2248);
or U4433 (N_4433,N_3858,N_2246);
or U4434 (N_4434,N_2003,N_3560);
or U4435 (N_4435,N_3283,N_2025);
nand U4436 (N_4436,N_3603,N_3111);
and U4437 (N_4437,N_2310,N_3501);
nand U4438 (N_4438,N_3650,N_2008);
nor U4439 (N_4439,N_3069,N_3341);
nand U4440 (N_4440,N_3739,N_2364);
xnor U4441 (N_4441,N_3995,N_3315);
and U4442 (N_4442,N_2932,N_2758);
nor U4443 (N_4443,N_3760,N_3602);
nor U4444 (N_4444,N_3012,N_3887);
and U4445 (N_4445,N_3477,N_2222);
and U4446 (N_4446,N_2753,N_3961);
nor U4447 (N_4447,N_2865,N_3438);
nor U4448 (N_4448,N_2546,N_2745);
and U4449 (N_4449,N_3989,N_2900);
or U4450 (N_4450,N_2293,N_3197);
nand U4451 (N_4451,N_3590,N_2301);
or U4452 (N_4452,N_3863,N_2988);
xor U4453 (N_4453,N_3476,N_3294);
nor U4454 (N_4454,N_2360,N_3549);
or U4455 (N_4455,N_2618,N_2555);
nand U4456 (N_4456,N_2960,N_2890);
xnor U4457 (N_4457,N_2641,N_3325);
xor U4458 (N_4458,N_2703,N_2326);
or U4459 (N_4459,N_3368,N_2270);
and U4460 (N_4460,N_3996,N_2731);
and U4461 (N_4461,N_2348,N_2621);
and U4462 (N_4462,N_3869,N_3484);
nor U4463 (N_4463,N_2678,N_3479);
or U4464 (N_4464,N_2245,N_2530);
nand U4465 (N_4465,N_2685,N_3797);
xor U4466 (N_4466,N_2299,N_3122);
and U4467 (N_4467,N_2998,N_2814);
or U4468 (N_4468,N_2218,N_3308);
nand U4469 (N_4469,N_2239,N_2214);
and U4470 (N_4470,N_3142,N_3396);
or U4471 (N_4471,N_3968,N_2092);
xnor U4472 (N_4472,N_2478,N_2919);
or U4473 (N_4473,N_2343,N_3369);
xnor U4474 (N_4474,N_3450,N_2359);
or U4475 (N_4475,N_3401,N_2943);
nor U4476 (N_4476,N_2501,N_2184);
or U4477 (N_4477,N_2696,N_3265);
nor U4478 (N_4478,N_3339,N_2079);
and U4479 (N_4479,N_3463,N_3443);
or U4480 (N_4480,N_3319,N_2937);
or U4481 (N_4481,N_2642,N_2472);
and U4482 (N_4482,N_2262,N_3029);
nand U4483 (N_4483,N_3868,N_3002);
or U4484 (N_4484,N_3536,N_2559);
and U4485 (N_4485,N_2399,N_2477);
nand U4486 (N_4486,N_2271,N_2429);
nor U4487 (N_4487,N_2964,N_2143);
and U4488 (N_4488,N_2282,N_3730);
nor U4489 (N_4489,N_3673,N_2834);
or U4490 (N_4490,N_3026,N_2309);
nor U4491 (N_4491,N_2439,N_3962);
nor U4492 (N_4492,N_3778,N_2511);
nand U4493 (N_4493,N_2283,N_3828);
nor U4494 (N_4494,N_3839,N_2949);
xnor U4495 (N_4495,N_3147,N_3449);
nor U4496 (N_4496,N_2251,N_2043);
and U4497 (N_4497,N_2197,N_2017);
and U4498 (N_4498,N_3216,N_2846);
or U4499 (N_4499,N_3033,N_2080);
nor U4500 (N_4500,N_2355,N_3277);
or U4501 (N_4501,N_3145,N_3718);
nand U4502 (N_4502,N_2206,N_2707);
nand U4503 (N_4503,N_3900,N_2543);
nand U4504 (N_4504,N_2198,N_3862);
nor U4505 (N_4505,N_3926,N_3930);
nor U4506 (N_4506,N_2215,N_3787);
xnor U4507 (N_4507,N_3007,N_3011);
nor U4508 (N_4508,N_2319,N_3374);
nor U4509 (N_4509,N_2275,N_3909);
and U4510 (N_4510,N_2414,N_3546);
or U4511 (N_4511,N_3818,N_3589);
xor U4512 (N_4512,N_3991,N_2930);
nand U4513 (N_4513,N_2350,N_2713);
xor U4514 (N_4514,N_2438,N_2372);
and U4515 (N_4515,N_3257,N_2592);
xor U4516 (N_4516,N_2103,N_2207);
nor U4517 (N_4517,N_3986,N_2662);
nor U4518 (N_4518,N_3902,N_2661);
nor U4519 (N_4519,N_3747,N_2339);
and U4520 (N_4520,N_2385,N_3076);
or U4521 (N_4521,N_3520,N_2422);
nor U4522 (N_4522,N_2503,N_3458);
nand U4523 (N_4523,N_2912,N_2940);
nor U4524 (N_4524,N_2055,N_2909);
nand U4525 (N_4525,N_2435,N_3203);
xnor U4526 (N_4526,N_3113,N_3690);
nor U4527 (N_4527,N_2852,N_2626);
xor U4528 (N_4528,N_2697,N_2322);
nand U4529 (N_4529,N_2737,N_3040);
nor U4530 (N_4530,N_3667,N_3936);
nor U4531 (N_4531,N_2973,N_3206);
or U4532 (N_4532,N_2327,N_2281);
nor U4533 (N_4533,N_3228,N_2951);
nor U4534 (N_4534,N_2323,N_3175);
xnor U4535 (N_4535,N_3623,N_3731);
nand U4536 (N_4536,N_3865,N_3979);
nor U4537 (N_4537,N_2856,N_2108);
or U4538 (N_4538,N_3434,N_3352);
xnor U4539 (N_4539,N_2462,N_2779);
xnor U4540 (N_4540,N_2466,N_2314);
xnor U4541 (N_4541,N_2668,N_3134);
xor U4542 (N_4542,N_3170,N_2223);
and U4543 (N_4543,N_2138,N_2513);
and U4544 (N_4544,N_3377,N_3183);
xnor U4545 (N_4545,N_3736,N_2924);
and U4546 (N_4546,N_3402,N_2591);
xor U4547 (N_4547,N_3439,N_3104);
nand U4548 (N_4548,N_3763,N_2871);
nand U4549 (N_4549,N_3855,N_2392);
and U4550 (N_4550,N_2303,N_2378);
nor U4551 (N_4551,N_2720,N_2724);
nor U4552 (N_4552,N_3030,N_3558);
nor U4553 (N_4553,N_2224,N_2061);
nor U4554 (N_4554,N_2063,N_2574);
and U4555 (N_4555,N_2370,N_3131);
xnor U4556 (N_4556,N_2191,N_2256);
and U4557 (N_4557,N_2027,N_3181);
and U4558 (N_4558,N_2780,N_2644);
nor U4559 (N_4559,N_3749,N_2089);
nor U4560 (N_4560,N_3846,N_3432);
or U4561 (N_4561,N_3360,N_2892);
nand U4562 (N_4562,N_3538,N_2633);
or U4563 (N_4563,N_2086,N_3775);
xnor U4564 (N_4564,N_2404,N_3159);
xnor U4565 (N_4565,N_3629,N_3074);
nor U4566 (N_4566,N_3218,N_3761);
xor U4567 (N_4567,N_3059,N_2151);
nand U4568 (N_4568,N_2539,N_3753);
nor U4569 (N_4569,N_3129,N_3656);
or U4570 (N_4570,N_2529,N_3692);
and U4571 (N_4571,N_2155,N_2965);
and U4572 (N_4572,N_3204,N_2171);
and U4573 (N_4573,N_2811,N_2550);
nand U4574 (N_4574,N_3496,N_2212);
xor U4575 (N_4575,N_2526,N_3017);
or U4576 (N_4576,N_3082,N_2725);
xor U4577 (N_4577,N_2910,N_3503);
xor U4578 (N_4578,N_2795,N_3684);
nor U4579 (N_4579,N_2185,N_2578);
or U4580 (N_4580,N_2084,N_2577);
xnor U4581 (N_4581,N_2157,N_3722);
nand U4582 (N_4582,N_3654,N_3896);
nand U4583 (N_4583,N_2274,N_3953);
xnor U4584 (N_4584,N_2190,N_3247);
xnor U4585 (N_4585,N_2317,N_3934);
and U4586 (N_4586,N_3221,N_2220);
nor U4587 (N_4587,N_2444,N_2719);
xnor U4588 (N_4588,N_3830,N_3389);
nand U4589 (N_4589,N_2593,N_2554);
nor U4590 (N_4590,N_2419,N_2552);
and U4591 (N_4591,N_2532,N_3630);
or U4592 (N_4592,N_3313,N_2933);
and U4593 (N_4593,N_2427,N_2805);
or U4594 (N_4594,N_2606,N_2163);
nor U4595 (N_4595,N_2367,N_2032);
or U4596 (N_4596,N_3250,N_3337);
nand U4597 (N_4597,N_2494,N_3189);
or U4598 (N_4598,N_3751,N_3620);
or U4599 (N_4599,N_3475,N_2244);
or U4600 (N_4600,N_3604,N_3665);
nand U4601 (N_4601,N_3586,N_2046);
xor U4602 (N_4602,N_2706,N_2300);
xnor U4603 (N_4603,N_2204,N_2766);
and U4604 (N_4604,N_2144,N_2572);
and U4605 (N_4605,N_3408,N_2769);
nand U4606 (N_4606,N_3364,N_3019);
xnor U4607 (N_4607,N_2672,N_2786);
and U4608 (N_4608,N_2149,N_2895);
nor U4609 (N_4609,N_3252,N_3322);
nor U4610 (N_4610,N_3946,N_3912);
xor U4611 (N_4611,N_2291,N_3361);
nor U4612 (N_4612,N_2800,N_3504);
xor U4613 (N_4613,N_2148,N_2566);
nand U4614 (N_4614,N_2159,N_3022);
nand U4615 (N_4615,N_3126,N_3655);
nand U4616 (N_4616,N_2732,N_3821);
or U4617 (N_4617,N_2738,N_3305);
and U4618 (N_4618,N_3103,N_2240);
nand U4619 (N_4619,N_3072,N_2961);
nor U4620 (N_4620,N_3622,N_2772);
nand U4621 (N_4621,N_2921,N_2018);
xor U4622 (N_4622,N_2727,N_3465);
or U4623 (N_4623,N_2916,N_3080);
and U4624 (N_4624,N_2957,N_2225);
nor U4625 (N_4625,N_3160,N_2363);
and U4626 (N_4626,N_2573,N_2037);
nand U4627 (N_4627,N_3611,N_2742);
nor U4628 (N_4628,N_2615,N_3836);
nor U4629 (N_4629,N_3416,N_3564);
nor U4630 (N_4630,N_3246,N_2522);
or U4631 (N_4631,N_2826,N_2237);
and U4632 (N_4632,N_2808,N_3421);
nand U4633 (N_4633,N_2926,N_3226);
or U4634 (N_4634,N_2019,N_3202);
nor U4635 (N_4635,N_2156,N_3972);
nor U4636 (N_4636,N_3988,N_3640);
or U4637 (N_4637,N_2879,N_3290);
and U4638 (N_4638,N_2400,N_3963);
nand U4639 (N_4639,N_2982,N_3317);
and U4640 (N_4640,N_3825,N_3916);
nand U4641 (N_4641,N_3805,N_3492);
nor U4642 (N_4642,N_3286,N_3645);
nand U4643 (N_4643,N_2883,N_2857);
nand U4644 (N_4644,N_2352,N_3249);
and U4645 (N_4645,N_3253,N_3509);
nand U4646 (N_4646,N_3370,N_2170);
and U4647 (N_4647,N_3494,N_2855);
and U4648 (N_4648,N_2100,N_3537);
and U4649 (N_4649,N_3239,N_3563);
or U4650 (N_4650,N_3282,N_2030);
and U4651 (N_4651,N_3708,N_2415);
nand U4652 (N_4652,N_2763,N_2124);
or U4653 (N_4653,N_3340,N_2996);
nand U4654 (N_4654,N_2451,N_3659);
or U4655 (N_4655,N_2297,N_3025);
nand U4656 (N_4656,N_3456,N_3671);
nand U4657 (N_4657,N_2867,N_2515);
nor U4658 (N_4658,N_2632,N_2006);
nand U4659 (N_4659,N_2213,N_3162);
xor U4660 (N_4660,N_3312,N_2947);
nor U4661 (N_4661,N_2073,N_3299);
and U4662 (N_4662,N_2434,N_2296);
nor U4663 (N_4663,N_2898,N_3444);
nand U4664 (N_4664,N_3351,N_3750);
nor U4665 (N_4665,N_3061,N_2454);
nor U4666 (N_4666,N_2506,N_2835);
nand U4667 (N_4667,N_3661,N_2768);
or U4668 (N_4668,N_3944,N_3461);
xor U4669 (N_4669,N_2946,N_2102);
nor U4670 (N_4670,N_2749,N_3499);
nand U4671 (N_4671,N_2628,N_3093);
nor U4672 (N_4672,N_2624,N_2817);
nor U4673 (N_4673,N_3567,N_2967);
and U4674 (N_4674,N_3929,N_2760);
xor U4675 (N_4675,N_2699,N_3446);
and U4676 (N_4676,N_3848,N_3154);
nor U4677 (N_4677,N_3945,N_3353);
xor U4678 (N_4678,N_2831,N_3195);
and U4679 (N_4679,N_2258,N_3384);
nand U4680 (N_4680,N_3663,N_3035);
or U4681 (N_4681,N_2995,N_3383);
or U4682 (N_4682,N_3888,N_3937);
and U4683 (N_4683,N_2923,N_2839);
nand U4684 (N_4684,N_2955,N_2196);
and U4685 (N_4685,N_2292,N_2402);
xnor U4686 (N_4686,N_2636,N_2803);
nor U4687 (N_4687,N_3877,N_3316);
nand U4688 (N_4688,N_3091,N_2362);
xnor U4689 (N_4689,N_2041,N_3267);
nor U4690 (N_4690,N_2674,N_3884);
and U4691 (N_4691,N_3380,N_2648);
or U4692 (N_4692,N_3338,N_2690);
nor U4693 (N_4693,N_3445,N_3583);
or U4694 (N_4694,N_2962,N_2784);
nand U4695 (N_4695,N_2169,N_2544);
and U4696 (N_4696,N_3559,N_2026);
xor U4697 (N_4697,N_2971,N_2825);
nand U4698 (N_4698,N_2774,N_2423);
or U4699 (N_4699,N_2268,N_2409);
xor U4700 (N_4700,N_2767,N_2465);
nand U4701 (N_4701,N_2217,N_3801);
xor U4702 (N_4702,N_3870,N_2531);
or U4703 (N_4703,N_2781,N_3482);
nor U4704 (N_4704,N_3320,N_2905);
or U4705 (N_4705,N_2864,N_2984);
xnor U4706 (N_4706,N_2754,N_3447);
xnor U4707 (N_4707,N_3298,N_3448);
and U4708 (N_4708,N_3978,N_2376);
xor U4709 (N_4709,N_3741,N_3756);
nand U4710 (N_4710,N_3209,N_3964);
and U4711 (N_4711,N_2712,N_2448);
nor U4712 (N_4712,N_3638,N_3528);
or U4713 (N_4713,N_2071,N_3244);
nor U4714 (N_4714,N_3117,N_2173);
xor U4715 (N_4715,N_3983,N_2771);
or U4716 (N_4716,N_3403,N_3232);
nor U4717 (N_4717,N_2266,N_2175);
xor U4718 (N_4718,N_3526,N_3168);
and U4719 (N_4719,N_2778,N_3779);
and U4720 (N_4720,N_2822,N_3392);
xor U4721 (N_4721,N_2235,N_3417);
nor U4722 (N_4722,N_3347,N_2432);
or U4723 (N_4723,N_2261,N_3053);
and U4724 (N_4724,N_2783,N_2928);
or U4725 (N_4725,N_3153,N_2596);
and U4726 (N_4726,N_2576,N_3495);
xor U4727 (N_4727,N_2394,N_2403);
and U4728 (N_4728,N_2655,N_3165);
xnor U4729 (N_4729,N_3457,N_2230);
nor U4730 (N_4730,N_2387,N_2241);
xor U4731 (N_4731,N_2316,N_3755);
nor U4732 (N_4732,N_3651,N_3594);
nand U4733 (N_4733,N_2999,N_2186);
xor U4734 (N_4734,N_2622,N_3174);
nor U4735 (N_4735,N_2723,N_3211);
or U4736 (N_4736,N_2751,N_3087);
xor U4737 (N_4737,N_2524,N_3767);
nand U4738 (N_4738,N_2390,N_2117);
xnor U4739 (N_4739,N_3544,N_2610);
nor U4740 (N_4740,N_3088,N_3179);
xnor U4741 (N_4741,N_2195,N_2761);
or U4742 (N_4742,N_2336,N_3006);
xnor U4743 (N_4743,N_3342,N_3772);
xor U4744 (N_4744,N_3302,N_2950);
and U4745 (N_4745,N_3804,N_2743);
xor U4746 (N_4746,N_3123,N_3346);
xnor U4747 (N_4747,N_2801,N_2176);
or U4748 (N_4748,N_2849,N_3139);
xor U4749 (N_4749,N_2116,N_3835);
xnor U4750 (N_4750,N_3171,N_2558);
and U4751 (N_4751,N_2837,N_3920);
and U4752 (N_4752,N_2346,N_2044);
and U4753 (N_4753,N_2094,N_2059);
or U4754 (N_4754,N_2236,N_2320);
nor U4755 (N_4755,N_3387,N_3157);
xnor U4756 (N_4756,N_3856,N_3591);
nor U4757 (N_4757,N_2009,N_2053);
and U4758 (N_4758,N_2509,N_3534);
and U4759 (N_4759,N_2252,N_2970);
nor U4760 (N_4760,N_3442,N_2646);
xor U4761 (N_4761,N_3031,N_2111);
nand U4762 (N_4762,N_3809,N_3672);
nor U4763 (N_4763,N_2201,N_2874);
or U4764 (N_4764,N_2829,N_3177);
nor U4765 (N_4765,N_3350,N_2756);
nand U4766 (N_4766,N_2455,N_2823);
nand U4767 (N_4767,N_3275,N_3938);
xor U4768 (N_4768,N_2715,N_2384);
and U4769 (N_4769,N_3234,N_2265);
xnor U4770 (N_4770,N_2872,N_3288);
xnor U4771 (N_4771,N_3083,N_2174);
nor U4772 (N_4772,N_2901,N_2827);
nor U4773 (N_4773,N_3734,N_3893);
and U4774 (N_4774,N_2125,N_2904);
nand U4775 (N_4775,N_2866,N_2945);
nor U4776 (N_4776,N_3085,N_2659);
nand U4777 (N_4777,N_2925,N_2410);
or U4778 (N_4778,N_3379,N_2977);
and U4779 (N_4779,N_2722,N_2499);
nand U4780 (N_4780,N_2562,N_2850);
xnor U4781 (N_4781,N_3950,N_2306);
and U4782 (N_4782,N_3429,N_2088);
and U4783 (N_4783,N_3580,N_3859);
or U4784 (N_4784,N_3506,N_2510);
nor U4785 (N_4785,N_2437,N_3737);
and U4786 (N_4786,N_3310,N_3515);
and U4787 (N_4787,N_3261,N_3518);
xnor U4788 (N_4788,N_3343,N_2782);
nand U4789 (N_4789,N_3982,N_2612);
or U4790 (N_4790,N_3844,N_3222);
nand U4791 (N_4791,N_2485,N_2519);
and U4792 (N_4792,N_3829,N_3984);
xor U4793 (N_4793,N_2269,N_3273);
xor U4794 (N_4794,N_2024,N_2167);
or U4795 (N_4795,N_3212,N_2630);
nor U4796 (N_4796,N_3853,N_3454);
or U4797 (N_4797,N_3119,N_2603);
xor U4798 (N_4798,N_2548,N_2639);
nand U4799 (N_4799,N_3128,N_3124);
nor U4800 (N_4800,N_3776,N_3291);
and U4801 (N_4801,N_2653,N_2168);
or U4802 (N_4802,N_3106,N_2656);
nand U4803 (N_4803,N_2804,N_2087);
or U4804 (N_4804,N_2594,N_3264);
xor U4805 (N_4805,N_2383,N_3550);
or U4806 (N_4806,N_2516,N_2939);
xnor U4807 (N_4807,N_2750,N_3245);
and U4808 (N_4808,N_3786,N_3386);
nor U4809 (N_4809,N_2673,N_3815);
and U4810 (N_4810,N_3144,N_2042);
xnor U4811 (N_4811,N_3453,N_3354);
and U4812 (N_4812,N_3561,N_2077);
xor U4813 (N_4813,N_2730,N_3757);
xor U4814 (N_4814,N_3079,N_2398);
xor U4815 (N_4815,N_3798,N_2250);
xnor U4816 (N_4816,N_3592,N_3508);
or U4817 (N_4817,N_2989,N_3947);
xnor U4818 (N_4818,N_2475,N_3715);
xor U4819 (N_4819,N_2335,N_2941);
xnor U4820 (N_4820,N_3918,N_3178);
nor U4821 (N_4821,N_2986,N_2396);
or U4822 (N_4822,N_3304,N_3649);
nand U4823 (N_4823,N_3680,N_3702);
nand U4824 (N_4824,N_3150,N_2338);
xor U4825 (N_4825,N_3270,N_2911);
and U4826 (N_4826,N_3703,N_3138);
xor U4827 (N_4827,N_2405,N_2838);
nor U4828 (N_4828,N_3977,N_3180);
and U4829 (N_4829,N_3441,N_3552);
nand U4830 (N_4830,N_2836,N_2936);
nand U4831 (N_4831,N_3788,N_3585);
nand U4832 (N_4832,N_2770,N_2746);
and U4833 (N_4833,N_3688,N_3857);
or U4834 (N_4834,N_3607,N_2638);
xor U4835 (N_4835,N_2365,N_3669);
nand U4836 (N_4836,N_2040,N_2347);
xor U4837 (N_4837,N_3793,N_3581);
nor U4838 (N_4838,N_2953,N_3309);
and U4839 (N_4839,N_2873,N_2020);
and U4840 (N_4840,N_3897,N_2875);
and U4841 (N_4841,N_3198,N_3385);
and U4842 (N_4842,N_3301,N_3791);
nor U4843 (N_4843,N_2067,N_2227);
xnor U4844 (N_4844,N_3810,N_2969);
or U4845 (N_4845,N_3691,N_3096);
xor U4846 (N_4846,N_2934,N_3626);
or U4847 (N_4847,N_3792,N_3711);
xor U4848 (N_4848,N_3428,N_2885);
nor U4849 (N_4849,N_2038,N_2076);
xnor U4850 (N_4850,N_3296,N_3579);
xor U4851 (N_4851,N_3430,N_3207);
xor U4852 (N_4852,N_2062,N_2881);
nor U4853 (N_4853,N_2878,N_2884);
or U4854 (N_4854,N_2487,N_2948);
xor U4855 (N_4855,N_3733,N_3554);
nor U4856 (N_4856,N_2264,N_2607);
nand U4857 (N_4857,N_3187,N_2469);
xnor U4858 (N_4858,N_2468,N_2608);
nor U4859 (N_4859,N_2031,N_3904);
nand U4860 (N_4860,N_3958,N_3488);
nand U4861 (N_4861,N_3148,N_2605);
or U4862 (N_4862,N_2294,N_3381);
nor U4863 (N_4863,N_3391,N_2141);
nor U4864 (N_4864,N_3530,N_3576);
or U4865 (N_4865,N_2681,N_3922);
nor U4866 (N_4866,N_2081,N_3820);
xnor U4867 (N_4867,N_2629,N_3008);
xor U4868 (N_4868,N_3959,N_2147);
nand U4869 (N_4869,N_2908,N_3875);
nor U4870 (N_4870,N_2739,N_3227);
nor U4871 (N_4871,N_2728,N_2765);
xnor U4872 (N_4872,N_2560,N_3539);
nor U4873 (N_4873,N_3784,N_2830);
or U4874 (N_4874,N_3378,N_3467);
or U4875 (N_4875,N_3486,N_3754);
nor U4876 (N_4876,N_2595,N_2844);
nor U4877 (N_4877,N_2616,N_2650);
xnor U4878 (N_4878,N_2122,N_2651);
nand U4879 (N_4879,N_2806,N_3230);
xnor U4880 (N_4880,N_3612,N_2922);
xnor U4881 (N_4881,N_2066,N_2357);
or U4882 (N_4882,N_3547,N_3213);
xnor U4883 (N_4883,N_3427,N_3271);
nor U4884 (N_4884,N_3071,N_2015);
nor U4885 (N_4885,N_2710,N_3957);
nand U4886 (N_4886,N_2479,N_3163);
xor U4887 (N_4887,N_3220,N_2824);
or U4888 (N_4888,N_3658,N_2868);
nor U4889 (N_4889,N_3460,N_3971);
and U4890 (N_4890,N_3606,N_3287);
nor U4891 (N_4891,N_3169,N_2082);
xnor U4892 (N_4892,N_3452,N_3525);
nor U4893 (N_4893,N_3051,N_2140);
nor U4894 (N_4894,N_2459,N_3635);
nand U4895 (N_4895,N_2449,N_3132);
nor U4896 (N_4896,N_3114,N_2280);
and U4897 (N_4897,N_2627,N_2764);
xor U4898 (N_4898,N_2497,N_2379);
nand U4899 (N_4899,N_3047,N_2484);
and U4900 (N_4900,N_3424,N_3272);
and U4901 (N_4901,N_2012,N_2203);
nand U4902 (N_4902,N_2679,N_3344);
or U4903 (N_4903,N_3852,N_3330);
xor U4904 (N_4904,N_3027,N_3431);
nand U4905 (N_4905,N_3701,N_3363);
or U4906 (N_4906,N_3765,N_2705);
and U4907 (N_4907,N_3090,N_2146);
and U4908 (N_4908,N_3039,N_3248);
and U4909 (N_4909,N_2311,N_2345);
or U4910 (N_4910,N_3956,N_2888);
nor U4911 (N_4911,N_3413,N_2016);
and U4912 (N_4912,N_2064,N_2537);
nand U4913 (N_4913,N_2480,N_3999);
and U4914 (N_4914,N_2033,N_2585);
or U4915 (N_4915,N_3570,N_2571);
and U4916 (N_4916,N_3985,N_2216);
nor U4917 (N_4917,N_3158,N_2121);
nor U4918 (N_4918,N_3556,N_2413);
nand U4919 (N_4919,N_3824,N_3885);
or U4920 (N_4920,N_3084,N_3874);
nand U4921 (N_4921,N_2704,N_3331);
nor U4922 (N_4922,N_2640,N_3018);
nor U4923 (N_4923,N_2790,N_3533);
nand U4924 (N_4924,N_3725,N_3664);
nor U4925 (N_4925,N_2461,N_3049);
or U4926 (N_4926,N_2004,N_2194);
nor U4927 (N_4927,N_3861,N_2897);
nor U4928 (N_4928,N_3849,N_3067);
and U4929 (N_4929,N_2935,N_2787);
or U4930 (N_4930,N_3704,N_3057);
nor U4931 (N_4931,N_2153,N_3238);
and U4932 (N_4932,N_3833,N_3941);
and U4933 (N_4933,N_3662,N_2231);
nand U4934 (N_4934,N_3328,N_3437);
nor U4935 (N_4935,N_2104,N_2162);
xnor U4936 (N_4936,N_2386,N_2072);
xor U4937 (N_4937,N_2702,N_3365);
or U4938 (N_4938,N_2547,N_3473);
nor U4939 (N_4939,N_3060,N_2456);
xor U4940 (N_4940,N_2060,N_2886);
nand U4941 (N_4941,N_3192,N_2333);
nand U4942 (N_4942,N_3644,N_3728);
xnor U4943 (N_4943,N_3323,N_2614);
nor U4944 (N_4944,N_3115,N_3511);
nand U4945 (N_4945,N_2843,N_3795);
and U4946 (N_4946,N_3913,N_2717);
xnor U4947 (N_4947,N_3882,N_2927);
xnor U4948 (N_4948,N_3489,N_3796);
nor U4949 (N_4949,N_2183,N_3813);
and U4950 (N_4950,N_2132,N_2369);
nor U4951 (N_4951,N_3300,N_3412);
nor U4952 (N_4952,N_3108,N_3847);
nand U4953 (N_4953,N_3601,N_3697);
or U4954 (N_4954,N_3372,N_2287);
nor U4955 (N_4955,N_3954,N_2762);
and U4956 (N_4956,N_2467,N_3532);
or U4957 (N_4957,N_2473,N_2505);
nand U4958 (N_4958,N_3973,N_3349);
xor U4959 (N_4959,N_2997,N_3919);
nand U4960 (N_4960,N_2993,N_3910);
nor U4961 (N_4961,N_3455,N_3172);
nor U4962 (N_4962,N_3744,N_3199);
xnor U4963 (N_4963,N_3293,N_2118);
nand U4964 (N_4964,N_3497,N_2166);
and U4965 (N_4965,N_2818,N_2193);
and U4966 (N_4966,N_2446,N_2324);
nand U4967 (N_4967,N_3745,N_3698);
nor U4968 (N_4968,N_3571,N_3613);
nand U4969 (N_4969,N_2815,N_2408);
or U4970 (N_4970,N_2126,N_3036);
nand U4971 (N_4971,N_3770,N_3965);
or U4972 (N_4972,N_3531,N_3418);
and U4973 (N_4973,N_3840,N_2528);
xor U4974 (N_4974,N_3105,N_3274);
xnor U4975 (N_4975,N_2353,N_2045);
nand U4976 (N_4976,N_3201,N_2816);
xor U4977 (N_4977,N_3540,N_2671);
nor U4978 (N_4978,N_2502,N_2721);
nor U4979 (N_4979,N_2377,N_3566);
nand U4980 (N_4980,N_2109,N_3895);
xor U4981 (N_4981,N_3070,N_3125);
and U4982 (N_4982,N_2375,N_3769);
nand U4983 (N_4983,N_3674,N_2709);
xnor U4984 (N_4984,N_2777,N_3598);
nand U4985 (N_4985,N_2321,N_2490);
and U4986 (N_4986,N_3834,N_2542);
and U4987 (N_4987,N_3336,N_3625);
nor U4988 (N_4988,N_3321,N_2069);
nand U4989 (N_4989,N_2304,N_3599);
nor U4990 (N_4990,N_2342,N_3610);
nand U4991 (N_4991,N_3976,N_2441);
nand U4992 (N_4992,N_3675,N_3578);
nand U4993 (N_4993,N_3433,N_2669);
and U4994 (N_4994,N_3367,N_2538);
nand U4995 (N_4995,N_3268,N_3969);
nor U4996 (N_4996,N_2035,N_2735);
or U4997 (N_4997,N_3615,N_3666);
and U4998 (N_4998,N_2130,N_2569);
or U4999 (N_4999,N_3643,N_2187);
nor U5000 (N_5000,N_3549,N_3146);
xnor U5001 (N_5001,N_2331,N_2186);
or U5002 (N_5002,N_3328,N_2470);
or U5003 (N_5003,N_3326,N_2694);
xnor U5004 (N_5004,N_2786,N_3171);
nand U5005 (N_5005,N_2794,N_3723);
or U5006 (N_5006,N_3307,N_3117);
and U5007 (N_5007,N_2540,N_3948);
xor U5008 (N_5008,N_3239,N_3292);
and U5009 (N_5009,N_3340,N_2656);
xnor U5010 (N_5010,N_3245,N_2379);
and U5011 (N_5011,N_3864,N_3513);
and U5012 (N_5012,N_2041,N_3974);
and U5013 (N_5013,N_2045,N_3461);
nor U5014 (N_5014,N_3285,N_3342);
nand U5015 (N_5015,N_3664,N_2713);
nand U5016 (N_5016,N_2052,N_2097);
nor U5017 (N_5017,N_2024,N_2060);
xnor U5018 (N_5018,N_3466,N_3638);
xnor U5019 (N_5019,N_3888,N_2891);
xor U5020 (N_5020,N_3720,N_2937);
nor U5021 (N_5021,N_2500,N_2076);
xnor U5022 (N_5022,N_2871,N_3158);
nand U5023 (N_5023,N_3641,N_3545);
xor U5024 (N_5024,N_3733,N_3608);
nand U5025 (N_5025,N_3536,N_2188);
and U5026 (N_5026,N_2121,N_2822);
nor U5027 (N_5027,N_2009,N_3501);
nor U5028 (N_5028,N_3874,N_3079);
xnor U5029 (N_5029,N_3125,N_3823);
nand U5030 (N_5030,N_3770,N_3056);
nor U5031 (N_5031,N_2475,N_2737);
and U5032 (N_5032,N_3327,N_2008);
or U5033 (N_5033,N_2125,N_2894);
or U5034 (N_5034,N_2934,N_2854);
or U5035 (N_5035,N_3803,N_3949);
nor U5036 (N_5036,N_3420,N_2372);
nor U5037 (N_5037,N_3308,N_3546);
nor U5038 (N_5038,N_3858,N_2108);
nand U5039 (N_5039,N_3073,N_3264);
nand U5040 (N_5040,N_2753,N_2163);
or U5041 (N_5041,N_2683,N_3074);
xnor U5042 (N_5042,N_3113,N_2676);
and U5043 (N_5043,N_2669,N_3016);
nand U5044 (N_5044,N_3352,N_3145);
nand U5045 (N_5045,N_2656,N_2983);
xor U5046 (N_5046,N_2008,N_2401);
and U5047 (N_5047,N_3471,N_2229);
and U5048 (N_5048,N_3604,N_2900);
and U5049 (N_5049,N_3760,N_2189);
nor U5050 (N_5050,N_2003,N_3119);
or U5051 (N_5051,N_2757,N_2936);
nand U5052 (N_5052,N_2437,N_2818);
or U5053 (N_5053,N_2798,N_2511);
xnor U5054 (N_5054,N_2780,N_3320);
and U5055 (N_5055,N_3322,N_3636);
or U5056 (N_5056,N_2401,N_2571);
or U5057 (N_5057,N_3004,N_3748);
nor U5058 (N_5058,N_2529,N_2419);
and U5059 (N_5059,N_2911,N_3204);
and U5060 (N_5060,N_2426,N_2679);
and U5061 (N_5061,N_3992,N_2765);
or U5062 (N_5062,N_3009,N_3807);
and U5063 (N_5063,N_3238,N_3190);
nor U5064 (N_5064,N_2143,N_2296);
or U5065 (N_5065,N_2041,N_3871);
nand U5066 (N_5066,N_3740,N_3337);
nand U5067 (N_5067,N_3520,N_2727);
xor U5068 (N_5068,N_3539,N_3596);
and U5069 (N_5069,N_3274,N_3029);
xnor U5070 (N_5070,N_3014,N_3176);
nand U5071 (N_5071,N_2242,N_2053);
and U5072 (N_5072,N_3102,N_2708);
nor U5073 (N_5073,N_3208,N_3113);
xor U5074 (N_5074,N_2306,N_2991);
xnor U5075 (N_5075,N_3910,N_3980);
or U5076 (N_5076,N_3975,N_2045);
nor U5077 (N_5077,N_3785,N_2740);
nand U5078 (N_5078,N_2883,N_2350);
or U5079 (N_5079,N_3591,N_2800);
nand U5080 (N_5080,N_2794,N_3738);
or U5081 (N_5081,N_2401,N_3697);
nor U5082 (N_5082,N_3628,N_3483);
nor U5083 (N_5083,N_3212,N_2272);
xnor U5084 (N_5084,N_3084,N_3217);
or U5085 (N_5085,N_2496,N_3762);
nand U5086 (N_5086,N_3704,N_2694);
xor U5087 (N_5087,N_2569,N_2339);
and U5088 (N_5088,N_3261,N_2625);
nand U5089 (N_5089,N_3456,N_3643);
xnor U5090 (N_5090,N_3390,N_2182);
and U5091 (N_5091,N_3731,N_3686);
xnor U5092 (N_5092,N_2422,N_3420);
nand U5093 (N_5093,N_2658,N_2900);
and U5094 (N_5094,N_2145,N_3961);
or U5095 (N_5095,N_3585,N_3929);
and U5096 (N_5096,N_2637,N_3513);
and U5097 (N_5097,N_3503,N_3496);
and U5098 (N_5098,N_3352,N_3229);
xnor U5099 (N_5099,N_3276,N_2202);
and U5100 (N_5100,N_3543,N_2642);
xnor U5101 (N_5101,N_2861,N_2909);
nand U5102 (N_5102,N_3184,N_2894);
or U5103 (N_5103,N_2483,N_3330);
nand U5104 (N_5104,N_3530,N_3400);
and U5105 (N_5105,N_2724,N_2381);
or U5106 (N_5106,N_3214,N_2456);
nor U5107 (N_5107,N_3192,N_2425);
nand U5108 (N_5108,N_3025,N_3680);
xnor U5109 (N_5109,N_3824,N_3841);
or U5110 (N_5110,N_2071,N_2833);
xnor U5111 (N_5111,N_3585,N_3363);
and U5112 (N_5112,N_3219,N_2784);
and U5113 (N_5113,N_3070,N_2754);
nand U5114 (N_5114,N_3670,N_3119);
or U5115 (N_5115,N_3439,N_2060);
nor U5116 (N_5116,N_3096,N_3194);
nor U5117 (N_5117,N_2597,N_3580);
xnor U5118 (N_5118,N_2840,N_2682);
and U5119 (N_5119,N_3726,N_3499);
or U5120 (N_5120,N_3217,N_2185);
and U5121 (N_5121,N_3897,N_3314);
and U5122 (N_5122,N_3062,N_2176);
nor U5123 (N_5123,N_2839,N_3273);
xnor U5124 (N_5124,N_2452,N_3562);
xor U5125 (N_5125,N_2006,N_2048);
xor U5126 (N_5126,N_2572,N_2185);
or U5127 (N_5127,N_2081,N_2666);
nand U5128 (N_5128,N_2405,N_2184);
nand U5129 (N_5129,N_2994,N_3615);
nor U5130 (N_5130,N_3898,N_2949);
nor U5131 (N_5131,N_3288,N_2477);
nor U5132 (N_5132,N_2441,N_2964);
nor U5133 (N_5133,N_3647,N_3983);
xnor U5134 (N_5134,N_2181,N_2899);
nand U5135 (N_5135,N_2126,N_2985);
xnor U5136 (N_5136,N_3342,N_2353);
nor U5137 (N_5137,N_3165,N_3752);
nor U5138 (N_5138,N_3851,N_3657);
xor U5139 (N_5139,N_3131,N_2658);
or U5140 (N_5140,N_2299,N_3636);
and U5141 (N_5141,N_2397,N_3919);
nor U5142 (N_5142,N_2998,N_3848);
or U5143 (N_5143,N_3804,N_2533);
xnor U5144 (N_5144,N_2451,N_3781);
nand U5145 (N_5145,N_3719,N_2813);
xnor U5146 (N_5146,N_2451,N_3137);
nand U5147 (N_5147,N_3805,N_3738);
nand U5148 (N_5148,N_3210,N_2578);
and U5149 (N_5149,N_3269,N_2697);
nor U5150 (N_5150,N_2821,N_2492);
nor U5151 (N_5151,N_2084,N_2136);
nand U5152 (N_5152,N_3081,N_2725);
xnor U5153 (N_5153,N_2008,N_3185);
or U5154 (N_5154,N_3073,N_2155);
or U5155 (N_5155,N_2744,N_3203);
nand U5156 (N_5156,N_3898,N_3038);
or U5157 (N_5157,N_2724,N_3411);
nand U5158 (N_5158,N_3612,N_2342);
and U5159 (N_5159,N_2513,N_2420);
nand U5160 (N_5160,N_2564,N_3786);
or U5161 (N_5161,N_2295,N_3961);
and U5162 (N_5162,N_2556,N_3684);
and U5163 (N_5163,N_3025,N_2399);
nor U5164 (N_5164,N_3960,N_2254);
nor U5165 (N_5165,N_3866,N_2441);
nor U5166 (N_5166,N_3580,N_3814);
xor U5167 (N_5167,N_3717,N_3837);
xnor U5168 (N_5168,N_2487,N_3782);
nand U5169 (N_5169,N_3155,N_3759);
xor U5170 (N_5170,N_3788,N_2691);
xnor U5171 (N_5171,N_3752,N_3271);
and U5172 (N_5172,N_2007,N_2270);
or U5173 (N_5173,N_2262,N_3696);
nor U5174 (N_5174,N_2762,N_2367);
xnor U5175 (N_5175,N_2409,N_3236);
nor U5176 (N_5176,N_3994,N_3573);
or U5177 (N_5177,N_3432,N_2868);
xnor U5178 (N_5178,N_2586,N_2050);
xor U5179 (N_5179,N_2858,N_3950);
nor U5180 (N_5180,N_3033,N_3853);
and U5181 (N_5181,N_3813,N_3742);
or U5182 (N_5182,N_2657,N_2500);
or U5183 (N_5183,N_3567,N_3190);
and U5184 (N_5184,N_2899,N_2534);
and U5185 (N_5185,N_2557,N_2180);
nor U5186 (N_5186,N_2109,N_2682);
nand U5187 (N_5187,N_2305,N_2513);
or U5188 (N_5188,N_3328,N_2699);
xnor U5189 (N_5189,N_2924,N_2840);
or U5190 (N_5190,N_2255,N_3622);
xnor U5191 (N_5191,N_2689,N_3613);
nor U5192 (N_5192,N_3919,N_2751);
xnor U5193 (N_5193,N_2712,N_2354);
xor U5194 (N_5194,N_2332,N_3232);
nand U5195 (N_5195,N_2195,N_2243);
or U5196 (N_5196,N_3815,N_2635);
nand U5197 (N_5197,N_3826,N_2146);
or U5198 (N_5198,N_3501,N_3165);
xnor U5199 (N_5199,N_3974,N_2987);
xnor U5200 (N_5200,N_2223,N_3991);
or U5201 (N_5201,N_2946,N_2362);
and U5202 (N_5202,N_3952,N_2879);
xnor U5203 (N_5203,N_3747,N_3773);
nor U5204 (N_5204,N_3791,N_3029);
and U5205 (N_5205,N_2164,N_3880);
nor U5206 (N_5206,N_3995,N_2678);
nand U5207 (N_5207,N_2781,N_3178);
and U5208 (N_5208,N_3975,N_3021);
or U5209 (N_5209,N_3607,N_2275);
nand U5210 (N_5210,N_3914,N_2299);
xor U5211 (N_5211,N_2770,N_3225);
nand U5212 (N_5212,N_2659,N_3930);
nand U5213 (N_5213,N_2884,N_3309);
and U5214 (N_5214,N_2726,N_3000);
or U5215 (N_5215,N_2973,N_2593);
nand U5216 (N_5216,N_3573,N_3921);
and U5217 (N_5217,N_3068,N_2635);
nor U5218 (N_5218,N_2369,N_2628);
and U5219 (N_5219,N_2694,N_2141);
nand U5220 (N_5220,N_3688,N_3824);
xnor U5221 (N_5221,N_3582,N_3203);
nor U5222 (N_5222,N_3150,N_3201);
nor U5223 (N_5223,N_3047,N_3284);
nor U5224 (N_5224,N_2449,N_3996);
xnor U5225 (N_5225,N_3701,N_2358);
and U5226 (N_5226,N_2659,N_2543);
nor U5227 (N_5227,N_2909,N_3510);
or U5228 (N_5228,N_2272,N_3426);
nand U5229 (N_5229,N_3310,N_2159);
nor U5230 (N_5230,N_2331,N_2934);
nor U5231 (N_5231,N_2744,N_3772);
and U5232 (N_5232,N_3142,N_3249);
and U5233 (N_5233,N_2277,N_2597);
xnor U5234 (N_5234,N_3815,N_2432);
and U5235 (N_5235,N_3018,N_2352);
nor U5236 (N_5236,N_2730,N_2252);
or U5237 (N_5237,N_2122,N_2478);
and U5238 (N_5238,N_3192,N_3992);
nand U5239 (N_5239,N_3904,N_3272);
and U5240 (N_5240,N_3493,N_2978);
xnor U5241 (N_5241,N_3235,N_2095);
xor U5242 (N_5242,N_3629,N_2236);
and U5243 (N_5243,N_3313,N_2992);
nand U5244 (N_5244,N_3214,N_2057);
or U5245 (N_5245,N_3115,N_2618);
xnor U5246 (N_5246,N_2456,N_3414);
nand U5247 (N_5247,N_3400,N_2616);
nand U5248 (N_5248,N_2122,N_3944);
and U5249 (N_5249,N_2259,N_2347);
nand U5250 (N_5250,N_3330,N_3297);
nand U5251 (N_5251,N_3363,N_3533);
and U5252 (N_5252,N_2214,N_3135);
nor U5253 (N_5253,N_3380,N_2525);
and U5254 (N_5254,N_3657,N_2158);
and U5255 (N_5255,N_2023,N_2875);
or U5256 (N_5256,N_2539,N_2651);
nor U5257 (N_5257,N_3123,N_2003);
or U5258 (N_5258,N_2499,N_2580);
nor U5259 (N_5259,N_2815,N_3721);
or U5260 (N_5260,N_3100,N_2145);
nor U5261 (N_5261,N_3367,N_2419);
xor U5262 (N_5262,N_2070,N_2155);
nor U5263 (N_5263,N_2896,N_2261);
nor U5264 (N_5264,N_3604,N_2308);
nor U5265 (N_5265,N_3947,N_2445);
or U5266 (N_5266,N_2310,N_2325);
or U5267 (N_5267,N_2229,N_2310);
or U5268 (N_5268,N_2242,N_2363);
xnor U5269 (N_5269,N_2499,N_2329);
and U5270 (N_5270,N_3943,N_2101);
and U5271 (N_5271,N_2133,N_3387);
or U5272 (N_5272,N_2651,N_2801);
or U5273 (N_5273,N_3443,N_3339);
nand U5274 (N_5274,N_3422,N_2718);
xor U5275 (N_5275,N_2845,N_2914);
or U5276 (N_5276,N_2529,N_2192);
and U5277 (N_5277,N_2141,N_3622);
or U5278 (N_5278,N_3937,N_2826);
nand U5279 (N_5279,N_3520,N_3566);
nor U5280 (N_5280,N_3365,N_2219);
nor U5281 (N_5281,N_3635,N_3042);
and U5282 (N_5282,N_2673,N_2920);
xor U5283 (N_5283,N_2370,N_2904);
or U5284 (N_5284,N_2566,N_3466);
xor U5285 (N_5285,N_3519,N_2290);
nand U5286 (N_5286,N_3856,N_2626);
xnor U5287 (N_5287,N_3161,N_2041);
nand U5288 (N_5288,N_3876,N_2431);
xor U5289 (N_5289,N_3523,N_2259);
or U5290 (N_5290,N_2804,N_3484);
nand U5291 (N_5291,N_2439,N_3296);
xnor U5292 (N_5292,N_3519,N_3599);
nor U5293 (N_5293,N_3421,N_2899);
and U5294 (N_5294,N_2906,N_2985);
nand U5295 (N_5295,N_3721,N_2511);
and U5296 (N_5296,N_2327,N_3452);
nand U5297 (N_5297,N_3441,N_3163);
or U5298 (N_5298,N_3552,N_2845);
xor U5299 (N_5299,N_2582,N_3637);
and U5300 (N_5300,N_3724,N_3462);
and U5301 (N_5301,N_2290,N_2977);
xnor U5302 (N_5302,N_2128,N_3931);
xnor U5303 (N_5303,N_2204,N_3836);
nand U5304 (N_5304,N_3798,N_2822);
or U5305 (N_5305,N_2584,N_3941);
or U5306 (N_5306,N_3532,N_3654);
nor U5307 (N_5307,N_2239,N_2412);
or U5308 (N_5308,N_3058,N_3495);
or U5309 (N_5309,N_3727,N_2198);
nor U5310 (N_5310,N_3429,N_2356);
nand U5311 (N_5311,N_3763,N_3442);
or U5312 (N_5312,N_3104,N_3081);
nor U5313 (N_5313,N_3618,N_2619);
and U5314 (N_5314,N_3328,N_3489);
and U5315 (N_5315,N_3107,N_2136);
nand U5316 (N_5316,N_2878,N_3516);
nand U5317 (N_5317,N_3635,N_2769);
xnor U5318 (N_5318,N_2794,N_2576);
xor U5319 (N_5319,N_2626,N_2725);
or U5320 (N_5320,N_2020,N_3492);
xnor U5321 (N_5321,N_2076,N_3895);
xnor U5322 (N_5322,N_3499,N_2413);
and U5323 (N_5323,N_3763,N_2776);
xnor U5324 (N_5324,N_2877,N_2908);
nor U5325 (N_5325,N_2654,N_3428);
nand U5326 (N_5326,N_3832,N_2073);
and U5327 (N_5327,N_3215,N_3821);
xor U5328 (N_5328,N_2066,N_3025);
nand U5329 (N_5329,N_2496,N_3108);
nand U5330 (N_5330,N_3234,N_3324);
xor U5331 (N_5331,N_2173,N_2158);
and U5332 (N_5332,N_3891,N_2031);
and U5333 (N_5333,N_3912,N_3586);
nand U5334 (N_5334,N_2779,N_2485);
or U5335 (N_5335,N_3710,N_2549);
xnor U5336 (N_5336,N_2378,N_2546);
nand U5337 (N_5337,N_3064,N_2103);
and U5338 (N_5338,N_3408,N_3962);
nor U5339 (N_5339,N_2345,N_2121);
or U5340 (N_5340,N_2837,N_2418);
and U5341 (N_5341,N_3378,N_2767);
nand U5342 (N_5342,N_2272,N_3226);
nor U5343 (N_5343,N_3844,N_3864);
nand U5344 (N_5344,N_2317,N_3515);
nor U5345 (N_5345,N_3491,N_2143);
xor U5346 (N_5346,N_3577,N_3614);
nand U5347 (N_5347,N_3546,N_3146);
nor U5348 (N_5348,N_2765,N_3647);
nand U5349 (N_5349,N_2629,N_3827);
nand U5350 (N_5350,N_2952,N_3924);
or U5351 (N_5351,N_2442,N_3170);
nand U5352 (N_5352,N_2669,N_2046);
nand U5353 (N_5353,N_2600,N_3216);
nor U5354 (N_5354,N_2342,N_2111);
nand U5355 (N_5355,N_2010,N_3317);
and U5356 (N_5356,N_3366,N_3910);
and U5357 (N_5357,N_2396,N_3631);
nor U5358 (N_5358,N_3108,N_3927);
nor U5359 (N_5359,N_3658,N_2874);
nor U5360 (N_5360,N_3808,N_3346);
or U5361 (N_5361,N_2003,N_3096);
and U5362 (N_5362,N_3920,N_2824);
xnor U5363 (N_5363,N_3145,N_3026);
nor U5364 (N_5364,N_2269,N_2186);
or U5365 (N_5365,N_3179,N_2567);
xnor U5366 (N_5366,N_3088,N_2789);
or U5367 (N_5367,N_3868,N_2575);
nand U5368 (N_5368,N_2987,N_2798);
nand U5369 (N_5369,N_2963,N_2516);
nor U5370 (N_5370,N_2608,N_3420);
and U5371 (N_5371,N_3803,N_3493);
or U5372 (N_5372,N_2626,N_3961);
xor U5373 (N_5373,N_2800,N_3139);
nor U5374 (N_5374,N_2020,N_2622);
nor U5375 (N_5375,N_3941,N_2047);
and U5376 (N_5376,N_2777,N_3661);
nor U5377 (N_5377,N_3138,N_2756);
or U5378 (N_5378,N_3205,N_3752);
and U5379 (N_5379,N_3565,N_3797);
nand U5380 (N_5380,N_2607,N_2938);
nor U5381 (N_5381,N_2437,N_3268);
nand U5382 (N_5382,N_2838,N_2658);
nand U5383 (N_5383,N_3763,N_3043);
xnor U5384 (N_5384,N_2454,N_2363);
or U5385 (N_5385,N_3709,N_2051);
or U5386 (N_5386,N_2817,N_2753);
xnor U5387 (N_5387,N_3508,N_2200);
and U5388 (N_5388,N_3930,N_3913);
nor U5389 (N_5389,N_2243,N_2761);
nor U5390 (N_5390,N_3731,N_3448);
or U5391 (N_5391,N_2206,N_2559);
xor U5392 (N_5392,N_3103,N_3295);
nand U5393 (N_5393,N_2569,N_3851);
or U5394 (N_5394,N_2481,N_3695);
or U5395 (N_5395,N_2291,N_3523);
nand U5396 (N_5396,N_3822,N_3173);
nor U5397 (N_5397,N_2609,N_3000);
nor U5398 (N_5398,N_2777,N_3755);
xor U5399 (N_5399,N_3365,N_3610);
nor U5400 (N_5400,N_3018,N_3940);
nor U5401 (N_5401,N_2935,N_3920);
xnor U5402 (N_5402,N_3887,N_2625);
and U5403 (N_5403,N_3241,N_2053);
nand U5404 (N_5404,N_3800,N_3397);
and U5405 (N_5405,N_2678,N_3845);
and U5406 (N_5406,N_3657,N_3081);
nand U5407 (N_5407,N_3440,N_2718);
nor U5408 (N_5408,N_3904,N_2184);
nor U5409 (N_5409,N_3892,N_3482);
nor U5410 (N_5410,N_3923,N_2246);
or U5411 (N_5411,N_2375,N_2366);
or U5412 (N_5412,N_2486,N_2301);
and U5413 (N_5413,N_3699,N_2892);
and U5414 (N_5414,N_2458,N_3495);
xor U5415 (N_5415,N_3060,N_3961);
or U5416 (N_5416,N_2258,N_2472);
or U5417 (N_5417,N_3089,N_3534);
nor U5418 (N_5418,N_2956,N_3270);
xnor U5419 (N_5419,N_2514,N_3989);
and U5420 (N_5420,N_2335,N_2417);
nand U5421 (N_5421,N_2405,N_2076);
nor U5422 (N_5422,N_3011,N_3944);
nor U5423 (N_5423,N_3686,N_2492);
nor U5424 (N_5424,N_3459,N_3085);
nand U5425 (N_5425,N_3978,N_2482);
xnor U5426 (N_5426,N_3952,N_3558);
xor U5427 (N_5427,N_2580,N_2521);
xor U5428 (N_5428,N_3003,N_3193);
or U5429 (N_5429,N_3530,N_3744);
xor U5430 (N_5430,N_2098,N_2840);
or U5431 (N_5431,N_3023,N_3137);
or U5432 (N_5432,N_3427,N_3604);
xnor U5433 (N_5433,N_3163,N_2512);
xor U5434 (N_5434,N_2220,N_2921);
or U5435 (N_5435,N_2494,N_3650);
xor U5436 (N_5436,N_2649,N_3747);
xor U5437 (N_5437,N_3962,N_2591);
xor U5438 (N_5438,N_3930,N_2711);
xor U5439 (N_5439,N_3266,N_2245);
xnor U5440 (N_5440,N_3241,N_3398);
and U5441 (N_5441,N_2558,N_2212);
xnor U5442 (N_5442,N_2234,N_2747);
xor U5443 (N_5443,N_2063,N_2633);
nor U5444 (N_5444,N_3385,N_3912);
nor U5445 (N_5445,N_3344,N_2449);
or U5446 (N_5446,N_3559,N_3038);
and U5447 (N_5447,N_2845,N_3056);
or U5448 (N_5448,N_2884,N_2611);
and U5449 (N_5449,N_2904,N_3784);
nand U5450 (N_5450,N_3542,N_3206);
or U5451 (N_5451,N_3858,N_3372);
and U5452 (N_5452,N_3407,N_3022);
xor U5453 (N_5453,N_2365,N_3810);
nand U5454 (N_5454,N_2975,N_2796);
nand U5455 (N_5455,N_2458,N_2942);
nand U5456 (N_5456,N_3615,N_3402);
nand U5457 (N_5457,N_2015,N_2136);
nand U5458 (N_5458,N_2375,N_2940);
or U5459 (N_5459,N_2945,N_3628);
or U5460 (N_5460,N_2072,N_3054);
and U5461 (N_5461,N_3154,N_2020);
and U5462 (N_5462,N_3233,N_2091);
nor U5463 (N_5463,N_2079,N_3205);
nand U5464 (N_5464,N_2295,N_2735);
and U5465 (N_5465,N_2152,N_3836);
and U5466 (N_5466,N_2173,N_2296);
nand U5467 (N_5467,N_3778,N_2192);
nor U5468 (N_5468,N_2992,N_3664);
xor U5469 (N_5469,N_2730,N_3527);
xor U5470 (N_5470,N_2083,N_3058);
and U5471 (N_5471,N_3146,N_2023);
nand U5472 (N_5472,N_3856,N_2434);
nand U5473 (N_5473,N_2144,N_2831);
nor U5474 (N_5474,N_2531,N_2648);
nor U5475 (N_5475,N_2711,N_3147);
and U5476 (N_5476,N_2634,N_2405);
or U5477 (N_5477,N_3227,N_2514);
and U5478 (N_5478,N_3105,N_3834);
xor U5479 (N_5479,N_3627,N_2497);
or U5480 (N_5480,N_2334,N_3493);
nand U5481 (N_5481,N_3687,N_2682);
xor U5482 (N_5482,N_2353,N_2028);
and U5483 (N_5483,N_3885,N_2456);
nor U5484 (N_5484,N_3402,N_2837);
nor U5485 (N_5485,N_2290,N_2630);
and U5486 (N_5486,N_3798,N_2513);
nand U5487 (N_5487,N_3088,N_2493);
nand U5488 (N_5488,N_2336,N_2013);
nand U5489 (N_5489,N_2115,N_3335);
nand U5490 (N_5490,N_3551,N_2450);
nor U5491 (N_5491,N_3032,N_2717);
nand U5492 (N_5492,N_2543,N_2519);
nand U5493 (N_5493,N_3312,N_3284);
nor U5494 (N_5494,N_2955,N_2953);
nor U5495 (N_5495,N_3460,N_2037);
xnor U5496 (N_5496,N_2849,N_2802);
or U5497 (N_5497,N_3162,N_2064);
and U5498 (N_5498,N_3508,N_3463);
and U5499 (N_5499,N_2169,N_3392);
nor U5500 (N_5500,N_2088,N_2796);
or U5501 (N_5501,N_3166,N_2077);
xor U5502 (N_5502,N_2269,N_2849);
nand U5503 (N_5503,N_2842,N_3875);
nor U5504 (N_5504,N_3885,N_2465);
xnor U5505 (N_5505,N_3895,N_3178);
or U5506 (N_5506,N_3195,N_2538);
xnor U5507 (N_5507,N_3970,N_3805);
or U5508 (N_5508,N_2979,N_2066);
xnor U5509 (N_5509,N_2688,N_2260);
xnor U5510 (N_5510,N_2854,N_3300);
or U5511 (N_5511,N_2570,N_2913);
xnor U5512 (N_5512,N_3214,N_3287);
xnor U5513 (N_5513,N_3216,N_3954);
nand U5514 (N_5514,N_2967,N_2734);
or U5515 (N_5515,N_3612,N_2312);
and U5516 (N_5516,N_2893,N_3948);
and U5517 (N_5517,N_3320,N_2453);
and U5518 (N_5518,N_3306,N_3144);
and U5519 (N_5519,N_3188,N_3584);
xor U5520 (N_5520,N_2166,N_2679);
and U5521 (N_5521,N_3143,N_2508);
or U5522 (N_5522,N_2286,N_3973);
and U5523 (N_5523,N_2283,N_3447);
or U5524 (N_5524,N_3180,N_2613);
nand U5525 (N_5525,N_2263,N_2151);
nand U5526 (N_5526,N_2309,N_2136);
nand U5527 (N_5527,N_3866,N_3434);
xnor U5528 (N_5528,N_3888,N_2077);
xor U5529 (N_5529,N_2538,N_3112);
xor U5530 (N_5530,N_2003,N_3976);
nand U5531 (N_5531,N_3834,N_3049);
or U5532 (N_5532,N_3517,N_3057);
and U5533 (N_5533,N_2665,N_3848);
or U5534 (N_5534,N_2863,N_2317);
xor U5535 (N_5535,N_2273,N_2894);
and U5536 (N_5536,N_2729,N_3599);
nand U5537 (N_5537,N_3780,N_2524);
xnor U5538 (N_5538,N_2097,N_3684);
nand U5539 (N_5539,N_3201,N_3076);
nand U5540 (N_5540,N_3196,N_2045);
nand U5541 (N_5541,N_2734,N_2175);
xor U5542 (N_5542,N_2425,N_2021);
xnor U5543 (N_5543,N_2637,N_2202);
xor U5544 (N_5544,N_3872,N_2454);
xor U5545 (N_5545,N_3420,N_3071);
nand U5546 (N_5546,N_3207,N_2503);
and U5547 (N_5547,N_2236,N_2577);
nand U5548 (N_5548,N_2941,N_2957);
or U5549 (N_5549,N_2433,N_2411);
xnor U5550 (N_5550,N_3613,N_3251);
nand U5551 (N_5551,N_3067,N_2859);
xor U5552 (N_5552,N_3910,N_3063);
nor U5553 (N_5553,N_2726,N_3802);
xor U5554 (N_5554,N_3982,N_2030);
xor U5555 (N_5555,N_2512,N_3079);
nand U5556 (N_5556,N_3230,N_2324);
or U5557 (N_5557,N_2861,N_3433);
nor U5558 (N_5558,N_2184,N_3650);
and U5559 (N_5559,N_2932,N_3728);
and U5560 (N_5560,N_2494,N_2943);
nor U5561 (N_5561,N_2759,N_2129);
xnor U5562 (N_5562,N_2804,N_2271);
and U5563 (N_5563,N_3641,N_2539);
xnor U5564 (N_5564,N_3003,N_3433);
nor U5565 (N_5565,N_2272,N_2310);
nand U5566 (N_5566,N_3326,N_2484);
and U5567 (N_5567,N_2316,N_2354);
or U5568 (N_5568,N_2794,N_3336);
nand U5569 (N_5569,N_2872,N_2851);
xor U5570 (N_5570,N_2610,N_2198);
nor U5571 (N_5571,N_3224,N_2256);
nor U5572 (N_5572,N_3042,N_3274);
and U5573 (N_5573,N_2789,N_3024);
or U5574 (N_5574,N_3342,N_3549);
and U5575 (N_5575,N_3700,N_2865);
nor U5576 (N_5576,N_3590,N_3705);
or U5577 (N_5577,N_3347,N_2757);
nand U5578 (N_5578,N_2360,N_2642);
nand U5579 (N_5579,N_3367,N_3507);
xor U5580 (N_5580,N_3167,N_2826);
xnor U5581 (N_5581,N_2508,N_2731);
or U5582 (N_5582,N_3158,N_3400);
and U5583 (N_5583,N_3318,N_2434);
or U5584 (N_5584,N_3852,N_2315);
xnor U5585 (N_5585,N_3343,N_2980);
or U5586 (N_5586,N_2100,N_2854);
nand U5587 (N_5587,N_3308,N_2742);
or U5588 (N_5588,N_3828,N_2517);
nor U5589 (N_5589,N_2990,N_2626);
xnor U5590 (N_5590,N_3784,N_2853);
nand U5591 (N_5591,N_2996,N_3192);
or U5592 (N_5592,N_2477,N_3065);
and U5593 (N_5593,N_3772,N_2416);
nor U5594 (N_5594,N_2763,N_2855);
nand U5595 (N_5595,N_3668,N_2257);
or U5596 (N_5596,N_2533,N_3885);
or U5597 (N_5597,N_3802,N_2653);
xnor U5598 (N_5598,N_2164,N_3943);
and U5599 (N_5599,N_2253,N_2536);
or U5600 (N_5600,N_3472,N_2891);
or U5601 (N_5601,N_3469,N_3314);
nand U5602 (N_5602,N_2895,N_2044);
nor U5603 (N_5603,N_2092,N_2920);
and U5604 (N_5604,N_2060,N_2257);
xor U5605 (N_5605,N_3828,N_2163);
nand U5606 (N_5606,N_2222,N_2923);
nand U5607 (N_5607,N_2151,N_3387);
or U5608 (N_5608,N_3557,N_3255);
xnor U5609 (N_5609,N_3200,N_3450);
and U5610 (N_5610,N_3115,N_3679);
xor U5611 (N_5611,N_2221,N_3842);
nand U5612 (N_5612,N_3906,N_2351);
nor U5613 (N_5613,N_3032,N_2466);
nand U5614 (N_5614,N_3929,N_3050);
xor U5615 (N_5615,N_3971,N_3668);
xnor U5616 (N_5616,N_2814,N_2107);
xnor U5617 (N_5617,N_3685,N_2234);
and U5618 (N_5618,N_3117,N_2409);
nand U5619 (N_5619,N_3553,N_2846);
or U5620 (N_5620,N_2040,N_3789);
nor U5621 (N_5621,N_3332,N_3772);
nor U5622 (N_5622,N_2781,N_2003);
xor U5623 (N_5623,N_2976,N_3453);
nor U5624 (N_5624,N_3047,N_3732);
xor U5625 (N_5625,N_3970,N_2712);
nand U5626 (N_5626,N_3353,N_3501);
and U5627 (N_5627,N_3183,N_2619);
or U5628 (N_5628,N_3796,N_3297);
nand U5629 (N_5629,N_2021,N_2431);
nor U5630 (N_5630,N_2355,N_2233);
xor U5631 (N_5631,N_2173,N_2090);
xnor U5632 (N_5632,N_2485,N_2143);
nand U5633 (N_5633,N_2504,N_3997);
or U5634 (N_5634,N_3667,N_3195);
nand U5635 (N_5635,N_2859,N_2268);
and U5636 (N_5636,N_3982,N_2802);
nor U5637 (N_5637,N_3564,N_3637);
xor U5638 (N_5638,N_3335,N_3665);
nand U5639 (N_5639,N_3050,N_3421);
nor U5640 (N_5640,N_2348,N_3965);
xnor U5641 (N_5641,N_3380,N_2596);
nor U5642 (N_5642,N_3791,N_2699);
xor U5643 (N_5643,N_2674,N_2718);
xnor U5644 (N_5644,N_3100,N_2849);
or U5645 (N_5645,N_2356,N_3146);
and U5646 (N_5646,N_3244,N_3205);
nor U5647 (N_5647,N_2094,N_3785);
nand U5648 (N_5648,N_2676,N_2675);
xor U5649 (N_5649,N_2109,N_2375);
nor U5650 (N_5650,N_2706,N_3008);
or U5651 (N_5651,N_2970,N_2098);
nand U5652 (N_5652,N_2640,N_3621);
or U5653 (N_5653,N_3598,N_2609);
nand U5654 (N_5654,N_2967,N_2178);
xnor U5655 (N_5655,N_3055,N_3314);
nor U5656 (N_5656,N_2639,N_2210);
nor U5657 (N_5657,N_3815,N_3157);
or U5658 (N_5658,N_2826,N_2366);
and U5659 (N_5659,N_2308,N_3349);
nand U5660 (N_5660,N_3958,N_3891);
xor U5661 (N_5661,N_2535,N_2736);
and U5662 (N_5662,N_3986,N_3502);
nor U5663 (N_5663,N_3296,N_3892);
xnor U5664 (N_5664,N_2280,N_3522);
xor U5665 (N_5665,N_3352,N_3808);
nand U5666 (N_5666,N_3519,N_3274);
and U5667 (N_5667,N_2122,N_2064);
or U5668 (N_5668,N_3051,N_2106);
nor U5669 (N_5669,N_2901,N_2968);
xor U5670 (N_5670,N_3348,N_2221);
xnor U5671 (N_5671,N_3458,N_3440);
or U5672 (N_5672,N_2218,N_2880);
or U5673 (N_5673,N_2792,N_3362);
or U5674 (N_5674,N_2341,N_3245);
or U5675 (N_5675,N_2291,N_3959);
xor U5676 (N_5676,N_2428,N_3061);
nand U5677 (N_5677,N_3194,N_2639);
or U5678 (N_5678,N_3070,N_2229);
xnor U5679 (N_5679,N_3087,N_3743);
nor U5680 (N_5680,N_3844,N_3954);
nand U5681 (N_5681,N_2173,N_3417);
and U5682 (N_5682,N_2728,N_3830);
or U5683 (N_5683,N_2927,N_2021);
nor U5684 (N_5684,N_3532,N_3485);
xnor U5685 (N_5685,N_3956,N_3208);
nor U5686 (N_5686,N_2440,N_2157);
nand U5687 (N_5687,N_2661,N_3397);
nor U5688 (N_5688,N_2213,N_3568);
nand U5689 (N_5689,N_3400,N_3076);
xor U5690 (N_5690,N_2616,N_2798);
or U5691 (N_5691,N_2803,N_2503);
nand U5692 (N_5692,N_3518,N_2842);
and U5693 (N_5693,N_2609,N_2645);
xor U5694 (N_5694,N_2576,N_3993);
nand U5695 (N_5695,N_2242,N_2902);
nand U5696 (N_5696,N_2680,N_3284);
and U5697 (N_5697,N_3361,N_2448);
nor U5698 (N_5698,N_2243,N_3422);
or U5699 (N_5699,N_2668,N_3993);
nor U5700 (N_5700,N_2617,N_3887);
xor U5701 (N_5701,N_3430,N_3937);
xor U5702 (N_5702,N_2305,N_3681);
nor U5703 (N_5703,N_2209,N_2758);
xnor U5704 (N_5704,N_2987,N_3671);
xnor U5705 (N_5705,N_2143,N_2001);
nor U5706 (N_5706,N_2301,N_2900);
and U5707 (N_5707,N_2167,N_2981);
nor U5708 (N_5708,N_3925,N_3494);
or U5709 (N_5709,N_3483,N_3010);
or U5710 (N_5710,N_3630,N_3066);
or U5711 (N_5711,N_3253,N_2503);
or U5712 (N_5712,N_3491,N_3634);
nor U5713 (N_5713,N_2904,N_3843);
or U5714 (N_5714,N_2454,N_2790);
xnor U5715 (N_5715,N_3674,N_2676);
and U5716 (N_5716,N_3304,N_3237);
nand U5717 (N_5717,N_3909,N_3682);
or U5718 (N_5718,N_2920,N_3953);
xnor U5719 (N_5719,N_2634,N_3177);
nand U5720 (N_5720,N_3401,N_3722);
nor U5721 (N_5721,N_3853,N_3328);
nor U5722 (N_5722,N_3511,N_3937);
nand U5723 (N_5723,N_3313,N_3478);
or U5724 (N_5724,N_2563,N_2352);
xor U5725 (N_5725,N_2672,N_2021);
or U5726 (N_5726,N_3910,N_3952);
and U5727 (N_5727,N_2080,N_3784);
or U5728 (N_5728,N_2945,N_3253);
nand U5729 (N_5729,N_3137,N_2390);
xor U5730 (N_5730,N_2716,N_2762);
and U5731 (N_5731,N_3329,N_2541);
nor U5732 (N_5732,N_3407,N_3864);
nor U5733 (N_5733,N_2991,N_3133);
nor U5734 (N_5734,N_3818,N_3428);
xnor U5735 (N_5735,N_2850,N_2313);
nand U5736 (N_5736,N_2867,N_3476);
and U5737 (N_5737,N_2652,N_2998);
or U5738 (N_5738,N_3917,N_2096);
nand U5739 (N_5739,N_3879,N_3147);
nor U5740 (N_5740,N_3471,N_2529);
xnor U5741 (N_5741,N_3298,N_3398);
and U5742 (N_5742,N_2479,N_2113);
or U5743 (N_5743,N_2738,N_3809);
or U5744 (N_5744,N_2279,N_3685);
xnor U5745 (N_5745,N_3446,N_2736);
or U5746 (N_5746,N_2175,N_3323);
or U5747 (N_5747,N_2241,N_2296);
or U5748 (N_5748,N_3134,N_3960);
nand U5749 (N_5749,N_3249,N_2288);
nor U5750 (N_5750,N_3989,N_2193);
nor U5751 (N_5751,N_3657,N_3173);
or U5752 (N_5752,N_2723,N_3468);
nor U5753 (N_5753,N_3266,N_2900);
or U5754 (N_5754,N_2432,N_3360);
and U5755 (N_5755,N_2829,N_3004);
or U5756 (N_5756,N_3571,N_3377);
or U5757 (N_5757,N_2038,N_3406);
or U5758 (N_5758,N_2368,N_2621);
and U5759 (N_5759,N_2185,N_2394);
xor U5760 (N_5760,N_3618,N_3774);
nand U5761 (N_5761,N_2248,N_3647);
and U5762 (N_5762,N_3723,N_2689);
nand U5763 (N_5763,N_2410,N_2794);
or U5764 (N_5764,N_3346,N_3655);
xor U5765 (N_5765,N_3424,N_2430);
or U5766 (N_5766,N_2974,N_3033);
and U5767 (N_5767,N_3859,N_3916);
nor U5768 (N_5768,N_3757,N_2316);
xor U5769 (N_5769,N_2783,N_3289);
and U5770 (N_5770,N_2297,N_3962);
nand U5771 (N_5771,N_2139,N_2588);
xnor U5772 (N_5772,N_3711,N_3256);
nand U5773 (N_5773,N_3023,N_2581);
nand U5774 (N_5774,N_3396,N_2553);
xor U5775 (N_5775,N_2814,N_2308);
xor U5776 (N_5776,N_2145,N_3181);
nand U5777 (N_5777,N_2040,N_2050);
and U5778 (N_5778,N_3014,N_2941);
nand U5779 (N_5779,N_3522,N_2894);
and U5780 (N_5780,N_3365,N_2940);
or U5781 (N_5781,N_2743,N_2796);
nor U5782 (N_5782,N_2556,N_3795);
nand U5783 (N_5783,N_2851,N_2214);
nand U5784 (N_5784,N_3661,N_3581);
or U5785 (N_5785,N_3446,N_2230);
nand U5786 (N_5786,N_2430,N_2933);
xnor U5787 (N_5787,N_2165,N_3799);
nor U5788 (N_5788,N_2744,N_2817);
and U5789 (N_5789,N_3473,N_2220);
xnor U5790 (N_5790,N_3570,N_3120);
or U5791 (N_5791,N_2636,N_3584);
nor U5792 (N_5792,N_2556,N_2048);
nor U5793 (N_5793,N_3407,N_3609);
nor U5794 (N_5794,N_2809,N_2968);
and U5795 (N_5795,N_2210,N_3076);
and U5796 (N_5796,N_3262,N_2403);
xor U5797 (N_5797,N_3051,N_2918);
and U5798 (N_5798,N_2700,N_3336);
nor U5799 (N_5799,N_3146,N_3847);
xnor U5800 (N_5800,N_3936,N_2951);
nor U5801 (N_5801,N_3364,N_2582);
xor U5802 (N_5802,N_2037,N_2348);
nor U5803 (N_5803,N_3794,N_3434);
and U5804 (N_5804,N_3667,N_2960);
nor U5805 (N_5805,N_2172,N_2896);
xor U5806 (N_5806,N_2121,N_3475);
nand U5807 (N_5807,N_2404,N_3069);
nand U5808 (N_5808,N_3888,N_2703);
nor U5809 (N_5809,N_3099,N_2803);
nand U5810 (N_5810,N_2582,N_2636);
xnor U5811 (N_5811,N_3345,N_2991);
nor U5812 (N_5812,N_3819,N_3522);
nand U5813 (N_5813,N_2988,N_3537);
xor U5814 (N_5814,N_3430,N_2570);
or U5815 (N_5815,N_3838,N_3065);
and U5816 (N_5816,N_2708,N_2931);
nor U5817 (N_5817,N_2215,N_2766);
nor U5818 (N_5818,N_3109,N_2181);
and U5819 (N_5819,N_2302,N_2919);
nor U5820 (N_5820,N_2832,N_2544);
nor U5821 (N_5821,N_2458,N_3831);
or U5822 (N_5822,N_2804,N_3576);
and U5823 (N_5823,N_2931,N_2337);
xor U5824 (N_5824,N_2631,N_2732);
xor U5825 (N_5825,N_2594,N_3065);
nor U5826 (N_5826,N_3785,N_3642);
nand U5827 (N_5827,N_3761,N_3191);
nor U5828 (N_5828,N_3662,N_2760);
nor U5829 (N_5829,N_3092,N_3018);
xor U5830 (N_5830,N_3175,N_2162);
or U5831 (N_5831,N_3792,N_3577);
xnor U5832 (N_5832,N_3242,N_2465);
xnor U5833 (N_5833,N_3707,N_3437);
and U5834 (N_5834,N_3636,N_2620);
nand U5835 (N_5835,N_3073,N_2521);
xor U5836 (N_5836,N_2805,N_2807);
and U5837 (N_5837,N_3534,N_3262);
xnor U5838 (N_5838,N_2554,N_2414);
nand U5839 (N_5839,N_3465,N_2625);
xnor U5840 (N_5840,N_2672,N_2050);
xnor U5841 (N_5841,N_2368,N_2289);
or U5842 (N_5842,N_2018,N_2668);
or U5843 (N_5843,N_2431,N_3600);
nand U5844 (N_5844,N_2536,N_3494);
or U5845 (N_5845,N_2792,N_3952);
xnor U5846 (N_5846,N_3653,N_3656);
or U5847 (N_5847,N_2983,N_3887);
nor U5848 (N_5848,N_2040,N_3545);
xnor U5849 (N_5849,N_3883,N_3736);
or U5850 (N_5850,N_3652,N_3720);
and U5851 (N_5851,N_2023,N_3653);
nor U5852 (N_5852,N_2824,N_3086);
nand U5853 (N_5853,N_2307,N_3785);
or U5854 (N_5854,N_2040,N_2256);
nand U5855 (N_5855,N_3263,N_3351);
xnor U5856 (N_5856,N_3969,N_3033);
nand U5857 (N_5857,N_2157,N_2099);
and U5858 (N_5858,N_3365,N_3337);
or U5859 (N_5859,N_2435,N_2995);
nor U5860 (N_5860,N_2171,N_2749);
xor U5861 (N_5861,N_2360,N_2197);
xor U5862 (N_5862,N_3961,N_3679);
xnor U5863 (N_5863,N_2570,N_3434);
or U5864 (N_5864,N_3284,N_2329);
nand U5865 (N_5865,N_3546,N_2214);
xnor U5866 (N_5866,N_3527,N_3916);
xor U5867 (N_5867,N_3609,N_3448);
and U5868 (N_5868,N_3501,N_2584);
nand U5869 (N_5869,N_3753,N_3885);
and U5870 (N_5870,N_2300,N_3715);
nand U5871 (N_5871,N_3396,N_2088);
nand U5872 (N_5872,N_3494,N_3976);
nor U5873 (N_5873,N_2449,N_3163);
nor U5874 (N_5874,N_2470,N_2858);
nand U5875 (N_5875,N_2229,N_2398);
or U5876 (N_5876,N_3218,N_3314);
xnor U5877 (N_5877,N_3012,N_3856);
nand U5878 (N_5878,N_2518,N_2166);
nand U5879 (N_5879,N_2573,N_3233);
nand U5880 (N_5880,N_3137,N_3066);
nand U5881 (N_5881,N_2893,N_3697);
xor U5882 (N_5882,N_2276,N_2275);
and U5883 (N_5883,N_2298,N_3478);
nand U5884 (N_5884,N_3732,N_2371);
nor U5885 (N_5885,N_3072,N_3446);
xor U5886 (N_5886,N_2887,N_3101);
nand U5887 (N_5887,N_3734,N_2580);
or U5888 (N_5888,N_3205,N_3907);
xnor U5889 (N_5889,N_2896,N_3820);
nor U5890 (N_5890,N_3560,N_3127);
xnor U5891 (N_5891,N_2361,N_2983);
nand U5892 (N_5892,N_3114,N_2620);
nand U5893 (N_5893,N_3839,N_3558);
nor U5894 (N_5894,N_2952,N_3197);
xor U5895 (N_5895,N_3631,N_3661);
and U5896 (N_5896,N_2559,N_2538);
nor U5897 (N_5897,N_2350,N_3530);
and U5898 (N_5898,N_2203,N_2417);
nor U5899 (N_5899,N_3193,N_2520);
nor U5900 (N_5900,N_3861,N_3205);
nand U5901 (N_5901,N_3902,N_2358);
xor U5902 (N_5902,N_2047,N_3306);
nand U5903 (N_5903,N_2374,N_2686);
nand U5904 (N_5904,N_3871,N_2771);
nor U5905 (N_5905,N_3781,N_3104);
nand U5906 (N_5906,N_2350,N_3562);
nor U5907 (N_5907,N_3396,N_2521);
xor U5908 (N_5908,N_2635,N_2073);
nand U5909 (N_5909,N_2830,N_2808);
xor U5910 (N_5910,N_3394,N_3279);
nor U5911 (N_5911,N_3408,N_3564);
xnor U5912 (N_5912,N_3208,N_3601);
xor U5913 (N_5913,N_3435,N_3959);
xnor U5914 (N_5914,N_2761,N_2945);
nand U5915 (N_5915,N_2404,N_2304);
nand U5916 (N_5916,N_2623,N_2706);
xnor U5917 (N_5917,N_2686,N_2630);
nor U5918 (N_5918,N_2315,N_3014);
and U5919 (N_5919,N_3152,N_3818);
xnor U5920 (N_5920,N_3549,N_2958);
nand U5921 (N_5921,N_3585,N_2597);
xor U5922 (N_5922,N_2136,N_3821);
nand U5923 (N_5923,N_2708,N_3667);
nand U5924 (N_5924,N_2011,N_3925);
nand U5925 (N_5925,N_3798,N_2373);
or U5926 (N_5926,N_2335,N_2671);
nor U5927 (N_5927,N_3680,N_2943);
or U5928 (N_5928,N_2687,N_2248);
or U5929 (N_5929,N_2757,N_2717);
nand U5930 (N_5930,N_2021,N_3341);
or U5931 (N_5931,N_3511,N_3790);
xor U5932 (N_5932,N_2563,N_3495);
nor U5933 (N_5933,N_3864,N_3345);
nand U5934 (N_5934,N_2394,N_2054);
nor U5935 (N_5935,N_3193,N_3194);
xnor U5936 (N_5936,N_2697,N_2068);
or U5937 (N_5937,N_3125,N_3887);
or U5938 (N_5938,N_3648,N_3662);
nor U5939 (N_5939,N_3338,N_3023);
nand U5940 (N_5940,N_3827,N_3910);
nor U5941 (N_5941,N_3572,N_3632);
nand U5942 (N_5942,N_3417,N_2504);
xor U5943 (N_5943,N_3161,N_3778);
nor U5944 (N_5944,N_3699,N_3392);
nor U5945 (N_5945,N_3926,N_3652);
xor U5946 (N_5946,N_3650,N_2070);
or U5947 (N_5947,N_3198,N_2973);
xor U5948 (N_5948,N_2642,N_2909);
or U5949 (N_5949,N_3897,N_2083);
nand U5950 (N_5950,N_3263,N_2649);
nor U5951 (N_5951,N_2542,N_3460);
nor U5952 (N_5952,N_2043,N_2924);
or U5953 (N_5953,N_2923,N_3330);
nand U5954 (N_5954,N_2313,N_2679);
xor U5955 (N_5955,N_2956,N_2381);
xor U5956 (N_5956,N_2188,N_3714);
xnor U5957 (N_5957,N_2400,N_3154);
or U5958 (N_5958,N_3459,N_2257);
nor U5959 (N_5959,N_2199,N_3931);
xor U5960 (N_5960,N_2931,N_3568);
and U5961 (N_5961,N_2587,N_3240);
and U5962 (N_5962,N_3296,N_2405);
and U5963 (N_5963,N_3493,N_3005);
nor U5964 (N_5964,N_3419,N_3934);
nor U5965 (N_5965,N_3189,N_2303);
nand U5966 (N_5966,N_3685,N_2984);
nand U5967 (N_5967,N_2031,N_2956);
and U5968 (N_5968,N_3883,N_2567);
and U5969 (N_5969,N_2031,N_2544);
nand U5970 (N_5970,N_3495,N_3788);
nor U5971 (N_5971,N_2512,N_2830);
nor U5972 (N_5972,N_2724,N_2858);
and U5973 (N_5973,N_3475,N_3886);
and U5974 (N_5974,N_2453,N_3112);
nand U5975 (N_5975,N_2628,N_3306);
nor U5976 (N_5976,N_3102,N_3468);
nor U5977 (N_5977,N_2586,N_3674);
nand U5978 (N_5978,N_3508,N_2216);
xor U5979 (N_5979,N_3154,N_2428);
nor U5980 (N_5980,N_3975,N_3723);
and U5981 (N_5981,N_2968,N_2233);
and U5982 (N_5982,N_3423,N_3144);
xor U5983 (N_5983,N_3384,N_2234);
nor U5984 (N_5984,N_3919,N_3256);
and U5985 (N_5985,N_2918,N_2239);
nor U5986 (N_5986,N_3382,N_3278);
nand U5987 (N_5987,N_2730,N_3990);
nand U5988 (N_5988,N_3559,N_2819);
nand U5989 (N_5989,N_2301,N_2073);
nand U5990 (N_5990,N_2726,N_2193);
or U5991 (N_5991,N_2162,N_3968);
nand U5992 (N_5992,N_2475,N_3518);
nor U5993 (N_5993,N_3449,N_2461);
nand U5994 (N_5994,N_2818,N_2404);
or U5995 (N_5995,N_3777,N_3270);
nand U5996 (N_5996,N_2150,N_2951);
and U5997 (N_5997,N_2763,N_3649);
or U5998 (N_5998,N_3094,N_3359);
xor U5999 (N_5999,N_2552,N_2963);
and U6000 (N_6000,N_5094,N_5436);
nor U6001 (N_6001,N_5832,N_4160);
xnor U6002 (N_6002,N_4737,N_5230);
nor U6003 (N_6003,N_4570,N_4510);
and U6004 (N_6004,N_4715,N_5614);
and U6005 (N_6005,N_5948,N_4261);
nor U6006 (N_6006,N_4871,N_4013);
and U6007 (N_6007,N_5619,N_4545);
nor U6008 (N_6008,N_4957,N_5982);
nand U6009 (N_6009,N_5695,N_5186);
xnor U6010 (N_6010,N_4842,N_4472);
nand U6011 (N_6011,N_5689,N_4869);
or U6012 (N_6012,N_4723,N_5262);
or U6013 (N_6013,N_4027,N_5008);
xnor U6014 (N_6014,N_4788,N_5355);
nor U6015 (N_6015,N_5173,N_5768);
nor U6016 (N_6016,N_5212,N_4091);
or U6017 (N_6017,N_5057,N_5681);
and U6018 (N_6018,N_5941,N_5775);
xnor U6019 (N_6019,N_4121,N_4523);
and U6020 (N_6020,N_4868,N_4475);
nor U6021 (N_6021,N_5688,N_5122);
xnor U6022 (N_6022,N_4144,N_4150);
nand U6023 (N_6023,N_5964,N_5333);
nand U6024 (N_6024,N_4700,N_4867);
and U6025 (N_6025,N_4255,N_4011);
nor U6026 (N_6026,N_5923,N_5540);
nor U6027 (N_6027,N_5610,N_4456);
or U6028 (N_6028,N_4736,N_5164);
xor U6029 (N_6029,N_4607,N_5208);
xnor U6030 (N_6030,N_5550,N_4098);
xnor U6031 (N_6031,N_4816,N_5836);
and U6032 (N_6032,N_5332,N_4429);
nand U6033 (N_6033,N_4229,N_5406);
or U6034 (N_6034,N_5274,N_5384);
xnor U6035 (N_6035,N_4647,N_5558);
xor U6036 (N_6036,N_4330,N_4390);
and U6037 (N_6037,N_4014,N_4666);
nand U6038 (N_6038,N_4288,N_5883);
and U6039 (N_6039,N_5142,N_4833);
xor U6040 (N_6040,N_5930,N_5628);
nand U6041 (N_6041,N_5335,N_5416);
and U6042 (N_6042,N_5320,N_4382);
nand U6043 (N_6043,N_5859,N_4830);
nor U6044 (N_6044,N_4460,N_4521);
xnor U6045 (N_6045,N_4032,N_5962);
xor U6046 (N_6046,N_5397,N_4694);
xnor U6047 (N_6047,N_5503,N_4758);
or U6048 (N_6048,N_5507,N_5059);
and U6049 (N_6049,N_4861,N_4777);
nand U6050 (N_6050,N_5828,N_4507);
nor U6051 (N_6051,N_4753,N_4086);
xor U6052 (N_6052,N_4481,N_4944);
or U6053 (N_6053,N_4346,N_5322);
and U6054 (N_6054,N_5519,N_4299);
nor U6055 (N_6055,N_4768,N_4360);
xnor U6056 (N_6056,N_5666,N_4359);
nor U6057 (N_6057,N_4953,N_5724);
nand U6058 (N_6058,N_5065,N_5109);
xnor U6059 (N_6059,N_4034,N_5647);
or U6060 (N_6060,N_5382,N_5917);
or U6061 (N_6061,N_5307,N_4470);
and U6062 (N_6062,N_4015,N_4030);
or U6063 (N_6063,N_4931,N_5099);
nor U6064 (N_6064,N_4985,N_4639);
nand U6065 (N_6065,N_4566,N_5734);
nor U6066 (N_6066,N_4041,N_5310);
and U6067 (N_6067,N_5353,N_5650);
or U6068 (N_6068,N_4722,N_5232);
and U6069 (N_6069,N_5165,N_4688);
nor U6070 (N_6070,N_4162,N_4929);
nand U6071 (N_6071,N_4266,N_4231);
nor U6072 (N_6072,N_4386,N_4284);
nand U6073 (N_6073,N_5601,N_5330);
and U6074 (N_6074,N_5638,N_4571);
xnor U6075 (N_6075,N_5779,N_5717);
and U6076 (N_6076,N_4474,N_5398);
xnor U6077 (N_6077,N_5953,N_4214);
or U6078 (N_6078,N_4449,N_5418);
or U6079 (N_6079,N_4002,N_4614);
nand U6080 (N_6080,N_5076,N_5067);
and U6081 (N_6081,N_4538,N_4010);
nor U6082 (N_6082,N_5357,N_5539);
nor U6083 (N_6083,N_4974,N_5053);
nor U6084 (N_6084,N_4468,N_4232);
nand U6085 (N_6085,N_4036,N_4493);
or U6086 (N_6086,N_5972,N_5872);
nand U6087 (N_6087,N_4218,N_5886);
and U6088 (N_6088,N_4683,N_5969);
nor U6089 (N_6089,N_4908,N_5462);
and U6090 (N_6090,N_4267,N_5482);
nor U6091 (N_6091,N_4824,N_4076);
nand U6092 (N_6092,N_5947,N_5551);
or U6093 (N_6093,N_4279,N_5248);
nor U6094 (N_6094,N_4919,N_5323);
nand U6095 (N_6095,N_4695,N_5119);
nand U6096 (N_6096,N_4463,N_4016);
or U6097 (N_6097,N_4602,N_5521);
nor U6098 (N_6098,N_4977,N_4033);
or U6099 (N_6099,N_5537,N_5765);
nor U6100 (N_6100,N_4565,N_4159);
or U6101 (N_6101,N_5863,N_4529);
xnor U6102 (N_6102,N_4771,N_5377);
xnor U6103 (N_6103,N_4125,N_4000);
and U6104 (N_6104,N_4772,N_4380);
nand U6105 (N_6105,N_4684,N_5280);
or U6106 (N_6106,N_5864,N_4747);
nand U6107 (N_6107,N_5279,N_4615);
nor U6108 (N_6108,N_4769,N_4462);
nand U6109 (N_6109,N_5691,N_4547);
nand U6110 (N_6110,N_4056,N_5706);
nor U6111 (N_6111,N_5895,N_4085);
and U6112 (N_6112,N_4573,N_4340);
or U6113 (N_6113,N_4294,N_4897);
nand U6114 (N_6114,N_4434,N_5233);
nand U6115 (N_6115,N_4689,N_4408);
xor U6116 (N_6116,N_4648,N_4223);
xor U6117 (N_6117,N_5791,N_5876);
xnor U6118 (N_6118,N_5531,N_5755);
or U6119 (N_6119,N_4329,N_5995);
nor U6120 (N_6120,N_4585,N_5254);
and U6121 (N_6121,N_5942,N_4618);
or U6122 (N_6122,N_5081,N_5754);
nor U6123 (N_6123,N_5480,N_5940);
nor U6124 (N_6124,N_5258,N_4438);
nor U6125 (N_6125,N_5799,N_5677);
xor U6126 (N_6126,N_5319,N_5805);
xnor U6127 (N_6127,N_4111,N_5066);
xor U6128 (N_6128,N_4937,N_5225);
nand U6129 (N_6129,N_5336,N_4652);
and U6130 (N_6130,N_5932,N_5401);
xnor U6131 (N_6131,N_4735,N_4038);
nor U6132 (N_6132,N_4691,N_4870);
or U6133 (N_6133,N_5998,N_4292);
or U6134 (N_6134,N_4854,N_5074);
nor U6135 (N_6135,N_4844,N_5556);
or U6136 (N_6136,N_4981,N_4806);
and U6137 (N_6137,N_5904,N_5635);
nor U6138 (N_6138,N_4675,N_4290);
or U6139 (N_6139,N_4809,N_4427);
or U6140 (N_6140,N_4793,N_4979);
or U6141 (N_6141,N_4881,N_4677);
and U6142 (N_6142,N_5420,N_4503);
or U6143 (N_6143,N_5375,N_4135);
nand U6144 (N_6144,N_4417,N_4062);
or U6145 (N_6145,N_4943,N_5169);
nand U6146 (N_6146,N_4370,N_4555);
and U6147 (N_6147,N_5300,N_4960);
and U6148 (N_6148,N_5349,N_5415);
and U6149 (N_6149,N_5644,N_4444);
nor U6150 (N_6150,N_5376,N_5546);
xor U6151 (N_6151,N_5427,N_5634);
nor U6152 (N_6152,N_4348,N_4423);
xor U6153 (N_6153,N_4966,N_5529);
or U6154 (N_6154,N_5712,N_4309);
xnor U6155 (N_6155,N_4012,N_5729);
and U6156 (N_6156,N_5661,N_5182);
nor U6157 (N_6157,N_5633,N_5704);
nand U6158 (N_6158,N_5602,N_5277);
nor U6159 (N_6159,N_4933,N_4873);
xnor U6160 (N_6160,N_5034,N_4625);
nor U6161 (N_6161,N_4197,N_4581);
xnor U6162 (N_6162,N_4513,N_5018);
and U6163 (N_6163,N_4781,N_4362);
or U6164 (N_6164,N_4709,N_5532);
xor U6165 (N_6165,N_5292,N_5272);
nand U6166 (N_6166,N_4894,N_4195);
or U6167 (N_6167,N_4318,N_4258);
and U6168 (N_6168,N_5874,N_5564);
nor U6169 (N_6169,N_4609,N_5815);
and U6170 (N_6170,N_5501,N_4484);
and U6171 (N_6171,N_4303,N_4754);
nand U6172 (N_6172,N_5327,N_4895);
nor U6173 (N_6173,N_4839,N_5266);
nor U6174 (N_6174,N_5334,N_4925);
and U6175 (N_6175,N_4997,N_5616);
nand U6176 (N_6176,N_4989,N_5234);
and U6177 (N_6177,N_4164,N_4240);
xnor U6178 (N_6178,N_5231,N_4316);
nand U6179 (N_6179,N_5425,N_5496);
nand U6180 (N_6180,N_5920,N_4070);
nand U6181 (N_6181,N_5002,N_5147);
nand U6182 (N_6182,N_5188,N_4331);
xor U6183 (N_6183,N_4275,N_4057);
and U6184 (N_6184,N_5820,N_4962);
xnor U6185 (N_6185,N_5346,N_4378);
or U6186 (N_6186,N_5987,N_4584);
or U6187 (N_6187,N_4577,N_4704);
and U6188 (N_6188,N_5983,N_4451);
or U6189 (N_6189,N_4559,N_5649);
or U6190 (N_6190,N_4716,N_4601);
xor U6191 (N_6191,N_5528,N_4950);
or U6192 (N_6192,N_5646,N_5851);
nor U6193 (N_6193,N_5299,N_4958);
or U6194 (N_6194,N_5429,N_5235);
or U6195 (N_6195,N_4471,N_4674);
xnor U6196 (N_6196,N_4798,N_5510);
nor U6197 (N_6197,N_4619,N_5451);
nand U6198 (N_6198,N_5329,N_4520);
and U6199 (N_6199,N_4439,N_5502);
or U6200 (N_6200,N_4221,N_5338);
nand U6201 (N_6201,N_4794,N_4101);
xnor U6202 (N_6202,N_4909,N_5887);
nor U6203 (N_6203,N_4608,N_5146);
and U6204 (N_6204,N_5985,N_4549);
nor U6205 (N_6205,N_5005,N_4915);
nand U6206 (N_6206,N_5727,N_4600);
xor U6207 (N_6207,N_4393,N_4560);
and U6208 (N_6208,N_4367,N_5504);
nand U6209 (N_6209,N_5197,N_4668);
nand U6210 (N_6210,N_4813,N_5888);
xor U6211 (N_6211,N_4385,N_5063);
nor U6212 (N_6212,N_4643,N_5276);
nand U6213 (N_6213,N_5780,N_5404);
nand U6214 (N_6214,N_4739,N_5555);
or U6215 (N_6215,N_5508,N_5162);
and U6216 (N_6216,N_4308,N_5183);
nor U6217 (N_6217,N_4506,N_4230);
xnor U6218 (N_6218,N_4219,N_5560);
nand U6219 (N_6219,N_4638,N_5424);
nand U6220 (N_6220,N_5512,N_4285);
or U6221 (N_6221,N_5345,N_5544);
xor U6222 (N_6222,N_5221,N_5267);
or U6223 (N_6223,N_4969,N_4263);
and U6224 (N_6224,N_5044,N_5839);
and U6225 (N_6225,N_4156,N_5494);
or U6226 (N_6226,N_5946,N_4744);
and U6227 (N_6227,N_4354,N_5670);
nor U6228 (N_6228,N_4073,N_5513);
and U6229 (N_6229,N_5976,N_5924);
or U6230 (N_6230,N_5545,N_5070);
or U6231 (N_6231,N_4431,N_5667);
xor U6232 (N_6232,N_5001,N_5159);
xnor U6233 (N_6233,N_5093,N_5553);
nor U6234 (N_6234,N_5731,N_5500);
nand U6235 (N_6235,N_5552,N_4366);
and U6236 (N_6236,N_4687,N_5662);
nand U6237 (N_6237,N_5816,N_4406);
and U6238 (N_6238,N_4020,N_4572);
or U6239 (N_6239,N_4847,N_5652);
nor U6240 (N_6240,N_4727,N_5367);
nor U6241 (N_6241,N_4698,N_5868);
nor U6242 (N_6242,N_4200,N_4405);
xor U6243 (N_6243,N_4826,N_5936);
or U6244 (N_6244,N_4259,N_5723);
or U6245 (N_6245,N_4106,N_4514);
or U6246 (N_6246,N_4412,N_4669);
nor U6247 (N_6247,N_4097,N_4814);
nand U6248 (N_6248,N_5378,N_4662);
nand U6249 (N_6249,N_4055,N_5852);
xor U6250 (N_6250,N_4006,N_4483);
nor U6251 (N_6251,N_5682,N_4530);
xnor U6252 (N_6252,N_4300,N_5933);
xnor U6253 (N_6253,N_5243,N_4850);
or U6254 (N_6254,N_4488,N_5938);
and U6255 (N_6255,N_4629,N_4673);
and U6256 (N_6256,N_4084,N_4174);
xnor U6257 (N_6257,N_4594,N_4682);
and U6258 (N_6258,N_5153,N_5675);
nor U6259 (N_6259,N_5697,N_5132);
and U6260 (N_6260,N_5928,N_4029);
nor U6261 (N_6261,N_5037,N_5641);
and U6262 (N_6262,N_5862,N_4732);
nor U6263 (N_6263,N_4022,N_4880);
and U6264 (N_6264,N_5447,N_4372);
and U6265 (N_6265,N_4835,N_5577);
nor U6266 (N_6266,N_4227,N_5793);
nand U6267 (N_6267,N_5111,N_5477);
nand U6268 (N_6268,N_4409,N_4719);
or U6269 (N_6269,N_4587,N_4323);
and U6270 (N_6270,N_4315,N_4075);
nor U6271 (N_6271,N_4001,N_4552);
or U6272 (N_6272,N_4211,N_5522);
and U6273 (N_6273,N_5700,N_4112);
nor U6274 (N_6274,N_4857,N_4155);
nand U6275 (N_6275,N_4243,N_4117);
and U6276 (N_6276,N_4454,N_5584);
nand U6277 (N_6277,N_4993,N_4636);
and U6278 (N_6278,N_5549,N_4654);
and U6279 (N_6279,N_4916,N_5204);
nor U6280 (N_6280,N_4305,N_5390);
nor U6281 (N_6281,N_5051,N_4199);
and U6282 (N_6282,N_5802,N_5955);
xor U6283 (N_6283,N_4216,N_5830);
nor U6284 (N_6284,N_5726,N_5324);
nand U6285 (N_6285,N_4491,N_4047);
and U6286 (N_6286,N_4147,N_4217);
xor U6287 (N_6287,N_4238,N_4762);
and U6288 (N_6288,N_4283,N_4186);
nand U6289 (N_6289,N_5224,N_5640);
or U6290 (N_6290,N_5632,N_5219);
or U6291 (N_6291,N_5304,N_5170);
nor U6292 (N_6292,N_4890,N_5321);
and U6293 (N_6293,N_4310,N_5603);
xnor U6294 (N_6294,N_4208,N_4495);
xor U6295 (N_6295,N_5855,N_4942);
or U6296 (N_6296,N_4326,N_4096);
or U6297 (N_6297,N_5607,N_5210);
nand U6298 (N_6298,N_4436,N_5489);
or U6299 (N_6299,N_4987,N_4465);
xor U6300 (N_6300,N_5259,N_4836);
nor U6301 (N_6301,N_5898,N_4918);
and U6302 (N_6302,N_4063,N_4332);
or U6303 (N_6303,N_5363,N_4141);
nand U6304 (N_6304,N_5903,N_5128);
nor U6305 (N_6305,N_4963,N_4902);
nor U6306 (N_6306,N_4784,N_4834);
and U6307 (N_6307,N_5297,N_4361);
xor U6308 (N_6308,N_5368,N_4265);
and U6309 (N_6309,N_4742,N_4729);
nor U6310 (N_6310,N_5387,N_5934);
or U6311 (N_6311,N_4100,N_5288);
and U6312 (N_6312,N_4224,N_5800);
xor U6313 (N_6313,N_5708,N_4637);
nor U6314 (N_6314,N_5270,N_5386);
nor U6315 (N_6315,N_4856,N_4557);
xor U6316 (N_6316,N_4035,N_5639);
and U6317 (N_6317,N_4166,N_4140);
nand U6318 (N_6318,N_5604,N_4368);
xor U6319 (N_6319,N_5705,N_5314);
nand U6320 (N_6320,N_4975,N_5589);
nor U6321 (N_6321,N_5988,N_4593);
xor U6322 (N_6322,N_5752,N_4352);
or U6323 (N_6323,N_5140,N_5020);
nor U6324 (N_6324,N_4228,N_4109);
nand U6325 (N_6325,N_4801,N_4982);
and U6326 (N_6326,N_4277,N_5956);
nand U6327 (N_6327,N_5557,N_5264);
and U6328 (N_6328,N_5719,N_4537);
nor U6329 (N_6329,N_5035,N_4752);
xnor U6330 (N_6330,N_5295,N_5108);
xor U6331 (N_6331,N_4865,N_4247);
and U6332 (N_6332,N_5472,N_5658);
or U6333 (N_6333,N_4328,N_5915);
or U6334 (N_6334,N_4779,N_4885);
and U6335 (N_6335,N_5905,N_5468);
xor U6336 (N_6336,N_4980,N_4226);
and U6337 (N_6337,N_4442,N_5252);
xor U6338 (N_6338,N_5757,N_4952);
nor U6339 (N_6339,N_5913,N_4680);
xnor U6340 (N_6340,N_4517,N_5251);
or U6341 (N_6341,N_5442,N_4357);
and U6342 (N_6342,N_4212,N_5478);
nand U6343 (N_6343,N_5331,N_4251);
nand U6344 (N_6344,N_5736,N_4270);
and U6345 (N_6345,N_5075,N_4911);
and U6346 (N_6346,N_5511,N_4432);
nand U6347 (N_6347,N_5725,N_5306);
nand U6348 (N_6348,N_5016,N_5694);
nor U6349 (N_6349,N_5533,N_4973);
nand U6350 (N_6350,N_4042,N_5202);
and U6351 (N_6351,N_4148,N_5696);
and U6352 (N_6352,N_5509,N_4198);
xor U6353 (N_6353,N_4910,N_4089);
nand U6354 (N_6354,N_4878,N_5654);
nand U6355 (N_6355,N_5271,N_4416);
nor U6356 (N_6356,N_4302,N_5908);
and U6357 (N_6357,N_5894,N_5643);
and U6358 (N_6358,N_4664,N_5834);
nand U6359 (N_6359,N_4518,N_4397);
and U6360 (N_6360,N_5699,N_4934);
nand U6361 (N_6361,N_4921,N_5303);
or U6362 (N_6362,N_5817,N_5713);
and U6363 (N_6363,N_5179,N_4964);
nand U6364 (N_6364,N_5396,N_5124);
xor U6365 (N_6365,N_5139,N_5975);
and U6366 (N_6366,N_4782,N_4525);
xnor U6367 (N_6367,N_5150,N_5721);
and U6368 (N_6368,N_5444,N_5841);
nor U6369 (N_6369,N_4939,N_4787);
and U6370 (N_6370,N_4296,N_4268);
or U6371 (N_6371,N_4457,N_4443);
xor U6372 (N_6372,N_5580,N_4676);
nor U6373 (N_6373,N_5530,N_4641);
xor U6374 (N_6374,N_5163,N_4774);
and U6375 (N_6375,N_4114,N_5152);
nor U6376 (N_6376,N_4505,N_4235);
xnor U6377 (N_6377,N_4196,N_4971);
nor U6378 (N_6378,N_4522,N_5958);
nor U6379 (N_6379,N_5045,N_4635);
nand U6380 (N_6380,N_4564,N_5901);
xnor U6381 (N_6381,N_5538,N_5223);
nor U6382 (N_6382,N_4215,N_5655);
and U6383 (N_6383,N_4134,N_5753);
or U6384 (N_6384,N_4879,N_4343);
or U6385 (N_6385,N_4129,N_4995);
and U6386 (N_6386,N_5980,N_4575);
nor U6387 (N_6387,N_5965,N_5608);
and U6388 (N_6388,N_4800,N_5850);
nand U6389 (N_6389,N_5842,N_4171);
xnor U6390 (N_6390,N_4342,N_4253);
nor U6391 (N_6391,N_4394,N_4967);
xnor U6392 (N_6392,N_4213,N_5474);
nor U6393 (N_6393,N_4461,N_4225);
nand U6394 (N_6394,N_5029,N_5428);
nand U6395 (N_6395,N_4656,N_4621);
nand U6396 (N_6396,N_4623,N_5824);
nor U6397 (N_6397,N_5648,N_4546);
and U6398 (N_6398,N_4353,N_5337);
or U6399 (N_6399,N_5592,N_5144);
nor U6400 (N_6400,N_5026,N_5437);
or U6401 (N_6401,N_4074,N_4170);
xor U6402 (N_6402,N_4886,N_5056);
xor U6403 (N_6403,N_5772,N_5285);
nor U6404 (N_6404,N_4061,N_5636);
nand U6405 (N_6405,N_5090,N_4976);
nand U6406 (N_6406,N_4720,N_4025);
nand U6407 (N_6407,N_4877,N_5910);
or U6408 (N_6408,N_4912,N_4616);
xor U6409 (N_6409,N_5205,N_4401);
and U6410 (N_6410,N_4756,N_4080);
or U6411 (N_6411,N_5354,N_4802);
or U6412 (N_6412,N_5215,N_4092);
nor U6413 (N_6413,N_4951,N_5242);
xnor U6414 (N_6414,N_5989,N_5679);
nor U6415 (N_6415,N_5819,N_5372);
nand U6416 (N_6416,N_4613,N_5916);
or U6417 (N_6417,N_5740,N_4708);
nor U6418 (N_6418,N_4103,N_4748);
and U6419 (N_6419,N_4078,N_4207);
and U6420 (N_6420,N_4863,N_4578);
nor U6421 (N_6421,N_4740,N_5228);
nand U6422 (N_6422,N_5893,N_5684);
and U6423 (N_6423,N_5061,N_5176);
xnor U6424 (N_6424,N_5878,N_5244);
nor U6425 (N_6425,N_4469,N_4822);
xnor U6426 (N_6426,N_5929,N_5195);
or U6427 (N_6427,N_5036,N_4105);
or U6428 (N_6428,N_5977,N_4496);
or U6429 (N_6429,N_5364,N_4743);
xor U6430 (N_6430,N_5356,N_5663);
or U6431 (N_6431,N_5410,N_5825);
nand U6432 (N_6432,N_5077,N_5973);
and U6433 (N_6433,N_4059,N_4838);
nor U6434 (N_6434,N_5073,N_5118);
xor U6435 (N_6435,N_4968,N_4428);
xor U6436 (N_6436,N_5268,N_4095);
nor U6437 (N_6437,N_5750,N_5698);
xnor U6438 (N_6438,N_4502,N_5344);
nor U6439 (N_6439,N_4580,N_5884);
nand U6440 (N_6440,N_4999,N_4701);
xor U6441 (N_6441,N_4563,N_4749);
xor U6442 (N_6442,N_5203,N_4524);
and U6443 (N_6443,N_4163,N_5823);
nor U6444 (N_6444,N_4930,N_5194);
nand U6445 (N_6445,N_5782,N_4811);
nor U6446 (N_6446,N_4418,N_5629);
nand U6447 (N_6447,N_5043,N_5253);
nand U6448 (N_6448,N_5595,N_4203);
nor U6449 (N_6449,N_4770,N_4551);
nor U6450 (N_6450,N_5459,N_5441);
nor U6451 (N_6451,N_4866,N_5918);
nor U6452 (N_6452,N_5542,N_4606);
xnor U6453 (N_6453,N_5520,N_4710);
xnor U6454 (N_6454,N_5787,N_5412);
xnor U6455 (N_6455,N_4480,N_5213);
nand U6456 (N_6456,N_5766,N_4333);
xor U6457 (N_6457,N_5426,N_4853);
nand U6458 (N_6458,N_4146,N_5283);
xor U6459 (N_6459,N_5984,N_5058);
nand U6460 (N_6460,N_5891,N_5088);
nand U6461 (N_6461,N_4825,N_5587);
or U6462 (N_6462,N_4685,N_4446);
nand U6463 (N_6463,N_5978,N_4659);
or U6464 (N_6464,N_4274,N_4287);
nor U6465 (N_6465,N_4077,N_5255);
and U6466 (N_6466,N_5720,N_5269);
xor U6467 (N_6467,N_4961,N_5590);
or U6468 (N_6468,N_4313,N_4037);
nand U6469 (N_6469,N_5784,N_4874);
or U6470 (N_6470,N_4696,N_4193);
xor U6471 (N_6471,N_5952,N_5112);
nand U6472 (N_6472,N_4202,N_4139);
nor U6473 (N_6473,N_5767,N_4778);
nand U6474 (N_6474,N_5104,N_4317);
nor U6475 (N_6475,N_5814,N_4242);
or U6476 (N_6476,N_5072,N_4478);
and U6477 (N_6477,N_4048,N_5421);
nand U6478 (N_6478,N_4433,N_4067);
nor U6479 (N_6479,N_5417,N_4116);
and U6480 (N_6480,N_4031,N_5609);
and U6481 (N_6481,N_4812,N_4005);
nand U6482 (N_6482,N_4900,N_4728);
xor U6483 (N_6483,N_5102,N_5548);
nor U6484 (N_6484,N_5499,N_4426);
nor U6485 (N_6485,N_4239,N_4090);
nand U6486 (N_6486,N_5714,N_5380);
nand U6487 (N_6487,N_5914,N_4624);
and U6488 (N_6488,N_4837,N_4731);
nor U6489 (N_6489,N_5284,N_4590);
nand U6490 (N_6490,N_4887,N_5950);
nor U6491 (N_6491,N_5971,N_5711);
xor U6492 (N_6492,N_5460,N_5935);
and U6493 (N_6493,N_5856,N_4419);
nor U6494 (N_6494,N_5265,N_4786);
nor U6495 (N_6495,N_5113,N_5240);
nor U6496 (N_6496,N_4248,N_5209);
xor U6497 (N_6497,N_5087,N_5857);
nand U6498 (N_6498,N_4998,N_5732);
nand U6499 (N_6499,N_5457,N_4371);
and U6500 (N_6500,N_5844,N_5690);
or U6501 (N_6501,N_4548,N_5671);
xor U6502 (N_6502,N_5031,N_4791);
or U6503 (N_6503,N_5214,N_4425);
nor U6504 (N_6504,N_4322,N_4028);
or U6505 (N_6505,N_5797,N_5136);
nor U6506 (N_6506,N_5615,N_5000);
nand U6507 (N_6507,N_5086,N_5525);
or U6508 (N_6508,N_4860,N_5833);
and U6509 (N_6509,N_4745,N_5217);
xor U6510 (N_6510,N_4633,N_4190);
and U6511 (N_6511,N_4003,N_5536);
nand U6512 (N_6512,N_4707,N_4252);
or U6513 (N_6513,N_5445,N_4447);
and U6514 (N_6514,N_5116,N_5569);
and U6515 (N_6515,N_4249,N_4663);
xnor U6516 (N_6516,N_5049,N_4905);
and U6517 (N_6517,N_4051,N_4927);
nor U6518 (N_6518,N_5506,N_5858);
xor U6519 (N_6519,N_5096,N_5229);
nand U6520 (N_6520,N_5909,N_5190);
nand U6521 (N_6521,N_4402,N_5350);
and U6522 (N_6522,N_4516,N_4917);
or U6523 (N_6523,N_5911,N_4640);
and U6524 (N_6524,N_5715,N_4714);
and U6525 (N_6525,N_4759,N_4901);
or U6526 (N_6526,N_5207,N_4388);
nor U6527 (N_6527,N_4645,N_4320);
and U6528 (N_6528,N_4490,N_4938);
or U6529 (N_6529,N_5341,N_4173);
or U6530 (N_6530,N_4374,N_4489);
and U6531 (N_6531,N_4576,N_4986);
nor U6532 (N_6532,N_4650,N_4829);
nor U6533 (N_6533,N_4533,N_5452);
nor U6534 (N_6534,N_4932,N_4542);
or U6535 (N_6535,N_4876,N_5089);
and U6536 (N_6536,N_5741,N_5879);
nor U6537 (N_6537,N_4941,N_5673);
nor U6538 (N_6538,N_4053,N_4702);
or U6539 (N_6539,N_4424,N_4903);
and U6540 (N_6540,N_4237,N_5826);
xor U6541 (N_6541,N_4697,N_5737);
xnor U6542 (N_6542,N_4693,N_4773);
xor U6543 (N_6543,N_5747,N_5517);
or U6544 (N_6544,N_5758,N_5004);
nor U6545 (N_6545,N_4004,N_5483);
nor U6546 (N_6546,N_5172,N_4792);
xnor U6547 (N_6547,N_5585,N_4143);
and U6548 (N_6548,N_5716,N_4068);
or U6549 (N_6549,N_4177,N_5885);
nand U6550 (N_6550,N_4415,N_5620);
or U6551 (N_6551,N_5311,N_4928);
and U6552 (N_6552,N_5762,N_5669);
and U6553 (N_6553,N_5598,N_4864);
or U6554 (N_6554,N_5015,N_4381);
nand U6555 (N_6555,N_4690,N_4622);
nor U6556 (N_6556,N_4087,N_5399);
or U6557 (N_6557,N_5430,N_4334);
nand U6558 (N_6558,N_5794,N_4845);
or U6559 (N_6559,N_4898,N_5582);
or U6560 (N_6560,N_5524,N_4169);
xnor U6561 (N_6561,N_4120,N_4420);
nand U6562 (N_6562,N_4404,N_4515);
or U6563 (N_6563,N_5490,N_5157);
or U6564 (N_6564,N_5906,N_5481);
nand U6565 (N_6565,N_4459,N_5039);
or U6566 (N_6566,N_4487,N_4083);
xnor U6567 (N_6567,N_5796,N_4464);
or U6568 (N_6568,N_5438,N_5448);
nor U6569 (N_6569,N_4052,N_5294);
or U6570 (N_6570,N_5873,N_4627);
nand U6571 (N_6571,N_5318,N_5155);
nand U6572 (N_6572,N_5064,N_5046);
nand U6573 (N_6573,N_4808,N_5701);
xor U6574 (N_6574,N_5042,N_5931);
or U6575 (N_6575,N_4046,N_5054);
and U6576 (N_6576,N_5686,N_4254);
and U6577 (N_6577,N_4205,N_4192);
xnor U6578 (N_6578,N_5660,N_4498);
and U6579 (N_6579,N_4764,N_5392);
nand U6580 (N_6580,N_5678,N_4717);
nor U6581 (N_6581,N_4597,N_5078);
or U6582 (N_6582,N_5835,N_5352);
nor U6583 (N_6583,N_4008,N_5707);
xor U6584 (N_6584,N_4306,N_4021);
xnor U6585 (N_6585,N_5882,N_5487);
and U6586 (N_6586,N_4775,N_5896);
or U6587 (N_6587,N_4123,N_5298);
or U6588 (N_6588,N_4763,N_4926);
xor U6589 (N_6589,N_4282,N_5110);
nand U6590 (N_6590,N_5591,N_4734);
or U6591 (N_6591,N_4984,N_4554);
nor U6592 (N_6592,N_5994,N_4526);
nor U6593 (N_6593,N_4992,N_5358);
nor U6594 (N_6594,N_4050,N_4325);
and U6595 (N_6595,N_5581,N_5583);
or U6596 (N_6596,N_5154,N_4539);
nand U6597 (N_6597,N_4841,N_5469);
nand U6598 (N_6598,N_4724,N_4154);
and U6599 (N_6599,N_5811,N_5317);
xor U6600 (N_6600,N_4389,N_4586);
xor U6601 (N_6601,N_4532,N_4113);
nor U6602 (N_6602,N_5211,N_4617);
or U6603 (N_6603,N_5803,N_5239);
nand U6604 (N_6604,N_5339,N_5105);
nor U6605 (N_6605,N_5778,N_4188);
nor U6606 (N_6606,N_4907,N_5351);
or U6607 (N_6607,N_5756,N_4181);
xor U6608 (N_6608,N_4776,N_5312);
nand U6609 (N_6609,N_5579,N_4651);
or U6610 (N_6610,N_5818,N_4176);
and U6611 (N_6611,N_5388,N_5129);
xnor U6612 (N_6612,N_5991,N_4145);
nor U6613 (N_6613,N_5846,N_4556);
nor U6614 (N_6614,N_4398,N_4127);
and U6615 (N_6615,N_5222,N_5561);
xor U6616 (N_6616,N_5296,N_4108);
nor U6617 (N_6617,N_4628,N_5305);
nand U6618 (N_6618,N_5455,N_5301);
nor U6619 (N_6619,N_4441,N_5246);
xor U6620 (N_6620,N_5187,N_5505);
or U6621 (N_6621,N_4721,N_4307);
xnor U6622 (N_6622,N_4923,N_4082);
or U6623 (N_6623,N_5742,N_4375);
nor U6624 (N_6624,N_5680,N_5365);
nand U6625 (N_6625,N_4567,N_4713);
nand U6626 (N_6626,N_4588,N_4828);
or U6627 (N_6627,N_5912,N_4272);
nor U6628 (N_6628,N_4094,N_4725);
nor U6629 (N_6629,N_4497,N_4153);
nor U6630 (N_6630,N_4591,N_5925);
and U6631 (N_6631,N_4804,N_4644);
xor U6632 (N_6632,N_4440,N_4805);
and U6633 (N_6633,N_5937,N_5514);
xor U6634 (N_6634,N_4007,N_4437);
xnor U6635 (N_6635,N_5781,N_5759);
nand U6636 (N_6636,N_5189,N_5566);
and U6637 (N_6637,N_5009,N_4209);
nor U6638 (N_6638,N_4273,N_4583);
and U6639 (N_6639,N_4045,N_4589);
and U6640 (N_6640,N_5097,N_4276);
and U6641 (N_6641,N_5907,N_5161);
or U6642 (N_6642,N_5071,N_5570);
xor U6643 (N_6643,N_4298,N_4954);
or U6644 (N_6644,N_5287,N_5423);
nand U6645 (N_6645,N_4665,N_5683);
nor U6646 (N_6646,N_4899,N_4492);
nor U6647 (N_6647,N_4072,N_5196);
or U6648 (N_6648,N_5963,N_5393);
or U6649 (N_6649,N_4946,N_5454);
nand U6650 (N_6650,N_5434,N_4301);
nand U6651 (N_6651,N_5069,N_5014);
and U6652 (N_6652,N_4043,N_5880);
xnor U6653 (N_6653,N_5156,N_5273);
xnor U6654 (N_6654,N_5735,N_5055);
nor U6655 (N_6655,N_5627,N_5534);
or U6656 (N_6656,N_4335,N_5199);
or U6657 (N_6657,N_5178,N_5185);
xnor U6658 (N_6658,N_4054,N_5739);
nand U6659 (N_6659,N_5369,N_4679);
or U6660 (N_6660,N_4349,N_5191);
nand U6661 (N_6661,N_4102,N_5656);
and U6662 (N_6662,N_4796,N_5746);
nor U6663 (N_6663,N_4858,N_4568);
xor U6664 (N_6664,N_4377,N_5138);
or U6665 (N_6665,N_5866,N_5151);
or U6666 (N_6666,N_5038,N_4528);
xnor U6667 (N_6667,N_4922,N_5959);
nor U6668 (N_6668,N_4327,N_5944);
xnor U6669 (N_6669,N_5659,N_4840);
nand U6670 (N_6670,N_4476,N_4194);
or U6671 (N_6671,N_5710,N_5177);
or U6672 (N_6672,N_5807,N_4686);
nor U6673 (N_6673,N_5999,N_5518);
nor U6674 (N_6674,N_5326,N_4264);
nor U6675 (N_6675,N_5484,N_4039);
xor U6676 (N_6676,N_4115,N_4531);
nor U6677 (N_6677,N_5006,N_4363);
nor U6678 (N_6678,N_5422,N_4620);
nand U6679 (N_6679,N_5095,N_5764);
xor U6680 (N_6680,N_4244,N_4599);
and U6681 (N_6681,N_5411,N_4852);
nand U6682 (N_6682,N_4741,N_5922);
and U6683 (N_6683,N_5745,N_5131);
nor U6684 (N_6684,N_4473,N_5275);
or U6685 (N_6685,N_4262,N_4040);
nor U6686 (N_6686,N_5871,N_5491);
and U6687 (N_6687,N_4935,N_4827);
xnor U6688 (N_6688,N_4494,N_5760);
or U6689 (N_6689,N_4295,N_5473);
or U6690 (N_6690,N_5611,N_5565);
or U6691 (N_6691,N_4338,N_4978);
nand U6692 (N_6692,N_4819,N_4391);
and U6693 (N_6693,N_5083,N_5370);
or U6694 (N_6694,N_5193,N_5012);
nor U6695 (N_6695,N_4064,N_4124);
xor U6696 (N_6696,N_5672,N_4184);
or U6697 (N_6697,N_4574,N_5769);
nor U6698 (N_6698,N_4582,N_4182);
nand U6699 (N_6699,N_4803,N_5653);
xor U6700 (N_6700,N_5403,N_5515);
xor U6701 (N_6701,N_5847,N_5927);
nor U6702 (N_6702,N_4807,N_5709);
nand U6703 (N_6703,N_5622,N_4511);
nor U6704 (N_6704,N_5313,N_4324);
nor U6705 (N_6705,N_4185,N_5889);
or U6706 (N_6706,N_5777,N_5167);
xnor U6707 (N_6707,N_5899,N_5106);
or U6708 (N_6708,N_5776,N_4256);
or U6709 (N_6709,N_4630,N_4384);
nand U6710 (N_6710,N_5160,N_4534);
xnor U6711 (N_6711,N_4562,N_4988);
nor U6712 (N_6712,N_5685,N_5703);
and U6713 (N_6713,N_5062,N_5149);
and U6714 (N_6714,N_4107,N_5860);
xnor U6715 (N_6715,N_5048,N_5461);
xnor U6716 (N_6716,N_4940,N_4983);
or U6717 (N_6717,N_5801,N_5371);
xor U6718 (N_6718,N_5361,N_5135);
nor U6719 (N_6719,N_4234,N_4733);
xnor U6720 (N_6720,N_5821,N_5030);
xnor U6721 (N_6721,N_4395,N_5527);
nor U6722 (N_6722,N_5467,N_5578);
nor U6723 (N_6723,N_4445,N_5032);
nor U6724 (N_6724,N_4790,N_4817);
nor U6725 (N_6725,N_4286,N_5789);
or U6726 (N_6726,N_5291,N_5730);
xnor U6727 (N_6727,N_4632,N_5554);
or U6728 (N_6728,N_5881,N_4018);
xnor U6729 (N_6729,N_5822,N_5379);
nor U6730 (N_6730,N_4920,N_5687);
nand U6731 (N_6731,N_5261,N_4947);
nor U6732 (N_6732,N_5806,N_5475);
nor U6733 (N_6733,N_4670,N_4499);
and U6734 (N_6734,N_5413,N_4726);
and U6735 (N_6735,N_5625,N_5786);
nor U6736 (N_6736,N_4751,N_4132);
nor U6737 (N_6737,N_5645,N_4843);
xor U6738 (N_6738,N_4411,N_5409);
nor U6739 (N_6739,N_4757,N_4681);
and U6740 (N_6740,N_4855,N_4509);
nor U6741 (N_6741,N_4746,N_5385);
or U6742 (N_6742,N_4138,N_5443);
nor U6743 (N_6743,N_5668,N_4634);
xor U6744 (N_6744,N_4785,N_4604);
nor U6745 (N_6745,N_5366,N_4157);
and U6746 (N_6746,N_5867,N_5060);
xor U6747 (N_6747,N_5612,N_5464);
xnor U6748 (N_6748,N_5516,N_4889);
xor U6749 (N_6749,N_5079,N_5599);
xnor U6750 (N_6750,N_5892,N_4891);
and U6751 (N_6751,N_5237,N_4172);
nand U6752 (N_6752,N_5693,N_5181);
xnor U6753 (N_6753,N_4904,N_4168);
nor U6754 (N_6754,N_5843,N_5325);
nor U6755 (N_6755,N_4851,N_5440);
xor U6756 (N_6756,N_4356,N_4099);
and U6757 (N_6757,N_5574,N_5115);
xor U6758 (N_6758,N_5951,N_4118);
or U6759 (N_6759,N_5771,N_5100);
nor U6760 (N_6760,N_4718,N_5795);
nand U6761 (N_6761,N_4738,N_5117);
nor U6762 (N_6762,N_5630,N_4278);
nor U6763 (N_6763,N_5875,N_4789);
or U6764 (N_6764,N_4339,N_5328);
xnor U6765 (N_6765,N_5206,N_4712);
or U6766 (N_6766,N_5256,N_5342);
or U6767 (N_6767,N_4820,N_4414);
nor U6768 (N_6768,N_4821,N_5408);
xor U6769 (N_6769,N_5347,N_4241);
and U6770 (N_6770,N_4093,N_5981);
xor U6771 (N_6771,N_4399,N_4996);
nor U6772 (N_6772,N_4760,N_4152);
and U6773 (N_6773,N_5238,N_4527);
nand U6774 (N_6774,N_4705,N_4161);
xor U6775 (N_6775,N_4500,N_4452);
xor U6776 (N_6776,N_4104,N_5919);
and U6777 (N_6777,N_5471,N_4355);
and U6778 (N_6778,N_5068,N_4017);
or U6779 (N_6779,N_5605,N_4610);
or U6780 (N_6780,N_4672,N_4403);
and U6781 (N_6781,N_5028,N_5970);
and U6782 (N_6782,N_4311,N_5626);
xnor U6783 (N_6783,N_4831,N_5141);
nor U6784 (N_6784,N_5383,N_5114);
xor U6785 (N_6785,N_4544,N_5798);
or U6786 (N_6786,N_5022,N_4347);
nor U6787 (N_6787,N_5809,N_5674);
xor U6788 (N_6788,N_5123,N_4959);
xor U6789 (N_6789,N_4896,N_5492);
nand U6790 (N_6790,N_5125,N_5348);
and U6791 (N_6791,N_4605,N_4373);
or U6792 (N_6792,N_5495,N_5362);
xnor U6793 (N_6793,N_5979,N_5853);
xor U6794 (N_6794,N_5617,N_5902);
nor U6795 (N_6795,N_4646,N_4945);
and U6796 (N_6796,N_5535,N_5526);
and U6797 (N_6797,N_4280,N_5389);
nor U6798 (N_6798,N_5192,N_4421);
nor U6799 (N_6799,N_4413,N_5961);
nand U6800 (N_6800,N_5479,N_4026);
xnor U6801 (N_6801,N_4882,N_5174);
xor U6802 (N_6802,N_5047,N_5547);
xnor U6803 (N_6803,N_4955,N_5562);
nand U6804 (N_6804,N_4376,N_4019);
and U6805 (N_6805,N_5642,N_5664);
nand U6806 (N_6806,N_4058,N_5498);
or U6807 (N_6807,N_5017,N_4949);
xor U6808 (N_6808,N_5749,N_5394);
nor U6809 (N_6809,N_5575,N_5175);
nand U6810 (N_6810,N_5568,N_4579);
or U6811 (N_6811,N_5260,N_5761);
nor U6812 (N_6812,N_5957,N_4448);
nor U6813 (N_6813,N_4888,N_5184);
xor U6814 (N_6814,N_5869,N_5281);
and U6815 (N_6815,N_4297,N_5637);
nand U6816 (N_6816,N_4994,N_4233);
nor U6817 (N_6817,N_5945,N_4849);
nor U6818 (N_6818,N_5665,N_4482);
xor U6819 (N_6819,N_5227,N_4750);
or U6820 (N_6820,N_5773,N_5463);
and U6821 (N_6821,N_4818,N_5597);
xnor U6822 (N_6822,N_4914,N_5126);
or U6823 (N_6823,N_4553,N_5309);
or U6824 (N_6824,N_5402,N_4337);
or U6825 (N_6825,N_4653,N_4970);
xnor U6826 (N_6826,N_4936,N_5360);
or U6827 (N_6827,N_4455,N_4180);
nand U6828 (N_6828,N_5813,N_4088);
nor U6829 (N_6829,N_4304,N_5023);
or U6830 (N_6830,N_5143,N_4965);
nand U6831 (N_6831,N_5439,N_5837);
and U6832 (N_6832,N_5391,N_4344);
nand U6833 (N_6833,N_4236,N_4795);
xor U6834 (N_6834,N_4222,N_5245);
and U6835 (N_6835,N_4543,N_5966);
or U6836 (N_6836,N_4023,N_5137);
xor U6837 (N_6837,N_4612,N_4631);
nand U6838 (N_6838,N_5618,N_4948);
or U6839 (N_6839,N_4703,N_5007);
nand U6840 (N_6840,N_4009,N_5586);
nor U6841 (N_6841,N_4924,N_4667);
xor U6842 (N_6842,N_5316,N_5458);
nand U6843 (N_6843,N_5241,N_4875);
nand U6844 (N_6844,N_4024,N_5198);
nand U6845 (N_6845,N_5011,N_5967);
xnor U6846 (N_6846,N_4178,N_4312);
nand U6847 (N_6847,N_4130,N_4069);
xor U6848 (N_6848,N_5249,N_5289);
or U6849 (N_6849,N_5861,N_5804);
or U6850 (N_6850,N_5278,N_4220);
nand U6851 (N_6851,N_5840,N_4453);
nor U6852 (N_6852,N_5865,N_4260);
or U6853 (N_6853,N_5293,N_5052);
xnor U6854 (N_6854,N_4400,N_5168);
nand U6855 (N_6855,N_4071,N_5098);
and U6856 (N_6856,N_5808,N_5783);
xnor U6857 (N_6857,N_4179,N_4846);
nor U6858 (N_6858,N_5343,N_5900);
nor U6859 (N_6859,N_4410,N_4892);
nand U6860 (N_6860,N_4823,N_5286);
xnor U6861 (N_6861,N_4519,N_5373);
nand U6862 (N_6862,N_5340,N_5788);
and U6863 (N_6863,N_5145,N_5435);
nand U6864 (N_6864,N_5158,N_5003);
nor U6865 (N_6865,N_4289,N_4561);
nand U6866 (N_6866,N_4699,N_4044);
or U6867 (N_6867,N_5453,N_5559);
xor U6868 (N_6868,N_5381,N_4246);
nand U6869 (N_6869,N_5282,N_5216);
or U6870 (N_6870,N_4596,N_4508);
xor U6871 (N_6871,N_4815,N_4365);
or U6872 (N_6872,N_5476,N_4136);
xor U6873 (N_6873,N_5623,N_5082);
xnor U6874 (N_6874,N_4783,N_5166);
and U6875 (N_6875,N_4550,N_4119);
nor U6876 (N_6876,N_4450,N_5571);
xor U6877 (N_6877,N_4191,N_5827);
nand U6878 (N_6878,N_4859,N_5021);
nand U6879 (N_6879,N_4848,N_5870);
or U6880 (N_6880,N_5594,N_4458);
or U6881 (N_6881,N_5849,N_5041);
or U6882 (N_6882,N_5497,N_5593);
nor U6883 (N_6883,N_5103,N_5419);
nand U6884 (N_6884,N_5877,N_4049);
nor U6885 (N_6885,N_4504,N_5456);
or U6886 (N_6886,N_5848,N_5949);
or U6887 (N_6887,N_5738,N_4396);
and U6888 (N_6888,N_5040,N_4131);
and U6889 (N_6889,N_4321,N_4319);
nand U6890 (N_6890,N_5250,N_5359);
nand U6891 (N_6891,N_5120,N_5954);
nor U6892 (N_6892,N_4060,N_4810);
nand U6893 (N_6893,N_4137,N_5133);
nor U6894 (N_6894,N_4657,N_5400);
nand U6895 (N_6895,N_4485,N_5290);
xnor U6896 (N_6896,N_5890,N_5829);
xor U6897 (N_6897,N_4187,N_5431);
or U6898 (N_6898,N_4956,N_5567);
and U6899 (N_6899,N_4345,N_5200);
xnor U6900 (N_6900,N_4883,N_4466);
nand U6901 (N_6901,N_5939,N_4158);
xnor U6902 (N_6902,N_4780,N_5702);
nor U6903 (N_6903,N_4430,N_4872);
or U6904 (N_6904,N_5263,N_5302);
and U6905 (N_6905,N_4183,N_4435);
or U6906 (N_6906,N_4189,N_4671);
nand U6907 (N_6907,N_5743,N_4206);
or U6908 (N_6908,N_4706,N_4122);
xnor U6909 (N_6909,N_5050,N_5180);
or U6910 (N_6910,N_5130,N_5572);
xnor U6911 (N_6911,N_5080,N_5024);
xor U6912 (N_6912,N_4512,N_5405);
and U6913 (N_6913,N_4369,N_5993);
and U6914 (N_6914,N_5220,N_5470);
and U6915 (N_6915,N_5774,N_5084);
or U6916 (N_6916,N_4133,N_4598);
and U6917 (N_6917,N_4293,N_5121);
or U6918 (N_6918,N_5450,N_4541);
nand U6919 (N_6919,N_4336,N_4972);
or U6920 (N_6920,N_5657,N_5374);
nand U6921 (N_6921,N_4755,N_4642);
and U6922 (N_6922,N_5465,N_4486);
or U6923 (N_6923,N_4765,N_5997);
and U6924 (N_6924,N_5019,N_5631);
nor U6925 (N_6925,N_5573,N_5446);
nand U6926 (N_6926,N_4392,N_5236);
nor U6927 (N_6927,N_4558,N_4799);
or U6928 (N_6928,N_5010,N_4569);
or U6929 (N_6929,N_4832,N_5576);
nor U6930 (N_6930,N_4341,N_4661);
and U6931 (N_6931,N_5613,N_5606);
and U6932 (N_6932,N_5621,N_4797);
nand U6933 (N_6933,N_5433,N_4422);
nand U6934 (N_6934,N_5974,N_5485);
nand U6935 (N_6935,N_5247,N_5395);
or U6936 (N_6936,N_4730,N_5921);
or U6937 (N_6937,N_4350,N_5792);
xor U6938 (N_6938,N_4314,N_5541);
nor U6939 (N_6939,N_4467,N_4884);
and U6940 (N_6940,N_5770,N_4204);
nor U6941 (N_6941,N_4257,N_5897);
or U6942 (N_6942,N_5600,N_5488);
nor U6943 (N_6943,N_4358,N_5226);
nand U6944 (N_6944,N_4477,N_4649);
xnor U6945 (N_6945,N_4893,N_5845);
nand U6946 (N_6946,N_4407,N_4678);
xor U6947 (N_6947,N_5810,N_4660);
xnor U6948 (N_6948,N_5733,N_4595);
xor U6949 (N_6949,N_4379,N_4065);
xor U6950 (N_6950,N_4269,N_4165);
xnor U6951 (N_6951,N_4536,N_4535);
xnor U6952 (N_6952,N_5854,N_4387);
xor U6953 (N_6953,N_4611,N_4658);
and U6954 (N_6954,N_5751,N_4692);
or U6955 (N_6955,N_5449,N_5722);
xor U6956 (N_6956,N_4766,N_5134);
nor U6957 (N_6957,N_4592,N_5523);
nand U6958 (N_6958,N_5943,N_5588);
xor U6959 (N_6959,N_5257,N_5091);
or U6960 (N_6960,N_4066,N_4110);
nand U6961 (N_6961,N_5486,N_5107);
xor U6962 (N_6962,N_4862,N_5432);
nor U6963 (N_6963,N_4079,N_5315);
nor U6964 (N_6964,N_4364,N_5101);
nor U6965 (N_6965,N_4291,N_5744);
nand U6966 (N_6966,N_5218,N_5414);
xnor U6967 (N_6967,N_5728,N_4281);
nand U6968 (N_6968,N_5025,N_5624);
nor U6969 (N_6969,N_4210,N_4151);
or U6970 (N_6970,N_5201,N_5563);
or U6971 (N_6971,N_5308,N_5676);
and U6972 (N_6972,N_5812,N_4991);
and U6973 (N_6973,N_4126,N_4479);
xor U6974 (N_6974,N_4655,N_5968);
nand U6975 (N_6975,N_5748,N_5838);
nor U6976 (N_6976,N_4913,N_4761);
and U6977 (N_6977,N_4603,N_4128);
or U6978 (N_6978,N_4711,N_4767);
nand U6979 (N_6979,N_5692,N_4201);
and U6980 (N_6980,N_5996,N_4250);
or U6981 (N_6981,N_5596,N_4142);
nand U6982 (N_6982,N_4501,N_5990);
and U6983 (N_6983,N_5790,N_5493);
or U6984 (N_6984,N_5148,N_4167);
nor U6985 (N_6985,N_5785,N_4906);
nor U6986 (N_6986,N_4175,N_4081);
and U6987 (N_6987,N_5926,N_5986);
xnor U6988 (N_6988,N_5992,N_5651);
nand U6989 (N_6989,N_4271,N_4990);
and U6990 (N_6990,N_5085,N_5033);
or U6991 (N_6991,N_5127,N_5543);
and U6992 (N_6992,N_4149,N_5407);
nor U6993 (N_6993,N_5092,N_5831);
xor U6994 (N_6994,N_5718,N_5960);
or U6995 (N_6995,N_5027,N_4245);
and U6996 (N_6996,N_5013,N_5171);
and U6997 (N_6997,N_4540,N_4383);
xnor U6998 (N_6998,N_5763,N_4626);
nor U6999 (N_6999,N_5466,N_4351);
nor U7000 (N_7000,N_4078,N_4334);
nor U7001 (N_7001,N_4154,N_5716);
xnor U7002 (N_7002,N_5583,N_4018);
nand U7003 (N_7003,N_4131,N_5589);
and U7004 (N_7004,N_5718,N_5655);
and U7005 (N_7005,N_4498,N_5031);
nand U7006 (N_7006,N_5891,N_5808);
xor U7007 (N_7007,N_4345,N_4383);
nor U7008 (N_7008,N_5938,N_4215);
and U7009 (N_7009,N_4338,N_4245);
xnor U7010 (N_7010,N_4578,N_4098);
or U7011 (N_7011,N_4872,N_5251);
nor U7012 (N_7012,N_4885,N_4627);
xnor U7013 (N_7013,N_5518,N_4503);
nand U7014 (N_7014,N_5972,N_5218);
nand U7015 (N_7015,N_5224,N_4248);
nor U7016 (N_7016,N_4995,N_4482);
and U7017 (N_7017,N_4983,N_5717);
and U7018 (N_7018,N_4251,N_4551);
and U7019 (N_7019,N_5693,N_4271);
nor U7020 (N_7020,N_5015,N_5436);
or U7021 (N_7021,N_4653,N_4662);
nor U7022 (N_7022,N_5598,N_4307);
or U7023 (N_7023,N_4522,N_5952);
and U7024 (N_7024,N_4131,N_4602);
or U7025 (N_7025,N_4850,N_4730);
nor U7026 (N_7026,N_5276,N_5246);
and U7027 (N_7027,N_4473,N_4524);
nand U7028 (N_7028,N_4498,N_4513);
nand U7029 (N_7029,N_4785,N_5167);
or U7030 (N_7030,N_5991,N_5774);
nor U7031 (N_7031,N_5420,N_4144);
or U7032 (N_7032,N_4440,N_4701);
xnor U7033 (N_7033,N_5496,N_5122);
nand U7034 (N_7034,N_4935,N_4966);
and U7035 (N_7035,N_5688,N_4625);
nand U7036 (N_7036,N_5987,N_4708);
xnor U7037 (N_7037,N_5373,N_4109);
and U7038 (N_7038,N_4612,N_5082);
or U7039 (N_7039,N_5365,N_4621);
nor U7040 (N_7040,N_5251,N_4476);
or U7041 (N_7041,N_4520,N_4462);
or U7042 (N_7042,N_4789,N_4394);
nand U7043 (N_7043,N_5536,N_4382);
and U7044 (N_7044,N_5926,N_4197);
xor U7045 (N_7045,N_4588,N_5606);
nor U7046 (N_7046,N_4509,N_4234);
xnor U7047 (N_7047,N_5799,N_5050);
xor U7048 (N_7048,N_4439,N_5831);
or U7049 (N_7049,N_5029,N_4585);
nor U7050 (N_7050,N_4461,N_4437);
nor U7051 (N_7051,N_4645,N_5536);
and U7052 (N_7052,N_5702,N_5069);
and U7053 (N_7053,N_5533,N_5423);
xnor U7054 (N_7054,N_4427,N_4220);
or U7055 (N_7055,N_4937,N_4453);
and U7056 (N_7056,N_5297,N_4855);
nand U7057 (N_7057,N_5704,N_5831);
and U7058 (N_7058,N_5539,N_5383);
xnor U7059 (N_7059,N_4132,N_5125);
nand U7060 (N_7060,N_4950,N_4744);
and U7061 (N_7061,N_4661,N_4455);
or U7062 (N_7062,N_5041,N_4933);
and U7063 (N_7063,N_5300,N_5530);
nand U7064 (N_7064,N_4128,N_4131);
nor U7065 (N_7065,N_4966,N_4980);
xor U7066 (N_7066,N_5119,N_5079);
nor U7067 (N_7067,N_4913,N_5139);
nand U7068 (N_7068,N_4724,N_4038);
nand U7069 (N_7069,N_4652,N_5225);
xor U7070 (N_7070,N_5490,N_5064);
nor U7071 (N_7071,N_5207,N_5420);
nand U7072 (N_7072,N_5734,N_5087);
and U7073 (N_7073,N_4401,N_5627);
nand U7074 (N_7074,N_5539,N_4857);
xor U7075 (N_7075,N_4230,N_5684);
nand U7076 (N_7076,N_5639,N_4806);
or U7077 (N_7077,N_5897,N_4209);
or U7078 (N_7078,N_5626,N_5627);
and U7079 (N_7079,N_4455,N_5093);
nor U7080 (N_7080,N_4775,N_5465);
and U7081 (N_7081,N_5332,N_4851);
and U7082 (N_7082,N_5691,N_5778);
xor U7083 (N_7083,N_5598,N_4787);
xnor U7084 (N_7084,N_5603,N_5981);
and U7085 (N_7085,N_5372,N_5262);
nor U7086 (N_7086,N_5046,N_5683);
or U7087 (N_7087,N_5052,N_5698);
xnor U7088 (N_7088,N_4760,N_5661);
nor U7089 (N_7089,N_4294,N_5189);
and U7090 (N_7090,N_5818,N_5841);
nand U7091 (N_7091,N_4175,N_4415);
xor U7092 (N_7092,N_5974,N_5356);
nand U7093 (N_7093,N_4750,N_4623);
or U7094 (N_7094,N_5684,N_4327);
or U7095 (N_7095,N_5035,N_5630);
or U7096 (N_7096,N_5549,N_4445);
or U7097 (N_7097,N_5400,N_4870);
nor U7098 (N_7098,N_4195,N_4229);
xor U7099 (N_7099,N_5177,N_4135);
and U7100 (N_7100,N_4065,N_4252);
xor U7101 (N_7101,N_4750,N_4388);
nor U7102 (N_7102,N_4216,N_4328);
or U7103 (N_7103,N_5872,N_4587);
xnor U7104 (N_7104,N_5769,N_5484);
nand U7105 (N_7105,N_4035,N_5943);
xnor U7106 (N_7106,N_4403,N_4162);
nor U7107 (N_7107,N_4148,N_4186);
and U7108 (N_7108,N_5722,N_5106);
and U7109 (N_7109,N_4670,N_5894);
or U7110 (N_7110,N_5994,N_4342);
or U7111 (N_7111,N_5028,N_5411);
or U7112 (N_7112,N_5828,N_5895);
nand U7113 (N_7113,N_4492,N_4019);
nor U7114 (N_7114,N_5960,N_5980);
or U7115 (N_7115,N_5744,N_4714);
xnor U7116 (N_7116,N_5981,N_5556);
nand U7117 (N_7117,N_4500,N_4384);
xnor U7118 (N_7118,N_4462,N_5322);
nand U7119 (N_7119,N_4324,N_4628);
xor U7120 (N_7120,N_5611,N_5498);
and U7121 (N_7121,N_4476,N_5605);
nor U7122 (N_7122,N_4628,N_5192);
nor U7123 (N_7123,N_4901,N_5382);
nor U7124 (N_7124,N_5437,N_4406);
nor U7125 (N_7125,N_4387,N_5238);
and U7126 (N_7126,N_4365,N_4811);
and U7127 (N_7127,N_4595,N_4585);
and U7128 (N_7128,N_4442,N_5197);
xor U7129 (N_7129,N_5112,N_5669);
and U7130 (N_7130,N_4550,N_4783);
nand U7131 (N_7131,N_4211,N_5530);
xor U7132 (N_7132,N_5588,N_4804);
and U7133 (N_7133,N_5314,N_4659);
nor U7134 (N_7134,N_4817,N_5063);
or U7135 (N_7135,N_4990,N_4216);
nor U7136 (N_7136,N_5926,N_4052);
nor U7137 (N_7137,N_4723,N_4895);
nand U7138 (N_7138,N_5926,N_5623);
nor U7139 (N_7139,N_4315,N_5127);
nand U7140 (N_7140,N_4074,N_5501);
nand U7141 (N_7141,N_5616,N_5514);
xnor U7142 (N_7142,N_4862,N_4121);
or U7143 (N_7143,N_4106,N_5947);
and U7144 (N_7144,N_4935,N_4404);
or U7145 (N_7145,N_4951,N_5435);
nand U7146 (N_7146,N_4015,N_4816);
xor U7147 (N_7147,N_4451,N_5798);
or U7148 (N_7148,N_5811,N_4909);
nor U7149 (N_7149,N_5327,N_4535);
or U7150 (N_7150,N_4295,N_4356);
xnor U7151 (N_7151,N_5889,N_5478);
nor U7152 (N_7152,N_4269,N_5271);
and U7153 (N_7153,N_5033,N_5715);
nor U7154 (N_7154,N_5082,N_4653);
or U7155 (N_7155,N_5591,N_4974);
xnor U7156 (N_7156,N_5930,N_5351);
xor U7157 (N_7157,N_5662,N_5472);
nand U7158 (N_7158,N_4917,N_5201);
and U7159 (N_7159,N_5793,N_4797);
and U7160 (N_7160,N_5640,N_4142);
nand U7161 (N_7161,N_4281,N_4177);
nor U7162 (N_7162,N_5396,N_5620);
nor U7163 (N_7163,N_5786,N_5578);
nor U7164 (N_7164,N_5483,N_5819);
or U7165 (N_7165,N_5083,N_4101);
xor U7166 (N_7166,N_4486,N_4168);
and U7167 (N_7167,N_5301,N_5188);
or U7168 (N_7168,N_4153,N_4994);
nor U7169 (N_7169,N_5696,N_5446);
and U7170 (N_7170,N_4719,N_5791);
xor U7171 (N_7171,N_5968,N_4526);
and U7172 (N_7172,N_4667,N_4009);
nor U7173 (N_7173,N_4167,N_4886);
xor U7174 (N_7174,N_5855,N_5501);
nand U7175 (N_7175,N_4504,N_4506);
nor U7176 (N_7176,N_4559,N_5516);
or U7177 (N_7177,N_5520,N_4212);
and U7178 (N_7178,N_5936,N_4474);
xnor U7179 (N_7179,N_4764,N_4674);
xnor U7180 (N_7180,N_5427,N_5602);
and U7181 (N_7181,N_4673,N_5463);
and U7182 (N_7182,N_5185,N_4970);
xnor U7183 (N_7183,N_5827,N_5801);
or U7184 (N_7184,N_4065,N_5631);
xnor U7185 (N_7185,N_5239,N_4201);
nor U7186 (N_7186,N_4598,N_5212);
or U7187 (N_7187,N_5625,N_5624);
nand U7188 (N_7188,N_5988,N_5987);
nor U7189 (N_7189,N_5714,N_4371);
xnor U7190 (N_7190,N_5660,N_4650);
xnor U7191 (N_7191,N_4302,N_4426);
and U7192 (N_7192,N_5715,N_5131);
xor U7193 (N_7193,N_4355,N_4925);
and U7194 (N_7194,N_5776,N_5785);
or U7195 (N_7195,N_4935,N_4062);
xor U7196 (N_7196,N_4220,N_4734);
xnor U7197 (N_7197,N_4952,N_4995);
and U7198 (N_7198,N_5199,N_4977);
nor U7199 (N_7199,N_5024,N_4915);
xnor U7200 (N_7200,N_4573,N_4090);
nor U7201 (N_7201,N_5013,N_4996);
and U7202 (N_7202,N_4564,N_4330);
and U7203 (N_7203,N_4164,N_4635);
nor U7204 (N_7204,N_5844,N_4015);
xor U7205 (N_7205,N_5118,N_4127);
nand U7206 (N_7206,N_4951,N_4572);
or U7207 (N_7207,N_4489,N_4638);
nand U7208 (N_7208,N_4094,N_5970);
or U7209 (N_7209,N_5419,N_5895);
and U7210 (N_7210,N_4559,N_5358);
or U7211 (N_7211,N_5173,N_5921);
xor U7212 (N_7212,N_4034,N_5165);
nand U7213 (N_7213,N_5392,N_5000);
nor U7214 (N_7214,N_4910,N_5543);
and U7215 (N_7215,N_5476,N_5394);
or U7216 (N_7216,N_5102,N_4572);
or U7217 (N_7217,N_4714,N_5504);
and U7218 (N_7218,N_5618,N_5702);
nor U7219 (N_7219,N_4730,N_5848);
and U7220 (N_7220,N_4621,N_4078);
and U7221 (N_7221,N_5305,N_4575);
nand U7222 (N_7222,N_4545,N_5287);
nand U7223 (N_7223,N_5825,N_4664);
or U7224 (N_7224,N_4850,N_4515);
nor U7225 (N_7225,N_5015,N_5861);
xnor U7226 (N_7226,N_4756,N_5459);
nor U7227 (N_7227,N_5724,N_4243);
xor U7228 (N_7228,N_5601,N_5287);
and U7229 (N_7229,N_4947,N_4837);
nor U7230 (N_7230,N_4439,N_4768);
xor U7231 (N_7231,N_4343,N_4756);
and U7232 (N_7232,N_4751,N_5123);
nand U7233 (N_7233,N_5531,N_5708);
xor U7234 (N_7234,N_5341,N_5196);
nand U7235 (N_7235,N_5277,N_4501);
xor U7236 (N_7236,N_4502,N_5969);
and U7237 (N_7237,N_5559,N_5177);
and U7238 (N_7238,N_4757,N_4229);
and U7239 (N_7239,N_5843,N_5014);
nand U7240 (N_7240,N_4499,N_4696);
or U7241 (N_7241,N_4959,N_4912);
or U7242 (N_7242,N_4599,N_4699);
and U7243 (N_7243,N_4005,N_4627);
nor U7244 (N_7244,N_4572,N_5234);
or U7245 (N_7245,N_5564,N_4282);
and U7246 (N_7246,N_5955,N_5548);
or U7247 (N_7247,N_5371,N_4601);
or U7248 (N_7248,N_4973,N_5514);
and U7249 (N_7249,N_4093,N_4617);
nor U7250 (N_7250,N_5654,N_5315);
nor U7251 (N_7251,N_4651,N_4072);
nand U7252 (N_7252,N_4866,N_4658);
xnor U7253 (N_7253,N_5370,N_5913);
nor U7254 (N_7254,N_5742,N_4248);
xnor U7255 (N_7255,N_5735,N_5451);
or U7256 (N_7256,N_4953,N_5113);
or U7257 (N_7257,N_4652,N_5628);
xor U7258 (N_7258,N_4372,N_5722);
or U7259 (N_7259,N_4803,N_5982);
nor U7260 (N_7260,N_5339,N_5619);
nor U7261 (N_7261,N_4795,N_5800);
or U7262 (N_7262,N_5737,N_4035);
nor U7263 (N_7263,N_5195,N_5085);
and U7264 (N_7264,N_4117,N_4905);
nand U7265 (N_7265,N_5704,N_4940);
or U7266 (N_7266,N_4894,N_4147);
xnor U7267 (N_7267,N_4527,N_5248);
or U7268 (N_7268,N_4962,N_5306);
nor U7269 (N_7269,N_5188,N_5866);
nor U7270 (N_7270,N_5324,N_4142);
xor U7271 (N_7271,N_4824,N_4069);
xor U7272 (N_7272,N_5984,N_4128);
and U7273 (N_7273,N_4885,N_4436);
nand U7274 (N_7274,N_5749,N_4837);
or U7275 (N_7275,N_5280,N_4589);
and U7276 (N_7276,N_4147,N_5410);
nand U7277 (N_7277,N_5078,N_5026);
or U7278 (N_7278,N_4073,N_5590);
or U7279 (N_7279,N_4853,N_5818);
nand U7280 (N_7280,N_4319,N_5281);
or U7281 (N_7281,N_5665,N_4767);
or U7282 (N_7282,N_4400,N_4715);
nand U7283 (N_7283,N_5395,N_4351);
nor U7284 (N_7284,N_4048,N_5957);
xor U7285 (N_7285,N_5392,N_4126);
and U7286 (N_7286,N_5907,N_4367);
nand U7287 (N_7287,N_4796,N_5374);
and U7288 (N_7288,N_5415,N_5820);
xor U7289 (N_7289,N_4276,N_5004);
nor U7290 (N_7290,N_5243,N_5579);
nand U7291 (N_7291,N_5068,N_4018);
or U7292 (N_7292,N_4641,N_4776);
nor U7293 (N_7293,N_5491,N_4982);
xnor U7294 (N_7294,N_5947,N_4247);
nor U7295 (N_7295,N_5413,N_4009);
xnor U7296 (N_7296,N_4329,N_4708);
and U7297 (N_7297,N_5712,N_4879);
nand U7298 (N_7298,N_4591,N_4180);
and U7299 (N_7299,N_5201,N_5864);
nand U7300 (N_7300,N_4897,N_4374);
or U7301 (N_7301,N_4175,N_4011);
nor U7302 (N_7302,N_4066,N_4914);
nand U7303 (N_7303,N_5844,N_5855);
nand U7304 (N_7304,N_5842,N_4792);
nand U7305 (N_7305,N_5394,N_4756);
and U7306 (N_7306,N_5445,N_5725);
nand U7307 (N_7307,N_5302,N_4136);
nor U7308 (N_7308,N_4460,N_5317);
or U7309 (N_7309,N_5601,N_4105);
nand U7310 (N_7310,N_5830,N_5027);
nand U7311 (N_7311,N_4810,N_4154);
or U7312 (N_7312,N_4851,N_5716);
nand U7313 (N_7313,N_5228,N_5173);
and U7314 (N_7314,N_4233,N_4253);
nor U7315 (N_7315,N_4549,N_4150);
nand U7316 (N_7316,N_4095,N_5027);
nand U7317 (N_7317,N_5617,N_5518);
and U7318 (N_7318,N_5993,N_4125);
nand U7319 (N_7319,N_4201,N_5312);
and U7320 (N_7320,N_4249,N_4416);
nand U7321 (N_7321,N_4265,N_4473);
or U7322 (N_7322,N_4193,N_4598);
or U7323 (N_7323,N_4740,N_4631);
or U7324 (N_7324,N_5236,N_5549);
and U7325 (N_7325,N_5742,N_4913);
nor U7326 (N_7326,N_4364,N_5126);
and U7327 (N_7327,N_4277,N_5795);
or U7328 (N_7328,N_5110,N_5808);
nor U7329 (N_7329,N_4832,N_4027);
and U7330 (N_7330,N_5957,N_4543);
xor U7331 (N_7331,N_4563,N_4880);
or U7332 (N_7332,N_4644,N_4822);
and U7333 (N_7333,N_4764,N_5838);
and U7334 (N_7334,N_4050,N_5711);
nand U7335 (N_7335,N_4541,N_4171);
or U7336 (N_7336,N_5900,N_5586);
xnor U7337 (N_7337,N_4941,N_4451);
or U7338 (N_7338,N_5421,N_5280);
nor U7339 (N_7339,N_4424,N_5067);
and U7340 (N_7340,N_4469,N_4630);
nor U7341 (N_7341,N_4331,N_4021);
xnor U7342 (N_7342,N_5325,N_4315);
nand U7343 (N_7343,N_5230,N_5779);
nand U7344 (N_7344,N_5753,N_4975);
nand U7345 (N_7345,N_4429,N_4926);
and U7346 (N_7346,N_4660,N_5840);
nor U7347 (N_7347,N_5088,N_5838);
and U7348 (N_7348,N_4185,N_4271);
nor U7349 (N_7349,N_4047,N_5134);
nor U7350 (N_7350,N_4094,N_5997);
nor U7351 (N_7351,N_5803,N_4929);
xor U7352 (N_7352,N_5087,N_4458);
nand U7353 (N_7353,N_4887,N_4721);
nand U7354 (N_7354,N_5129,N_5316);
or U7355 (N_7355,N_5942,N_5913);
and U7356 (N_7356,N_4888,N_5927);
xnor U7357 (N_7357,N_4816,N_5116);
xor U7358 (N_7358,N_4433,N_4514);
or U7359 (N_7359,N_4959,N_4585);
and U7360 (N_7360,N_4434,N_4399);
xor U7361 (N_7361,N_5152,N_4328);
or U7362 (N_7362,N_4755,N_4031);
nand U7363 (N_7363,N_4396,N_5741);
or U7364 (N_7364,N_4088,N_4862);
nor U7365 (N_7365,N_5421,N_4323);
xor U7366 (N_7366,N_5566,N_5816);
xor U7367 (N_7367,N_4160,N_5261);
nand U7368 (N_7368,N_4662,N_5125);
and U7369 (N_7369,N_5687,N_4725);
or U7370 (N_7370,N_4263,N_5637);
and U7371 (N_7371,N_5423,N_4775);
nand U7372 (N_7372,N_5078,N_4744);
and U7373 (N_7373,N_5142,N_4819);
xor U7374 (N_7374,N_5512,N_5171);
xor U7375 (N_7375,N_4760,N_4889);
and U7376 (N_7376,N_5509,N_5490);
or U7377 (N_7377,N_5093,N_5228);
or U7378 (N_7378,N_4280,N_5823);
xnor U7379 (N_7379,N_5982,N_4714);
nand U7380 (N_7380,N_4007,N_4908);
and U7381 (N_7381,N_5852,N_4764);
nand U7382 (N_7382,N_4392,N_5604);
or U7383 (N_7383,N_5404,N_4570);
nand U7384 (N_7384,N_5630,N_5726);
xnor U7385 (N_7385,N_5524,N_5206);
nand U7386 (N_7386,N_4536,N_4841);
nand U7387 (N_7387,N_4491,N_5449);
or U7388 (N_7388,N_5341,N_5794);
nor U7389 (N_7389,N_4014,N_4860);
xor U7390 (N_7390,N_4897,N_4989);
nor U7391 (N_7391,N_4334,N_5502);
or U7392 (N_7392,N_5201,N_5900);
nor U7393 (N_7393,N_5362,N_4724);
xnor U7394 (N_7394,N_5281,N_5651);
and U7395 (N_7395,N_4916,N_5659);
and U7396 (N_7396,N_4335,N_4841);
xnor U7397 (N_7397,N_4943,N_5164);
nor U7398 (N_7398,N_5350,N_5745);
nand U7399 (N_7399,N_4449,N_5376);
and U7400 (N_7400,N_4752,N_4268);
or U7401 (N_7401,N_5898,N_5940);
xor U7402 (N_7402,N_4380,N_4543);
nand U7403 (N_7403,N_5482,N_5562);
and U7404 (N_7404,N_5027,N_5977);
and U7405 (N_7405,N_5959,N_5215);
nand U7406 (N_7406,N_4308,N_4170);
and U7407 (N_7407,N_5000,N_5342);
nor U7408 (N_7408,N_5315,N_4746);
or U7409 (N_7409,N_5757,N_5122);
nand U7410 (N_7410,N_5332,N_4247);
xnor U7411 (N_7411,N_4684,N_4203);
xnor U7412 (N_7412,N_4542,N_4606);
xnor U7413 (N_7413,N_5097,N_5298);
nor U7414 (N_7414,N_4667,N_4581);
and U7415 (N_7415,N_5957,N_5435);
nor U7416 (N_7416,N_4634,N_4927);
or U7417 (N_7417,N_5921,N_5281);
or U7418 (N_7418,N_5086,N_4459);
or U7419 (N_7419,N_4062,N_5531);
or U7420 (N_7420,N_5150,N_5552);
and U7421 (N_7421,N_5841,N_4777);
and U7422 (N_7422,N_5997,N_4712);
nor U7423 (N_7423,N_5050,N_5591);
nor U7424 (N_7424,N_4485,N_5840);
or U7425 (N_7425,N_4244,N_4187);
and U7426 (N_7426,N_4627,N_4689);
xor U7427 (N_7427,N_5406,N_4042);
xor U7428 (N_7428,N_4339,N_4942);
and U7429 (N_7429,N_4303,N_4276);
and U7430 (N_7430,N_5118,N_5652);
xnor U7431 (N_7431,N_5670,N_4963);
nor U7432 (N_7432,N_4272,N_5385);
nor U7433 (N_7433,N_5264,N_5840);
and U7434 (N_7434,N_5349,N_4522);
or U7435 (N_7435,N_5336,N_4840);
xnor U7436 (N_7436,N_4407,N_4322);
xor U7437 (N_7437,N_5357,N_5844);
nand U7438 (N_7438,N_4896,N_5989);
or U7439 (N_7439,N_5548,N_4920);
nor U7440 (N_7440,N_5777,N_5871);
or U7441 (N_7441,N_5984,N_4076);
or U7442 (N_7442,N_4211,N_4596);
or U7443 (N_7443,N_5523,N_4197);
xnor U7444 (N_7444,N_4578,N_4657);
and U7445 (N_7445,N_4467,N_4403);
or U7446 (N_7446,N_5520,N_5733);
or U7447 (N_7447,N_5304,N_5415);
xnor U7448 (N_7448,N_5099,N_4394);
or U7449 (N_7449,N_5372,N_5661);
or U7450 (N_7450,N_5890,N_5834);
nor U7451 (N_7451,N_5632,N_5688);
xnor U7452 (N_7452,N_5297,N_4557);
nand U7453 (N_7453,N_5022,N_5725);
nor U7454 (N_7454,N_4907,N_5894);
nand U7455 (N_7455,N_5076,N_4163);
xor U7456 (N_7456,N_4982,N_4246);
or U7457 (N_7457,N_5707,N_4198);
nor U7458 (N_7458,N_5699,N_4130);
nor U7459 (N_7459,N_4476,N_5501);
xnor U7460 (N_7460,N_5564,N_4118);
or U7461 (N_7461,N_5164,N_4303);
nor U7462 (N_7462,N_4696,N_4230);
and U7463 (N_7463,N_4613,N_5101);
nor U7464 (N_7464,N_4839,N_4431);
and U7465 (N_7465,N_5954,N_4910);
or U7466 (N_7466,N_5300,N_5127);
xnor U7467 (N_7467,N_4427,N_4549);
or U7468 (N_7468,N_4006,N_4754);
nand U7469 (N_7469,N_4462,N_4850);
nor U7470 (N_7470,N_5960,N_4482);
nand U7471 (N_7471,N_4105,N_4304);
nor U7472 (N_7472,N_5654,N_5753);
or U7473 (N_7473,N_4624,N_5685);
nor U7474 (N_7474,N_4636,N_5985);
nand U7475 (N_7475,N_5157,N_4400);
xnor U7476 (N_7476,N_4636,N_5983);
and U7477 (N_7477,N_5589,N_4423);
nor U7478 (N_7478,N_4424,N_5573);
and U7479 (N_7479,N_5060,N_5870);
nor U7480 (N_7480,N_5799,N_5703);
or U7481 (N_7481,N_5207,N_4660);
xnor U7482 (N_7482,N_5982,N_5403);
nor U7483 (N_7483,N_4169,N_5292);
nand U7484 (N_7484,N_4378,N_4646);
nand U7485 (N_7485,N_5158,N_4241);
nand U7486 (N_7486,N_4151,N_5023);
nand U7487 (N_7487,N_5571,N_5568);
nand U7488 (N_7488,N_4282,N_5970);
or U7489 (N_7489,N_4312,N_5564);
and U7490 (N_7490,N_5391,N_4766);
xor U7491 (N_7491,N_5389,N_4707);
nand U7492 (N_7492,N_5785,N_4259);
nor U7493 (N_7493,N_5774,N_4563);
and U7494 (N_7494,N_5961,N_4478);
xnor U7495 (N_7495,N_4133,N_4057);
or U7496 (N_7496,N_4368,N_5183);
or U7497 (N_7497,N_5376,N_5262);
nor U7498 (N_7498,N_5863,N_4149);
xor U7499 (N_7499,N_4393,N_5760);
and U7500 (N_7500,N_4604,N_4336);
xor U7501 (N_7501,N_5193,N_5529);
nor U7502 (N_7502,N_5659,N_5480);
xor U7503 (N_7503,N_5714,N_4915);
and U7504 (N_7504,N_4831,N_5132);
nor U7505 (N_7505,N_4974,N_4474);
nand U7506 (N_7506,N_4392,N_5883);
nand U7507 (N_7507,N_4200,N_5813);
or U7508 (N_7508,N_5459,N_4635);
xor U7509 (N_7509,N_4550,N_4092);
and U7510 (N_7510,N_5076,N_4675);
nor U7511 (N_7511,N_5714,N_4788);
or U7512 (N_7512,N_4100,N_4448);
nand U7513 (N_7513,N_4489,N_5988);
xor U7514 (N_7514,N_5845,N_4100);
xor U7515 (N_7515,N_5462,N_5477);
or U7516 (N_7516,N_5697,N_4579);
xor U7517 (N_7517,N_5258,N_5009);
and U7518 (N_7518,N_5697,N_4131);
or U7519 (N_7519,N_5858,N_5895);
or U7520 (N_7520,N_4080,N_4382);
and U7521 (N_7521,N_5040,N_4148);
xor U7522 (N_7522,N_4722,N_5029);
nand U7523 (N_7523,N_5681,N_5656);
xor U7524 (N_7524,N_4590,N_4889);
nor U7525 (N_7525,N_5111,N_4300);
nor U7526 (N_7526,N_4137,N_5879);
nand U7527 (N_7527,N_5215,N_5158);
xnor U7528 (N_7528,N_5339,N_5215);
nor U7529 (N_7529,N_4964,N_5258);
nor U7530 (N_7530,N_4983,N_5304);
or U7531 (N_7531,N_4521,N_4438);
nand U7532 (N_7532,N_5543,N_4452);
or U7533 (N_7533,N_4832,N_4517);
xor U7534 (N_7534,N_4368,N_5023);
and U7535 (N_7535,N_5850,N_5478);
nand U7536 (N_7536,N_4979,N_4698);
nand U7537 (N_7537,N_5520,N_4981);
or U7538 (N_7538,N_5660,N_5981);
and U7539 (N_7539,N_5121,N_5440);
xnor U7540 (N_7540,N_5998,N_5467);
nor U7541 (N_7541,N_5595,N_4631);
nand U7542 (N_7542,N_4252,N_4204);
nor U7543 (N_7543,N_4117,N_5914);
nor U7544 (N_7544,N_5992,N_5492);
or U7545 (N_7545,N_5883,N_4933);
or U7546 (N_7546,N_4269,N_4279);
nand U7547 (N_7547,N_5380,N_5770);
nor U7548 (N_7548,N_5304,N_5787);
and U7549 (N_7549,N_5956,N_4180);
or U7550 (N_7550,N_4416,N_4687);
xor U7551 (N_7551,N_4276,N_4213);
nand U7552 (N_7552,N_5872,N_5738);
or U7553 (N_7553,N_5156,N_5085);
xnor U7554 (N_7554,N_4256,N_4805);
xor U7555 (N_7555,N_4781,N_5322);
or U7556 (N_7556,N_5271,N_4760);
nor U7557 (N_7557,N_4310,N_4317);
xnor U7558 (N_7558,N_5788,N_4139);
nor U7559 (N_7559,N_4149,N_5806);
nand U7560 (N_7560,N_4945,N_4699);
nor U7561 (N_7561,N_5877,N_4096);
or U7562 (N_7562,N_5529,N_4160);
and U7563 (N_7563,N_5785,N_5809);
nand U7564 (N_7564,N_5152,N_4047);
and U7565 (N_7565,N_4553,N_4528);
nor U7566 (N_7566,N_5997,N_4012);
nor U7567 (N_7567,N_4125,N_4966);
xor U7568 (N_7568,N_4563,N_5878);
nor U7569 (N_7569,N_4144,N_4726);
nand U7570 (N_7570,N_4239,N_5763);
nand U7571 (N_7571,N_4503,N_4120);
and U7572 (N_7572,N_4739,N_4954);
xor U7573 (N_7573,N_5534,N_5328);
and U7574 (N_7574,N_4849,N_4395);
nand U7575 (N_7575,N_4439,N_5061);
nand U7576 (N_7576,N_4113,N_4328);
xor U7577 (N_7577,N_5273,N_4708);
nand U7578 (N_7578,N_5411,N_5344);
or U7579 (N_7579,N_4446,N_5915);
and U7580 (N_7580,N_5838,N_4544);
and U7581 (N_7581,N_5653,N_4979);
and U7582 (N_7582,N_5255,N_4889);
xor U7583 (N_7583,N_4076,N_4081);
nor U7584 (N_7584,N_5562,N_5872);
nand U7585 (N_7585,N_5663,N_4490);
or U7586 (N_7586,N_4019,N_5180);
xnor U7587 (N_7587,N_4433,N_5146);
nand U7588 (N_7588,N_5365,N_4911);
nand U7589 (N_7589,N_4282,N_5679);
xor U7590 (N_7590,N_4969,N_4518);
nor U7591 (N_7591,N_5147,N_4902);
or U7592 (N_7592,N_4299,N_5468);
xnor U7593 (N_7593,N_4070,N_5869);
and U7594 (N_7594,N_4963,N_4074);
xor U7595 (N_7595,N_4608,N_5748);
nand U7596 (N_7596,N_4225,N_4406);
nand U7597 (N_7597,N_4837,N_4049);
and U7598 (N_7598,N_5827,N_5226);
and U7599 (N_7599,N_4535,N_5641);
and U7600 (N_7600,N_5603,N_4071);
nor U7601 (N_7601,N_5514,N_4474);
and U7602 (N_7602,N_5075,N_4375);
or U7603 (N_7603,N_5774,N_5958);
or U7604 (N_7604,N_4350,N_4748);
nand U7605 (N_7605,N_4135,N_5110);
nand U7606 (N_7606,N_5875,N_5297);
nor U7607 (N_7607,N_4364,N_4214);
and U7608 (N_7608,N_5959,N_4598);
xor U7609 (N_7609,N_5518,N_4874);
nand U7610 (N_7610,N_4600,N_4247);
and U7611 (N_7611,N_5662,N_5309);
xnor U7612 (N_7612,N_4567,N_5210);
and U7613 (N_7613,N_4552,N_4792);
nand U7614 (N_7614,N_5519,N_5235);
xor U7615 (N_7615,N_5511,N_4660);
and U7616 (N_7616,N_4036,N_5396);
and U7617 (N_7617,N_4811,N_4241);
xnor U7618 (N_7618,N_5575,N_5492);
or U7619 (N_7619,N_4901,N_4929);
xnor U7620 (N_7620,N_4250,N_5633);
or U7621 (N_7621,N_4785,N_4090);
and U7622 (N_7622,N_5124,N_5375);
and U7623 (N_7623,N_5148,N_5784);
or U7624 (N_7624,N_4523,N_5509);
xnor U7625 (N_7625,N_5500,N_4225);
and U7626 (N_7626,N_4358,N_5634);
xor U7627 (N_7627,N_5535,N_4034);
xnor U7628 (N_7628,N_4923,N_4950);
and U7629 (N_7629,N_5335,N_5166);
nor U7630 (N_7630,N_5645,N_5151);
nand U7631 (N_7631,N_5169,N_5590);
xor U7632 (N_7632,N_5507,N_5629);
and U7633 (N_7633,N_5150,N_5202);
nor U7634 (N_7634,N_5020,N_5776);
nand U7635 (N_7635,N_4840,N_5790);
or U7636 (N_7636,N_5641,N_4367);
xor U7637 (N_7637,N_4843,N_4801);
nor U7638 (N_7638,N_5083,N_4269);
and U7639 (N_7639,N_5859,N_4598);
xnor U7640 (N_7640,N_5021,N_4979);
or U7641 (N_7641,N_4671,N_4580);
nand U7642 (N_7642,N_4051,N_5976);
and U7643 (N_7643,N_5773,N_4485);
xnor U7644 (N_7644,N_4265,N_5133);
nor U7645 (N_7645,N_5399,N_4248);
nand U7646 (N_7646,N_5592,N_5428);
and U7647 (N_7647,N_4294,N_4645);
and U7648 (N_7648,N_5671,N_5348);
or U7649 (N_7649,N_4549,N_4784);
nand U7650 (N_7650,N_4049,N_5829);
and U7651 (N_7651,N_4796,N_4088);
nand U7652 (N_7652,N_4809,N_5889);
nor U7653 (N_7653,N_5480,N_4454);
or U7654 (N_7654,N_5263,N_5201);
and U7655 (N_7655,N_4007,N_4637);
nand U7656 (N_7656,N_5241,N_4694);
or U7657 (N_7657,N_5316,N_5930);
and U7658 (N_7658,N_4021,N_4985);
or U7659 (N_7659,N_4299,N_4487);
and U7660 (N_7660,N_4486,N_4699);
nor U7661 (N_7661,N_5564,N_4821);
nand U7662 (N_7662,N_5302,N_4724);
nand U7663 (N_7663,N_5280,N_4687);
and U7664 (N_7664,N_4372,N_4706);
xor U7665 (N_7665,N_4108,N_4809);
xor U7666 (N_7666,N_5592,N_5230);
nor U7667 (N_7667,N_5744,N_4957);
nand U7668 (N_7668,N_5289,N_4454);
xnor U7669 (N_7669,N_4006,N_4806);
xor U7670 (N_7670,N_5766,N_5914);
nand U7671 (N_7671,N_4276,N_5325);
nand U7672 (N_7672,N_4490,N_5425);
xnor U7673 (N_7673,N_4219,N_4535);
xor U7674 (N_7674,N_5602,N_5847);
and U7675 (N_7675,N_4698,N_4776);
nor U7676 (N_7676,N_5260,N_4742);
nor U7677 (N_7677,N_5361,N_4710);
xnor U7678 (N_7678,N_4248,N_5344);
and U7679 (N_7679,N_4498,N_4834);
nor U7680 (N_7680,N_4046,N_4465);
xor U7681 (N_7681,N_4746,N_4329);
or U7682 (N_7682,N_5761,N_5722);
or U7683 (N_7683,N_5546,N_4795);
and U7684 (N_7684,N_5987,N_5391);
nand U7685 (N_7685,N_5390,N_5533);
nand U7686 (N_7686,N_4232,N_4202);
nand U7687 (N_7687,N_4767,N_4020);
nor U7688 (N_7688,N_4599,N_5847);
or U7689 (N_7689,N_5523,N_4230);
and U7690 (N_7690,N_4243,N_5711);
nor U7691 (N_7691,N_5813,N_4265);
nand U7692 (N_7692,N_4060,N_5657);
and U7693 (N_7693,N_5496,N_4001);
and U7694 (N_7694,N_5851,N_4768);
xnor U7695 (N_7695,N_4834,N_5536);
and U7696 (N_7696,N_5664,N_5195);
and U7697 (N_7697,N_4256,N_5464);
nand U7698 (N_7698,N_5440,N_4969);
xor U7699 (N_7699,N_4677,N_5039);
and U7700 (N_7700,N_5676,N_5938);
or U7701 (N_7701,N_5916,N_5572);
and U7702 (N_7702,N_4127,N_5130);
nor U7703 (N_7703,N_5512,N_4608);
or U7704 (N_7704,N_5428,N_5577);
nor U7705 (N_7705,N_5652,N_5962);
nand U7706 (N_7706,N_4485,N_5490);
or U7707 (N_7707,N_4204,N_5805);
nor U7708 (N_7708,N_5871,N_5102);
and U7709 (N_7709,N_5243,N_5528);
and U7710 (N_7710,N_5493,N_5752);
or U7711 (N_7711,N_5475,N_5348);
or U7712 (N_7712,N_5297,N_4261);
or U7713 (N_7713,N_4532,N_5492);
xor U7714 (N_7714,N_4772,N_5275);
or U7715 (N_7715,N_5958,N_4580);
or U7716 (N_7716,N_4135,N_4606);
and U7717 (N_7717,N_5052,N_5389);
nor U7718 (N_7718,N_5256,N_5832);
nor U7719 (N_7719,N_5424,N_4878);
and U7720 (N_7720,N_4713,N_4991);
xor U7721 (N_7721,N_4634,N_4291);
nand U7722 (N_7722,N_4520,N_5602);
xnor U7723 (N_7723,N_5792,N_5299);
or U7724 (N_7724,N_4585,N_5008);
nand U7725 (N_7725,N_5687,N_4235);
nand U7726 (N_7726,N_4558,N_4949);
xor U7727 (N_7727,N_5771,N_4591);
nor U7728 (N_7728,N_4085,N_4541);
and U7729 (N_7729,N_5262,N_5456);
nand U7730 (N_7730,N_4514,N_5945);
nor U7731 (N_7731,N_5795,N_5606);
nand U7732 (N_7732,N_4441,N_5060);
or U7733 (N_7733,N_4356,N_4364);
xnor U7734 (N_7734,N_4566,N_4142);
xor U7735 (N_7735,N_5259,N_5384);
or U7736 (N_7736,N_5804,N_4848);
or U7737 (N_7737,N_4742,N_5302);
nand U7738 (N_7738,N_4690,N_5339);
xnor U7739 (N_7739,N_5022,N_4024);
xnor U7740 (N_7740,N_4696,N_5439);
and U7741 (N_7741,N_4519,N_5191);
xor U7742 (N_7742,N_5015,N_4839);
or U7743 (N_7743,N_4261,N_5557);
nand U7744 (N_7744,N_5881,N_5981);
nor U7745 (N_7745,N_5459,N_5324);
xnor U7746 (N_7746,N_5991,N_4341);
nor U7747 (N_7747,N_4713,N_5641);
xor U7748 (N_7748,N_4303,N_5569);
or U7749 (N_7749,N_5417,N_5095);
or U7750 (N_7750,N_4249,N_4642);
nand U7751 (N_7751,N_4546,N_5357);
nor U7752 (N_7752,N_5928,N_5979);
xor U7753 (N_7753,N_5910,N_5168);
or U7754 (N_7754,N_5981,N_4673);
or U7755 (N_7755,N_4256,N_4970);
nand U7756 (N_7756,N_5422,N_4428);
and U7757 (N_7757,N_4580,N_4973);
xor U7758 (N_7758,N_4561,N_4341);
and U7759 (N_7759,N_5051,N_5220);
nand U7760 (N_7760,N_5986,N_4157);
nand U7761 (N_7761,N_5442,N_4273);
nor U7762 (N_7762,N_4618,N_4397);
nand U7763 (N_7763,N_5405,N_5243);
and U7764 (N_7764,N_5464,N_4447);
nand U7765 (N_7765,N_5671,N_4719);
nor U7766 (N_7766,N_4842,N_4880);
xor U7767 (N_7767,N_4245,N_5259);
nand U7768 (N_7768,N_5221,N_5716);
nor U7769 (N_7769,N_5759,N_4384);
and U7770 (N_7770,N_5859,N_4796);
nor U7771 (N_7771,N_5283,N_5722);
or U7772 (N_7772,N_4464,N_4478);
xnor U7773 (N_7773,N_4214,N_5967);
and U7774 (N_7774,N_4785,N_4788);
or U7775 (N_7775,N_5993,N_4152);
xor U7776 (N_7776,N_5935,N_4566);
nand U7777 (N_7777,N_4852,N_4306);
nand U7778 (N_7778,N_4268,N_5552);
or U7779 (N_7779,N_5878,N_5503);
or U7780 (N_7780,N_4910,N_5217);
xor U7781 (N_7781,N_5842,N_4680);
nor U7782 (N_7782,N_5718,N_5684);
and U7783 (N_7783,N_4845,N_5529);
nand U7784 (N_7784,N_5241,N_5681);
nand U7785 (N_7785,N_4228,N_4825);
and U7786 (N_7786,N_5131,N_5513);
and U7787 (N_7787,N_5728,N_5908);
nor U7788 (N_7788,N_4525,N_4479);
xor U7789 (N_7789,N_4016,N_5122);
nand U7790 (N_7790,N_4549,N_4905);
and U7791 (N_7791,N_4470,N_5620);
nand U7792 (N_7792,N_4788,N_4657);
nand U7793 (N_7793,N_4225,N_5033);
nand U7794 (N_7794,N_5504,N_4623);
and U7795 (N_7795,N_5500,N_5552);
nand U7796 (N_7796,N_5139,N_4411);
xnor U7797 (N_7797,N_4827,N_5210);
nand U7798 (N_7798,N_4264,N_4702);
or U7799 (N_7799,N_5978,N_4674);
or U7800 (N_7800,N_4665,N_5226);
nand U7801 (N_7801,N_5743,N_4594);
and U7802 (N_7802,N_4303,N_5700);
nand U7803 (N_7803,N_4673,N_4156);
and U7804 (N_7804,N_5905,N_4458);
and U7805 (N_7805,N_5252,N_5932);
or U7806 (N_7806,N_4893,N_4308);
xnor U7807 (N_7807,N_5381,N_5613);
and U7808 (N_7808,N_5307,N_4154);
nand U7809 (N_7809,N_5392,N_4356);
nor U7810 (N_7810,N_4399,N_4617);
and U7811 (N_7811,N_5044,N_4164);
nor U7812 (N_7812,N_4063,N_5031);
nand U7813 (N_7813,N_4635,N_4249);
nand U7814 (N_7814,N_5149,N_4153);
nand U7815 (N_7815,N_5035,N_4697);
nand U7816 (N_7816,N_4922,N_4756);
or U7817 (N_7817,N_5700,N_5175);
nand U7818 (N_7818,N_4080,N_4653);
and U7819 (N_7819,N_4311,N_4759);
or U7820 (N_7820,N_5679,N_5039);
nor U7821 (N_7821,N_4853,N_5689);
and U7822 (N_7822,N_4457,N_4368);
nand U7823 (N_7823,N_4096,N_4885);
and U7824 (N_7824,N_4142,N_5630);
and U7825 (N_7825,N_4362,N_4254);
nor U7826 (N_7826,N_4864,N_4535);
and U7827 (N_7827,N_5060,N_4400);
nand U7828 (N_7828,N_5587,N_5069);
nor U7829 (N_7829,N_4063,N_4635);
and U7830 (N_7830,N_5672,N_4906);
xnor U7831 (N_7831,N_4186,N_5893);
nand U7832 (N_7832,N_4569,N_4344);
and U7833 (N_7833,N_4241,N_5873);
nor U7834 (N_7834,N_5918,N_5178);
or U7835 (N_7835,N_4583,N_4581);
xor U7836 (N_7836,N_4147,N_4886);
xnor U7837 (N_7837,N_5366,N_4752);
nand U7838 (N_7838,N_5720,N_4799);
nor U7839 (N_7839,N_5004,N_5539);
or U7840 (N_7840,N_4023,N_4427);
nor U7841 (N_7841,N_4551,N_4068);
nand U7842 (N_7842,N_4120,N_4150);
and U7843 (N_7843,N_4279,N_5523);
or U7844 (N_7844,N_5987,N_4310);
nor U7845 (N_7845,N_4180,N_5038);
xnor U7846 (N_7846,N_5953,N_4140);
nor U7847 (N_7847,N_4680,N_4087);
nor U7848 (N_7848,N_4958,N_5891);
xor U7849 (N_7849,N_5487,N_5526);
xnor U7850 (N_7850,N_5458,N_5543);
and U7851 (N_7851,N_4226,N_5563);
or U7852 (N_7852,N_4686,N_5048);
xor U7853 (N_7853,N_4995,N_4887);
nand U7854 (N_7854,N_5170,N_5996);
xor U7855 (N_7855,N_5224,N_4752);
or U7856 (N_7856,N_4216,N_4479);
and U7857 (N_7857,N_4836,N_4346);
nand U7858 (N_7858,N_4587,N_5123);
nand U7859 (N_7859,N_4938,N_4476);
or U7860 (N_7860,N_5733,N_5064);
or U7861 (N_7861,N_5233,N_5597);
nor U7862 (N_7862,N_5269,N_4578);
and U7863 (N_7863,N_5099,N_4188);
and U7864 (N_7864,N_4325,N_4633);
nor U7865 (N_7865,N_4311,N_5760);
xnor U7866 (N_7866,N_4135,N_4524);
xor U7867 (N_7867,N_4501,N_4453);
and U7868 (N_7868,N_5287,N_5433);
xor U7869 (N_7869,N_5903,N_4180);
nor U7870 (N_7870,N_5343,N_5988);
and U7871 (N_7871,N_5445,N_4169);
nand U7872 (N_7872,N_5955,N_4264);
or U7873 (N_7873,N_5783,N_5135);
nor U7874 (N_7874,N_5983,N_4190);
nand U7875 (N_7875,N_4390,N_4454);
nand U7876 (N_7876,N_5916,N_4257);
or U7877 (N_7877,N_4550,N_4672);
and U7878 (N_7878,N_4108,N_5867);
xnor U7879 (N_7879,N_4065,N_4426);
nand U7880 (N_7880,N_5001,N_5278);
nand U7881 (N_7881,N_4203,N_5230);
xnor U7882 (N_7882,N_4554,N_5092);
xnor U7883 (N_7883,N_5305,N_5461);
nor U7884 (N_7884,N_4279,N_4772);
and U7885 (N_7885,N_5456,N_4236);
xor U7886 (N_7886,N_5276,N_5061);
and U7887 (N_7887,N_5873,N_4619);
nand U7888 (N_7888,N_5946,N_4278);
and U7889 (N_7889,N_5292,N_4130);
xnor U7890 (N_7890,N_5407,N_4197);
and U7891 (N_7891,N_5388,N_4411);
and U7892 (N_7892,N_5954,N_5402);
nor U7893 (N_7893,N_5894,N_5627);
nand U7894 (N_7894,N_5973,N_5028);
nand U7895 (N_7895,N_4351,N_4979);
nand U7896 (N_7896,N_5429,N_5456);
nand U7897 (N_7897,N_5953,N_5515);
nor U7898 (N_7898,N_4838,N_4525);
and U7899 (N_7899,N_4667,N_5116);
and U7900 (N_7900,N_5884,N_5886);
xnor U7901 (N_7901,N_5517,N_5617);
nand U7902 (N_7902,N_4242,N_5908);
nor U7903 (N_7903,N_4657,N_4095);
or U7904 (N_7904,N_5193,N_5202);
nor U7905 (N_7905,N_5147,N_4289);
and U7906 (N_7906,N_5272,N_5337);
nor U7907 (N_7907,N_4912,N_4416);
xnor U7908 (N_7908,N_5759,N_4805);
nor U7909 (N_7909,N_4078,N_4738);
xor U7910 (N_7910,N_4537,N_4598);
xor U7911 (N_7911,N_4054,N_5958);
or U7912 (N_7912,N_4937,N_5215);
nand U7913 (N_7913,N_5553,N_5251);
and U7914 (N_7914,N_4954,N_4035);
or U7915 (N_7915,N_5177,N_4841);
nor U7916 (N_7916,N_5706,N_5532);
nand U7917 (N_7917,N_4588,N_5627);
or U7918 (N_7918,N_5507,N_5065);
or U7919 (N_7919,N_5512,N_5594);
and U7920 (N_7920,N_4683,N_5316);
nand U7921 (N_7921,N_4658,N_5077);
nand U7922 (N_7922,N_4898,N_4838);
nand U7923 (N_7923,N_5571,N_5493);
xnor U7924 (N_7924,N_4928,N_4219);
nand U7925 (N_7925,N_4540,N_5571);
nand U7926 (N_7926,N_5196,N_5579);
or U7927 (N_7927,N_5282,N_5206);
xor U7928 (N_7928,N_4945,N_5131);
nand U7929 (N_7929,N_5143,N_5718);
or U7930 (N_7930,N_4046,N_5619);
xnor U7931 (N_7931,N_5123,N_4738);
nand U7932 (N_7932,N_4084,N_4869);
nor U7933 (N_7933,N_5952,N_5942);
xor U7934 (N_7934,N_4219,N_4828);
xnor U7935 (N_7935,N_5648,N_5274);
nor U7936 (N_7936,N_5104,N_5633);
and U7937 (N_7937,N_4941,N_4472);
nand U7938 (N_7938,N_4289,N_5611);
nand U7939 (N_7939,N_4050,N_4201);
and U7940 (N_7940,N_5083,N_5866);
nand U7941 (N_7941,N_4272,N_5604);
and U7942 (N_7942,N_5831,N_4060);
or U7943 (N_7943,N_5934,N_4949);
or U7944 (N_7944,N_4216,N_4231);
xor U7945 (N_7945,N_5625,N_5031);
or U7946 (N_7946,N_5144,N_5575);
nor U7947 (N_7947,N_4483,N_4953);
xnor U7948 (N_7948,N_5229,N_4005);
or U7949 (N_7949,N_5285,N_4170);
xor U7950 (N_7950,N_5634,N_5948);
nor U7951 (N_7951,N_4717,N_4154);
and U7952 (N_7952,N_4667,N_5948);
nand U7953 (N_7953,N_5668,N_4903);
or U7954 (N_7954,N_4850,N_5692);
nor U7955 (N_7955,N_4257,N_5680);
nand U7956 (N_7956,N_4020,N_4615);
xor U7957 (N_7957,N_4920,N_5465);
and U7958 (N_7958,N_4692,N_5724);
xnor U7959 (N_7959,N_4969,N_5916);
and U7960 (N_7960,N_5493,N_5512);
xnor U7961 (N_7961,N_4948,N_5742);
nor U7962 (N_7962,N_5001,N_5345);
xor U7963 (N_7963,N_4455,N_4105);
or U7964 (N_7964,N_5658,N_4533);
and U7965 (N_7965,N_5830,N_5102);
nand U7966 (N_7966,N_4274,N_4354);
xnor U7967 (N_7967,N_5795,N_5070);
nand U7968 (N_7968,N_5721,N_5365);
nor U7969 (N_7969,N_4483,N_4631);
nor U7970 (N_7970,N_4061,N_4758);
xnor U7971 (N_7971,N_5837,N_5976);
nand U7972 (N_7972,N_4362,N_5537);
and U7973 (N_7973,N_5870,N_4931);
and U7974 (N_7974,N_5080,N_4743);
and U7975 (N_7975,N_5407,N_5916);
and U7976 (N_7976,N_5541,N_4723);
nand U7977 (N_7977,N_5602,N_5439);
xor U7978 (N_7978,N_4764,N_4857);
nor U7979 (N_7979,N_5802,N_5500);
nor U7980 (N_7980,N_5214,N_4113);
and U7981 (N_7981,N_4753,N_4612);
nand U7982 (N_7982,N_4692,N_5903);
or U7983 (N_7983,N_5054,N_5493);
and U7984 (N_7984,N_5671,N_5323);
and U7985 (N_7985,N_5669,N_4416);
nor U7986 (N_7986,N_5683,N_5949);
nand U7987 (N_7987,N_4521,N_5350);
or U7988 (N_7988,N_5340,N_4600);
nand U7989 (N_7989,N_5241,N_5058);
nand U7990 (N_7990,N_4323,N_4035);
xor U7991 (N_7991,N_4748,N_5082);
and U7992 (N_7992,N_5950,N_4412);
nor U7993 (N_7993,N_5698,N_5049);
xor U7994 (N_7994,N_4692,N_4140);
nand U7995 (N_7995,N_4753,N_5839);
or U7996 (N_7996,N_5374,N_4742);
or U7997 (N_7997,N_4314,N_5989);
or U7998 (N_7998,N_4185,N_4550);
nor U7999 (N_7999,N_4726,N_5382);
and U8000 (N_8000,N_6288,N_7888);
nand U8001 (N_8001,N_7722,N_6051);
xnor U8002 (N_8002,N_6322,N_6742);
xnor U8003 (N_8003,N_7474,N_6090);
xor U8004 (N_8004,N_7876,N_7564);
nand U8005 (N_8005,N_7924,N_7251);
nor U8006 (N_8006,N_6161,N_7245);
nand U8007 (N_8007,N_6219,N_6457);
nand U8008 (N_8008,N_6330,N_6080);
and U8009 (N_8009,N_7543,N_7059);
nand U8010 (N_8010,N_6493,N_6429);
xor U8011 (N_8011,N_6842,N_7110);
and U8012 (N_8012,N_7552,N_7829);
or U8013 (N_8013,N_6784,N_7470);
or U8014 (N_8014,N_7666,N_7003);
nand U8015 (N_8015,N_6936,N_6922);
and U8016 (N_8016,N_7312,N_7200);
and U8017 (N_8017,N_7280,N_7426);
xnor U8018 (N_8018,N_6260,N_7535);
nand U8019 (N_8019,N_6271,N_6082);
nor U8020 (N_8020,N_7310,N_6924);
or U8021 (N_8021,N_7771,N_6024);
or U8022 (N_8022,N_6737,N_6909);
xor U8023 (N_8023,N_7658,N_6932);
xor U8024 (N_8024,N_6587,N_7826);
nand U8025 (N_8025,N_6549,N_6809);
nor U8026 (N_8026,N_6362,N_7659);
and U8027 (N_8027,N_7051,N_7174);
or U8028 (N_8028,N_6403,N_6767);
nor U8029 (N_8029,N_6116,N_6751);
nor U8030 (N_8030,N_6861,N_6658);
nand U8031 (N_8031,N_7612,N_6480);
or U8032 (N_8032,N_7592,N_6631);
or U8033 (N_8033,N_6278,N_6426);
or U8034 (N_8034,N_7134,N_6298);
nor U8035 (N_8035,N_7387,N_6018);
nand U8036 (N_8036,N_6764,N_7299);
xnor U8037 (N_8037,N_7754,N_6409);
xor U8038 (N_8038,N_7716,N_6999);
nor U8039 (N_8039,N_6202,N_6665);
xnor U8040 (N_8040,N_7024,N_7480);
and U8041 (N_8041,N_7711,N_7545);
xor U8042 (N_8042,N_6092,N_7979);
nor U8043 (N_8043,N_6551,N_7911);
nor U8044 (N_8044,N_7842,N_7295);
xnor U8045 (N_8045,N_6319,N_6828);
nand U8046 (N_8046,N_6451,N_7331);
xor U8047 (N_8047,N_7550,N_7120);
and U8048 (N_8048,N_6006,N_7640);
xor U8049 (N_8049,N_6688,N_7524);
nor U8050 (N_8050,N_6479,N_7297);
or U8051 (N_8051,N_7585,N_7157);
and U8052 (N_8052,N_6944,N_7928);
nand U8053 (N_8053,N_7981,N_6912);
xnor U8054 (N_8054,N_6898,N_7663);
nor U8055 (N_8055,N_6388,N_6340);
or U8056 (N_8056,N_7142,N_6647);
nand U8057 (N_8057,N_6789,N_6565);
and U8058 (N_8058,N_7737,N_6685);
or U8059 (N_8059,N_7149,N_7267);
and U8060 (N_8060,N_7109,N_6946);
nor U8061 (N_8061,N_6947,N_6572);
xnor U8062 (N_8062,N_7909,N_6763);
or U8063 (N_8063,N_7094,N_7869);
nand U8064 (N_8064,N_7424,N_6229);
xor U8065 (N_8065,N_7671,N_6239);
nor U8066 (N_8066,N_7069,N_7063);
nor U8067 (N_8067,N_7496,N_7043);
nand U8068 (N_8068,N_7313,N_6207);
xnor U8069 (N_8069,N_6821,N_7165);
nand U8070 (N_8070,N_7817,N_6435);
nand U8071 (N_8071,N_6610,N_6150);
and U8072 (N_8072,N_6183,N_7664);
nor U8073 (N_8073,N_7115,N_6738);
nor U8074 (N_8074,N_6146,N_7974);
nand U8075 (N_8075,N_6920,N_7554);
xor U8076 (N_8076,N_7400,N_6145);
xnor U8077 (N_8077,N_6848,N_7561);
nor U8078 (N_8078,N_6530,N_6351);
and U8079 (N_8079,N_7744,N_6277);
or U8080 (N_8080,N_7401,N_7616);
xor U8081 (N_8081,N_7361,N_7795);
and U8082 (N_8082,N_7075,N_7908);
and U8083 (N_8083,N_6299,N_6078);
xnor U8084 (N_8084,N_6667,N_7672);
and U8085 (N_8085,N_6108,N_7014);
nor U8086 (N_8086,N_7727,N_7673);
and U8087 (N_8087,N_6783,N_6566);
or U8088 (N_8088,N_6683,N_7526);
nand U8089 (N_8089,N_7559,N_7090);
and U8090 (N_8090,N_6378,N_6881);
nor U8091 (N_8091,N_7775,N_7904);
and U8092 (N_8092,N_7358,N_6490);
xnor U8093 (N_8093,N_7648,N_6645);
xnor U8094 (N_8094,N_7499,N_6653);
or U8095 (N_8095,N_6470,N_7718);
nor U8096 (N_8096,N_6517,N_7475);
xnor U8097 (N_8097,N_6335,N_7293);
or U8098 (N_8098,N_7380,N_6682);
nand U8099 (N_8099,N_6484,N_6372);
nand U8100 (N_8100,N_6338,N_6437);
and U8101 (N_8101,N_7485,N_6670);
or U8102 (N_8102,N_7717,N_7969);
and U8103 (N_8103,N_6215,N_7001);
and U8104 (N_8104,N_7121,N_7598);
nand U8105 (N_8105,N_6355,N_7335);
and U8106 (N_8106,N_6963,N_6140);
xor U8107 (N_8107,N_7099,N_7871);
nand U8108 (N_8108,N_7960,N_7541);
and U8109 (N_8109,N_7926,N_6010);
or U8110 (N_8110,N_6544,N_6833);
or U8111 (N_8111,N_7140,N_6040);
nand U8112 (N_8112,N_6538,N_7206);
nand U8113 (N_8113,N_6777,N_7084);
xnor U8114 (N_8114,N_6272,N_7371);
and U8115 (N_8115,N_6890,N_7827);
and U8116 (N_8116,N_6804,N_7081);
nor U8117 (N_8117,N_7621,N_6615);
xnor U8118 (N_8118,N_7383,N_7311);
or U8119 (N_8119,N_7837,N_6240);
or U8120 (N_8120,N_7581,N_6443);
or U8121 (N_8121,N_7456,N_6268);
nor U8122 (N_8122,N_7253,N_6884);
nor U8123 (N_8123,N_6353,N_6560);
xnor U8124 (N_8124,N_7430,N_7505);
or U8125 (N_8125,N_6919,N_7935);
or U8126 (N_8126,N_6053,N_6706);
and U8127 (N_8127,N_6279,N_7560);
nor U8128 (N_8128,N_7836,N_7420);
and U8129 (N_8129,N_7025,N_6213);
or U8130 (N_8130,N_7828,N_6387);
or U8131 (N_8131,N_7962,N_7344);
xnor U8132 (N_8132,N_6988,N_7213);
nor U8133 (N_8133,N_6510,N_7154);
xnor U8134 (N_8134,N_6328,N_7534);
xnor U8135 (N_8135,N_6996,N_7998);
nor U8136 (N_8136,N_6147,N_6694);
or U8137 (N_8137,N_7947,N_7649);
or U8138 (N_8138,N_6636,N_7864);
nor U8139 (N_8139,N_6546,N_6370);
nor U8140 (N_8140,N_7186,N_6313);
nor U8141 (N_8141,N_6612,N_6605);
nand U8142 (N_8142,N_6839,N_6344);
or U8143 (N_8143,N_7602,N_7324);
xnor U8144 (N_8144,N_7569,N_6392);
or U8145 (N_8145,N_7891,N_7368);
or U8146 (N_8146,N_6730,N_6280);
or U8147 (N_8147,N_6169,N_7333);
xnor U8148 (N_8148,N_6453,N_6628);
and U8149 (N_8149,N_6698,N_7385);
and U8150 (N_8150,N_7571,N_6716);
xor U8151 (N_8151,N_6166,N_7991);
and U8152 (N_8152,N_6862,N_7896);
nor U8153 (N_8153,N_7751,N_6914);
xnor U8154 (N_8154,N_7282,N_6652);
nand U8155 (N_8155,N_7123,N_7857);
and U8156 (N_8156,N_6185,N_7493);
nand U8157 (N_8157,N_7866,N_6649);
and U8158 (N_8158,N_6432,N_7214);
nand U8159 (N_8159,N_6921,N_7670);
or U8160 (N_8160,N_6485,N_7172);
or U8161 (N_8161,N_6261,N_6941);
and U8162 (N_8162,N_7375,N_6635);
or U8163 (N_8163,N_6476,N_7779);
nor U8164 (N_8164,N_6427,N_7920);
nand U8165 (N_8165,N_6592,N_7799);
nand U8166 (N_8166,N_7409,N_7347);
or U8167 (N_8167,N_7317,N_7085);
or U8168 (N_8168,N_7049,N_7968);
xnor U8169 (N_8169,N_7390,N_6979);
nor U8170 (N_8170,N_6282,N_6002);
or U8171 (N_8171,N_6269,N_6130);
or U8172 (N_8172,N_7989,N_7013);
and U8173 (N_8173,N_7575,N_7017);
and U8174 (N_8174,N_6622,N_7147);
and U8175 (N_8175,N_6243,N_6015);
or U8176 (N_8176,N_6124,N_7296);
and U8177 (N_8177,N_7429,N_6527);
nand U8178 (N_8178,N_7281,N_6225);
nor U8179 (N_8179,N_7990,N_7018);
xor U8180 (N_8180,N_6115,N_6585);
nor U8181 (N_8181,N_6822,N_7111);
nor U8182 (N_8182,N_7848,N_7396);
nor U8183 (N_8183,N_6501,N_7563);
and U8184 (N_8184,N_6702,N_7788);
xor U8185 (N_8185,N_6324,N_7494);
or U8186 (N_8186,N_7381,N_6749);
nand U8187 (N_8187,N_7301,N_6188);
or U8188 (N_8188,N_7678,N_6664);
nor U8189 (N_8189,N_6109,N_6302);
xor U8190 (N_8190,N_6630,N_7635);
xnor U8191 (N_8191,N_6060,N_6720);
nand U8192 (N_8192,N_7416,N_6036);
nor U8193 (N_8193,N_7778,N_7468);
nand U8194 (N_8194,N_7167,N_7000);
and U8195 (N_8195,N_6295,N_7133);
or U8196 (N_8196,N_7441,N_6153);
nand U8197 (N_8197,N_6900,N_7425);
nand U8198 (N_8198,N_6383,N_6112);
xor U8199 (N_8199,N_6352,N_6699);
or U8200 (N_8200,N_7939,N_6047);
nand U8201 (N_8201,N_6791,N_7058);
nor U8202 (N_8202,N_7726,N_6850);
nand U8203 (N_8203,N_6314,N_7511);
nor U8204 (N_8204,N_6014,N_7961);
and U8205 (N_8205,N_6765,N_6257);
and U8206 (N_8206,N_6304,N_6766);
nor U8207 (N_8207,N_7700,N_7275);
xor U8208 (N_8208,N_6747,N_6677);
or U8209 (N_8209,N_6462,N_7184);
or U8210 (N_8210,N_7801,N_6512);
and U8211 (N_8211,N_6465,N_6985);
nor U8212 (N_8212,N_7764,N_6398);
nand U8213 (N_8213,N_6062,N_6461);
and U8214 (N_8214,N_6671,N_6906);
or U8215 (N_8215,N_7596,N_7162);
xor U8216 (N_8216,N_7048,N_6498);
nand U8217 (N_8217,N_7798,N_6315);
or U8218 (N_8218,N_7542,N_7374);
and U8219 (N_8219,N_7784,N_6537);
nand U8220 (N_8220,N_7752,N_6980);
nor U8221 (N_8221,N_6829,N_6399);
nor U8222 (N_8222,N_7417,N_6275);
and U8223 (N_8223,N_7254,N_7931);
or U8224 (N_8224,N_6928,N_6540);
nor U8225 (N_8225,N_7975,N_6633);
and U8226 (N_8226,N_7323,N_7644);
xnor U8227 (N_8227,N_7285,N_7040);
nor U8228 (N_8228,N_6144,N_6876);
xor U8229 (N_8229,N_6923,N_7087);
xnor U8230 (N_8230,N_6503,N_6475);
and U8231 (N_8231,N_6638,N_6669);
or U8232 (N_8232,N_7767,N_6696);
nand U8233 (N_8233,N_6323,N_7166);
nand U8234 (N_8234,N_7078,N_7508);
or U8235 (N_8235,N_7590,N_7587);
nor U8236 (N_8236,N_7124,N_7382);
xor U8237 (N_8237,N_6575,N_7356);
and U8238 (N_8238,N_6186,N_7062);
nand U8239 (N_8239,N_6569,N_6746);
xnor U8240 (N_8240,N_7039,N_6864);
nor U8241 (N_8241,N_7810,N_6588);
and U8242 (N_8242,N_7354,N_6818);
xnor U8243 (N_8243,N_6792,N_7704);
nand U8244 (N_8244,N_7580,N_7414);
nand U8245 (N_8245,N_6235,N_7620);
nand U8246 (N_8246,N_7258,N_6846);
nor U8247 (N_8247,N_7469,N_6254);
and U8248 (N_8248,N_7957,N_7811);
nand U8249 (N_8249,N_6369,N_6859);
nand U8250 (N_8250,N_6995,N_7540);
or U8251 (N_8251,N_6043,N_7209);
nor U8252 (N_8252,N_6386,N_7273);
xor U8253 (N_8253,N_7660,N_7854);
and U8254 (N_8254,N_6056,N_7797);
nor U8255 (N_8255,N_7309,N_7789);
and U8256 (N_8256,N_7431,N_6439);
or U8257 (N_8257,N_7755,N_6567);
nor U8258 (N_8258,N_7367,N_7965);
nand U8259 (N_8259,N_7045,N_7098);
xor U8260 (N_8260,N_7723,N_6438);
or U8261 (N_8261,N_6545,N_6477);
nor U8262 (N_8262,N_7632,N_7650);
xor U8263 (N_8263,N_7201,N_7225);
nand U8264 (N_8264,N_7447,N_6838);
xor U8265 (N_8265,N_6954,N_7230);
xnor U8266 (N_8266,N_7195,N_6899);
and U8267 (N_8267,N_6558,N_7473);
or U8268 (N_8268,N_7925,N_7052);
nand U8269 (N_8269,N_7370,N_7694);
and U8270 (N_8270,N_7365,N_7476);
nor U8271 (N_8271,N_7182,N_6578);
nor U8272 (N_8272,N_6896,N_6776);
xor U8273 (N_8273,N_6226,N_7963);
xnor U8274 (N_8274,N_7178,N_7086);
or U8275 (N_8275,N_7122,N_6561);
nand U8276 (N_8276,N_7608,N_6986);
and U8277 (N_8277,N_7146,N_6740);
and U8278 (N_8278,N_6486,N_6548);
and U8279 (N_8279,N_7967,N_7114);
nand U8280 (N_8280,N_6786,N_6916);
xnor U8281 (N_8281,N_7372,N_7002);
nand U8282 (N_8282,N_6155,N_7418);
or U8283 (N_8283,N_6371,N_7440);
xnor U8284 (N_8284,N_7988,N_6945);
nand U8285 (N_8285,N_7696,N_7405);
nand U8286 (N_8286,N_6469,N_6083);
xnor U8287 (N_8287,N_7046,N_7833);
nand U8288 (N_8288,N_6759,N_7710);
and U8289 (N_8289,N_7287,N_6431);
xor U8290 (N_8290,N_6423,N_7242);
or U8291 (N_8291,N_7248,N_7465);
or U8292 (N_8292,N_6031,N_6249);
or U8293 (N_8293,N_7738,N_7362);
or U8294 (N_8294,N_7645,N_6719);
nor U8295 (N_8295,N_7005,N_7319);
and U8296 (N_8296,N_6576,N_6606);
xnor U8297 (N_8297,N_7872,N_7748);
or U8298 (N_8298,N_7647,N_7408);
and U8299 (N_8299,N_6700,N_6368);
and U8300 (N_8300,N_7867,N_7132);
or U8301 (N_8301,N_7610,N_6672);
nand U8302 (N_8302,N_7224,N_7819);
nor U8303 (N_8303,N_7089,N_7633);
or U8304 (N_8304,N_7606,N_6200);
or U8305 (N_8305,N_7035,N_6528);
nand U8306 (N_8306,N_7237,N_6741);
nand U8307 (N_8307,N_7274,N_6289);
nor U8308 (N_8308,N_7830,N_6693);
or U8309 (N_8309,N_6726,N_6495);
and U8310 (N_8310,N_6970,N_6220);
nor U8311 (N_8311,N_7613,N_7011);
xor U8312 (N_8312,N_6563,N_6897);
nand U8313 (N_8313,N_6869,N_7502);
nand U8314 (N_8314,N_7812,N_7603);
or U8315 (N_8315,N_7906,N_7010);
or U8316 (N_8316,N_7392,N_6055);
nand U8317 (N_8317,N_6464,N_6400);
and U8318 (N_8318,N_7403,N_6711);
and U8319 (N_8319,N_7539,N_7655);
and U8320 (N_8320,N_7525,N_6070);
and U8321 (N_8321,N_6170,N_7774);
nand U8322 (N_8322,N_6136,N_6005);
nor U8323 (N_8323,N_7781,N_6831);
nor U8324 (N_8324,N_6904,N_7315);
nand U8325 (N_8325,N_7236,N_6487);
nor U8326 (N_8326,N_6404,N_7958);
xnor U8327 (N_8327,N_7160,N_6364);
nand U8328 (N_8328,N_7643,N_6889);
or U8329 (N_8329,N_6039,N_6595);
nand U8330 (N_8330,N_6874,N_7890);
nand U8331 (N_8331,N_6069,N_6953);
and U8332 (N_8332,N_7169,N_6074);
xnor U8333 (N_8333,N_7841,N_7853);
xor U8334 (N_8334,N_7294,N_7984);
xnor U8335 (N_8335,N_6625,N_6250);
and U8336 (N_8336,N_6163,N_6009);
and U8337 (N_8337,N_7923,N_6659);
nor U8338 (N_8338,N_7103,N_7264);
nand U8339 (N_8339,N_7067,N_6910);
or U8340 (N_8340,N_7060,N_7118);
xnor U8341 (N_8341,N_6772,N_7451);
xnor U8342 (N_8342,N_7638,N_6231);
xnor U8343 (N_8343,N_7221,N_6264);
or U8344 (N_8344,N_6046,N_7292);
and U8345 (N_8345,N_7152,N_7674);
nand U8346 (N_8346,N_7352,N_7604);
nand U8347 (N_8347,N_6968,N_6008);
and U8348 (N_8348,N_7577,N_6637);
or U8349 (N_8349,N_7459,N_7500);
and U8350 (N_8350,N_7936,N_7556);
and U8351 (N_8351,N_7956,N_6311);
xnor U8352 (N_8352,N_7846,N_6158);
and U8353 (N_8353,N_7743,N_6316);
or U8354 (N_8354,N_6514,N_7432);
and U8355 (N_8355,N_6027,N_7233);
and U8356 (N_8356,N_6866,N_7472);
or U8357 (N_8357,N_6781,N_7588);
nand U8358 (N_8358,N_6895,N_7676);
nor U8359 (N_8359,N_7145,N_6458);
or U8360 (N_8360,N_6455,N_7506);
nand U8361 (N_8361,N_6396,N_7803);
nand U8362 (N_8362,N_6126,N_6623);
or U8363 (N_8363,N_7265,N_7977);
nor U8364 (N_8364,N_7023,N_6661);
or U8365 (N_8365,N_6836,N_6680);
nor U8366 (N_8366,N_7343,N_6875);
nand U8367 (N_8367,N_7180,N_7599);
or U8368 (N_8368,N_7983,N_6138);
nor U8369 (N_8369,N_7657,N_6444);
or U8370 (N_8370,N_7422,N_6957);
nor U8371 (N_8371,N_7821,N_7745);
nor U8372 (N_8372,N_6173,N_6463);
nor U8373 (N_8373,N_7735,N_7646);
or U8374 (N_8374,N_7088,N_7291);
or U8375 (N_8375,N_6782,N_7339);
nand U8376 (N_8376,N_7814,N_7636);
nand U8377 (N_8377,N_7807,N_6419);
or U8378 (N_8378,N_7216,N_7820);
nand U8379 (N_8379,N_6382,N_6216);
and U8380 (N_8380,N_7030,N_7859);
xor U8381 (N_8381,N_7720,N_6291);
xor U8382 (N_8382,N_7079,N_7521);
nand U8383 (N_8383,N_7702,N_7379);
or U8384 (N_8384,N_7491,N_7028);
xor U8385 (N_8385,N_6882,N_6969);
or U8386 (N_8386,N_7458,N_7758);
nor U8387 (N_8387,N_7813,N_7567);
or U8388 (N_8388,N_6509,N_6381);
or U8389 (N_8389,N_6714,N_6978);
xor U8390 (N_8390,N_6739,N_6228);
or U8391 (N_8391,N_6021,N_6066);
nand U8392 (N_8392,N_6870,N_7877);
and U8393 (N_8393,N_6196,N_6184);
and U8394 (N_8394,N_6640,N_6194);
nand U8395 (N_8395,N_7398,N_6390);
and U8396 (N_8396,N_6843,N_6731);
xnor U8397 (N_8397,N_6327,N_7192);
and U8398 (N_8398,N_6948,N_7303);
nor U8399 (N_8399,N_7625,N_6918);
xnor U8400 (N_8400,N_6643,N_6832);
xnor U8401 (N_8401,N_7661,N_6245);
or U8402 (N_8402,N_7626,N_7047);
or U8403 (N_8403,N_7937,N_6408);
or U8404 (N_8404,N_7260,N_6019);
nand U8405 (N_8405,N_6888,N_6703);
nand U8406 (N_8406,N_6241,N_6004);
or U8407 (N_8407,N_7949,N_6613);
nor U8408 (N_8408,N_7349,N_7749);
xor U8409 (N_8409,N_6134,N_7982);
and U8410 (N_8410,N_7341,N_7822);
nand U8411 (N_8411,N_7056,N_6013);
or U8412 (N_8412,N_7113,N_7766);
xnor U8413 (N_8413,N_6445,N_6391);
nand U8414 (N_8414,N_6321,N_6655);
nand U8415 (N_8415,N_6413,N_6529);
nand U8416 (N_8416,N_6041,N_6908);
and U8417 (N_8417,N_6333,N_6814);
nor U8418 (N_8418,N_7695,N_7986);
nor U8419 (N_8419,N_6165,N_7955);
nand U8420 (N_8420,N_6262,N_6286);
nand U8421 (N_8421,N_7792,N_7689);
nor U8422 (N_8422,N_6000,N_6117);
nor U8423 (N_8423,N_6865,N_7389);
nand U8424 (N_8424,N_7662,N_7393);
xnor U8425 (N_8425,N_6405,N_6937);
and U8426 (N_8426,N_7104,N_6057);
nor U8427 (N_8427,N_7844,N_7318);
or U8428 (N_8428,N_6195,N_7536);
xnor U8429 (N_8429,N_7615,N_7915);
xor U8430 (N_8430,N_7164,N_7574);
xor U8431 (N_8431,N_7693,N_6096);
xor U8432 (N_8432,N_7747,N_6841);
and U8433 (N_8433,N_7868,N_7402);
nand U8434 (N_8434,N_6297,N_6679);
nand U8435 (N_8435,N_6306,N_7997);
or U8436 (N_8436,N_7641,N_7449);
and U8437 (N_8437,N_7483,N_6374);
nand U8438 (N_8438,N_6877,N_6692);
nand U8439 (N_8439,N_7435,N_7562);
nand U8440 (N_8440,N_6071,N_7460);
nor U8441 (N_8441,N_7816,N_6744);
and U8442 (N_8442,N_6522,N_6815);
nor U8443 (N_8443,N_7482,N_6849);
xnor U8444 (N_8444,N_7345,N_7815);
nand U8445 (N_8445,N_7021,N_6760);
nor U8446 (N_8446,N_6903,N_7307);
nand U8447 (N_8447,N_7019,N_7376);
xor U8448 (N_8448,N_6237,N_6085);
nand U8449 (N_8449,N_6925,N_7746);
and U8450 (N_8450,N_6030,N_6505);
xnor U8451 (N_8451,N_7218,N_6796);
or U8452 (N_8452,N_7407,N_6054);
or U8453 (N_8453,N_7091,N_6975);
nand U8454 (N_8454,N_6705,N_7825);
or U8455 (N_8455,N_6729,N_6813);
and U8456 (N_8456,N_6580,N_7457);
nand U8457 (N_8457,N_6583,N_6913);
and U8458 (N_8458,N_6617,N_7940);
nand U8459 (N_8459,N_6830,N_6139);
nor U8460 (N_8460,N_6511,N_7546);
and U8461 (N_8461,N_7442,N_6375);
nand U8462 (N_8462,N_7994,N_6212);
xor U8463 (N_8463,N_6748,N_6806);
or U8464 (N_8464,N_7041,N_6964);
nor U8465 (N_8465,N_6265,N_6406);
nor U8466 (N_8466,N_6065,N_7314);
xnor U8467 (N_8467,N_7597,N_6536);
or U8468 (N_8468,N_6255,N_6539);
and U8469 (N_8469,N_7589,N_7034);
nor U8470 (N_8470,N_7721,N_6556);
or U8471 (N_8471,N_6557,N_7576);
and U8472 (N_8472,N_6417,N_7437);
and U8473 (N_8473,N_7929,N_6500);
nor U8474 (N_8474,N_7913,N_7675);
or U8475 (N_8475,N_7032,N_7304);
nor U8476 (N_8476,N_6320,N_6780);
nor U8477 (N_8477,N_6076,N_6482);
nor U8478 (N_8478,N_7850,N_6525);
xnor U8479 (N_8479,N_7255,N_6981);
or U8480 (N_8480,N_6210,N_7707);
xor U8481 (N_8481,N_7072,N_6542);
nor U8482 (N_8482,N_6835,N_6393);
nor U8483 (N_8483,N_6614,N_7252);
nor U8484 (N_8484,N_6436,N_6707);
or U8485 (N_8485,N_7763,N_7061);
and U8486 (N_8486,N_6142,N_7634);
nor U8487 (N_8487,N_6329,N_6803);
nor U8488 (N_8488,N_7557,N_6950);
nand U8489 (N_8489,N_6414,N_6757);
and U8490 (N_8490,N_7719,N_6502);
nor U8491 (N_8491,N_6524,N_6411);
nor U8492 (N_8492,N_6853,N_6801);
nand U8493 (N_8493,N_7870,N_7731);
or U8494 (N_8494,N_6590,N_6581);
nand U8495 (N_8495,N_6026,N_7584);
xnor U8496 (N_8496,N_7100,N_7223);
xor U8497 (N_8497,N_7858,N_6127);
nor U8498 (N_8498,N_6206,N_6296);
and U8499 (N_8499,N_7847,N_7461);
and U8500 (N_8500,N_6363,N_7455);
nand U8501 (N_8501,N_6564,N_7009);
nor U8502 (N_8502,N_7619,N_7845);
xnor U8503 (N_8503,N_6449,N_7630);
nor U8504 (N_8504,N_7985,N_6506);
nor U8505 (N_8505,N_6293,N_6025);
nand U8506 (N_8506,N_6307,N_6952);
nand U8507 (N_8507,N_6167,N_7185);
or U8508 (N_8508,N_7951,N_6562);
nor U8509 (N_8509,N_6943,N_7733);
or U8510 (N_8510,N_6029,N_7016);
xor U8511 (N_8511,N_7210,N_6191);
and U8512 (N_8512,N_6994,N_6067);
nor U8513 (N_8513,N_7183,N_7302);
xor U8514 (N_8514,N_6099,N_7736);
nor U8515 (N_8515,N_7912,N_7427);
or U8516 (N_8516,N_7112,N_6883);
and U8517 (N_8517,N_6708,N_6892);
or U8518 (N_8518,N_7107,N_6385);
nor U8519 (N_8519,N_7863,N_6602);
xnor U8520 (N_8520,N_6110,N_6086);
or U8521 (N_8521,N_7471,N_6174);
and U8522 (N_8522,N_6122,N_6657);
nor U8523 (N_8523,N_6586,N_6073);
nand U8524 (N_8524,N_6798,N_6035);
or U8525 (N_8525,N_6162,N_7537);
or U8526 (N_8526,N_7840,N_6519);
or U8527 (N_8527,N_6450,N_7498);
nand U8528 (N_8528,N_7391,N_7517);
nand U8529 (N_8529,N_7512,N_7808);
or U8530 (N_8530,N_7806,N_7108);
and U8531 (N_8531,N_7609,N_6294);
nor U8532 (N_8532,N_6011,N_7703);
xnor U8533 (N_8533,N_6724,N_6424);
nand U8534 (N_8534,N_6935,N_7346);
nand U8535 (N_8535,N_6591,N_6104);
and U8536 (N_8536,N_7369,N_6769);
nand U8537 (N_8537,N_7691,N_7579);
and U8538 (N_8538,N_6609,N_7478);
nand U8539 (N_8539,N_7305,N_6395);
nor U8540 (N_8540,N_7623,N_7922);
or U8541 (N_8541,N_6440,N_7793);
nor U8542 (N_8542,N_6492,N_7235);
nor U8543 (N_8543,N_6365,N_7943);
xnor U8544 (N_8544,N_6872,N_7914);
and U8545 (N_8545,N_7151,N_7092);
and U8546 (N_8546,N_7757,N_6459);
and U8547 (N_8547,N_6644,N_6001);
nor U8548 (N_8548,N_6755,N_6422);
xnor U8549 (N_8549,N_6825,N_6513);
nor U8550 (N_8550,N_6958,N_7289);
xnor U8551 (N_8551,N_7682,N_7203);
or U8552 (N_8552,N_6331,N_7971);
and U8553 (N_8553,N_6712,N_6050);
nor U8554 (N_8554,N_7071,N_6263);
and U8555 (N_8555,N_7095,N_6878);
or U8556 (N_8556,N_7688,N_7593);
xnor U8557 (N_8557,N_6159,N_7669);
and U8558 (N_8558,N_7783,N_7578);
nor U8559 (N_8559,N_6577,N_6735);
nand U8560 (N_8560,N_6128,N_7794);
or U8561 (N_8561,N_6301,N_6193);
or U8562 (N_8562,N_7353,N_7462);
or U8563 (N_8563,N_7637,N_7917);
nand U8564 (N_8564,N_6497,N_6971);
nand U8565 (N_8565,N_7042,N_6753);
nor U8566 (N_8566,N_7777,N_6626);
xnor U8567 (N_8567,N_6654,N_7741);
nand U8568 (N_8568,N_7681,N_7229);
nand U8569 (N_8569,N_6627,N_7600);
nand U8570 (N_8570,N_7568,N_6389);
xnor U8571 (N_8571,N_7805,N_6176);
xor U8572 (N_8572,N_7851,N_6619);
nor U8573 (N_8573,N_6348,N_6550);
and U8574 (N_8574,N_6733,N_6152);
or U8575 (N_8575,N_7729,N_6118);
or U8576 (N_8576,N_7320,N_6533);
nand U8577 (N_8577,N_6181,N_7954);
and U8578 (N_8578,N_7905,N_6603);
nor U8579 (N_8579,N_7787,N_6885);
nor U8580 (N_8580,N_6559,N_7330);
xor U8581 (N_8581,N_6285,N_7874);
or U8582 (N_8582,N_7993,N_6190);
nand U8583 (N_8583,N_7439,N_7933);
nor U8584 (N_8584,N_6534,N_7119);
nand U8585 (N_8585,N_6929,N_7444);
xor U8586 (N_8586,N_7910,N_7428);
nor U8587 (N_8587,N_7549,N_7900);
or U8588 (N_8588,N_6758,N_7181);
nand U8589 (N_8589,N_7290,N_6721);
nor U8590 (N_8590,N_7668,N_7515);
nand U8591 (N_8591,N_6624,N_7279);
or U8592 (N_8592,N_7448,N_7187);
nand U8593 (N_8593,N_7008,N_6998);
xnor U8594 (N_8594,N_7168,N_7776);
nand U8595 (N_8595,N_7796,N_6102);
xnor U8596 (N_8596,N_6646,N_7855);
or U8597 (N_8597,N_6632,N_6817);
nand U8598 (N_8598,N_7366,N_7271);
or U8599 (N_8599,N_6982,N_7135);
and U8600 (N_8600,N_6662,N_7327);
or U8601 (N_8601,N_7831,N_7873);
and U8602 (N_8602,N_7463,N_6725);
nor U8603 (N_8603,N_6068,N_6508);
and U8604 (N_8604,N_6778,N_7927);
nor U8605 (N_8605,N_6499,N_6133);
nor U8606 (N_8606,N_7126,N_7244);
xnor U8607 (N_8607,N_6666,N_7329);
nand U8608 (N_8608,N_6023,N_7809);
and U8609 (N_8609,N_7227,N_7211);
nand U8610 (N_8610,N_7004,N_7143);
and U8611 (N_8611,N_6038,N_7879);
nor U8612 (N_8612,N_7839,N_7156);
or U8613 (N_8613,N_6570,N_6734);
and U8614 (N_8614,N_6164,N_6361);
nand U8615 (N_8615,N_6907,N_6687);
nand U8616 (N_8616,N_6977,N_7708);
and U8617 (N_8617,N_6281,N_7903);
or U8618 (N_8618,N_6198,N_7823);
nor U8619 (N_8619,N_6252,N_7538);
or U8620 (N_8620,N_7742,N_7438);
nand U8621 (N_8621,N_7328,N_6081);
xnor U8622 (N_8622,N_7053,N_6873);
and U8623 (N_8623,N_7007,N_7363);
or U8624 (N_8624,N_6790,N_7768);
nor U8625 (N_8625,N_6468,N_7531);
or U8626 (N_8626,N_6397,N_7734);
nor U8627 (N_8627,N_7131,N_7680);
or U8628 (N_8628,N_6345,N_6349);
and U8629 (N_8629,N_7247,N_6143);
and U8630 (N_8630,N_6648,N_7205);
nand U8631 (N_8631,N_6531,N_6905);
or U8632 (N_8632,N_7523,N_7208);
or U8633 (N_8633,N_6336,N_6132);
xnor U8634 (N_8634,N_7946,N_6826);
nor U8635 (N_8635,N_7753,N_7885);
xor U8636 (N_8636,N_7665,N_7860);
xor U8637 (N_8637,N_7212,N_6723);
nor U8638 (N_8638,N_7406,N_6879);
or U8639 (N_8639,N_7504,N_7486);
or U8640 (N_8640,N_7130,N_6805);
nor U8641 (N_8641,N_6059,N_7878);
nand U8642 (N_8642,N_7893,N_6808);
nor U8643 (N_8643,N_6227,N_7194);
nand U8644 (N_8644,N_6845,N_6474);
or U8645 (N_8645,N_7155,N_7012);
nand U8646 (N_8646,N_7980,N_6160);
or U8647 (N_8647,N_7261,N_6774);
nor U8648 (N_8648,N_7892,N_6660);
nand U8649 (N_8649,N_7532,N_6812);
or U8650 (N_8650,N_6416,N_7529);
xor U8651 (N_8651,N_7677,N_7786);
nor U8652 (N_8652,N_6718,N_6446);
or U8653 (N_8653,N_6420,N_7898);
or U8654 (N_8654,N_7683,N_6634);
nand U8655 (N_8655,N_7516,N_6251);
or U8656 (N_8656,N_6489,N_6203);
or U8657 (N_8657,N_6218,N_6430);
xor U8658 (N_8658,N_7953,N_6488);
and U8659 (N_8659,N_7800,N_6871);
and U8660 (N_8660,N_6032,N_6433);
or U8661 (N_8661,N_6787,N_7919);
and U8662 (N_8662,N_7631,N_6715);
xnor U8663 (N_8663,N_7232,N_6287);
and U8664 (N_8664,N_7082,N_6105);
xnor U8665 (N_8665,N_6171,N_7566);
nor U8666 (N_8666,N_7101,N_6217);
or U8667 (N_8667,N_6290,N_6880);
or U8668 (N_8668,N_7074,N_6574);
and U8669 (N_8669,N_6111,N_7642);
nor U8670 (N_8670,N_7583,N_7501);
nor U8671 (N_8671,N_7730,N_6042);
or U8672 (N_8672,N_6274,N_7137);
or U8673 (N_8673,N_7544,N_7412);
or U8674 (N_8674,N_7276,N_6754);
xor U8675 (N_8675,N_7607,N_7692);
or U8676 (N_8676,N_6902,N_7782);
nor U8677 (N_8677,N_7732,N_7340);
nand U8678 (N_8678,N_7163,N_6061);
and U8679 (N_8679,N_6141,N_7654);
nor U8680 (N_8680,N_6938,N_7785);
and U8681 (N_8681,N_7740,N_7503);
nor U8682 (N_8682,N_7373,N_7802);
xnor U8683 (N_8683,N_7728,N_7959);
and U8684 (N_8684,N_6410,N_6553);
xnor U8685 (N_8685,N_7686,N_7322);
or U8686 (N_8686,N_7179,N_7193);
nand U8687 (N_8687,N_6418,N_7175);
nand U8688 (N_8688,N_7266,N_6959);
or U8689 (N_8689,N_6891,N_6867);
nand U8690 (N_8690,N_7513,N_7605);
nor U8691 (N_8691,N_6017,N_7945);
or U8692 (N_8692,N_7278,N_7818);
or U8693 (N_8693,N_6926,N_6415);
or U8694 (N_8694,N_7725,N_6121);
nand U8695 (N_8695,N_7941,N_6854);
and U8696 (N_8696,N_6594,N_7780);
xnor U8697 (N_8697,N_7932,N_7530);
nor U8698 (N_8698,N_7228,N_6611);
nand U8699 (N_8699,N_6816,N_6337);
nor U8700 (N_8700,N_6616,N_6394);
nor U8701 (N_8701,N_7591,N_7054);
nor U8702 (N_8702,N_7762,N_7551);
xor U8703 (N_8703,N_7076,N_6827);
nor U8704 (N_8704,N_7217,N_6182);
xnor U8705 (N_8705,N_6837,N_6761);
nand U8706 (N_8706,N_7127,N_7966);
xnor U8707 (N_8707,N_7445,N_7548);
xnor U8708 (N_8708,N_7907,N_7177);
nand U8709 (N_8709,N_7300,N_6598);
nor U8710 (N_8710,N_6359,N_6949);
xnor U8711 (N_8711,N_7332,N_6599);
or U8712 (N_8712,N_6593,N_7357);
or U8713 (N_8713,N_6601,N_6855);
or U8714 (N_8714,N_7191,N_6684);
nand U8715 (N_8715,N_7066,N_6927);
nand U8716 (N_8716,N_7083,N_7765);
and U8717 (N_8717,N_7378,N_6481);
or U8718 (N_8718,N_7570,N_7895);
nor U8719 (N_8719,N_6491,N_6496);
and U8720 (N_8720,N_6175,N_6911);
nand U8721 (N_8721,N_6253,N_6852);
nor U8722 (N_8722,N_7518,N_6442);
and U8723 (N_8723,N_7308,N_7150);
or U8724 (N_8724,N_7653,N_6589);
or U8725 (N_8725,N_6441,N_7934);
and U8726 (N_8726,N_6515,N_7243);
nand U8727 (N_8727,N_6097,N_6189);
or U8728 (N_8728,N_6743,N_7769);
nor U8729 (N_8729,N_6756,N_6917);
xnor U8730 (N_8730,N_6341,N_6360);
nand U8731 (N_8731,N_6283,N_6728);
nand U8732 (N_8732,N_6230,N_7176);
nand U8733 (N_8733,N_7699,N_6868);
or U8734 (N_8734,N_7601,N_6965);
nor U8735 (N_8735,N_7651,N_6993);
nand U8736 (N_8736,N_7097,N_7404);
and U8737 (N_8737,N_7246,N_6084);
or U8738 (N_8738,N_7286,N_7106);
nand U8739 (N_8739,N_7159,N_7972);
or U8740 (N_8740,N_7902,N_6123);
nand U8741 (N_8741,N_6149,N_7849);
and U8742 (N_8742,N_6673,N_7618);
nand U8743 (N_8743,N_7899,N_7930);
and U8744 (N_8744,N_7865,N_7999);
or U8745 (N_8745,N_6732,N_6332);
nor U8746 (N_8746,N_6072,N_7887);
and U8747 (N_8747,N_7948,N_7477);
or U8748 (N_8748,N_6930,N_6309);
or U8749 (N_8749,N_7886,N_6119);
nor U8750 (N_8750,N_7533,N_7269);
nor U8751 (N_8751,N_7288,N_7622);
and U8752 (N_8752,N_6992,N_7141);
nor U8753 (N_8753,N_7697,N_6197);
and U8754 (N_8754,N_6270,N_7219);
nor U8755 (N_8755,N_6379,N_7015);
and U8756 (N_8756,N_7055,N_6401);
and U8757 (N_8757,N_6095,N_7701);
xor U8758 (N_8758,N_7284,N_7249);
nor U8759 (N_8759,N_6428,N_7558);
xor U8760 (N_8760,N_6120,N_6607);
nor U8761 (N_8761,N_7553,N_6604);
nand U8762 (N_8762,N_7750,N_6997);
and U8763 (N_8763,N_7038,N_6775);
nor U8764 (N_8764,N_7944,N_6678);
nor U8765 (N_8765,N_7950,N_7519);
xor U8766 (N_8766,N_7337,N_6087);
or U8767 (N_8767,N_6292,N_7384);
nand U8768 (N_8768,N_7804,N_6942);
xnor U8769 (N_8769,N_6350,N_6022);
or U8770 (N_8770,N_6367,N_7453);
nand U8771 (N_8771,N_6233,N_6342);
or U8772 (N_8772,N_7334,N_6794);
nor U8773 (N_8773,N_6582,N_7897);
nand U8774 (N_8774,N_6310,N_6052);
xor U8775 (N_8775,N_7360,N_7202);
nor U8776 (N_8776,N_6701,N_7628);
or U8777 (N_8777,N_6058,N_7880);
xor U8778 (N_8778,N_6088,N_7835);
or U8779 (N_8779,N_6131,N_7388);
nand U8780 (N_8780,N_6211,N_6223);
and U8781 (N_8781,N_6238,N_6471);
and U8782 (N_8782,N_7020,N_7283);
or U8783 (N_8783,N_6955,N_7894);
or U8784 (N_8784,N_7148,N_7627);
or U8785 (N_8785,N_6717,N_7884);
xnor U8786 (N_8786,N_7022,N_7006);
and U8787 (N_8787,N_7852,N_6709);
or U8788 (N_8788,N_6208,N_7756);
or U8789 (N_8789,N_7359,N_7144);
xnor U8790 (N_8790,N_6114,N_6802);
or U8791 (N_8791,N_7454,N_7262);
xor U8792 (N_8792,N_6961,N_6939);
nand U8793 (N_8793,N_6915,N_6454);
and U8794 (N_8794,N_7987,N_6045);
nand U8795 (N_8795,N_6460,N_6221);
nand U8796 (N_8796,N_7973,N_7068);
and U8797 (N_8797,N_7434,N_7096);
xor U8798 (N_8798,N_6412,N_7773);
nor U8799 (N_8799,N_6276,N_6799);
and U8800 (N_8800,N_6113,N_6180);
nand U8801 (N_8801,N_6049,N_6077);
and U8802 (N_8802,N_7759,N_6676);
xor U8803 (N_8803,N_6156,N_7881);
nand U8804 (N_8804,N_7709,N_6931);
nand U8805 (N_8805,N_6811,N_6447);
nand U8806 (N_8806,N_6695,N_6722);
nor U8807 (N_8807,N_7510,N_6745);
or U8808 (N_8808,N_6356,N_6573);
and U8809 (N_8809,N_6172,N_7250);
nor U8810 (N_8810,N_7639,N_7490);
nor U8811 (N_8811,N_6376,N_7555);
nor U8812 (N_8812,N_7497,N_6668);
and U8813 (N_8813,N_6650,N_7364);
or U8814 (N_8814,N_6554,N_7528);
xor U8815 (N_8815,N_7481,N_7464);
xor U8816 (N_8816,N_6847,N_7685);
xor U8817 (N_8817,N_6247,N_7105);
nor U8818 (N_8818,N_6028,N_6256);
xor U8819 (N_8819,N_7624,N_7450);
and U8820 (N_8820,N_6547,N_7706);
xor U8821 (N_8821,N_6820,N_7489);
nor U8822 (N_8822,N_6984,N_7916);
or U8823 (N_8823,N_6354,N_6860);
or U8824 (N_8824,N_7713,N_7739);
or U8825 (N_8825,N_7350,N_7080);
and U8826 (N_8826,N_7861,N_7595);
and U8827 (N_8827,N_6168,N_7466);
nor U8828 (N_8828,N_6148,N_6305);
nor U8829 (N_8829,N_7484,N_6242);
nor U8830 (N_8830,N_6137,N_6857);
nor U8831 (N_8831,N_7129,N_7306);
nand U8832 (N_8832,N_6317,N_6863);
nor U8833 (N_8833,N_6020,N_7889);
xnor U8834 (N_8834,N_7547,N_7207);
nand U8835 (N_8835,N_6819,N_7514);
xnor U8836 (N_8836,N_6834,N_6248);
or U8837 (N_8837,N_6956,N_7399);
xor U8838 (N_8838,N_6674,N_6518);
xnor U8839 (N_8839,N_6473,N_7705);
nand U8840 (N_8840,N_7565,N_6541);
xor U8841 (N_8841,N_7419,N_7918);
and U8842 (N_8842,N_7698,N_6691);
xor U8843 (N_8843,N_7509,N_6178);
or U8844 (N_8844,N_7687,N_7348);
and U8845 (N_8845,N_6303,N_7978);
and U8846 (N_8846,N_7158,N_7196);
nand U8847 (N_8847,N_6003,N_6974);
nor U8848 (N_8848,N_6044,N_7198);
and U8849 (N_8849,N_7862,N_7772);
or U8850 (N_8850,N_6258,N_6224);
xnor U8851 (N_8851,N_6618,N_6532);
nor U8852 (N_8852,N_7522,N_7336);
xnor U8853 (N_8853,N_6504,N_7197);
nand U8854 (N_8854,N_7171,N_6107);
nand U8855 (N_8855,N_6101,N_6663);
and U8856 (N_8856,N_6568,N_6689);
nand U8857 (N_8857,N_6407,N_6523);
and U8858 (N_8858,N_6346,N_6103);
nor U8859 (N_8859,N_6308,N_6064);
nand U8860 (N_8860,N_6179,N_7970);
nand U8861 (N_8861,N_6967,N_6893);
nor U8862 (N_8862,N_7065,N_7263);
or U8863 (N_8863,N_7433,N_6771);
xnor U8864 (N_8864,N_7976,N_6284);
nand U8865 (N_8865,N_6157,N_7234);
or U8866 (N_8866,N_6713,N_7952);
nand U8867 (N_8867,N_6651,N_7724);
xor U8868 (N_8868,N_7394,N_7325);
and U8869 (N_8869,N_6037,N_7342);
nand U8870 (N_8870,N_6034,N_6770);
nand U8871 (N_8871,N_6421,N_6151);
xor U8872 (N_8872,N_7220,N_6199);
or U8873 (N_8873,N_6079,N_6456);
or U8874 (N_8874,N_6526,N_6552);
nor U8875 (N_8875,N_7791,N_7077);
nand U8876 (N_8876,N_6266,N_7832);
nor U8877 (N_8877,N_6762,N_7684);
nand U8878 (N_8878,N_7415,N_6989);
and U8879 (N_8879,N_6800,N_6373);
nand U8880 (N_8880,N_7277,N_6452);
nor U8881 (N_8881,N_6326,N_6543);
nand U8882 (N_8882,N_7964,N_7760);
nor U8883 (N_8883,N_7834,N_7188);
or U8884 (N_8884,N_6016,N_6259);
nor U8885 (N_8885,N_7883,N_6768);
or U8886 (N_8886,N_6007,N_7520);
and U8887 (N_8887,N_7173,N_6048);
and U8888 (N_8888,N_7824,N_7189);
nand U8889 (N_8889,N_7652,N_7073);
nor U8890 (N_8890,N_6033,N_6697);
xor U8891 (N_8891,N_6177,N_6951);
or U8892 (N_8892,N_6571,N_6187);
and U8893 (N_8893,N_7270,N_6347);
and U8894 (N_8894,N_6325,N_6629);
and U8895 (N_8895,N_7992,N_6106);
and U8896 (N_8896,N_6793,N_7995);
and U8897 (N_8897,N_6990,N_7875);
or U8898 (N_8898,N_6201,N_6267);
nor U8899 (N_8899,N_6466,N_6894);
and U8900 (N_8900,N_7492,N_6823);
xor U8901 (N_8901,N_6940,N_7938);
nor U8902 (N_8902,N_6222,N_6448);
nand U8903 (N_8903,N_7467,N_6100);
or U8904 (N_8904,N_6752,N_6232);
and U8905 (N_8905,N_6535,N_6991);
and U8906 (N_8906,N_7222,N_7026);
nand U8907 (N_8907,N_7443,N_7321);
nand U8908 (N_8908,N_6204,N_6960);
and U8909 (N_8909,N_7856,N_6339);
nand U8910 (N_8910,N_7452,N_6621);
and U8911 (N_8911,N_7355,N_6472);
xnor U8912 (N_8912,N_6933,N_7714);
nand U8913 (N_8913,N_6727,N_7901);
or U8914 (N_8914,N_6012,N_7268);
and U8915 (N_8915,N_7240,N_6856);
or U8916 (N_8916,N_6334,N_6579);
or U8917 (N_8917,N_7215,N_6797);
xnor U8918 (N_8918,N_6642,N_6824);
and U8919 (N_8919,N_6192,N_7351);
and U8920 (N_8920,N_7395,N_7617);
and U8921 (N_8921,N_6318,N_6366);
nand U8922 (N_8922,N_7770,N_6384);
nand U8923 (N_8923,N_7027,N_6840);
nor U8924 (N_8924,N_7256,N_7479);
nor U8925 (N_8925,N_7397,N_7064);
or U8926 (N_8926,N_6795,N_7656);
nand U8927 (N_8927,N_7031,N_6478);
and U8928 (N_8928,N_6639,N_6788);
nand U8929 (N_8929,N_7316,N_6098);
and U8930 (N_8930,N_6135,N_6273);
xor U8931 (N_8931,N_6597,N_6214);
nor U8932 (N_8932,N_6656,N_7128);
xnor U8933 (N_8933,N_6750,N_6973);
and U8934 (N_8934,N_6600,N_7411);
xnor U8935 (N_8935,N_6234,N_7033);
nand U8936 (N_8936,N_7594,N_6584);
xnor U8937 (N_8937,N_7921,N_6312);
nand U8938 (N_8938,N_6377,N_7377);
nand U8939 (N_8939,N_7117,N_6205);
xor U8940 (N_8940,N_7715,N_7326);
nor U8941 (N_8941,N_6690,N_7057);
or U8942 (N_8942,N_6675,N_6987);
nand U8943 (N_8943,N_6425,N_6209);
xor U8944 (N_8944,N_6357,N_7679);
and U8945 (N_8945,N_6434,N_7029);
nand U8946 (N_8946,N_7572,N_7199);
or U8947 (N_8947,N_6236,N_6244);
and U8948 (N_8948,N_7070,N_6704);
nand U8949 (N_8949,N_6516,N_6520);
or U8950 (N_8950,N_6246,N_7446);
and U8951 (N_8951,N_6596,N_6343);
xor U8952 (N_8952,N_6736,N_7611);
nand U8953 (N_8953,N_6934,N_6810);
or U8954 (N_8954,N_6129,N_6681);
nor U8955 (N_8955,N_7116,N_6483);
nand U8956 (N_8956,N_6686,N_7037);
nor U8957 (N_8957,N_6710,N_7436);
xor U8958 (N_8958,N_7586,N_6380);
nand U8959 (N_8959,N_7102,N_6858);
and U8960 (N_8960,N_7125,N_7153);
nand U8961 (N_8961,N_7838,N_6887);
nand U8962 (N_8962,N_7712,N_7231);
xnor U8963 (N_8963,N_6125,N_6089);
or U8964 (N_8964,N_6093,N_6608);
xor U8965 (N_8965,N_6773,N_6358);
xnor U8966 (N_8966,N_6300,N_7050);
nor U8967 (N_8967,N_6091,N_7298);
xor U8968 (N_8968,N_6094,N_6402);
and U8969 (N_8969,N_7790,N_7582);
or U8970 (N_8970,N_6972,N_6555);
nor U8971 (N_8971,N_7204,N_7527);
and U8972 (N_8972,N_7138,N_6901);
and U8973 (N_8973,N_7036,N_6154);
xnor U8974 (N_8974,N_7942,N_7241);
and U8975 (N_8975,N_7761,N_7996);
or U8976 (N_8976,N_6886,N_7226);
nand U8977 (N_8977,N_6467,N_6521);
and U8978 (N_8978,N_7413,N_6063);
and U8979 (N_8979,N_7239,N_6779);
nand U8980 (N_8980,N_7093,N_7488);
nor U8981 (N_8981,N_7487,N_6962);
xnor U8982 (N_8982,N_6976,N_7259);
xnor U8983 (N_8983,N_7170,N_6807);
or U8984 (N_8984,N_6620,N_7386);
or U8985 (N_8985,N_7257,N_7667);
xnor U8986 (N_8986,N_7843,N_7573);
nand U8987 (N_8987,N_6507,N_6966);
nand U8988 (N_8988,N_7690,N_7495);
and U8989 (N_8989,N_6983,N_7238);
and U8990 (N_8990,N_7190,N_6851);
nor U8991 (N_8991,N_7272,N_6785);
nor U8992 (N_8992,N_7421,N_6075);
nand U8993 (N_8993,N_7139,N_7882);
and U8994 (N_8994,N_7614,N_7338);
nor U8995 (N_8995,N_6641,N_7507);
nand U8996 (N_8996,N_7161,N_7410);
nand U8997 (N_8997,N_6844,N_7136);
nor U8998 (N_8998,N_7423,N_7629);
and U8999 (N_8999,N_7044,N_6494);
nand U9000 (N_9000,N_6757,N_6217);
nor U9001 (N_9001,N_7262,N_6362);
xor U9002 (N_9002,N_6429,N_7315);
or U9003 (N_9003,N_6460,N_6072);
or U9004 (N_9004,N_7634,N_7158);
or U9005 (N_9005,N_6467,N_6076);
nand U9006 (N_9006,N_7904,N_7169);
or U9007 (N_9007,N_7834,N_7343);
or U9008 (N_9008,N_6097,N_7721);
xnor U9009 (N_9009,N_6287,N_7677);
and U9010 (N_9010,N_7789,N_6881);
nand U9011 (N_9011,N_7036,N_7102);
and U9012 (N_9012,N_7221,N_7942);
or U9013 (N_9013,N_7454,N_7014);
nor U9014 (N_9014,N_7273,N_6211);
nand U9015 (N_9015,N_7225,N_7410);
and U9016 (N_9016,N_6884,N_6576);
or U9017 (N_9017,N_7229,N_7588);
or U9018 (N_9018,N_6037,N_6425);
and U9019 (N_9019,N_6336,N_7479);
nor U9020 (N_9020,N_6422,N_6883);
and U9021 (N_9021,N_6866,N_6707);
or U9022 (N_9022,N_6762,N_7492);
nor U9023 (N_9023,N_7150,N_7120);
nand U9024 (N_9024,N_6963,N_7922);
nand U9025 (N_9025,N_6881,N_7980);
and U9026 (N_9026,N_7903,N_7931);
xnor U9027 (N_9027,N_6773,N_7758);
xnor U9028 (N_9028,N_7710,N_7758);
or U9029 (N_9029,N_7725,N_7881);
nand U9030 (N_9030,N_7089,N_7709);
nor U9031 (N_9031,N_7771,N_6212);
nand U9032 (N_9032,N_7367,N_7420);
and U9033 (N_9033,N_6572,N_7400);
nand U9034 (N_9034,N_6524,N_6161);
xor U9035 (N_9035,N_7247,N_7675);
and U9036 (N_9036,N_6560,N_6036);
nor U9037 (N_9037,N_7985,N_6072);
nand U9038 (N_9038,N_6755,N_7721);
or U9039 (N_9039,N_7589,N_6475);
nor U9040 (N_9040,N_7537,N_6691);
and U9041 (N_9041,N_7442,N_6026);
xnor U9042 (N_9042,N_6174,N_7269);
nand U9043 (N_9043,N_7588,N_6563);
nand U9044 (N_9044,N_7073,N_7090);
and U9045 (N_9045,N_6483,N_7332);
and U9046 (N_9046,N_7344,N_6272);
nand U9047 (N_9047,N_6867,N_6323);
xnor U9048 (N_9048,N_7900,N_7300);
nand U9049 (N_9049,N_6654,N_6143);
nand U9050 (N_9050,N_6881,N_6118);
nand U9051 (N_9051,N_6331,N_7378);
nand U9052 (N_9052,N_6951,N_6157);
xor U9053 (N_9053,N_6490,N_6820);
nand U9054 (N_9054,N_7228,N_7852);
xnor U9055 (N_9055,N_7256,N_6882);
nand U9056 (N_9056,N_7317,N_7230);
and U9057 (N_9057,N_7586,N_6412);
nor U9058 (N_9058,N_6176,N_6319);
or U9059 (N_9059,N_6782,N_7970);
nand U9060 (N_9060,N_7489,N_7866);
nand U9061 (N_9061,N_7976,N_7769);
xnor U9062 (N_9062,N_6565,N_6715);
and U9063 (N_9063,N_6841,N_7592);
nand U9064 (N_9064,N_7324,N_6140);
and U9065 (N_9065,N_6254,N_7838);
xnor U9066 (N_9066,N_7953,N_6546);
xor U9067 (N_9067,N_6282,N_7572);
or U9068 (N_9068,N_7783,N_7895);
nand U9069 (N_9069,N_7274,N_7968);
and U9070 (N_9070,N_7346,N_7696);
xnor U9071 (N_9071,N_6836,N_6755);
nand U9072 (N_9072,N_6861,N_7839);
and U9073 (N_9073,N_6951,N_7001);
and U9074 (N_9074,N_7942,N_6020);
nand U9075 (N_9075,N_6675,N_7934);
or U9076 (N_9076,N_6590,N_6907);
nor U9077 (N_9077,N_6186,N_6064);
nor U9078 (N_9078,N_7611,N_7082);
and U9079 (N_9079,N_6744,N_6922);
and U9080 (N_9080,N_6085,N_7694);
and U9081 (N_9081,N_6086,N_7369);
and U9082 (N_9082,N_6117,N_7828);
nand U9083 (N_9083,N_7871,N_6375);
or U9084 (N_9084,N_6009,N_6988);
nor U9085 (N_9085,N_6308,N_6657);
and U9086 (N_9086,N_7930,N_7521);
nand U9087 (N_9087,N_6439,N_6578);
or U9088 (N_9088,N_7321,N_6044);
and U9089 (N_9089,N_7680,N_6993);
nor U9090 (N_9090,N_6502,N_6919);
nand U9091 (N_9091,N_7910,N_7918);
xnor U9092 (N_9092,N_6320,N_7971);
or U9093 (N_9093,N_7581,N_6709);
or U9094 (N_9094,N_7743,N_6995);
and U9095 (N_9095,N_7542,N_6098);
xor U9096 (N_9096,N_7775,N_6209);
xor U9097 (N_9097,N_7297,N_6878);
or U9098 (N_9098,N_6944,N_7579);
or U9099 (N_9099,N_6809,N_6750);
nand U9100 (N_9100,N_7245,N_7879);
nor U9101 (N_9101,N_7409,N_6395);
and U9102 (N_9102,N_6658,N_7844);
xor U9103 (N_9103,N_7791,N_6405);
nand U9104 (N_9104,N_7587,N_6490);
and U9105 (N_9105,N_7859,N_6812);
and U9106 (N_9106,N_6393,N_6050);
or U9107 (N_9107,N_7562,N_6551);
nor U9108 (N_9108,N_7949,N_6574);
nand U9109 (N_9109,N_6771,N_6430);
nand U9110 (N_9110,N_6276,N_7015);
xor U9111 (N_9111,N_7364,N_7667);
xor U9112 (N_9112,N_7856,N_7869);
nor U9113 (N_9113,N_6472,N_7047);
or U9114 (N_9114,N_7704,N_7513);
or U9115 (N_9115,N_6842,N_6883);
nand U9116 (N_9116,N_6761,N_7229);
nand U9117 (N_9117,N_7430,N_7353);
or U9118 (N_9118,N_7009,N_6084);
nor U9119 (N_9119,N_7329,N_7656);
xnor U9120 (N_9120,N_6156,N_7948);
and U9121 (N_9121,N_7932,N_6156);
nor U9122 (N_9122,N_6485,N_7634);
and U9123 (N_9123,N_7073,N_6286);
nor U9124 (N_9124,N_7842,N_6742);
nand U9125 (N_9125,N_6750,N_7994);
and U9126 (N_9126,N_7063,N_7029);
nor U9127 (N_9127,N_7129,N_7778);
nor U9128 (N_9128,N_6438,N_6944);
nor U9129 (N_9129,N_7069,N_6761);
xor U9130 (N_9130,N_7178,N_7284);
or U9131 (N_9131,N_7837,N_7515);
nor U9132 (N_9132,N_7052,N_6349);
xor U9133 (N_9133,N_6610,N_7440);
nand U9134 (N_9134,N_6262,N_6110);
and U9135 (N_9135,N_6150,N_7492);
xor U9136 (N_9136,N_7956,N_7677);
and U9137 (N_9137,N_7899,N_6806);
xnor U9138 (N_9138,N_6367,N_6190);
nor U9139 (N_9139,N_6415,N_7918);
xnor U9140 (N_9140,N_6941,N_7972);
xor U9141 (N_9141,N_7815,N_6702);
xnor U9142 (N_9142,N_6847,N_6667);
and U9143 (N_9143,N_7775,N_6684);
nor U9144 (N_9144,N_7773,N_6633);
nor U9145 (N_9145,N_6969,N_6125);
or U9146 (N_9146,N_7945,N_6080);
or U9147 (N_9147,N_7374,N_7280);
and U9148 (N_9148,N_6972,N_6495);
nor U9149 (N_9149,N_6145,N_6561);
xor U9150 (N_9150,N_7643,N_7907);
and U9151 (N_9151,N_7469,N_7636);
or U9152 (N_9152,N_6784,N_6194);
xnor U9153 (N_9153,N_7352,N_7325);
nand U9154 (N_9154,N_7204,N_7754);
xor U9155 (N_9155,N_6483,N_7439);
nor U9156 (N_9156,N_7951,N_6421);
xor U9157 (N_9157,N_7300,N_6548);
nor U9158 (N_9158,N_7049,N_6237);
nand U9159 (N_9159,N_6769,N_7766);
nor U9160 (N_9160,N_7302,N_7515);
xnor U9161 (N_9161,N_7851,N_6011);
xor U9162 (N_9162,N_6867,N_7743);
nor U9163 (N_9163,N_6615,N_7066);
xor U9164 (N_9164,N_6693,N_6730);
or U9165 (N_9165,N_6544,N_7783);
nand U9166 (N_9166,N_7794,N_7834);
nand U9167 (N_9167,N_7230,N_6633);
nor U9168 (N_9168,N_6991,N_6433);
nor U9169 (N_9169,N_6987,N_7051);
xnor U9170 (N_9170,N_7893,N_6288);
and U9171 (N_9171,N_6824,N_7219);
and U9172 (N_9172,N_6849,N_6368);
or U9173 (N_9173,N_7693,N_6000);
and U9174 (N_9174,N_6117,N_6612);
nand U9175 (N_9175,N_7054,N_7708);
or U9176 (N_9176,N_7245,N_6969);
nand U9177 (N_9177,N_7751,N_7218);
nand U9178 (N_9178,N_6850,N_6687);
nand U9179 (N_9179,N_6777,N_6368);
nand U9180 (N_9180,N_6339,N_7433);
xnor U9181 (N_9181,N_7974,N_6320);
xor U9182 (N_9182,N_7429,N_7033);
or U9183 (N_9183,N_7845,N_6739);
xor U9184 (N_9184,N_6987,N_6306);
or U9185 (N_9185,N_7127,N_7550);
nor U9186 (N_9186,N_7917,N_7958);
xor U9187 (N_9187,N_7483,N_6530);
nor U9188 (N_9188,N_6442,N_7950);
nor U9189 (N_9189,N_6221,N_7378);
xnor U9190 (N_9190,N_7872,N_7860);
or U9191 (N_9191,N_6467,N_6011);
nor U9192 (N_9192,N_6865,N_7521);
or U9193 (N_9193,N_6463,N_6468);
or U9194 (N_9194,N_7361,N_7119);
nand U9195 (N_9195,N_6825,N_6071);
or U9196 (N_9196,N_7504,N_7724);
nand U9197 (N_9197,N_6708,N_6446);
nor U9198 (N_9198,N_6499,N_7450);
and U9199 (N_9199,N_7314,N_7823);
nand U9200 (N_9200,N_7310,N_6399);
and U9201 (N_9201,N_6045,N_6359);
nor U9202 (N_9202,N_6364,N_6014);
nand U9203 (N_9203,N_6272,N_7825);
and U9204 (N_9204,N_7807,N_6907);
or U9205 (N_9205,N_6023,N_6789);
xor U9206 (N_9206,N_7726,N_6950);
or U9207 (N_9207,N_7912,N_6778);
xor U9208 (N_9208,N_7678,N_6963);
or U9209 (N_9209,N_6175,N_7517);
nand U9210 (N_9210,N_6879,N_6877);
and U9211 (N_9211,N_7707,N_6709);
nand U9212 (N_9212,N_6094,N_7299);
and U9213 (N_9213,N_7836,N_7673);
or U9214 (N_9214,N_6575,N_6735);
nand U9215 (N_9215,N_6893,N_7661);
nand U9216 (N_9216,N_6904,N_7395);
and U9217 (N_9217,N_7896,N_7902);
or U9218 (N_9218,N_7441,N_6037);
nand U9219 (N_9219,N_7263,N_6741);
nor U9220 (N_9220,N_7648,N_7808);
xor U9221 (N_9221,N_7880,N_7452);
nor U9222 (N_9222,N_6689,N_7207);
and U9223 (N_9223,N_7397,N_7805);
nand U9224 (N_9224,N_7036,N_7567);
nor U9225 (N_9225,N_7602,N_6995);
nand U9226 (N_9226,N_7760,N_6937);
and U9227 (N_9227,N_7384,N_7642);
xnor U9228 (N_9228,N_6622,N_6588);
nand U9229 (N_9229,N_7779,N_7249);
or U9230 (N_9230,N_7685,N_7610);
and U9231 (N_9231,N_7690,N_7492);
or U9232 (N_9232,N_7180,N_6479);
and U9233 (N_9233,N_6543,N_6626);
xnor U9234 (N_9234,N_7834,N_7731);
and U9235 (N_9235,N_6451,N_7599);
xor U9236 (N_9236,N_7473,N_6365);
nor U9237 (N_9237,N_7663,N_7473);
nand U9238 (N_9238,N_7913,N_7870);
nand U9239 (N_9239,N_7996,N_6178);
and U9240 (N_9240,N_6436,N_7217);
nand U9241 (N_9241,N_7993,N_6821);
and U9242 (N_9242,N_6261,N_6442);
nand U9243 (N_9243,N_7827,N_7844);
and U9244 (N_9244,N_6955,N_6752);
or U9245 (N_9245,N_6485,N_6938);
nand U9246 (N_9246,N_6738,N_6933);
or U9247 (N_9247,N_7301,N_7902);
and U9248 (N_9248,N_6797,N_7011);
nor U9249 (N_9249,N_6486,N_7743);
or U9250 (N_9250,N_7945,N_6506);
xor U9251 (N_9251,N_6669,N_6152);
xor U9252 (N_9252,N_7200,N_7641);
xor U9253 (N_9253,N_6905,N_7385);
nor U9254 (N_9254,N_6874,N_7730);
and U9255 (N_9255,N_6599,N_6780);
or U9256 (N_9256,N_6853,N_6092);
nand U9257 (N_9257,N_7950,N_6148);
nand U9258 (N_9258,N_6637,N_6014);
nand U9259 (N_9259,N_7403,N_7702);
or U9260 (N_9260,N_6986,N_6957);
nand U9261 (N_9261,N_7797,N_7435);
or U9262 (N_9262,N_7235,N_7886);
nor U9263 (N_9263,N_6844,N_6434);
nand U9264 (N_9264,N_7911,N_7174);
nor U9265 (N_9265,N_6324,N_6066);
and U9266 (N_9266,N_6011,N_6756);
nand U9267 (N_9267,N_6605,N_7440);
xnor U9268 (N_9268,N_7740,N_6431);
nor U9269 (N_9269,N_7553,N_6799);
and U9270 (N_9270,N_6368,N_7001);
nand U9271 (N_9271,N_7041,N_7778);
xnor U9272 (N_9272,N_7494,N_7072);
xnor U9273 (N_9273,N_7414,N_6022);
or U9274 (N_9274,N_6539,N_7745);
xor U9275 (N_9275,N_6741,N_7264);
and U9276 (N_9276,N_6802,N_7667);
and U9277 (N_9277,N_7942,N_6370);
nand U9278 (N_9278,N_6318,N_7859);
nor U9279 (N_9279,N_7914,N_7523);
or U9280 (N_9280,N_6261,N_7940);
nor U9281 (N_9281,N_7715,N_6886);
xnor U9282 (N_9282,N_7026,N_6088);
nor U9283 (N_9283,N_6534,N_7631);
or U9284 (N_9284,N_7034,N_7551);
and U9285 (N_9285,N_6357,N_7670);
nand U9286 (N_9286,N_6856,N_7652);
nand U9287 (N_9287,N_7734,N_6505);
and U9288 (N_9288,N_6743,N_6496);
and U9289 (N_9289,N_6731,N_6010);
or U9290 (N_9290,N_7709,N_7552);
or U9291 (N_9291,N_7588,N_7764);
nor U9292 (N_9292,N_7718,N_6490);
and U9293 (N_9293,N_6832,N_6048);
nor U9294 (N_9294,N_7471,N_6431);
xnor U9295 (N_9295,N_7842,N_6489);
or U9296 (N_9296,N_7893,N_7567);
and U9297 (N_9297,N_6779,N_6924);
and U9298 (N_9298,N_6118,N_7586);
nand U9299 (N_9299,N_7927,N_7979);
nand U9300 (N_9300,N_7888,N_6444);
and U9301 (N_9301,N_6419,N_7264);
and U9302 (N_9302,N_6246,N_6763);
nand U9303 (N_9303,N_6440,N_7056);
nand U9304 (N_9304,N_7660,N_6688);
or U9305 (N_9305,N_7306,N_7163);
and U9306 (N_9306,N_6235,N_7979);
nor U9307 (N_9307,N_7624,N_7957);
nor U9308 (N_9308,N_7948,N_6098);
nand U9309 (N_9309,N_7300,N_6908);
nand U9310 (N_9310,N_6241,N_7152);
or U9311 (N_9311,N_6402,N_6572);
and U9312 (N_9312,N_7996,N_7976);
and U9313 (N_9313,N_6083,N_6443);
nor U9314 (N_9314,N_6910,N_7802);
nand U9315 (N_9315,N_7510,N_6837);
and U9316 (N_9316,N_7775,N_7988);
xor U9317 (N_9317,N_7758,N_6998);
nand U9318 (N_9318,N_7376,N_6030);
xor U9319 (N_9319,N_6827,N_7029);
or U9320 (N_9320,N_7712,N_7664);
xnor U9321 (N_9321,N_6746,N_6158);
nor U9322 (N_9322,N_7757,N_6722);
and U9323 (N_9323,N_6039,N_6411);
xnor U9324 (N_9324,N_7857,N_7125);
nand U9325 (N_9325,N_7958,N_7933);
or U9326 (N_9326,N_7033,N_6739);
or U9327 (N_9327,N_6525,N_7885);
and U9328 (N_9328,N_7746,N_7287);
nand U9329 (N_9329,N_7167,N_7606);
nor U9330 (N_9330,N_6028,N_6495);
nand U9331 (N_9331,N_7068,N_7655);
or U9332 (N_9332,N_7961,N_6000);
nor U9333 (N_9333,N_7202,N_6753);
nor U9334 (N_9334,N_6827,N_7685);
or U9335 (N_9335,N_6166,N_6886);
nor U9336 (N_9336,N_7458,N_6261);
xnor U9337 (N_9337,N_6519,N_6228);
and U9338 (N_9338,N_6613,N_6540);
nor U9339 (N_9339,N_6562,N_7208);
nand U9340 (N_9340,N_7967,N_7655);
xnor U9341 (N_9341,N_6315,N_6144);
nor U9342 (N_9342,N_6476,N_6962);
or U9343 (N_9343,N_6235,N_6313);
nand U9344 (N_9344,N_7751,N_6214);
nand U9345 (N_9345,N_7375,N_6490);
xnor U9346 (N_9346,N_6694,N_6625);
nor U9347 (N_9347,N_7028,N_6932);
nand U9348 (N_9348,N_6163,N_6187);
xnor U9349 (N_9349,N_7803,N_6290);
xnor U9350 (N_9350,N_6555,N_6694);
xor U9351 (N_9351,N_6994,N_6099);
nand U9352 (N_9352,N_7852,N_6056);
or U9353 (N_9353,N_6063,N_6206);
or U9354 (N_9354,N_6939,N_6106);
xnor U9355 (N_9355,N_7636,N_7053);
or U9356 (N_9356,N_7046,N_6483);
or U9357 (N_9357,N_7415,N_7600);
xor U9358 (N_9358,N_7404,N_6437);
xnor U9359 (N_9359,N_7797,N_6578);
nor U9360 (N_9360,N_6975,N_7689);
or U9361 (N_9361,N_6607,N_7765);
or U9362 (N_9362,N_7885,N_7974);
xnor U9363 (N_9363,N_7368,N_6486);
and U9364 (N_9364,N_6572,N_7653);
nor U9365 (N_9365,N_7476,N_6431);
or U9366 (N_9366,N_7704,N_6868);
nand U9367 (N_9367,N_6687,N_6652);
or U9368 (N_9368,N_6508,N_7170);
or U9369 (N_9369,N_7478,N_6628);
and U9370 (N_9370,N_7186,N_6909);
xnor U9371 (N_9371,N_6297,N_6837);
nor U9372 (N_9372,N_6236,N_7733);
xor U9373 (N_9373,N_6475,N_6432);
nor U9374 (N_9374,N_7353,N_7223);
nand U9375 (N_9375,N_7837,N_7616);
and U9376 (N_9376,N_6104,N_6272);
nand U9377 (N_9377,N_6196,N_6303);
xnor U9378 (N_9378,N_7883,N_7134);
nor U9379 (N_9379,N_7413,N_7615);
and U9380 (N_9380,N_6260,N_7651);
nand U9381 (N_9381,N_6921,N_6623);
and U9382 (N_9382,N_6018,N_7920);
nand U9383 (N_9383,N_6288,N_6197);
or U9384 (N_9384,N_7605,N_7726);
xnor U9385 (N_9385,N_7449,N_6451);
and U9386 (N_9386,N_6574,N_7613);
nand U9387 (N_9387,N_6815,N_6021);
nand U9388 (N_9388,N_6844,N_6153);
and U9389 (N_9389,N_6791,N_6388);
nand U9390 (N_9390,N_7704,N_6573);
nand U9391 (N_9391,N_6311,N_7112);
and U9392 (N_9392,N_6128,N_7910);
nand U9393 (N_9393,N_7413,N_6982);
xnor U9394 (N_9394,N_6195,N_6732);
nand U9395 (N_9395,N_7458,N_7515);
and U9396 (N_9396,N_7435,N_7927);
nor U9397 (N_9397,N_7139,N_6062);
and U9398 (N_9398,N_7014,N_6207);
and U9399 (N_9399,N_7504,N_6646);
nand U9400 (N_9400,N_7853,N_6107);
nor U9401 (N_9401,N_6454,N_7079);
xor U9402 (N_9402,N_7273,N_6543);
nand U9403 (N_9403,N_7793,N_7923);
xnor U9404 (N_9404,N_7990,N_6944);
and U9405 (N_9405,N_6090,N_7581);
or U9406 (N_9406,N_7684,N_6722);
and U9407 (N_9407,N_7379,N_6878);
and U9408 (N_9408,N_6025,N_7638);
nand U9409 (N_9409,N_7566,N_6093);
nand U9410 (N_9410,N_7446,N_7263);
nand U9411 (N_9411,N_7563,N_7365);
nand U9412 (N_9412,N_7221,N_7575);
or U9413 (N_9413,N_6587,N_6464);
nor U9414 (N_9414,N_7684,N_6153);
nand U9415 (N_9415,N_7656,N_7888);
nor U9416 (N_9416,N_6684,N_6916);
or U9417 (N_9417,N_7673,N_7419);
and U9418 (N_9418,N_7856,N_6135);
and U9419 (N_9419,N_7790,N_6902);
and U9420 (N_9420,N_7392,N_6238);
nand U9421 (N_9421,N_7177,N_6002);
or U9422 (N_9422,N_6055,N_7789);
nand U9423 (N_9423,N_6984,N_7019);
or U9424 (N_9424,N_6042,N_6940);
or U9425 (N_9425,N_7241,N_6192);
or U9426 (N_9426,N_6481,N_7278);
or U9427 (N_9427,N_6392,N_7631);
and U9428 (N_9428,N_7402,N_6922);
xnor U9429 (N_9429,N_7313,N_7226);
nor U9430 (N_9430,N_6332,N_6206);
xnor U9431 (N_9431,N_6320,N_7458);
or U9432 (N_9432,N_6353,N_6146);
nor U9433 (N_9433,N_7891,N_6346);
nor U9434 (N_9434,N_6674,N_7510);
and U9435 (N_9435,N_7852,N_7182);
and U9436 (N_9436,N_6314,N_6029);
and U9437 (N_9437,N_7482,N_7261);
nor U9438 (N_9438,N_6250,N_6174);
nand U9439 (N_9439,N_6015,N_7122);
nand U9440 (N_9440,N_7200,N_7664);
nor U9441 (N_9441,N_6036,N_7627);
xnor U9442 (N_9442,N_6997,N_7819);
or U9443 (N_9443,N_6535,N_7844);
or U9444 (N_9444,N_7327,N_6468);
or U9445 (N_9445,N_7223,N_7663);
xnor U9446 (N_9446,N_6855,N_7167);
nor U9447 (N_9447,N_6912,N_7917);
and U9448 (N_9448,N_6220,N_6674);
xnor U9449 (N_9449,N_7075,N_6533);
and U9450 (N_9450,N_6278,N_6911);
nand U9451 (N_9451,N_7271,N_7608);
xnor U9452 (N_9452,N_7605,N_6281);
and U9453 (N_9453,N_7717,N_6278);
nor U9454 (N_9454,N_6168,N_6908);
nor U9455 (N_9455,N_6312,N_7701);
nor U9456 (N_9456,N_7598,N_6175);
and U9457 (N_9457,N_6079,N_6483);
or U9458 (N_9458,N_6072,N_7431);
xnor U9459 (N_9459,N_6947,N_6784);
xor U9460 (N_9460,N_6246,N_7112);
and U9461 (N_9461,N_6506,N_7175);
and U9462 (N_9462,N_6862,N_7352);
xor U9463 (N_9463,N_6120,N_7469);
xor U9464 (N_9464,N_7593,N_7135);
and U9465 (N_9465,N_7308,N_6639);
or U9466 (N_9466,N_6759,N_7164);
nand U9467 (N_9467,N_6790,N_7399);
and U9468 (N_9468,N_6819,N_7808);
and U9469 (N_9469,N_7950,N_7106);
or U9470 (N_9470,N_7817,N_6249);
nor U9471 (N_9471,N_7015,N_6356);
xor U9472 (N_9472,N_7643,N_6003);
nor U9473 (N_9473,N_7244,N_6679);
and U9474 (N_9474,N_7850,N_6518);
or U9475 (N_9475,N_7590,N_7044);
nand U9476 (N_9476,N_6169,N_7982);
and U9477 (N_9477,N_6539,N_7172);
xor U9478 (N_9478,N_7856,N_6953);
and U9479 (N_9479,N_6761,N_7333);
or U9480 (N_9480,N_7846,N_6787);
nor U9481 (N_9481,N_7735,N_7055);
nand U9482 (N_9482,N_7624,N_7190);
and U9483 (N_9483,N_7952,N_7490);
and U9484 (N_9484,N_6602,N_6764);
or U9485 (N_9485,N_7898,N_6879);
nor U9486 (N_9486,N_6345,N_6928);
or U9487 (N_9487,N_7310,N_7513);
and U9488 (N_9488,N_6020,N_6758);
or U9489 (N_9489,N_7645,N_6963);
and U9490 (N_9490,N_6665,N_7606);
xor U9491 (N_9491,N_6488,N_6524);
and U9492 (N_9492,N_7295,N_6676);
or U9493 (N_9493,N_6664,N_7930);
nor U9494 (N_9494,N_7831,N_6116);
xnor U9495 (N_9495,N_6266,N_7459);
xnor U9496 (N_9496,N_7966,N_6759);
nor U9497 (N_9497,N_7792,N_7467);
or U9498 (N_9498,N_7823,N_6248);
and U9499 (N_9499,N_6508,N_7996);
xnor U9500 (N_9500,N_6944,N_7897);
xor U9501 (N_9501,N_6171,N_6704);
and U9502 (N_9502,N_7101,N_7566);
and U9503 (N_9503,N_7219,N_7581);
nor U9504 (N_9504,N_7205,N_7216);
nand U9505 (N_9505,N_7833,N_7908);
nor U9506 (N_9506,N_6732,N_7348);
nand U9507 (N_9507,N_6040,N_6261);
nand U9508 (N_9508,N_6399,N_7994);
xnor U9509 (N_9509,N_7102,N_6358);
xor U9510 (N_9510,N_7982,N_7224);
nand U9511 (N_9511,N_6345,N_6573);
nor U9512 (N_9512,N_6839,N_6047);
and U9513 (N_9513,N_7850,N_7151);
and U9514 (N_9514,N_6706,N_7707);
nor U9515 (N_9515,N_6311,N_6987);
and U9516 (N_9516,N_7125,N_6610);
xor U9517 (N_9517,N_7526,N_7849);
or U9518 (N_9518,N_6697,N_6159);
and U9519 (N_9519,N_7510,N_7027);
nand U9520 (N_9520,N_6586,N_6985);
xor U9521 (N_9521,N_6023,N_6719);
or U9522 (N_9522,N_6149,N_6571);
nor U9523 (N_9523,N_6921,N_6486);
xnor U9524 (N_9524,N_6413,N_6811);
nand U9525 (N_9525,N_6002,N_6086);
nand U9526 (N_9526,N_6252,N_6565);
xnor U9527 (N_9527,N_7854,N_6853);
nand U9528 (N_9528,N_7259,N_6929);
nand U9529 (N_9529,N_7169,N_6666);
xnor U9530 (N_9530,N_6757,N_6065);
and U9531 (N_9531,N_6361,N_7465);
nor U9532 (N_9532,N_7445,N_7794);
nor U9533 (N_9533,N_7204,N_7068);
and U9534 (N_9534,N_6006,N_7897);
nor U9535 (N_9535,N_7251,N_7845);
and U9536 (N_9536,N_7137,N_7344);
nor U9537 (N_9537,N_7380,N_7842);
nor U9538 (N_9538,N_6597,N_6333);
or U9539 (N_9539,N_7260,N_7280);
and U9540 (N_9540,N_6395,N_6677);
xor U9541 (N_9541,N_7827,N_6381);
nor U9542 (N_9542,N_6100,N_6652);
nor U9543 (N_9543,N_6449,N_7865);
xnor U9544 (N_9544,N_6147,N_6888);
nand U9545 (N_9545,N_7059,N_7921);
or U9546 (N_9546,N_7735,N_6955);
nand U9547 (N_9547,N_6310,N_6404);
nand U9548 (N_9548,N_6323,N_6640);
and U9549 (N_9549,N_6102,N_6886);
and U9550 (N_9550,N_6130,N_7735);
nor U9551 (N_9551,N_7087,N_7614);
and U9552 (N_9552,N_7064,N_7647);
nor U9553 (N_9553,N_6027,N_6260);
or U9554 (N_9554,N_6602,N_6269);
nand U9555 (N_9555,N_6761,N_6144);
and U9556 (N_9556,N_7997,N_6732);
xor U9557 (N_9557,N_7942,N_7243);
nand U9558 (N_9558,N_7811,N_7042);
and U9559 (N_9559,N_6577,N_6263);
xor U9560 (N_9560,N_6154,N_7624);
or U9561 (N_9561,N_6789,N_7535);
or U9562 (N_9562,N_7562,N_7240);
and U9563 (N_9563,N_6467,N_6709);
nor U9564 (N_9564,N_6512,N_7072);
nand U9565 (N_9565,N_7548,N_7262);
nor U9566 (N_9566,N_7222,N_7010);
and U9567 (N_9567,N_6328,N_7120);
xnor U9568 (N_9568,N_7392,N_7919);
nor U9569 (N_9569,N_6664,N_7057);
xnor U9570 (N_9570,N_7523,N_7408);
or U9571 (N_9571,N_6957,N_7130);
or U9572 (N_9572,N_6396,N_7073);
xnor U9573 (N_9573,N_7455,N_6500);
nand U9574 (N_9574,N_6661,N_7650);
and U9575 (N_9575,N_6992,N_6296);
or U9576 (N_9576,N_6965,N_6850);
nand U9577 (N_9577,N_6720,N_6078);
and U9578 (N_9578,N_6714,N_6271);
and U9579 (N_9579,N_6346,N_7018);
and U9580 (N_9580,N_7223,N_6835);
or U9581 (N_9581,N_6744,N_6550);
and U9582 (N_9582,N_6976,N_7970);
nand U9583 (N_9583,N_6813,N_7742);
nor U9584 (N_9584,N_7527,N_7914);
or U9585 (N_9585,N_6924,N_6032);
nor U9586 (N_9586,N_6739,N_7821);
and U9587 (N_9587,N_7894,N_7311);
xor U9588 (N_9588,N_7772,N_6888);
nand U9589 (N_9589,N_7713,N_6671);
nand U9590 (N_9590,N_6891,N_7602);
nand U9591 (N_9591,N_7083,N_7900);
and U9592 (N_9592,N_6687,N_6813);
or U9593 (N_9593,N_7537,N_7584);
nand U9594 (N_9594,N_7695,N_7480);
nor U9595 (N_9595,N_7864,N_6662);
or U9596 (N_9596,N_7243,N_7282);
or U9597 (N_9597,N_7577,N_7982);
and U9598 (N_9598,N_7985,N_6876);
xnor U9599 (N_9599,N_6706,N_7713);
xnor U9600 (N_9600,N_6429,N_6795);
xor U9601 (N_9601,N_6869,N_7014);
or U9602 (N_9602,N_6798,N_7658);
nor U9603 (N_9603,N_7016,N_6775);
nor U9604 (N_9604,N_7863,N_6883);
or U9605 (N_9605,N_7514,N_7819);
nor U9606 (N_9606,N_7895,N_7076);
or U9607 (N_9607,N_7238,N_6977);
nand U9608 (N_9608,N_6872,N_7503);
nand U9609 (N_9609,N_6655,N_7645);
nand U9610 (N_9610,N_6894,N_7905);
and U9611 (N_9611,N_6021,N_6508);
and U9612 (N_9612,N_7749,N_6570);
and U9613 (N_9613,N_6621,N_6393);
or U9614 (N_9614,N_6522,N_7112);
xor U9615 (N_9615,N_7439,N_7826);
nor U9616 (N_9616,N_6545,N_6891);
nor U9617 (N_9617,N_6354,N_6968);
or U9618 (N_9618,N_6850,N_7901);
nand U9619 (N_9619,N_6274,N_6556);
nand U9620 (N_9620,N_6077,N_7452);
xnor U9621 (N_9621,N_7705,N_7579);
nand U9622 (N_9622,N_7370,N_7063);
xnor U9623 (N_9623,N_7737,N_6635);
or U9624 (N_9624,N_7774,N_7112);
nand U9625 (N_9625,N_6970,N_7492);
or U9626 (N_9626,N_7210,N_7055);
nor U9627 (N_9627,N_7236,N_6477);
nand U9628 (N_9628,N_6145,N_6284);
nand U9629 (N_9629,N_6895,N_7708);
xor U9630 (N_9630,N_6873,N_6027);
and U9631 (N_9631,N_7885,N_6881);
or U9632 (N_9632,N_7525,N_7709);
or U9633 (N_9633,N_6586,N_7202);
and U9634 (N_9634,N_7053,N_7021);
nor U9635 (N_9635,N_6449,N_7993);
or U9636 (N_9636,N_6970,N_7648);
nor U9637 (N_9637,N_6640,N_6011);
xor U9638 (N_9638,N_7908,N_7326);
xor U9639 (N_9639,N_6514,N_6973);
and U9640 (N_9640,N_7722,N_7091);
or U9641 (N_9641,N_7494,N_6452);
nand U9642 (N_9642,N_6962,N_7813);
nand U9643 (N_9643,N_7382,N_7978);
or U9644 (N_9644,N_6671,N_7090);
nor U9645 (N_9645,N_6260,N_7859);
xnor U9646 (N_9646,N_7033,N_6110);
nor U9647 (N_9647,N_7661,N_7920);
or U9648 (N_9648,N_7069,N_6760);
nand U9649 (N_9649,N_6459,N_6728);
and U9650 (N_9650,N_7881,N_7940);
and U9651 (N_9651,N_7604,N_7996);
and U9652 (N_9652,N_6707,N_7460);
and U9653 (N_9653,N_7878,N_7772);
and U9654 (N_9654,N_6096,N_7309);
xor U9655 (N_9655,N_6382,N_7167);
or U9656 (N_9656,N_6181,N_7083);
or U9657 (N_9657,N_7788,N_6972);
nor U9658 (N_9658,N_7816,N_6801);
or U9659 (N_9659,N_7665,N_7444);
or U9660 (N_9660,N_7744,N_6114);
xor U9661 (N_9661,N_6662,N_6563);
nand U9662 (N_9662,N_7230,N_6559);
and U9663 (N_9663,N_6037,N_7868);
nand U9664 (N_9664,N_6949,N_6577);
nand U9665 (N_9665,N_7113,N_6078);
or U9666 (N_9666,N_7185,N_6629);
xnor U9667 (N_9667,N_7749,N_6402);
nand U9668 (N_9668,N_6706,N_7170);
xnor U9669 (N_9669,N_7777,N_6943);
xnor U9670 (N_9670,N_6024,N_7612);
xor U9671 (N_9671,N_7096,N_6424);
and U9672 (N_9672,N_6087,N_7282);
nand U9673 (N_9673,N_6583,N_6877);
nand U9674 (N_9674,N_7226,N_6577);
nand U9675 (N_9675,N_7012,N_7306);
or U9676 (N_9676,N_7083,N_7784);
or U9677 (N_9677,N_7373,N_6380);
and U9678 (N_9678,N_6116,N_7243);
nand U9679 (N_9679,N_7900,N_6533);
nand U9680 (N_9680,N_6569,N_7144);
xor U9681 (N_9681,N_7635,N_7868);
xnor U9682 (N_9682,N_6598,N_6527);
nand U9683 (N_9683,N_6973,N_7773);
nor U9684 (N_9684,N_6050,N_6052);
xor U9685 (N_9685,N_6027,N_6425);
nor U9686 (N_9686,N_6481,N_7416);
nor U9687 (N_9687,N_6813,N_7168);
and U9688 (N_9688,N_7972,N_7890);
nand U9689 (N_9689,N_6156,N_7712);
nand U9690 (N_9690,N_6140,N_6149);
and U9691 (N_9691,N_6620,N_6354);
or U9692 (N_9692,N_7025,N_6263);
nand U9693 (N_9693,N_7230,N_6741);
and U9694 (N_9694,N_6602,N_7658);
nand U9695 (N_9695,N_6200,N_7177);
or U9696 (N_9696,N_7300,N_6641);
or U9697 (N_9697,N_7909,N_6956);
nand U9698 (N_9698,N_6037,N_6751);
or U9699 (N_9699,N_6160,N_6352);
nor U9700 (N_9700,N_7590,N_7523);
xnor U9701 (N_9701,N_7945,N_7546);
and U9702 (N_9702,N_6285,N_6448);
nand U9703 (N_9703,N_6690,N_6900);
xor U9704 (N_9704,N_6743,N_7931);
xor U9705 (N_9705,N_7694,N_6491);
nand U9706 (N_9706,N_7706,N_6670);
nor U9707 (N_9707,N_6684,N_7046);
nand U9708 (N_9708,N_6073,N_6222);
and U9709 (N_9709,N_7997,N_7284);
and U9710 (N_9710,N_7674,N_6150);
nor U9711 (N_9711,N_7635,N_7713);
or U9712 (N_9712,N_7936,N_6549);
nor U9713 (N_9713,N_6610,N_6941);
nor U9714 (N_9714,N_6547,N_6486);
and U9715 (N_9715,N_6306,N_7089);
or U9716 (N_9716,N_6826,N_7288);
nand U9717 (N_9717,N_6626,N_6783);
and U9718 (N_9718,N_7080,N_6277);
and U9719 (N_9719,N_7776,N_7353);
nor U9720 (N_9720,N_6803,N_7006);
nor U9721 (N_9721,N_7338,N_7070);
nand U9722 (N_9722,N_7738,N_7764);
or U9723 (N_9723,N_7467,N_6116);
or U9724 (N_9724,N_6081,N_6297);
nor U9725 (N_9725,N_6934,N_7925);
nand U9726 (N_9726,N_6562,N_6883);
or U9727 (N_9727,N_7146,N_7159);
or U9728 (N_9728,N_6324,N_7232);
xnor U9729 (N_9729,N_7262,N_7842);
or U9730 (N_9730,N_7815,N_7273);
xor U9731 (N_9731,N_7819,N_6731);
xor U9732 (N_9732,N_7275,N_6945);
xor U9733 (N_9733,N_7881,N_6847);
or U9734 (N_9734,N_6179,N_6255);
xor U9735 (N_9735,N_6857,N_6344);
xnor U9736 (N_9736,N_6450,N_6283);
nand U9737 (N_9737,N_6294,N_7891);
or U9738 (N_9738,N_6586,N_7858);
xor U9739 (N_9739,N_7644,N_6860);
and U9740 (N_9740,N_6978,N_7120);
xnor U9741 (N_9741,N_6989,N_7131);
and U9742 (N_9742,N_7091,N_7375);
xor U9743 (N_9743,N_7828,N_7036);
and U9744 (N_9744,N_6703,N_6370);
and U9745 (N_9745,N_7080,N_7468);
and U9746 (N_9746,N_7324,N_6449);
nor U9747 (N_9747,N_6411,N_7399);
and U9748 (N_9748,N_7408,N_6010);
nor U9749 (N_9749,N_6268,N_6673);
xnor U9750 (N_9750,N_6102,N_7554);
nand U9751 (N_9751,N_6893,N_7913);
nand U9752 (N_9752,N_6710,N_6848);
nor U9753 (N_9753,N_7614,N_6989);
xnor U9754 (N_9754,N_7383,N_7555);
nor U9755 (N_9755,N_6891,N_6877);
or U9756 (N_9756,N_7182,N_7274);
nand U9757 (N_9757,N_7947,N_7754);
nand U9758 (N_9758,N_7662,N_6620);
or U9759 (N_9759,N_6447,N_6007);
or U9760 (N_9760,N_7874,N_7975);
and U9761 (N_9761,N_6588,N_7196);
nand U9762 (N_9762,N_7754,N_7771);
and U9763 (N_9763,N_6855,N_6432);
and U9764 (N_9764,N_6312,N_6310);
and U9765 (N_9765,N_7052,N_7756);
or U9766 (N_9766,N_7381,N_6058);
nand U9767 (N_9767,N_6546,N_7693);
nand U9768 (N_9768,N_7654,N_7061);
or U9769 (N_9769,N_7961,N_7970);
nand U9770 (N_9770,N_7187,N_6710);
and U9771 (N_9771,N_7632,N_7598);
nand U9772 (N_9772,N_6683,N_7093);
xnor U9773 (N_9773,N_7719,N_7375);
nor U9774 (N_9774,N_7513,N_7107);
nand U9775 (N_9775,N_7971,N_6797);
nor U9776 (N_9776,N_7865,N_7623);
nor U9777 (N_9777,N_7399,N_6987);
and U9778 (N_9778,N_6927,N_6425);
xor U9779 (N_9779,N_6303,N_7974);
and U9780 (N_9780,N_6790,N_7211);
nor U9781 (N_9781,N_6722,N_6757);
nor U9782 (N_9782,N_6171,N_6773);
xnor U9783 (N_9783,N_6757,N_7399);
nor U9784 (N_9784,N_6952,N_7818);
nor U9785 (N_9785,N_6933,N_6548);
or U9786 (N_9786,N_7555,N_6861);
and U9787 (N_9787,N_7702,N_7427);
and U9788 (N_9788,N_7293,N_6697);
nand U9789 (N_9789,N_7359,N_6930);
or U9790 (N_9790,N_7475,N_6561);
nor U9791 (N_9791,N_7101,N_6766);
xnor U9792 (N_9792,N_6242,N_7361);
or U9793 (N_9793,N_7813,N_7062);
or U9794 (N_9794,N_7008,N_6272);
nor U9795 (N_9795,N_6437,N_6784);
or U9796 (N_9796,N_7682,N_6503);
nor U9797 (N_9797,N_7227,N_6857);
nor U9798 (N_9798,N_7431,N_6728);
nor U9799 (N_9799,N_6330,N_7420);
nand U9800 (N_9800,N_7240,N_7741);
nor U9801 (N_9801,N_7558,N_7157);
and U9802 (N_9802,N_6181,N_6300);
xor U9803 (N_9803,N_6411,N_6439);
nand U9804 (N_9804,N_6426,N_6991);
or U9805 (N_9805,N_7152,N_6760);
and U9806 (N_9806,N_6696,N_6641);
nor U9807 (N_9807,N_6725,N_7558);
and U9808 (N_9808,N_7296,N_7869);
or U9809 (N_9809,N_7519,N_6844);
nor U9810 (N_9810,N_6528,N_7100);
and U9811 (N_9811,N_7022,N_6403);
or U9812 (N_9812,N_6831,N_7883);
xnor U9813 (N_9813,N_6500,N_6924);
nor U9814 (N_9814,N_6354,N_6548);
or U9815 (N_9815,N_7165,N_6096);
or U9816 (N_9816,N_7933,N_6480);
nand U9817 (N_9817,N_6207,N_7314);
and U9818 (N_9818,N_7369,N_6291);
or U9819 (N_9819,N_7595,N_6002);
and U9820 (N_9820,N_7374,N_6724);
nand U9821 (N_9821,N_6397,N_6916);
xnor U9822 (N_9822,N_6733,N_7893);
and U9823 (N_9823,N_7197,N_7682);
nand U9824 (N_9824,N_7852,N_7366);
and U9825 (N_9825,N_7106,N_7458);
nand U9826 (N_9826,N_6777,N_6196);
nand U9827 (N_9827,N_6656,N_6530);
xnor U9828 (N_9828,N_7144,N_7840);
and U9829 (N_9829,N_7539,N_7694);
or U9830 (N_9830,N_7630,N_6224);
or U9831 (N_9831,N_6054,N_6826);
nand U9832 (N_9832,N_7826,N_6553);
and U9833 (N_9833,N_6136,N_6920);
nand U9834 (N_9834,N_7445,N_7649);
or U9835 (N_9835,N_6747,N_7573);
xnor U9836 (N_9836,N_6653,N_6718);
xor U9837 (N_9837,N_7835,N_6192);
or U9838 (N_9838,N_6804,N_6381);
nand U9839 (N_9839,N_7039,N_6457);
xnor U9840 (N_9840,N_7277,N_7539);
or U9841 (N_9841,N_7059,N_7663);
or U9842 (N_9842,N_7429,N_7811);
xor U9843 (N_9843,N_7246,N_6437);
nor U9844 (N_9844,N_7014,N_6210);
xor U9845 (N_9845,N_6150,N_6588);
nor U9846 (N_9846,N_7644,N_7967);
or U9847 (N_9847,N_7448,N_6691);
and U9848 (N_9848,N_7707,N_6017);
and U9849 (N_9849,N_6299,N_7815);
or U9850 (N_9850,N_6411,N_7520);
nor U9851 (N_9851,N_7724,N_6403);
xor U9852 (N_9852,N_7752,N_7765);
or U9853 (N_9853,N_7654,N_7894);
and U9854 (N_9854,N_6262,N_7653);
and U9855 (N_9855,N_7305,N_6213);
and U9856 (N_9856,N_7024,N_7462);
or U9857 (N_9857,N_6988,N_7743);
nand U9858 (N_9858,N_6454,N_6939);
and U9859 (N_9859,N_7599,N_7160);
nor U9860 (N_9860,N_6520,N_6193);
nor U9861 (N_9861,N_7050,N_7296);
nor U9862 (N_9862,N_6356,N_7021);
nand U9863 (N_9863,N_7261,N_7417);
xor U9864 (N_9864,N_7731,N_6185);
or U9865 (N_9865,N_7788,N_7465);
nand U9866 (N_9866,N_7886,N_6342);
or U9867 (N_9867,N_6245,N_6503);
or U9868 (N_9868,N_6632,N_7925);
or U9869 (N_9869,N_7128,N_6627);
xor U9870 (N_9870,N_6142,N_6006);
nor U9871 (N_9871,N_7964,N_7379);
nor U9872 (N_9872,N_6848,N_7659);
and U9873 (N_9873,N_6573,N_6628);
xor U9874 (N_9874,N_7649,N_6771);
or U9875 (N_9875,N_7734,N_6357);
and U9876 (N_9876,N_6760,N_6014);
nand U9877 (N_9877,N_7384,N_6212);
nor U9878 (N_9878,N_7549,N_6484);
and U9879 (N_9879,N_6963,N_7794);
and U9880 (N_9880,N_7894,N_7677);
xor U9881 (N_9881,N_6503,N_6152);
nor U9882 (N_9882,N_6521,N_7160);
or U9883 (N_9883,N_7621,N_7962);
or U9884 (N_9884,N_7482,N_6650);
nand U9885 (N_9885,N_7717,N_7860);
nor U9886 (N_9886,N_6514,N_7793);
or U9887 (N_9887,N_7421,N_7288);
nand U9888 (N_9888,N_6035,N_7467);
or U9889 (N_9889,N_7474,N_7113);
nor U9890 (N_9890,N_6487,N_7735);
nor U9891 (N_9891,N_6761,N_7523);
nor U9892 (N_9892,N_7303,N_6886);
or U9893 (N_9893,N_6829,N_6084);
nand U9894 (N_9894,N_6458,N_7864);
and U9895 (N_9895,N_6851,N_7668);
nand U9896 (N_9896,N_7238,N_6604);
and U9897 (N_9897,N_6431,N_6158);
xnor U9898 (N_9898,N_6176,N_6587);
nor U9899 (N_9899,N_6297,N_7263);
xor U9900 (N_9900,N_7714,N_6387);
xnor U9901 (N_9901,N_6868,N_6290);
and U9902 (N_9902,N_6461,N_6714);
xnor U9903 (N_9903,N_7315,N_6440);
or U9904 (N_9904,N_6641,N_6811);
or U9905 (N_9905,N_6037,N_6624);
and U9906 (N_9906,N_6197,N_7786);
nor U9907 (N_9907,N_6287,N_6867);
nor U9908 (N_9908,N_6390,N_6391);
nand U9909 (N_9909,N_7634,N_6473);
or U9910 (N_9910,N_6539,N_6455);
and U9911 (N_9911,N_6517,N_6368);
nor U9912 (N_9912,N_7807,N_7310);
or U9913 (N_9913,N_7507,N_6473);
nand U9914 (N_9914,N_7358,N_6266);
nand U9915 (N_9915,N_7088,N_7613);
xnor U9916 (N_9916,N_6590,N_7175);
and U9917 (N_9917,N_7659,N_6004);
or U9918 (N_9918,N_7980,N_6293);
nor U9919 (N_9919,N_7969,N_7906);
and U9920 (N_9920,N_7758,N_7990);
nand U9921 (N_9921,N_7097,N_6313);
and U9922 (N_9922,N_6308,N_7035);
nand U9923 (N_9923,N_7417,N_6716);
xnor U9924 (N_9924,N_7125,N_6419);
xnor U9925 (N_9925,N_7879,N_7648);
nor U9926 (N_9926,N_6438,N_6984);
xnor U9927 (N_9927,N_6454,N_6914);
xor U9928 (N_9928,N_7928,N_7222);
xor U9929 (N_9929,N_7692,N_6579);
nor U9930 (N_9930,N_7120,N_7035);
xor U9931 (N_9931,N_7275,N_6275);
and U9932 (N_9932,N_7529,N_6548);
xnor U9933 (N_9933,N_6135,N_7973);
and U9934 (N_9934,N_6806,N_6922);
or U9935 (N_9935,N_7373,N_7317);
or U9936 (N_9936,N_6776,N_6664);
and U9937 (N_9937,N_6924,N_7573);
and U9938 (N_9938,N_7215,N_7392);
nand U9939 (N_9939,N_6664,N_7907);
xor U9940 (N_9940,N_7829,N_6466);
or U9941 (N_9941,N_7950,N_6706);
and U9942 (N_9942,N_7916,N_6777);
nand U9943 (N_9943,N_6307,N_7613);
nor U9944 (N_9944,N_7690,N_6980);
nand U9945 (N_9945,N_6932,N_7417);
nor U9946 (N_9946,N_7063,N_6535);
nor U9947 (N_9947,N_7216,N_6979);
nand U9948 (N_9948,N_7933,N_6331);
or U9949 (N_9949,N_6572,N_7625);
nor U9950 (N_9950,N_6666,N_7132);
nand U9951 (N_9951,N_6631,N_7350);
nand U9952 (N_9952,N_6373,N_7947);
xnor U9953 (N_9953,N_7074,N_7738);
nor U9954 (N_9954,N_7555,N_6470);
nor U9955 (N_9955,N_7353,N_6318);
and U9956 (N_9956,N_7987,N_7745);
and U9957 (N_9957,N_6167,N_6381);
xnor U9958 (N_9958,N_6543,N_6993);
or U9959 (N_9959,N_6819,N_7579);
and U9960 (N_9960,N_6670,N_7301);
and U9961 (N_9961,N_6499,N_7968);
nor U9962 (N_9962,N_7041,N_6122);
nor U9963 (N_9963,N_6567,N_7001);
and U9964 (N_9964,N_7688,N_7600);
nand U9965 (N_9965,N_6742,N_6342);
nor U9966 (N_9966,N_7349,N_6869);
nand U9967 (N_9967,N_7325,N_6175);
and U9968 (N_9968,N_7124,N_6042);
and U9969 (N_9969,N_6250,N_6058);
nand U9970 (N_9970,N_7959,N_7338);
nor U9971 (N_9971,N_7352,N_7626);
xnor U9972 (N_9972,N_6927,N_7816);
xnor U9973 (N_9973,N_6216,N_7446);
xor U9974 (N_9974,N_7496,N_6627);
nand U9975 (N_9975,N_6891,N_6799);
and U9976 (N_9976,N_6721,N_7462);
nand U9977 (N_9977,N_6888,N_6448);
and U9978 (N_9978,N_7529,N_7274);
xor U9979 (N_9979,N_7332,N_6148);
xnor U9980 (N_9980,N_7735,N_7691);
or U9981 (N_9981,N_7586,N_7119);
nand U9982 (N_9982,N_7807,N_7194);
and U9983 (N_9983,N_7464,N_7323);
xnor U9984 (N_9984,N_7673,N_6647);
nand U9985 (N_9985,N_7870,N_7201);
and U9986 (N_9986,N_7805,N_6813);
nand U9987 (N_9987,N_7961,N_6044);
nand U9988 (N_9988,N_7747,N_6712);
or U9989 (N_9989,N_6049,N_7116);
or U9990 (N_9990,N_7082,N_6348);
xor U9991 (N_9991,N_6078,N_6485);
and U9992 (N_9992,N_6910,N_6318);
or U9993 (N_9993,N_6093,N_6477);
nor U9994 (N_9994,N_6570,N_7607);
xor U9995 (N_9995,N_6258,N_6194);
nor U9996 (N_9996,N_6946,N_7857);
xnor U9997 (N_9997,N_6463,N_6471);
xor U9998 (N_9998,N_6452,N_6244);
and U9999 (N_9999,N_7811,N_7586);
nor U10000 (N_10000,N_9896,N_9010);
nor U10001 (N_10001,N_9854,N_8298);
xnor U10002 (N_10002,N_8573,N_8687);
nor U10003 (N_10003,N_9929,N_8086);
or U10004 (N_10004,N_9055,N_8362);
nor U10005 (N_10005,N_8945,N_9869);
xor U10006 (N_10006,N_8004,N_9718);
xnor U10007 (N_10007,N_8404,N_9085);
nand U10008 (N_10008,N_9362,N_8775);
and U10009 (N_10009,N_8593,N_8091);
and U10010 (N_10010,N_9924,N_9438);
and U10011 (N_10011,N_8802,N_9948);
xor U10012 (N_10012,N_8729,N_9781);
and U10013 (N_10013,N_8030,N_8027);
nand U10014 (N_10014,N_9427,N_9301);
nand U10015 (N_10015,N_9588,N_8385);
xor U10016 (N_10016,N_8604,N_8549);
and U10017 (N_10017,N_8466,N_9864);
and U10018 (N_10018,N_8267,N_9537);
and U10019 (N_10019,N_8672,N_8890);
nand U10020 (N_10020,N_8705,N_9753);
and U10021 (N_10021,N_9455,N_8182);
xnor U10022 (N_10022,N_8011,N_9098);
nor U10023 (N_10023,N_9934,N_8543);
nor U10024 (N_10024,N_8499,N_8081);
xor U10025 (N_10025,N_8761,N_9442);
or U10026 (N_10026,N_8072,N_9075);
xnor U10027 (N_10027,N_8542,N_9740);
and U10028 (N_10028,N_9120,N_8850);
or U10029 (N_10029,N_8896,N_9001);
and U10030 (N_10030,N_9474,N_8119);
and U10031 (N_10031,N_8155,N_9020);
nand U10032 (N_10032,N_8619,N_9198);
nand U10033 (N_10033,N_8796,N_9480);
and U10034 (N_10034,N_8765,N_9618);
and U10035 (N_10035,N_9830,N_9583);
xor U10036 (N_10036,N_8185,N_9628);
and U10037 (N_10037,N_9802,N_9617);
or U10038 (N_10038,N_9141,N_9481);
xor U10039 (N_10039,N_8352,N_9789);
nor U10040 (N_10040,N_9733,N_8618);
or U10041 (N_10041,N_8620,N_9265);
or U10042 (N_10042,N_9756,N_9182);
nor U10043 (N_10043,N_9408,N_9709);
or U10044 (N_10044,N_9521,N_8795);
xnor U10045 (N_10045,N_9766,N_9243);
and U10046 (N_10046,N_9181,N_9205);
or U10047 (N_10047,N_9834,N_9707);
or U10048 (N_10048,N_8962,N_8503);
or U10049 (N_10049,N_8410,N_8506);
xnor U10050 (N_10050,N_8422,N_9042);
and U10051 (N_10051,N_9108,N_9998);
or U10052 (N_10052,N_9147,N_9426);
nand U10053 (N_10053,N_9551,N_8184);
xor U10054 (N_10054,N_8942,N_8674);
nor U10055 (N_10055,N_8012,N_8288);
and U10056 (N_10056,N_8317,N_9953);
and U10057 (N_10057,N_9563,N_8412);
or U10058 (N_10058,N_8002,N_9876);
nor U10059 (N_10059,N_9549,N_8121);
nor U10060 (N_10060,N_9992,N_8148);
nor U10061 (N_10061,N_9890,N_9956);
and U10062 (N_10062,N_8658,N_8242);
or U10063 (N_10063,N_9463,N_8174);
xnor U10064 (N_10064,N_8591,N_9732);
and U10065 (N_10065,N_9107,N_8472);
and U10066 (N_10066,N_8290,N_9639);
and U10067 (N_10067,N_8846,N_8274);
xnor U10068 (N_10068,N_8331,N_9871);
xor U10069 (N_10069,N_9931,N_9633);
xnor U10070 (N_10070,N_9849,N_9882);
nand U10071 (N_10071,N_9449,N_9926);
nand U10072 (N_10072,N_8966,N_8793);
nand U10073 (N_10073,N_8143,N_9716);
xor U10074 (N_10074,N_8414,N_8068);
or U10075 (N_10075,N_9823,N_8758);
xor U10076 (N_10076,N_8611,N_8695);
and U10077 (N_10077,N_9545,N_8233);
nor U10078 (N_10078,N_9084,N_8101);
and U10079 (N_10079,N_8361,N_8296);
or U10080 (N_10080,N_9596,N_9105);
xnor U10081 (N_10081,N_8433,N_8189);
nor U10082 (N_10082,N_9217,N_8925);
nand U10083 (N_10083,N_8652,N_9996);
nand U10084 (N_10084,N_8548,N_8640);
and U10085 (N_10085,N_9782,N_9865);
and U10086 (N_10086,N_9062,N_9662);
or U10087 (N_10087,N_8228,N_8043);
or U10088 (N_10088,N_9570,N_8704);
and U10089 (N_10089,N_8938,N_9467);
nor U10090 (N_10090,N_8998,N_8161);
xnor U10091 (N_10091,N_9283,N_9257);
xnor U10092 (N_10092,N_8493,N_8328);
nand U10093 (N_10093,N_8500,N_8715);
xnor U10094 (N_10094,N_9347,N_9309);
xor U10095 (N_10095,N_9158,N_9542);
and U10096 (N_10096,N_9312,N_9398);
xnor U10097 (N_10097,N_8713,N_9341);
nor U10098 (N_10098,N_8368,N_9884);
nor U10099 (N_10099,N_9514,N_9820);
and U10100 (N_10100,N_9544,N_9389);
nand U10101 (N_10101,N_8755,N_8416);
or U10102 (N_10102,N_8044,N_8747);
nand U10103 (N_10103,N_8608,N_9152);
nor U10104 (N_10104,N_8558,N_8092);
or U10105 (N_10105,N_8862,N_9693);
xor U10106 (N_10106,N_8502,N_9028);
or U10107 (N_10107,N_9349,N_8532);
nand U10108 (N_10108,N_9614,N_9836);
nand U10109 (N_10109,N_8753,N_9813);
nor U10110 (N_10110,N_8899,N_9457);
or U10111 (N_10111,N_8306,N_9183);
and U10112 (N_10112,N_9985,N_9172);
nand U10113 (N_10113,N_8347,N_8431);
or U10114 (N_10114,N_8975,N_8964);
and U10115 (N_10115,N_9278,N_8486);
or U10116 (N_10116,N_9149,N_9047);
or U10117 (N_10117,N_8418,N_8078);
xnor U10118 (N_10118,N_8007,N_8401);
or U10119 (N_10119,N_8234,N_8988);
nor U10120 (N_10120,N_9798,N_9790);
nand U10121 (N_10121,N_8398,N_9477);
or U10122 (N_10122,N_8784,N_8151);
or U10123 (N_10123,N_9728,N_8733);
nand U10124 (N_10124,N_8671,N_8740);
or U10125 (N_10125,N_8047,N_9143);
xnor U10126 (N_10126,N_8179,N_8650);
nor U10127 (N_10127,N_8446,N_8224);
nor U10128 (N_10128,N_9529,N_9666);
nand U10129 (N_10129,N_9388,N_8302);
nor U10130 (N_10130,N_8874,N_8886);
and U10131 (N_10131,N_9987,N_9167);
nand U10132 (N_10132,N_9220,N_8336);
or U10133 (N_10133,N_8280,N_8842);
xor U10134 (N_10134,N_9346,N_8538);
xor U10135 (N_10135,N_8096,N_9195);
or U10136 (N_10136,N_9337,N_9280);
nand U10137 (N_10137,N_9074,N_8451);
or U10138 (N_10138,N_9725,N_8448);
nor U10139 (N_10139,N_9032,N_9510);
nand U10140 (N_10140,N_9527,N_9441);
and U10141 (N_10141,N_8763,N_9974);
or U10142 (N_10142,N_9784,N_9496);
nor U10143 (N_10143,N_8138,N_8498);
nand U10144 (N_10144,N_8567,N_9810);
and U10145 (N_10145,N_9684,N_8746);
xor U10146 (N_10146,N_9212,N_8948);
xor U10147 (N_10147,N_8635,N_8929);
and U10148 (N_10148,N_9952,N_9640);
nor U10149 (N_10149,N_8655,N_8140);
or U10150 (N_10150,N_8726,N_8191);
xor U10151 (N_10151,N_9921,N_8927);
nor U10152 (N_10152,N_9531,N_9980);
xor U10153 (N_10153,N_9720,N_8820);
and U10154 (N_10154,N_9623,N_8495);
nor U10155 (N_10155,N_9236,N_9609);
and U10156 (N_10156,N_8154,N_9373);
xnor U10157 (N_10157,N_9444,N_9904);
nor U10158 (N_10158,N_9995,N_8894);
or U10159 (N_10159,N_9885,N_8137);
and U10160 (N_10160,N_9254,N_9958);
nand U10161 (N_10161,N_8760,N_8623);
nor U10162 (N_10162,N_8196,N_9769);
nor U10163 (N_10163,N_8455,N_9848);
and U10164 (N_10164,N_9197,N_8617);
nand U10165 (N_10165,N_9306,N_8583);
xnor U10166 (N_10166,N_8314,N_9384);
nor U10167 (N_10167,N_8933,N_8207);
xnor U10168 (N_10168,N_8229,N_9487);
nor U10169 (N_10169,N_9997,N_9140);
nand U10170 (N_10170,N_9646,N_9196);
xor U10171 (N_10171,N_8491,N_9076);
and U10172 (N_10172,N_9380,N_8218);
xor U10173 (N_10173,N_9626,N_9523);
nor U10174 (N_10174,N_9379,N_9788);
and U10175 (N_10175,N_9376,N_9942);
or U10176 (N_10176,N_9004,N_8301);
and U10177 (N_10177,N_9819,N_9261);
and U10178 (N_10178,N_9967,N_9225);
xnor U10179 (N_10179,N_9550,N_9895);
xor U10180 (N_10180,N_9516,N_8434);
or U10181 (N_10181,N_9497,N_8510);
xor U10182 (N_10182,N_9951,N_9025);
nor U10183 (N_10183,N_9371,N_8065);
or U10184 (N_10184,N_8831,N_8147);
xnor U10185 (N_10185,N_9123,N_8197);
or U10186 (N_10186,N_8193,N_8996);
or U10187 (N_10187,N_8450,N_8585);
or U10188 (N_10188,N_9066,N_8642);
or U10189 (N_10189,N_8651,N_8947);
or U10190 (N_10190,N_8621,N_9354);
nand U10191 (N_10191,N_9378,N_9701);
nor U10192 (N_10192,N_8323,N_9223);
nor U10193 (N_10193,N_8406,N_8355);
xor U10194 (N_10194,N_9852,N_8615);
nor U10195 (N_10195,N_9695,N_9827);
xnor U10196 (N_10196,N_8093,N_8860);
or U10197 (N_10197,N_9824,N_9587);
and U10198 (N_10198,N_9641,N_9330);
and U10199 (N_10199,N_8958,N_9856);
xnor U10200 (N_10200,N_9901,N_8198);
nor U10201 (N_10201,N_9201,N_8142);
and U10202 (N_10202,N_8659,N_9174);
and U10203 (N_10203,N_9717,N_9161);
nor U10204 (N_10204,N_9858,N_8767);
nor U10205 (N_10205,N_8253,N_9874);
nor U10206 (N_10206,N_8054,N_9271);
nor U10207 (N_10207,N_8055,N_9667);
nor U10208 (N_10208,N_9375,N_8354);
or U10209 (N_10209,N_8042,N_9679);
and U10210 (N_10210,N_9590,N_9611);
xnor U10211 (N_10211,N_8985,N_9580);
nor U10212 (N_10212,N_8104,N_8235);
nor U10213 (N_10213,N_9336,N_8698);
and U10214 (N_10214,N_8654,N_9699);
xor U10215 (N_10215,N_8807,N_9381);
xnor U10216 (N_10216,N_8100,N_8186);
or U10217 (N_10217,N_8830,N_9139);
or U10218 (N_10218,N_8626,N_9232);
xor U10219 (N_10219,N_8968,N_9060);
xor U10220 (N_10220,N_8735,N_8483);
nor U10221 (N_10221,N_8381,N_9035);
nand U10222 (N_10222,N_9277,N_9739);
nor U10223 (N_10223,N_9959,N_8800);
nand U10224 (N_10224,N_8930,N_9897);
nand U10225 (N_10225,N_8809,N_9413);
nand U10226 (N_10226,N_8397,N_9994);
or U10227 (N_10227,N_9601,N_8478);
nor U10228 (N_10228,N_8969,N_9582);
and U10229 (N_10229,N_8117,N_9835);
nor U10230 (N_10230,N_8633,N_8613);
nor U10231 (N_10231,N_9267,N_8026);
nand U10232 (N_10232,N_8534,N_8308);
or U10233 (N_10233,N_9234,N_9476);
nand U10234 (N_10234,N_9268,N_9420);
nor U10235 (N_10235,N_8889,N_9907);
xnor U10236 (N_10236,N_8989,N_8006);
and U10237 (N_10237,N_9759,N_9841);
and U10238 (N_10238,N_9593,N_9465);
and U10239 (N_10239,N_8073,N_9272);
nand U10240 (N_10240,N_8520,N_9009);
xor U10241 (N_10241,N_9114,N_9129);
nand U10242 (N_10242,N_8089,N_9171);
xnor U10243 (N_10243,N_9654,N_9137);
xor U10244 (N_10244,N_8220,N_8700);
nor U10245 (N_10245,N_9644,N_9748);
nand U10246 (N_10246,N_8575,N_9540);
xnor U10247 (N_10247,N_9034,N_9318);
and U10248 (N_10248,N_8881,N_9089);
xnor U10249 (N_10249,N_9965,N_8772);
or U10250 (N_10250,N_9266,N_9344);
nor U10251 (N_10251,N_8984,N_9231);
or U10252 (N_10252,N_8821,N_8734);
nand U10253 (N_10253,N_9228,N_9579);
and U10254 (N_10254,N_9925,N_8826);
or U10255 (N_10255,N_9193,N_8957);
nor U10256 (N_10256,N_8946,N_8108);
and U10257 (N_10257,N_8653,N_8022);
nor U10258 (N_10258,N_8986,N_8497);
xor U10259 (N_10259,N_9533,N_9736);
xor U10260 (N_10260,N_9729,N_9303);
xor U10261 (N_10261,N_9064,N_9957);
and U10262 (N_10262,N_8808,N_9989);
nand U10263 (N_10263,N_9621,N_8438);
nand U10264 (N_10264,N_9585,N_8219);
nand U10265 (N_10265,N_9063,N_9316);
and U10266 (N_10266,N_8914,N_9770);
and U10267 (N_10267,N_8771,N_9829);
nand U10268 (N_10268,N_8514,N_8541);
and U10269 (N_10269,N_9675,N_9363);
xnor U10270 (N_10270,N_9356,N_9334);
xor U10271 (N_10271,N_9136,N_9061);
xor U10272 (N_10272,N_9397,N_8214);
xor U10273 (N_10273,N_8295,N_9902);
or U10274 (N_10274,N_8384,N_8134);
xnor U10275 (N_10275,N_9115,N_8291);
or U10276 (N_10276,N_8221,N_8344);
nand U10277 (N_10277,N_9661,N_9021);
and U10278 (N_10278,N_9660,N_8678);
or U10279 (N_10279,N_9711,N_8646);
or U10280 (N_10280,N_8085,N_8343);
xor U10281 (N_10281,N_8389,N_8243);
xnor U10282 (N_10282,N_8318,N_9875);
nor U10283 (N_10283,N_9048,N_8609);
nand U10284 (N_10284,N_9599,N_9778);
or U10285 (N_10285,N_9470,N_8892);
and U10286 (N_10286,N_8175,N_9504);
xor U10287 (N_10287,N_9619,N_8827);
xnor U10288 (N_10288,N_9905,N_9226);
or U10289 (N_10289,N_8013,N_9402);
nor U10290 (N_10290,N_8424,N_9863);
or U10291 (N_10291,N_9304,N_9148);
or U10292 (N_10292,N_9180,N_8511);
nand U10293 (N_10293,N_9743,N_9710);
nand U10294 (N_10294,N_9012,N_9393);
nor U10295 (N_10295,N_8828,N_9469);
or U10296 (N_10296,N_9530,N_8790);
xor U10297 (N_10297,N_9305,N_8870);
nor U10298 (N_10298,N_8634,N_9811);
xor U10299 (N_10299,N_9322,N_9664);
or U10300 (N_10300,N_9809,N_9534);
nor U10301 (N_10301,N_8132,N_8074);
nand U10302 (N_10302,N_8387,N_9451);
or U10303 (N_10303,N_8866,N_8492);
nor U10304 (N_10304,N_9401,N_9296);
and U10305 (N_10305,N_9093,N_9622);
nor U10306 (N_10306,N_8061,N_8029);
xnor U10307 (N_10307,N_8904,N_9883);
and U10308 (N_10308,N_9574,N_8107);
nand U10309 (N_10309,N_9763,N_8550);
nand U10310 (N_10310,N_8601,N_8912);
and U10311 (N_10311,N_9691,N_8690);
nor U10312 (N_10312,N_9165,N_9100);
xnor U10313 (N_10313,N_8409,N_9216);
or U10314 (N_10314,N_9391,N_8120);
or U10315 (N_10315,N_9635,N_8786);
nor U10316 (N_10316,N_9466,N_8701);
xnor U10317 (N_10317,N_9026,N_9104);
or U10318 (N_10318,N_8403,N_8041);
xnor U10319 (N_10319,N_9122,N_9124);
nand U10320 (N_10320,N_9353,N_8832);
and U10321 (N_10321,N_8162,N_8415);
or U10322 (N_10322,N_9742,N_8390);
nor U10323 (N_10323,N_9630,N_8526);
and U10324 (N_10324,N_8366,N_8359);
and U10325 (N_10325,N_9478,N_8803);
xnor U10326 (N_10326,N_8512,N_9366);
xor U10327 (N_10327,N_8707,N_8867);
xor U10328 (N_10328,N_9979,N_8702);
and U10329 (N_10329,N_8363,N_9650);
or U10330 (N_10330,N_9258,N_8452);
nand U10331 (N_10331,N_9482,N_9433);
xor U10332 (N_10332,N_8321,N_8970);
or U10333 (N_10333,N_8113,N_9252);
nor U10334 (N_10334,N_8139,N_9773);
xnor U10335 (N_10335,N_8494,N_8563);
xor U10336 (N_10336,N_8126,N_9735);
or U10337 (N_10337,N_8895,N_8313);
and U10338 (N_10338,N_9595,N_8241);
nor U10339 (N_10339,N_8232,N_8835);
or U10340 (N_10340,N_9826,N_9439);
nand U10341 (N_10341,N_8782,N_9051);
xor U10342 (N_10342,N_9991,N_8001);
nor U10343 (N_10343,N_8873,N_8961);
xnor U10344 (N_10344,N_9150,N_8552);
xnor U10345 (N_10345,N_9390,N_9135);
or U10346 (N_10346,N_8884,N_9270);
and U10347 (N_10347,N_9333,N_8710);
nand U10348 (N_10348,N_8776,N_8923);
nor U10349 (N_10349,N_8407,N_9737);
or U10350 (N_10350,N_9815,N_9919);
nand U10351 (N_10351,N_9357,N_9799);
nor U10352 (N_10352,N_8838,N_9249);
or U10353 (N_10353,N_9112,N_8067);
and U10354 (N_10354,N_9768,N_9604);
and U10355 (N_10355,N_9538,N_9638);
or U10356 (N_10356,N_8736,N_8666);
nand U10357 (N_10357,N_8906,N_9414);
or U10358 (N_10358,N_9543,N_8168);
or U10359 (N_10359,N_9524,N_8281);
xor U10360 (N_10360,N_8667,N_9065);
nand U10361 (N_10361,N_8977,N_9264);
and U10362 (N_10362,N_9282,N_8237);
nand U10363 (N_10363,N_8665,N_9396);
xnor U10364 (N_10364,N_8245,N_8156);
nand U10365 (N_10365,N_8587,N_8683);
nor U10366 (N_10366,N_8825,N_9208);
or U10367 (N_10367,N_8584,N_8792);
xor U10368 (N_10368,N_8829,N_8423);
xor U10369 (N_10369,N_9289,N_9800);
nor U10370 (N_10370,N_8400,N_9307);
nand U10371 (N_10371,N_8568,N_9687);
nand U10372 (N_10372,N_8950,N_9801);
and U10373 (N_10373,N_9950,N_8959);
xnor U10374 (N_10374,N_9636,N_8066);
nand U10375 (N_10375,N_9475,N_8031);
nor U10376 (N_10376,N_9456,N_8656);
nor U10377 (N_10377,N_8059,N_8339);
nand U10378 (N_10378,N_8489,N_8124);
and U10379 (N_10379,N_9116,N_8668);
and U10380 (N_10380,N_9555,N_8730);
nand U10381 (N_10381,N_8071,N_9059);
and U10382 (N_10382,N_9041,N_9765);
or U10383 (N_10383,N_8170,N_8684);
nand U10384 (N_10384,N_8246,N_8614);
and U10385 (N_10385,N_8277,N_9647);
nor U10386 (N_10386,N_9435,N_9715);
nand U10387 (N_10387,N_9440,N_8266);
and U10388 (N_10388,N_9859,N_9088);
nand U10389 (N_10389,N_8859,N_9620);
nor U10390 (N_10390,N_8610,N_9941);
nor U10391 (N_10391,N_9973,N_8202);
xnor U10392 (N_10392,N_8356,N_8588);
nor U10393 (N_10393,N_9525,N_9081);
and U10394 (N_10394,N_9315,N_8643);
or U10395 (N_10395,N_9052,N_8109);
xnor U10396 (N_10396,N_9351,N_8582);
nor U10397 (N_10397,N_8284,N_9955);
or U10398 (N_10398,N_9079,N_9177);
nand U10399 (N_10399,N_8783,N_8180);
or U10400 (N_10400,N_8675,N_8084);
and U10401 (N_10401,N_9526,N_9787);
and U10402 (N_10402,N_8806,N_9567);
xnor U10403 (N_10403,N_8262,N_8839);
nor U10404 (N_10404,N_8509,N_8199);
nor U10405 (N_10405,N_9923,N_9259);
and U10406 (N_10406,N_9888,N_9310);
nor U10407 (N_10407,N_8903,N_8380);
nor U10408 (N_10408,N_8905,N_9731);
nand U10409 (N_10409,N_8854,N_9886);
and U10410 (N_10410,N_9983,N_8299);
nand U10411 (N_10411,N_9853,N_9803);
and U10412 (N_10412,N_8333,N_8158);
or U10413 (N_10413,N_9215,N_9324);
nand U10414 (N_10414,N_8539,N_8015);
nand U10415 (N_10415,N_8943,N_8141);
or U10416 (N_10416,N_9460,N_8670);
xnor U10417 (N_10417,N_9067,N_9068);
xor U10418 (N_10418,N_8562,N_8097);
xor U10419 (N_10419,N_9860,N_8038);
or U10420 (N_10420,N_9719,N_8394);
nand U10421 (N_10421,N_9038,N_8797);
nor U10422 (N_10422,N_9007,N_8627);
and U10423 (N_10423,N_9539,N_9916);
or U10424 (N_10424,N_9155,N_9263);
nand U10425 (N_10425,N_9328,N_8016);
xor U10426 (N_10426,N_9429,N_9502);
xnor U10427 (N_10427,N_8953,N_8122);
and U10428 (N_10428,N_9677,N_8293);
nor U10429 (N_10429,N_9615,N_9222);
xor U10430 (N_10430,N_9818,N_8467);
and U10431 (N_10431,N_9253,N_8883);
nor U10432 (N_10432,N_9764,N_8470);
xor U10433 (N_10433,N_9031,N_9127);
nand U10434 (N_10434,N_9045,N_8928);
xor U10435 (N_10435,N_9757,N_9900);
nor U10436 (N_10436,N_9168,N_8559);
nand U10437 (N_10437,N_8282,N_8723);
xor U10438 (N_10438,N_8738,N_9332);
xnor U10439 (N_10439,N_9117,N_8863);
or U10440 (N_10440,N_8367,N_9977);
or U10441 (N_10441,N_9912,N_8206);
xor U10442 (N_10442,N_9369,N_9988);
and U10443 (N_10443,N_8128,N_8993);
or U10444 (N_10444,N_9483,N_8980);
nor U10445 (N_10445,N_8247,N_8442);
nor U10446 (N_10446,N_8999,N_8307);
nor U10447 (N_10447,N_8173,N_9937);
xor U10448 (N_10448,N_9505,N_8851);
nand U10449 (N_10449,N_9187,N_8264);
xor U10450 (N_10450,N_9632,N_8459);
or U10451 (N_10451,N_8521,N_8664);
nand U10452 (N_10452,N_9339,N_9491);
and U10453 (N_10453,N_9598,N_9683);
and U10454 (N_10454,N_9688,N_8660);
nor U10455 (N_10455,N_8836,N_9434);
nor U10456 (N_10456,N_8069,N_9454);
or U10457 (N_10457,N_9606,N_8531);
nand U10458 (N_10458,N_8337,N_8032);
nor U10459 (N_10459,N_9960,N_8437);
and U10460 (N_10460,N_9793,N_8145);
nand U10461 (N_10461,N_8960,N_8703);
and U10462 (N_10462,N_9040,N_8425);
or U10463 (N_10463,N_9892,N_9610);
and U10464 (N_10464,N_9692,N_9109);
nor U10465 (N_10465,N_9473,N_9602);
nor U10466 (N_10466,N_9246,N_9706);
nor U10467 (N_10467,N_8922,N_8597);
nand U10468 (N_10468,N_9338,N_8223);
or U10469 (N_10469,N_9943,N_9909);
nand U10470 (N_10470,N_9893,N_9290);
xor U10471 (N_10471,N_9839,N_9548);
xor U10472 (N_10472,N_9984,N_9930);
nand U10473 (N_10473,N_9325,N_8956);
xor U10474 (N_10474,N_8877,N_9377);
nand U10475 (N_10475,N_9961,N_8458);
or U10476 (N_10476,N_8350,N_8129);
nand U10477 (N_10477,N_9682,N_8050);
nand U10478 (N_10478,N_8560,N_9520);
or U10479 (N_10479,N_8523,N_8464);
nor U10480 (N_10480,N_9121,N_9592);
or U10481 (N_10481,N_9918,N_9308);
or U10482 (N_10482,N_8209,N_9698);
nor U10483 (N_10483,N_9986,N_8334);
nand U10484 (N_10484,N_9843,N_8212);
and U10485 (N_10485,N_9690,N_9094);
nand U10486 (N_10486,N_8114,N_8987);
nor U10487 (N_10487,N_9877,N_9229);
nand U10488 (N_10488,N_9828,N_9284);
or U10489 (N_10489,N_8752,N_9237);
or U10490 (N_10490,N_9898,N_8739);
xor U10491 (N_10491,N_9411,N_9847);
nor U10492 (N_10492,N_9087,N_8990);
or U10493 (N_10493,N_9816,N_9342);
nor U10494 (N_10494,N_9297,N_9144);
or U10495 (N_10495,N_9071,N_8477);
nand U10496 (N_10496,N_8023,N_8110);
xor U10497 (N_10497,N_9131,N_8595);
nor U10498 (N_10498,N_8537,N_9436);
nor U10499 (N_10499,N_8324,N_9355);
xnor U10500 (N_10500,N_8577,N_9517);
and U10501 (N_10501,N_8332,N_9755);
nand U10502 (N_10502,N_9335,N_8978);
nand U10503 (N_10503,N_9151,N_9910);
nor U10504 (N_10504,N_8913,N_9671);
or U10505 (N_10505,N_9247,N_8471);
nand U10506 (N_10506,N_9488,N_8000);
and U10507 (N_10507,N_9947,N_9866);
and U10508 (N_10508,N_9037,N_8005);
or U10509 (N_10509,N_9724,N_9385);
xor U10510 (N_10510,N_8682,N_8391);
nor U10511 (N_10511,N_9792,N_9233);
and U10512 (N_10512,N_8364,N_9591);
nor U10513 (N_10513,N_8309,N_8811);
xnor U10514 (N_10514,N_8045,N_8845);
and U10515 (N_10515,N_8578,N_9288);
xor U10516 (N_10516,N_9565,N_9082);
and U10517 (N_10517,N_9039,N_9564);
nor U10518 (N_10518,N_9605,N_8529);
nor U10519 (N_10519,N_8728,N_9726);
and U10520 (N_10520,N_8625,N_9915);
or U10521 (N_10521,N_9668,N_9023);
xor U10522 (N_10522,N_8461,N_8791);
or U10523 (N_10523,N_9553,N_9777);
nor U10524 (N_10524,N_9224,N_8231);
and U10525 (N_10525,N_8430,N_9971);
xnor U10526 (N_10526,N_9556,N_8566);
nor U10527 (N_10527,N_8488,N_9722);
nand U10528 (N_10528,N_8751,N_9350);
and U10529 (N_10529,N_8112,N_8270);
or U10530 (N_10530,N_9513,N_9370);
xnor U10531 (N_10531,N_9500,N_9207);
xnor U10532 (N_10532,N_8051,N_8327);
and U10533 (N_10533,N_8505,N_9368);
nor U10534 (N_10534,N_9101,N_8632);
xor U10535 (N_10535,N_9821,N_9982);
and U10536 (N_10536,N_9273,N_9978);
nor U10537 (N_10537,N_9464,N_8516);
xor U10538 (N_10538,N_9184,N_9817);
xor U10539 (N_10539,N_8465,N_8688);
nand U10540 (N_10540,N_8580,N_8673);
nand U10541 (N_10541,N_8908,N_8369);
xor U10542 (N_10542,N_8581,N_9703);
nand U10543 (N_10543,N_9423,N_8160);
nor U10544 (N_10544,N_8133,N_9532);
xnor U10545 (N_10545,N_8440,N_9613);
nand U10546 (N_10546,N_8216,N_9281);
or U10547 (N_10547,N_9758,N_9577);
nor U10548 (N_10548,N_8794,N_8441);
or U10549 (N_10549,N_9881,N_8589);
or U10550 (N_10550,N_8320,N_9573);
nand U10551 (N_10551,N_8527,N_9558);
or U10552 (N_10552,N_9407,N_9714);
and U10553 (N_10553,N_8824,N_9750);
nand U10554 (N_10554,N_9844,N_8941);
xor U10555 (N_10555,N_8476,N_9586);
and U10556 (N_10556,N_8785,N_8463);
xor U10557 (N_10557,N_9576,N_9091);
xor U10558 (N_10558,N_9416,N_8427);
nand U10559 (N_10559,N_9199,N_8586);
or U10560 (N_10560,N_8818,N_9256);
or U10561 (N_10561,N_8856,N_9319);
xnor U10562 (N_10562,N_8094,N_9607);
or U10563 (N_10563,N_9134,N_9648);
xor U10564 (N_10564,N_9017,N_9867);
xnor U10565 (N_10565,N_8420,N_9169);
and U10566 (N_10566,N_8533,N_8303);
or U10567 (N_10567,N_8408,N_9846);
nand U10568 (N_10568,N_8484,N_8766);
nor U10569 (N_10569,N_8781,N_9498);
and U10570 (N_10570,N_9191,N_8816);
xnor U10571 (N_10571,N_9240,N_9862);
and U10572 (N_10572,N_9913,N_9230);
xor U10573 (N_10573,N_9645,N_9425);
or U10574 (N_10574,N_9033,N_9594);
or U10575 (N_10575,N_8706,N_9873);
or U10576 (N_10576,N_8965,N_8663);
or U10577 (N_10577,N_9200,N_8777);
and U10578 (N_10578,N_9430,N_8686);
nor U10579 (N_10579,N_8694,N_9751);
and U10580 (N_10580,N_9779,N_9581);
or U10581 (N_10581,N_8287,N_8770);
nor U10582 (N_10582,N_8208,N_8540);
xor U10583 (N_10583,N_9559,N_8024);
and U10584 (N_10584,N_8040,N_9861);
or U10585 (N_10585,N_8592,N_9145);
or U10586 (N_10586,N_9928,N_8457);
nand U10587 (N_10587,N_9894,N_8952);
nand U10588 (N_10588,N_8305,N_8572);
nor U10589 (N_10589,N_9340,N_8879);
nor U10590 (N_10590,N_9358,N_9651);
nor U10591 (N_10591,N_8149,N_9320);
nand U10592 (N_10592,N_8130,N_8021);
nand U10593 (N_10593,N_9406,N_8436);
nor U10594 (N_10594,N_9851,N_9327);
xor U10595 (N_10595,N_9727,N_9238);
or U10596 (N_10596,N_9070,N_8150);
xnor U10597 (N_10597,N_9431,N_9365);
xnor U10598 (N_10598,N_8865,N_8273);
nor U10599 (N_10599,N_9495,N_8915);
and U10600 (N_10600,N_9044,N_8555);
nand U10601 (N_10601,N_9274,N_8316);
or U10602 (N_10602,N_8157,N_8039);
or U10603 (N_10603,N_8501,N_9160);
or U10604 (N_10604,N_9612,N_8239);
nand U10605 (N_10605,N_8528,N_8429);
nand U10606 (N_10606,N_8916,N_9708);
nor U10607 (N_10607,N_8911,N_8371);
xnor U10608 (N_10608,N_8376,N_9383);
xor U10609 (N_10609,N_9786,N_8940);
or U10610 (N_10610,N_9410,N_9700);
or U10611 (N_10611,N_8153,N_9251);
or U10612 (N_10612,N_9119,N_9003);
or U10613 (N_10613,N_8750,N_9616);
xnor U10614 (N_10614,N_8090,N_9812);
or U10615 (N_10615,N_9569,N_8742);
nor U10616 (N_10616,N_9162,N_9014);
or U10617 (N_10617,N_8432,N_9775);
and U10618 (N_10618,N_9448,N_8982);
xnor U10619 (N_10619,N_8019,N_9872);
nand U10620 (N_10620,N_8530,N_9484);
or U10621 (N_10621,N_8382,N_9019);
nand U10622 (N_10622,N_8607,N_9073);
xor U10623 (N_10623,N_8645,N_9981);
nor U10624 (N_10624,N_8181,N_8857);
and U10625 (N_10625,N_9157,N_8649);
and U10626 (N_10626,N_8475,N_9054);
or U10627 (N_10627,N_8691,N_9494);
and U10628 (N_10628,N_8692,N_8056);
or U10629 (N_10629,N_8413,N_8574);
nand U10630 (N_10630,N_8435,N_9214);
xor U10631 (N_10631,N_9712,N_8256);
nor U10632 (N_10632,N_9964,N_9676);
or U10633 (N_10633,N_8377,N_9186);
and U10634 (N_10634,N_8631,N_8553);
and U10635 (N_10635,N_9221,N_9462);
nand U10636 (N_10636,N_8696,N_9395);
nor U10637 (N_10637,N_9642,N_9572);
xor U10638 (N_10638,N_9927,N_9702);
and U10639 (N_10639,N_8834,N_9512);
nor U10640 (N_10640,N_8762,N_9050);
or U10641 (N_10641,N_9036,N_9653);
nor U10642 (N_10642,N_9880,N_8351);
xor U10643 (N_10643,N_8748,N_8010);
or U10644 (N_10644,N_9805,N_9043);
and U10645 (N_10645,N_9949,N_8099);
nand U10646 (N_10646,N_8257,N_8576);
nor U10647 (N_10647,N_9946,N_8136);
xnor U10648 (N_10648,N_8028,N_9176);
nor U10649 (N_10649,N_9552,N_8310);
or U10650 (N_10650,N_8681,N_8373);
xnor U10651 (N_10651,N_8460,N_9673);
xnor U10652 (N_10652,N_9113,N_8647);
or U10653 (N_10653,N_9343,N_9891);
xnor U10654 (N_10654,N_9090,N_9118);
and U10655 (N_10655,N_9747,N_9663);
xor U10656 (N_10656,N_8712,N_9665);
and U10657 (N_10657,N_8773,N_8346);
nand U10658 (N_10658,N_9568,N_8033);
or U10659 (N_10659,N_8036,N_8893);
nor U10660 (N_10660,N_8272,N_8570);
or U10661 (N_10661,N_9903,N_9686);
nor U10662 (N_10662,N_9963,N_8624);
nor U10663 (N_10663,N_8685,N_9024);
nor U10664 (N_10664,N_8918,N_9298);
nand U10665 (N_10665,N_8187,N_8731);
nand U10666 (N_10666,N_9561,N_9990);
nor U10667 (N_10667,N_9293,N_9428);
and U10668 (N_10668,N_8909,N_9999);
and U10669 (N_10669,N_8115,N_9013);
nand U10670 (N_10670,N_8034,N_8172);
nand U10671 (N_10671,N_8462,N_8340);
or U10672 (N_10672,N_8891,N_8276);
and U10673 (N_10673,N_9814,N_9331);
and U10674 (N_10674,N_9235,N_8525);
and U10675 (N_10675,N_8983,N_8258);
and U10676 (N_10676,N_9400,N_9970);
and U10677 (N_10677,N_9213,N_9795);
or U10678 (N_10678,N_8518,N_9202);
or U10679 (N_10679,N_8222,N_8579);
xor U10680 (N_10680,N_9486,N_9908);
xor U10681 (N_10681,N_8545,N_9132);
nand U10682 (N_10682,N_9468,N_9417);
or U10683 (N_10683,N_8260,N_9920);
xnor U10684 (N_10684,N_8014,N_8439);
xor U10685 (N_10685,N_8285,N_9387);
and U10686 (N_10686,N_8289,N_8165);
nor U10687 (N_10687,N_9218,N_9130);
nand U10688 (N_10688,N_9503,N_9780);
xor U10689 (N_10689,N_8083,N_9656);
nand U10690 (N_10690,N_9248,N_9159);
nand U10691 (N_10691,N_8569,N_8819);
and U10692 (N_10692,N_8600,N_9072);
or U10693 (N_10693,N_9680,N_9437);
nand U10694 (N_10694,N_9399,N_9806);
nand U10695 (N_10695,N_8813,N_8662);
nor U10696 (N_10696,N_9099,N_9352);
or U10697 (N_10697,N_8453,N_9518);
and U10698 (N_10698,N_9364,N_8759);
or U10699 (N_10699,N_8861,N_8676);
nor U10700 (N_10700,N_9360,N_8716);
and U10701 (N_10701,N_8872,N_8805);
or U10702 (N_10702,N_9833,N_8236);
nor U10703 (N_10703,N_8955,N_8278);
nor U10704 (N_10704,N_8123,N_8190);
or U10705 (N_10705,N_9741,N_9655);
xor U10706 (N_10706,N_8561,N_8192);
xnor U10707 (N_10707,N_9562,N_9674);
and U10708 (N_10708,N_9153,N_8456);
nor U10709 (N_10709,N_8106,N_9783);
nor U10710 (N_10710,N_8204,N_9192);
nor U10711 (N_10711,N_8917,N_8974);
and U10712 (N_10712,N_8251,N_8379);
and U10713 (N_10713,N_9292,N_9685);
nor U10714 (N_10714,N_8639,N_9771);
nor U10715 (N_10715,N_8799,N_8375);
xor U10716 (N_10716,N_9713,N_9689);
and U10717 (N_10717,N_8727,N_9694);
nor U10718 (N_10718,N_8060,N_9111);
nor U10719 (N_10719,N_9855,N_9767);
xnor U10720 (N_10720,N_8546,N_9443);
and U10721 (N_10721,N_8932,N_9672);
and U10722 (N_10722,N_9637,N_9760);
nor U10723 (N_10723,N_8603,N_8823);
xnor U10724 (N_10724,N_8949,N_9681);
and U10725 (N_10725,N_9796,N_9000);
xnor U10726 (N_10726,N_9492,N_8907);
and U10727 (N_10727,N_8386,N_8564);
or U10728 (N_10728,N_8937,N_9403);
nand U10729 (N_10729,N_9629,N_9287);
and U10730 (N_10730,N_9125,N_8517);
xor U10731 (N_10731,N_8598,N_9831);
and U10732 (N_10732,N_9506,N_8176);
nor U10733 (N_10733,N_8769,N_9878);
nand U10734 (N_10734,N_8405,N_9286);
or U10735 (N_10735,N_9600,N_8383);
nand U10736 (N_10736,N_9348,N_9938);
or U10737 (N_10737,N_8049,N_9077);
nand U10738 (N_10738,N_8812,N_8490);
nor U10739 (N_10739,N_9627,N_8778);
nand U10740 (N_10740,N_9730,N_8205);
or U10741 (N_10741,N_8638,N_8326);
nor U10742 (N_10742,N_8971,N_8342);
xor U10743 (N_10743,N_8822,N_8070);
nand U10744 (N_10744,N_8315,N_8250);
nand U10745 (N_10745,N_9049,N_8473);
nor U10746 (N_10746,N_8304,N_8009);
nor U10747 (N_10747,N_9857,N_9940);
nor U10748 (N_10748,N_9933,N_9625);
nand U10749 (N_10749,N_9547,N_8211);
nor U10750 (N_10750,N_9461,N_9203);
and U10751 (N_10751,N_9170,N_9657);
nand U10752 (N_10752,N_8754,N_9005);
nor U10753 (N_10753,N_8920,N_8058);
nor U10754 (N_10754,N_8926,N_9432);
or U10755 (N_10755,N_8853,N_9842);
and U10756 (N_10756,N_9501,N_8098);
xnor U10757 (N_10757,N_8648,N_9794);
xor U10758 (N_10758,N_8732,N_8426);
nor U10759 (N_10759,N_9490,N_9749);
nor U10760 (N_10760,N_9670,N_9329);
nor U10761 (N_10761,N_9519,N_8240);
nor U10762 (N_10762,N_9138,N_9311);
and U10763 (N_10763,N_8325,N_9027);
or U10764 (N_10764,N_9096,N_8018);
xor U10765 (N_10765,N_8417,N_8201);
nand U10766 (N_10766,N_9156,N_8628);
or U10767 (N_10767,N_9571,N_8744);
nor U10768 (N_10768,N_8810,N_9825);
nor U10769 (N_10769,N_8319,N_8227);
nand U10770 (N_10770,N_8641,N_8921);
and U10771 (N_10771,N_8411,N_9011);
and U10772 (N_10772,N_9206,N_9807);
and U10773 (N_10773,N_9269,N_9785);
xnor U10774 (N_10774,N_8163,N_8322);
and U10775 (N_10775,N_8102,N_8428);
xnor U10776 (N_10776,N_8848,N_9968);
nand U10777 (N_10777,N_9744,N_8677);
xnor U10778 (N_10778,N_8841,N_8252);
xor U10779 (N_10779,N_8474,N_8513);
xor U10780 (N_10780,N_9511,N_8052);
or U10781 (N_10781,N_9424,N_8901);
or U10782 (N_10782,N_9584,N_8745);
or U10783 (N_10783,N_9106,N_8479);
nor U10784 (N_10784,N_8481,N_9313);
and U10785 (N_10785,N_9057,N_8402);
and U10786 (N_10786,N_9018,N_9421);
and U10787 (N_10787,N_8843,N_8844);
and U10788 (N_10788,N_9911,N_9275);
and U10789 (N_10789,N_9499,N_8294);
xnor U10790 (N_10790,N_9575,N_8225);
nand U10791 (N_10791,N_9314,N_9557);
nand U10792 (N_10792,N_8419,N_8374);
nor U10793 (N_10793,N_8348,N_9761);
nand U10794 (N_10794,N_8329,N_8504);
nand U10795 (N_10795,N_9255,N_8178);
xor U10796 (N_10796,N_8482,N_8697);
nand U10797 (N_10797,N_8210,N_8875);
and U10798 (N_10798,N_9015,N_9535);
nand U10799 (N_10799,N_8077,N_9321);
or U10800 (N_10800,N_8720,N_9359);
nor U10801 (N_10801,N_9972,N_9485);
and U10802 (N_10802,N_8605,N_9472);
nand U10803 (N_10803,N_9190,N_9083);
xor U10804 (N_10804,N_8847,N_8888);
nand U10805 (N_10805,N_8020,N_8230);
nand U10806 (N_10806,N_8717,N_8764);
or U10807 (N_10807,N_8622,N_9868);
nor U10808 (N_10808,N_8292,N_8963);
or U10809 (N_10809,N_9696,N_8166);
xnor U10810 (N_10810,N_8508,N_9723);
nand U10811 (N_10811,N_9419,N_8741);
nor U10812 (N_10812,N_8599,N_9914);
xor U10813 (N_10813,N_8392,N_9631);
nand U10814 (N_10814,N_8017,N_8215);
xnor U10815 (N_10815,N_8064,N_9489);
nor U10816 (N_10816,N_8519,N_9838);
xnor U10817 (N_10817,N_8311,N_9133);
nand U10818 (N_10818,N_9374,N_8722);
nand U10819 (N_10819,N_8345,N_9086);
or U10820 (N_10820,N_9295,N_8254);
xnor U10821 (N_10821,N_8037,N_8082);
or U10822 (N_10822,N_8936,N_9797);
nand U10823 (N_10823,N_8768,N_9734);
nor U10824 (N_10824,N_9746,N_8689);
and U10825 (N_10825,N_9658,N_9762);
and U10826 (N_10826,N_9541,N_8357);
and U10827 (N_10827,N_8217,N_9453);
xor U10828 (N_10828,N_8330,N_9046);
or U10829 (N_10829,N_9932,N_8725);
or U10830 (N_10830,N_9659,N_8248);
nor U10831 (N_10831,N_8737,N_8393);
nand U10832 (N_10832,N_8468,N_8779);
xor U10833 (N_10833,N_8255,N_9652);
xnor U10834 (N_10834,N_8973,N_9804);
or U10835 (N_10835,N_8275,N_8596);
and U10836 (N_10836,N_9966,N_8135);
or U10837 (N_10837,N_9323,N_9095);
or U10838 (N_10838,N_9752,N_9936);
or U10839 (N_10839,N_8787,N_8931);
xor U10840 (N_10840,N_8195,N_8743);
xor U10841 (N_10841,N_9879,N_8616);
xor U10842 (N_10842,N_9906,N_8399);
xnor U10843 (N_10843,N_8048,N_8902);
nand U10844 (N_10844,N_8111,N_8335);
nor U10845 (N_10845,N_8341,N_9608);
nand U10846 (N_10846,N_8469,N_8487);
or U10847 (N_10847,N_8855,N_8088);
nor U10848 (N_10848,N_8719,N_9603);
xnor U10849 (N_10849,N_8062,N_8876);
xor U10850 (N_10850,N_8076,N_8788);
nor U10851 (N_10851,N_8485,N_8388);
nor U10852 (N_10852,N_9146,N_9845);
xnor U10853 (N_10853,N_8080,N_8699);
nor U10854 (N_10854,N_9078,N_8131);
xnor U10855 (N_10855,N_9887,N_9697);
xor U10856 (N_10856,N_8571,N_8159);
nor U10857 (N_10857,N_9808,N_9418);
nand U10858 (N_10858,N_9006,N_8900);
nor U10859 (N_10859,N_8991,N_8780);
or U10860 (N_10860,N_9242,N_8125);
and U10861 (N_10861,N_8118,N_8551);
and U10862 (N_10862,N_8370,N_9210);
and U10863 (N_10863,N_9445,N_9945);
xnor U10864 (N_10864,N_9589,N_8536);
or U10865 (N_10865,N_9126,N_9479);
nor U10866 (N_10866,N_9209,N_8935);
or U10867 (N_10867,N_9554,N_8372);
nand U10868 (N_10868,N_8449,N_8063);
xnor U10869 (N_10869,N_9528,N_8053);
or U10870 (N_10870,N_8919,N_9097);
or U10871 (N_10871,N_9917,N_8833);
nor U10872 (N_10872,N_9969,N_8167);
and U10873 (N_10873,N_8849,N_9110);
and U10874 (N_10874,N_8967,N_9446);
or U10875 (N_10875,N_8263,N_9597);
or U10876 (N_10876,N_9244,N_9300);
and U10877 (N_10877,N_8556,N_8554);
nor U10878 (N_10878,N_8944,N_8756);
or U10879 (N_10879,N_8522,N_8757);
nor U10880 (N_10880,N_9372,N_8798);
and U10881 (N_10881,N_8801,N_9245);
nand U10882 (N_10882,N_9163,N_9382);
nand U10883 (N_10883,N_8507,N_8924);
and U10884 (N_10884,N_8565,N_8594);
nand U10885 (N_10885,N_9889,N_9837);
or U10886 (N_10886,N_8515,N_8606);
and U10887 (N_10887,N_9738,N_9069);
and U10888 (N_10888,N_9791,N_9822);
and U10889 (N_10889,N_8261,N_9016);
and U10890 (N_10890,N_9976,N_8268);
xor U10891 (N_10891,N_9669,N_8360);
nor U10892 (N_10892,N_9279,N_8116);
or U10893 (N_10893,N_9219,N_9241);
and U10894 (N_10894,N_9002,N_9705);
nor U10895 (N_10895,N_8353,N_9250);
and U10896 (N_10896,N_8679,N_9409);
nand U10897 (N_10897,N_9030,N_8378);
and U10898 (N_10898,N_9211,N_9508);
xor U10899 (N_10899,N_8864,N_9493);
and U10900 (N_10900,N_8283,N_9173);
and U10901 (N_10901,N_9164,N_8338);
xor U10902 (N_10902,N_8524,N_8164);
or U10903 (N_10903,N_8815,N_8868);
nand U10904 (N_10904,N_8721,N_8557);
nor U10905 (N_10905,N_9507,N_8897);
or U10906 (N_10906,N_8194,N_8711);
or U10907 (N_10907,N_8238,N_9522);
and U10908 (N_10908,N_9774,N_8259);
xor U10909 (N_10909,N_9850,N_8188);
nand U10910 (N_10910,N_8365,N_9029);
nor U10911 (N_10911,N_9053,N_8008);
nand U10912 (N_10912,N_9546,N_8286);
and U10913 (N_10913,N_8035,N_9361);
nand U10914 (N_10914,N_9939,N_9008);
nand U10915 (N_10915,N_8910,N_8693);
nand U10916 (N_10916,N_9649,N_8445);
and U10917 (N_10917,N_8075,N_8661);
and U10918 (N_10918,N_8997,N_8869);
nand U10919 (N_10919,N_8265,N_9056);
or U10920 (N_10920,N_8177,N_9386);
xor U10921 (N_10921,N_8669,N_9103);
or U10922 (N_10922,N_8709,N_9993);
nand U10923 (N_10923,N_8547,N_9634);
nor U10924 (N_10924,N_9128,N_8095);
and U10925 (N_10925,N_9317,N_8312);
xor U10926 (N_10926,N_8544,N_8749);
or U10927 (N_10927,N_9175,N_8249);
nor U10928 (N_10928,N_8882,N_8146);
or U10929 (N_10929,N_8602,N_9954);
or U10930 (N_10930,N_8590,N_9840);
nor U10931 (N_10931,N_9704,N_8954);
and U10932 (N_10932,N_8269,N_9058);
or U10933 (N_10933,N_9185,N_9870);
nand U10934 (N_10934,N_9276,N_9745);
or U10935 (N_10935,N_8480,N_9643);
nand U10936 (N_10936,N_8203,N_9294);
and U10937 (N_10937,N_9447,N_8657);
or U10938 (N_10938,N_9092,N_8804);
nor U10939 (N_10939,N_9405,N_9262);
or U10940 (N_10940,N_8979,N_8858);
xor U10941 (N_10941,N_8421,N_8817);
nand U10942 (N_10942,N_8840,N_9285);
xor U10943 (N_10943,N_9227,N_8680);
nand U10944 (N_10944,N_8887,N_8103);
nand U10945 (N_10945,N_9260,N_8939);
nand U10946 (N_10946,N_8454,N_9392);
and U10947 (N_10947,N_8644,N_9189);
nand U10948 (N_10948,N_8629,N_8358);
and U10949 (N_10949,N_8127,N_9471);
xor U10950 (N_10950,N_9291,N_9962);
nand U10951 (N_10951,N_8995,N_9299);
nand U10952 (N_10952,N_9509,N_8718);
or U10953 (N_10953,N_8496,N_9179);
nor U10954 (N_10954,N_9178,N_8636);
nor U10955 (N_10955,N_8878,N_8852);
xor U10956 (N_10956,N_8144,N_8297);
nand U10957 (N_10957,N_9142,N_9404);
xnor U10958 (N_10958,N_8789,N_9776);
xor U10959 (N_10959,N_9975,N_9415);
xnor U10960 (N_10960,N_8271,N_9536);
and U10961 (N_10961,N_9560,N_9458);
nor U10962 (N_10962,N_9935,N_9944);
and U10963 (N_10963,N_8213,N_8183);
or U10964 (N_10964,N_9678,N_9922);
or U10965 (N_10965,N_9204,N_9566);
and U10966 (N_10966,N_8814,N_9899);
nand U10967 (N_10967,N_8300,N_8171);
nor U10968 (N_10968,N_8079,N_8003);
nor U10969 (N_10969,N_9188,N_8992);
nor U10970 (N_10970,N_8395,N_8637);
xor U10971 (N_10971,N_9450,N_8105);
nor U10972 (N_10972,N_9367,N_9452);
nor U10973 (N_10973,N_8152,N_8714);
and U10974 (N_10974,N_8885,N_8774);
nor U10975 (N_10975,N_9022,N_9302);
or U10976 (N_10976,N_8244,N_8200);
nand U10977 (N_10977,N_9772,N_9459);
or U10978 (N_10978,N_8057,N_8025);
xnor U10979 (N_10979,N_8612,N_8279);
nand U10980 (N_10980,N_8951,N_8880);
nor U10981 (N_10981,N_8708,N_8087);
and U10982 (N_10982,N_8349,N_9412);
nand U10983 (N_10983,N_8535,N_9166);
nor U10984 (N_10984,N_9080,N_9624);
nand U10985 (N_10985,N_8837,N_9394);
xor U10986 (N_10986,N_8724,N_8976);
or U10987 (N_10987,N_9326,N_8396);
nor U10988 (N_10988,N_8226,N_9754);
and U10989 (N_10989,N_9422,N_9578);
nor U10990 (N_10990,N_9102,N_9154);
or U10991 (N_10991,N_8443,N_9345);
and U10992 (N_10992,N_8981,N_8994);
and U10993 (N_10993,N_9239,N_9832);
and U10994 (N_10994,N_8871,N_8444);
or U10995 (N_10995,N_9721,N_8630);
xor U10996 (N_10996,N_8934,N_8169);
or U10997 (N_10997,N_8447,N_8972);
nand U10998 (N_10998,N_8046,N_9194);
xnor U10999 (N_10999,N_9515,N_8898);
and U11000 (N_11000,N_9924,N_8861);
nand U11001 (N_11001,N_8609,N_8708);
xor U11002 (N_11002,N_9699,N_9790);
and U11003 (N_11003,N_9911,N_8399);
nor U11004 (N_11004,N_8857,N_9545);
nor U11005 (N_11005,N_9193,N_8684);
and U11006 (N_11006,N_9649,N_9470);
or U11007 (N_11007,N_8053,N_9225);
or U11008 (N_11008,N_9526,N_8113);
or U11009 (N_11009,N_9114,N_9032);
and U11010 (N_11010,N_9596,N_9505);
nand U11011 (N_11011,N_8464,N_8175);
or U11012 (N_11012,N_9336,N_8574);
and U11013 (N_11013,N_8835,N_9450);
xnor U11014 (N_11014,N_8517,N_9848);
and U11015 (N_11015,N_9651,N_9846);
or U11016 (N_11016,N_9668,N_9229);
nand U11017 (N_11017,N_8661,N_8471);
xnor U11018 (N_11018,N_9352,N_8002);
or U11019 (N_11019,N_9016,N_9758);
and U11020 (N_11020,N_9649,N_8832);
and U11021 (N_11021,N_8451,N_8859);
nand U11022 (N_11022,N_9267,N_9537);
xnor U11023 (N_11023,N_8998,N_8293);
and U11024 (N_11024,N_9164,N_8482);
xor U11025 (N_11025,N_8121,N_9245);
nor U11026 (N_11026,N_8827,N_8469);
xnor U11027 (N_11027,N_9231,N_9195);
or U11028 (N_11028,N_9377,N_9936);
or U11029 (N_11029,N_9816,N_8636);
or U11030 (N_11030,N_9748,N_9407);
nor U11031 (N_11031,N_9158,N_9966);
xnor U11032 (N_11032,N_8568,N_9583);
and U11033 (N_11033,N_9858,N_9380);
nor U11034 (N_11034,N_9120,N_9840);
nand U11035 (N_11035,N_9325,N_8573);
nor U11036 (N_11036,N_8690,N_8493);
nand U11037 (N_11037,N_9819,N_8641);
nor U11038 (N_11038,N_8697,N_8376);
or U11039 (N_11039,N_9098,N_8308);
nand U11040 (N_11040,N_9490,N_9531);
nand U11041 (N_11041,N_9769,N_8796);
nor U11042 (N_11042,N_9542,N_9365);
or U11043 (N_11043,N_8961,N_9513);
xor U11044 (N_11044,N_8902,N_8365);
xnor U11045 (N_11045,N_9922,N_8190);
and U11046 (N_11046,N_8051,N_8765);
or U11047 (N_11047,N_9913,N_9272);
nor U11048 (N_11048,N_8034,N_8913);
nor U11049 (N_11049,N_9036,N_8363);
or U11050 (N_11050,N_9828,N_8715);
nand U11051 (N_11051,N_9409,N_8944);
and U11052 (N_11052,N_9938,N_8444);
nand U11053 (N_11053,N_9101,N_9994);
xor U11054 (N_11054,N_9052,N_9688);
nor U11055 (N_11055,N_9802,N_8858);
or U11056 (N_11056,N_9505,N_8218);
and U11057 (N_11057,N_9230,N_9268);
or U11058 (N_11058,N_8107,N_9143);
and U11059 (N_11059,N_8803,N_8129);
or U11060 (N_11060,N_9534,N_8052);
xnor U11061 (N_11061,N_8444,N_8486);
nand U11062 (N_11062,N_8276,N_8105);
xor U11063 (N_11063,N_8170,N_9991);
nor U11064 (N_11064,N_8828,N_9987);
or U11065 (N_11065,N_9807,N_8000);
xor U11066 (N_11066,N_8839,N_9862);
nand U11067 (N_11067,N_9053,N_9083);
and U11068 (N_11068,N_8999,N_8774);
nor U11069 (N_11069,N_8605,N_9966);
and U11070 (N_11070,N_9811,N_9812);
xnor U11071 (N_11071,N_8490,N_8986);
and U11072 (N_11072,N_9718,N_9642);
nor U11073 (N_11073,N_8414,N_8406);
xnor U11074 (N_11074,N_9426,N_8604);
or U11075 (N_11075,N_8061,N_8770);
or U11076 (N_11076,N_8227,N_8188);
and U11077 (N_11077,N_8301,N_9829);
xor U11078 (N_11078,N_9126,N_9138);
nand U11079 (N_11079,N_8791,N_8852);
nor U11080 (N_11080,N_8206,N_8553);
or U11081 (N_11081,N_8379,N_9822);
nor U11082 (N_11082,N_9185,N_8309);
or U11083 (N_11083,N_8952,N_8081);
nor U11084 (N_11084,N_9669,N_8336);
xor U11085 (N_11085,N_8838,N_8934);
or U11086 (N_11086,N_8018,N_9853);
nand U11087 (N_11087,N_8022,N_9333);
nor U11088 (N_11088,N_8523,N_8948);
or U11089 (N_11089,N_9483,N_8046);
nor U11090 (N_11090,N_8520,N_8590);
nor U11091 (N_11091,N_9845,N_8694);
or U11092 (N_11092,N_8712,N_9994);
and U11093 (N_11093,N_9136,N_9793);
xor U11094 (N_11094,N_8653,N_8414);
and U11095 (N_11095,N_9589,N_9054);
or U11096 (N_11096,N_8757,N_8094);
nand U11097 (N_11097,N_9113,N_8868);
nand U11098 (N_11098,N_9561,N_8301);
and U11099 (N_11099,N_9141,N_8616);
nand U11100 (N_11100,N_8147,N_8932);
xnor U11101 (N_11101,N_8948,N_8729);
nand U11102 (N_11102,N_8433,N_8490);
nand U11103 (N_11103,N_8662,N_8529);
or U11104 (N_11104,N_9786,N_8118);
xor U11105 (N_11105,N_9805,N_9440);
and U11106 (N_11106,N_8036,N_8105);
xnor U11107 (N_11107,N_8748,N_8180);
or U11108 (N_11108,N_8673,N_9201);
nor U11109 (N_11109,N_9340,N_9482);
or U11110 (N_11110,N_8505,N_9890);
and U11111 (N_11111,N_9354,N_8287);
nand U11112 (N_11112,N_9915,N_8314);
or U11113 (N_11113,N_8090,N_9032);
nand U11114 (N_11114,N_8381,N_8334);
nor U11115 (N_11115,N_8440,N_9589);
xnor U11116 (N_11116,N_8608,N_9111);
nand U11117 (N_11117,N_9501,N_8525);
xor U11118 (N_11118,N_9501,N_9221);
nand U11119 (N_11119,N_9757,N_9534);
nor U11120 (N_11120,N_8288,N_8370);
nor U11121 (N_11121,N_8396,N_8613);
and U11122 (N_11122,N_8310,N_8240);
or U11123 (N_11123,N_8698,N_8996);
or U11124 (N_11124,N_8229,N_9414);
xor U11125 (N_11125,N_8701,N_9503);
nand U11126 (N_11126,N_8595,N_8852);
and U11127 (N_11127,N_8301,N_9957);
nand U11128 (N_11128,N_8802,N_9657);
nor U11129 (N_11129,N_9861,N_8530);
and U11130 (N_11130,N_9934,N_8997);
or U11131 (N_11131,N_9408,N_8336);
nand U11132 (N_11132,N_8367,N_8223);
nor U11133 (N_11133,N_8437,N_9163);
and U11134 (N_11134,N_8245,N_9307);
and U11135 (N_11135,N_8472,N_9522);
nand U11136 (N_11136,N_9736,N_9960);
xnor U11137 (N_11137,N_8736,N_8555);
nand U11138 (N_11138,N_8013,N_8044);
nor U11139 (N_11139,N_9894,N_9184);
nor U11140 (N_11140,N_8038,N_8139);
xor U11141 (N_11141,N_9440,N_8058);
and U11142 (N_11142,N_8236,N_8273);
and U11143 (N_11143,N_9308,N_8834);
or U11144 (N_11144,N_8134,N_8876);
nand U11145 (N_11145,N_8201,N_9972);
xor U11146 (N_11146,N_9269,N_8003);
and U11147 (N_11147,N_8208,N_8596);
nand U11148 (N_11148,N_9126,N_9442);
or U11149 (N_11149,N_9756,N_9492);
nor U11150 (N_11150,N_8498,N_8737);
xnor U11151 (N_11151,N_8366,N_9070);
or U11152 (N_11152,N_9617,N_9880);
nor U11153 (N_11153,N_8942,N_9416);
or U11154 (N_11154,N_9134,N_8480);
xor U11155 (N_11155,N_8611,N_8635);
nor U11156 (N_11156,N_9337,N_8630);
xor U11157 (N_11157,N_9118,N_8417);
nand U11158 (N_11158,N_8668,N_9881);
or U11159 (N_11159,N_9371,N_9225);
nor U11160 (N_11160,N_8548,N_8777);
nor U11161 (N_11161,N_9155,N_8245);
nor U11162 (N_11162,N_9128,N_9486);
xnor U11163 (N_11163,N_9196,N_8574);
nor U11164 (N_11164,N_9352,N_8021);
xnor U11165 (N_11165,N_9650,N_9303);
and U11166 (N_11166,N_9552,N_9831);
nand U11167 (N_11167,N_8200,N_9751);
and U11168 (N_11168,N_8545,N_8204);
and U11169 (N_11169,N_8036,N_8063);
nor U11170 (N_11170,N_9200,N_8857);
nor U11171 (N_11171,N_8188,N_9228);
and U11172 (N_11172,N_9136,N_9957);
and U11173 (N_11173,N_9572,N_8608);
or U11174 (N_11174,N_9843,N_8362);
and U11175 (N_11175,N_8422,N_8066);
and U11176 (N_11176,N_9381,N_9915);
nand U11177 (N_11177,N_8022,N_9082);
or U11178 (N_11178,N_8349,N_9770);
or U11179 (N_11179,N_9349,N_9976);
or U11180 (N_11180,N_8303,N_9635);
nor U11181 (N_11181,N_8605,N_9978);
and U11182 (N_11182,N_9114,N_9424);
nand U11183 (N_11183,N_9633,N_9617);
and U11184 (N_11184,N_9368,N_8426);
or U11185 (N_11185,N_8370,N_8416);
nand U11186 (N_11186,N_8279,N_9605);
nand U11187 (N_11187,N_9959,N_8548);
or U11188 (N_11188,N_9599,N_9551);
or U11189 (N_11189,N_8283,N_8777);
and U11190 (N_11190,N_9997,N_8141);
nor U11191 (N_11191,N_9492,N_9082);
nor U11192 (N_11192,N_8820,N_9753);
and U11193 (N_11193,N_8364,N_8309);
or U11194 (N_11194,N_8521,N_9451);
xnor U11195 (N_11195,N_9071,N_9415);
and U11196 (N_11196,N_9160,N_8798);
nor U11197 (N_11197,N_9389,N_9489);
nor U11198 (N_11198,N_8533,N_8364);
or U11199 (N_11199,N_9496,N_9075);
nor U11200 (N_11200,N_8673,N_9223);
or U11201 (N_11201,N_9687,N_9274);
or U11202 (N_11202,N_8013,N_8370);
and U11203 (N_11203,N_8170,N_9450);
and U11204 (N_11204,N_8467,N_8302);
nand U11205 (N_11205,N_9532,N_9436);
nor U11206 (N_11206,N_8824,N_9826);
nand U11207 (N_11207,N_8579,N_8701);
xor U11208 (N_11208,N_8404,N_9412);
and U11209 (N_11209,N_8969,N_8644);
or U11210 (N_11210,N_9988,N_9950);
or U11211 (N_11211,N_9915,N_8327);
nor U11212 (N_11212,N_9992,N_9679);
nor U11213 (N_11213,N_9412,N_9789);
xnor U11214 (N_11214,N_8176,N_8723);
nor U11215 (N_11215,N_8278,N_9768);
xnor U11216 (N_11216,N_8749,N_9422);
or U11217 (N_11217,N_9206,N_9115);
nor U11218 (N_11218,N_9418,N_8669);
and U11219 (N_11219,N_8437,N_8953);
and U11220 (N_11220,N_9549,N_8890);
or U11221 (N_11221,N_9816,N_8460);
or U11222 (N_11222,N_9498,N_8149);
or U11223 (N_11223,N_9041,N_8048);
nor U11224 (N_11224,N_8428,N_9415);
nand U11225 (N_11225,N_8118,N_8030);
xnor U11226 (N_11226,N_8359,N_9413);
xnor U11227 (N_11227,N_9715,N_8340);
or U11228 (N_11228,N_9713,N_9188);
and U11229 (N_11229,N_9516,N_8225);
and U11230 (N_11230,N_8537,N_8242);
or U11231 (N_11231,N_8230,N_9601);
and U11232 (N_11232,N_9946,N_9983);
xnor U11233 (N_11233,N_8557,N_9599);
nor U11234 (N_11234,N_8025,N_8102);
and U11235 (N_11235,N_8959,N_9072);
nor U11236 (N_11236,N_8815,N_9817);
nand U11237 (N_11237,N_9033,N_9188);
xor U11238 (N_11238,N_8773,N_8191);
xor U11239 (N_11239,N_9251,N_8145);
xnor U11240 (N_11240,N_8846,N_8259);
nand U11241 (N_11241,N_8779,N_9238);
xnor U11242 (N_11242,N_8701,N_8464);
xor U11243 (N_11243,N_9086,N_9576);
nand U11244 (N_11244,N_8795,N_9748);
nor U11245 (N_11245,N_9411,N_8320);
and U11246 (N_11246,N_8578,N_8568);
nor U11247 (N_11247,N_8411,N_8046);
and U11248 (N_11248,N_9023,N_9971);
or U11249 (N_11249,N_8073,N_9210);
or U11250 (N_11250,N_8282,N_8892);
nand U11251 (N_11251,N_9152,N_8494);
xor U11252 (N_11252,N_8347,N_9813);
and U11253 (N_11253,N_9830,N_8520);
nor U11254 (N_11254,N_9199,N_8143);
and U11255 (N_11255,N_8290,N_9281);
and U11256 (N_11256,N_8313,N_8344);
nand U11257 (N_11257,N_8601,N_9533);
and U11258 (N_11258,N_8643,N_9740);
nor U11259 (N_11259,N_8806,N_9383);
or U11260 (N_11260,N_9220,N_8018);
or U11261 (N_11261,N_8893,N_9969);
nor U11262 (N_11262,N_8720,N_9718);
and U11263 (N_11263,N_8176,N_9184);
or U11264 (N_11264,N_8816,N_8181);
or U11265 (N_11265,N_9203,N_8147);
nand U11266 (N_11266,N_8654,N_9152);
or U11267 (N_11267,N_9319,N_9487);
xnor U11268 (N_11268,N_9653,N_8393);
or U11269 (N_11269,N_8140,N_9443);
and U11270 (N_11270,N_9490,N_9413);
xnor U11271 (N_11271,N_9226,N_8114);
nor U11272 (N_11272,N_9892,N_8645);
or U11273 (N_11273,N_8174,N_9592);
nand U11274 (N_11274,N_8772,N_8062);
nand U11275 (N_11275,N_8105,N_8601);
nor U11276 (N_11276,N_8823,N_8161);
xor U11277 (N_11277,N_9726,N_8879);
xor U11278 (N_11278,N_8832,N_9074);
or U11279 (N_11279,N_9153,N_8235);
and U11280 (N_11280,N_9768,N_9760);
and U11281 (N_11281,N_8751,N_8371);
or U11282 (N_11282,N_9026,N_8229);
xor U11283 (N_11283,N_9615,N_9112);
or U11284 (N_11284,N_9907,N_8593);
and U11285 (N_11285,N_8201,N_9248);
nor U11286 (N_11286,N_8665,N_9042);
or U11287 (N_11287,N_8570,N_8650);
xor U11288 (N_11288,N_9898,N_9477);
and U11289 (N_11289,N_9502,N_9641);
and U11290 (N_11290,N_8666,N_9961);
and U11291 (N_11291,N_9577,N_9412);
xnor U11292 (N_11292,N_8559,N_8527);
or U11293 (N_11293,N_8000,N_8047);
or U11294 (N_11294,N_8413,N_8372);
nor U11295 (N_11295,N_9619,N_9902);
nand U11296 (N_11296,N_9790,N_9163);
xnor U11297 (N_11297,N_8149,N_8860);
and U11298 (N_11298,N_8850,N_8877);
or U11299 (N_11299,N_9419,N_8343);
or U11300 (N_11300,N_8476,N_9079);
or U11301 (N_11301,N_9845,N_9203);
and U11302 (N_11302,N_8906,N_9573);
and U11303 (N_11303,N_8817,N_9732);
xor U11304 (N_11304,N_9010,N_8605);
or U11305 (N_11305,N_9622,N_8253);
or U11306 (N_11306,N_8022,N_8004);
xnor U11307 (N_11307,N_9570,N_8559);
and U11308 (N_11308,N_9051,N_8718);
xor U11309 (N_11309,N_9336,N_9832);
nand U11310 (N_11310,N_9547,N_9430);
and U11311 (N_11311,N_9811,N_8674);
xnor U11312 (N_11312,N_8327,N_9739);
or U11313 (N_11313,N_9199,N_8974);
nor U11314 (N_11314,N_8225,N_8224);
nor U11315 (N_11315,N_8910,N_8250);
nor U11316 (N_11316,N_9360,N_9856);
and U11317 (N_11317,N_9765,N_8492);
and U11318 (N_11318,N_8787,N_8571);
xor U11319 (N_11319,N_8398,N_9769);
nor U11320 (N_11320,N_9165,N_9444);
and U11321 (N_11321,N_9094,N_9931);
nand U11322 (N_11322,N_9593,N_9533);
or U11323 (N_11323,N_9051,N_8464);
or U11324 (N_11324,N_8394,N_8593);
nand U11325 (N_11325,N_9033,N_8884);
nor U11326 (N_11326,N_9512,N_8528);
nor U11327 (N_11327,N_9609,N_9582);
nand U11328 (N_11328,N_9174,N_9332);
and U11329 (N_11329,N_9653,N_9836);
nor U11330 (N_11330,N_9372,N_8971);
and U11331 (N_11331,N_8032,N_8242);
nor U11332 (N_11332,N_8675,N_9007);
xor U11333 (N_11333,N_8971,N_9863);
nor U11334 (N_11334,N_8058,N_8226);
and U11335 (N_11335,N_8795,N_8645);
nor U11336 (N_11336,N_9867,N_8103);
or U11337 (N_11337,N_8948,N_9546);
or U11338 (N_11338,N_8716,N_9272);
xor U11339 (N_11339,N_9950,N_8949);
and U11340 (N_11340,N_9095,N_9113);
xor U11341 (N_11341,N_9313,N_9772);
nor U11342 (N_11342,N_8067,N_8213);
or U11343 (N_11343,N_9490,N_8819);
nand U11344 (N_11344,N_9881,N_8859);
and U11345 (N_11345,N_9651,N_8380);
or U11346 (N_11346,N_9972,N_8343);
and U11347 (N_11347,N_8876,N_8495);
or U11348 (N_11348,N_9343,N_8641);
and U11349 (N_11349,N_8280,N_9707);
nor U11350 (N_11350,N_9789,N_9073);
or U11351 (N_11351,N_8692,N_8577);
or U11352 (N_11352,N_8903,N_8721);
nor U11353 (N_11353,N_9452,N_9282);
and U11354 (N_11354,N_9046,N_9893);
and U11355 (N_11355,N_8001,N_9160);
or U11356 (N_11356,N_9986,N_8336);
or U11357 (N_11357,N_8477,N_9920);
or U11358 (N_11358,N_8474,N_9122);
nor U11359 (N_11359,N_8488,N_9861);
nand U11360 (N_11360,N_8241,N_8083);
nor U11361 (N_11361,N_9735,N_8987);
xor U11362 (N_11362,N_8980,N_8195);
and U11363 (N_11363,N_8392,N_8007);
and U11364 (N_11364,N_9709,N_9174);
nand U11365 (N_11365,N_9189,N_8661);
nand U11366 (N_11366,N_8013,N_8158);
nand U11367 (N_11367,N_8330,N_8548);
or U11368 (N_11368,N_9321,N_9176);
or U11369 (N_11369,N_8969,N_8383);
and U11370 (N_11370,N_9211,N_8353);
xnor U11371 (N_11371,N_9979,N_9144);
nor U11372 (N_11372,N_9642,N_8884);
xnor U11373 (N_11373,N_9820,N_9687);
and U11374 (N_11374,N_9352,N_8298);
and U11375 (N_11375,N_8110,N_9972);
or U11376 (N_11376,N_8805,N_9841);
nand U11377 (N_11377,N_8266,N_8979);
or U11378 (N_11378,N_8368,N_9564);
xor U11379 (N_11379,N_8691,N_8604);
and U11380 (N_11380,N_8751,N_8675);
or U11381 (N_11381,N_9381,N_9551);
nand U11382 (N_11382,N_8920,N_8756);
or U11383 (N_11383,N_8444,N_8757);
nand U11384 (N_11384,N_8376,N_9055);
nor U11385 (N_11385,N_8052,N_8939);
xnor U11386 (N_11386,N_8588,N_8151);
nand U11387 (N_11387,N_9399,N_8483);
nor U11388 (N_11388,N_9555,N_9015);
and U11389 (N_11389,N_9724,N_8535);
or U11390 (N_11390,N_8407,N_9455);
and U11391 (N_11391,N_9727,N_8269);
xor U11392 (N_11392,N_8146,N_8039);
nor U11393 (N_11393,N_9649,N_8355);
xor U11394 (N_11394,N_8455,N_9468);
nor U11395 (N_11395,N_8168,N_8637);
nor U11396 (N_11396,N_8972,N_9601);
and U11397 (N_11397,N_8741,N_8141);
xnor U11398 (N_11398,N_9372,N_9307);
nor U11399 (N_11399,N_9868,N_8950);
xnor U11400 (N_11400,N_8686,N_8620);
nor U11401 (N_11401,N_8581,N_8061);
xor U11402 (N_11402,N_9313,N_9350);
nand U11403 (N_11403,N_9165,N_9548);
nor U11404 (N_11404,N_8660,N_8407);
xnor U11405 (N_11405,N_9896,N_8599);
or U11406 (N_11406,N_8152,N_8834);
nor U11407 (N_11407,N_8018,N_9107);
and U11408 (N_11408,N_8218,N_9522);
or U11409 (N_11409,N_8055,N_9694);
xnor U11410 (N_11410,N_8570,N_9791);
nor U11411 (N_11411,N_8819,N_8700);
and U11412 (N_11412,N_9634,N_9834);
nand U11413 (N_11413,N_8363,N_9256);
nor U11414 (N_11414,N_8093,N_9579);
xor U11415 (N_11415,N_9558,N_8169);
or U11416 (N_11416,N_9437,N_9075);
nor U11417 (N_11417,N_9706,N_8210);
or U11418 (N_11418,N_8739,N_9701);
or U11419 (N_11419,N_9437,N_9417);
xnor U11420 (N_11420,N_9447,N_9499);
xnor U11421 (N_11421,N_9889,N_9034);
and U11422 (N_11422,N_9174,N_9504);
xor U11423 (N_11423,N_8375,N_8029);
or U11424 (N_11424,N_9029,N_9988);
or U11425 (N_11425,N_9698,N_9968);
or U11426 (N_11426,N_9843,N_8132);
or U11427 (N_11427,N_9872,N_8757);
nor U11428 (N_11428,N_8585,N_8654);
and U11429 (N_11429,N_8839,N_8920);
xnor U11430 (N_11430,N_9650,N_9048);
nand U11431 (N_11431,N_9201,N_8911);
and U11432 (N_11432,N_8320,N_9456);
or U11433 (N_11433,N_9819,N_9245);
or U11434 (N_11434,N_9201,N_8119);
nand U11435 (N_11435,N_9848,N_8082);
and U11436 (N_11436,N_8084,N_9937);
or U11437 (N_11437,N_8550,N_8840);
or U11438 (N_11438,N_9148,N_9006);
nor U11439 (N_11439,N_9840,N_9891);
nor U11440 (N_11440,N_8754,N_8125);
or U11441 (N_11441,N_8874,N_8547);
nand U11442 (N_11442,N_9985,N_8361);
xor U11443 (N_11443,N_8289,N_9015);
xnor U11444 (N_11444,N_8753,N_8179);
nand U11445 (N_11445,N_8189,N_9502);
or U11446 (N_11446,N_9482,N_8676);
or U11447 (N_11447,N_9391,N_8005);
xor U11448 (N_11448,N_9861,N_8218);
nand U11449 (N_11449,N_8474,N_8231);
nor U11450 (N_11450,N_8496,N_8841);
and U11451 (N_11451,N_8583,N_8790);
nand U11452 (N_11452,N_8932,N_8873);
nand U11453 (N_11453,N_8592,N_9126);
nor U11454 (N_11454,N_9536,N_9724);
and U11455 (N_11455,N_9670,N_9160);
xor U11456 (N_11456,N_8267,N_8512);
nand U11457 (N_11457,N_8264,N_9272);
or U11458 (N_11458,N_8485,N_8122);
and U11459 (N_11459,N_9341,N_8904);
nor U11460 (N_11460,N_9773,N_8843);
and U11461 (N_11461,N_9453,N_9812);
and U11462 (N_11462,N_8038,N_8105);
or U11463 (N_11463,N_9087,N_9497);
or U11464 (N_11464,N_9727,N_9985);
nand U11465 (N_11465,N_9051,N_9821);
nor U11466 (N_11466,N_9313,N_8820);
xor U11467 (N_11467,N_9007,N_8583);
or U11468 (N_11468,N_8937,N_9642);
xnor U11469 (N_11469,N_9638,N_8272);
and U11470 (N_11470,N_9842,N_9064);
and U11471 (N_11471,N_9775,N_8983);
nand U11472 (N_11472,N_8566,N_9216);
nor U11473 (N_11473,N_9957,N_8630);
or U11474 (N_11474,N_9133,N_9201);
or U11475 (N_11475,N_8087,N_8605);
xnor U11476 (N_11476,N_8847,N_8172);
nor U11477 (N_11477,N_8378,N_8492);
xor U11478 (N_11478,N_8973,N_8407);
and U11479 (N_11479,N_9319,N_8058);
xnor U11480 (N_11480,N_8693,N_9323);
nor U11481 (N_11481,N_8732,N_8910);
nand U11482 (N_11482,N_8706,N_8543);
nand U11483 (N_11483,N_9642,N_8020);
nor U11484 (N_11484,N_9152,N_9118);
nor U11485 (N_11485,N_8400,N_9449);
xnor U11486 (N_11486,N_9147,N_8151);
or U11487 (N_11487,N_8563,N_8842);
and U11488 (N_11488,N_9493,N_8555);
xor U11489 (N_11489,N_9100,N_9328);
or U11490 (N_11490,N_9784,N_9566);
or U11491 (N_11491,N_9768,N_9585);
nor U11492 (N_11492,N_8806,N_9952);
or U11493 (N_11493,N_8622,N_8074);
xor U11494 (N_11494,N_8500,N_8471);
or U11495 (N_11495,N_9096,N_8456);
nor U11496 (N_11496,N_9118,N_9496);
nand U11497 (N_11497,N_9516,N_9222);
nor U11498 (N_11498,N_8562,N_8251);
or U11499 (N_11499,N_9191,N_9454);
or U11500 (N_11500,N_9408,N_8130);
xnor U11501 (N_11501,N_9357,N_8119);
nor U11502 (N_11502,N_8043,N_8808);
nor U11503 (N_11503,N_8201,N_9428);
nand U11504 (N_11504,N_9108,N_8642);
xor U11505 (N_11505,N_8533,N_8436);
xor U11506 (N_11506,N_8204,N_8988);
nor U11507 (N_11507,N_9414,N_9391);
and U11508 (N_11508,N_9734,N_8961);
or U11509 (N_11509,N_9362,N_9086);
nor U11510 (N_11510,N_8592,N_9896);
and U11511 (N_11511,N_9116,N_9489);
nor U11512 (N_11512,N_9111,N_8581);
nand U11513 (N_11513,N_9657,N_8259);
and U11514 (N_11514,N_9237,N_9372);
nor U11515 (N_11515,N_9222,N_8026);
xor U11516 (N_11516,N_9563,N_8903);
or U11517 (N_11517,N_9436,N_8064);
xnor U11518 (N_11518,N_8713,N_9569);
xor U11519 (N_11519,N_8950,N_8834);
nor U11520 (N_11520,N_8001,N_8317);
and U11521 (N_11521,N_9948,N_9849);
nand U11522 (N_11522,N_8030,N_9949);
nand U11523 (N_11523,N_8032,N_9467);
and U11524 (N_11524,N_9936,N_8775);
and U11525 (N_11525,N_9682,N_9447);
nand U11526 (N_11526,N_8563,N_8829);
and U11527 (N_11527,N_8022,N_8342);
nor U11528 (N_11528,N_8719,N_8383);
nor U11529 (N_11529,N_8949,N_8973);
or U11530 (N_11530,N_9368,N_9827);
xor U11531 (N_11531,N_9249,N_8092);
nand U11532 (N_11532,N_8131,N_9121);
nor U11533 (N_11533,N_9095,N_9206);
or U11534 (N_11534,N_9814,N_9829);
and U11535 (N_11535,N_8642,N_9791);
xor U11536 (N_11536,N_8048,N_9602);
xnor U11537 (N_11537,N_9735,N_8960);
and U11538 (N_11538,N_8615,N_9404);
and U11539 (N_11539,N_8826,N_9853);
nor U11540 (N_11540,N_8952,N_9283);
nand U11541 (N_11541,N_9864,N_8162);
and U11542 (N_11542,N_8599,N_9642);
or U11543 (N_11543,N_8487,N_8667);
or U11544 (N_11544,N_9274,N_9506);
nand U11545 (N_11545,N_8178,N_9347);
nor U11546 (N_11546,N_9827,N_8878);
or U11547 (N_11547,N_8508,N_9664);
xnor U11548 (N_11548,N_9218,N_8134);
nor U11549 (N_11549,N_8765,N_8707);
or U11550 (N_11550,N_8843,N_8592);
nand U11551 (N_11551,N_8716,N_8815);
and U11552 (N_11552,N_8254,N_9947);
nor U11553 (N_11553,N_9116,N_8930);
or U11554 (N_11554,N_8430,N_8746);
and U11555 (N_11555,N_8730,N_8821);
nand U11556 (N_11556,N_9583,N_9294);
and U11557 (N_11557,N_9773,N_8235);
xor U11558 (N_11558,N_8367,N_9371);
or U11559 (N_11559,N_9234,N_9629);
nand U11560 (N_11560,N_8089,N_8341);
and U11561 (N_11561,N_9239,N_9790);
or U11562 (N_11562,N_9651,N_8927);
and U11563 (N_11563,N_8668,N_8030);
xnor U11564 (N_11564,N_9628,N_8569);
or U11565 (N_11565,N_8697,N_9813);
nand U11566 (N_11566,N_9143,N_8191);
nand U11567 (N_11567,N_8104,N_9545);
nor U11568 (N_11568,N_8855,N_8166);
xor U11569 (N_11569,N_9414,N_8662);
nand U11570 (N_11570,N_9556,N_9487);
or U11571 (N_11571,N_8001,N_9002);
xor U11572 (N_11572,N_9926,N_9869);
and U11573 (N_11573,N_8892,N_9504);
xor U11574 (N_11574,N_8131,N_9511);
nor U11575 (N_11575,N_9791,N_9051);
nor U11576 (N_11576,N_9191,N_9020);
or U11577 (N_11577,N_8398,N_8004);
xor U11578 (N_11578,N_8843,N_9430);
nand U11579 (N_11579,N_8252,N_9160);
xnor U11580 (N_11580,N_8002,N_8989);
xor U11581 (N_11581,N_8712,N_8404);
and U11582 (N_11582,N_9261,N_8303);
xor U11583 (N_11583,N_9357,N_9955);
nand U11584 (N_11584,N_9651,N_8140);
or U11585 (N_11585,N_8195,N_8994);
and U11586 (N_11586,N_8185,N_9576);
and U11587 (N_11587,N_9567,N_8952);
nor U11588 (N_11588,N_9332,N_9485);
xor U11589 (N_11589,N_9434,N_8715);
or U11590 (N_11590,N_9251,N_9580);
and U11591 (N_11591,N_8400,N_8355);
nand U11592 (N_11592,N_9468,N_8843);
nand U11593 (N_11593,N_9496,N_9138);
and U11594 (N_11594,N_8524,N_8682);
nand U11595 (N_11595,N_9624,N_8539);
xnor U11596 (N_11596,N_9871,N_8450);
nand U11597 (N_11597,N_8745,N_9906);
or U11598 (N_11598,N_8036,N_8202);
nor U11599 (N_11599,N_8191,N_9122);
nand U11600 (N_11600,N_8235,N_9543);
or U11601 (N_11601,N_9138,N_8502);
xor U11602 (N_11602,N_8026,N_8244);
and U11603 (N_11603,N_9947,N_9709);
nor U11604 (N_11604,N_9491,N_9876);
nand U11605 (N_11605,N_8610,N_8905);
xor U11606 (N_11606,N_8184,N_9677);
and U11607 (N_11607,N_8317,N_8799);
xnor U11608 (N_11608,N_9801,N_9856);
and U11609 (N_11609,N_9714,N_9693);
nand U11610 (N_11610,N_9677,N_8354);
and U11611 (N_11611,N_8090,N_9950);
or U11612 (N_11612,N_8723,N_9925);
or U11613 (N_11613,N_9753,N_9482);
and U11614 (N_11614,N_8689,N_9335);
nand U11615 (N_11615,N_8284,N_9611);
xnor U11616 (N_11616,N_9403,N_9959);
nand U11617 (N_11617,N_9413,N_9172);
nand U11618 (N_11618,N_8540,N_9949);
or U11619 (N_11619,N_9232,N_8913);
xor U11620 (N_11620,N_9750,N_9248);
nand U11621 (N_11621,N_9476,N_9278);
xor U11622 (N_11622,N_8997,N_9702);
nand U11623 (N_11623,N_8025,N_8592);
or U11624 (N_11624,N_9594,N_8605);
nand U11625 (N_11625,N_8234,N_9516);
and U11626 (N_11626,N_9891,N_9686);
nand U11627 (N_11627,N_9462,N_9212);
nor U11628 (N_11628,N_9385,N_9801);
nor U11629 (N_11629,N_8877,N_9527);
and U11630 (N_11630,N_8597,N_8497);
and U11631 (N_11631,N_8902,N_9588);
or U11632 (N_11632,N_8213,N_9214);
xor U11633 (N_11633,N_9643,N_9160);
or U11634 (N_11634,N_8889,N_8184);
nand U11635 (N_11635,N_9006,N_8656);
nor U11636 (N_11636,N_9305,N_9577);
and U11637 (N_11637,N_8136,N_8905);
and U11638 (N_11638,N_8330,N_8229);
nand U11639 (N_11639,N_8336,N_8519);
or U11640 (N_11640,N_8152,N_8329);
and U11641 (N_11641,N_9107,N_8154);
xnor U11642 (N_11642,N_8035,N_9915);
or U11643 (N_11643,N_9933,N_9738);
nor U11644 (N_11644,N_9597,N_9643);
nor U11645 (N_11645,N_8313,N_8684);
and U11646 (N_11646,N_8816,N_9135);
xor U11647 (N_11647,N_9305,N_9413);
and U11648 (N_11648,N_9185,N_9110);
or U11649 (N_11649,N_8075,N_9636);
xor U11650 (N_11650,N_9743,N_8865);
nor U11651 (N_11651,N_9801,N_9354);
nor U11652 (N_11652,N_8412,N_8835);
nand U11653 (N_11653,N_8480,N_9262);
and U11654 (N_11654,N_8480,N_9978);
xor U11655 (N_11655,N_8760,N_9506);
and U11656 (N_11656,N_9847,N_8300);
nor U11657 (N_11657,N_8526,N_8788);
or U11658 (N_11658,N_9444,N_9079);
nand U11659 (N_11659,N_8412,N_8183);
nor U11660 (N_11660,N_9385,N_9844);
xnor U11661 (N_11661,N_9602,N_9625);
xor U11662 (N_11662,N_8361,N_9362);
xnor U11663 (N_11663,N_8367,N_8904);
xor U11664 (N_11664,N_9210,N_9831);
nand U11665 (N_11665,N_8487,N_9160);
or U11666 (N_11666,N_8900,N_9576);
or U11667 (N_11667,N_8441,N_9103);
nor U11668 (N_11668,N_9452,N_9534);
nor U11669 (N_11669,N_9069,N_9752);
or U11670 (N_11670,N_8365,N_8919);
xor U11671 (N_11671,N_9226,N_9851);
nand U11672 (N_11672,N_8331,N_9010);
or U11673 (N_11673,N_9465,N_9541);
xnor U11674 (N_11674,N_8061,N_8920);
xor U11675 (N_11675,N_8178,N_8664);
nand U11676 (N_11676,N_9032,N_9027);
nor U11677 (N_11677,N_8783,N_9146);
and U11678 (N_11678,N_9809,N_8840);
nand U11679 (N_11679,N_8215,N_8966);
xor U11680 (N_11680,N_9932,N_8105);
nand U11681 (N_11681,N_9143,N_8211);
nand U11682 (N_11682,N_8454,N_8580);
nor U11683 (N_11683,N_9554,N_8904);
xnor U11684 (N_11684,N_9900,N_8936);
or U11685 (N_11685,N_8271,N_8651);
nand U11686 (N_11686,N_8657,N_9675);
xnor U11687 (N_11687,N_8148,N_9242);
xor U11688 (N_11688,N_8878,N_8295);
and U11689 (N_11689,N_9105,N_8085);
and U11690 (N_11690,N_9154,N_9767);
and U11691 (N_11691,N_8055,N_9370);
and U11692 (N_11692,N_8027,N_9081);
xor U11693 (N_11693,N_8513,N_8468);
nor U11694 (N_11694,N_8604,N_9677);
nor U11695 (N_11695,N_9210,N_8001);
or U11696 (N_11696,N_8041,N_9160);
or U11697 (N_11697,N_9465,N_9090);
nand U11698 (N_11698,N_9342,N_9793);
nor U11699 (N_11699,N_8295,N_9616);
nor U11700 (N_11700,N_9179,N_9694);
and U11701 (N_11701,N_9419,N_9512);
xnor U11702 (N_11702,N_9993,N_8763);
and U11703 (N_11703,N_8620,N_9762);
nor U11704 (N_11704,N_8964,N_8993);
and U11705 (N_11705,N_8726,N_9215);
xnor U11706 (N_11706,N_8614,N_9536);
and U11707 (N_11707,N_8468,N_8469);
xnor U11708 (N_11708,N_8096,N_8477);
nand U11709 (N_11709,N_8095,N_9294);
nand U11710 (N_11710,N_8516,N_8256);
nand U11711 (N_11711,N_9995,N_8677);
nor U11712 (N_11712,N_9024,N_8121);
nand U11713 (N_11713,N_8045,N_8235);
and U11714 (N_11714,N_9652,N_8480);
or U11715 (N_11715,N_9233,N_9822);
nand U11716 (N_11716,N_9719,N_8306);
and U11717 (N_11717,N_8846,N_8546);
nand U11718 (N_11718,N_8258,N_8704);
and U11719 (N_11719,N_9531,N_9069);
xnor U11720 (N_11720,N_8287,N_9405);
nand U11721 (N_11721,N_9363,N_8714);
or U11722 (N_11722,N_8703,N_9309);
xnor U11723 (N_11723,N_8039,N_8059);
or U11724 (N_11724,N_9786,N_9157);
and U11725 (N_11725,N_8143,N_8442);
nand U11726 (N_11726,N_9943,N_9988);
or U11727 (N_11727,N_8626,N_8198);
xor U11728 (N_11728,N_8793,N_8004);
nor U11729 (N_11729,N_9000,N_8571);
or U11730 (N_11730,N_9621,N_8733);
xor U11731 (N_11731,N_8753,N_8915);
or U11732 (N_11732,N_9843,N_8198);
nor U11733 (N_11733,N_9591,N_8051);
xnor U11734 (N_11734,N_8258,N_9971);
nor U11735 (N_11735,N_9320,N_9253);
nand U11736 (N_11736,N_8633,N_9271);
or U11737 (N_11737,N_9945,N_8771);
xnor U11738 (N_11738,N_9343,N_8262);
nor U11739 (N_11739,N_8577,N_8185);
and U11740 (N_11740,N_8348,N_8460);
and U11741 (N_11741,N_9140,N_8171);
and U11742 (N_11742,N_8138,N_8272);
nor U11743 (N_11743,N_8918,N_9079);
nand U11744 (N_11744,N_9067,N_8880);
and U11745 (N_11745,N_8389,N_9676);
and U11746 (N_11746,N_8153,N_8252);
and U11747 (N_11747,N_9069,N_8507);
or U11748 (N_11748,N_8882,N_9207);
or U11749 (N_11749,N_9108,N_9149);
xnor U11750 (N_11750,N_8431,N_9507);
and U11751 (N_11751,N_9190,N_9995);
and U11752 (N_11752,N_8540,N_8560);
or U11753 (N_11753,N_8413,N_9834);
xnor U11754 (N_11754,N_8610,N_8536);
and U11755 (N_11755,N_8599,N_8383);
nand U11756 (N_11756,N_8195,N_9590);
nor U11757 (N_11757,N_8388,N_9504);
xnor U11758 (N_11758,N_9588,N_9526);
nor U11759 (N_11759,N_9201,N_8547);
or U11760 (N_11760,N_8925,N_9226);
xnor U11761 (N_11761,N_8161,N_8316);
or U11762 (N_11762,N_9928,N_9764);
xnor U11763 (N_11763,N_9810,N_8707);
xor U11764 (N_11764,N_9110,N_9621);
xor U11765 (N_11765,N_9617,N_8347);
or U11766 (N_11766,N_8381,N_9529);
xnor U11767 (N_11767,N_9909,N_9999);
xor U11768 (N_11768,N_8814,N_8636);
nand U11769 (N_11769,N_8667,N_8807);
and U11770 (N_11770,N_9696,N_9429);
nor U11771 (N_11771,N_9911,N_8516);
nand U11772 (N_11772,N_8670,N_8851);
nand U11773 (N_11773,N_9138,N_9977);
xor U11774 (N_11774,N_9449,N_8151);
nand U11775 (N_11775,N_8321,N_8692);
nor U11776 (N_11776,N_8661,N_9348);
nand U11777 (N_11777,N_8719,N_8032);
and U11778 (N_11778,N_8494,N_9686);
xnor U11779 (N_11779,N_9616,N_8274);
xnor U11780 (N_11780,N_8047,N_9391);
xnor U11781 (N_11781,N_8701,N_8914);
nand U11782 (N_11782,N_9144,N_8914);
xnor U11783 (N_11783,N_8888,N_9858);
nor U11784 (N_11784,N_9072,N_8586);
nor U11785 (N_11785,N_8842,N_9678);
xnor U11786 (N_11786,N_9264,N_9334);
xnor U11787 (N_11787,N_8441,N_8111);
xor U11788 (N_11788,N_9614,N_8599);
xor U11789 (N_11789,N_8220,N_9123);
or U11790 (N_11790,N_8680,N_8804);
nor U11791 (N_11791,N_8564,N_8951);
nor U11792 (N_11792,N_8821,N_8787);
or U11793 (N_11793,N_8789,N_9675);
nand U11794 (N_11794,N_9592,N_8850);
nor U11795 (N_11795,N_8350,N_8786);
or U11796 (N_11796,N_9549,N_8945);
nand U11797 (N_11797,N_8656,N_9972);
and U11798 (N_11798,N_9088,N_9068);
nor U11799 (N_11799,N_9806,N_9504);
or U11800 (N_11800,N_9533,N_8837);
nor U11801 (N_11801,N_8323,N_9823);
nand U11802 (N_11802,N_8625,N_9904);
and U11803 (N_11803,N_8225,N_8981);
or U11804 (N_11804,N_9620,N_8578);
or U11805 (N_11805,N_9504,N_8630);
xnor U11806 (N_11806,N_8767,N_8816);
nand U11807 (N_11807,N_8605,N_9088);
and U11808 (N_11808,N_8181,N_9490);
nor U11809 (N_11809,N_9396,N_8891);
xor U11810 (N_11810,N_8321,N_8706);
or U11811 (N_11811,N_9312,N_9818);
nand U11812 (N_11812,N_8998,N_8197);
and U11813 (N_11813,N_9455,N_8675);
xnor U11814 (N_11814,N_8612,N_8809);
xor U11815 (N_11815,N_9385,N_9691);
and U11816 (N_11816,N_9862,N_8923);
nor U11817 (N_11817,N_8212,N_9910);
and U11818 (N_11818,N_9892,N_9885);
xor U11819 (N_11819,N_8207,N_9290);
or U11820 (N_11820,N_8945,N_9360);
nor U11821 (N_11821,N_8918,N_9270);
or U11822 (N_11822,N_9902,N_8334);
or U11823 (N_11823,N_8526,N_8346);
nand U11824 (N_11824,N_8513,N_9055);
xnor U11825 (N_11825,N_9653,N_9850);
nand U11826 (N_11826,N_8012,N_8624);
nand U11827 (N_11827,N_9715,N_8674);
nand U11828 (N_11828,N_9366,N_8773);
nor U11829 (N_11829,N_8447,N_9170);
nor U11830 (N_11830,N_9828,N_9586);
and U11831 (N_11831,N_9577,N_9434);
nor U11832 (N_11832,N_8416,N_9766);
and U11833 (N_11833,N_9894,N_8309);
or U11834 (N_11834,N_8005,N_9687);
nor U11835 (N_11835,N_9322,N_9896);
or U11836 (N_11836,N_9596,N_8120);
nor U11837 (N_11837,N_9277,N_8980);
and U11838 (N_11838,N_8910,N_9995);
xnor U11839 (N_11839,N_9980,N_9815);
nor U11840 (N_11840,N_9193,N_9891);
xor U11841 (N_11841,N_9810,N_9213);
xnor U11842 (N_11842,N_8872,N_9699);
nand U11843 (N_11843,N_8404,N_9335);
nand U11844 (N_11844,N_8105,N_9282);
nor U11845 (N_11845,N_8504,N_8877);
nor U11846 (N_11846,N_8992,N_8079);
and U11847 (N_11847,N_8968,N_9939);
nor U11848 (N_11848,N_9936,N_9360);
xor U11849 (N_11849,N_9619,N_9293);
xor U11850 (N_11850,N_8997,N_8542);
or U11851 (N_11851,N_9668,N_8355);
nand U11852 (N_11852,N_9986,N_9062);
and U11853 (N_11853,N_8047,N_9922);
and U11854 (N_11854,N_9439,N_9302);
or U11855 (N_11855,N_9022,N_8448);
or U11856 (N_11856,N_8905,N_8437);
xnor U11857 (N_11857,N_9622,N_8080);
nand U11858 (N_11858,N_9363,N_9310);
nor U11859 (N_11859,N_9566,N_9233);
xor U11860 (N_11860,N_9259,N_8843);
nor U11861 (N_11861,N_8552,N_8038);
or U11862 (N_11862,N_8545,N_9715);
nor U11863 (N_11863,N_8331,N_9721);
nor U11864 (N_11864,N_8143,N_8963);
or U11865 (N_11865,N_9730,N_8889);
and U11866 (N_11866,N_9809,N_8430);
and U11867 (N_11867,N_9831,N_9941);
or U11868 (N_11868,N_8980,N_8201);
nor U11869 (N_11869,N_9495,N_8675);
nor U11870 (N_11870,N_8118,N_8156);
nor U11871 (N_11871,N_8037,N_8031);
nor U11872 (N_11872,N_9235,N_9533);
and U11873 (N_11873,N_9691,N_8267);
xor U11874 (N_11874,N_9918,N_9230);
nand U11875 (N_11875,N_8309,N_9023);
nand U11876 (N_11876,N_9637,N_8483);
nand U11877 (N_11877,N_8604,N_8627);
nor U11878 (N_11878,N_8902,N_8503);
nand U11879 (N_11879,N_8901,N_8698);
and U11880 (N_11880,N_9913,N_8891);
and U11881 (N_11881,N_9650,N_8958);
nand U11882 (N_11882,N_9749,N_9401);
xor U11883 (N_11883,N_8855,N_8564);
nand U11884 (N_11884,N_8943,N_9592);
nand U11885 (N_11885,N_8886,N_8930);
or U11886 (N_11886,N_9600,N_9011);
and U11887 (N_11887,N_8618,N_9943);
or U11888 (N_11888,N_8537,N_9166);
or U11889 (N_11889,N_9994,N_9444);
and U11890 (N_11890,N_9586,N_9425);
xnor U11891 (N_11891,N_9466,N_9613);
nand U11892 (N_11892,N_9569,N_8971);
xnor U11893 (N_11893,N_9767,N_9539);
nand U11894 (N_11894,N_8107,N_9920);
xor U11895 (N_11895,N_9835,N_8675);
or U11896 (N_11896,N_9151,N_8475);
nor U11897 (N_11897,N_9476,N_8678);
nand U11898 (N_11898,N_9072,N_9696);
and U11899 (N_11899,N_8666,N_9153);
and U11900 (N_11900,N_9140,N_8978);
xor U11901 (N_11901,N_9843,N_8207);
or U11902 (N_11902,N_9138,N_8255);
nand U11903 (N_11903,N_8105,N_9355);
and U11904 (N_11904,N_9787,N_8075);
and U11905 (N_11905,N_9615,N_8846);
xor U11906 (N_11906,N_8936,N_9050);
or U11907 (N_11907,N_9436,N_8576);
or U11908 (N_11908,N_8768,N_9642);
xor U11909 (N_11909,N_8877,N_8635);
xor U11910 (N_11910,N_9888,N_9660);
or U11911 (N_11911,N_9052,N_9356);
nor U11912 (N_11912,N_8140,N_9043);
xnor U11913 (N_11913,N_9572,N_8402);
nand U11914 (N_11914,N_8848,N_8255);
nor U11915 (N_11915,N_8417,N_9683);
nor U11916 (N_11916,N_8165,N_8328);
or U11917 (N_11917,N_8067,N_8884);
nor U11918 (N_11918,N_8184,N_8232);
or U11919 (N_11919,N_8728,N_8709);
and U11920 (N_11920,N_9591,N_9830);
and U11921 (N_11921,N_9108,N_8881);
xnor U11922 (N_11922,N_8022,N_9663);
nand U11923 (N_11923,N_8022,N_9522);
xnor U11924 (N_11924,N_8372,N_8680);
nand U11925 (N_11925,N_8023,N_8200);
xnor U11926 (N_11926,N_8687,N_8352);
or U11927 (N_11927,N_9761,N_8917);
and U11928 (N_11928,N_8946,N_8327);
nand U11929 (N_11929,N_9820,N_8762);
xor U11930 (N_11930,N_9787,N_9075);
nor U11931 (N_11931,N_8386,N_8760);
or U11932 (N_11932,N_8583,N_9273);
or U11933 (N_11933,N_8174,N_9150);
nand U11934 (N_11934,N_9569,N_8301);
or U11935 (N_11935,N_9104,N_8980);
xor U11936 (N_11936,N_9630,N_9607);
xor U11937 (N_11937,N_8389,N_9408);
xnor U11938 (N_11938,N_9048,N_8522);
nor U11939 (N_11939,N_9352,N_9318);
nand U11940 (N_11940,N_8954,N_9471);
xor U11941 (N_11941,N_8848,N_8168);
nand U11942 (N_11942,N_9069,N_8080);
or U11943 (N_11943,N_8954,N_9048);
nor U11944 (N_11944,N_8212,N_9083);
or U11945 (N_11945,N_9927,N_8798);
nand U11946 (N_11946,N_8307,N_8095);
or U11947 (N_11947,N_8667,N_9717);
and U11948 (N_11948,N_9899,N_8888);
and U11949 (N_11949,N_9379,N_8297);
nor U11950 (N_11950,N_8983,N_9028);
or U11951 (N_11951,N_8719,N_8232);
xor U11952 (N_11952,N_8334,N_8177);
or U11953 (N_11953,N_9134,N_8634);
and U11954 (N_11954,N_8865,N_8597);
or U11955 (N_11955,N_9031,N_8882);
and U11956 (N_11956,N_8122,N_8432);
xor U11957 (N_11957,N_8769,N_9028);
xnor U11958 (N_11958,N_9063,N_9626);
nor U11959 (N_11959,N_8868,N_8499);
nand U11960 (N_11960,N_8510,N_9116);
nand U11961 (N_11961,N_8212,N_9462);
xnor U11962 (N_11962,N_8466,N_8796);
nor U11963 (N_11963,N_8418,N_9601);
nor U11964 (N_11964,N_8832,N_8542);
or U11965 (N_11965,N_9077,N_9549);
xor U11966 (N_11966,N_9596,N_9419);
and U11967 (N_11967,N_8808,N_8145);
or U11968 (N_11968,N_8525,N_8014);
or U11969 (N_11969,N_8613,N_9346);
or U11970 (N_11970,N_9672,N_8253);
nand U11971 (N_11971,N_9097,N_8528);
and U11972 (N_11972,N_8927,N_8395);
and U11973 (N_11973,N_9535,N_8285);
nand U11974 (N_11974,N_8665,N_9028);
nor U11975 (N_11975,N_8424,N_9426);
or U11976 (N_11976,N_9123,N_8942);
or U11977 (N_11977,N_9494,N_8579);
nor U11978 (N_11978,N_8445,N_8405);
or U11979 (N_11979,N_9108,N_9595);
or U11980 (N_11980,N_9555,N_9315);
and U11981 (N_11981,N_9661,N_9622);
or U11982 (N_11982,N_9938,N_9278);
and U11983 (N_11983,N_8693,N_8610);
or U11984 (N_11984,N_9399,N_9195);
xor U11985 (N_11985,N_9849,N_8474);
and U11986 (N_11986,N_8935,N_8750);
or U11987 (N_11987,N_9330,N_9116);
nand U11988 (N_11988,N_9626,N_9141);
and U11989 (N_11989,N_9175,N_8817);
nor U11990 (N_11990,N_8003,N_8563);
nor U11991 (N_11991,N_8626,N_9762);
nor U11992 (N_11992,N_8578,N_8149);
xor U11993 (N_11993,N_8333,N_8024);
nand U11994 (N_11994,N_9468,N_9388);
nand U11995 (N_11995,N_8979,N_8664);
and U11996 (N_11996,N_8776,N_9364);
nor U11997 (N_11997,N_9484,N_9296);
or U11998 (N_11998,N_9030,N_8411);
and U11999 (N_11999,N_8013,N_9927);
or U12000 (N_12000,N_11737,N_10242);
and U12001 (N_12001,N_10597,N_11527);
xnor U12002 (N_12002,N_10924,N_10295);
nand U12003 (N_12003,N_10887,N_10133);
and U12004 (N_12004,N_11670,N_11101);
or U12005 (N_12005,N_10021,N_10656);
nor U12006 (N_12006,N_10284,N_11439);
nor U12007 (N_12007,N_10640,N_10759);
xnor U12008 (N_12008,N_11650,N_10197);
and U12009 (N_12009,N_11074,N_10010);
xnor U12010 (N_12010,N_10661,N_10081);
xnor U12011 (N_12011,N_11771,N_11192);
nor U12012 (N_12012,N_11788,N_11599);
or U12013 (N_12013,N_11346,N_11573);
nand U12014 (N_12014,N_11172,N_10884);
nand U12015 (N_12015,N_10613,N_10076);
nand U12016 (N_12016,N_11732,N_10317);
nor U12017 (N_12017,N_10020,N_11994);
or U12018 (N_12018,N_10904,N_11025);
nand U12019 (N_12019,N_10420,N_11225);
and U12020 (N_12020,N_10775,N_11575);
xor U12021 (N_12021,N_10356,N_11106);
nand U12022 (N_12022,N_10294,N_11161);
or U12023 (N_12023,N_10310,N_10390);
nor U12024 (N_12024,N_11468,N_11924);
nand U12025 (N_12025,N_11780,N_11905);
or U12026 (N_12026,N_11504,N_11474);
or U12027 (N_12027,N_10678,N_10374);
and U12028 (N_12028,N_11729,N_11019);
or U12029 (N_12029,N_10771,N_10537);
nand U12030 (N_12030,N_11001,N_10458);
and U12031 (N_12031,N_11785,N_11290);
xor U12032 (N_12032,N_10515,N_10077);
or U12033 (N_12033,N_10300,N_10140);
nor U12034 (N_12034,N_11404,N_11183);
nand U12035 (N_12035,N_11082,N_10146);
and U12036 (N_12036,N_11093,N_10422);
nand U12037 (N_12037,N_10083,N_11634);
nor U12038 (N_12038,N_11327,N_10933);
nor U12039 (N_12039,N_10974,N_11740);
nor U12040 (N_12040,N_11015,N_11537);
nand U12041 (N_12041,N_11297,N_11705);
nand U12042 (N_12042,N_11651,N_10061);
nor U12043 (N_12043,N_10565,N_10522);
nand U12044 (N_12044,N_10503,N_11062);
or U12045 (N_12045,N_11837,N_11039);
or U12046 (N_12046,N_10105,N_10059);
nand U12047 (N_12047,N_10423,N_11860);
or U12048 (N_12048,N_11099,N_10915);
or U12049 (N_12049,N_10783,N_10540);
xor U12050 (N_12050,N_10641,N_11684);
nand U12051 (N_12051,N_11311,N_10844);
and U12052 (N_12052,N_11380,N_10541);
xnor U12053 (N_12053,N_10559,N_10820);
and U12054 (N_12054,N_10680,N_11129);
nor U12055 (N_12055,N_11087,N_10840);
or U12056 (N_12056,N_10101,N_11445);
or U12057 (N_12057,N_11350,N_10389);
nor U12058 (N_12058,N_11796,N_10094);
or U12059 (N_12059,N_10033,N_11133);
or U12060 (N_12060,N_10250,N_11873);
and U12061 (N_12061,N_10634,N_10037);
or U12062 (N_12062,N_11438,N_11772);
or U12063 (N_12063,N_11384,N_10040);
xnor U12064 (N_12064,N_10695,N_10428);
xor U12065 (N_12065,N_10504,N_10028);
xor U12066 (N_12066,N_11122,N_11556);
and U12067 (N_12067,N_11261,N_11549);
or U12068 (N_12068,N_11823,N_11826);
nor U12069 (N_12069,N_11482,N_10062);
xnor U12070 (N_12070,N_11494,N_10237);
xor U12071 (N_12071,N_11375,N_11031);
nand U12072 (N_12072,N_10805,N_10139);
or U12073 (N_12073,N_10404,N_10756);
xnor U12074 (N_12074,N_11601,N_10829);
and U12075 (N_12075,N_10411,N_10527);
xnor U12076 (N_12076,N_10311,N_10777);
nand U12077 (N_12077,N_10985,N_11047);
or U12078 (N_12078,N_10425,N_10681);
nand U12079 (N_12079,N_10211,N_11876);
or U12080 (N_12080,N_11509,N_10700);
nor U12081 (N_12081,N_10757,N_11703);
xnor U12082 (N_12082,N_10267,N_10693);
nor U12083 (N_12083,N_10470,N_11529);
and U12084 (N_12084,N_10176,N_10270);
and U12085 (N_12085,N_11927,N_10705);
and U12086 (N_12086,N_10684,N_11888);
nand U12087 (N_12087,N_11516,N_10457);
nor U12088 (N_12088,N_11535,N_11464);
nor U12089 (N_12089,N_10851,N_10203);
or U12090 (N_12090,N_11953,N_10223);
nand U12091 (N_12091,N_11950,N_11797);
nor U12092 (N_12092,N_10943,N_11802);
nor U12093 (N_12093,N_11613,N_10058);
nand U12094 (N_12094,N_11263,N_10654);
or U12095 (N_12095,N_11518,N_10660);
and U12096 (N_12096,N_10912,N_10630);
or U12097 (N_12097,N_10362,N_11248);
and U12098 (N_12098,N_10750,N_10898);
or U12099 (N_12099,N_10536,N_10408);
nand U12100 (N_12100,N_11429,N_10120);
nor U12101 (N_12101,N_10792,N_11783);
xor U12102 (N_12102,N_11661,N_11965);
nand U12103 (N_12103,N_11760,N_10970);
nand U12104 (N_12104,N_11154,N_10627);
nand U12105 (N_12105,N_11774,N_10967);
xnor U12106 (N_12106,N_11954,N_11228);
or U12107 (N_12107,N_11368,N_11523);
xnor U12108 (N_12108,N_10254,N_11997);
xnor U12109 (N_12109,N_10155,N_10670);
xor U12110 (N_12110,N_10762,N_10834);
nor U12111 (N_12111,N_10372,N_10165);
or U12112 (N_12112,N_10196,N_11461);
and U12113 (N_12113,N_10490,N_10174);
nand U12114 (N_12114,N_11653,N_11528);
nor U12115 (N_12115,N_11621,N_10566);
and U12116 (N_12116,N_11815,N_11757);
nor U12117 (N_12117,N_11726,N_11655);
xor U12118 (N_12118,N_11937,N_11483);
and U12119 (N_12119,N_11071,N_11289);
nor U12120 (N_12120,N_10357,N_10532);
nor U12121 (N_12121,N_11394,N_10774);
nand U12122 (N_12122,N_11120,N_10012);
or U12123 (N_12123,N_11301,N_11676);
nor U12124 (N_12124,N_10817,N_10316);
nor U12125 (N_12125,N_10547,N_11486);
xnor U12126 (N_12126,N_11484,N_11711);
nor U12127 (N_12127,N_11681,N_10217);
nor U12128 (N_12128,N_10482,N_10781);
nor U12129 (N_12129,N_10534,N_10494);
nand U12130 (N_12130,N_11582,N_11677);
and U12131 (N_12131,N_10341,N_10475);
and U12132 (N_12132,N_10415,N_11807);
or U12133 (N_12133,N_10264,N_10115);
xor U12134 (N_12134,N_11231,N_11918);
nor U12135 (N_12135,N_10876,N_10618);
and U12136 (N_12136,N_11512,N_10994);
xnor U12137 (N_12137,N_11616,N_11948);
xor U12138 (N_12138,N_10435,N_11595);
nor U12139 (N_12139,N_11869,N_11018);
nor U12140 (N_12140,N_11324,N_10936);
and U12141 (N_12141,N_10694,N_11958);
and U12142 (N_12142,N_11214,N_10995);
xnor U12143 (N_12143,N_10241,N_10896);
nor U12144 (N_12144,N_10327,N_10863);
nor U12145 (N_12145,N_10309,N_11686);
or U12146 (N_12146,N_11383,N_11405);
nand U12147 (N_12147,N_11316,N_11193);
nor U12148 (N_12148,N_11447,N_11952);
nand U12149 (N_12149,N_11855,N_11386);
nand U12150 (N_12150,N_10321,N_10639);
xor U12151 (N_12151,N_11401,N_10208);
nand U12152 (N_12152,N_11020,N_10818);
nand U12153 (N_12153,N_11822,N_11237);
or U12154 (N_12154,N_11936,N_11072);
xnor U12155 (N_12155,N_10811,N_10557);
nand U12156 (N_12156,N_10132,N_11999);
nand U12157 (N_12157,N_10642,N_10170);
nand U12158 (N_12158,N_11075,N_10746);
nand U12159 (N_12159,N_10265,N_11603);
nand U12160 (N_12160,N_10438,N_10379);
nand U12161 (N_12161,N_11699,N_11867);
or U12162 (N_12162,N_10479,N_11446);
xnor U12163 (N_12163,N_10668,N_11792);
xor U12164 (N_12164,N_10652,N_11751);
and U12165 (N_12165,N_11450,N_10378);
nand U12166 (N_12166,N_10891,N_10748);
xor U12167 (N_12167,N_10214,N_10722);
and U12168 (N_12168,N_10005,N_11896);
and U12169 (N_12169,N_11803,N_10339);
xnor U12170 (N_12170,N_10169,N_11043);
xnor U12171 (N_12171,N_11479,N_11007);
nand U12172 (N_12172,N_11764,N_10869);
or U12173 (N_12173,N_11269,N_11627);
and U12174 (N_12174,N_11592,N_10688);
and U12175 (N_12175,N_10032,N_11735);
or U12176 (N_12176,N_10745,N_11647);
nand U12177 (N_12177,N_11648,N_11041);
xnor U12178 (N_12178,N_10441,N_10674);
nor U12179 (N_12179,N_10500,N_11293);
and U12180 (N_12180,N_10712,N_11220);
xor U12181 (N_12181,N_11545,N_10822);
nor U12182 (N_12182,N_10643,N_11402);
xor U12183 (N_12183,N_11755,N_11819);
nand U12184 (N_12184,N_10109,N_10809);
and U12185 (N_12185,N_11742,N_11276);
nor U12186 (N_12186,N_11871,N_11770);
or U12187 (N_12187,N_11949,N_11884);
nor U12188 (N_12188,N_10666,N_11798);
xnor U12189 (N_12189,N_10445,N_11761);
or U12190 (N_12190,N_11779,N_10434);
nand U12191 (N_12191,N_10131,N_10478);
nand U12192 (N_12192,N_10865,N_11235);
nor U12193 (N_12193,N_10864,N_10839);
and U12194 (N_12194,N_11738,N_10052);
or U12195 (N_12195,N_10355,N_10244);
or U12196 (N_12196,N_11051,N_11663);
nand U12197 (N_12197,N_11283,N_10723);
or U12198 (N_12198,N_11196,N_11310);
or U12199 (N_12199,N_11496,N_10160);
and U12200 (N_12200,N_10448,N_10766);
xnor U12201 (N_12201,N_11899,N_10859);
or U12202 (N_12202,N_10855,N_11393);
nand U12203 (N_12203,N_11672,N_10554);
nand U12204 (N_12204,N_10204,N_10392);
and U12205 (N_12205,N_10516,N_10779);
or U12206 (N_12206,N_11233,N_10591);
nand U12207 (N_12207,N_10182,N_10215);
or U12208 (N_12208,N_10477,N_11594);
nor U12209 (N_12209,N_11268,N_11136);
nand U12210 (N_12210,N_11983,N_10138);
nand U12211 (N_12211,N_10535,N_10741);
or U12212 (N_12212,N_10041,N_11178);
nand U12213 (N_12213,N_11148,N_10826);
nand U12214 (N_12214,N_10524,N_10736);
or U12215 (N_12215,N_10509,N_10137);
or U12216 (N_12216,N_10075,N_11448);
or U12217 (N_12217,N_11305,N_11959);
nand U12218 (N_12218,N_11619,N_10773);
or U12219 (N_12219,N_11636,N_10605);
and U12220 (N_12220,N_11414,N_10624);
or U12221 (N_12221,N_10397,N_11841);
xor U12222 (N_12222,N_11804,N_11278);
and U12223 (N_12223,N_10272,N_10814);
and U12224 (N_12224,N_11548,N_11546);
and U12225 (N_12225,N_11578,N_11799);
xnor U12226 (N_12226,N_10786,N_11832);
or U12227 (N_12227,N_11107,N_11462);
nand U12228 (N_12228,N_11519,N_10025);
and U12229 (N_12229,N_11165,N_10417);
and U12230 (N_12230,N_10584,N_11333);
or U12231 (N_12231,N_10134,N_11789);
xnor U12232 (N_12232,N_10628,N_10108);
nor U12233 (N_12233,N_11100,N_10953);
nor U12234 (N_12234,N_10796,N_11622);
nand U12235 (N_12235,N_10276,N_10446);
nand U12236 (N_12236,N_10269,N_11849);
or U12237 (N_12237,N_11715,N_11662);
nor U12238 (N_12238,N_10709,N_11469);
nand U12239 (N_12239,N_11682,N_11530);
and U12240 (N_12240,N_11141,N_10489);
nand U12241 (N_12241,N_11270,N_11877);
nand U12242 (N_12242,N_11978,N_10246);
nand U12243 (N_12243,N_10332,N_10292);
and U12244 (N_12244,N_11168,N_11149);
nand U12245 (N_12245,N_10699,N_10400);
and U12246 (N_12246,N_11294,N_10258);
nor U12247 (N_12247,N_10171,N_10381);
or U12248 (N_12248,N_11862,N_11046);
xnor U12249 (N_12249,N_10523,N_10430);
nor U12250 (N_12250,N_11554,N_10533);
or U12251 (N_12251,N_11126,N_11265);
and U12252 (N_12252,N_11252,N_11159);
nand U12253 (N_12253,N_11188,N_11880);
or U12254 (N_12254,N_11315,N_10572);
nand U12255 (N_12255,N_10049,N_10401);
xor U12256 (N_12256,N_10825,N_10560);
xnor U12257 (N_12257,N_10222,N_10191);
nand U12258 (N_12258,N_11692,N_11369);
or U12259 (N_12259,N_10180,N_11810);
nor U12260 (N_12260,N_10949,N_11531);
nor U12261 (N_12261,N_10626,N_11202);
nand U12262 (N_12262,N_11969,N_10439);
nor U12263 (N_12263,N_11717,N_10307);
xnor U12264 (N_12264,N_11045,N_11274);
nand U12265 (N_12265,N_10261,N_10177);
nand U12266 (N_12266,N_11646,N_10073);
nand U12267 (N_12267,N_10271,N_11396);
xor U12268 (N_12268,N_10905,N_10658);
nand U12269 (N_12269,N_10808,N_11164);
nor U12270 (N_12270,N_10645,N_10892);
xnor U12271 (N_12271,N_11190,N_11702);
or U12272 (N_12272,N_11088,N_10333);
or U12273 (N_12273,N_10277,N_11866);
nor U12274 (N_12274,N_11977,N_11037);
or U12275 (N_12275,N_10606,N_11221);
or U12276 (N_12276,N_10361,N_11749);
nand U12277 (N_12277,N_11288,N_11187);
xnor U12278 (N_12278,N_10729,N_10455);
xnor U12279 (N_12279,N_11304,N_10351);
or U12280 (N_12280,N_11710,N_11539);
nand U12281 (N_12281,N_11060,N_11895);
or U12282 (N_12282,N_11160,N_10064);
xor U12283 (N_12283,N_11624,N_11114);
nor U12284 (N_12284,N_10952,N_10143);
nand U12285 (N_12285,N_11961,N_11836);
nand U12286 (N_12286,N_11914,N_10459);
nand U12287 (N_12287,N_11437,N_10245);
xnor U12288 (N_12288,N_10274,N_10162);
xnor U12289 (N_12289,N_10424,N_11344);
nand U12290 (N_12290,N_11442,N_11666);
xnor U12291 (N_12291,N_10402,N_11412);
nor U12292 (N_12292,N_10019,N_10836);
nor U12293 (N_12293,N_11628,N_10440);
nor U12294 (N_12294,N_11626,N_10004);
nor U12295 (N_12295,N_10570,N_11951);
and U12296 (N_12296,N_11911,N_11434);
nor U12297 (N_12297,N_11066,N_10293);
xnor U12298 (N_12298,N_10733,N_11424);
and U12299 (N_12299,N_11495,N_11169);
nor U12300 (N_12300,N_11562,N_11750);
nor U12301 (N_12301,N_10249,N_11985);
xnor U12302 (N_12302,N_11559,N_10319);
nor U12303 (N_12303,N_11463,N_11557);
nor U12304 (N_12304,N_10785,N_11759);
or U12305 (N_12305,N_11851,N_10828);
xor U12306 (N_12306,N_10708,N_10493);
and U12307 (N_12307,N_10291,N_10972);
and U12308 (N_12308,N_10734,N_11491);
xor U12309 (N_12309,N_10954,N_10145);
xnor U12310 (N_12310,N_11381,N_10384);
nand U12311 (N_12311,N_10585,N_11362);
nand U12312 (N_12312,N_11000,N_11435);
or U12313 (N_12313,N_10703,N_10740);
and U12314 (N_12314,N_10982,N_10797);
xor U12315 (N_12315,N_11245,N_11781);
and U12316 (N_12316,N_10322,N_10821);
and U12317 (N_12317,N_11206,N_11579);
or U12318 (N_12318,N_11935,N_11318);
xnor U12319 (N_12319,N_10168,N_11285);
or U12320 (N_12320,N_11080,N_11932);
nand U12321 (N_12321,N_11820,N_10443);
xor U12322 (N_12322,N_11864,N_11189);
xor U12323 (N_12323,N_10528,N_11922);
and U12324 (N_12324,N_11923,N_11859);
or U12325 (N_12325,N_11838,N_10095);
and U12326 (N_12326,N_10488,N_10248);
or U12327 (N_12327,N_11758,N_10043);
or U12328 (N_12328,N_11185,N_10984);
xnor U12329 (N_12329,N_11552,N_10749);
and U12330 (N_12330,N_11124,N_11320);
nand U12331 (N_12331,N_11128,N_10056);
or U12332 (N_12332,N_11162,N_10702);
and U12333 (N_12333,N_10697,N_10935);
nor U12334 (N_12334,N_11373,N_10496);
or U12335 (N_12335,N_10675,N_11883);
nor U12336 (N_12336,N_11611,N_10414);
xnor U12337 (N_12337,N_10027,N_11191);
nor U12338 (N_12338,N_10367,N_11700);
or U12339 (N_12339,N_10370,N_10858);
or U12340 (N_12340,N_11390,N_10718);
xor U12341 (N_12341,N_11553,N_10857);
xnor U12342 (N_12342,N_11704,N_11081);
or U12343 (N_12343,N_10364,N_11480);
nor U12344 (N_12344,N_10832,N_10382);
xnor U12345 (N_12345,N_10098,N_11846);
nand U12346 (N_12346,N_11481,N_11085);
or U12347 (N_12347,N_10848,N_10612);
nand U12348 (N_12348,N_10525,N_10882);
xor U12349 (N_12349,N_10011,N_11021);
nand U12350 (N_12350,N_10268,N_10616);
xnor U12351 (N_12351,N_11615,N_10758);
and U12352 (N_12352,N_11112,N_11492);
xnor U12353 (N_12353,N_11378,N_11395);
or U12354 (N_12354,N_11002,N_11551);
xnor U12355 (N_12355,N_11925,N_10406);
nand U12356 (N_12356,N_11223,N_10153);
xnor U12357 (N_12357,N_11990,N_11255);
nor U12358 (N_12358,N_10205,N_10588);
xnor U12359 (N_12359,N_11543,N_11649);
and U12360 (N_12360,N_11510,N_11853);
xor U12361 (N_12361,N_11904,N_11029);
nand U12362 (N_12362,N_10615,N_11282);
nor U12363 (N_12363,N_10117,N_10992);
nor U12364 (N_12364,N_11065,N_10754);
nand U12365 (N_12365,N_10039,N_10136);
nand U12366 (N_12366,N_10454,N_11251);
or U12367 (N_12367,N_11891,N_11054);
and U12368 (N_12368,N_11008,N_10129);
and U12369 (N_12369,N_10546,N_11302);
nand U12370 (N_12370,N_10599,N_10505);
or U12371 (N_12371,N_10167,N_11787);
and U12372 (N_12372,N_11377,N_11299);
xnor U12373 (N_12373,N_11897,N_10476);
nand U12374 (N_12374,N_10706,N_11391);
or U12375 (N_12375,N_10763,N_11581);
nand U12376 (N_12376,N_10328,N_10663);
and U12377 (N_12377,N_11894,N_10259);
or U12378 (N_12378,N_11730,N_11308);
and U12379 (N_12379,N_11242,N_11868);
and U12380 (N_12380,N_10358,N_11407);
nor U12381 (N_12381,N_10673,N_10085);
xor U12382 (N_12382,N_10199,N_11878);
or U12383 (N_12383,N_11389,N_10472);
or U12384 (N_12384,N_10562,N_11669);
or U12385 (N_12385,N_10239,N_11680);
xnor U12386 (N_12386,N_10683,N_10667);
nand U12387 (N_12387,N_10150,N_11170);
nor U12388 (N_12388,N_11125,N_10412);
nor U12389 (N_12389,N_11219,N_10078);
nand U12390 (N_12390,N_10352,N_11709);
or U12391 (N_12391,N_10147,N_10499);
and U12392 (N_12392,N_11275,N_10116);
xor U12393 (N_12393,N_11598,N_11295);
nor U12394 (N_12394,N_11336,N_11410);
xnor U12395 (N_12395,N_10042,N_10187);
and U12396 (N_12396,N_11207,N_10976);
xnor U12397 (N_12397,N_11226,N_10803);
nand U12398 (N_12398,N_10800,N_11840);
and U12399 (N_12399,N_11113,N_11560);
and U12400 (N_12400,N_10051,N_11667);
or U12401 (N_12401,N_10583,N_11536);
nor U12402 (N_12402,N_10433,N_11406);
xor U12403 (N_12403,N_10671,N_10784);
nor U12404 (N_12404,N_10354,N_10514);
and U12405 (N_12405,N_11693,N_11341);
nand U12406 (N_12406,N_10462,N_10569);
nand U12407 (N_12407,N_11623,N_11307);
nor U12408 (N_12408,N_11179,N_10679);
xnor U12409 (N_12409,N_10770,N_10790);
and U12410 (N_12410,N_11416,N_11177);
or U12411 (N_12411,N_11131,N_10827);
or U12412 (N_12412,N_10469,N_11351);
or U12413 (N_12413,N_10054,N_10538);
and U12414 (N_12414,N_11142,N_10486);
xor U12415 (N_12415,N_10996,N_10919);
or U12416 (N_12416,N_10655,N_10166);
nand U12417 (N_12417,N_11777,N_11229);
or U12418 (N_12418,N_11879,N_11724);
or U12419 (N_12419,N_10934,N_10927);
and U12420 (N_12420,N_10631,N_10113);
nand U12421 (N_12421,N_10909,N_11791);
nand U12422 (N_12422,N_10066,N_10184);
nor U12423 (N_12423,N_11813,N_11532);
nor U12424 (N_12424,N_10638,N_11067);
xnor U12425 (N_12425,N_11091,N_10951);
or U12426 (N_12426,N_10347,N_11262);
or U12427 (N_12427,N_10346,N_10252);
nor U12428 (N_12428,N_10920,N_11762);
nor U12429 (N_12429,N_11205,N_11590);
nor U12430 (N_12430,N_11645,N_10518);
xor U12431 (N_12431,N_10045,N_11903);
nor U12432 (N_12432,N_11986,N_10387);
xor U12433 (N_12433,N_10152,N_10968);
nand U12434 (N_12434,N_11583,N_10226);
nand U12435 (N_12435,N_11123,N_11631);
or U12436 (N_12436,N_10001,N_10592);
nor U12437 (N_12437,N_10238,N_11356);
nor U12438 (N_12438,N_11303,N_11250);
or U12439 (N_12439,N_10502,N_11477);
or U12440 (N_12440,N_10961,N_11111);
xor U12441 (N_12441,N_10938,N_10281);
nand U12442 (N_12442,N_11259,N_10305);
xor U12443 (N_12443,N_10647,N_11174);
xor U12444 (N_12444,N_11921,N_10416);
xor U12445 (N_12445,N_10487,N_10900);
or U12446 (N_12446,N_10672,N_11143);
and U12447 (N_12447,N_10926,N_10034);
xnor U12448 (N_12448,N_10210,N_10383);
nor U12449 (N_12449,N_11280,N_11423);
nor U12450 (N_12450,N_11073,N_10835);
nand U12451 (N_12451,N_11249,N_10236);
and U12452 (N_12452,N_11361,N_10833);
nand U12453 (N_12453,N_11963,N_10772);
nand U12454 (N_12454,N_10731,N_10280);
or U12455 (N_12455,N_10429,N_10092);
or U12456 (N_12456,N_11465,N_11558);
xnor U12457 (N_12457,N_10312,N_11264);
nor U12458 (N_12458,N_10508,N_10188);
xor U12459 (N_12459,N_10366,N_10313);
or U12460 (N_12460,N_11728,N_11833);
or U12461 (N_12461,N_11063,N_11171);
and U12462 (N_12462,N_11042,N_11872);
or U12463 (N_12463,N_10190,N_11277);
nand U12464 (N_12464,N_10742,N_11794);
nor U12465 (N_12465,N_10460,N_11561);
or U12466 (N_12466,N_11003,N_11366);
nor U12467 (N_12467,N_11654,N_11014);
nand U12468 (N_12468,N_10009,N_10183);
or U12469 (N_12469,N_10320,N_10517);
or U12470 (N_12470,N_10633,N_11182);
and U12471 (N_12471,N_11520,N_10752);
nor U12472 (N_12472,N_11917,N_11156);
nor U12473 (N_12473,N_11947,N_10452);
nor U12474 (N_12474,N_10539,N_11313);
and U12475 (N_12475,N_10450,N_10388);
or U12476 (N_12476,N_11083,N_11753);
xor U12477 (N_12477,N_11471,N_11588);
and U12478 (N_12478,N_10815,N_11906);
and U12479 (N_12479,N_10813,N_10125);
and U12480 (N_12480,N_10956,N_10224);
xor U12481 (N_12481,N_10053,N_10594);
nor U12482 (N_12482,N_10993,N_10192);
and U12483 (N_12483,N_10287,N_10449);
and U12484 (N_12484,N_10256,N_11204);
xor U12485 (N_12485,N_11584,N_11077);
and U12486 (N_12486,N_11852,N_10046);
nand U12487 (N_12487,N_11865,N_11828);
and U12488 (N_12488,N_10596,N_11151);
xnor U12489 (N_12489,N_11033,N_10093);
nand U12490 (N_12490,N_10218,N_11570);
or U12491 (N_12491,N_11337,N_10977);
nor U12492 (N_12492,N_10929,N_11150);
nand U12493 (N_12493,N_11514,N_11665);
nor U12494 (N_12494,N_11524,N_11596);
or U12495 (N_12495,N_11587,N_11574);
nor U12496 (N_12496,N_10315,N_10604);
or U12497 (N_12497,N_11712,N_10945);
xor U12498 (N_12498,N_11022,N_10589);
and U12499 (N_12499,N_11805,N_10971);
xor U12500 (N_12500,N_10251,N_11517);
and U12501 (N_12501,N_10906,N_11966);
nand U12502 (N_12502,N_11769,N_11475);
nor U12503 (N_12503,N_10471,N_10057);
nand U12504 (N_12504,N_10714,N_10850);
xnor U12505 (N_12505,N_10883,N_10365);
nor U12506 (N_12506,N_10942,N_11364);
or U12507 (N_12507,N_10577,N_11254);
and U12508 (N_12508,N_11834,N_10713);
and U12509 (N_12509,N_10127,N_11260);
or U12510 (N_12510,N_11035,N_10304);
and U12511 (N_12511,N_10761,N_10229);
and U12512 (N_12512,N_11147,N_10621);
nand U12513 (N_12513,N_11768,N_11490);
and U12514 (N_12514,N_11097,N_11690);
and U12515 (N_12515,N_10873,N_10881);
and U12516 (N_12516,N_11882,N_11577);
and U12517 (N_12517,N_10531,N_10202);
nor U12518 (N_12518,N_11830,N_11069);
nand U12519 (N_12519,N_10262,N_10944);
and U12520 (N_12520,N_11773,N_11635);
nand U12521 (N_12521,N_11211,N_10903);
xnor U12522 (N_12522,N_11752,N_11352);
and U12523 (N_12523,N_11466,N_10879);
xnor U12524 (N_12524,N_10744,N_10644);
nor U12525 (N_12525,N_11784,N_10323);
xor U12526 (N_12526,N_11698,N_10568);
or U12527 (N_12527,N_11061,N_10751);
and U12528 (N_12528,N_10664,N_10794);
xor U12529 (N_12529,N_11854,N_10485);
nand U12530 (N_12530,N_11230,N_11971);
nor U12531 (N_12531,N_10501,N_11733);
xor U12532 (N_12532,N_11722,N_11683);
and U12533 (N_12533,N_11139,N_10158);
nor U12534 (N_12534,N_10923,N_11421);
xnor U12535 (N_12535,N_10474,N_10483);
nor U12536 (N_12536,N_11359,N_10877);
nand U12537 (N_12537,N_11140,N_11084);
or U12538 (N_12538,N_11610,N_10220);
or U12539 (N_12539,N_10393,N_10185);
or U12540 (N_12540,N_10636,N_11342);
nand U12541 (N_12541,N_11354,N_11374);
nand U12542 (N_12542,N_10888,N_10016);
or U12543 (N_12543,N_10089,N_11326);
or U12544 (N_12544,N_10657,N_11795);
nor U12545 (N_12545,N_10087,N_11236);
or U12546 (N_12546,N_10691,N_11488);
nor U12547 (N_12547,N_11885,N_11630);
nor U12548 (N_12548,N_11203,N_11417);
and U12549 (N_12549,N_11155,N_10593);
or U12550 (N_12550,N_11267,N_11708);
nor U12551 (N_12551,N_10157,N_10824);
nor U12552 (N_12552,N_10289,N_10843);
and U12553 (N_12553,N_10875,N_10055);
nand U12554 (N_12554,N_11887,N_10413);
and U12555 (N_12555,N_10716,N_10632);
xor U12556 (N_12556,N_10975,N_11109);
and U12557 (N_12557,N_11555,N_11565);
or U12558 (N_12558,N_10273,N_11606);
nand U12559 (N_12559,N_11674,N_10526);
or U12560 (N_12560,N_10648,N_11597);
nor U12561 (N_12561,N_10651,N_10542);
nand U12562 (N_12562,N_10932,N_10780);
nand U12563 (N_12563,N_11279,N_10595);
nor U12564 (N_12564,N_11258,N_11898);
or U12565 (N_12565,N_11526,N_10247);
nor U12566 (N_12566,N_11814,N_11821);
or U12567 (N_12567,N_10189,N_10620);
nor U12568 (N_12568,N_10296,N_11335);
nor U12569 (N_12569,N_10897,N_10981);
nor U12570 (N_12570,N_10957,N_10960);
and U12571 (N_12571,N_10895,N_11993);
nand U12572 (N_12572,N_11643,N_10581);
and U12573 (N_12573,N_10867,N_10928);
and U12574 (N_12574,N_11247,N_11782);
or U12575 (N_12575,N_10907,N_10925);
or U12576 (N_12576,N_11968,N_11272);
or U12577 (N_12577,N_10846,N_10149);
nor U12578 (N_12578,N_10561,N_11974);
xor U12579 (N_12579,N_11012,N_11544);
or U12580 (N_12580,N_11433,N_11132);
nor U12581 (N_12581,N_10911,N_10436);
or U12582 (N_12582,N_11827,N_10082);
nand U12583 (N_12583,N_10860,N_10194);
nor U12584 (N_12584,N_10737,N_11050);
and U12585 (N_12585,N_10368,N_10091);
or U12586 (N_12586,N_10856,N_11585);
xnor U12587 (N_12587,N_11376,N_11355);
nor U12588 (N_12588,N_11503,N_10939);
xor U12589 (N_12589,N_10442,N_10257);
xnor U12590 (N_12590,N_10070,N_10573);
or U12591 (N_12591,N_11453,N_11678);
or U12592 (N_12592,N_11281,N_11506);
nor U12593 (N_12593,N_11919,N_10791);
xnor U12594 (N_12594,N_11756,N_11875);
nand U12595 (N_12595,N_11507,N_11322);
and U12596 (N_12596,N_11658,N_11625);
xnor U12597 (N_12597,N_10886,N_10159);
xnor U12598 (N_12598,N_10854,N_11425);
xor U12599 (N_12599,N_10206,N_11199);
or U12600 (N_12600,N_10650,N_11210);
or U12601 (N_12601,N_11744,N_11027);
nand U12602 (N_12602,N_11467,N_11298);
xnor U12603 (N_12603,N_11786,N_11902);
xor U12604 (N_12604,N_10776,N_11673);
nand U12605 (N_12605,N_11982,N_11640);
xor U12606 (N_12606,N_10403,N_11056);
or U12607 (N_12607,N_10349,N_11808);
nand U12608 (N_12608,N_11538,N_10359);
xnor U12609 (N_12609,N_10444,N_10161);
nand U12610 (N_12610,N_10299,N_11920);
nor U12611 (N_12611,N_11909,N_10795);
and U12612 (N_12612,N_11734,N_10659);
or U12613 (N_12613,N_10520,N_11478);
nor U12614 (N_12614,N_10175,N_11642);
and U12615 (N_12615,N_10614,N_10555);
xnor U12616 (N_12616,N_10243,N_11096);
nor U12617 (N_12617,N_11397,N_10209);
xor U12618 (N_12618,N_11420,N_11502);
nand U12619 (N_12619,N_11400,N_10629);
nand U12620 (N_12620,N_10104,N_11367);
xnor U12621 (N_12621,N_11153,N_11004);
or U12622 (N_12622,N_10964,N_10765);
xor U12623 (N_12623,N_11317,N_11212);
or U12624 (N_12624,N_10580,N_11970);
xor U12625 (N_12625,N_11144,N_11508);
and U12626 (N_12626,N_10306,N_11487);
nor U12627 (N_12627,N_10872,N_10492);
xor U12628 (N_12628,N_10980,N_11257);
nor U12629 (N_12629,N_10017,N_10297);
or U12630 (N_12630,N_10456,N_10350);
or U12631 (N_12631,N_10348,N_11745);
and U12632 (N_12632,N_10622,N_10986);
xor U12633 (N_12633,N_10698,N_10603);
or U12634 (N_12634,N_10506,N_10015);
or U12635 (N_12635,N_10468,N_11286);
or U12636 (N_12636,N_11348,N_10038);
nor U12637 (N_12637,N_10653,N_11955);
nand U12638 (N_12638,N_11515,N_10035);
and U12639 (N_12639,N_11567,N_11960);
and U12640 (N_12640,N_11842,N_11240);
and U12641 (N_12641,N_11563,N_11609);
xnor U12642 (N_12642,N_11409,N_11701);
xnor U12643 (N_12643,N_11824,N_11428);
nor U12644 (N_12644,N_10344,N_11271);
nand U12645 (N_12645,N_11194,N_11201);
nor U12646 (N_12646,N_11940,N_10067);
nor U12647 (N_12647,N_10314,N_11694);
nor U12648 (N_12648,N_10578,N_11934);
xor U12649 (N_12649,N_11331,N_10118);
and U12650 (N_12650,N_10548,N_10849);
xor U12651 (N_12651,N_11103,N_11411);
nand U12652 (N_12652,N_11967,N_11607);
xnor U12653 (N_12653,N_10724,N_10894);
nand U12654 (N_12654,N_11736,N_11413);
xnor U12655 (N_12655,N_11957,N_10979);
nand U12656 (N_12656,N_10495,N_11614);
or U12657 (N_12657,N_11456,N_10099);
nor U12658 (N_12658,N_11550,N_11806);
or U12659 (N_12659,N_11408,N_11273);
xor U12660 (N_12660,N_11979,N_10611);
nand U12661 (N_12661,N_10704,N_10507);
nand U12662 (N_12662,N_11659,N_10156);
and U12663 (N_12663,N_10385,N_11266);
nor U12664 (N_12664,N_10178,N_11928);
nand U12665 (N_12665,N_11962,N_11501);
or U12666 (N_12666,N_11239,N_11011);
or U12667 (N_12667,N_10807,N_11725);
and U12668 (N_12668,N_11716,N_11198);
xnor U12669 (N_12669,N_10847,N_10409);
or U12670 (N_12670,N_11330,N_10519);
nand U12671 (N_12671,N_11184,N_11811);
or U12672 (N_12672,N_11403,N_10419);
nor U12673 (N_12673,N_11357,N_10334);
and U12674 (N_12674,N_10014,N_11092);
and U12675 (N_12675,N_10338,N_11432);
xor U12676 (N_12676,N_10669,N_11926);
xnor U12677 (N_12677,N_10181,N_10787);
nand U12678 (N_12678,N_11108,N_11347);
xor U12679 (N_12679,N_10360,N_11419);
and U12680 (N_12680,N_11440,N_11166);
or U12681 (N_12681,N_10103,N_10233);
and U12682 (N_12682,N_11987,N_10998);
or U12683 (N_12683,N_11576,N_11321);
xnor U12684 (N_12684,N_11024,N_11098);
and U12685 (N_12685,N_11118,N_10122);
and U12686 (N_12686,N_10601,N_10260);
and U12687 (N_12687,N_10030,N_10121);
nand U12688 (N_12688,N_11687,N_11195);
and U12689 (N_12689,N_10088,N_10151);
xnor U12690 (N_12690,N_10600,N_10637);
and U12691 (N_12691,N_11387,N_10080);
or U12692 (N_12692,N_11743,N_10031);
and U12693 (N_12693,N_11441,N_11675);
xor U12694 (N_12694,N_11089,N_10710);
and U12695 (N_12695,N_11130,N_10687);
or U12696 (N_12696,N_10084,N_10767);
and U12697 (N_12697,N_10739,N_11964);
xnor U12698 (N_12698,N_10484,N_11637);
or U12699 (N_12699,N_11644,N_11858);
or U12700 (N_12700,N_10608,N_10579);
nand U12701 (N_12701,N_10022,N_10255);
xor U12702 (N_12702,N_11110,N_10686);
nand U12703 (N_12703,N_11668,N_11253);
nand U12704 (N_12704,N_11312,N_10721);
or U12705 (N_12705,N_11988,N_11870);
xor U12706 (N_12706,N_11723,N_10373);
or U12707 (N_12707,N_10172,N_10962);
xnor U12708 (N_12708,N_11158,N_10336);
or U12709 (N_12709,N_11426,N_10941);
nand U12710 (N_12710,N_10831,N_11076);
or U12711 (N_12711,N_11829,N_10902);
nand U12712 (N_12712,N_11863,N_11765);
nor U12713 (N_12713,N_10391,N_10154);
or U12714 (N_12714,N_11608,N_11117);
and U12715 (N_12715,N_10649,N_11006);
and U12716 (N_12716,N_10193,N_11339);
xor U12717 (N_12717,N_10586,N_10574);
and U12718 (N_12718,N_10282,N_10768);
or U12719 (N_12719,N_10868,N_11319);
or U12720 (N_12720,N_10195,N_11040);
and U12721 (N_12721,N_11455,N_11222);
xor U12722 (N_12722,N_11541,N_10173);
nor U12723 (N_12723,N_11910,N_11292);
nand U12724 (N_12724,N_11633,N_10006);
nand U12725 (N_12725,N_10728,N_10511);
or U12726 (N_12726,N_10144,N_10326);
xor U12727 (N_12727,N_10862,N_10623);
or U12728 (N_12728,N_10026,N_11119);
xnor U12729 (N_12729,N_10845,N_11436);
nor U12730 (N_12730,N_10065,N_10963);
nand U12731 (N_12731,N_10617,N_10318);
xor U12732 (N_12732,N_10405,N_11095);
or U12733 (N_12733,N_10590,N_11457);
xnor U12734 (N_12734,N_11843,N_10000);
nor U12735 (N_12735,N_11767,N_11038);
or U12736 (N_12736,N_10689,N_11741);
xnor U12737 (N_12737,N_10386,N_10029);
xnor U12738 (N_12738,N_11525,N_11766);
and U12739 (N_12739,N_10213,N_11566);
xnor U12740 (N_12740,N_11094,N_10102);
xnor U12741 (N_12741,N_10755,N_11748);
xnor U12742 (N_12742,N_10163,N_11731);
xor U12743 (N_12743,N_10111,N_11754);
or U12744 (N_12744,N_11881,N_10778);
nand U12745 (N_12745,N_11998,N_10720);
and U12746 (N_12746,N_10788,N_10007);
nand U12747 (N_12747,N_10421,N_11976);
xnor U12748 (N_12748,N_10946,N_10725);
and U12749 (N_12749,N_11431,N_11306);
and U12750 (N_12750,N_11521,N_10050);
or U12751 (N_12751,N_10880,N_11652);
or U12752 (N_12752,N_11300,N_11540);
or U12753 (N_12753,N_11511,N_11399);
nor U12754 (N_12754,N_10735,N_10186);
xnor U12755 (N_12755,N_11946,N_11942);
or U12756 (N_12756,N_10002,N_11427);
and U12757 (N_12757,N_10227,N_10838);
or U12758 (N_12758,N_10551,N_11656);
xnor U12759 (N_12759,N_10587,N_11209);
or U12760 (N_12760,N_11564,N_11746);
nand U12761 (N_12761,N_10071,N_10931);
xor U12762 (N_12762,N_10753,N_11032);
or U12763 (N_12763,N_11370,N_11790);
xnor U12764 (N_12764,N_11016,N_11679);
nor U12765 (N_12765,N_10047,N_11984);
nand U12766 (N_12766,N_10003,N_10285);
nand U12767 (N_12767,N_10711,N_10090);
or U12768 (N_12768,N_11028,N_11844);
xnor U12769 (N_12769,N_11422,N_11493);
nor U12770 (N_12770,N_11589,N_10464);
and U12771 (N_12771,N_11618,N_11513);
nor U12772 (N_12772,N_11070,N_10676);
and U12773 (N_12773,N_10369,N_11721);
nand U12774 (N_12774,N_11688,N_11036);
and U12775 (N_12775,N_11102,N_10018);
and U12776 (N_12776,N_11079,N_10225);
or U12777 (N_12777,N_11956,N_10969);
nand U12778 (N_12778,N_11931,N_10878);
nand U12779 (N_12779,N_11569,N_10013);
or U12780 (N_12780,N_11542,N_10842);
nand U12781 (N_12781,N_11215,N_11105);
nand U12782 (N_12782,N_10453,N_11135);
xnor U12783 (N_12783,N_10837,N_11992);
or U12784 (N_12784,N_10437,N_11793);
nand U12785 (N_12785,N_11499,N_10852);
or U12786 (N_12786,N_11945,N_11291);
and U12787 (N_12787,N_11009,N_11451);
nor U12788 (N_12788,N_11371,N_11382);
nor U12789 (N_12789,N_10418,N_10481);
nor U12790 (N_12790,N_11816,N_10918);
nor U12791 (N_12791,N_11332,N_10008);
xnor U12792 (N_12792,N_10426,N_10989);
nor U12793 (N_12793,N_10069,N_11718);
and U12794 (N_12794,N_11660,N_10216);
nand U12795 (N_12795,N_11137,N_11861);
nor U12796 (N_12796,N_11418,N_11460);
nor U12797 (N_12797,N_10123,N_10096);
xnor U12798 (N_12798,N_10999,N_10063);
nand U12799 (N_12799,N_11586,N_10910);
nand U12800 (N_12800,N_10988,N_11817);
nand U12801 (N_12801,N_10230,N_10353);
xnor U12802 (N_12802,N_10997,N_10619);
nor U12803 (N_12803,N_10544,N_10853);
or U12804 (N_12804,N_10921,N_11200);
and U12805 (N_12805,N_11638,N_11090);
or U12806 (N_12806,N_11163,N_10130);
nor U12807 (N_12807,N_10760,N_10552);
and U12808 (N_12808,N_10219,N_10682);
nand U12809 (N_12809,N_11430,N_10983);
nand U12810 (N_12810,N_10602,N_11127);
nor U12811 (N_12811,N_11695,N_10816);
xnor U12812 (N_12812,N_10889,N_11706);
nand U12813 (N_12813,N_10124,N_11916);
or U12814 (N_12814,N_11053,N_10549);
or U12815 (N_12815,N_11800,N_11234);
nor U12816 (N_12816,N_10575,N_11547);
nor U12817 (N_12817,N_11005,N_10079);
nand U12818 (N_12818,N_11892,N_11522);
nand U12819 (N_12819,N_10991,N_11358);
or U12820 (N_12820,N_11329,N_10266);
xor U12821 (N_12821,N_11901,N_11629);
and U12822 (N_12822,N_11727,N_11604);
nand U12823 (N_12823,N_11747,N_10913);
or U12824 (N_12824,N_10543,N_10610);
or U12825 (N_12825,N_10135,N_10556);
and U12826 (N_12826,N_10690,N_11048);
xor U12827 (N_12827,N_10396,N_10513);
nor U12828 (N_12828,N_10890,N_11939);
xnor U12829 (N_12829,N_11930,N_10467);
xor U12830 (N_12830,N_11145,N_11739);
nor U12831 (N_12831,N_10498,N_11121);
and U12832 (N_12832,N_11845,N_11058);
nand U12833 (N_12833,N_10717,N_10303);
or U12834 (N_12834,N_10451,N_10940);
and U12835 (N_12835,N_11044,N_11385);
and U12836 (N_12836,N_11620,N_11167);
xor U12837 (N_12837,N_10461,N_10376);
or U12838 (N_12838,N_11533,N_11497);
xor U12839 (N_12839,N_10812,N_11847);
nor U12840 (N_12840,N_10337,N_10512);
nand U12841 (N_12841,N_11208,N_10491);
nor U12842 (N_12842,N_10288,N_11889);
xor U12843 (N_12843,N_10363,N_11068);
and U12844 (N_12844,N_11505,N_11991);
nor U12845 (N_12845,N_10112,N_11839);
xor U12846 (N_12846,N_10044,N_11900);
nand U12847 (N_12847,N_10730,N_11340);
nor U12848 (N_12848,N_11372,N_10861);
or U12849 (N_12849,N_11685,N_10380);
or U12850 (N_12850,N_10696,N_10329);
or U12851 (N_12851,N_11186,N_11572);
or U12852 (N_12852,N_11972,N_10086);
and U12853 (N_12853,N_10719,N_10298);
xnor U12854 (N_12854,N_11995,N_10407);
or U12855 (N_12855,N_10283,N_11055);
or U12856 (N_12856,N_10072,N_11775);
and U12857 (N_12857,N_10738,N_11933);
and U12858 (N_12858,N_10107,N_11857);
and U12859 (N_12859,N_10874,N_11449);
nor U12860 (N_12860,N_10119,N_10893);
nand U12861 (N_12861,N_11580,N_11848);
and U12862 (N_12862,N_10340,N_10871);
nor U12863 (N_12863,N_11173,N_11498);
and U12864 (N_12864,N_10563,N_10830);
or U12865 (N_12865,N_11571,N_11915);
nand U12866 (N_12866,N_11349,N_10263);
nor U12867 (N_12867,N_11328,N_11023);
xor U12868 (N_12868,N_10324,N_10793);
or U12869 (N_12869,N_11296,N_10609);
or U12870 (N_12870,N_10959,N_11146);
nor U12871 (N_12871,N_11938,N_10607);
or U12872 (N_12872,N_11593,N_10036);
or U12873 (N_12873,N_11657,N_10799);
nor U12874 (N_12874,N_11338,N_10823);
nor U12875 (N_12875,N_11443,N_11452);
nand U12876 (N_12876,N_10802,N_10715);
nand U12877 (N_12877,N_11500,N_10097);
and U12878 (N_12878,N_10023,N_10290);
nand U12879 (N_12879,N_10068,N_10427);
or U12880 (N_12880,N_10234,N_10901);
or U12881 (N_12881,N_11227,N_10646);
or U12882 (N_12882,N_11907,N_11287);
nor U12883 (N_12883,N_10550,N_11602);
or U12884 (N_12884,N_11473,N_11689);
or U12885 (N_12885,N_10377,N_10480);
and U12886 (N_12886,N_11763,N_10024);
and U12887 (N_12887,N_10908,N_11224);
xor U12888 (N_12888,N_11944,N_11030);
and U12889 (N_12889,N_10335,N_11835);
nand U12890 (N_12890,N_11713,N_10463);
and U12891 (N_12891,N_10553,N_11476);
or U12892 (N_12892,N_10279,N_11568);
nand U12893 (N_12893,N_10275,N_11485);
or U12894 (N_12894,N_11246,N_10231);
and U12895 (N_12895,N_11256,N_10278);
nand U12896 (N_12896,N_11360,N_11034);
xor U12897 (N_12897,N_11334,N_10769);
or U12898 (N_12898,N_11707,N_11989);
or U12899 (N_12899,N_11365,N_11908);
xor U12900 (N_12900,N_10567,N_10937);
nor U12901 (N_12901,N_11197,N_11818);
or U12902 (N_12902,N_11157,N_10571);
xor U12903 (N_12903,N_11013,N_11691);
nand U12904 (N_12904,N_10955,N_10074);
xnor U12905 (N_12905,N_10253,N_10465);
nand U12906 (N_12906,N_11238,N_10576);
or U12907 (N_12907,N_11353,N_10870);
or U12908 (N_12908,N_10819,N_11134);
or U12909 (N_12909,N_10164,N_10625);
nand U12910 (N_12910,N_11639,N_10286);
xor U12911 (N_12911,N_11913,N_10965);
xor U12912 (N_12912,N_10410,N_11181);
nor U12913 (N_12913,N_10497,N_10885);
nor U12914 (N_12914,N_10325,N_10917);
nor U12915 (N_12915,N_10431,N_10394);
and U12916 (N_12916,N_11632,N_10301);
nand U12917 (N_12917,N_11176,N_10564);
nand U12918 (N_12918,N_10530,N_10582);
nor U12919 (N_12919,N_11388,N_10342);
and U12920 (N_12920,N_10990,N_10529);
nor U12921 (N_12921,N_10100,N_11444);
and U12922 (N_12922,N_10179,N_10343);
and U12923 (N_12923,N_11874,N_10914);
xnor U12924 (N_12924,N_11175,N_10692);
nand U12925 (N_12925,N_10048,N_10947);
nand U12926 (N_12926,N_11392,N_11104);
nand U12927 (N_12927,N_10345,N_11244);
nor U12928 (N_12928,N_10398,N_10395);
xnor U12929 (N_12929,N_10198,N_11809);
or U12930 (N_12930,N_11059,N_10447);
or U12931 (N_12931,N_10789,N_10240);
nor U12932 (N_12932,N_11825,N_11890);
xnor U12933 (N_12933,N_10221,N_10810);
nor U12934 (N_12934,N_10782,N_10375);
or U12935 (N_12935,N_10148,N_10806);
or U12936 (N_12936,N_10510,N_10726);
and U12937 (N_12937,N_11534,N_11975);
nor U12938 (N_12938,N_11241,N_10743);
xor U12939 (N_12939,N_10200,N_10432);
xor U12940 (N_12940,N_10665,N_11856);
nor U12941 (N_12941,N_11323,N_11489);
xor U12942 (N_12942,N_10727,N_11026);
nand U12943 (N_12943,N_11981,N_11325);
and U12944 (N_12944,N_10966,N_11010);
and U12945 (N_12945,N_11213,N_10922);
or U12946 (N_12946,N_11115,N_11218);
nand U12947 (N_12947,N_11086,N_10201);
nor U12948 (N_12948,N_11612,N_10685);
xnor U12949 (N_12949,N_11980,N_11152);
and U12950 (N_12950,N_11801,N_11398);
nor U12951 (N_12951,N_11049,N_11217);
nor U12952 (N_12952,N_10308,N_11591);
or U12953 (N_12953,N_10141,N_11929);
nor U12954 (N_12954,N_11017,N_10399);
and U12955 (N_12955,N_11776,N_10707);
and U12956 (N_12956,N_11831,N_11996);
nand U12957 (N_12957,N_11714,N_11116);
or U12958 (N_12958,N_11941,N_11605);
nor U12959 (N_12959,N_10128,N_10142);
nor U12960 (N_12960,N_10114,N_11617);
or U12961 (N_12961,N_10747,N_11232);
nand U12962 (N_12962,N_11415,N_10841);
or U12963 (N_12963,N_10106,N_11345);
xnor U12964 (N_12964,N_10958,N_10677);
and U12965 (N_12965,N_11180,N_11379);
xnor U12966 (N_12966,N_11057,N_11886);
or U12967 (N_12967,N_11052,N_10899);
nand U12968 (N_12968,N_10598,N_10866);
nand U12969 (N_12969,N_10930,N_10916);
xor U12970 (N_12970,N_10987,N_10060);
nand U12971 (N_12971,N_11284,N_10302);
nand U12972 (N_12972,N_11454,N_10973);
nor U12973 (N_12973,N_10331,N_11309);
and U12974 (N_12974,N_11472,N_11600);
nor U12975 (N_12975,N_11459,N_10212);
xnor U12976 (N_12976,N_10764,N_10948);
xor U12977 (N_12977,N_11243,N_10804);
and U12978 (N_12978,N_11216,N_11078);
and U12979 (N_12979,N_10473,N_11778);
xor U12980 (N_12980,N_11719,N_10235);
nor U12981 (N_12981,N_11343,N_10371);
or U12982 (N_12982,N_10950,N_10978);
nand U12983 (N_12983,N_10701,N_11671);
and U12984 (N_12984,N_10798,N_11470);
or U12985 (N_12985,N_10330,N_11912);
or U12986 (N_12986,N_11812,N_10110);
nand U12987 (N_12987,N_11664,N_11893);
nor U12988 (N_12988,N_11973,N_11641);
nor U12989 (N_12989,N_10228,N_11458);
nand U12990 (N_12990,N_11943,N_11314);
and U12991 (N_12991,N_10732,N_11850);
or U12992 (N_12992,N_10521,N_11696);
nand U12993 (N_12993,N_10662,N_10466);
or U12994 (N_12994,N_10126,N_10232);
and U12995 (N_12995,N_11064,N_11697);
or U12996 (N_12996,N_10558,N_11720);
nor U12997 (N_12997,N_11138,N_10207);
nor U12998 (N_12998,N_10635,N_10545);
and U12999 (N_12999,N_11363,N_10801);
or U13000 (N_13000,N_10986,N_11562);
nand U13001 (N_13001,N_11124,N_10394);
xor U13002 (N_13002,N_10050,N_11425);
nand U13003 (N_13003,N_11036,N_11789);
or U13004 (N_13004,N_10332,N_11978);
xnor U13005 (N_13005,N_11998,N_10641);
and U13006 (N_13006,N_10749,N_10381);
nand U13007 (N_13007,N_10491,N_10195);
and U13008 (N_13008,N_10885,N_10992);
nor U13009 (N_13009,N_10785,N_11975);
nand U13010 (N_13010,N_10178,N_10411);
and U13011 (N_13011,N_11968,N_11632);
or U13012 (N_13012,N_11127,N_11796);
or U13013 (N_13013,N_11733,N_10935);
or U13014 (N_13014,N_10869,N_11689);
and U13015 (N_13015,N_11976,N_11746);
nor U13016 (N_13016,N_11382,N_11773);
xnor U13017 (N_13017,N_11128,N_10515);
nand U13018 (N_13018,N_11355,N_10366);
or U13019 (N_13019,N_11683,N_11569);
nor U13020 (N_13020,N_11054,N_11162);
nand U13021 (N_13021,N_11861,N_11826);
or U13022 (N_13022,N_10991,N_11112);
or U13023 (N_13023,N_11636,N_10211);
xnor U13024 (N_13024,N_11012,N_11642);
or U13025 (N_13025,N_11262,N_11243);
or U13026 (N_13026,N_10714,N_10343);
nand U13027 (N_13027,N_11341,N_10634);
or U13028 (N_13028,N_11822,N_10291);
and U13029 (N_13029,N_10554,N_11933);
nand U13030 (N_13030,N_11886,N_10895);
xnor U13031 (N_13031,N_11749,N_11204);
and U13032 (N_13032,N_10048,N_11388);
xor U13033 (N_13033,N_10930,N_10064);
and U13034 (N_13034,N_11804,N_10856);
nand U13035 (N_13035,N_10957,N_10666);
xnor U13036 (N_13036,N_11826,N_10639);
nor U13037 (N_13037,N_10296,N_10421);
and U13038 (N_13038,N_11098,N_11732);
or U13039 (N_13039,N_10523,N_10598);
xnor U13040 (N_13040,N_10387,N_11795);
nand U13041 (N_13041,N_10814,N_11511);
or U13042 (N_13042,N_10376,N_11394);
xnor U13043 (N_13043,N_11422,N_10044);
xnor U13044 (N_13044,N_10681,N_11588);
and U13045 (N_13045,N_10458,N_10417);
or U13046 (N_13046,N_10104,N_10200);
and U13047 (N_13047,N_10063,N_10422);
nand U13048 (N_13048,N_10303,N_11626);
nand U13049 (N_13049,N_10361,N_10842);
and U13050 (N_13050,N_11680,N_10312);
nor U13051 (N_13051,N_11892,N_11470);
and U13052 (N_13052,N_10539,N_11358);
nand U13053 (N_13053,N_11343,N_10786);
nand U13054 (N_13054,N_10985,N_10503);
nand U13055 (N_13055,N_10835,N_11286);
and U13056 (N_13056,N_11609,N_10290);
nor U13057 (N_13057,N_10729,N_11752);
nand U13058 (N_13058,N_10089,N_11566);
and U13059 (N_13059,N_11036,N_11259);
nand U13060 (N_13060,N_11792,N_10651);
nand U13061 (N_13061,N_10131,N_11101);
nand U13062 (N_13062,N_10761,N_11019);
nand U13063 (N_13063,N_10392,N_10566);
and U13064 (N_13064,N_10482,N_11980);
nor U13065 (N_13065,N_11400,N_11127);
xor U13066 (N_13066,N_11604,N_10687);
and U13067 (N_13067,N_10181,N_10990);
and U13068 (N_13068,N_11682,N_10441);
xnor U13069 (N_13069,N_10107,N_11139);
xnor U13070 (N_13070,N_10480,N_10774);
nor U13071 (N_13071,N_11492,N_10258);
nor U13072 (N_13072,N_10907,N_10800);
nor U13073 (N_13073,N_10973,N_11316);
and U13074 (N_13074,N_10896,N_10219);
xor U13075 (N_13075,N_11180,N_11325);
nand U13076 (N_13076,N_11614,N_10284);
nor U13077 (N_13077,N_10069,N_11432);
and U13078 (N_13078,N_11102,N_11363);
or U13079 (N_13079,N_11305,N_10685);
nand U13080 (N_13080,N_10956,N_10355);
or U13081 (N_13081,N_10940,N_10738);
xor U13082 (N_13082,N_10438,N_10646);
or U13083 (N_13083,N_11345,N_10517);
nor U13084 (N_13084,N_11047,N_10151);
and U13085 (N_13085,N_11187,N_10670);
xor U13086 (N_13086,N_10027,N_11832);
nand U13087 (N_13087,N_10070,N_11671);
nand U13088 (N_13088,N_10166,N_11698);
xor U13089 (N_13089,N_10874,N_10415);
xor U13090 (N_13090,N_11554,N_11573);
nand U13091 (N_13091,N_11782,N_11801);
nor U13092 (N_13092,N_11035,N_11765);
or U13093 (N_13093,N_10507,N_11414);
or U13094 (N_13094,N_11513,N_11205);
nor U13095 (N_13095,N_11909,N_10863);
and U13096 (N_13096,N_10424,N_11622);
or U13097 (N_13097,N_11785,N_11331);
or U13098 (N_13098,N_11283,N_11108);
xnor U13099 (N_13099,N_11288,N_10910);
or U13100 (N_13100,N_11938,N_10648);
xnor U13101 (N_13101,N_11085,N_11934);
or U13102 (N_13102,N_10964,N_11314);
nor U13103 (N_13103,N_11715,N_11408);
nor U13104 (N_13104,N_11455,N_11246);
or U13105 (N_13105,N_11151,N_10225);
xnor U13106 (N_13106,N_11203,N_10729);
xor U13107 (N_13107,N_11364,N_11727);
nor U13108 (N_13108,N_10543,N_11560);
nand U13109 (N_13109,N_10575,N_11158);
and U13110 (N_13110,N_11483,N_11125);
xor U13111 (N_13111,N_11542,N_11577);
nand U13112 (N_13112,N_11360,N_10989);
nor U13113 (N_13113,N_10825,N_11156);
nor U13114 (N_13114,N_10664,N_10295);
xnor U13115 (N_13115,N_10010,N_11669);
and U13116 (N_13116,N_10884,N_10110);
or U13117 (N_13117,N_11683,N_11296);
and U13118 (N_13118,N_11469,N_10992);
and U13119 (N_13119,N_10127,N_11486);
or U13120 (N_13120,N_10386,N_10211);
xnor U13121 (N_13121,N_11730,N_11575);
or U13122 (N_13122,N_11552,N_10232);
and U13123 (N_13123,N_11187,N_10609);
and U13124 (N_13124,N_11579,N_11199);
and U13125 (N_13125,N_11902,N_11269);
and U13126 (N_13126,N_11039,N_10767);
or U13127 (N_13127,N_11604,N_11414);
and U13128 (N_13128,N_10824,N_10773);
nand U13129 (N_13129,N_11630,N_10122);
xnor U13130 (N_13130,N_11511,N_10060);
nor U13131 (N_13131,N_10722,N_10083);
and U13132 (N_13132,N_11257,N_10932);
xor U13133 (N_13133,N_10546,N_11439);
and U13134 (N_13134,N_10993,N_10350);
xnor U13135 (N_13135,N_10591,N_11003);
or U13136 (N_13136,N_11787,N_11385);
and U13137 (N_13137,N_10219,N_10370);
or U13138 (N_13138,N_11293,N_10501);
and U13139 (N_13139,N_10839,N_10521);
nand U13140 (N_13140,N_10016,N_11057);
nor U13141 (N_13141,N_10043,N_11506);
xnor U13142 (N_13142,N_11311,N_11051);
nor U13143 (N_13143,N_10187,N_10808);
or U13144 (N_13144,N_10915,N_10182);
nand U13145 (N_13145,N_10047,N_10738);
or U13146 (N_13146,N_10327,N_10887);
and U13147 (N_13147,N_11411,N_10975);
nor U13148 (N_13148,N_10056,N_10534);
or U13149 (N_13149,N_11412,N_10585);
or U13150 (N_13150,N_10088,N_11254);
or U13151 (N_13151,N_10878,N_10927);
or U13152 (N_13152,N_10362,N_11272);
or U13153 (N_13153,N_11322,N_10930);
nand U13154 (N_13154,N_10256,N_10349);
and U13155 (N_13155,N_11678,N_11051);
and U13156 (N_13156,N_10230,N_10041);
and U13157 (N_13157,N_10004,N_11568);
xor U13158 (N_13158,N_10355,N_11663);
nor U13159 (N_13159,N_10374,N_10840);
and U13160 (N_13160,N_10487,N_10250);
xor U13161 (N_13161,N_11460,N_11294);
xor U13162 (N_13162,N_11503,N_10768);
nor U13163 (N_13163,N_10486,N_10982);
nor U13164 (N_13164,N_11742,N_10092);
or U13165 (N_13165,N_10433,N_11500);
or U13166 (N_13166,N_10693,N_11580);
nor U13167 (N_13167,N_11391,N_10899);
nand U13168 (N_13168,N_10639,N_11122);
xnor U13169 (N_13169,N_11446,N_10533);
or U13170 (N_13170,N_10951,N_11271);
nand U13171 (N_13171,N_11328,N_11797);
nand U13172 (N_13172,N_11722,N_11007);
xor U13173 (N_13173,N_10462,N_11983);
and U13174 (N_13174,N_11618,N_10437);
nand U13175 (N_13175,N_11223,N_10480);
and U13176 (N_13176,N_10828,N_10145);
and U13177 (N_13177,N_11362,N_10848);
nor U13178 (N_13178,N_10736,N_10020);
xor U13179 (N_13179,N_11174,N_11173);
nor U13180 (N_13180,N_10594,N_11974);
or U13181 (N_13181,N_11318,N_11710);
or U13182 (N_13182,N_11424,N_10022);
xor U13183 (N_13183,N_10694,N_10116);
or U13184 (N_13184,N_10183,N_11218);
or U13185 (N_13185,N_11822,N_11306);
nor U13186 (N_13186,N_11374,N_10036);
xor U13187 (N_13187,N_10344,N_10915);
and U13188 (N_13188,N_11215,N_11493);
nor U13189 (N_13189,N_11319,N_11983);
and U13190 (N_13190,N_11770,N_10935);
xnor U13191 (N_13191,N_11732,N_10767);
nor U13192 (N_13192,N_10070,N_11522);
and U13193 (N_13193,N_11040,N_11228);
nor U13194 (N_13194,N_10561,N_11014);
nor U13195 (N_13195,N_11390,N_11272);
nand U13196 (N_13196,N_11003,N_11761);
nor U13197 (N_13197,N_11735,N_10766);
nand U13198 (N_13198,N_10190,N_10154);
nor U13199 (N_13199,N_10379,N_10206);
nor U13200 (N_13200,N_11557,N_11151);
or U13201 (N_13201,N_11800,N_11480);
nand U13202 (N_13202,N_10062,N_10079);
nand U13203 (N_13203,N_10778,N_11777);
and U13204 (N_13204,N_11012,N_10884);
or U13205 (N_13205,N_10312,N_10000);
or U13206 (N_13206,N_11214,N_11053);
xor U13207 (N_13207,N_11802,N_11129);
nand U13208 (N_13208,N_10600,N_10074);
nand U13209 (N_13209,N_11714,N_11419);
and U13210 (N_13210,N_10397,N_10542);
nor U13211 (N_13211,N_10063,N_10770);
and U13212 (N_13212,N_10242,N_11297);
xnor U13213 (N_13213,N_11654,N_10625);
or U13214 (N_13214,N_10545,N_10622);
or U13215 (N_13215,N_10002,N_11568);
or U13216 (N_13216,N_10665,N_11508);
nor U13217 (N_13217,N_10648,N_10454);
nand U13218 (N_13218,N_10825,N_11992);
xor U13219 (N_13219,N_10628,N_11825);
and U13220 (N_13220,N_10911,N_10635);
or U13221 (N_13221,N_11853,N_10296);
nand U13222 (N_13222,N_10377,N_10444);
and U13223 (N_13223,N_11958,N_11897);
or U13224 (N_13224,N_10372,N_10700);
nor U13225 (N_13225,N_11016,N_11119);
nand U13226 (N_13226,N_10069,N_10563);
xnor U13227 (N_13227,N_10367,N_10441);
or U13228 (N_13228,N_11183,N_10827);
xnor U13229 (N_13229,N_10541,N_10959);
nand U13230 (N_13230,N_11911,N_10836);
nor U13231 (N_13231,N_10609,N_10263);
xnor U13232 (N_13232,N_11734,N_10657);
and U13233 (N_13233,N_10625,N_10867);
nand U13234 (N_13234,N_11326,N_10240);
or U13235 (N_13235,N_11179,N_10576);
nor U13236 (N_13236,N_10953,N_10619);
nand U13237 (N_13237,N_11861,N_11480);
or U13238 (N_13238,N_10399,N_10991);
or U13239 (N_13239,N_11986,N_11233);
or U13240 (N_13240,N_11499,N_11971);
nand U13241 (N_13241,N_10533,N_10258);
xnor U13242 (N_13242,N_10462,N_10916);
nor U13243 (N_13243,N_10317,N_11021);
and U13244 (N_13244,N_10127,N_11977);
and U13245 (N_13245,N_11469,N_10042);
nor U13246 (N_13246,N_10800,N_10654);
or U13247 (N_13247,N_10947,N_10893);
nand U13248 (N_13248,N_10560,N_10899);
or U13249 (N_13249,N_10341,N_10820);
nand U13250 (N_13250,N_11235,N_10720);
nand U13251 (N_13251,N_11394,N_11104);
xnor U13252 (N_13252,N_11640,N_11291);
xnor U13253 (N_13253,N_10840,N_10386);
or U13254 (N_13254,N_11955,N_10781);
and U13255 (N_13255,N_10619,N_10225);
or U13256 (N_13256,N_10513,N_11699);
xnor U13257 (N_13257,N_10643,N_11342);
xnor U13258 (N_13258,N_10028,N_11410);
nor U13259 (N_13259,N_10960,N_11176);
and U13260 (N_13260,N_10764,N_11687);
nand U13261 (N_13261,N_10130,N_11538);
nand U13262 (N_13262,N_10342,N_11367);
xnor U13263 (N_13263,N_10768,N_10239);
and U13264 (N_13264,N_10155,N_11997);
xnor U13265 (N_13265,N_11657,N_11078);
nor U13266 (N_13266,N_10816,N_10058);
or U13267 (N_13267,N_10927,N_10602);
xnor U13268 (N_13268,N_11165,N_10106);
nor U13269 (N_13269,N_11980,N_10213);
xor U13270 (N_13270,N_10565,N_11978);
xor U13271 (N_13271,N_10954,N_11102);
nand U13272 (N_13272,N_11200,N_11985);
or U13273 (N_13273,N_11672,N_10590);
nand U13274 (N_13274,N_11444,N_11624);
and U13275 (N_13275,N_11799,N_10911);
and U13276 (N_13276,N_11068,N_11844);
and U13277 (N_13277,N_10426,N_11846);
or U13278 (N_13278,N_11886,N_10317);
and U13279 (N_13279,N_11523,N_11631);
or U13280 (N_13280,N_10486,N_11178);
xor U13281 (N_13281,N_10196,N_10930);
or U13282 (N_13282,N_11237,N_11665);
nand U13283 (N_13283,N_11769,N_11400);
xor U13284 (N_13284,N_10470,N_11410);
and U13285 (N_13285,N_11699,N_11209);
nand U13286 (N_13286,N_10686,N_10974);
and U13287 (N_13287,N_10554,N_11758);
nand U13288 (N_13288,N_10854,N_11206);
nand U13289 (N_13289,N_10241,N_10294);
nand U13290 (N_13290,N_10227,N_10755);
and U13291 (N_13291,N_10717,N_11144);
xor U13292 (N_13292,N_11193,N_11140);
xor U13293 (N_13293,N_11824,N_11054);
xor U13294 (N_13294,N_11825,N_11899);
or U13295 (N_13295,N_11522,N_11836);
and U13296 (N_13296,N_11716,N_11496);
and U13297 (N_13297,N_11649,N_11346);
nor U13298 (N_13298,N_10141,N_10206);
or U13299 (N_13299,N_11720,N_10960);
nand U13300 (N_13300,N_10462,N_10029);
nand U13301 (N_13301,N_10562,N_11135);
and U13302 (N_13302,N_11518,N_11741);
or U13303 (N_13303,N_10565,N_10230);
or U13304 (N_13304,N_10986,N_10491);
or U13305 (N_13305,N_11862,N_11728);
and U13306 (N_13306,N_10565,N_11946);
nor U13307 (N_13307,N_10860,N_10102);
nor U13308 (N_13308,N_10408,N_10048);
or U13309 (N_13309,N_11840,N_11706);
nor U13310 (N_13310,N_10185,N_10325);
nor U13311 (N_13311,N_10175,N_10000);
nor U13312 (N_13312,N_10519,N_11936);
nor U13313 (N_13313,N_11815,N_10038);
nand U13314 (N_13314,N_11290,N_11693);
nand U13315 (N_13315,N_10958,N_10194);
and U13316 (N_13316,N_11272,N_10124);
or U13317 (N_13317,N_10337,N_11550);
or U13318 (N_13318,N_10046,N_11568);
nand U13319 (N_13319,N_11907,N_11025);
xor U13320 (N_13320,N_11261,N_10847);
and U13321 (N_13321,N_10423,N_10687);
xnor U13322 (N_13322,N_11199,N_10986);
xor U13323 (N_13323,N_10594,N_10476);
and U13324 (N_13324,N_11917,N_10316);
and U13325 (N_13325,N_10692,N_10706);
nand U13326 (N_13326,N_11898,N_10409);
xnor U13327 (N_13327,N_10066,N_11706);
xnor U13328 (N_13328,N_11081,N_10299);
nand U13329 (N_13329,N_11679,N_10039);
nand U13330 (N_13330,N_10527,N_10128);
xor U13331 (N_13331,N_11468,N_10960);
nor U13332 (N_13332,N_10304,N_11849);
nand U13333 (N_13333,N_10074,N_10107);
and U13334 (N_13334,N_10203,N_10586);
or U13335 (N_13335,N_11200,N_11962);
nand U13336 (N_13336,N_10473,N_10062);
nand U13337 (N_13337,N_10216,N_11558);
nand U13338 (N_13338,N_10216,N_11419);
xnor U13339 (N_13339,N_10514,N_11813);
or U13340 (N_13340,N_11264,N_10288);
xnor U13341 (N_13341,N_10891,N_10616);
nand U13342 (N_13342,N_10246,N_11237);
nand U13343 (N_13343,N_10504,N_10943);
nand U13344 (N_13344,N_10048,N_10171);
nand U13345 (N_13345,N_10774,N_10117);
or U13346 (N_13346,N_11291,N_10491);
and U13347 (N_13347,N_10843,N_10533);
xnor U13348 (N_13348,N_10338,N_11254);
nor U13349 (N_13349,N_11428,N_10419);
nand U13350 (N_13350,N_10701,N_10358);
nor U13351 (N_13351,N_11859,N_10629);
xor U13352 (N_13352,N_10251,N_11871);
xnor U13353 (N_13353,N_10032,N_10133);
nor U13354 (N_13354,N_11739,N_11843);
or U13355 (N_13355,N_10761,N_10427);
xnor U13356 (N_13356,N_10328,N_11557);
nor U13357 (N_13357,N_10489,N_11423);
or U13358 (N_13358,N_11619,N_11622);
xnor U13359 (N_13359,N_11651,N_11875);
and U13360 (N_13360,N_10636,N_10065);
nor U13361 (N_13361,N_11251,N_11438);
or U13362 (N_13362,N_11771,N_10420);
xnor U13363 (N_13363,N_10676,N_10205);
nor U13364 (N_13364,N_10951,N_10126);
nand U13365 (N_13365,N_11495,N_11625);
nand U13366 (N_13366,N_10660,N_11791);
nand U13367 (N_13367,N_11760,N_10282);
nor U13368 (N_13368,N_11241,N_10312);
xor U13369 (N_13369,N_11407,N_11841);
and U13370 (N_13370,N_11044,N_10770);
xor U13371 (N_13371,N_10265,N_11936);
nand U13372 (N_13372,N_10769,N_11227);
nand U13373 (N_13373,N_10208,N_11668);
or U13374 (N_13374,N_11828,N_11111);
nor U13375 (N_13375,N_10622,N_11296);
nor U13376 (N_13376,N_10805,N_10432);
nor U13377 (N_13377,N_11065,N_11548);
nor U13378 (N_13378,N_11581,N_10206);
xnor U13379 (N_13379,N_11563,N_10439);
nor U13380 (N_13380,N_11562,N_11576);
nor U13381 (N_13381,N_11903,N_11083);
xor U13382 (N_13382,N_11197,N_11815);
nor U13383 (N_13383,N_10712,N_10818);
nand U13384 (N_13384,N_11347,N_10578);
nor U13385 (N_13385,N_10629,N_11488);
nand U13386 (N_13386,N_11454,N_10695);
and U13387 (N_13387,N_11098,N_11467);
nor U13388 (N_13388,N_11264,N_10701);
or U13389 (N_13389,N_10792,N_11401);
nor U13390 (N_13390,N_10881,N_11851);
or U13391 (N_13391,N_11327,N_10610);
nor U13392 (N_13392,N_11367,N_10719);
xor U13393 (N_13393,N_11563,N_11851);
or U13394 (N_13394,N_11064,N_11425);
and U13395 (N_13395,N_11793,N_10855);
xor U13396 (N_13396,N_10794,N_11888);
xor U13397 (N_13397,N_10679,N_10657);
nor U13398 (N_13398,N_10888,N_10098);
nand U13399 (N_13399,N_11720,N_10842);
nor U13400 (N_13400,N_11543,N_11224);
or U13401 (N_13401,N_11546,N_11912);
nand U13402 (N_13402,N_11594,N_11595);
nand U13403 (N_13403,N_10178,N_11630);
and U13404 (N_13404,N_11092,N_10661);
nand U13405 (N_13405,N_11529,N_10269);
nand U13406 (N_13406,N_10842,N_10990);
xor U13407 (N_13407,N_11838,N_10143);
nor U13408 (N_13408,N_11145,N_11502);
nand U13409 (N_13409,N_11782,N_10260);
and U13410 (N_13410,N_10642,N_11027);
xnor U13411 (N_13411,N_10415,N_10504);
xor U13412 (N_13412,N_11161,N_11417);
or U13413 (N_13413,N_11118,N_10407);
or U13414 (N_13414,N_11510,N_10577);
xor U13415 (N_13415,N_11423,N_11061);
or U13416 (N_13416,N_11696,N_11525);
or U13417 (N_13417,N_10203,N_11832);
nor U13418 (N_13418,N_10749,N_11805);
xnor U13419 (N_13419,N_10111,N_10195);
or U13420 (N_13420,N_10882,N_11926);
xnor U13421 (N_13421,N_10532,N_11367);
or U13422 (N_13422,N_10317,N_10070);
nand U13423 (N_13423,N_11277,N_11024);
xnor U13424 (N_13424,N_10750,N_11726);
nand U13425 (N_13425,N_11008,N_10955);
nor U13426 (N_13426,N_10253,N_10122);
xor U13427 (N_13427,N_10928,N_10208);
and U13428 (N_13428,N_10634,N_11363);
or U13429 (N_13429,N_11729,N_11871);
and U13430 (N_13430,N_11872,N_10016);
nor U13431 (N_13431,N_10560,N_10430);
nand U13432 (N_13432,N_10617,N_10019);
and U13433 (N_13433,N_10447,N_10101);
and U13434 (N_13434,N_11189,N_11580);
or U13435 (N_13435,N_11032,N_11514);
xnor U13436 (N_13436,N_11307,N_11539);
xor U13437 (N_13437,N_11067,N_11987);
nor U13438 (N_13438,N_10143,N_10867);
nand U13439 (N_13439,N_11795,N_10831);
xnor U13440 (N_13440,N_10125,N_11426);
xnor U13441 (N_13441,N_11114,N_10678);
or U13442 (N_13442,N_10003,N_11207);
and U13443 (N_13443,N_11449,N_10560);
nand U13444 (N_13444,N_11335,N_11580);
nand U13445 (N_13445,N_10943,N_11262);
and U13446 (N_13446,N_11777,N_11096);
xor U13447 (N_13447,N_10800,N_11225);
or U13448 (N_13448,N_10381,N_11234);
or U13449 (N_13449,N_10804,N_10263);
nor U13450 (N_13450,N_10181,N_11915);
nor U13451 (N_13451,N_10783,N_11023);
or U13452 (N_13452,N_11893,N_10402);
nand U13453 (N_13453,N_10579,N_11067);
and U13454 (N_13454,N_10520,N_10921);
xnor U13455 (N_13455,N_10478,N_11057);
nand U13456 (N_13456,N_11923,N_11703);
xor U13457 (N_13457,N_11052,N_10798);
nand U13458 (N_13458,N_11713,N_11474);
or U13459 (N_13459,N_11703,N_10422);
nor U13460 (N_13460,N_11165,N_10094);
or U13461 (N_13461,N_11064,N_11658);
or U13462 (N_13462,N_11116,N_11260);
or U13463 (N_13463,N_10445,N_10458);
and U13464 (N_13464,N_10144,N_10275);
nor U13465 (N_13465,N_11168,N_11000);
or U13466 (N_13466,N_11795,N_10761);
nor U13467 (N_13467,N_11538,N_11261);
nand U13468 (N_13468,N_11796,N_11211);
and U13469 (N_13469,N_11661,N_11403);
nor U13470 (N_13470,N_10774,N_11967);
nor U13471 (N_13471,N_10484,N_10504);
xor U13472 (N_13472,N_10027,N_11460);
and U13473 (N_13473,N_11960,N_10443);
nand U13474 (N_13474,N_11546,N_11542);
nand U13475 (N_13475,N_10371,N_10243);
and U13476 (N_13476,N_11886,N_10160);
xnor U13477 (N_13477,N_10109,N_10451);
xor U13478 (N_13478,N_10086,N_10668);
nand U13479 (N_13479,N_10938,N_11375);
xnor U13480 (N_13480,N_11334,N_11372);
xor U13481 (N_13481,N_11628,N_10009);
nor U13482 (N_13482,N_11486,N_10041);
nor U13483 (N_13483,N_11185,N_10029);
and U13484 (N_13484,N_11400,N_10903);
or U13485 (N_13485,N_10624,N_11413);
xor U13486 (N_13486,N_11026,N_10959);
xnor U13487 (N_13487,N_10848,N_11114);
nand U13488 (N_13488,N_11797,N_10470);
nand U13489 (N_13489,N_11610,N_10963);
nand U13490 (N_13490,N_11203,N_11550);
nand U13491 (N_13491,N_10229,N_10567);
nand U13492 (N_13492,N_10844,N_11626);
nand U13493 (N_13493,N_10993,N_11435);
nand U13494 (N_13494,N_10728,N_11940);
nand U13495 (N_13495,N_10254,N_11010);
xor U13496 (N_13496,N_10343,N_10166);
xor U13497 (N_13497,N_10945,N_10535);
or U13498 (N_13498,N_11772,N_10607);
or U13499 (N_13499,N_10182,N_10918);
xnor U13500 (N_13500,N_11310,N_11980);
xnor U13501 (N_13501,N_10790,N_10587);
xor U13502 (N_13502,N_10193,N_10092);
xor U13503 (N_13503,N_10669,N_10849);
nand U13504 (N_13504,N_11883,N_10271);
nor U13505 (N_13505,N_10787,N_11501);
nand U13506 (N_13506,N_10691,N_10698);
or U13507 (N_13507,N_10280,N_11009);
or U13508 (N_13508,N_11079,N_10846);
nand U13509 (N_13509,N_10068,N_10704);
or U13510 (N_13510,N_11850,N_10761);
nor U13511 (N_13511,N_10738,N_11246);
xor U13512 (N_13512,N_10350,N_11421);
xnor U13513 (N_13513,N_11416,N_10298);
nor U13514 (N_13514,N_10311,N_11658);
or U13515 (N_13515,N_10886,N_10661);
or U13516 (N_13516,N_11098,N_11406);
and U13517 (N_13517,N_10545,N_11224);
xor U13518 (N_13518,N_10661,N_10617);
and U13519 (N_13519,N_11478,N_11381);
and U13520 (N_13520,N_11152,N_11003);
xnor U13521 (N_13521,N_11646,N_10315);
nor U13522 (N_13522,N_11980,N_10906);
nor U13523 (N_13523,N_11735,N_10658);
nor U13524 (N_13524,N_10578,N_11434);
or U13525 (N_13525,N_11170,N_10042);
and U13526 (N_13526,N_11521,N_11416);
or U13527 (N_13527,N_10287,N_10649);
nand U13528 (N_13528,N_11755,N_10834);
or U13529 (N_13529,N_10066,N_10806);
xnor U13530 (N_13530,N_11461,N_11656);
and U13531 (N_13531,N_10782,N_11982);
nand U13532 (N_13532,N_10387,N_10787);
nor U13533 (N_13533,N_11556,N_10374);
nand U13534 (N_13534,N_11242,N_10725);
xor U13535 (N_13535,N_10727,N_11992);
and U13536 (N_13536,N_11300,N_10939);
nor U13537 (N_13537,N_10069,N_11765);
or U13538 (N_13538,N_11348,N_11017);
xor U13539 (N_13539,N_10024,N_10445);
xnor U13540 (N_13540,N_10617,N_10570);
nand U13541 (N_13541,N_11364,N_11716);
nand U13542 (N_13542,N_11354,N_11361);
and U13543 (N_13543,N_11070,N_10980);
nor U13544 (N_13544,N_10025,N_10378);
xor U13545 (N_13545,N_10917,N_11152);
nand U13546 (N_13546,N_10168,N_10307);
nor U13547 (N_13547,N_10367,N_10506);
and U13548 (N_13548,N_11727,N_11939);
or U13549 (N_13549,N_11472,N_10900);
xor U13550 (N_13550,N_11855,N_11843);
or U13551 (N_13551,N_11666,N_10557);
and U13552 (N_13552,N_11040,N_10787);
or U13553 (N_13553,N_11430,N_10140);
xnor U13554 (N_13554,N_11777,N_11947);
nand U13555 (N_13555,N_11154,N_11695);
xor U13556 (N_13556,N_10231,N_10483);
nand U13557 (N_13557,N_10219,N_11821);
xor U13558 (N_13558,N_11173,N_11314);
and U13559 (N_13559,N_10735,N_10187);
xor U13560 (N_13560,N_11541,N_10081);
nor U13561 (N_13561,N_10726,N_10927);
or U13562 (N_13562,N_10393,N_10674);
xor U13563 (N_13563,N_10191,N_11524);
or U13564 (N_13564,N_10171,N_10244);
or U13565 (N_13565,N_11609,N_10882);
or U13566 (N_13566,N_11394,N_10843);
xnor U13567 (N_13567,N_11645,N_10482);
and U13568 (N_13568,N_11553,N_10701);
or U13569 (N_13569,N_10710,N_10069);
or U13570 (N_13570,N_11209,N_10931);
and U13571 (N_13571,N_10659,N_11230);
nor U13572 (N_13572,N_11970,N_11516);
or U13573 (N_13573,N_11121,N_11746);
xnor U13574 (N_13574,N_10242,N_10240);
xnor U13575 (N_13575,N_11559,N_11663);
nor U13576 (N_13576,N_11043,N_11359);
and U13577 (N_13577,N_10316,N_11991);
nand U13578 (N_13578,N_10568,N_10333);
nor U13579 (N_13579,N_10481,N_11323);
nand U13580 (N_13580,N_11464,N_11471);
or U13581 (N_13581,N_11498,N_10103);
and U13582 (N_13582,N_11339,N_10471);
and U13583 (N_13583,N_11555,N_10387);
nor U13584 (N_13584,N_10658,N_11662);
and U13585 (N_13585,N_11943,N_10548);
nor U13586 (N_13586,N_10920,N_11928);
and U13587 (N_13587,N_11143,N_11111);
or U13588 (N_13588,N_11877,N_10289);
or U13589 (N_13589,N_10624,N_10269);
nand U13590 (N_13590,N_11959,N_11757);
or U13591 (N_13591,N_10614,N_11152);
and U13592 (N_13592,N_11456,N_10388);
or U13593 (N_13593,N_10846,N_10596);
xnor U13594 (N_13594,N_10776,N_11473);
or U13595 (N_13595,N_11706,N_11458);
nand U13596 (N_13596,N_10848,N_11533);
xnor U13597 (N_13597,N_11836,N_11856);
xor U13598 (N_13598,N_11568,N_10754);
nor U13599 (N_13599,N_10879,N_11170);
nand U13600 (N_13600,N_11466,N_11097);
or U13601 (N_13601,N_11896,N_11125);
and U13602 (N_13602,N_10390,N_11919);
nor U13603 (N_13603,N_11506,N_10641);
nor U13604 (N_13604,N_11030,N_10011);
or U13605 (N_13605,N_11239,N_11511);
nor U13606 (N_13606,N_10590,N_10894);
and U13607 (N_13607,N_11883,N_11611);
or U13608 (N_13608,N_10582,N_10735);
nor U13609 (N_13609,N_10075,N_10806);
nor U13610 (N_13610,N_10605,N_11424);
nand U13611 (N_13611,N_10691,N_10147);
nor U13612 (N_13612,N_10905,N_11110);
nand U13613 (N_13613,N_11364,N_11623);
nor U13614 (N_13614,N_10341,N_11601);
nand U13615 (N_13615,N_10451,N_10831);
nor U13616 (N_13616,N_11903,N_11283);
nor U13617 (N_13617,N_11732,N_11573);
nand U13618 (N_13618,N_11670,N_11699);
and U13619 (N_13619,N_10658,N_10614);
nor U13620 (N_13620,N_10869,N_10991);
nor U13621 (N_13621,N_10313,N_10469);
nand U13622 (N_13622,N_10364,N_11489);
xor U13623 (N_13623,N_10570,N_11867);
and U13624 (N_13624,N_11985,N_10942);
nor U13625 (N_13625,N_10582,N_11615);
xor U13626 (N_13626,N_10602,N_10829);
and U13627 (N_13627,N_10172,N_10291);
xor U13628 (N_13628,N_10148,N_11828);
xnor U13629 (N_13629,N_11379,N_10537);
nor U13630 (N_13630,N_10161,N_11927);
xor U13631 (N_13631,N_11371,N_11124);
nor U13632 (N_13632,N_11273,N_10489);
or U13633 (N_13633,N_10692,N_11425);
nand U13634 (N_13634,N_11273,N_11114);
xnor U13635 (N_13635,N_10933,N_11317);
xnor U13636 (N_13636,N_11359,N_11181);
nor U13637 (N_13637,N_10959,N_10551);
nand U13638 (N_13638,N_11743,N_11521);
and U13639 (N_13639,N_11948,N_11420);
or U13640 (N_13640,N_11211,N_10906);
nor U13641 (N_13641,N_11471,N_10936);
or U13642 (N_13642,N_11109,N_10596);
nand U13643 (N_13643,N_10364,N_11868);
nand U13644 (N_13644,N_11920,N_11382);
and U13645 (N_13645,N_10855,N_11547);
and U13646 (N_13646,N_10681,N_11088);
nor U13647 (N_13647,N_10816,N_11323);
or U13648 (N_13648,N_11768,N_11649);
nor U13649 (N_13649,N_10514,N_10981);
or U13650 (N_13650,N_10924,N_10876);
nor U13651 (N_13651,N_10941,N_10043);
xnor U13652 (N_13652,N_11173,N_11911);
xnor U13653 (N_13653,N_10527,N_10387);
or U13654 (N_13654,N_10503,N_10289);
xor U13655 (N_13655,N_10190,N_11141);
nor U13656 (N_13656,N_10244,N_10132);
nand U13657 (N_13657,N_10631,N_10478);
nand U13658 (N_13658,N_10906,N_11175);
nor U13659 (N_13659,N_11062,N_10098);
nor U13660 (N_13660,N_10606,N_11415);
and U13661 (N_13661,N_11994,N_10982);
nand U13662 (N_13662,N_10452,N_11331);
and U13663 (N_13663,N_10311,N_10667);
or U13664 (N_13664,N_11868,N_10204);
or U13665 (N_13665,N_10447,N_11982);
nand U13666 (N_13666,N_10732,N_10102);
and U13667 (N_13667,N_11371,N_11545);
nor U13668 (N_13668,N_10493,N_10205);
nand U13669 (N_13669,N_11127,N_10939);
or U13670 (N_13670,N_11402,N_11917);
nor U13671 (N_13671,N_10094,N_10541);
or U13672 (N_13672,N_11477,N_10803);
nor U13673 (N_13673,N_10262,N_10499);
xor U13674 (N_13674,N_11670,N_11746);
or U13675 (N_13675,N_10750,N_11762);
and U13676 (N_13676,N_10199,N_10128);
nor U13677 (N_13677,N_11558,N_11287);
and U13678 (N_13678,N_10215,N_11818);
and U13679 (N_13679,N_11351,N_11070);
xnor U13680 (N_13680,N_11155,N_10107);
xnor U13681 (N_13681,N_11366,N_10180);
nand U13682 (N_13682,N_10711,N_11015);
or U13683 (N_13683,N_11375,N_10046);
or U13684 (N_13684,N_10087,N_10065);
and U13685 (N_13685,N_10991,N_10551);
and U13686 (N_13686,N_10285,N_11138);
and U13687 (N_13687,N_11043,N_11548);
or U13688 (N_13688,N_10887,N_10804);
or U13689 (N_13689,N_10058,N_11786);
nor U13690 (N_13690,N_10739,N_10305);
nor U13691 (N_13691,N_11309,N_11978);
or U13692 (N_13692,N_10335,N_11290);
and U13693 (N_13693,N_10088,N_11161);
xor U13694 (N_13694,N_10404,N_10601);
or U13695 (N_13695,N_11420,N_11427);
or U13696 (N_13696,N_11063,N_11277);
and U13697 (N_13697,N_11464,N_10291);
and U13698 (N_13698,N_11805,N_10201);
nor U13699 (N_13699,N_10595,N_11803);
nand U13700 (N_13700,N_10146,N_10672);
xnor U13701 (N_13701,N_10229,N_10930);
xnor U13702 (N_13702,N_11982,N_10369);
or U13703 (N_13703,N_10427,N_10992);
or U13704 (N_13704,N_10690,N_10293);
xnor U13705 (N_13705,N_10793,N_10660);
nor U13706 (N_13706,N_10963,N_10169);
and U13707 (N_13707,N_11826,N_11497);
nor U13708 (N_13708,N_11919,N_10397);
and U13709 (N_13709,N_10394,N_11004);
nor U13710 (N_13710,N_11219,N_11728);
xor U13711 (N_13711,N_11495,N_10539);
nand U13712 (N_13712,N_11425,N_10275);
nor U13713 (N_13713,N_11357,N_11460);
xnor U13714 (N_13714,N_11553,N_10886);
or U13715 (N_13715,N_11141,N_11262);
nand U13716 (N_13716,N_11485,N_10720);
nor U13717 (N_13717,N_11977,N_10451);
and U13718 (N_13718,N_11843,N_10569);
nor U13719 (N_13719,N_10820,N_11093);
xnor U13720 (N_13720,N_11074,N_10946);
nor U13721 (N_13721,N_11403,N_10110);
and U13722 (N_13722,N_11344,N_10609);
and U13723 (N_13723,N_10114,N_10311);
nand U13724 (N_13724,N_11986,N_11434);
nor U13725 (N_13725,N_10251,N_11402);
xnor U13726 (N_13726,N_11279,N_10283);
nor U13727 (N_13727,N_10858,N_10320);
or U13728 (N_13728,N_11311,N_11298);
nand U13729 (N_13729,N_10523,N_10559);
xnor U13730 (N_13730,N_11234,N_10056);
nor U13731 (N_13731,N_11960,N_10846);
nor U13732 (N_13732,N_10264,N_10019);
and U13733 (N_13733,N_11606,N_10371);
xor U13734 (N_13734,N_11346,N_11837);
nand U13735 (N_13735,N_11032,N_11408);
nand U13736 (N_13736,N_10746,N_11811);
and U13737 (N_13737,N_10452,N_10165);
xnor U13738 (N_13738,N_11116,N_11622);
xnor U13739 (N_13739,N_11801,N_11745);
nand U13740 (N_13740,N_10335,N_11502);
and U13741 (N_13741,N_10329,N_10700);
nor U13742 (N_13742,N_11141,N_11632);
xnor U13743 (N_13743,N_11253,N_11601);
and U13744 (N_13744,N_11730,N_10721);
nor U13745 (N_13745,N_10191,N_10479);
and U13746 (N_13746,N_10681,N_11197);
or U13747 (N_13747,N_11878,N_10585);
or U13748 (N_13748,N_10549,N_10225);
nand U13749 (N_13749,N_11033,N_10665);
nand U13750 (N_13750,N_10318,N_11534);
nor U13751 (N_13751,N_11405,N_10809);
or U13752 (N_13752,N_10428,N_10034);
nor U13753 (N_13753,N_10154,N_10355);
xor U13754 (N_13754,N_10538,N_11989);
nand U13755 (N_13755,N_10023,N_10846);
and U13756 (N_13756,N_10859,N_11129);
xnor U13757 (N_13757,N_10503,N_10291);
or U13758 (N_13758,N_11826,N_11343);
xnor U13759 (N_13759,N_10306,N_10023);
or U13760 (N_13760,N_10502,N_11845);
nor U13761 (N_13761,N_11414,N_11317);
nor U13762 (N_13762,N_10159,N_10846);
nand U13763 (N_13763,N_11303,N_11931);
and U13764 (N_13764,N_11541,N_10717);
xor U13765 (N_13765,N_11433,N_11499);
nand U13766 (N_13766,N_11213,N_10506);
nor U13767 (N_13767,N_11098,N_11902);
xor U13768 (N_13768,N_11236,N_10061);
nand U13769 (N_13769,N_10305,N_10905);
nor U13770 (N_13770,N_10815,N_11953);
nand U13771 (N_13771,N_10110,N_10546);
xor U13772 (N_13772,N_10258,N_10291);
nand U13773 (N_13773,N_10967,N_10302);
nand U13774 (N_13774,N_11238,N_11879);
and U13775 (N_13775,N_11204,N_10649);
or U13776 (N_13776,N_10135,N_10427);
nor U13777 (N_13777,N_11803,N_11940);
or U13778 (N_13778,N_10134,N_11935);
nor U13779 (N_13779,N_11779,N_10347);
nor U13780 (N_13780,N_10259,N_11432);
or U13781 (N_13781,N_11798,N_10822);
nor U13782 (N_13782,N_10841,N_10580);
xnor U13783 (N_13783,N_11570,N_10131);
nor U13784 (N_13784,N_10905,N_10323);
nor U13785 (N_13785,N_11159,N_10780);
nor U13786 (N_13786,N_10293,N_10264);
nand U13787 (N_13787,N_11072,N_11480);
nor U13788 (N_13788,N_10282,N_10992);
and U13789 (N_13789,N_10955,N_10719);
and U13790 (N_13790,N_10395,N_11169);
or U13791 (N_13791,N_10290,N_11852);
xor U13792 (N_13792,N_11639,N_10406);
and U13793 (N_13793,N_11584,N_11591);
or U13794 (N_13794,N_10776,N_10959);
or U13795 (N_13795,N_11231,N_10462);
xor U13796 (N_13796,N_10605,N_11463);
nand U13797 (N_13797,N_11465,N_11243);
xnor U13798 (N_13798,N_10533,N_11753);
or U13799 (N_13799,N_10581,N_10368);
nor U13800 (N_13800,N_11700,N_10647);
nand U13801 (N_13801,N_10525,N_10553);
nor U13802 (N_13802,N_11440,N_10409);
xor U13803 (N_13803,N_10453,N_11463);
nand U13804 (N_13804,N_11973,N_10208);
and U13805 (N_13805,N_10459,N_11438);
nand U13806 (N_13806,N_10490,N_11048);
and U13807 (N_13807,N_10485,N_11599);
and U13808 (N_13808,N_11037,N_10549);
or U13809 (N_13809,N_11211,N_10708);
xnor U13810 (N_13810,N_10782,N_10441);
xor U13811 (N_13811,N_10027,N_11582);
xnor U13812 (N_13812,N_10911,N_11875);
nand U13813 (N_13813,N_11984,N_10536);
nor U13814 (N_13814,N_10839,N_10677);
nor U13815 (N_13815,N_11133,N_10468);
and U13816 (N_13816,N_11119,N_11662);
and U13817 (N_13817,N_11756,N_10894);
or U13818 (N_13818,N_10965,N_10401);
and U13819 (N_13819,N_11032,N_10713);
or U13820 (N_13820,N_11988,N_11336);
xnor U13821 (N_13821,N_11922,N_11672);
and U13822 (N_13822,N_10894,N_10412);
or U13823 (N_13823,N_10471,N_11447);
xor U13824 (N_13824,N_11208,N_10740);
and U13825 (N_13825,N_10525,N_10000);
and U13826 (N_13826,N_11374,N_10616);
or U13827 (N_13827,N_11328,N_10786);
or U13828 (N_13828,N_10088,N_10033);
and U13829 (N_13829,N_11337,N_11770);
nor U13830 (N_13830,N_11090,N_11286);
nand U13831 (N_13831,N_10150,N_11275);
and U13832 (N_13832,N_10260,N_11744);
or U13833 (N_13833,N_10724,N_11790);
nand U13834 (N_13834,N_10256,N_10149);
nand U13835 (N_13835,N_10208,N_11313);
and U13836 (N_13836,N_10925,N_10884);
and U13837 (N_13837,N_10837,N_10366);
and U13838 (N_13838,N_11609,N_10551);
or U13839 (N_13839,N_11173,N_10569);
and U13840 (N_13840,N_11225,N_10265);
nor U13841 (N_13841,N_11941,N_10172);
or U13842 (N_13842,N_10326,N_10630);
or U13843 (N_13843,N_11892,N_10820);
nor U13844 (N_13844,N_11294,N_10225);
nor U13845 (N_13845,N_10428,N_10680);
xnor U13846 (N_13846,N_11035,N_11763);
and U13847 (N_13847,N_10417,N_11805);
or U13848 (N_13848,N_10977,N_10744);
xor U13849 (N_13849,N_11726,N_10860);
nor U13850 (N_13850,N_10813,N_11169);
xor U13851 (N_13851,N_10074,N_10723);
and U13852 (N_13852,N_11027,N_11926);
nand U13853 (N_13853,N_10202,N_10806);
xnor U13854 (N_13854,N_10779,N_10345);
nand U13855 (N_13855,N_10975,N_10622);
and U13856 (N_13856,N_10393,N_10975);
and U13857 (N_13857,N_11577,N_11993);
xor U13858 (N_13858,N_11531,N_11649);
xnor U13859 (N_13859,N_10694,N_11456);
or U13860 (N_13860,N_11636,N_10034);
or U13861 (N_13861,N_10763,N_10865);
and U13862 (N_13862,N_10062,N_10366);
and U13863 (N_13863,N_10450,N_11770);
or U13864 (N_13864,N_10260,N_10659);
nor U13865 (N_13865,N_10228,N_10029);
nor U13866 (N_13866,N_11746,N_11797);
and U13867 (N_13867,N_10679,N_10099);
nand U13868 (N_13868,N_11334,N_11434);
nand U13869 (N_13869,N_11897,N_10087);
nor U13870 (N_13870,N_10500,N_11517);
nor U13871 (N_13871,N_11424,N_10825);
and U13872 (N_13872,N_11625,N_10033);
nor U13873 (N_13873,N_11805,N_10603);
xnor U13874 (N_13874,N_11980,N_10260);
or U13875 (N_13875,N_10771,N_11969);
xnor U13876 (N_13876,N_10344,N_11226);
xnor U13877 (N_13877,N_11786,N_10093);
or U13878 (N_13878,N_11359,N_11538);
or U13879 (N_13879,N_10812,N_10426);
nand U13880 (N_13880,N_11708,N_11401);
or U13881 (N_13881,N_11966,N_10683);
and U13882 (N_13882,N_11456,N_10405);
nor U13883 (N_13883,N_11178,N_10169);
xnor U13884 (N_13884,N_10835,N_11374);
nand U13885 (N_13885,N_11124,N_11087);
nand U13886 (N_13886,N_10520,N_11041);
nor U13887 (N_13887,N_10341,N_10639);
and U13888 (N_13888,N_10736,N_10626);
nand U13889 (N_13889,N_10450,N_10513);
nor U13890 (N_13890,N_11122,N_11010);
or U13891 (N_13891,N_10315,N_11623);
and U13892 (N_13892,N_11095,N_11756);
nand U13893 (N_13893,N_10056,N_10161);
and U13894 (N_13894,N_10204,N_10677);
or U13895 (N_13895,N_10712,N_11644);
xnor U13896 (N_13896,N_10817,N_10592);
and U13897 (N_13897,N_11303,N_11819);
nand U13898 (N_13898,N_10838,N_10336);
or U13899 (N_13899,N_10431,N_10612);
xnor U13900 (N_13900,N_11177,N_11657);
nand U13901 (N_13901,N_10458,N_10337);
xor U13902 (N_13902,N_11340,N_10937);
nor U13903 (N_13903,N_10406,N_11465);
xor U13904 (N_13904,N_11331,N_11096);
xnor U13905 (N_13905,N_10081,N_11683);
and U13906 (N_13906,N_11644,N_10910);
xor U13907 (N_13907,N_11112,N_10491);
nand U13908 (N_13908,N_11703,N_10539);
or U13909 (N_13909,N_11412,N_11907);
nor U13910 (N_13910,N_10798,N_10805);
and U13911 (N_13911,N_10989,N_11309);
xnor U13912 (N_13912,N_11728,N_11122);
xor U13913 (N_13913,N_10033,N_11304);
nor U13914 (N_13914,N_11574,N_10677);
xor U13915 (N_13915,N_11170,N_11914);
nand U13916 (N_13916,N_11578,N_11607);
or U13917 (N_13917,N_10173,N_10780);
nor U13918 (N_13918,N_11911,N_10887);
nand U13919 (N_13919,N_10103,N_11041);
nor U13920 (N_13920,N_11039,N_11534);
nor U13921 (N_13921,N_10308,N_10521);
and U13922 (N_13922,N_11931,N_11895);
and U13923 (N_13923,N_11115,N_10604);
and U13924 (N_13924,N_11238,N_11212);
or U13925 (N_13925,N_11318,N_11007);
nor U13926 (N_13926,N_10169,N_11223);
xor U13927 (N_13927,N_11835,N_10608);
nand U13928 (N_13928,N_11609,N_11109);
or U13929 (N_13929,N_11943,N_11338);
or U13930 (N_13930,N_10190,N_10049);
nand U13931 (N_13931,N_11902,N_10477);
nor U13932 (N_13932,N_10604,N_10176);
and U13933 (N_13933,N_10499,N_10440);
and U13934 (N_13934,N_11013,N_10182);
xor U13935 (N_13935,N_10578,N_10198);
nand U13936 (N_13936,N_10917,N_10528);
nor U13937 (N_13937,N_11282,N_11850);
or U13938 (N_13938,N_11209,N_10778);
xnor U13939 (N_13939,N_11345,N_10061);
xor U13940 (N_13940,N_11733,N_10473);
or U13941 (N_13941,N_11394,N_10736);
or U13942 (N_13942,N_10761,N_11493);
nor U13943 (N_13943,N_10370,N_10491);
nor U13944 (N_13944,N_10808,N_11834);
and U13945 (N_13945,N_10739,N_11548);
nor U13946 (N_13946,N_10584,N_10449);
nand U13947 (N_13947,N_10289,N_10759);
xnor U13948 (N_13948,N_10240,N_11030);
and U13949 (N_13949,N_10915,N_11517);
and U13950 (N_13950,N_11373,N_10720);
and U13951 (N_13951,N_10169,N_11994);
nor U13952 (N_13952,N_11570,N_10935);
or U13953 (N_13953,N_10315,N_10741);
nand U13954 (N_13954,N_11443,N_11240);
xnor U13955 (N_13955,N_10135,N_11534);
and U13956 (N_13956,N_10672,N_11672);
nand U13957 (N_13957,N_11379,N_10675);
nand U13958 (N_13958,N_10945,N_11513);
nand U13959 (N_13959,N_11688,N_11678);
or U13960 (N_13960,N_11033,N_11048);
or U13961 (N_13961,N_10350,N_11992);
and U13962 (N_13962,N_11141,N_10568);
nor U13963 (N_13963,N_11250,N_11654);
nor U13964 (N_13964,N_11658,N_10168);
nor U13965 (N_13965,N_11160,N_11050);
xnor U13966 (N_13966,N_10146,N_10046);
and U13967 (N_13967,N_11591,N_11483);
nand U13968 (N_13968,N_10496,N_10332);
or U13969 (N_13969,N_10712,N_11882);
nand U13970 (N_13970,N_10929,N_10216);
nand U13971 (N_13971,N_10995,N_10480);
and U13972 (N_13972,N_10676,N_11145);
or U13973 (N_13973,N_11968,N_11038);
xor U13974 (N_13974,N_10484,N_10692);
or U13975 (N_13975,N_10388,N_10934);
nor U13976 (N_13976,N_10160,N_10688);
nor U13977 (N_13977,N_10737,N_10519);
or U13978 (N_13978,N_10047,N_10450);
or U13979 (N_13979,N_11887,N_11531);
xnor U13980 (N_13980,N_10199,N_11623);
xnor U13981 (N_13981,N_11876,N_11217);
xor U13982 (N_13982,N_11422,N_10927);
and U13983 (N_13983,N_10255,N_11851);
or U13984 (N_13984,N_11843,N_11052);
and U13985 (N_13985,N_11057,N_10684);
xnor U13986 (N_13986,N_11347,N_11456);
and U13987 (N_13987,N_10275,N_11072);
nand U13988 (N_13988,N_10119,N_10094);
and U13989 (N_13989,N_10625,N_11598);
nor U13990 (N_13990,N_10957,N_11400);
xor U13991 (N_13991,N_11833,N_10763);
xnor U13992 (N_13992,N_10453,N_11214);
xor U13993 (N_13993,N_10926,N_10610);
or U13994 (N_13994,N_11121,N_10323);
nor U13995 (N_13995,N_11687,N_11617);
or U13996 (N_13996,N_11184,N_11358);
nand U13997 (N_13997,N_10467,N_10507);
xor U13998 (N_13998,N_11399,N_10383);
nor U13999 (N_13999,N_11698,N_10286);
and U14000 (N_14000,N_12133,N_12493);
nor U14001 (N_14001,N_12809,N_12629);
and U14002 (N_14002,N_13407,N_13727);
or U14003 (N_14003,N_13570,N_13314);
or U14004 (N_14004,N_13410,N_13749);
nand U14005 (N_14005,N_12881,N_13213);
and U14006 (N_14006,N_13331,N_12300);
xnor U14007 (N_14007,N_12069,N_13211);
nor U14008 (N_14008,N_12323,N_12696);
nor U14009 (N_14009,N_13506,N_12174);
xnor U14010 (N_14010,N_13345,N_12984);
nand U14011 (N_14011,N_13724,N_13029);
and U14012 (N_14012,N_12238,N_12622);
or U14013 (N_14013,N_12105,N_13043);
xor U14014 (N_14014,N_12660,N_12306);
and U14015 (N_14015,N_13040,N_12876);
and U14016 (N_14016,N_13937,N_12945);
nor U14017 (N_14017,N_12823,N_12920);
and U14018 (N_14018,N_13542,N_13698);
xnor U14019 (N_14019,N_13150,N_12373);
nor U14020 (N_14020,N_13223,N_12036);
or U14021 (N_14021,N_12934,N_13630);
and U14022 (N_14022,N_13028,N_13057);
nor U14023 (N_14023,N_13599,N_12387);
xor U14024 (N_14024,N_13725,N_12588);
nor U14025 (N_14025,N_12040,N_12969);
nand U14026 (N_14026,N_13188,N_12748);
xor U14027 (N_14027,N_12094,N_13585);
nor U14028 (N_14028,N_12200,N_13397);
xor U14029 (N_14029,N_13647,N_13851);
nor U14030 (N_14030,N_13025,N_13549);
nor U14031 (N_14031,N_13837,N_13988);
or U14032 (N_14032,N_13858,N_12634);
nor U14033 (N_14033,N_13998,N_13751);
nor U14034 (N_14034,N_13127,N_12194);
or U14035 (N_14035,N_12366,N_12245);
nand U14036 (N_14036,N_12569,N_13203);
and U14037 (N_14037,N_12193,N_12861);
and U14038 (N_14038,N_12271,N_12162);
or U14039 (N_14039,N_12883,N_12107);
nand U14040 (N_14040,N_13441,N_13867);
nor U14041 (N_14041,N_13960,N_12348);
or U14042 (N_14042,N_12285,N_13856);
and U14043 (N_14043,N_13604,N_12740);
or U14044 (N_14044,N_12335,N_12146);
or U14045 (N_14045,N_13050,N_13058);
xnor U14046 (N_14046,N_12466,N_13174);
or U14047 (N_14047,N_12835,N_13182);
xor U14048 (N_14048,N_12307,N_12381);
nor U14049 (N_14049,N_13201,N_12134);
nor U14050 (N_14050,N_13202,N_13635);
xor U14051 (N_14051,N_13034,N_13171);
xnor U14052 (N_14052,N_13242,N_12706);
nor U14053 (N_14053,N_13634,N_13500);
or U14054 (N_14054,N_12091,N_12982);
nand U14055 (N_14055,N_12743,N_12456);
nand U14056 (N_14056,N_13009,N_13513);
nor U14057 (N_14057,N_12216,N_13421);
or U14058 (N_14058,N_13085,N_12243);
nor U14059 (N_14059,N_12824,N_13146);
xor U14060 (N_14060,N_13437,N_13245);
xnor U14061 (N_14061,N_12154,N_12548);
or U14062 (N_14062,N_13673,N_12914);
and U14063 (N_14063,N_13183,N_12848);
nor U14064 (N_14064,N_12668,N_12693);
or U14065 (N_14065,N_12630,N_13566);
xor U14066 (N_14066,N_12450,N_12050);
nand U14067 (N_14067,N_13319,N_13024);
nand U14068 (N_14068,N_13655,N_12111);
nand U14069 (N_14069,N_13498,N_12645);
nand U14070 (N_14070,N_13853,N_12427);
or U14071 (N_14071,N_13115,N_12151);
or U14072 (N_14072,N_12714,N_13310);
xor U14073 (N_14073,N_12556,N_12142);
nor U14074 (N_14074,N_13576,N_13370);
or U14075 (N_14075,N_13790,N_12175);
and U14076 (N_14076,N_12022,N_13265);
and U14077 (N_14077,N_13446,N_12061);
or U14078 (N_14078,N_13989,N_13660);
nor U14079 (N_14079,N_12892,N_13362);
or U14080 (N_14080,N_12447,N_13518);
nor U14081 (N_14081,N_13160,N_12899);
nor U14082 (N_14082,N_13677,N_12426);
nand U14083 (N_14083,N_13237,N_12415);
xor U14084 (N_14084,N_13470,N_12709);
nor U14085 (N_14085,N_13328,N_12988);
xor U14086 (N_14086,N_13391,N_12430);
nor U14087 (N_14087,N_12698,N_13944);
nand U14088 (N_14088,N_13194,N_12993);
nand U14089 (N_14089,N_12636,N_13846);
and U14090 (N_14090,N_13109,N_12078);
or U14091 (N_14091,N_12852,N_13266);
nand U14092 (N_14092,N_12670,N_13772);
nor U14093 (N_14093,N_13783,N_13735);
or U14094 (N_14094,N_13015,N_13017);
nand U14095 (N_14095,N_12128,N_12541);
or U14096 (N_14096,N_12785,N_13209);
and U14097 (N_14097,N_13049,N_13950);
or U14098 (N_14098,N_12972,N_13756);
nor U14099 (N_14099,N_13426,N_12839);
nor U14100 (N_14100,N_12788,N_13807);
xnor U14101 (N_14101,N_13380,N_13584);
or U14102 (N_14102,N_12955,N_13385);
xor U14103 (N_14103,N_13167,N_12429);
or U14104 (N_14104,N_12234,N_13369);
and U14105 (N_14105,N_12321,N_12408);
nor U14106 (N_14106,N_13704,N_12318);
nand U14107 (N_14107,N_12682,N_13792);
nor U14108 (N_14108,N_13555,N_12518);
nand U14109 (N_14109,N_13102,N_13991);
xor U14110 (N_14110,N_13767,N_13639);
or U14111 (N_14111,N_12544,N_12815);
nor U14112 (N_14112,N_12363,N_12560);
nand U14113 (N_14113,N_13198,N_13350);
nor U14114 (N_14114,N_12991,N_12229);
xor U14115 (N_14115,N_12747,N_12741);
or U14116 (N_14116,N_13746,N_13948);
nand U14117 (N_14117,N_13092,N_13341);
xor U14118 (N_14118,N_12762,N_12946);
nor U14119 (N_14119,N_12202,N_12821);
and U14120 (N_14120,N_12566,N_13803);
xnor U14121 (N_14121,N_13912,N_13308);
nor U14122 (N_14122,N_13804,N_12587);
xor U14123 (N_14123,N_13327,N_13760);
or U14124 (N_14124,N_13149,N_13762);
nor U14125 (N_14125,N_13221,N_12517);
xnor U14126 (N_14126,N_12780,N_13687);
xnor U14127 (N_14127,N_12547,N_13436);
nand U14128 (N_14128,N_12010,N_13931);
or U14129 (N_14129,N_12656,N_12840);
and U14130 (N_14130,N_12025,N_12642);
and U14131 (N_14131,N_13911,N_13489);
nand U14132 (N_14132,N_13935,N_12192);
nor U14133 (N_14133,N_12973,N_12394);
xor U14134 (N_14134,N_13039,N_12330);
or U14135 (N_14135,N_13228,N_13965);
and U14136 (N_14136,N_13486,N_12295);
xnor U14137 (N_14137,N_13164,N_13121);
xnor U14138 (N_14138,N_13631,N_12378);
and U14139 (N_14139,N_12451,N_13514);
or U14140 (N_14140,N_13206,N_12879);
or U14141 (N_14141,N_13439,N_13882);
nand U14142 (N_14142,N_13993,N_13154);
nor U14143 (N_14143,N_13306,N_12964);
xor U14144 (N_14144,N_12958,N_12008);
and U14145 (N_14145,N_12506,N_12737);
or U14146 (N_14146,N_13929,N_13877);
xor U14147 (N_14147,N_12292,N_13214);
xor U14148 (N_14148,N_12145,N_13204);
or U14149 (N_14149,N_13754,N_12853);
or U14150 (N_14150,N_13969,N_12789);
nor U14151 (N_14151,N_12500,N_13716);
nor U14152 (N_14152,N_13387,N_12303);
and U14153 (N_14153,N_13384,N_12716);
xor U14154 (N_14154,N_13855,N_13609);
nand U14155 (N_14155,N_13823,N_13278);
and U14156 (N_14156,N_13822,N_12819);
xor U14157 (N_14157,N_13842,N_13197);
nand U14158 (N_14158,N_12441,N_13689);
and U14159 (N_14159,N_12023,N_13508);
and U14160 (N_14160,N_13685,N_13818);
nor U14161 (N_14161,N_13707,N_13742);
xor U14162 (N_14162,N_12087,N_13545);
and U14163 (N_14163,N_13006,N_12607);
or U14164 (N_14164,N_13693,N_12404);
nand U14165 (N_14165,N_12974,N_12294);
nor U14166 (N_14166,N_13982,N_12293);
xor U14167 (N_14167,N_12123,N_12051);
nor U14168 (N_14168,N_13699,N_12334);
and U14169 (N_14169,N_12116,N_13868);
nor U14170 (N_14170,N_13761,N_13475);
and U14171 (N_14171,N_12906,N_12227);
xnor U14172 (N_14172,N_13431,N_13927);
nand U14173 (N_14173,N_13451,N_13744);
and U14174 (N_14174,N_13591,N_12398);
and U14175 (N_14175,N_13193,N_12726);
xnor U14176 (N_14176,N_12802,N_13554);
and U14177 (N_14177,N_12437,N_12937);
or U14178 (N_14178,N_12392,N_13984);
nor U14179 (N_14179,N_13978,N_13658);
nand U14180 (N_14180,N_12113,N_12921);
or U14181 (N_14181,N_13524,N_13357);
and U14182 (N_14182,N_12522,N_12046);
nor U14183 (N_14183,N_13255,N_12230);
nand U14184 (N_14184,N_12895,N_13659);
nor U14185 (N_14185,N_13074,N_12118);
or U14186 (N_14186,N_12777,N_12073);
xor U14187 (N_14187,N_12922,N_12729);
nor U14188 (N_14188,N_13187,N_13117);
nor U14189 (N_14189,N_12834,N_13657);
nand U14190 (N_14190,N_13540,N_13709);
nor U14191 (N_14191,N_12664,N_13428);
or U14192 (N_14192,N_12890,N_13128);
nor U14193 (N_14193,N_12244,N_13963);
and U14194 (N_14194,N_13987,N_13483);
and U14195 (N_14195,N_12672,N_12844);
xnor U14196 (N_14196,N_13056,N_12505);
nand U14197 (N_14197,N_13316,N_13132);
nor U14198 (N_14198,N_12658,N_12106);
xnor U14199 (N_14199,N_13741,N_12951);
xnor U14200 (N_14200,N_13063,N_13095);
xnor U14201 (N_14201,N_13184,N_12024);
and U14202 (N_14202,N_12822,N_12529);
and U14203 (N_14203,N_13977,N_13442);
or U14204 (N_14204,N_12894,N_12346);
nand U14205 (N_14205,N_13682,N_13841);
xor U14206 (N_14206,N_12110,N_12643);
xor U14207 (N_14207,N_12851,N_13324);
nand U14208 (N_14208,N_13582,N_13898);
or U14209 (N_14209,N_12262,N_13493);
nand U14210 (N_14210,N_13053,N_12979);
nand U14211 (N_14211,N_12268,N_12021);
xnor U14212 (N_14212,N_12962,N_12764);
or U14213 (N_14213,N_13669,N_13852);
xor U14214 (N_14214,N_13145,N_12459);
or U14215 (N_14215,N_12273,N_12076);
and U14216 (N_14216,N_13798,N_12157);
nand U14217 (N_14217,N_13601,N_12872);
and U14218 (N_14218,N_12375,N_13219);
nor U14219 (N_14219,N_13408,N_12768);
or U14220 (N_14220,N_13967,N_13976);
nand U14221 (N_14221,N_12240,N_12396);
and U14222 (N_14222,N_13051,N_12058);
or U14223 (N_14223,N_13847,N_13358);
or U14224 (N_14224,N_13482,N_13100);
nor U14225 (N_14225,N_13861,N_12035);
nand U14226 (N_14226,N_12164,N_13487);
xor U14227 (N_14227,N_13550,N_12970);
nor U14228 (N_14228,N_13586,N_12703);
nand U14229 (N_14229,N_12910,N_13398);
or U14230 (N_14230,N_12549,N_12885);
and U14231 (N_14231,N_13654,N_13535);
xor U14232 (N_14232,N_13173,N_13259);
xnor U14233 (N_14233,N_13481,N_13089);
or U14234 (N_14234,N_12976,N_13721);
nand U14235 (N_14235,N_12032,N_12722);
nor U14236 (N_14236,N_13318,N_12911);
nor U14237 (N_14237,N_12048,N_12516);
nand U14238 (N_14238,N_12416,N_12180);
or U14239 (N_14239,N_13008,N_12362);
or U14240 (N_14240,N_13539,N_12096);
nor U14241 (N_14241,N_13466,N_12018);
or U14242 (N_14242,N_13180,N_13469);
and U14243 (N_14243,N_13404,N_13645);
nand U14244 (N_14244,N_12614,N_12882);
or U14245 (N_14245,N_12915,N_13175);
nand U14246 (N_14246,N_13621,N_13217);
or U14247 (N_14247,N_12567,N_12613);
nand U14248 (N_14248,N_13885,N_13515);
or U14249 (N_14249,N_13904,N_13311);
nor U14250 (N_14250,N_12543,N_13819);
or U14251 (N_14251,N_12397,N_12940);
xnor U14252 (N_14252,N_12648,N_12455);
xnor U14253 (N_14253,N_12454,N_12521);
or U14254 (N_14254,N_12558,N_13956);
nand U14255 (N_14255,N_13951,N_12044);
xnor U14256 (N_14256,N_12575,N_13365);
or U14257 (N_14257,N_12790,N_12236);
and U14258 (N_14258,N_13247,N_12152);
nor U14259 (N_14259,N_12727,N_12410);
or U14260 (N_14260,N_12460,N_12043);
and U14261 (N_14261,N_13480,N_13608);
nor U14262 (N_14262,N_12472,N_12352);
or U14263 (N_14263,N_12507,N_12843);
or U14264 (N_14264,N_13892,N_13364);
nand U14265 (N_14265,N_13422,N_13569);
xnor U14266 (N_14266,N_12367,N_12857);
nand U14267 (N_14267,N_12919,N_13523);
xor U14268 (N_14268,N_12605,N_12226);
xor U14269 (N_14269,N_13717,N_12286);
xor U14270 (N_14270,N_12150,N_13884);
nor U14271 (N_14271,N_13771,N_12850);
nor U14272 (N_14272,N_13079,N_12277);
nand U14273 (N_14273,N_13665,N_13003);
and U14274 (N_14274,N_12228,N_12184);
xnor U14275 (N_14275,N_13081,N_12205);
nand U14276 (N_14276,N_13455,N_13135);
xor U14277 (N_14277,N_13828,N_12978);
nor U14278 (N_14278,N_13134,N_12148);
nand U14279 (N_14279,N_12719,N_12807);
nor U14280 (N_14280,N_13919,N_13254);
and U14281 (N_14281,N_13983,N_12222);
nand U14282 (N_14282,N_12684,N_13210);
and U14283 (N_14283,N_13473,N_13690);
xor U14284 (N_14284,N_12440,N_13458);
nor U14285 (N_14285,N_13097,N_13080);
nor U14286 (N_14286,N_12435,N_13276);
nand U14287 (N_14287,N_13200,N_12756);
and U14288 (N_14288,N_12084,N_13383);
nor U14289 (N_14289,N_13844,N_12877);
nor U14290 (N_14290,N_13177,N_13010);
xor U14291 (N_14291,N_13652,N_13970);
and U14292 (N_14292,N_12469,N_12612);
or U14293 (N_14293,N_12386,N_12369);
nand U14294 (N_14294,N_12583,N_12923);
nor U14295 (N_14295,N_13416,N_12312);
or U14296 (N_14296,N_13333,N_12031);
xor U14297 (N_14297,N_12213,N_13857);
xor U14298 (N_14298,N_12482,N_13131);
or U14299 (N_14299,N_13434,N_12565);
and U14300 (N_14300,N_13529,N_12093);
nor U14301 (N_14301,N_12204,N_13577);
nor U14302 (N_14302,N_12220,N_13954);
nand U14303 (N_14303,N_12399,N_13390);
and U14304 (N_14304,N_12675,N_12590);
or U14305 (N_14305,N_13953,N_13959);
nand U14306 (N_14306,N_12977,N_13465);
nand U14307 (N_14307,N_12153,N_12704);
nor U14308 (N_14308,N_13291,N_13873);
xor U14309 (N_14309,N_12795,N_13507);
nand U14310 (N_14310,N_12579,N_13054);
or U14311 (N_14311,N_13438,N_13943);
or U14312 (N_14312,N_13999,N_12715);
and U14313 (N_14313,N_13531,N_13517);
nand U14314 (N_14314,N_12424,N_13763);
nor U14315 (N_14315,N_12752,N_12199);
nor U14316 (N_14316,N_12208,N_13157);
and U14317 (N_14317,N_12169,N_12284);
and U14318 (N_14318,N_13662,N_12718);
and U14319 (N_14319,N_12739,N_13298);
or U14320 (N_14320,N_13033,N_13290);
nand U14321 (N_14321,N_12866,N_12818);
nand U14322 (N_14322,N_13525,N_13702);
and U14323 (N_14323,N_12797,N_13229);
and U14324 (N_14324,N_12738,N_12075);
or U14325 (N_14325,N_13457,N_12928);
and U14326 (N_14326,N_13589,N_13322);
nand U14327 (N_14327,N_13047,N_13252);
nor U14328 (N_14328,N_12388,N_13321);
and U14329 (N_14329,N_13061,N_13440);
nor U14330 (N_14330,N_12997,N_13083);
xnor U14331 (N_14331,N_12480,N_13547);
nor U14332 (N_14332,N_13107,N_13267);
and U14333 (N_14333,N_12038,N_12837);
nand U14334 (N_14334,N_12808,N_13670);
xor U14335 (N_14335,N_12086,N_12604);
nor U14336 (N_14336,N_13072,N_13530);
or U14337 (N_14337,N_13084,N_13142);
nor U14338 (N_14338,N_13124,N_13594);
nand U14339 (N_14339,N_13274,N_13087);
and U14340 (N_14340,N_12931,N_13691);
and U14341 (N_14341,N_13575,N_12813);
or U14342 (N_14342,N_13845,N_13059);
or U14343 (N_14343,N_13729,N_13166);
xnor U14344 (N_14344,N_12520,N_13941);
nand U14345 (N_14345,N_13747,N_13700);
or U14346 (N_14346,N_12536,N_13165);
or U14347 (N_14347,N_13031,N_13838);
nand U14348 (N_14348,N_12555,N_12327);
or U14349 (N_14349,N_12135,N_13494);
xor U14350 (N_14350,N_13632,N_13300);
nor U14351 (N_14351,N_13579,N_12471);
xnor U14352 (N_14352,N_12765,N_13249);
xor U14353 (N_14353,N_12485,N_12310);
xor U14354 (N_14354,N_12641,N_13307);
and U14355 (N_14355,N_12836,N_12695);
or U14356 (N_14356,N_13938,N_12418);
nor U14357 (N_14357,N_12535,N_13069);
xor U14358 (N_14358,N_12224,N_13713);
and U14359 (N_14359,N_13342,N_12619);
or U14360 (N_14360,N_13222,N_12030);
and U14361 (N_14361,N_13836,N_13817);
nand U14362 (N_14362,N_12633,N_12314);
and U14363 (N_14363,N_12854,N_12372);
nor U14364 (N_14364,N_12239,N_13101);
or U14365 (N_14365,N_12568,N_13411);
and U14366 (N_14366,N_12787,N_12782);
and U14367 (N_14367,N_13811,N_12610);
nor U14368 (N_14368,N_12481,N_13215);
xnor U14369 (N_14369,N_12602,N_13692);
nor U14370 (N_14370,N_13789,N_13663);
nand U14371 (N_14371,N_12763,N_12863);
nor U14372 (N_14372,N_12419,N_12724);
or U14373 (N_14373,N_13366,N_12734);
nand U14374 (N_14374,N_12144,N_13800);
and U14375 (N_14375,N_12640,N_13376);
and U14376 (N_14376,N_12733,N_13042);
nand U14377 (N_14377,N_13026,N_13295);
xor U14378 (N_14378,N_12859,N_13377);
xor U14379 (N_14379,N_13456,N_12932);
nor U14380 (N_14380,N_13347,N_12995);
nand U14381 (N_14381,N_12319,N_13289);
nand U14382 (N_14382,N_12954,N_12476);
xnor U14383 (N_14383,N_12420,N_13368);
nand U14384 (N_14384,N_12596,N_12356);
nor U14385 (N_14385,N_13910,N_13253);
or U14386 (N_14386,N_12912,N_12589);
and U14387 (N_14387,N_12552,N_13233);
or U14388 (N_14388,N_13181,N_13907);
nand U14389 (N_14389,N_13002,N_12831);
nand U14390 (N_14390,N_13330,N_12725);
xnor U14391 (N_14391,N_13924,N_12513);
or U14392 (N_14392,N_13472,N_12407);
xor U14393 (N_14393,N_12677,N_13810);
nor U14394 (N_14394,N_13750,N_12779);
nor U14395 (N_14395,N_13179,N_13520);
nor U14396 (N_14396,N_12647,N_12163);
xnor U14397 (N_14397,N_12728,N_12311);
and U14398 (N_14398,N_13212,N_12936);
or U14399 (N_14399,N_13258,N_12699);
nand U14400 (N_14400,N_12102,N_12122);
and U14401 (N_14401,N_13723,N_12203);
and U14402 (N_14402,N_13161,N_12503);
and U14403 (N_14403,N_13032,N_13612);
nor U14404 (N_14404,N_13070,N_13769);
or U14405 (N_14405,N_13045,N_12924);
or U14406 (N_14406,N_12067,N_13133);
and U14407 (N_14407,N_13137,N_13393);
xnor U14408 (N_14408,N_12248,N_13900);
nor U14409 (N_14409,N_13894,N_12712);
or U14410 (N_14410,N_12364,N_12121);
and U14411 (N_14411,N_13415,N_13400);
and U14412 (N_14412,N_12434,N_12283);
or U14413 (N_14413,N_13373,N_13583);
xor U14414 (N_14414,N_12414,N_12406);
nor U14415 (N_14415,N_12573,N_12315);
and U14416 (N_14416,N_12950,N_12975);
nor U14417 (N_14417,N_12452,N_13711);
xor U14418 (N_14418,N_12898,N_13737);
or U14419 (N_14419,N_13353,N_12411);
or U14420 (N_14420,N_12794,N_12099);
nor U14421 (N_14421,N_12745,N_13664);
nand U14422 (N_14422,N_12376,N_13499);
and U14423 (N_14423,N_13801,N_12159);
xor U14424 (N_14424,N_13269,N_13496);
nand U14425 (N_14425,N_12125,N_13629);
nand U14426 (N_14426,N_12527,N_12717);
or U14427 (N_14427,N_13285,N_12280);
and U14428 (N_14428,N_13934,N_13831);
xor U14429 (N_14429,N_13277,N_12097);
nor U14430 (N_14430,N_13464,N_12006);
or U14431 (N_14431,N_13860,N_13288);
or U14432 (N_14432,N_13371,N_13420);
or U14433 (N_14433,N_13765,N_12005);
and U14434 (N_14434,N_12066,N_12956);
and U14435 (N_14435,N_13256,N_13883);
or U14436 (N_14436,N_13809,N_12731);
nor U14437 (N_14437,N_12949,N_12971);
xor U14438 (N_14438,N_12033,N_12723);
xnor U14439 (N_14439,N_13519,N_13016);
nand U14440 (N_14440,N_13827,N_12351);
nand U14441 (N_14441,N_13299,N_12887);
or U14442 (N_14442,N_13304,N_12172);
nand U14443 (N_14443,N_13261,N_12943);
nor U14444 (N_14444,N_13879,N_13593);
nor U14445 (N_14445,N_13610,N_12063);
and U14446 (N_14446,N_13773,N_12553);
nand U14447 (N_14447,N_13551,N_12720);
nor U14448 (N_14448,N_12258,N_12333);
xnor U14449 (N_14449,N_12344,N_13615);
xnor U14450 (N_14450,N_13315,N_13497);
xnor U14451 (N_14451,N_12120,N_12494);
or U14452 (N_14452,N_12247,N_13778);
or U14453 (N_14453,N_13379,N_13932);
xor U14454 (N_14454,N_13962,N_13019);
and U14455 (N_14455,N_12860,N_13147);
or U14456 (N_14456,N_13556,N_13375);
and U14457 (N_14457,N_13787,N_12680);
nor U14458 (N_14458,N_13666,N_13105);
or U14459 (N_14459,N_12804,N_12170);
nor U14460 (N_14460,N_13012,N_12037);
xor U14461 (N_14461,N_12379,N_13425);
nor U14462 (N_14462,N_12358,N_13168);
xnor U14463 (N_14463,N_13292,N_12453);
nor U14464 (N_14464,N_12833,N_13445);
or U14465 (N_14465,N_13196,N_13000);
nor U14466 (N_14466,N_12187,N_12221);
xnor U14467 (N_14467,N_12847,N_12391);
xor U14468 (N_14468,N_13865,N_12353);
nand U14469 (N_14469,N_13429,N_12137);
or U14470 (N_14470,N_13283,N_12811);
and U14471 (N_14471,N_13185,N_12669);
nand U14472 (N_14472,N_12626,N_13917);
nor U14473 (N_14473,N_13768,N_13122);
and U14474 (N_14474,N_12104,N_12231);
or U14475 (N_14475,N_12328,N_12502);
and U14476 (N_14476,N_12986,N_12774);
and U14477 (N_14477,N_12160,N_13985);
or U14478 (N_14478,N_13602,N_12905);
and U14479 (N_14479,N_12927,N_13646);
nand U14480 (N_14480,N_13071,N_12161);
nand U14481 (N_14481,N_12100,N_12652);
or U14482 (N_14482,N_13543,N_13432);
nor U14483 (N_14483,N_13826,N_12028);
nor U14484 (N_14484,N_12759,N_12241);
and U14485 (N_14485,N_13323,N_12291);
xnor U14486 (N_14486,N_13903,N_12422);
nor U14487 (N_14487,N_13571,N_13064);
and U14488 (N_14488,N_13325,N_12409);
nor U14489 (N_14489,N_12068,N_12868);
nand U14490 (N_14490,N_12983,N_12212);
or U14491 (N_14491,N_12994,N_13676);
or U14492 (N_14492,N_13011,N_13973);
nor U14493 (N_14493,N_13078,N_13624);
nor U14494 (N_14494,N_13094,N_12631);
nor U14495 (N_14495,N_12697,N_12665);
or U14496 (N_14496,N_13997,N_13915);
and U14497 (N_14497,N_12771,N_12805);
xor U14498 (N_14498,N_12989,N_12215);
and U14499 (N_14499,N_13536,N_12329);
nor U14500 (N_14500,N_12926,N_12252);
xor U14501 (N_14501,N_13159,N_13423);
xor U14502 (N_14502,N_12784,N_12929);
or U14503 (N_14503,N_12758,N_13348);
nand U14504 (N_14504,N_12683,N_13981);
or U14505 (N_14505,N_13799,N_12276);
xnor U14506 (N_14506,N_12711,N_12263);
nand U14507 (N_14507,N_12968,N_12431);
nand U14508 (N_14508,N_13820,N_12581);
and U14509 (N_14509,N_12269,N_13471);
or U14510 (N_14510,N_13896,N_12045);
nand U14511 (N_14511,N_12916,N_12462);
xor U14512 (N_14512,N_13337,N_12532);
xnor U14513 (N_14513,N_12206,N_12165);
or U14514 (N_14514,N_13093,N_13313);
nand U14515 (N_14515,N_12735,N_12694);
nor U14516 (N_14516,N_12289,N_12057);
xor U14517 (N_14517,N_12448,N_13541);
and U14518 (N_14518,N_13854,N_13552);
and U14519 (N_14519,N_13829,N_13022);
or U14520 (N_14520,N_13005,N_12401);
xor U14521 (N_14521,N_13296,N_12413);
and U14522 (N_14522,N_13027,N_12799);
nand U14523 (N_14523,N_13082,N_13246);
and U14524 (N_14524,N_12235,N_13980);
and U14525 (N_14525,N_13759,N_13479);
or U14526 (N_14526,N_13151,N_13887);
nand U14527 (N_14527,N_13516,N_12948);
and U14528 (N_14528,N_13433,N_13123);
nor U14529 (N_14529,N_13220,N_13459);
or U14530 (N_14530,N_12542,N_12960);
or U14531 (N_14531,N_13839,N_13719);
or U14532 (N_14532,N_12083,N_13484);
nor U14533 (N_14533,N_12504,N_12374);
or U14534 (N_14534,N_13671,N_12512);
or U14535 (N_14535,N_12049,N_12776);
xor U14536 (N_14536,N_12755,N_12039);
or U14537 (N_14537,N_12925,N_13728);
and U14538 (N_14538,N_13399,N_12708);
and U14539 (N_14539,N_12621,N_13235);
nor U14540 (N_14540,N_13782,N_13779);
or U14541 (N_14541,N_13835,N_13443);
and U14542 (N_14542,N_12690,N_12592);
nor U14543 (N_14543,N_13816,N_13925);
nor U14544 (N_14544,N_12060,N_12878);
and U14545 (N_14545,N_12889,N_13260);
nor U14546 (N_14546,N_12339,N_13753);
xnor U14547 (N_14547,N_12479,N_12828);
xor U14548 (N_14548,N_12691,N_13355);
and U14549 (N_14549,N_12838,N_12685);
xor U14550 (N_14550,N_13871,N_13733);
and U14551 (N_14551,N_13512,N_12841);
and U14552 (N_14552,N_12223,N_13866);
or U14553 (N_14553,N_12939,N_13192);
nand U14554 (N_14554,N_12830,N_12564);
and U14555 (N_14555,N_13344,N_12845);
or U14556 (N_14556,N_13986,N_12446);
and U14557 (N_14557,N_12562,N_13644);
nor U14558 (N_14558,N_13041,N_13401);
and U14559 (N_14559,N_13994,N_13562);
xnor U14560 (N_14560,N_13686,N_12242);
or U14561 (N_14561,N_12519,N_13065);
xor U14562 (N_14562,N_12508,N_13156);
or U14563 (N_14563,N_13743,N_13503);
and U14564 (N_14564,N_13067,N_13573);
and U14565 (N_14565,N_13784,N_12015);
nor U14566 (N_14566,N_13730,N_12705);
xor U14567 (N_14567,N_13485,N_13731);
nand U14568 (N_14568,N_13338,N_13030);
xor U14569 (N_14569,N_13326,N_13849);
nor U14570 (N_14570,N_13597,N_12679);
xnor U14571 (N_14571,N_12721,N_13170);
nand U14572 (N_14572,N_13450,N_12488);
or U14573 (N_14573,N_13815,N_12139);
nor U14574 (N_14574,N_13734,N_12112);
nor U14575 (N_14575,N_12017,N_12089);
nor U14576 (N_14576,N_12405,N_13234);
nor U14577 (N_14577,N_12412,N_13491);
or U14578 (N_14578,N_13418,N_12109);
nor U14579 (N_14579,N_13103,N_13395);
xnor U14580 (N_14580,N_13961,N_12158);
and U14581 (N_14581,N_12769,N_12255);
or U14582 (N_14582,N_12064,N_12131);
xnor U14583 (N_14583,N_12016,N_13568);
nand U14584 (N_14584,N_12499,N_13975);
nand U14585 (N_14585,N_13918,N_13830);
nand U14586 (N_14586,N_13618,N_12918);
nand U14587 (N_14587,N_13683,N_13488);
and U14588 (N_14588,N_13718,N_12766);
nor U14589 (N_14589,N_13895,N_12001);
xnor U14590 (N_14590,N_12267,N_13694);
nand U14591 (N_14591,N_12383,N_13679);
xnor U14592 (N_14592,N_12143,N_12457);
or U14593 (N_14593,N_13020,N_13565);
xor U14594 (N_14594,N_13334,N_12189);
or U14595 (N_14595,N_12281,N_12528);
or U14596 (N_14596,N_13638,N_13195);
and U14597 (N_14597,N_12609,N_12871);
nand U14598 (N_14598,N_13651,N_13386);
nor U14599 (N_14599,N_12253,N_12663);
nor U14600 (N_14600,N_13557,N_12644);
and U14601 (N_14601,N_12132,N_12775);
and U14602 (N_14602,N_12341,N_13340);
nand U14603 (N_14603,N_13559,N_13495);
xor U14604 (N_14604,N_13257,N_12261);
or U14605 (N_14605,N_12210,N_12115);
xnor U14606 (N_14606,N_12167,N_12757);
xor U14607 (N_14607,N_12004,N_13876);
nand U14608 (N_14608,N_13720,N_12019);
nor U14609 (N_14609,N_12662,N_13774);
or U14610 (N_14610,N_12129,N_12209);
nand U14611 (N_14611,N_12687,N_13748);
xor U14612 (N_14612,N_13435,N_12029);
nor U14613 (N_14613,N_13587,N_12305);
nand U14614 (N_14614,N_13505,N_12585);
nor U14615 (N_14615,N_13474,N_13138);
nand U14616 (N_14616,N_12870,N_12326);
and U14617 (N_14617,N_12337,N_12700);
or U14618 (N_14618,N_12054,N_13271);
xor U14619 (N_14619,N_13561,N_13172);
and U14620 (N_14620,N_13263,N_12746);
nand U14621 (N_14621,N_13412,N_12639);
nor U14622 (N_14622,N_13546,N_13477);
nand U14623 (N_14623,N_13814,N_12179);
xnor U14624 (N_14624,N_13044,N_12561);
nand U14625 (N_14625,N_13813,N_13878);
nor U14626 (N_14626,N_12108,N_13037);
and U14627 (N_14627,N_13448,N_13141);
or U14628 (N_14628,N_13712,N_13476);
and U14629 (N_14629,N_12384,N_13899);
xor U14630 (N_14630,N_12599,N_12119);
nand U14631 (N_14631,N_12615,N_13626);
nand U14632 (N_14632,N_12380,N_12584);
xnor U14633 (N_14633,N_12888,N_13363);
nand U14634 (N_14634,N_12468,N_13755);
nor U14635 (N_14635,N_13381,N_13705);
and U14636 (N_14636,N_13293,N_12980);
xnor U14637 (N_14637,N_12361,N_12623);
xnor U14638 (N_14638,N_13528,N_13282);
or U14639 (N_14639,N_12540,N_12686);
or U14640 (N_14640,N_12689,N_12027);
or U14641 (N_14641,N_13625,N_13936);
xor U14642 (N_14642,N_12470,N_12603);
and U14643 (N_14643,N_13359,N_13305);
xor U14644 (N_14644,N_13656,N_12781);
and U14645 (N_14645,N_12168,N_12730);
xnor U14646 (N_14646,N_12702,N_13805);
xor U14647 (N_14647,N_12900,N_12654);
or U14648 (N_14648,N_13850,N_13869);
xor U14649 (N_14649,N_12347,N_12014);
nor U14650 (N_14650,N_13921,N_12961);
and U14651 (N_14651,N_13616,N_12858);
nor U14652 (N_14652,N_12842,N_12188);
xnor U14653 (N_14653,N_12331,N_13231);
xor U14654 (N_14654,N_12586,N_13414);
nor U14655 (N_14655,N_13974,N_13600);
or U14656 (N_14656,N_12829,N_12963);
nor U14657 (N_14657,N_13802,N_13343);
nand U14658 (N_14658,N_13068,N_12967);
xnor U14659 (N_14659,N_13939,N_13928);
and U14660 (N_14660,N_13788,N_13757);
nor U14661 (N_14661,N_12657,N_13378);
nand U14662 (N_14662,N_12421,N_13367);
or U14663 (N_14663,N_12439,N_12893);
or U14664 (N_14664,N_13332,N_12272);
nand U14665 (N_14665,N_12249,N_13360);
xnor U14666 (N_14666,N_12959,N_13945);
nand U14667 (N_14667,N_12511,N_13906);
or U14668 (N_14668,N_12627,N_12140);
xor U14669 (N_14669,N_13592,N_13226);
xor U14670 (N_14670,N_12869,N_12744);
nor U14671 (N_14671,N_12077,N_13736);
xnor U14672 (N_14672,N_13199,N_13126);
and U14673 (N_14673,N_13661,N_13875);
nand U14674 (N_14674,N_12792,N_13406);
or U14675 (N_14675,N_12933,N_12638);
xnor U14676 (N_14676,N_12810,N_13162);
and U14677 (N_14677,N_13952,N_13272);
nand U14678 (N_14678,N_13780,N_13806);
and U14679 (N_14679,N_13232,N_13511);
nor U14680 (N_14680,N_13297,N_12403);
or U14681 (N_14681,N_12987,N_12778);
xor U14682 (N_14682,N_13302,N_13560);
or U14683 (N_14683,N_13158,N_12875);
nor U14684 (N_14684,N_12732,N_12901);
and U14685 (N_14685,N_12081,N_12601);
nor U14686 (N_14686,N_13708,N_13427);
nor U14687 (N_14687,N_13112,N_13125);
nor U14688 (N_14688,N_13796,N_12177);
or U14689 (N_14689,N_13870,N_13317);
and U14690 (N_14690,N_13396,N_12320);
or U14691 (N_14691,N_13014,N_12103);
nor U14692 (N_14692,N_12676,N_13038);
and U14693 (N_14693,N_13091,N_13913);
or U14694 (N_14694,N_13758,N_12577);
nand U14695 (N_14695,N_13098,N_12806);
xor U14696 (N_14696,N_12126,N_13957);
and U14697 (N_14697,N_12282,N_12692);
xnor U14698 (N_14698,N_13273,N_13275);
and U14699 (N_14699,N_13888,N_13681);
nor U14700 (N_14700,N_12436,N_12322);
nor U14701 (N_14701,N_12445,N_12996);
nor U14702 (N_14702,N_12902,N_12886);
and U14703 (N_14703,N_13270,N_13207);
or U14704 (N_14704,N_12428,N_13564);
or U14705 (N_14705,N_13678,N_12297);
nand U14706 (N_14706,N_12316,N_12572);
nand U14707 (N_14707,N_12130,N_12138);
nor U14708 (N_14708,N_13598,N_13889);
nor U14709 (N_14709,N_13930,N_13419);
nor U14710 (N_14710,N_12891,N_13178);
or U14711 (N_14711,N_12365,N_13490);
and U14712 (N_14712,N_12265,N_13144);
nand U14713 (N_14713,N_13971,N_12938);
and U14714 (N_14714,N_13620,N_12935);
and U14715 (N_14715,N_13824,N_13793);
nor U14716 (N_14716,N_12178,N_12114);
xnor U14717 (N_14717,N_12085,N_12608);
or U14718 (N_14718,N_13216,N_13964);
nor U14719 (N_14719,N_13764,N_12880);
nand U14720 (N_14720,N_12826,N_12578);
and U14721 (N_14721,N_12537,N_12944);
and U14722 (N_14722,N_13886,N_12012);
and U14723 (N_14723,N_13463,N_13833);
xnor U14724 (N_14724,N_13143,N_13449);
or U14725 (N_14725,N_12801,N_12072);
or U14726 (N_14726,N_13848,N_13680);
nor U14727 (N_14727,N_13905,N_12338);
nor U14728 (N_14728,N_12304,N_13920);
nand U14729 (N_14729,N_12800,N_12171);
or U14730 (N_14730,N_13120,N_13697);
nor U14731 (N_14731,N_12632,N_13077);
and U14732 (N_14732,N_13264,N_12793);
xor U14733 (N_14733,N_12655,N_13902);
xor U14734 (N_14734,N_13336,N_13553);
nand U14735 (N_14735,N_12141,N_12359);
nor U14736 (N_14736,N_13786,N_12155);
and U14737 (N_14737,N_13502,N_13374);
and U14738 (N_14738,N_12127,N_12301);
nor U14739 (N_14739,N_13908,N_12308);
nand U14740 (N_14740,N_13739,N_12490);
nand U14741 (N_14741,N_13023,N_12628);
nand U14742 (N_14742,N_13268,N_12947);
or U14743 (N_14743,N_13239,N_13361);
xor U14744 (N_14744,N_13354,N_12290);
or U14745 (N_14745,N_13346,N_13169);
or U14746 (N_14746,N_12913,N_12343);
and U14747 (N_14747,N_13812,N_13893);
and U14748 (N_14748,N_12237,N_12849);
xnor U14749 (N_14749,N_12368,N_13897);
nand U14750 (N_14750,N_12713,N_13116);
and U14751 (N_14751,N_13111,N_12791);
xor U14752 (N_14752,N_13752,N_13864);
or U14753 (N_14753,N_13710,N_12070);
xnor U14754 (N_14754,N_13230,N_13106);
and U14755 (N_14755,N_13832,N_13521);
or U14756 (N_14756,N_13715,N_13738);
nor U14757 (N_14757,N_12197,N_12884);
xor U14758 (N_14758,N_13461,N_13301);
or U14759 (N_14759,N_13726,N_13218);
xor U14760 (N_14760,N_12591,N_13189);
nand U14761 (N_14761,N_13606,N_12515);
and U14762 (N_14762,N_12497,N_12186);
nor U14763 (N_14763,N_12611,N_12659);
xnor U14764 (N_14764,N_13244,N_12260);
or U14765 (N_14765,N_12449,N_13405);
nand U14766 (N_14766,N_12232,N_13534);
or U14767 (N_14767,N_13544,N_12198);
nor U14768 (N_14768,N_12867,N_12071);
nand U14769 (N_14769,N_12814,N_13706);
and U14770 (N_14770,N_12501,N_12907);
nor U14771 (N_14771,N_12332,N_12266);
xor U14772 (N_14772,N_13130,N_13872);
nand U14773 (N_14773,N_13424,N_12530);
nand U14774 (N_14774,N_13190,N_13933);
or U14775 (N_14775,N_12559,N_12371);
xnor U14776 (N_14776,N_12056,N_12026);
and U14777 (N_14777,N_12701,N_12463);
nor U14778 (N_14778,N_13563,N_12007);
or U14779 (N_14779,N_12385,N_13075);
nand U14780 (N_14780,N_12079,N_12816);
xnor U14781 (N_14781,N_12279,N_12432);
and U14782 (N_14782,N_13732,N_13603);
nand U14783 (N_14783,N_12786,N_12798);
nand U14784 (N_14784,N_13335,N_13060);
and U14785 (N_14785,N_13046,N_13018);
nor U14786 (N_14786,N_12580,N_12966);
nor U14787 (N_14787,N_13250,N_12055);
xnor U14788 (N_14788,N_13636,N_13004);
and U14789 (N_14789,N_13834,N_12442);
or U14790 (N_14790,N_13096,N_12218);
and U14791 (N_14791,N_12423,N_13312);
or U14792 (N_14792,N_12182,N_13874);
xnor U14793 (N_14793,N_13262,N_12534);
or U14794 (N_14794,N_12395,N_13821);
nand U14795 (N_14795,N_12254,N_13372);
nor U14796 (N_14796,N_13766,N_12957);
nand U14797 (N_14797,N_13703,N_13674);
nor U14798 (N_14798,N_13251,N_13891);
or U14799 (N_14799,N_12302,N_13403);
nand U14800 (N_14800,N_13695,N_12563);
and U14801 (N_14801,N_12817,N_13862);
and U14802 (N_14802,N_13136,N_12256);
or U14803 (N_14803,N_13510,N_12117);
nand U14804 (N_14804,N_12176,N_13533);
xor U14805 (N_14805,N_12783,N_13791);
and U14806 (N_14806,N_12000,N_13303);
nand U14807 (N_14807,N_12173,N_13320);
nand U14808 (N_14808,N_12296,N_13241);
xnor U14809 (N_14809,N_13548,N_13248);
xnor U14810 (N_14810,N_12486,N_12620);
xor U14811 (N_14811,N_12524,N_12336);
and U14812 (N_14812,N_13522,N_12360);
xor U14813 (N_14813,N_12618,N_12487);
and U14814 (N_14814,N_12635,N_13224);
nand U14815 (N_14815,N_12616,N_12013);
nand U14816 (N_14816,N_12674,N_13650);
or U14817 (N_14817,N_12355,N_12598);
nor U14818 (N_14818,N_13825,N_13580);
and U14819 (N_14819,N_12090,N_12673);
nand U14820 (N_14820,N_13007,N_13581);
nor U14821 (N_14821,N_13148,N_13140);
xor U14822 (N_14822,N_13642,N_12812);
and U14823 (N_14823,N_12908,N_12370);
and U14824 (N_14824,N_12710,N_13538);
nor U14825 (N_14825,N_12443,N_12557);
and U14826 (N_14826,N_12571,N_12554);
xor U14827 (N_14827,N_13280,N_12325);
xor U14828 (N_14828,N_12594,N_13356);
xnor U14829 (N_14829,N_13890,N_13901);
xor U14830 (N_14830,N_12551,N_13176);
nor U14831 (N_14831,N_12653,N_12484);
and U14832 (N_14832,N_12667,N_12042);
or U14833 (N_14833,N_12903,N_13468);
or U14834 (N_14834,N_13501,N_13949);
nand U14835 (N_14835,N_13588,N_12475);
nand U14836 (N_14836,N_12474,N_13389);
and U14837 (N_14837,N_13595,N_12275);
and U14838 (N_14838,N_12904,N_13227);
nor U14839 (N_14839,N_13649,N_13607);
nand U14840 (N_14840,N_12350,N_12495);
xor U14841 (N_14841,N_13444,N_12473);
and U14842 (N_14842,N_12651,N_12349);
nor U14843 (N_14843,N_13532,N_13118);
xor U14844 (N_14844,N_12637,N_12417);
xor U14845 (N_14845,N_13996,N_13696);
nand U14846 (N_14846,N_12761,N_12593);
nand U14847 (N_14847,N_12523,N_12342);
or U14848 (N_14848,N_12832,N_12550);
nand U14849 (N_14849,N_12661,N_12124);
or U14850 (N_14850,N_13066,N_13714);
nand U14851 (N_14851,N_12278,N_13294);
nand U14852 (N_14852,N_12772,N_13923);
or U14853 (N_14853,N_13840,N_13942);
nor U14854 (N_14854,N_13958,N_12052);
and U14855 (N_14855,N_12546,N_12538);
or U14856 (N_14856,N_12354,N_13640);
nor U14857 (N_14857,N_13035,N_13995);
or U14858 (N_14858,N_13968,N_13240);
xor U14859 (N_14859,N_13611,N_13352);
or U14860 (N_14860,N_13740,N_12190);
nand U14861 (N_14861,N_13527,N_13055);
and U14862 (N_14862,N_12214,N_12751);
nand U14863 (N_14863,N_12952,N_13329);
or U14864 (N_14864,N_13955,N_13578);
xor U14865 (N_14865,N_12998,N_12201);
nand U14866 (N_14866,N_12489,N_13062);
or U14867 (N_14867,N_13947,N_13454);
xnor U14868 (N_14868,N_12299,N_12257);
nor U14869 (N_14869,N_13992,N_13284);
and U14870 (N_14870,N_12003,N_13940);
and U14871 (N_14871,N_12909,N_12953);
xnor U14872 (N_14872,N_13770,N_13225);
and U14873 (N_14873,N_13155,N_12082);
nor U14874 (N_14874,N_13776,N_12531);
xor U14875 (N_14875,N_12650,N_12181);
nand U14876 (N_14876,N_12274,N_13808);
nor U14877 (N_14877,N_12496,N_12357);
or U14878 (N_14878,N_12433,N_12156);
or U14879 (N_14879,N_12251,N_12570);
or U14880 (N_14880,N_13926,N_12770);
or U14881 (N_14881,N_13021,N_12597);
nand U14882 (N_14882,N_13013,N_13537);
nor U14883 (N_14883,N_13086,N_12533);
nand U14884 (N_14884,N_13972,N_12041);
nor U14885 (N_14885,N_13349,N_13675);
nor U14886 (N_14886,N_12582,N_12009);
xnor U14887 (N_14887,N_13467,N_12264);
or U14888 (N_14888,N_13627,N_12509);
or U14889 (N_14889,N_12101,N_13462);
or U14890 (N_14890,N_12681,N_12225);
and U14891 (N_14891,N_13623,N_13637);
xnor U14892 (N_14892,N_12270,N_12606);
xor U14893 (N_14893,N_12574,N_13382);
nand U14894 (N_14894,N_13775,N_13777);
xor U14895 (N_14895,N_13667,N_13191);
and U14896 (N_14896,N_13605,N_12400);
nand U14897 (N_14897,N_13243,N_12195);
xnor U14898 (N_14898,N_13881,N_13394);
xnor U14899 (N_14899,N_12990,N_13036);
nor U14900 (N_14900,N_12796,N_12803);
nor U14901 (N_14901,N_12941,N_12324);
or U14902 (N_14902,N_13339,N_12425);
xnor U14903 (N_14903,N_12053,N_12340);
or U14904 (N_14904,N_13990,N_12147);
xor U14905 (N_14905,N_12753,N_13452);
xnor U14906 (N_14906,N_12992,N_13286);
or U14907 (N_14907,N_12917,N_12625);
and U14908 (N_14908,N_12250,N_13684);
nand U14909 (N_14909,N_13163,N_12377);
or U14910 (N_14910,N_12595,N_12649);
nand U14911 (N_14911,N_13914,N_13567);
and U14912 (N_14912,N_12438,N_12217);
nor U14913 (N_14913,N_12166,N_13745);
or U14914 (N_14914,N_12011,N_12742);
nand U14915 (N_14915,N_12080,N_13643);
and U14916 (N_14916,N_13785,N_12047);
nand U14917 (N_14917,N_12491,N_12465);
nand U14918 (N_14918,N_12865,N_12020);
and U14919 (N_14919,N_12666,N_13076);
and U14920 (N_14920,N_13447,N_13843);
or U14921 (N_14921,N_13509,N_12896);
nor U14922 (N_14922,N_13628,N_13099);
and U14923 (N_14923,N_12345,N_13110);
xor U14924 (N_14924,N_12525,N_13641);
or U14925 (N_14925,N_12846,N_13596);
or U14926 (N_14926,N_12382,N_13946);
nand U14927 (N_14927,N_13279,N_13088);
xor U14928 (N_14928,N_13492,N_12287);
xor U14929 (N_14929,N_12483,N_12467);
or U14930 (N_14930,N_12402,N_12510);
nand U14931 (N_14931,N_13453,N_13402);
xor U14932 (N_14932,N_12897,N_12827);
and U14933 (N_14933,N_13614,N_13572);
or U14934 (N_14934,N_12514,N_13916);
and U14935 (N_14935,N_12749,N_13113);
nor U14936 (N_14936,N_12464,N_12825);
or U14937 (N_14937,N_13119,N_12942);
or U14938 (N_14938,N_13152,N_13073);
nand U14939 (N_14939,N_13281,N_12062);
nand U14940 (N_14940,N_13648,N_12688);
or U14941 (N_14941,N_13880,N_12624);
nand U14942 (N_14942,N_13238,N_12855);
nand U14943 (N_14943,N_13392,N_13388);
or U14944 (N_14944,N_12864,N_13504);
nand U14945 (N_14945,N_13966,N_12092);
xnor U14946 (N_14946,N_13114,N_12862);
or U14947 (N_14947,N_13795,N_13104);
nor U14948 (N_14948,N_12183,N_13351);
nor U14949 (N_14949,N_12288,N_13613);
or U14950 (N_14950,N_12965,N_12461);
nand U14951 (N_14951,N_12760,N_13526);
nor U14952 (N_14952,N_12219,N_13430);
xor U14953 (N_14953,N_12576,N_12059);
nand U14954 (N_14954,N_13460,N_12646);
nand U14955 (N_14955,N_13309,N_13909);
and U14956 (N_14956,N_12773,N_12981);
nor U14957 (N_14957,N_12313,N_13001);
nand U14958 (N_14958,N_12246,N_12736);
xnor U14959 (N_14959,N_13574,N_12874);
and U14960 (N_14960,N_13859,N_12999);
nand U14961 (N_14961,N_12750,N_12873);
nand U14962 (N_14962,N_13108,N_13781);
nand U14963 (N_14963,N_12985,N_13205);
or U14964 (N_14964,N_13668,N_12309);
and U14965 (N_14965,N_12767,N_13672);
xnor U14966 (N_14966,N_12034,N_12820);
xnor U14967 (N_14967,N_12196,N_12478);
nor U14968 (N_14968,N_12707,N_13701);
or U14969 (N_14969,N_13153,N_12754);
nand U14970 (N_14970,N_12600,N_13979);
xor U14971 (N_14971,N_12389,N_12259);
xnor U14972 (N_14972,N_12678,N_13619);
or U14973 (N_14973,N_12088,N_12191);
nand U14974 (N_14974,N_13090,N_13413);
nand U14975 (N_14975,N_12233,N_12136);
nand U14976 (N_14976,N_13688,N_12390);
nor U14977 (N_14977,N_12211,N_12477);
nand U14978 (N_14978,N_12065,N_12930);
nor U14979 (N_14979,N_12207,N_12185);
or U14980 (N_14980,N_13617,N_13558);
xnor U14981 (N_14981,N_13052,N_13139);
xor U14982 (N_14982,N_13797,N_13236);
or U14983 (N_14983,N_13417,N_12098);
xnor U14984 (N_14984,N_12539,N_12492);
nor U14985 (N_14985,N_13653,N_13922);
xnor U14986 (N_14986,N_12298,N_13478);
xnor U14987 (N_14987,N_13287,N_13722);
or U14988 (N_14988,N_13863,N_12444);
and U14989 (N_14989,N_13409,N_12095);
nand U14990 (N_14990,N_12458,N_13048);
nor U14991 (N_14991,N_12002,N_13794);
and U14992 (N_14992,N_13622,N_12617);
nand U14993 (N_14993,N_13129,N_13186);
xor U14994 (N_14994,N_12526,N_13590);
and U14995 (N_14995,N_13633,N_12317);
xor U14996 (N_14996,N_12671,N_12393);
xor U14997 (N_14997,N_13208,N_12856);
nand U14998 (N_14998,N_12074,N_12545);
nand U14999 (N_14999,N_12149,N_12498);
nor U15000 (N_15000,N_13453,N_12947);
or U15001 (N_15001,N_13589,N_12704);
xor U15002 (N_15002,N_12185,N_13237);
nand U15003 (N_15003,N_12004,N_12685);
and U15004 (N_15004,N_12584,N_13894);
nand U15005 (N_15005,N_13375,N_12232);
nor U15006 (N_15006,N_13655,N_12066);
xor U15007 (N_15007,N_12028,N_13873);
or U15008 (N_15008,N_12244,N_12982);
xor U15009 (N_15009,N_12240,N_12487);
or U15010 (N_15010,N_12299,N_12550);
and U15011 (N_15011,N_13763,N_13503);
nand U15012 (N_15012,N_13536,N_12883);
and U15013 (N_15013,N_12878,N_13582);
nand U15014 (N_15014,N_13410,N_13435);
and U15015 (N_15015,N_13791,N_12599);
and U15016 (N_15016,N_13362,N_13625);
and U15017 (N_15017,N_12977,N_12794);
xor U15018 (N_15018,N_12297,N_12551);
xnor U15019 (N_15019,N_12150,N_12962);
or U15020 (N_15020,N_13070,N_12801);
nor U15021 (N_15021,N_13616,N_13966);
xnor U15022 (N_15022,N_12579,N_13789);
and U15023 (N_15023,N_12222,N_13168);
nand U15024 (N_15024,N_12626,N_13119);
or U15025 (N_15025,N_13888,N_13030);
nor U15026 (N_15026,N_12381,N_12329);
nor U15027 (N_15027,N_13730,N_13796);
nor U15028 (N_15028,N_12295,N_12046);
xor U15029 (N_15029,N_12008,N_12128);
nand U15030 (N_15030,N_12228,N_13412);
nand U15031 (N_15031,N_13217,N_12292);
nor U15032 (N_15032,N_13044,N_13094);
nand U15033 (N_15033,N_13592,N_13066);
or U15034 (N_15034,N_13659,N_13691);
nand U15035 (N_15035,N_12540,N_13022);
nand U15036 (N_15036,N_12200,N_12387);
nor U15037 (N_15037,N_13426,N_13718);
or U15038 (N_15038,N_13679,N_12018);
nor U15039 (N_15039,N_12872,N_13455);
xor U15040 (N_15040,N_13835,N_12865);
nand U15041 (N_15041,N_12415,N_12793);
or U15042 (N_15042,N_13634,N_12815);
xor U15043 (N_15043,N_12538,N_12178);
or U15044 (N_15044,N_13279,N_13551);
nor U15045 (N_15045,N_12494,N_12035);
nand U15046 (N_15046,N_12018,N_12946);
and U15047 (N_15047,N_12225,N_12857);
nand U15048 (N_15048,N_13580,N_13142);
or U15049 (N_15049,N_13299,N_13312);
xor U15050 (N_15050,N_12411,N_13243);
nand U15051 (N_15051,N_13927,N_13332);
nand U15052 (N_15052,N_12123,N_12562);
or U15053 (N_15053,N_13623,N_12528);
nor U15054 (N_15054,N_12817,N_12660);
or U15055 (N_15055,N_12041,N_13134);
xnor U15056 (N_15056,N_12793,N_13437);
and U15057 (N_15057,N_13278,N_12653);
nand U15058 (N_15058,N_13461,N_12629);
nor U15059 (N_15059,N_12994,N_13437);
or U15060 (N_15060,N_12394,N_12066);
and U15061 (N_15061,N_12894,N_13983);
and U15062 (N_15062,N_13206,N_13652);
or U15063 (N_15063,N_12006,N_13508);
and U15064 (N_15064,N_12202,N_13889);
nand U15065 (N_15065,N_13979,N_13838);
and U15066 (N_15066,N_13540,N_12732);
nand U15067 (N_15067,N_13474,N_13559);
nand U15068 (N_15068,N_12543,N_13638);
nor U15069 (N_15069,N_13218,N_12918);
or U15070 (N_15070,N_12582,N_13097);
or U15071 (N_15071,N_12036,N_12125);
or U15072 (N_15072,N_13328,N_13781);
nand U15073 (N_15073,N_12835,N_12038);
and U15074 (N_15074,N_12782,N_13167);
or U15075 (N_15075,N_12681,N_13125);
nor U15076 (N_15076,N_12209,N_12259);
or U15077 (N_15077,N_12449,N_12325);
xnor U15078 (N_15078,N_12439,N_13197);
nor U15079 (N_15079,N_13147,N_13875);
nand U15080 (N_15080,N_12237,N_13407);
or U15081 (N_15081,N_13775,N_12499);
nand U15082 (N_15082,N_12752,N_13258);
or U15083 (N_15083,N_12255,N_13399);
xor U15084 (N_15084,N_13547,N_13302);
nor U15085 (N_15085,N_12852,N_12528);
and U15086 (N_15086,N_13866,N_13321);
nand U15087 (N_15087,N_12616,N_13594);
nand U15088 (N_15088,N_12905,N_13559);
xor U15089 (N_15089,N_12792,N_13838);
and U15090 (N_15090,N_13207,N_12409);
nor U15091 (N_15091,N_12924,N_13264);
nor U15092 (N_15092,N_13933,N_13132);
and U15093 (N_15093,N_13146,N_12762);
xnor U15094 (N_15094,N_12320,N_12026);
nor U15095 (N_15095,N_13737,N_13366);
nand U15096 (N_15096,N_12332,N_12440);
and U15097 (N_15097,N_12330,N_13972);
nor U15098 (N_15098,N_13758,N_13401);
or U15099 (N_15099,N_13447,N_12022);
or U15100 (N_15100,N_12531,N_12968);
and U15101 (N_15101,N_12795,N_12798);
xor U15102 (N_15102,N_13179,N_12516);
or U15103 (N_15103,N_12882,N_13481);
nand U15104 (N_15104,N_13824,N_12212);
or U15105 (N_15105,N_12728,N_13066);
xnor U15106 (N_15106,N_13201,N_13907);
or U15107 (N_15107,N_12502,N_13605);
nand U15108 (N_15108,N_13315,N_12588);
nand U15109 (N_15109,N_13808,N_13522);
xnor U15110 (N_15110,N_13650,N_12476);
xor U15111 (N_15111,N_13239,N_13100);
nor U15112 (N_15112,N_13450,N_12346);
xnor U15113 (N_15113,N_13437,N_13875);
xnor U15114 (N_15114,N_12036,N_13359);
and U15115 (N_15115,N_12173,N_12123);
xor U15116 (N_15116,N_12922,N_12106);
nor U15117 (N_15117,N_13815,N_12808);
and U15118 (N_15118,N_13468,N_13116);
and U15119 (N_15119,N_13908,N_13313);
xor U15120 (N_15120,N_13563,N_12712);
nor U15121 (N_15121,N_13354,N_12982);
nor U15122 (N_15122,N_13160,N_12734);
or U15123 (N_15123,N_12813,N_12030);
nand U15124 (N_15124,N_12666,N_13436);
nand U15125 (N_15125,N_12826,N_12719);
nor U15126 (N_15126,N_12199,N_13379);
and U15127 (N_15127,N_12328,N_13982);
nor U15128 (N_15128,N_13932,N_13159);
and U15129 (N_15129,N_13897,N_12288);
nor U15130 (N_15130,N_12095,N_12204);
nand U15131 (N_15131,N_13286,N_13435);
xor U15132 (N_15132,N_12706,N_12918);
nor U15133 (N_15133,N_13313,N_13575);
or U15134 (N_15134,N_12642,N_12519);
nor U15135 (N_15135,N_12946,N_12145);
nand U15136 (N_15136,N_12469,N_12373);
or U15137 (N_15137,N_12756,N_12705);
xnor U15138 (N_15138,N_12112,N_13311);
xnor U15139 (N_15139,N_12463,N_12357);
xor U15140 (N_15140,N_13646,N_13380);
xor U15141 (N_15141,N_12696,N_13435);
nand U15142 (N_15142,N_12336,N_13022);
or U15143 (N_15143,N_12354,N_13427);
or U15144 (N_15144,N_13886,N_13333);
nand U15145 (N_15145,N_12711,N_12957);
nor U15146 (N_15146,N_12346,N_12554);
nand U15147 (N_15147,N_13867,N_13090);
nand U15148 (N_15148,N_12604,N_13444);
xor U15149 (N_15149,N_13664,N_12228);
or U15150 (N_15150,N_12095,N_13319);
or U15151 (N_15151,N_13115,N_12195);
xor U15152 (N_15152,N_12561,N_12328);
nor U15153 (N_15153,N_12302,N_12508);
xnor U15154 (N_15154,N_12259,N_12757);
xor U15155 (N_15155,N_13356,N_13537);
xor U15156 (N_15156,N_13947,N_12874);
and U15157 (N_15157,N_13830,N_13420);
nor U15158 (N_15158,N_13693,N_12191);
or U15159 (N_15159,N_12751,N_13211);
nor U15160 (N_15160,N_13297,N_13146);
xor U15161 (N_15161,N_13920,N_13310);
nor U15162 (N_15162,N_12608,N_13382);
xor U15163 (N_15163,N_12703,N_12062);
nand U15164 (N_15164,N_12764,N_12495);
xnor U15165 (N_15165,N_12634,N_12590);
or U15166 (N_15166,N_13492,N_13541);
or U15167 (N_15167,N_12889,N_13962);
and U15168 (N_15168,N_13358,N_12200);
nand U15169 (N_15169,N_13517,N_13205);
and U15170 (N_15170,N_13337,N_12739);
nor U15171 (N_15171,N_13615,N_12587);
and U15172 (N_15172,N_13058,N_12496);
or U15173 (N_15173,N_13933,N_12043);
nand U15174 (N_15174,N_13244,N_13480);
and U15175 (N_15175,N_13227,N_12979);
nor U15176 (N_15176,N_12926,N_13365);
xor U15177 (N_15177,N_12784,N_12945);
xor U15178 (N_15178,N_13881,N_13446);
or U15179 (N_15179,N_12393,N_12268);
or U15180 (N_15180,N_13710,N_12282);
or U15181 (N_15181,N_12692,N_13005);
nor U15182 (N_15182,N_12151,N_13790);
or U15183 (N_15183,N_12315,N_13689);
nor U15184 (N_15184,N_12222,N_13543);
or U15185 (N_15185,N_13548,N_12093);
xor U15186 (N_15186,N_12253,N_12601);
nand U15187 (N_15187,N_12027,N_12269);
and U15188 (N_15188,N_12169,N_13756);
or U15189 (N_15189,N_12280,N_12568);
xor U15190 (N_15190,N_12843,N_13143);
xnor U15191 (N_15191,N_12828,N_13189);
and U15192 (N_15192,N_13300,N_12362);
nand U15193 (N_15193,N_13039,N_12592);
and U15194 (N_15194,N_13122,N_12715);
or U15195 (N_15195,N_12099,N_13537);
nor U15196 (N_15196,N_13922,N_13985);
nor U15197 (N_15197,N_13999,N_12865);
or U15198 (N_15198,N_12392,N_12331);
nand U15199 (N_15199,N_13264,N_13964);
xnor U15200 (N_15200,N_13047,N_13585);
nor U15201 (N_15201,N_12617,N_12277);
nor U15202 (N_15202,N_13231,N_12801);
and U15203 (N_15203,N_12176,N_13938);
nand U15204 (N_15204,N_12330,N_13698);
or U15205 (N_15205,N_12072,N_13763);
nand U15206 (N_15206,N_13386,N_12584);
nand U15207 (N_15207,N_12720,N_13518);
or U15208 (N_15208,N_13533,N_13941);
nand U15209 (N_15209,N_12004,N_13218);
nor U15210 (N_15210,N_13649,N_12480);
nor U15211 (N_15211,N_13022,N_12253);
or U15212 (N_15212,N_12208,N_13709);
xnor U15213 (N_15213,N_12042,N_12212);
xnor U15214 (N_15214,N_13884,N_12970);
xor U15215 (N_15215,N_12886,N_13920);
or U15216 (N_15216,N_13382,N_13109);
nor U15217 (N_15217,N_12813,N_12501);
or U15218 (N_15218,N_12093,N_13011);
xor U15219 (N_15219,N_12417,N_13093);
and U15220 (N_15220,N_12876,N_12691);
xnor U15221 (N_15221,N_12401,N_12606);
nand U15222 (N_15222,N_12947,N_13173);
nand U15223 (N_15223,N_12512,N_12944);
or U15224 (N_15224,N_13161,N_12594);
nor U15225 (N_15225,N_13971,N_13099);
nand U15226 (N_15226,N_13637,N_12365);
or U15227 (N_15227,N_12925,N_12504);
and U15228 (N_15228,N_12573,N_13437);
nand U15229 (N_15229,N_12271,N_13823);
nor U15230 (N_15230,N_12489,N_12943);
nor U15231 (N_15231,N_12449,N_13051);
nor U15232 (N_15232,N_13390,N_12828);
xnor U15233 (N_15233,N_13608,N_13523);
nor U15234 (N_15234,N_12776,N_13608);
or U15235 (N_15235,N_12033,N_12138);
or U15236 (N_15236,N_12164,N_12692);
nor U15237 (N_15237,N_12207,N_12151);
nand U15238 (N_15238,N_13811,N_12048);
or U15239 (N_15239,N_13196,N_13060);
or U15240 (N_15240,N_12636,N_13666);
xor U15241 (N_15241,N_13265,N_12460);
nand U15242 (N_15242,N_13892,N_13413);
nand U15243 (N_15243,N_12283,N_12803);
nor U15244 (N_15244,N_13270,N_12237);
or U15245 (N_15245,N_13881,N_13121);
xnor U15246 (N_15246,N_12564,N_13926);
nor U15247 (N_15247,N_13027,N_12367);
nor U15248 (N_15248,N_12086,N_12760);
or U15249 (N_15249,N_12889,N_12974);
nand U15250 (N_15250,N_13683,N_12066);
and U15251 (N_15251,N_13717,N_12837);
xor U15252 (N_15252,N_13319,N_12404);
or U15253 (N_15253,N_12337,N_12212);
xor U15254 (N_15254,N_13848,N_12769);
xor U15255 (N_15255,N_12812,N_13099);
xor U15256 (N_15256,N_13316,N_13840);
and U15257 (N_15257,N_13375,N_12977);
nor U15258 (N_15258,N_12676,N_13789);
nor U15259 (N_15259,N_13624,N_12647);
or U15260 (N_15260,N_13450,N_13271);
nor U15261 (N_15261,N_13205,N_13431);
and U15262 (N_15262,N_12464,N_12789);
nor U15263 (N_15263,N_13137,N_12237);
or U15264 (N_15264,N_13713,N_13131);
xnor U15265 (N_15265,N_12713,N_13145);
nand U15266 (N_15266,N_12112,N_13011);
and U15267 (N_15267,N_13776,N_13829);
and U15268 (N_15268,N_13405,N_13677);
xor U15269 (N_15269,N_13131,N_13938);
xnor U15270 (N_15270,N_12760,N_12454);
nand U15271 (N_15271,N_13091,N_13430);
and U15272 (N_15272,N_13689,N_12633);
xnor U15273 (N_15273,N_13956,N_12778);
and U15274 (N_15274,N_13906,N_13172);
xnor U15275 (N_15275,N_12274,N_13849);
and U15276 (N_15276,N_12022,N_12090);
nor U15277 (N_15277,N_13533,N_12564);
nand U15278 (N_15278,N_12258,N_12463);
xnor U15279 (N_15279,N_13255,N_13610);
nor U15280 (N_15280,N_13670,N_12709);
nor U15281 (N_15281,N_13843,N_13803);
or U15282 (N_15282,N_12500,N_13555);
and U15283 (N_15283,N_12383,N_12886);
and U15284 (N_15284,N_13851,N_13881);
or U15285 (N_15285,N_12556,N_12941);
xor U15286 (N_15286,N_13716,N_12701);
and U15287 (N_15287,N_13279,N_13726);
and U15288 (N_15288,N_13974,N_12902);
nor U15289 (N_15289,N_13077,N_13308);
nand U15290 (N_15290,N_12039,N_13253);
nor U15291 (N_15291,N_12629,N_13220);
or U15292 (N_15292,N_12628,N_13189);
and U15293 (N_15293,N_12172,N_13192);
and U15294 (N_15294,N_12947,N_12695);
nor U15295 (N_15295,N_13337,N_13189);
nand U15296 (N_15296,N_12768,N_13913);
nor U15297 (N_15297,N_12203,N_12429);
nand U15298 (N_15298,N_12283,N_12576);
and U15299 (N_15299,N_13588,N_13294);
xnor U15300 (N_15300,N_13903,N_13077);
nor U15301 (N_15301,N_12938,N_13769);
nand U15302 (N_15302,N_12819,N_13441);
or U15303 (N_15303,N_13132,N_13644);
and U15304 (N_15304,N_12291,N_12751);
or U15305 (N_15305,N_12450,N_13704);
and U15306 (N_15306,N_12357,N_12299);
or U15307 (N_15307,N_13733,N_12461);
nand U15308 (N_15308,N_12347,N_13177);
nand U15309 (N_15309,N_12003,N_13192);
xnor U15310 (N_15310,N_12573,N_12555);
xor U15311 (N_15311,N_12481,N_13736);
and U15312 (N_15312,N_13595,N_12199);
nand U15313 (N_15313,N_13220,N_13175);
xnor U15314 (N_15314,N_13640,N_12737);
xor U15315 (N_15315,N_12908,N_12398);
nand U15316 (N_15316,N_12400,N_13940);
or U15317 (N_15317,N_12330,N_12441);
nor U15318 (N_15318,N_13259,N_12713);
nor U15319 (N_15319,N_12808,N_12158);
and U15320 (N_15320,N_13218,N_13716);
or U15321 (N_15321,N_12830,N_12471);
or U15322 (N_15322,N_12268,N_12765);
nor U15323 (N_15323,N_12031,N_12599);
and U15324 (N_15324,N_12045,N_13836);
or U15325 (N_15325,N_12083,N_12877);
nor U15326 (N_15326,N_13805,N_12035);
and U15327 (N_15327,N_13762,N_12662);
xnor U15328 (N_15328,N_13098,N_12506);
or U15329 (N_15329,N_12110,N_13855);
and U15330 (N_15330,N_13665,N_12363);
nor U15331 (N_15331,N_12592,N_13674);
nand U15332 (N_15332,N_12248,N_12384);
and U15333 (N_15333,N_13821,N_13229);
xor U15334 (N_15334,N_12211,N_13894);
xnor U15335 (N_15335,N_12008,N_13078);
nand U15336 (N_15336,N_13251,N_12192);
nand U15337 (N_15337,N_12924,N_13433);
xnor U15338 (N_15338,N_12294,N_13599);
and U15339 (N_15339,N_13937,N_12539);
or U15340 (N_15340,N_12054,N_12665);
xor U15341 (N_15341,N_13920,N_12247);
or U15342 (N_15342,N_12104,N_12207);
or U15343 (N_15343,N_13080,N_13837);
nand U15344 (N_15344,N_12705,N_12452);
or U15345 (N_15345,N_13734,N_12568);
and U15346 (N_15346,N_13470,N_12900);
nor U15347 (N_15347,N_12498,N_13523);
nor U15348 (N_15348,N_13844,N_12412);
or U15349 (N_15349,N_12163,N_12405);
xnor U15350 (N_15350,N_13102,N_13545);
nor U15351 (N_15351,N_13305,N_13318);
or U15352 (N_15352,N_12027,N_13137);
nor U15353 (N_15353,N_13460,N_13651);
or U15354 (N_15354,N_13163,N_13501);
and U15355 (N_15355,N_13320,N_13967);
nor U15356 (N_15356,N_12542,N_12803);
nand U15357 (N_15357,N_12807,N_13045);
and U15358 (N_15358,N_13165,N_12826);
or U15359 (N_15359,N_13795,N_13887);
xnor U15360 (N_15360,N_13309,N_13333);
xnor U15361 (N_15361,N_12325,N_13870);
xor U15362 (N_15362,N_12140,N_12853);
nand U15363 (N_15363,N_12796,N_12687);
nand U15364 (N_15364,N_12947,N_13447);
xnor U15365 (N_15365,N_12299,N_13770);
xnor U15366 (N_15366,N_13944,N_12588);
nor U15367 (N_15367,N_13559,N_13231);
xor U15368 (N_15368,N_13619,N_12793);
xor U15369 (N_15369,N_12075,N_12874);
nand U15370 (N_15370,N_13285,N_12582);
nand U15371 (N_15371,N_12312,N_13523);
nor U15372 (N_15372,N_13148,N_12811);
or U15373 (N_15373,N_13564,N_12288);
xor U15374 (N_15374,N_12721,N_12263);
nor U15375 (N_15375,N_13897,N_12222);
xor U15376 (N_15376,N_13264,N_12499);
or U15377 (N_15377,N_12080,N_13668);
xnor U15378 (N_15378,N_12805,N_12341);
and U15379 (N_15379,N_12658,N_12089);
xnor U15380 (N_15380,N_13174,N_12096);
or U15381 (N_15381,N_12885,N_13838);
and U15382 (N_15382,N_13390,N_13967);
nor U15383 (N_15383,N_12123,N_12197);
or U15384 (N_15384,N_13669,N_12687);
nand U15385 (N_15385,N_13624,N_13959);
nor U15386 (N_15386,N_12089,N_13008);
nand U15387 (N_15387,N_12895,N_12484);
or U15388 (N_15388,N_12225,N_13343);
nor U15389 (N_15389,N_13678,N_13582);
and U15390 (N_15390,N_13189,N_13993);
xnor U15391 (N_15391,N_12471,N_13392);
xnor U15392 (N_15392,N_13678,N_13390);
and U15393 (N_15393,N_12540,N_13734);
nor U15394 (N_15394,N_13591,N_12726);
xnor U15395 (N_15395,N_13123,N_13521);
or U15396 (N_15396,N_13961,N_13642);
or U15397 (N_15397,N_12665,N_12260);
or U15398 (N_15398,N_12959,N_13195);
xor U15399 (N_15399,N_13471,N_13599);
nand U15400 (N_15400,N_13688,N_13845);
nand U15401 (N_15401,N_13011,N_13024);
or U15402 (N_15402,N_12492,N_13450);
nand U15403 (N_15403,N_12599,N_12267);
nor U15404 (N_15404,N_13174,N_13413);
nor U15405 (N_15405,N_12637,N_13804);
nand U15406 (N_15406,N_13045,N_12822);
nor U15407 (N_15407,N_12831,N_13590);
and U15408 (N_15408,N_12986,N_13690);
nand U15409 (N_15409,N_12794,N_12168);
nor U15410 (N_15410,N_12341,N_13184);
or U15411 (N_15411,N_13033,N_13776);
nor U15412 (N_15412,N_13445,N_13149);
xnor U15413 (N_15413,N_12283,N_12059);
nand U15414 (N_15414,N_13160,N_13255);
and U15415 (N_15415,N_12146,N_13113);
and U15416 (N_15416,N_13908,N_12108);
xnor U15417 (N_15417,N_13100,N_12471);
nor U15418 (N_15418,N_12690,N_13115);
nor U15419 (N_15419,N_13057,N_13544);
and U15420 (N_15420,N_12391,N_13631);
xnor U15421 (N_15421,N_12329,N_13910);
xnor U15422 (N_15422,N_12692,N_13172);
nand U15423 (N_15423,N_12968,N_13463);
or U15424 (N_15424,N_13756,N_12927);
xor U15425 (N_15425,N_12594,N_12025);
or U15426 (N_15426,N_13548,N_12770);
xor U15427 (N_15427,N_13000,N_13856);
and U15428 (N_15428,N_12741,N_12676);
nand U15429 (N_15429,N_12854,N_12022);
nor U15430 (N_15430,N_13045,N_13956);
or U15431 (N_15431,N_12790,N_12737);
or U15432 (N_15432,N_13727,N_12310);
or U15433 (N_15433,N_13965,N_13605);
nand U15434 (N_15434,N_13696,N_13512);
nand U15435 (N_15435,N_12767,N_13123);
or U15436 (N_15436,N_12435,N_13124);
nor U15437 (N_15437,N_13815,N_13900);
nor U15438 (N_15438,N_12792,N_12781);
nor U15439 (N_15439,N_12856,N_13952);
xor U15440 (N_15440,N_13624,N_13375);
xnor U15441 (N_15441,N_13933,N_12682);
or U15442 (N_15442,N_12230,N_13886);
or U15443 (N_15443,N_12987,N_13684);
and U15444 (N_15444,N_13639,N_13119);
or U15445 (N_15445,N_12374,N_13141);
and U15446 (N_15446,N_12714,N_13550);
or U15447 (N_15447,N_13783,N_12767);
nand U15448 (N_15448,N_12830,N_13308);
and U15449 (N_15449,N_13160,N_13724);
nand U15450 (N_15450,N_13698,N_13233);
xnor U15451 (N_15451,N_13957,N_12753);
xor U15452 (N_15452,N_12070,N_13358);
xnor U15453 (N_15453,N_13669,N_13437);
nand U15454 (N_15454,N_13613,N_12629);
xor U15455 (N_15455,N_13069,N_13048);
or U15456 (N_15456,N_12787,N_12713);
nand U15457 (N_15457,N_13405,N_13069);
or U15458 (N_15458,N_12759,N_13544);
and U15459 (N_15459,N_13276,N_12361);
nand U15460 (N_15460,N_13277,N_13537);
and U15461 (N_15461,N_12825,N_12419);
nor U15462 (N_15462,N_12366,N_12680);
and U15463 (N_15463,N_13361,N_12273);
nand U15464 (N_15464,N_13192,N_13594);
xnor U15465 (N_15465,N_13632,N_12496);
xnor U15466 (N_15466,N_13316,N_13387);
nor U15467 (N_15467,N_13043,N_13459);
and U15468 (N_15468,N_13071,N_13249);
xnor U15469 (N_15469,N_13288,N_13274);
or U15470 (N_15470,N_13950,N_13954);
or U15471 (N_15471,N_13136,N_13396);
or U15472 (N_15472,N_12256,N_13875);
nand U15473 (N_15473,N_12965,N_12417);
nor U15474 (N_15474,N_13119,N_12130);
or U15475 (N_15475,N_13713,N_13218);
nand U15476 (N_15476,N_13748,N_12920);
nor U15477 (N_15477,N_12318,N_12182);
or U15478 (N_15478,N_12803,N_12134);
and U15479 (N_15479,N_13456,N_12173);
and U15480 (N_15480,N_12080,N_12141);
xor U15481 (N_15481,N_12605,N_12257);
or U15482 (N_15482,N_12701,N_12970);
or U15483 (N_15483,N_12369,N_12156);
nor U15484 (N_15484,N_13278,N_13542);
nand U15485 (N_15485,N_12395,N_12907);
or U15486 (N_15486,N_13661,N_13726);
and U15487 (N_15487,N_13843,N_13321);
or U15488 (N_15488,N_13135,N_13346);
and U15489 (N_15489,N_13547,N_13608);
xor U15490 (N_15490,N_12805,N_13522);
nand U15491 (N_15491,N_13078,N_13901);
xor U15492 (N_15492,N_12241,N_12451);
nor U15493 (N_15493,N_12982,N_12314);
and U15494 (N_15494,N_13557,N_13207);
and U15495 (N_15495,N_13585,N_12135);
nor U15496 (N_15496,N_12693,N_12077);
xor U15497 (N_15497,N_13828,N_13841);
nand U15498 (N_15498,N_13655,N_13667);
and U15499 (N_15499,N_12299,N_13196);
nor U15500 (N_15500,N_12327,N_13578);
nand U15501 (N_15501,N_13360,N_13992);
nor U15502 (N_15502,N_13601,N_13457);
or U15503 (N_15503,N_13610,N_12903);
nand U15504 (N_15504,N_13220,N_13456);
nor U15505 (N_15505,N_12428,N_12812);
nor U15506 (N_15506,N_13919,N_12316);
xor U15507 (N_15507,N_12353,N_12522);
nor U15508 (N_15508,N_13160,N_13708);
nor U15509 (N_15509,N_13169,N_13368);
or U15510 (N_15510,N_12530,N_12322);
or U15511 (N_15511,N_12359,N_12319);
nor U15512 (N_15512,N_12028,N_12851);
and U15513 (N_15513,N_13861,N_12530);
and U15514 (N_15514,N_13537,N_12582);
and U15515 (N_15515,N_12053,N_13562);
xor U15516 (N_15516,N_12042,N_13322);
nand U15517 (N_15517,N_12936,N_13545);
nand U15518 (N_15518,N_12804,N_13770);
or U15519 (N_15519,N_12017,N_13201);
xnor U15520 (N_15520,N_13311,N_12296);
nor U15521 (N_15521,N_13252,N_13083);
xnor U15522 (N_15522,N_12605,N_13187);
and U15523 (N_15523,N_13460,N_13821);
nand U15524 (N_15524,N_12209,N_13494);
or U15525 (N_15525,N_12197,N_13516);
xor U15526 (N_15526,N_13098,N_12374);
xor U15527 (N_15527,N_13142,N_12913);
and U15528 (N_15528,N_12981,N_13127);
xnor U15529 (N_15529,N_12257,N_13688);
xnor U15530 (N_15530,N_12634,N_13762);
nand U15531 (N_15531,N_12491,N_12262);
nand U15532 (N_15532,N_12062,N_12747);
xor U15533 (N_15533,N_13241,N_12108);
nand U15534 (N_15534,N_12119,N_13024);
or U15535 (N_15535,N_12966,N_12786);
or U15536 (N_15536,N_12496,N_13648);
or U15537 (N_15537,N_12195,N_12608);
and U15538 (N_15538,N_12028,N_13130);
nand U15539 (N_15539,N_13988,N_12132);
nor U15540 (N_15540,N_12034,N_12975);
and U15541 (N_15541,N_12515,N_13279);
nor U15542 (N_15542,N_13674,N_13882);
and U15543 (N_15543,N_13504,N_13640);
nand U15544 (N_15544,N_12125,N_12899);
nor U15545 (N_15545,N_13988,N_12894);
xnor U15546 (N_15546,N_12279,N_13623);
and U15547 (N_15547,N_13949,N_12227);
or U15548 (N_15548,N_12539,N_12377);
or U15549 (N_15549,N_12553,N_12665);
or U15550 (N_15550,N_12203,N_13814);
and U15551 (N_15551,N_12522,N_13395);
xor U15552 (N_15552,N_13181,N_13723);
or U15553 (N_15553,N_13785,N_13067);
or U15554 (N_15554,N_13697,N_13611);
xnor U15555 (N_15555,N_12992,N_12386);
and U15556 (N_15556,N_13532,N_13912);
and U15557 (N_15557,N_12884,N_12965);
nand U15558 (N_15558,N_13121,N_13265);
or U15559 (N_15559,N_12186,N_13070);
or U15560 (N_15560,N_12669,N_12651);
nand U15561 (N_15561,N_12865,N_12915);
xor U15562 (N_15562,N_13297,N_12747);
and U15563 (N_15563,N_12834,N_12084);
and U15564 (N_15564,N_12216,N_12465);
nor U15565 (N_15565,N_12761,N_13769);
nor U15566 (N_15566,N_12271,N_13272);
nor U15567 (N_15567,N_13951,N_12333);
nand U15568 (N_15568,N_13696,N_13725);
and U15569 (N_15569,N_12044,N_13761);
and U15570 (N_15570,N_12585,N_13735);
nor U15571 (N_15571,N_13608,N_13306);
and U15572 (N_15572,N_12377,N_13680);
nand U15573 (N_15573,N_12098,N_13109);
or U15574 (N_15574,N_13925,N_13160);
xor U15575 (N_15575,N_12143,N_12232);
or U15576 (N_15576,N_12574,N_13417);
nand U15577 (N_15577,N_12208,N_13266);
nand U15578 (N_15578,N_13760,N_12621);
nor U15579 (N_15579,N_12192,N_12952);
and U15580 (N_15580,N_13683,N_12946);
and U15581 (N_15581,N_13412,N_13518);
and U15582 (N_15582,N_13031,N_12319);
or U15583 (N_15583,N_12634,N_13518);
or U15584 (N_15584,N_13742,N_13587);
nor U15585 (N_15585,N_13047,N_13136);
and U15586 (N_15586,N_13019,N_13878);
nand U15587 (N_15587,N_13984,N_12141);
or U15588 (N_15588,N_13861,N_13563);
nor U15589 (N_15589,N_13968,N_13429);
or U15590 (N_15590,N_12168,N_12135);
nor U15591 (N_15591,N_12618,N_13459);
nor U15592 (N_15592,N_13274,N_12350);
or U15593 (N_15593,N_12514,N_12785);
or U15594 (N_15594,N_13631,N_13251);
nand U15595 (N_15595,N_12829,N_12488);
and U15596 (N_15596,N_12832,N_12496);
and U15597 (N_15597,N_12059,N_13499);
nor U15598 (N_15598,N_13424,N_12525);
nand U15599 (N_15599,N_13957,N_13627);
and U15600 (N_15600,N_12699,N_12582);
or U15601 (N_15601,N_13698,N_13315);
xnor U15602 (N_15602,N_13024,N_13276);
nor U15603 (N_15603,N_12770,N_12811);
nor U15604 (N_15604,N_12193,N_13465);
xnor U15605 (N_15605,N_12562,N_12224);
nand U15606 (N_15606,N_12180,N_13209);
xnor U15607 (N_15607,N_13076,N_13097);
or U15608 (N_15608,N_12362,N_12440);
and U15609 (N_15609,N_12160,N_12866);
xnor U15610 (N_15610,N_12919,N_12131);
or U15611 (N_15611,N_12485,N_13707);
nor U15612 (N_15612,N_13057,N_13050);
nor U15613 (N_15613,N_12793,N_12432);
or U15614 (N_15614,N_12664,N_13224);
or U15615 (N_15615,N_12831,N_13835);
and U15616 (N_15616,N_13560,N_12244);
nand U15617 (N_15617,N_12699,N_12143);
and U15618 (N_15618,N_13890,N_12625);
xnor U15619 (N_15619,N_12774,N_13134);
nand U15620 (N_15620,N_13163,N_12470);
and U15621 (N_15621,N_13356,N_12342);
nor U15622 (N_15622,N_12444,N_12269);
and U15623 (N_15623,N_12207,N_13501);
and U15624 (N_15624,N_13341,N_12557);
or U15625 (N_15625,N_12030,N_12697);
or U15626 (N_15626,N_12032,N_13736);
xnor U15627 (N_15627,N_13746,N_12046);
xnor U15628 (N_15628,N_12581,N_13704);
xor U15629 (N_15629,N_13827,N_12787);
nor U15630 (N_15630,N_12876,N_13663);
and U15631 (N_15631,N_13871,N_12816);
nor U15632 (N_15632,N_13136,N_13254);
nand U15633 (N_15633,N_13567,N_13811);
or U15634 (N_15634,N_13425,N_12316);
nand U15635 (N_15635,N_12791,N_13270);
and U15636 (N_15636,N_13644,N_12534);
or U15637 (N_15637,N_13249,N_13000);
and U15638 (N_15638,N_13565,N_12742);
nand U15639 (N_15639,N_13282,N_12832);
or U15640 (N_15640,N_13938,N_12168);
or U15641 (N_15641,N_12540,N_12374);
nor U15642 (N_15642,N_13670,N_13866);
and U15643 (N_15643,N_12786,N_12124);
nor U15644 (N_15644,N_13977,N_13927);
or U15645 (N_15645,N_12403,N_13578);
xnor U15646 (N_15646,N_12488,N_13675);
xnor U15647 (N_15647,N_13120,N_12807);
xnor U15648 (N_15648,N_13995,N_13715);
nor U15649 (N_15649,N_13536,N_13725);
xor U15650 (N_15650,N_12285,N_13486);
xnor U15651 (N_15651,N_13512,N_12284);
nor U15652 (N_15652,N_13788,N_13954);
xor U15653 (N_15653,N_12311,N_12478);
or U15654 (N_15654,N_12756,N_12944);
nor U15655 (N_15655,N_13604,N_13091);
nor U15656 (N_15656,N_12703,N_12584);
nor U15657 (N_15657,N_13651,N_12440);
and U15658 (N_15658,N_13685,N_12364);
or U15659 (N_15659,N_12103,N_13231);
or U15660 (N_15660,N_12708,N_13557);
and U15661 (N_15661,N_13158,N_13634);
and U15662 (N_15662,N_12674,N_13160);
xnor U15663 (N_15663,N_13812,N_13561);
nor U15664 (N_15664,N_13339,N_13802);
nor U15665 (N_15665,N_12848,N_12010);
nand U15666 (N_15666,N_12088,N_13789);
xnor U15667 (N_15667,N_13176,N_12976);
or U15668 (N_15668,N_12902,N_13144);
nand U15669 (N_15669,N_13020,N_12233);
xnor U15670 (N_15670,N_13814,N_13566);
nand U15671 (N_15671,N_13114,N_13941);
nand U15672 (N_15672,N_12748,N_12319);
or U15673 (N_15673,N_13664,N_13338);
and U15674 (N_15674,N_12692,N_13148);
or U15675 (N_15675,N_12392,N_13478);
and U15676 (N_15676,N_12773,N_13266);
nand U15677 (N_15677,N_12863,N_12245);
or U15678 (N_15678,N_13570,N_12758);
xnor U15679 (N_15679,N_13343,N_12053);
and U15680 (N_15680,N_12821,N_12183);
or U15681 (N_15681,N_12223,N_12789);
nand U15682 (N_15682,N_12410,N_13269);
or U15683 (N_15683,N_12272,N_12095);
nand U15684 (N_15684,N_13519,N_13438);
xor U15685 (N_15685,N_13402,N_12629);
and U15686 (N_15686,N_13810,N_13663);
nor U15687 (N_15687,N_12490,N_13991);
and U15688 (N_15688,N_12061,N_13876);
and U15689 (N_15689,N_13283,N_13610);
xor U15690 (N_15690,N_12658,N_12475);
or U15691 (N_15691,N_12978,N_12439);
nor U15692 (N_15692,N_13883,N_12736);
and U15693 (N_15693,N_13208,N_12062);
xor U15694 (N_15694,N_12203,N_13509);
nand U15695 (N_15695,N_12618,N_13812);
xnor U15696 (N_15696,N_12214,N_12439);
nand U15697 (N_15697,N_12672,N_12053);
nor U15698 (N_15698,N_12607,N_13532);
and U15699 (N_15699,N_12164,N_12860);
nand U15700 (N_15700,N_12496,N_13872);
nor U15701 (N_15701,N_13578,N_13554);
nor U15702 (N_15702,N_12153,N_13286);
nand U15703 (N_15703,N_12265,N_13947);
nand U15704 (N_15704,N_13631,N_13868);
xnor U15705 (N_15705,N_12612,N_12273);
nor U15706 (N_15706,N_13286,N_13716);
or U15707 (N_15707,N_12742,N_12553);
xnor U15708 (N_15708,N_12882,N_13946);
nor U15709 (N_15709,N_12257,N_13310);
and U15710 (N_15710,N_13238,N_12151);
nor U15711 (N_15711,N_13603,N_12922);
nor U15712 (N_15712,N_13780,N_12368);
and U15713 (N_15713,N_13216,N_12792);
or U15714 (N_15714,N_13679,N_13645);
or U15715 (N_15715,N_12745,N_13036);
xnor U15716 (N_15716,N_12551,N_12715);
or U15717 (N_15717,N_13507,N_13863);
nor U15718 (N_15718,N_13095,N_12138);
xnor U15719 (N_15719,N_13169,N_13694);
and U15720 (N_15720,N_13320,N_12613);
nand U15721 (N_15721,N_13198,N_13342);
xor U15722 (N_15722,N_12859,N_12920);
and U15723 (N_15723,N_13228,N_13465);
nor U15724 (N_15724,N_12499,N_13443);
and U15725 (N_15725,N_13253,N_13663);
nor U15726 (N_15726,N_12241,N_12060);
nand U15727 (N_15727,N_12560,N_12652);
or U15728 (N_15728,N_12252,N_13278);
nor U15729 (N_15729,N_12165,N_12727);
or U15730 (N_15730,N_13051,N_12851);
nor U15731 (N_15731,N_12563,N_13495);
nand U15732 (N_15732,N_13724,N_13220);
and U15733 (N_15733,N_12877,N_12492);
nor U15734 (N_15734,N_13764,N_12420);
xnor U15735 (N_15735,N_13718,N_13182);
nor U15736 (N_15736,N_13540,N_12564);
nand U15737 (N_15737,N_13626,N_13670);
nand U15738 (N_15738,N_12177,N_12853);
nor U15739 (N_15739,N_12431,N_12475);
nand U15740 (N_15740,N_12180,N_13855);
nand U15741 (N_15741,N_12265,N_13476);
or U15742 (N_15742,N_12639,N_12498);
nand U15743 (N_15743,N_13197,N_12176);
nor U15744 (N_15744,N_13974,N_13464);
and U15745 (N_15745,N_12441,N_12351);
or U15746 (N_15746,N_12156,N_13999);
xnor U15747 (N_15747,N_13318,N_13289);
xor U15748 (N_15748,N_12801,N_12965);
or U15749 (N_15749,N_13005,N_13357);
nand U15750 (N_15750,N_13971,N_13557);
nor U15751 (N_15751,N_13647,N_13382);
or U15752 (N_15752,N_13495,N_12904);
xnor U15753 (N_15753,N_13421,N_12186);
or U15754 (N_15754,N_13183,N_13036);
or U15755 (N_15755,N_12231,N_13936);
or U15756 (N_15756,N_12119,N_13947);
nor U15757 (N_15757,N_13030,N_13123);
nor U15758 (N_15758,N_12483,N_13262);
or U15759 (N_15759,N_13589,N_12061);
nand U15760 (N_15760,N_13408,N_12898);
and U15761 (N_15761,N_12146,N_13772);
xnor U15762 (N_15762,N_13698,N_13786);
and U15763 (N_15763,N_13835,N_13793);
or U15764 (N_15764,N_12520,N_12109);
or U15765 (N_15765,N_13880,N_13564);
nor U15766 (N_15766,N_12765,N_13579);
or U15767 (N_15767,N_12482,N_12879);
nor U15768 (N_15768,N_13732,N_12116);
nor U15769 (N_15769,N_13743,N_12532);
and U15770 (N_15770,N_13406,N_13109);
nor U15771 (N_15771,N_13109,N_13015);
nand U15772 (N_15772,N_12450,N_12944);
nor U15773 (N_15773,N_12341,N_13305);
and U15774 (N_15774,N_12006,N_13623);
nand U15775 (N_15775,N_12281,N_12232);
and U15776 (N_15776,N_12699,N_12743);
nand U15777 (N_15777,N_12725,N_13349);
nand U15778 (N_15778,N_12067,N_13596);
or U15779 (N_15779,N_12045,N_12688);
xnor U15780 (N_15780,N_12837,N_13305);
or U15781 (N_15781,N_12944,N_13067);
or U15782 (N_15782,N_13297,N_12648);
and U15783 (N_15783,N_13493,N_12132);
and U15784 (N_15784,N_13186,N_13175);
nand U15785 (N_15785,N_13833,N_13254);
nor U15786 (N_15786,N_12036,N_13930);
or U15787 (N_15787,N_12060,N_13716);
or U15788 (N_15788,N_13145,N_12417);
nand U15789 (N_15789,N_12717,N_13309);
nor U15790 (N_15790,N_12938,N_13688);
xor U15791 (N_15791,N_13407,N_12432);
nand U15792 (N_15792,N_12228,N_12614);
or U15793 (N_15793,N_13078,N_13643);
nand U15794 (N_15794,N_12372,N_13572);
and U15795 (N_15795,N_13346,N_12927);
xnor U15796 (N_15796,N_12946,N_12775);
and U15797 (N_15797,N_12715,N_12396);
nand U15798 (N_15798,N_13110,N_13815);
xor U15799 (N_15799,N_12294,N_13467);
nand U15800 (N_15800,N_12779,N_13276);
nor U15801 (N_15801,N_12730,N_13748);
xor U15802 (N_15802,N_13490,N_12765);
nand U15803 (N_15803,N_13254,N_12224);
xnor U15804 (N_15804,N_13999,N_13370);
and U15805 (N_15805,N_13323,N_12887);
nand U15806 (N_15806,N_13938,N_13928);
nand U15807 (N_15807,N_13432,N_12973);
and U15808 (N_15808,N_12096,N_12592);
xor U15809 (N_15809,N_13425,N_13177);
nand U15810 (N_15810,N_13481,N_13088);
nor U15811 (N_15811,N_13515,N_12231);
nand U15812 (N_15812,N_13594,N_13525);
nor U15813 (N_15813,N_12859,N_13345);
xor U15814 (N_15814,N_13845,N_13066);
nor U15815 (N_15815,N_13009,N_12040);
and U15816 (N_15816,N_12482,N_13013);
nand U15817 (N_15817,N_12572,N_12684);
xnor U15818 (N_15818,N_12229,N_13332);
and U15819 (N_15819,N_12563,N_13511);
nor U15820 (N_15820,N_12222,N_13964);
xnor U15821 (N_15821,N_13900,N_13187);
or U15822 (N_15822,N_13757,N_13992);
and U15823 (N_15823,N_12980,N_12932);
and U15824 (N_15824,N_13521,N_12902);
nand U15825 (N_15825,N_12211,N_13628);
xnor U15826 (N_15826,N_12172,N_13266);
nand U15827 (N_15827,N_12533,N_13278);
nor U15828 (N_15828,N_13588,N_13503);
nand U15829 (N_15829,N_12424,N_13393);
xnor U15830 (N_15830,N_13215,N_13563);
nand U15831 (N_15831,N_12586,N_12712);
and U15832 (N_15832,N_12754,N_13958);
and U15833 (N_15833,N_13732,N_13130);
nor U15834 (N_15834,N_12542,N_12855);
or U15835 (N_15835,N_13690,N_13351);
or U15836 (N_15836,N_12284,N_12244);
or U15837 (N_15837,N_12013,N_13394);
and U15838 (N_15838,N_12016,N_13617);
nand U15839 (N_15839,N_13328,N_13128);
or U15840 (N_15840,N_12069,N_12995);
or U15841 (N_15841,N_13751,N_13049);
nor U15842 (N_15842,N_13102,N_12055);
xor U15843 (N_15843,N_12052,N_12059);
nor U15844 (N_15844,N_13910,N_13439);
or U15845 (N_15845,N_13282,N_12029);
or U15846 (N_15846,N_12539,N_13803);
nor U15847 (N_15847,N_13665,N_13677);
and U15848 (N_15848,N_12322,N_12567);
xor U15849 (N_15849,N_13068,N_13632);
or U15850 (N_15850,N_13720,N_12318);
nor U15851 (N_15851,N_12912,N_13570);
xnor U15852 (N_15852,N_12278,N_12551);
xor U15853 (N_15853,N_12566,N_12718);
xnor U15854 (N_15854,N_13608,N_13564);
nor U15855 (N_15855,N_13813,N_13949);
nand U15856 (N_15856,N_12083,N_13359);
nand U15857 (N_15857,N_12138,N_13165);
or U15858 (N_15858,N_13184,N_12309);
nor U15859 (N_15859,N_12557,N_13194);
xnor U15860 (N_15860,N_12712,N_12234);
and U15861 (N_15861,N_12400,N_13610);
or U15862 (N_15862,N_13267,N_12314);
xnor U15863 (N_15863,N_13410,N_12794);
nand U15864 (N_15864,N_12451,N_13063);
xnor U15865 (N_15865,N_12808,N_12340);
xnor U15866 (N_15866,N_12364,N_13037);
and U15867 (N_15867,N_12668,N_12424);
xnor U15868 (N_15868,N_12538,N_13257);
or U15869 (N_15869,N_13270,N_12160);
nand U15870 (N_15870,N_12363,N_13877);
nor U15871 (N_15871,N_13782,N_13296);
xnor U15872 (N_15872,N_13951,N_13572);
nor U15873 (N_15873,N_13436,N_12429);
nand U15874 (N_15874,N_13018,N_13440);
and U15875 (N_15875,N_13790,N_13354);
and U15876 (N_15876,N_13386,N_12949);
nand U15877 (N_15877,N_13710,N_12882);
or U15878 (N_15878,N_13306,N_13259);
nand U15879 (N_15879,N_12929,N_12409);
and U15880 (N_15880,N_13558,N_13175);
xor U15881 (N_15881,N_13941,N_12729);
nor U15882 (N_15882,N_13315,N_13939);
nor U15883 (N_15883,N_13620,N_13366);
or U15884 (N_15884,N_12771,N_13719);
xor U15885 (N_15885,N_13033,N_12238);
and U15886 (N_15886,N_12585,N_12499);
and U15887 (N_15887,N_13954,N_12040);
xor U15888 (N_15888,N_12485,N_13627);
and U15889 (N_15889,N_13590,N_12152);
or U15890 (N_15890,N_13803,N_12460);
and U15891 (N_15891,N_13159,N_12671);
xor U15892 (N_15892,N_13356,N_12584);
nor U15893 (N_15893,N_13374,N_13823);
nor U15894 (N_15894,N_12413,N_12314);
xnor U15895 (N_15895,N_12311,N_13327);
nand U15896 (N_15896,N_12566,N_12649);
nand U15897 (N_15897,N_12966,N_13481);
nor U15898 (N_15898,N_12544,N_13064);
or U15899 (N_15899,N_12718,N_12152);
nand U15900 (N_15900,N_13416,N_13612);
and U15901 (N_15901,N_12714,N_12699);
nand U15902 (N_15902,N_13157,N_12997);
or U15903 (N_15903,N_13711,N_12246);
xnor U15904 (N_15904,N_13964,N_12935);
nand U15905 (N_15905,N_12388,N_13565);
nor U15906 (N_15906,N_12878,N_13955);
nand U15907 (N_15907,N_13683,N_12879);
or U15908 (N_15908,N_12583,N_12006);
xor U15909 (N_15909,N_13580,N_13429);
nand U15910 (N_15910,N_13829,N_13076);
and U15911 (N_15911,N_13064,N_12015);
xnor U15912 (N_15912,N_13975,N_13168);
xnor U15913 (N_15913,N_12449,N_12210);
xor U15914 (N_15914,N_13236,N_12555);
xor U15915 (N_15915,N_12914,N_13209);
or U15916 (N_15916,N_12670,N_12058);
and U15917 (N_15917,N_12925,N_12773);
and U15918 (N_15918,N_13008,N_13834);
nand U15919 (N_15919,N_12106,N_13547);
xnor U15920 (N_15920,N_13786,N_13100);
or U15921 (N_15921,N_12268,N_12834);
or U15922 (N_15922,N_12765,N_13664);
nor U15923 (N_15923,N_12838,N_13638);
xor U15924 (N_15924,N_12062,N_12936);
nand U15925 (N_15925,N_12242,N_12330);
nor U15926 (N_15926,N_13045,N_12054);
or U15927 (N_15927,N_12596,N_12452);
or U15928 (N_15928,N_13702,N_13786);
xnor U15929 (N_15929,N_12044,N_12399);
or U15930 (N_15930,N_13426,N_12425);
or U15931 (N_15931,N_12425,N_12928);
or U15932 (N_15932,N_13549,N_13132);
or U15933 (N_15933,N_12129,N_13348);
or U15934 (N_15934,N_13488,N_13008);
nor U15935 (N_15935,N_12903,N_13653);
xor U15936 (N_15936,N_12567,N_13371);
xor U15937 (N_15937,N_13329,N_12546);
xnor U15938 (N_15938,N_13540,N_12733);
nand U15939 (N_15939,N_12368,N_13205);
nand U15940 (N_15940,N_13029,N_13186);
and U15941 (N_15941,N_13941,N_12087);
and U15942 (N_15942,N_13055,N_13940);
and U15943 (N_15943,N_12001,N_12951);
nand U15944 (N_15944,N_12844,N_13119);
xnor U15945 (N_15945,N_12963,N_12912);
or U15946 (N_15946,N_13080,N_13032);
nand U15947 (N_15947,N_13913,N_13716);
nor U15948 (N_15948,N_12226,N_12951);
nand U15949 (N_15949,N_13479,N_12033);
and U15950 (N_15950,N_12055,N_12563);
nand U15951 (N_15951,N_13465,N_13364);
nand U15952 (N_15952,N_12069,N_12382);
nand U15953 (N_15953,N_13247,N_13438);
and U15954 (N_15954,N_12216,N_13760);
xor U15955 (N_15955,N_12834,N_12174);
nor U15956 (N_15956,N_13454,N_12152);
nand U15957 (N_15957,N_12102,N_13481);
or U15958 (N_15958,N_13479,N_12129);
nor U15959 (N_15959,N_12602,N_12132);
xnor U15960 (N_15960,N_13891,N_12819);
and U15961 (N_15961,N_12662,N_12790);
nand U15962 (N_15962,N_13136,N_12921);
xor U15963 (N_15963,N_13103,N_12897);
xor U15964 (N_15964,N_12041,N_12366);
and U15965 (N_15965,N_13769,N_12553);
nor U15966 (N_15966,N_13071,N_12884);
nor U15967 (N_15967,N_13462,N_13851);
nand U15968 (N_15968,N_13472,N_12398);
xnor U15969 (N_15969,N_13954,N_12290);
nor U15970 (N_15970,N_13759,N_12229);
and U15971 (N_15971,N_13117,N_13703);
or U15972 (N_15972,N_13400,N_12151);
nor U15973 (N_15973,N_13351,N_12538);
or U15974 (N_15974,N_12424,N_12705);
nand U15975 (N_15975,N_13448,N_13701);
nand U15976 (N_15976,N_12108,N_12921);
and U15977 (N_15977,N_12850,N_12833);
nand U15978 (N_15978,N_12304,N_13448);
xor U15979 (N_15979,N_13263,N_13598);
nand U15980 (N_15980,N_12067,N_13593);
xnor U15981 (N_15981,N_12224,N_12693);
or U15982 (N_15982,N_13747,N_12185);
and U15983 (N_15983,N_12773,N_12615);
or U15984 (N_15984,N_13146,N_12480);
nor U15985 (N_15985,N_12968,N_13626);
nor U15986 (N_15986,N_12525,N_12578);
nor U15987 (N_15987,N_12708,N_13294);
xor U15988 (N_15988,N_12818,N_12548);
nand U15989 (N_15989,N_12958,N_12012);
nand U15990 (N_15990,N_12107,N_13595);
and U15991 (N_15991,N_13085,N_12206);
xnor U15992 (N_15992,N_12271,N_12553);
and U15993 (N_15993,N_13687,N_12615);
nand U15994 (N_15994,N_13484,N_13619);
nand U15995 (N_15995,N_12091,N_12182);
and U15996 (N_15996,N_12391,N_13649);
nand U15997 (N_15997,N_12454,N_12335);
xor U15998 (N_15998,N_13340,N_13079);
and U15999 (N_15999,N_13672,N_12865);
and U16000 (N_16000,N_15571,N_15377);
and U16001 (N_16001,N_15016,N_15359);
xor U16002 (N_16002,N_15372,N_14644);
xor U16003 (N_16003,N_15575,N_15945);
or U16004 (N_16004,N_15811,N_15090);
and U16005 (N_16005,N_15653,N_15005);
xnor U16006 (N_16006,N_15553,N_15710);
or U16007 (N_16007,N_14656,N_15364);
nand U16008 (N_16008,N_15983,N_15762);
nor U16009 (N_16009,N_14290,N_14127);
or U16010 (N_16010,N_15104,N_14960);
and U16011 (N_16011,N_15288,N_15332);
or U16012 (N_16012,N_15108,N_15084);
nand U16013 (N_16013,N_15486,N_15728);
xor U16014 (N_16014,N_15740,N_14162);
nand U16015 (N_16015,N_14748,N_14492);
nand U16016 (N_16016,N_15257,N_15695);
nand U16017 (N_16017,N_15944,N_14938);
xnor U16018 (N_16018,N_14347,N_15927);
and U16019 (N_16019,N_15252,N_14310);
xnor U16020 (N_16020,N_14045,N_15806);
and U16021 (N_16021,N_14589,N_15787);
and U16022 (N_16022,N_14762,N_14599);
nand U16023 (N_16023,N_15764,N_15441);
xnor U16024 (N_16024,N_15176,N_15069);
and U16025 (N_16025,N_14374,N_15092);
nor U16026 (N_16026,N_14072,N_15051);
nand U16027 (N_16027,N_15459,N_14533);
nor U16028 (N_16028,N_15131,N_15815);
xnor U16029 (N_16029,N_14726,N_14626);
xor U16030 (N_16030,N_15249,N_15211);
xnor U16031 (N_16031,N_15260,N_15151);
or U16032 (N_16032,N_14957,N_14517);
nor U16033 (N_16033,N_15192,N_15919);
xnor U16034 (N_16034,N_15129,N_14569);
and U16035 (N_16035,N_14897,N_14623);
xnor U16036 (N_16036,N_14831,N_15440);
and U16037 (N_16037,N_15873,N_14013);
and U16038 (N_16038,N_15573,N_14435);
and U16039 (N_16039,N_15296,N_15093);
or U16040 (N_16040,N_14051,N_15847);
nor U16041 (N_16041,N_15198,N_15253);
nor U16042 (N_16042,N_14036,N_15026);
or U16043 (N_16043,N_15742,N_15098);
nand U16044 (N_16044,N_14945,N_14886);
nor U16045 (N_16045,N_14033,N_14705);
xnor U16046 (N_16046,N_14559,N_14203);
nand U16047 (N_16047,N_14415,N_14075);
or U16048 (N_16048,N_15250,N_14985);
and U16049 (N_16049,N_14200,N_14242);
or U16050 (N_16050,N_15770,N_14329);
or U16051 (N_16051,N_14638,N_14506);
xnor U16052 (N_16052,N_14659,N_15791);
nor U16053 (N_16053,N_14970,N_14685);
xor U16054 (N_16054,N_14881,N_14229);
and U16055 (N_16055,N_14201,N_14025);
xor U16056 (N_16056,N_14912,N_14063);
and U16057 (N_16057,N_15401,N_14348);
nor U16058 (N_16058,N_14742,N_14512);
and U16059 (N_16059,N_14793,N_15236);
or U16060 (N_16060,N_14378,N_15545);
nand U16061 (N_16061,N_15813,N_14670);
or U16062 (N_16062,N_15772,N_15941);
nand U16063 (N_16063,N_15404,N_15608);
nand U16064 (N_16064,N_15088,N_14009);
nand U16065 (N_16065,N_15693,N_15833);
xnor U16066 (N_16066,N_14819,N_15230);
and U16067 (N_16067,N_15962,N_15706);
nor U16068 (N_16068,N_14604,N_14430);
nand U16069 (N_16069,N_15495,N_14543);
and U16070 (N_16070,N_14826,N_14947);
xor U16071 (N_16071,N_15938,N_14620);
nand U16072 (N_16072,N_14278,N_14151);
nor U16073 (N_16073,N_14707,N_15530);
xor U16074 (N_16074,N_14469,N_15474);
and U16075 (N_16075,N_14518,N_15515);
xnor U16076 (N_16076,N_14014,N_14850);
or U16077 (N_16077,N_14382,N_15000);
or U16078 (N_16078,N_14001,N_14528);
or U16079 (N_16079,N_15623,N_14885);
nand U16080 (N_16080,N_14916,N_14529);
nand U16081 (N_16081,N_15605,N_14178);
xor U16082 (N_16082,N_14183,N_14166);
and U16083 (N_16083,N_15760,N_15013);
or U16084 (N_16084,N_15731,N_14216);
nand U16085 (N_16085,N_14526,N_15353);
nand U16086 (N_16086,N_14769,N_14114);
nand U16087 (N_16087,N_15914,N_14069);
xnor U16088 (N_16088,N_14806,N_14925);
and U16089 (N_16089,N_14384,N_15067);
nand U16090 (N_16090,N_15113,N_15667);
nand U16091 (N_16091,N_15354,N_14611);
and U16092 (N_16092,N_15527,N_14699);
or U16093 (N_16093,N_15763,N_15326);
or U16094 (N_16094,N_14815,N_15507);
nand U16095 (N_16095,N_15876,N_14205);
xor U16096 (N_16096,N_14675,N_15334);
or U16097 (N_16097,N_14610,N_14580);
nor U16098 (N_16098,N_14505,N_14299);
or U16099 (N_16099,N_14591,N_14573);
and U16100 (N_16100,N_14787,N_14365);
xnor U16101 (N_16101,N_14551,N_15384);
and U16102 (N_16102,N_14639,N_14175);
xor U16103 (N_16103,N_15902,N_15532);
xnor U16104 (N_16104,N_14943,N_14406);
and U16105 (N_16105,N_14164,N_14437);
nor U16106 (N_16106,N_15061,N_14086);
or U16107 (N_16107,N_14463,N_15274);
xnor U16108 (N_16108,N_15637,N_15950);
and U16109 (N_16109,N_14373,N_14770);
nor U16110 (N_16110,N_15700,N_15598);
nor U16111 (N_16111,N_15947,N_14830);
or U16112 (N_16112,N_14750,N_14657);
and U16113 (N_16113,N_15294,N_14956);
xor U16114 (N_16114,N_14917,N_14153);
xnor U16115 (N_16115,N_15768,N_15738);
xor U16116 (N_16116,N_14377,N_14240);
nor U16117 (N_16117,N_14062,N_15814);
nand U16118 (N_16118,N_15722,N_14088);
nor U16119 (N_16119,N_15099,N_14444);
and U16120 (N_16120,N_14005,N_14673);
nor U16121 (N_16121,N_14050,N_14052);
or U16122 (N_16122,N_15704,N_15665);
nand U16123 (N_16123,N_14284,N_14157);
xor U16124 (N_16124,N_15786,N_14398);
nor U16125 (N_16125,N_14027,N_14358);
xnor U16126 (N_16126,N_14988,N_14309);
nand U16127 (N_16127,N_15759,N_15227);
nand U16128 (N_16128,N_15087,N_14766);
xor U16129 (N_16129,N_14434,N_14305);
nand U16130 (N_16130,N_15380,N_14801);
and U16131 (N_16131,N_15362,N_15702);
or U16132 (N_16132,N_15863,N_15984);
xor U16133 (N_16133,N_15389,N_14394);
nor U16134 (N_16134,N_14649,N_15855);
xor U16135 (N_16135,N_14385,N_14691);
nand U16136 (N_16136,N_15449,N_15106);
nand U16137 (N_16137,N_15552,N_14333);
or U16138 (N_16138,N_15986,N_15980);
or U16139 (N_16139,N_14308,N_15671);
or U16140 (N_16140,N_14828,N_15133);
or U16141 (N_16141,N_15295,N_15402);
xor U16142 (N_16142,N_14368,N_14584);
xnor U16143 (N_16143,N_15641,N_14570);
nand U16144 (N_16144,N_15497,N_15411);
or U16145 (N_16145,N_14028,N_15971);
nand U16146 (N_16146,N_15455,N_15164);
and U16147 (N_16147,N_14474,N_15679);
nor U16148 (N_16148,N_14379,N_14545);
nand U16149 (N_16149,N_15062,N_14091);
nor U16150 (N_16150,N_14338,N_15718);
nor U16151 (N_16151,N_14751,N_15564);
and U16152 (N_16152,N_14362,N_15270);
xnor U16153 (N_16153,N_15821,N_14058);
and U16154 (N_16154,N_15994,N_15419);
and U16155 (N_16155,N_15923,N_14558);
or U16156 (N_16156,N_15042,N_14195);
and U16157 (N_16157,N_15145,N_14143);
nor U16158 (N_16158,N_14919,N_14432);
xor U16159 (N_16159,N_15444,N_15720);
and U16160 (N_16160,N_15032,N_14140);
or U16161 (N_16161,N_15010,N_15550);
nand U16162 (N_16162,N_15559,N_14958);
or U16163 (N_16163,N_14120,N_14789);
or U16164 (N_16164,N_14171,N_15154);
nor U16165 (N_16165,N_15872,N_14856);
or U16166 (N_16166,N_15707,N_14461);
or U16167 (N_16167,N_15115,N_15511);
or U16168 (N_16168,N_15243,N_15796);
nand U16169 (N_16169,N_15029,N_14669);
or U16170 (N_16170,N_15551,N_15269);
nor U16171 (N_16171,N_14319,N_14079);
nor U16172 (N_16172,N_15325,N_14287);
or U16173 (N_16173,N_14540,N_15566);
nor U16174 (N_16174,N_14711,N_14668);
or U16175 (N_16175,N_14318,N_15186);
and U16176 (N_16176,N_15469,N_14489);
xor U16177 (N_16177,N_14070,N_15612);
nand U16178 (N_16178,N_15283,N_14633);
nor U16179 (N_16179,N_14129,N_15827);
nand U16180 (N_16180,N_14767,N_15057);
or U16181 (N_16181,N_15238,N_15157);
xor U16182 (N_16182,N_14927,N_15022);
nor U16183 (N_16183,N_15300,N_14900);
xor U16184 (N_16184,N_14262,N_15398);
nand U16185 (N_16185,N_14860,N_15340);
or U16186 (N_16186,N_14875,N_15691);
nand U16187 (N_16187,N_14614,N_14321);
and U16188 (N_16188,N_15975,N_15666);
or U16189 (N_16189,N_14781,N_14878);
nand U16190 (N_16190,N_15795,N_15174);
xnor U16191 (N_16191,N_15156,N_15989);
nor U16192 (N_16192,N_15820,N_15263);
nor U16193 (N_16193,N_15144,N_14500);
and U16194 (N_16194,N_14887,N_14953);
xnor U16195 (N_16195,N_15278,N_14547);
and U16196 (N_16196,N_15431,N_15554);
nor U16197 (N_16197,N_14335,N_14977);
nand U16198 (N_16198,N_14163,N_14986);
or U16199 (N_16199,N_15542,N_15500);
nor U16200 (N_16200,N_14983,N_15755);
nand U16201 (N_16201,N_14152,N_14752);
and U16202 (N_16202,N_14892,N_14672);
xnor U16203 (N_16203,N_14267,N_14316);
and U16204 (N_16204,N_15044,N_15118);
and U16205 (N_16205,N_15281,N_15990);
and U16206 (N_16206,N_14269,N_15737);
nand U16207 (N_16207,N_14150,N_14807);
nor U16208 (N_16208,N_15064,N_14293);
xnor U16209 (N_16209,N_14590,N_15675);
nor U16210 (N_16210,N_14544,N_15966);
and U16211 (N_16211,N_14468,N_15898);
nor U16212 (N_16212,N_15767,N_14303);
xor U16213 (N_16213,N_14835,N_14412);
nand U16214 (N_16214,N_14708,N_14930);
and U16215 (N_16215,N_15878,N_15529);
nor U16216 (N_16216,N_14342,N_14763);
nand U16217 (N_16217,N_14778,N_15881);
and U16218 (N_16218,N_15313,N_14627);
xnor U16219 (N_16219,N_15793,N_14901);
or U16220 (N_16220,N_14593,N_15732);
xor U16221 (N_16221,N_14966,N_15447);
or U16222 (N_16222,N_14999,N_14566);
xor U16223 (N_16223,N_15512,N_14660);
nand U16224 (N_16224,N_15925,N_15930);
xor U16225 (N_16225,N_14652,N_15960);
nor U16226 (N_16226,N_14263,N_15361);
and U16227 (N_16227,N_14124,N_14247);
nor U16228 (N_16228,N_15711,N_15785);
xor U16229 (N_16229,N_14509,N_15794);
and U16230 (N_16230,N_15972,N_14745);
nand U16231 (N_16231,N_14786,N_14926);
or U16232 (N_16232,N_14252,N_14243);
nor U16233 (N_16233,N_15482,N_14121);
nor U16234 (N_16234,N_15100,N_14940);
nor U16235 (N_16235,N_15163,N_14737);
nand U16236 (N_16236,N_14413,N_15579);
or U16237 (N_16237,N_15105,N_15019);
and U16238 (N_16238,N_15289,N_14702);
nor U16239 (N_16239,N_15286,N_14425);
xnor U16240 (N_16240,N_15309,N_15824);
and U16241 (N_16241,N_15913,N_15150);
xnor U16242 (N_16242,N_15287,N_14641);
and U16243 (N_16243,N_15611,N_14857);
or U16244 (N_16244,N_14426,N_14785);
or U16245 (N_16245,N_14775,N_15922);
nand U16246 (N_16246,N_14888,N_15991);
nand U16247 (N_16247,N_14055,N_14395);
or U16248 (N_16248,N_14113,N_14709);
nand U16249 (N_16249,N_15639,N_15981);
xnor U16250 (N_16250,N_14965,N_15357);
or U16251 (N_16251,N_15582,N_15304);
xor U16252 (N_16252,N_14992,N_14331);
and U16253 (N_16253,N_15436,N_15319);
or U16254 (N_16254,N_14496,N_14391);
nor U16255 (N_16255,N_15850,N_15382);
nand U16256 (N_16256,N_14019,N_15912);
and U16257 (N_16257,N_15077,N_14583);
nor U16258 (N_16258,N_15739,N_15298);
and U16259 (N_16259,N_15948,N_15830);
nand U16260 (N_16260,N_15617,N_14723);
or U16261 (N_16261,N_14248,N_14768);
xor U16262 (N_16262,N_15328,N_15640);
nand U16263 (N_16263,N_15125,N_14054);
nand U16264 (N_16264,N_15102,N_15951);
xor U16265 (N_16265,N_14771,N_14225);
nor U16266 (N_16266,N_14096,N_15807);
xnor U16267 (N_16267,N_14936,N_14400);
nand U16268 (N_16268,N_14681,N_15117);
nor U16269 (N_16269,N_14721,N_15883);
nand U16270 (N_16270,N_15537,N_14997);
nor U16271 (N_16271,N_14824,N_14695);
nor U16272 (N_16272,N_15668,N_15874);
xnor U16273 (N_16273,N_15909,N_15526);
xnor U16274 (N_16274,N_15674,N_14450);
nor U16275 (N_16275,N_14409,N_14845);
xor U16276 (N_16276,N_14217,N_14630);
nand U16277 (N_16277,N_15242,N_15413);
nor U16278 (N_16278,N_14613,N_14396);
and U16279 (N_16279,N_14577,N_15776);
nand U16280 (N_16280,N_14834,N_15757);
or U16281 (N_16281,N_15030,N_14250);
or U16282 (N_16282,N_14585,N_14112);
nand U16283 (N_16283,N_14967,N_14294);
nor U16284 (N_16284,N_15386,N_15730);
xor U16285 (N_16285,N_14792,N_14193);
nand U16286 (N_16286,N_14433,N_14061);
or U16287 (N_16287,N_15047,N_14292);
xnor U16288 (N_16288,N_15387,N_15200);
and U16289 (N_16289,N_15181,N_14109);
xor U16290 (N_16290,N_14740,N_14990);
or U16291 (N_16291,N_15426,N_15293);
xor U16292 (N_16292,N_15475,N_14441);
xnor U16293 (N_16293,N_15658,N_15222);
and U16294 (N_16294,N_14504,N_15725);
nor U16295 (N_16295,N_14950,N_14607);
and U16296 (N_16296,N_15819,N_14186);
nor U16297 (N_16297,N_14710,N_15462);
or U16298 (N_16298,N_14893,N_15086);
xor U16299 (N_16299,N_14224,N_15453);
nand U16300 (N_16300,N_15011,N_15204);
and U16301 (N_16301,N_14961,N_15081);
and U16302 (N_16302,N_15835,N_15631);
nor U16303 (N_16303,N_14363,N_14414);
or U16304 (N_16304,N_14475,N_15038);
nor U16305 (N_16305,N_15134,N_15318);
and U16306 (N_16306,N_14531,N_14882);
nand U16307 (N_16307,N_14905,N_14858);
nor U16308 (N_16308,N_15247,N_14431);
or U16309 (N_16309,N_14448,N_14773);
nand U16310 (N_16310,N_15258,N_14941);
or U16311 (N_16311,N_15660,N_14066);
xnor U16312 (N_16312,N_15729,N_15433);
nand U16313 (N_16313,N_14862,N_14827);
xnor U16314 (N_16314,N_14777,N_14865);
and U16315 (N_16315,N_15799,N_14389);
or U16316 (N_16316,N_14064,N_15329);
nand U16317 (N_16317,N_15977,N_15333);
xor U16318 (N_16318,N_15771,N_15607);
or U16319 (N_16319,N_15004,N_15632);
or U16320 (N_16320,N_15219,N_15544);
nor U16321 (N_16321,N_15306,N_14738);
nand U16322 (N_16322,N_14106,N_14562);
or U16323 (N_16323,N_15208,N_14408);
or U16324 (N_16324,N_15392,N_14549);
xnor U16325 (N_16325,N_15454,N_15993);
xnor U16326 (N_16326,N_15973,N_15369);
xor U16327 (N_16327,N_14800,N_15890);
or U16328 (N_16328,N_14780,N_14536);
and U16329 (N_16329,N_15533,N_14173);
xnor U16330 (N_16330,N_14954,N_15645);
nor U16331 (N_16331,N_14654,N_14497);
nor U16332 (N_16332,N_15160,N_15240);
xor U16333 (N_16333,N_14154,N_15578);
nor U16334 (N_16334,N_15390,N_14706);
nand U16335 (N_16335,N_15655,N_14077);
nand U16336 (N_16336,N_14161,N_15320);
nand U16337 (N_16337,N_14913,N_14510);
or U16338 (N_16338,N_15746,N_14747);
nand U16339 (N_16339,N_15373,N_15110);
and U16340 (N_16340,N_14067,N_14073);
nand U16341 (N_16341,N_14371,N_14796);
nor U16342 (N_16342,N_15498,N_15465);
xor U16343 (N_16343,N_14557,N_14976);
xnor U16344 (N_16344,N_14515,N_14390);
xnor U16345 (N_16345,N_15629,N_15792);
nor U16346 (N_16346,N_14920,N_15557);
xnor U16347 (N_16347,N_15625,N_15254);
xnor U16348 (N_16348,N_15997,N_14393);
xor U16349 (N_16349,N_14288,N_15080);
nor U16350 (N_16350,N_15502,N_15988);
or U16351 (N_16351,N_15280,N_14841);
xnor U16352 (N_16352,N_15014,N_15713);
and U16353 (N_16353,N_14023,N_14973);
or U16354 (N_16354,N_15568,N_14791);
or U16355 (N_16355,N_15403,N_15429);
and U16356 (N_16356,N_14816,N_14765);
xor U16357 (N_16357,N_14552,N_15324);
xor U16358 (N_16358,N_14174,N_14179);
nand U16359 (N_16359,N_14041,N_14687);
or U16360 (N_16360,N_14821,N_15936);
nand U16361 (N_16361,N_15107,N_15723);
or U16362 (N_16362,N_15538,N_15301);
nor U16363 (N_16363,N_15158,N_15268);
nor U16364 (N_16364,N_15717,N_14859);
and U16365 (N_16365,N_15052,N_15840);
nor U16366 (N_16366,N_15589,N_14658);
nor U16367 (N_16367,N_15170,N_15095);
xnor U16368 (N_16368,N_14218,N_15998);
or U16369 (N_16369,N_14651,N_14117);
xor U16370 (N_16370,N_15618,N_14251);
xor U16371 (N_16371,N_15416,N_14981);
nand U16372 (N_16372,N_15135,N_14429);
xor U16373 (N_16373,N_14728,N_15128);
or U16374 (N_16374,N_15017,N_14176);
or U16375 (N_16375,N_15173,N_15906);
nand U16376 (N_16376,N_14093,N_15490);
nand U16377 (N_16377,N_14724,N_14126);
and U16378 (N_16378,N_14447,N_15694);
or U16379 (N_16379,N_15692,N_14873);
or U16380 (N_16380,N_14714,N_15009);
xnor U16381 (N_16381,N_15569,N_15572);
xor U16382 (N_16382,N_15567,N_14397);
xor U16383 (N_16383,N_15116,N_14804);
nand U16384 (N_16384,N_14972,N_15060);
nand U16385 (N_16385,N_15335,N_15659);
xor U16386 (N_16386,N_14572,N_14107);
nor U16387 (N_16387,N_15120,N_15905);
and U16388 (N_16388,N_15514,N_15101);
or U16389 (N_16389,N_14494,N_15570);
xor U16390 (N_16390,N_14478,N_14629);
or U16391 (N_16391,N_14464,N_15122);
nor U16392 (N_16392,N_15933,N_14561);
and U16393 (N_16393,N_15834,N_15864);
nor U16394 (N_16394,N_14332,N_15483);
nor U16395 (N_16395,N_15442,N_15634);
and U16396 (N_16396,N_15904,N_14689);
xor U16397 (N_16397,N_14795,N_15037);
or U16398 (N_16398,N_14210,N_15065);
xnor U16399 (N_16399,N_14502,N_15276);
nand U16400 (N_16400,N_15344,N_14256);
nor U16401 (N_16401,N_15229,N_15615);
or U16402 (N_16402,N_14756,N_14291);
nor U16403 (N_16403,N_14460,N_15231);
nor U16404 (N_16404,N_14423,N_15430);
and U16405 (N_16405,N_14277,N_14234);
xor U16406 (N_16406,N_14004,N_14035);
or U16407 (N_16407,N_15210,N_15626);
nor U16408 (N_16408,N_14030,N_15509);
and U16409 (N_16409,N_15593,N_15188);
nor U16410 (N_16410,N_14187,N_15844);
nor U16411 (N_16411,N_14037,N_15916);
xor U16412 (N_16412,N_14046,N_14346);
nand U16413 (N_16413,N_14115,N_14586);
nand U16414 (N_16414,N_14522,N_15642);
and U16415 (N_16415,N_14244,N_15661);
or U16416 (N_16416,N_14898,N_15308);
xnor U16417 (N_16417,N_15696,N_15870);
nor U16418 (N_16418,N_14524,N_15915);
nand U16419 (N_16419,N_15924,N_14727);
or U16420 (N_16420,N_15446,N_15756);
xnor U16421 (N_16421,N_14231,N_15201);
nand U16422 (N_16422,N_15445,N_14190);
nand U16423 (N_16423,N_15149,N_14103);
xor U16424 (N_16424,N_14417,N_14220);
and U16425 (N_16425,N_14537,N_15264);
and U16426 (N_16426,N_15443,N_15487);
or U16427 (N_16427,N_14995,N_15234);
nand U16428 (N_16428,N_15698,N_15432);
or U16429 (N_16429,N_15458,N_14486);
nor U16430 (N_16430,N_15741,N_15506);
xnor U16431 (N_16431,N_15303,N_15745);
xor U16432 (N_16432,N_14717,N_14667);
nor U16433 (N_16433,N_14732,N_15775);
xnor U16434 (N_16434,N_14833,N_15327);
nand U16435 (N_16435,N_15235,N_15774);
nand U16436 (N_16436,N_15769,N_14184);
xnor U16437 (N_16437,N_14065,N_14784);
nand U16438 (N_16438,N_15202,N_15349);
nor U16439 (N_16439,N_15045,N_15932);
nand U16440 (N_16440,N_14158,N_15277);
nor U16441 (N_16441,N_15248,N_14753);
nor U16442 (N_16442,N_15082,N_14491);
and U16443 (N_16443,N_15177,N_15027);
nand U16444 (N_16444,N_14810,N_14105);
and U16445 (N_16445,N_15053,N_14214);
or U16446 (N_16446,N_15143,N_14894);
xor U16447 (N_16447,N_15148,N_14538);
nand U16448 (N_16448,N_15012,N_15321);
and U16449 (N_16449,N_15307,N_15832);
nand U16450 (N_16450,N_15220,N_14198);
nor U16451 (N_16451,N_14369,N_14655);
xnor U16452 (N_16452,N_15866,N_15341);
xor U16453 (N_16453,N_15068,N_15753);
nand U16454 (N_16454,N_14470,N_14471);
and U16455 (N_16455,N_14324,N_15839);
nand U16456 (N_16456,N_14439,N_14653);
nor U16457 (N_16457,N_15385,N_14625);
nor U16458 (N_16458,N_14053,N_15624);
nand U16459 (N_16459,N_14202,N_15501);
and U16460 (N_16460,N_14963,N_15197);
nand U16461 (N_16461,N_15937,N_15895);
xnor U16462 (N_16462,N_14914,N_14146);
xnor U16463 (N_16463,N_14642,N_14191);
nand U16464 (N_16464,N_15493,N_14402);
or U16465 (N_16465,N_15285,N_14133);
xor U16466 (N_16466,N_15338,N_14690);
nor U16467 (N_16467,N_15926,N_15376);
xnor U16468 (N_16468,N_14640,N_14832);
or U16469 (N_16469,N_14692,N_15112);
nor U16470 (N_16470,N_15427,N_14741);
and U16471 (N_16471,N_14836,N_15155);
nand U16472 (N_16472,N_15652,N_14022);
nor U16473 (N_16473,N_14455,N_14488);
nor U16474 (N_16474,N_14910,N_15360);
or U16475 (N_16475,N_14602,N_14869);
nor U16476 (N_16476,N_14301,N_15995);
nand U16477 (N_16477,N_15476,N_15585);
nor U16478 (N_16478,N_15055,N_14746);
nand U16479 (N_16479,N_14459,N_15831);
or U16480 (N_16480,N_15371,N_15588);
and U16481 (N_16481,N_15089,N_15805);
xor U16482 (N_16482,N_15168,N_14328);
nand U16483 (N_16483,N_15789,N_15196);
nand U16484 (N_16484,N_15628,N_15788);
or U16485 (N_16485,N_15302,N_14498);
or U16486 (N_16486,N_15417,N_15003);
or U16487 (N_16487,N_15524,N_14996);
nor U16488 (N_16488,N_15284,N_15246);
xnor U16489 (N_16489,N_14612,N_15630);
nand U16490 (N_16490,N_15072,N_14507);
nor U16491 (N_16491,N_14876,N_15643);
xnor U16492 (N_16492,N_15256,N_15784);
nand U16493 (N_16493,N_14286,N_14006);
or U16494 (N_16494,N_15456,N_15396);
or U16495 (N_16495,N_14405,N_15323);
nand U16496 (N_16496,N_15415,N_14846);
nor U16497 (N_16497,N_14123,N_14024);
nand U16498 (N_16498,N_14078,N_14421);
or U16499 (N_16499,N_15809,N_15565);
nand U16500 (N_16500,N_14131,N_15681);
and U16501 (N_16501,N_15031,N_15314);
xnor U16502 (N_16502,N_14352,N_14587);
nand U16503 (N_16503,N_14908,N_15059);
nand U16504 (N_16504,N_14194,N_15190);
nor U16505 (N_16505,N_14874,N_14386);
or U16506 (N_16506,N_14924,N_14624);
nor U16507 (N_16507,N_15516,N_14232);
or U16508 (N_16508,N_14317,N_14038);
xor U16509 (N_16509,N_15522,N_15315);
and U16510 (N_16510,N_14718,N_15508);
nand U16511 (N_16511,N_15467,N_14137);
and U16512 (N_16512,N_15818,N_15672);
or U16513 (N_16513,N_15407,N_14148);
nor U16514 (N_16514,N_15180,N_15119);
and U16515 (N_16515,N_15856,N_15886);
or U16516 (N_16516,N_14095,N_15383);
and U16517 (N_16517,N_14446,N_14048);
or U16518 (N_16518,N_14595,N_15195);
xnor U16519 (N_16519,N_15233,N_15472);
xnor U16520 (N_16520,N_14241,N_14918);
nor U16521 (N_16521,N_14381,N_14147);
or U16522 (N_16522,N_14661,N_14139);
xor U16523 (N_16523,N_14074,N_15510);
xor U16524 (N_16524,N_14141,N_15959);
or U16525 (N_16525,N_15563,N_15183);
xor U16526 (N_16526,N_15075,N_14090);
nand U16527 (N_16527,N_15751,N_15039);
xnor U16528 (N_16528,N_14853,N_15635);
nand U16529 (N_16529,N_15471,N_15215);
and U16530 (N_16530,N_14647,N_15903);
nand U16531 (N_16531,N_15209,N_14082);
xnor U16532 (N_16532,N_15900,N_15736);
and U16533 (N_16533,N_15169,N_15137);
nor U16534 (N_16534,N_14199,N_15410);
nand U16535 (N_16535,N_14458,N_15056);
nand U16536 (N_16536,N_15686,N_14783);
nand U16537 (N_16537,N_14399,N_15928);
and U16538 (N_16538,N_15034,N_14928);
or U16539 (N_16539,N_15779,N_15697);
or U16540 (N_16540,N_14863,N_15074);
and U16541 (N_16541,N_15644,N_14010);
xnor U16542 (N_16542,N_15648,N_15421);
nand U16543 (N_16543,N_15581,N_14012);
nand U16544 (N_16544,N_15422,N_15956);
nor U16545 (N_16545,N_15867,N_15292);
or U16546 (N_16546,N_15929,N_14160);
and U16547 (N_16547,N_14582,N_15549);
nor U16548 (N_16548,N_14110,N_15114);
nand U16549 (N_16549,N_14868,N_15586);
nor U16550 (N_16550,N_15040,N_14609);
and U16551 (N_16551,N_15152,N_14026);
and U16552 (N_16552,N_15669,N_14228);
nor U16553 (N_16553,N_14473,N_14177);
nor U16554 (N_16554,N_14743,N_15518);
or U16555 (N_16555,N_14635,N_15656);
or U16556 (N_16556,N_15857,N_14092);
or U16557 (N_16557,N_14563,N_14253);
and U16558 (N_16558,N_15712,N_15650);
nor U16559 (N_16559,N_15073,N_14116);
or U16560 (N_16560,N_14255,N_14805);
and U16561 (N_16561,N_14523,N_14731);
nand U16562 (N_16562,N_15761,N_15939);
xnor U16563 (N_16563,N_14196,N_14935);
xnor U16564 (N_16564,N_15002,N_15193);
nor U16565 (N_16565,N_14964,N_14895);
nor U16566 (N_16566,N_15555,N_15781);
and U16567 (N_16567,N_15838,N_14000);
or U16568 (N_16568,N_15802,N_15620);
and U16569 (N_16569,N_15845,N_14682);
nand U16570 (N_16570,N_14034,N_14275);
and U16571 (N_16571,N_14207,N_15424);
or U16572 (N_16572,N_15191,N_15871);
or U16573 (N_16573,N_15803,N_15083);
or U16574 (N_16574,N_14720,N_14168);
nand U16575 (N_16575,N_15893,N_14501);
nand U16576 (N_16576,N_14798,N_15214);
xor U16577 (N_16577,N_15400,N_15663);
and U16578 (N_16578,N_15897,N_14525);
or U16579 (N_16579,N_14605,N_14829);
nor U16580 (N_16580,N_15434,N_15601);
and U16581 (N_16581,N_14211,N_15224);
nor U16582 (N_16582,N_14325,N_14149);
nor U16583 (N_16583,N_15868,N_14678);
or U16584 (N_16584,N_14989,N_14933);
xnor U16585 (N_16585,N_15347,N_15633);
xor U16586 (N_16586,N_14648,N_14820);
nand U16587 (N_16587,N_14754,N_14861);
or U16588 (N_16588,N_15266,N_14703);
xor U16589 (N_16589,N_15790,N_15381);
and U16590 (N_16590,N_14099,N_15646);
nand U16591 (N_16591,N_15539,N_15172);
nor U16592 (N_16592,N_14264,N_14239);
xnor U16593 (N_16593,N_15954,N_14356);
and U16594 (N_16594,N_14080,N_15879);
or U16595 (N_16595,N_14730,N_14759);
nor U16596 (N_16596,N_14327,N_14764);
and U16597 (N_16597,N_14758,N_15141);
nor U16598 (N_16598,N_14962,N_14693);
or U16599 (N_16599,N_14307,N_15969);
and U16600 (N_16600,N_14003,N_15918);
or U16601 (N_16601,N_15379,N_15543);
nand U16602 (N_16602,N_15677,N_15931);
nor U16603 (N_16603,N_14454,N_15316);
xor U16604 (N_16604,N_15992,N_14939);
nor U16605 (N_16605,N_15018,N_14122);
and U16606 (N_16606,N_14987,N_15299);
and U16607 (N_16607,N_14296,N_14235);
nor U16608 (N_16608,N_15531,N_15079);
nand U16609 (N_16609,N_14380,N_15996);
xnor U16610 (N_16610,N_14283,N_15494);
or U16611 (N_16611,N_15780,N_15865);
nor U16612 (N_16612,N_14817,N_14411);
xor U16613 (N_16613,N_15735,N_15754);
xor U16614 (N_16614,N_15262,N_14679);
nand U16615 (N_16615,N_14392,N_15165);
xnor U16616 (N_16616,N_14980,N_15610);
or U16617 (N_16617,N_14039,N_14546);
or U16618 (N_16618,N_14233,N_15091);
nor U16619 (N_16619,N_14044,N_15232);
xnor U16620 (N_16620,N_15297,N_14744);
nand U16621 (N_16621,N_15979,N_14615);
or U16622 (N_16622,N_15752,N_14258);
and U16623 (N_16623,N_14257,N_15778);
and U16624 (N_16624,N_15273,N_14516);
nor U16625 (N_16625,N_15826,N_14755);
or U16626 (N_16626,N_14944,N_14213);
xnor U16627 (N_16627,N_15849,N_15967);
nor U16628 (N_16628,N_14948,N_14616);
nand U16629 (N_16629,N_14942,N_14946);
nor U16630 (N_16630,N_15346,N_14266);
or U16631 (N_16631,N_15690,N_15435);
and U16632 (N_16632,N_14734,N_15964);
and U16633 (N_16633,N_15428,N_15716);
or U16634 (N_16634,N_15008,N_14508);
and U16635 (N_16635,N_14029,N_15602);
nor U16636 (N_16636,N_15370,N_14729);
xor U16637 (N_16637,N_15337,N_14227);
and U16638 (N_16638,N_14937,N_14071);
nand U16639 (N_16639,N_15412,N_14237);
and U16640 (N_16640,N_15733,N_15048);
nand U16641 (N_16641,N_14883,N_15851);
xnor U16642 (N_16642,N_15636,N_14451);
nand U16643 (N_16643,N_14259,N_15758);
and U16644 (N_16644,N_15046,N_14539);
nand U16645 (N_16645,N_15199,N_15703);
and U16646 (N_16646,N_14366,N_14664);
or U16647 (N_16647,N_15466,N_14008);
and U16648 (N_16648,N_14111,N_14081);
or U16649 (N_16649,N_15399,N_15182);
nor U16650 (N_16650,N_14663,N_14031);
nand U16651 (N_16651,N_15899,N_15339);
or U16652 (N_16652,N_14636,N_15452);
or U16653 (N_16653,N_14355,N_15683);
or U16654 (N_16654,N_15734,N_14911);
or U16655 (N_16655,N_15662,N_15638);
nand U16656 (N_16656,N_14594,N_14297);
nand U16657 (N_16657,N_14165,N_14323);
nand U16658 (N_16658,N_14181,N_14312);
xnor U16659 (N_16659,N_14271,N_15358);
or U16660 (N_16660,N_15317,N_14493);
or U16661 (N_16661,N_14383,N_15041);
and U16662 (N_16662,N_14579,N_14298);
xor U16663 (N_16663,N_14733,N_14974);
or U16664 (N_16664,N_14223,N_15457);
nand U16665 (N_16665,N_14554,N_15974);
nand U16666 (N_16666,N_14484,N_14749);
nor U16667 (N_16667,N_14270,N_14467);
and U16668 (N_16668,N_14222,N_14206);
nand U16669 (N_16669,N_14360,N_15670);
nand U16670 (N_16670,N_14011,N_15875);
xnor U16671 (N_16671,N_15606,N_14866);
or U16672 (N_16672,N_15798,N_15351);
and U16673 (N_16673,N_15221,N_15547);
nand U16674 (N_16674,N_14979,N_14694);
or U16675 (N_16675,N_15217,N_14462);
xor U16676 (N_16676,N_15825,N_15777);
xnor U16677 (N_16677,N_14601,N_15955);
nand U16678 (N_16678,N_14404,N_14578);
xnor U16679 (N_16679,N_15271,N_14057);
xnor U16680 (N_16680,N_15085,N_14209);
nor U16681 (N_16681,N_14637,N_14565);
xor U16682 (N_16682,N_14279,N_15917);
and U16683 (N_16683,N_15921,N_15748);
nand U16684 (N_16684,N_15071,N_15305);
nor U16685 (N_16685,N_14597,N_15488);
and U16686 (N_16686,N_15477,N_15654);
xor U16687 (N_16687,N_15773,N_15783);
or U16688 (N_16688,N_14596,N_15935);
nor U16689 (N_16689,N_15721,N_15517);
nand U16690 (N_16690,N_14782,N_14169);
xor U16691 (N_16691,N_14238,N_14085);
or U16692 (N_16692,N_15536,N_15070);
or U16693 (N_16693,N_15212,N_14812);
and U16694 (N_16694,N_14097,N_15460);
and U16695 (N_16695,N_14289,N_14619);
and U16696 (N_16696,N_15616,N_15647);
or U16697 (N_16697,N_15860,N_15492);
and U16698 (N_16698,N_15479,N_14848);
nand U16699 (N_16699,N_15350,N_15395);
or U16700 (N_16700,N_15408,N_15907);
and U16701 (N_16701,N_14320,N_15365);
nor U16702 (N_16702,N_15583,N_14016);
xor U16703 (N_16703,N_15291,N_14847);
nor U16704 (N_16704,N_15884,N_14219);
xnor U16705 (N_16705,N_15049,N_14600);
and U16706 (N_16706,N_14631,N_15161);
nand U16707 (N_16707,N_14118,N_15020);
and U16708 (N_16708,N_15265,N_15021);
or U16709 (N_16709,N_14984,N_14959);
or U16710 (N_16710,N_15162,N_15226);
or U16711 (N_16711,N_15940,N_14719);
and U16712 (N_16712,N_14245,N_14811);
xor U16713 (N_16713,N_14440,N_14145);
nand U16714 (N_16714,N_14854,N_14666);
nand U16715 (N_16715,N_15343,N_15481);
or U16716 (N_16716,N_14665,N_15678);
nor U16717 (N_16717,N_14128,N_14345);
xnor U16718 (N_16718,N_15708,N_15808);
nor U16719 (N_16719,N_14645,N_15858);
xor U16720 (N_16720,N_15178,N_14872);
nand U16721 (N_16721,N_15147,N_14419);
nor U16722 (N_16722,N_15521,N_15574);
xor U16723 (N_16723,N_15078,N_14550);
or U16724 (N_16724,N_15368,N_14132);
nand U16725 (N_16725,N_14416,N_14443);
or U16726 (N_16726,N_14632,N_14825);
or U16727 (N_16727,N_14100,N_15239);
and U16728 (N_16728,N_15499,N_15136);
nor U16729 (N_16729,N_14880,N_14696);
and U16730 (N_16730,N_14592,N_15891);
xor U16731 (N_16731,N_15817,N_14490);
xor U16732 (N_16732,N_14172,N_15138);
nand U16733 (N_16733,N_15393,N_15609);
nand U16734 (N_16734,N_14688,N_14040);
and U16735 (N_16735,N_15461,N_15541);
nor U16736 (N_16736,N_15414,N_14104);
nor U16737 (N_16737,N_14330,N_14273);
xor U16738 (N_16738,N_15970,N_14527);
nand U16739 (N_16739,N_15920,N_14456);
or U16740 (N_16740,N_15999,N_15599);
nand U16741 (N_16741,N_15614,N_14725);
xor U16742 (N_16742,N_15171,N_14134);
nor U16743 (N_16743,N_14932,N_15591);
nor U16744 (N_16744,N_14282,N_14272);
nor U16745 (N_16745,N_14313,N_14891);
xnor U16746 (N_16746,N_14991,N_15418);
nor U16747 (N_16747,N_15709,N_15837);
or U16748 (N_16748,N_15649,N_15908);
nand U16749 (N_16749,N_14621,N_15237);
nand U16750 (N_16750,N_15076,N_14155);
or U16751 (N_16751,N_15958,N_15852);
or U16752 (N_16752,N_14698,N_15800);
and U16753 (N_16753,N_14797,N_15782);
xnor U16754 (N_16754,N_15063,N_15448);
or U16755 (N_16755,N_15103,N_14839);
nor U16756 (N_16756,N_15406,N_14560);
nand U16757 (N_16757,N_14466,N_14553);
and U16758 (N_16758,N_14418,N_15378);
nor U16759 (N_16759,N_15701,N_15175);
or U16760 (N_16760,N_15312,N_14555);
xnor U16761 (N_16761,N_15603,N_14715);
and U16762 (N_16762,N_15388,N_15882);
and U16763 (N_16763,N_14420,N_14364);
or U16764 (N_16764,N_15345,N_14424);
or U16765 (N_16765,N_14167,N_15535);
xnor U16766 (N_16766,N_14877,N_14520);
nand U16767 (N_16767,N_15025,N_15282);
xor U16768 (N_16768,N_14511,N_14341);
xnor U16769 (N_16769,N_15255,N_15841);
nor U16770 (N_16770,N_14903,N_15245);
nor U16771 (N_16771,N_15001,N_15853);
xnor U16772 (N_16772,N_15394,N_14949);
or U16773 (N_16773,N_15132,N_15153);
nand U16774 (N_16774,N_14968,N_14934);
and U16775 (N_16775,N_14774,N_14101);
or U16776 (N_16776,N_14436,N_14503);
nor U16777 (N_16777,N_14156,N_15259);
and U16778 (N_16778,N_15705,N_14842);
nand U16779 (N_16779,N_15952,N_15901);
and U16780 (N_16780,N_15146,N_14618);
nor U16781 (N_16781,N_15023,N_15889);
nor U16782 (N_16782,N_14388,N_15978);
nor U16783 (N_16783,N_15594,N_14068);
or U16784 (N_16784,N_14994,N_14662);
nor U16785 (N_16785,N_14015,N_15468);
and U16786 (N_16786,N_15223,N_14779);
and U16787 (N_16787,N_15965,N_14260);
xnor U16788 (N_16788,N_15478,N_14799);
and U16789 (N_16789,N_15528,N_14541);
or U16790 (N_16790,N_15592,N_14896);
nand U16791 (N_16791,N_14476,N_14513);
xnor U16792 (N_16792,N_15801,N_15126);
nand U16793 (N_16793,N_15525,N_14567);
nand U16794 (N_16794,N_14337,N_14683);
nor U16795 (N_16795,N_15534,N_15946);
nor U16796 (N_16796,N_15627,N_15207);
nand U16797 (N_16797,N_14280,N_15504);
nor U16798 (N_16798,N_14056,N_14226);
or U16799 (N_16799,N_14357,N_14098);
or U16800 (N_16800,N_14849,N_15310);
and U16801 (N_16801,N_14803,N_15621);
and U16802 (N_16802,N_14281,N_15836);
nand U16803 (N_16803,N_14581,N_15375);
and U16804 (N_16804,N_14864,N_14904);
nor U16805 (N_16805,N_14808,N_14410);
xnor U16806 (N_16806,N_15595,N_14844);
nand U16807 (N_16807,N_14757,N_15714);
nor U16808 (N_16808,N_14261,N_15189);
or U16809 (N_16809,N_15985,N_14170);
or U16810 (N_16810,N_15094,N_14838);
xnor U16811 (N_16811,N_15743,N_14643);
xnor U16812 (N_16812,N_14646,N_15139);
xor U16813 (N_16813,N_15726,N_15587);
or U16814 (N_16814,N_15050,N_15942);
nand U16815 (N_16815,N_14951,N_14343);
nand U16816 (N_16816,N_15374,N_14367);
nand U16817 (N_16817,N_14701,N_14532);
and U16818 (N_16818,N_15140,N_14144);
nor U16819 (N_16819,N_14813,N_14606);
or U16820 (N_16820,N_15953,N_14094);
nand U16821 (N_16821,N_14314,N_14480);
or U16822 (N_16822,N_14142,N_14761);
nand U16823 (N_16823,N_15976,N_14215);
or U16824 (N_16824,N_15036,N_14340);
nand U16825 (N_16825,N_15097,N_15861);
and U16826 (N_16826,N_15687,N_14089);
or U16827 (N_16827,N_14802,N_14884);
and U16828 (N_16828,N_15439,N_14867);
xnor U16829 (N_16829,N_14285,N_15397);
nand U16830 (N_16830,N_14840,N_15033);
xor U16831 (N_16831,N_15496,N_14276);
nand U16832 (N_16832,N_14274,N_15680);
nand U16833 (N_16833,N_15367,N_15885);
nand U16834 (N_16834,N_14180,N_14002);
and U16835 (N_16835,N_15859,N_14588);
nand U16836 (N_16836,N_14674,N_14130);
or U16837 (N_16837,N_14519,N_14676);
and U16838 (N_16838,N_15622,N_15194);
xnor U16839 (N_16839,N_14189,N_14542);
nand U16840 (N_16840,N_14372,N_15035);
xnor U16841 (N_16841,N_14349,N_15225);
and U16842 (N_16842,N_14534,N_15109);
and U16843 (N_16843,N_14978,N_15205);
and U16844 (N_16844,N_15275,N_15688);
or U16845 (N_16845,N_14576,N_14304);
nand U16846 (N_16846,N_15185,N_15719);
or U16847 (N_16847,N_15513,N_14634);
or U16848 (N_16848,N_15423,N_15420);
or U16849 (N_16849,N_14879,N_14776);
xor U16850 (N_16850,N_15470,N_14020);
nor U16851 (N_16851,N_14060,N_14246);
xor U16852 (N_16852,N_14955,N_15251);
or U16853 (N_16853,N_15519,N_15848);
and U16854 (N_16854,N_14686,N_14442);
or U16855 (N_16855,N_14353,N_15464);
or U16856 (N_16856,N_15887,N_14982);
or U16857 (N_16857,N_14136,N_15584);
xnor U16858 (N_16858,N_15963,N_15203);
or U16859 (N_16859,N_14017,N_15949);
nand U16860 (N_16860,N_15749,N_14574);
nand U16861 (N_16861,N_14375,N_14197);
and U16862 (N_16862,N_15505,N_15130);
nor U16863 (N_16863,N_15968,N_14837);
nand U16864 (N_16864,N_15982,N_14704);
xor U16865 (N_16865,N_14059,N_15261);
nand U16866 (N_16866,N_14403,N_15560);
xnor U16867 (N_16867,N_14125,N_15894);
or U16868 (N_16868,N_14530,N_14603);
xor U16869 (N_16869,N_15657,N_15843);
nand U16870 (N_16870,N_14344,N_14479);
nand U16871 (N_16871,N_15804,N_15028);
nand U16872 (N_16872,N_14326,N_14716);
xor U16873 (N_16873,N_14483,N_15810);
nand U16874 (N_16874,N_15043,N_15880);
nor U16875 (N_16875,N_14809,N_14485);
and U16876 (N_16876,N_14556,N_15473);
xor U16877 (N_16877,N_15685,N_15015);
nor U16878 (N_16878,N_14931,N_14315);
and U16879 (N_16879,N_15450,N_14457);
nand U16880 (N_16880,N_14482,N_14300);
or U16881 (N_16881,N_15480,N_14870);
nor U16882 (N_16882,N_15228,N_15409);
or U16883 (N_16883,N_15058,N_14119);
xnor U16884 (N_16884,N_15272,N_15366);
nand U16885 (N_16885,N_14915,N_14971);
xor U16886 (N_16886,N_14021,N_14007);
nand U16887 (N_16887,N_15279,N_15957);
or U16888 (N_16888,N_14427,N_14192);
xnor U16889 (N_16889,N_15491,N_14376);
nand U16890 (N_16890,N_14564,N_15744);
xnor U16891 (N_16891,N_14407,N_15869);
nor U16892 (N_16892,N_15892,N_14598);
or U16893 (N_16893,N_15822,N_14697);
or U16894 (N_16894,N_15218,N_14736);
xor U16895 (N_16895,N_14306,N_14350);
nor U16896 (N_16896,N_14822,N_15750);
xor U16897 (N_16897,N_15451,N_15267);
and U16898 (N_16898,N_15342,N_14387);
nand U16899 (N_16899,N_15943,N_15405);
xor U16900 (N_16900,N_15322,N_14249);
and U16901 (N_16901,N_14975,N_14018);
nor U16902 (N_16902,N_15391,N_15715);
or U16903 (N_16903,N_14608,N_14087);
xnor U16904 (N_16904,N_14735,N_14823);
or U16905 (N_16905,N_15356,N_15987);
or U16906 (N_16906,N_15437,N_14102);
nand U16907 (N_16907,N_14254,N_14680);
and U16908 (N_16908,N_14906,N_14188);
nor U16909 (N_16909,N_15862,N_15167);
nand U16910 (N_16910,N_15054,N_15546);
nand U16911 (N_16911,N_14265,N_14049);
xnor U16912 (N_16912,N_14790,N_14818);
nand U16913 (N_16913,N_14084,N_14032);
and U16914 (N_16914,N_15910,N_14311);
xor U16915 (N_16915,N_14083,N_14677);
nor U16916 (N_16916,N_14993,N_15520);
xnor U16917 (N_16917,N_14212,N_14208);
nor U16918 (N_16918,N_15355,N_15846);
xor U16919 (N_16919,N_14453,N_15684);
nand U16920 (N_16920,N_15727,N_14472);
xnor U16921 (N_16921,N_14568,N_15765);
and U16922 (N_16922,N_15179,N_15651);
or U16923 (N_16923,N_15425,N_14548);
xor U16924 (N_16924,N_15463,N_14890);
or U16925 (N_16925,N_15576,N_14514);
nand U16926 (N_16926,N_14495,N_14159);
or U16927 (N_16927,N_14923,N_14361);
nor U16928 (N_16928,N_15766,N_15124);
nand U16929 (N_16929,N_14998,N_14851);
nand U16930 (N_16930,N_14907,N_15888);
and U16931 (N_16931,N_15911,N_15142);
nand U16932 (N_16932,N_14499,N_14465);
xnor U16933 (N_16933,N_15123,N_14221);
nor U16934 (N_16934,N_15127,N_14445);
xor U16935 (N_16935,N_15613,N_15166);
nor U16936 (N_16936,N_15689,N_14047);
or U16937 (N_16937,N_14042,N_14575);
nor U16938 (N_16938,N_14617,N_15184);
nand U16939 (N_16939,N_15331,N_15206);
nor U16940 (N_16940,N_15600,N_14902);
xnor U16941 (N_16941,N_15604,N_15348);
nand U16942 (N_16942,N_15829,N_15673);
and U16943 (N_16943,N_14671,N_14043);
xor U16944 (N_16944,N_14351,N_14230);
xnor U16945 (N_16945,N_14909,N_15352);
and U16946 (N_16946,N_15489,N_15580);
xnor U16947 (N_16947,N_15896,N_15828);
nor U16948 (N_16948,N_14135,N_14268);
or U16949 (N_16949,N_14449,N_15438);
and U16950 (N_16950,N_14322,N_15556);
or U16951 (N_16951,N_14922,N_14339);
or U16952 (N_16952,N_14477,N_14302);
or U16953 (N_16953,N_15111,N_15961);
or U16954 (N_16954,N_14628,N_14772);
and U16955 (N_16955,N_15823,N_14929);
xor U16956 (N_16956,N_15523,N_14684);
or U16957 (N_16957,N_15216,N_15290);
and U16958 (N_16958,N_14739,N_15619);
and U16959 (N_16959,N_14185,N_15159);
xor U16960 (N_16960,N_15007,N_14370);
and U16961 (N_16961,N_15336,N_15724);
nor U16962 (N_16962,N_14334,N_15503);
or U16963 (N_16963,N_14722,N_14852);
nor U16964 (N_16964,N_14354,N_15096);
xnor U16965 (N_16965,N_14760,N_14899);
nand U16966 (N_16966,N_14401,N_14535);
nor U16967 (N_16967,N_15213,N_14108);
or U16968 (N_16968,N_14076,N_15577);
nand U16969 (N_16969,N_14700,N_15187);
nor U16970 (N_16970,N_15816,N_15024);
or U16971 (N_16971,N_14650,N_14487);
and U16972 (N_16972,N_15311,N_14871);
and U16973 (N_16973,N_14921,N_15596);
or U16974 (N_16974,N_14814,N_14843);
and U16975 (N_16975,N_15854,N_15485);
and U16976 (N_16976,N_15747,N_14481);
and U16977 (N_16977,N_15330,N_14969);
or U16978 (N_16978,N_15066,N_14855);
or U16979 (N_16979,N_14712,N_15797);
xor U16980 (N_16980,N_15590,N_14713);
nor U16981 (N_16981,N_14182,N_15562);
or U16982 (N_16982,N_15121,N_15676);
or U16983 (N_16983,N_15682,N_15006);
xor U16984 (N_16984,N_14428,N_15699);
nand U16985 (N_16985,N_15877,N_14794);
nor U16986 (N_16986,N_14295,N_15484);
and U16987 (N_16987,N_15664,N_15934);
nor U16988 (N_16988,N_15812,N_15244);
or U16989 (N_16989,N_15540,N_14138);
xor U16990 (N_16990,N_14521,N_15558);
nand U16991 (N_16991,N_14336,N_14452);
or U16992 (N_16992,N_15597,N_14236);
nor U16993 (N_16993,N_14571,N_15548);
and U16994 (N_16994,N_15842,N_15241);
nor U16995 (N_16995,N_14359,N_14788);
nand U16996 (N_16996,N_14889,N_14952);
nand U16997 (N_16997,N_14622,N_15363);
nand U16998 (N_16998,N_15561,N_14438);
and U16999 (N_16999,N_14422,N_14204);
xor U17000 (N_17000,N_14684,N_15231);
xnor U17001 (N_17001,N_14359,N_15874);
xor U17002 (N_17002,N_15297,N_15745);
xnor U17003 (N_17003,N_14362,N_14020);
and U17004 (N_17004,N_14502,N_15445);
and U17005 (N_17005,N_15720,N_15426);
nor U17006 (N_17006,N_14345,N_14185);
nor U17007 (N_17007,N_14288,N_15459);
nor U17008 (N_17008,N_15813,N_15197);
or U17009 (N_17009,N_15282,N_15073);
and U17010 (N_17010,N_15552,N_15551);
or U17011 (N_17011,N_15995,N_15964);
or U17012 (N_17012,N_15502,N_14480);
or U17013 (N_17013,N_15409,N_14618);
and U17014 (N_17014,N_15470,N_14584);
nand U17015 (N_17015,N_14543,N_14442);
nor U17016 (N_17016,N_14881,N_14987);
nor U17017 (N_17017,N_15914,N_15855);
and U17018 (N_17018,N_15119,N_15095);
nand U17019 (N_17019,N_14933,N_14239);
and U17020 (N_17020,N_15029,N_14928);
and U17021 (N_17021,N_15748,N_14130);
nand U17022 (N_17022,N_14614,N_15597);
or U17023 (N_17023,N_14079,N_14061);
nand U17024 (N_17024,N_14259,N_15383);
nor U17025 (N_17025,N_15839,N_14951);
nand U17026 (N_17026,N_14783,N_15568);
or U17027 (N_17027,N_14470,N_15824);
nand U17028 (N_17028,N_14670,N_15389);
xnor U17029 (N_17029,N_15151,N_15155);
and U17030 (N_17030,N_14635,N_14427);
xnor U17031 (N_17031,N_15740,N_15367);
xor U17032 (N_17032,N_14140,N_14075);
and U17033 (N_17033,N_14266,N_14155);
nor U17034 (N_17034,N_15903,N_14023);
or U17035 (N_17035,N_14101,N_14755);
nand U17036 (N_17036,N_14224,N_14717);
nand U17037 (N_17037,N_15680,N_14938);
nor U17038 (N_17038,N_15352,N_14211);
nand U17039 (N_17039,N_15586,N_14702);
nor U17040 (N_17040,N_15391,N_15018);
xnor U17041 (N_17041,N_15191,N_14927);
nor U17042 (N_17042,N_15254,N_15691);
nand U17043 (N_17043,N_15403,N_15301);
xor U17044 (N_17044,N_15995,N_15386);
nor U17045 (N_17045,N_14929,N_14855);
or U17046 (N_17046,N_14107,N_14689);
and U17047 (N_17047,N_15468,N_15130);
xor U17048 (N_17048,N_15026,N_14739);
and U17049 (N_17049,N_14485,N_14185);
xor U17050 (N_17050,N_15573,N_14638);
nor U17051 (N_17051,N_15173,N_14267);
nor U17052 (N_17052,N_14321,N_15111);
xor U17053 (N_17053,N_15042,N_14656);
xor U17054 (N_17054,N_15181,N_15340);
nand U17055 (N_17055,N_15300,N_15912);
xnor U17056 (N_17056,N_15033,N_15508);
and U17057 (N_17057,N_14270,N_14498);
and U17058 (N_17058,N_14651,N_15073);
or U17059 (N_17059,N_15361,N_15962);
xnor U17060 (N_17060,N_15857,N_15818);
nor U17061 (N_17061,N_15198,N_14112);
and U17062 (N_17062,N_14440,N_15466);
nor U17063 (N_17063,N_14552,N_15710);
and U17064 (N_17064,N_14184,N_15675);
xnor U17065 (N_17065,N_15413,N_15995);
nand U17066 (N_17066,N_15310,N_14208);
xnor U17067 (N_17067,N_15069,N_14504);
and U17068 (N_17068,N_14190,N_15180);
nor U17069 (N_17069,N_14743,N_15193);
nand U17070 (N_17070,N_15035,N_14720);
xor U17071 (N_17071,N_15761,N_14578);
nand U17072 (N_17072,N_15852,N_14315);
or U17073 (N_17073,N_14647,N_14195);
and U17074 (N_17074,N_15744,N_15109);
and U17075 (N_17075,N_15931,N_15530);
and U17076 (N_17076,N_15484,N_14826);
xnor U17077 (N_17077,N_14480,N_14704);
and U17078 (N_17078,N_14515,N_15392);
xnor U17079 (N_17079,N_15444,N_14058);
nand U17080 (N_17080,N_14050,N_14287);
and U17081 (N_17081,N_14291,N_14230);
nand U17082 (N_17082,N_15903,N_14440);
or U17083 (N_17083,N_14510,N_14610);
nand U17084 (N_17084,N_14232,N_14617);
xor U17085 (N_17085,N_14208,N_15280);
nor U17086 (N_17086,N_15935,N_14505);
nand U17087 (N_17087,N_14005,N_14286);
nand U17088 (N_17088,N_14619,N_14833);
nand U17089 (N_17089,N_14594,N_14707);
xor U17090 (N_17090,N_14595,N_14895);
nand U17091 (N_17091,N_14133,N_15968);
nor U17092 (N_17092,N_14427,N_14057);
and U17093 (N_17093,N_15452,N_14959);
nor U17094 (N_17094,N_15738,N_15490);
xnor U17095 (N_17095,N_15027,N_15155);
xnor U17096 (N_17096,N_14268,N_15791);
nor U17097 (N_17097,N_14843,N_15724);
nand U17098 (N_17098,N_14229,N_14891);
and U17099 (N_17099,N_14542,N_15318);
xnor U17100 (N_17100,N_14652,N_15931);
nand U17101 (N_17101,N_14955,N_15365);
nor U17102 (N_17102,N_15582,N_14282);
nand U17103 (N_17103,N_15263,N_14583);
nor U17104 (N_17104,N_14570,N_14111);
nor U17105 (N_17105,N_14194,N_15980);
and U17106 (N_17106,N_15415,N_15088);
nor U17107 (N_17107,N_14603,N_14646);
nor U17108 (N_17108,N_14588,N_14930);
nand U17109 (N_17109,N_15475,N_15739);
or U17110 (N_17110,N_15941,N_15853);
xnor U17111 (N_17111,N_14237,N_15569);
and U17112 (N_17112,N_15839,N_14538);
nor U17113 (N_17113,N_14791,N_15244);
nor U17114 (N_17114,N_14848,N_14612);
xnor U17115 (N_17115,N_14359,N_15640);
nand U17116 (N_17116,N_15906,N_14552);
nand U17117 (N_17117,N_15795,N_14350);
nand U17118 (N_17118,N_15834,N_15439);
nand U17119 (N_17119,N_15843,N_14049);
xor U17120 (N_17120,N_15498,N_15817);
and U17121 (N_17121,N_15700,N_14174);
nand U17122 (N_17122,N_15025,N_14998);
or U17123 (N_17123,N_14010,N_14655);
nor U17124 (N_17124,N_15036,N_15297);
nand U17125 (N_17125,N_14505,N_14267);
and U17126 (N_17126,N_14413,N_15097);
and U17127 (N_17127,N_14416,N_15770);
xnor U17128 (N_17128,N_15598,N_14603);
xor U17129 (N_17129,N_14688,N_15389);
xor U17130 (N_17130,N_15117,N_14329);
xor U17131 (N_17131,N_15041,N_15767);
nand U17132 (N_17132,N_14926,N_15276);
nand U17133 (N_17133,N_14796,N_15519);
or U17134 (N_17134,N_15533,N_14029);
nand U17135 (N_17135,N_15210,N_14708);
nor U17136 (N_17136,N_14622,N_14011);
nand U17137 (N_17137,N_15719,N_15560);
xnor U17138 (N_17138,N_15492,N_14907);
or U17139 (N_17139,N_14829,N_15017);
nand U17140 (N_17140,N_15400,N_15173);
nor U17141 (N_17141,N_14399,N_15728);
and U17142 (N_17142,N_15980,N_14629);
or U17143 (N_17143,N_15765,N_15020);
or U17144 (N_17144,N_14466,N_14440);
and U17145 (N_17145,N_15710,N_15256);
nand U17146 (N_17146,N_15267,N_14494);
or U17147 (N_17147,N_14322,N_14690);
and U17148 (N_17148,N_15449,N_14054);
nor U17149 (N_17149,N_15256,N_15864);
nand U17150 (N_17150,N_15725,N_15399);
or U17151 (N_17151,N_15325,N_15625);
and U17152 (N_17152,N_15445,N_15894);
or U17153 (N_17153,N_14117,N_15249);
or U17154 (N_17154,N_14724,N_14261);
nor U17155 (N_17155,N_14182,N_14856);
or U17156 (N_17156,N_15715,N_14262);
nand U17157 (N_17157,N_14699,N_15868);
or U17158 (N_17158,N_14259,N_15524);
nand U17159 (N_17159,N_14187,N_15029);
nor U17160 (N_17160,N_14814,N_15185);
and U17161 (N_17161,N_15972,N_14797);
xor U17162 (N_17162,N_14406,N_15706);
xnor U17163 (N_17163,N_14997,N_14097);
nand U17164 (N_17164,N_14887,N_15903);
or U17165 (N_17165,N_15882,N_14117);
or U17166 (N_17166,N_14065,N_15239);
xnor U17167 (N_17167,N_15275,N_15239);
and U17168 (N_17168,N_15774,N_15330);
and U17169 (N_17169,N_14222,N_15054);
nand U17170 (N_17170,N_14148,N_15046);
and U17171 (N_17171,N_15924,N_15184);
xor U17172 (N_17172,N_15005,N_14212);
xor U17173 (N_17173,N_15142,N_15151);
and U17174 (N_17174,N_14380,N_14143);
and U17175 (N_17175,N_15280,N_15927);
or U17176 (N_17176,N_15539,N_15171);
xnor U17177 (N_17177,N_15364,N_15903);
nor U17178 (N_17178,N_14613,N_14332);
or U17179 (N_17179,N_15596,N_14134);
nand U17180 (N_17180,N_15288,N_15882);
or U17181 (N_17181,N_14264,N_14727);
nand U17182 (N_17182,N_14619,N_14045);
xor U17183 (N_17183,N_14559,N_14471);
xnor U17184 (N_17184,N_14283,N_15204);
nand U17185 (N_17185,N_15510,N_14528);
and U17186 (N_17186,N_15389,N_15348);
or U17187 (N_17187,N_14737,N_14767);
or U17188 (N_17188,N_15021,N_15544);
and U17189 (N_17189,N_15167,N_15090);
nor U17190 (N_17190,N_14277,N_14712);
xnor U17191 (N_17191,N_14523,N_15090);
nor U17192 (N_17192,N_15236,N_14191);
nor U17193 (N_17193,N_15315,N_14151);
nand U17194 (N_17194,N_14636,N_15343);
nor U17195 (N_17195,N_15749,N_14047);
and U17196 (N_17196,N_14624,N_14294);
nor U17197 (N_17197,N_15091,N_15332);
xor U17198 (N_17198,N_14857,N_15520);
xnor U17199 (N_17199,N_15274,N_14791);
nand U17200 (N_17200,N_14116,N_14077);
nand U17201 (N_17201,N_15555,N_15059);
nand U17202 (N_17202,N_14271,N_14096);
nor U17203 (N_17203,N_15834,N_14696);
or U17204 (N_17204,N_15899,N_14012);
nand U17205 (N_17205,N_14222,N_15861);
and U17206 (N_17206,N_14012,N_14239);
nor U17207 (N_17207,N_15581,N_14714);
and U17208 (N_17208,N_14256,N_15513);
or U17209 (N_17209,N_14041,N_15417);
and U17210 (N_17210,N_15323,N_15417);
and U17211 (N_17211,N_14491,N_14359);
or U17212 (N_17212,N_14826,N_15674);
nand U17213 (N_17213,N_14414,N_14111);
xor U17214 (N_17214,N_15245,N_14704);
nor U17215 (N_17215,N_15041,N_15430);
or U17216 (N_17216,N_14148,N_14269);
nor U17217 (N_17217,N_14341,N_14163);
nand U17218 (N_17218,N_14420,N_14603);
and U17219 (N_17219,N_15907,N_14949);
nand U17220 (N_17220,N_14649,N_14091);
and U17221 (N_17221,N_14131,N_14677);
xor U17222 (N_17222,N_14199,N_14281);
xor U17223 (N_17223,N_14231,N_14661);
or U17224 (N_17224,N_14718,N_14324);
nor U17225 (N_17225,N_14252,N_15608);
and U17226 (N_17226,N_14961,N_14633);
xnor U17227 (N_17227,N_14180,N_14865);
nand U17228 (N_17228,N_14476,N_15730);
xnor U17229 (N_17229,N_15003,N_14285);
nand U17230 (N_17230,N_14993,N_14697);
nor U17231 (N_17231,N_15098,N_15253);
xnor U17232 (N_17232,N_15720,N_14619);
and U17233 (N_17233,N_15673,N_15090);
and U17234 (N_17234,N_15616,N_14436);
or U17235 (N_17235,N_15428,N_14680);
and U17236 (N_17236,N_14232,N_14678);
or U17237 (N_17237,N_14513,N_14511);
nand U17238 (N_17238,N_14972,N_15034);
and U17239 (N_17239,N_15839,N_15975);
and U17240 (N_17240,N_15159,N_15806);
xnor U17241 (N_17241,N_14875,N_15140);
or U17242 (N_17242,N_14869,N_15567);
xnor U17243 (N_17243,N_15992,N_14533);
nor U17244 (N_17244,N_15274,N_15374);
nor U17245 (N_17245,N_15696,N_14710);
nand U17246 (N_17246,N_14285,N_15534);
and U17247 (N_17247,N_14497,N_15356);
xor U17248 (N_17248,N_14233,N_14828);
or U17249 (N_17249,N_14111,N_14475);
nand U17250 (N_17250,N_14074,N_14941);
xor U17251 (N_17251,N_14120,N_14728);
or U17252 (N_17252,N_14693,N_14067);
nand U17253 (N_17253,N_15900,N_14280);
xnor U17254 (N_17254,N_15883,N_15421);
xnor U17255 (N_17255,N_15837,N_14391);
nor U17256 (N_17256,N_15303,N_15500);
xor U17257 (N_17257,N_14629,N_14462);
nor U17258 (N_17258,N_14280,N_15352);
and U17259 (N_17259,N_15633,N_15305);
xor U17260 (N_17260,N_15459,N_14928);
and U17261 (N_17261,N_14816,N_15250);
nand U17262 (N_17262,N_14485,N_14786);
nor U17263 (N_17263,N_14591,N_14660);
and U17264 (N_17264,N_14982,N_14148);
xor U17265 (N_17265,N_14219,N_15277);
and U17266 (N_17266,N_14657,N_14175);
and U17267 (N_17267,N_14855,N_15645);
nor U17268 (N_17268,N_14476,N_14964);
nand U17269 (N_17269,N_15504,N_15461);
or U17270 (N_17270,N_14848,N_15305);
or U17271 (N_17271,N_15784,N_15081);
nand U17272 (N_17272,N_15095,N_15142);
nor U17273 (N_17273,N_14842,N_15255);
and U17274 (N_17274,N_15387,N_14086);
xor U17275 (N_17275,N_14488,N_14112);
nand U17276 (N_17276,N_14357,N_15909);
and U17277 (N_17277,N_14113,N_15387);
and U17278 (N_17278,N_14120,N_15682);
nor U17279 (N_17279,N_14359,N_14522);
and U17280 (N_17280,N_14035,N_15593);
nand U17281 (N_17281,N_15803,N_15681);
xor U17282 (N_17282,N_14312,N_14369);
and U17283 (N_17283,N_15879,N_15435);
nor U17284 (N_17284,N_14985,N_15145);
and U17285 (N_17285,N_15585,N_14814);
nand U17286 (N_17286,N_14863,N_15718);
or U17287 (N_17287,N_14446,N_14034);
and U17288 (N_17288,N_15545,N_15071);
xnor U17289 (N_17289,N_15729,N_15588);
or U17290 (N_17290,N_14577,N_14402);
nand U17291 (N_17291,N_14295,N_15078);
nor U17292 (N_17292,N_15179,N_15693);
or U17293 (N_17293,N_14008,N_14791);
and U17294 (N_17294,N_15869,N_14092);
nand U17295 (N_17295,N_15822,N_15830);
xnor U17296 (N_17296,N_15692,N_15154);
nor U17297 (N_17297,N_14221,N_14375);
and U17298 (N_17298,N_15334,N_14376);
nor U17299 (N_17299,N_14671,N_14009);
nand U17300 (N_17300,N_15117,N_15219);
nor U17301 (N_17301,N_14696,N_15745);
and U17302 (N_17302,N_14075,N_14583);
nand U17303 (N_17303,N_14428,N_14913);
and U17304 (N_17304,N_14543,N_15101);
nand U17305 (N_17305,N_14944,N_14029);
xor U17306 (N_17306,N_15597,N_15840);
or U17307 (N_17307,N_14356,N_15771);
or U17308 (N_17308,N_14620,N_14362);
nand U17309 (N_17309,N_14909,N_14414);
and U17310 (N_17310,N_14971,N_14401);
nor U17311 (N_17311,N_14917,N_15577);
nor U17312 (N_17312,N_15703,N_14923);
or U17313 (N_17313,N_15654,N_14173);
or U17314 (N_17314,N_15591,N_14890);
xor U17315 (N_17315,N_15043,N_15182);
nand U17316 (N_17316,N_14131,N_15748);
and U17317 (N_17317,N_14018,N_15706);
or U17318 (N_17318,N_15144,N_14584);
xnor U17319 (N_17319,N_15260,N_14525);
and U17320 (N_17320,N_14099,N_15170);
xnor U17321 (N_17321,N_15448,N_14350);
nand U17322 (N_17322,N_15151,N_14066);
nor U17323 (N_17323,N_15441,N_15064);
or U17324 (N_17324,N_14318,N_14379);
nand U17325 (N_17325,N_15399,N_14102);
or U17326 (N_17326,N_14295,N_15530);
xnor U17327 (N_17327,N_15722,N_14105);
nand U17328 (N_17328,N_15356,N_14649);
and U17329 (N_17329,N_14784,N_15904);
and U17330 (N_17330,N_15626,N_14290);
nand U17331 (N_17331,N_15302,N_15140);
nand U17332 (N_17332,N_14104,N_14377);
xnor U17333 (N_17333,N_15730,N_14789);
and U17334 (N_17334,N_15143,N_14395);
nand U17335 (N_17335,N_14544,N_15687);
or U17336 (N_17336,N_15534,N_15685);
nand U17337 (N_17337,N_14687,N_15304);
or U17338 (N_17338,N_14272,N_15630);
or U17339 (N_17339,N_14366,N_14303);
nand U17340 (N_17340,N_15418,N_14581);
and U17341 (N_17341,N_15906,N_14430);
xnor U17342 (N_17342,N_14502,N_15120);
xnor U17343 (N_17343,N_14262,N_15099);
xnor U17344 (N_17344,N_15652,N_14057);
nand U17345 (N_17345,N_14033,N_15309);
nor U17346 (N_17346,N_14963,N_15929);
xor U17347 (N_17347,N_15442,N_14948);
nor U17348 (N_17348,N_15649,N_15415);
nor U17349 (N_17349,N_14753,N_15476);
nor U17350 (N_17350,N_15997,N_14140);
nand U17351 (N_17351,N_14881,N_15840);
nor U17352 (N_17352,N_14515,N_14788);
or U17353 (N_17353,N_14357,N_14922);
nor U17354 (N_17354,N_14893,N_15616);
nor U17355 (N_17355,N_15167,N_15074);
and U17356 (N_17356,N_15951,N_14910);
nor U17357 (N_17357,N_14265,N_15475);
nor U17358 (N_17358,N_15017,N_15289);
xnor U17359 (N_17359,N_14465,N_15679);
and U17360 (N_17360,N_14402,N_14576);
nand U17361 (N_17361,N_15171,N_15475);
and U17362 (N_17362,N_14175,N_15100);
nor U17363 (N_17363,N_14254,N_15213);
or U17364 (N_17364,N_15018,N_15773);
xnor U17365 (N_17365,N_14696,N_14544);
nand U17366 (N_17366,N_15745,N_14795);
nand U17367 (N_17367,N_14760,N_15277);
or U17368 (N_17368,N_15323,N_14638);
nor U17369 (N_17369,N_14858,N_15952);
and U17370 (N_17370,N_15911,N_15199);
nand U17371 (N_17371,N_15206,N_14964);
and U17372 (N_17372,N_14670,N_15160);
nor U17373 (N_17373,N_15241,N_15209);
nor U17374 (N_17374,N_15389,N_14278);
or U17375 (N_17375,N_14136,N_15581);
nand U17376 (N_17376,N_15773,N_15233);
nand U17377 (N_17377,N_15414,N_14746);
and U17378 (N_17378,N_14514,N_15227);
and U17379 (N_17379,N_15950,N_15627);
nand U17380 (N_17380,N_14082,N_15621);
nand U17381 (N_17381,N_15483,N_15933);
nand U17382 (N_17382,N_15502,N_15318);
and U17383 (N_17383,N_15322,N_14848);
and U17384 (N_17384,N_14888,N_14099);
nor U17385 (N_17385,N_15357,N_15625);
or U17386 (N_17386,N_15933,N_14372);
nor U17387 (N_17387,N_15429,N_15970);
xor U17388 (N_17388,N_15365,N_14270);
or U17389 (N_17389,N_14287,N_15563);
and U17390 (N_17390,N_15008,N_14978);
nor U17391 (N_17391,N_15541,N_14555);
nor U17392 (N_17392,N_15166,N_14482);
or U17393 (N_17393,N_14853,N_14656);
or U17394 (N_17394,N_14861,N_15343);
xor U17395 (N_17395,N_15653,N_15785);
nand U17396 (N_17396,N_15520,N_14835);
and U17397 (N_17397,N_14681,N_14294);
or U17398 (N_17398,N_14319,N_15995);
nand U17399 (N_17399,N_14990,N_15415);
nand U17400 (N_17400,N_15449,N_15275);
nor U17401 (N_17401,N_15915,N_14271);
and U17402 (N_17402,N_15760,N_14567);
nand U17403 (N_17403,N_14996,N_14289);
nand U17404 (N_17404,N_15529,N_14061);
and U17405 (N_17405,N_14391,N_15404);
nor U17406 (N_17406,N_15516,N_14522);
nand U17407 (N_17407,N_14324,N_14789);
or U17408 (N_17408,N_15348,N_14123);
or U17409 (N_17409,N_15132,N_15316);
nor U17410 (N_17410,N_15645,N_15841);
xnor U17411 (N_17411,N_15182,N_14958);
nor U17412 (N_17412,N_14146,N_14926);
nand U17413 (N_17413,N_15375,N_14047);
and U17414 (N_17414,N_15697,N_15880);
nor U17415 (N_17415,N_15073,N_15908);
nand U17416 (N_17416,N_15288,N_15890);
nand U17417 (N_17417,N_14985,N_14706);
nand U17418 (N_17418,N_15456,N_14763);
nand U17419 (N_17419,N_14468,N_15829);
or U17420 (N_17420,N_15709,N_14646);
xor U17421 (N_17421,N_14285,N_15905);
nand U17422 (N_17422,N_15557,N_15034);
and U17423 (N_17423,N_15771,N_14760);
and U17424 (N_17424,N_15454,N_15216);
nor U17425 (N_17425,N_15543,N_15044);
nand U17426 (N_17426,N_14081,N_15709);
and U17427 (N_17427,N_14576,N_14392);
and U17428 (N_17428,N_14659,N_14624);
nand U17429 (N_17429,N_14559,N_14402);
xor U17430 (N_17430,N_14107,N_15183);
and U17431 (N_17431,N_15573,N_15291);
and U17432 (N_17432,N_14020,N_14622);
or U17433 (N_17433,N_14570,N_15808);
nand U17434 (N_17434,N_14739,N_15237);
xor U17435 (N_17435,N_14718,N_14610);
and U17436 (N_17436,N_14483,N_14612);
and U17437 (N_17437,N_14353,N_15288);
or U17438 (N_17438,N_15744,N_14806);
and U17439 (N_17439,N_15812,N_15174);
or U17440 (N_17440,N_15471,N_15124);
nand U17441 (N_17441,N_14771,N_14741);
nor U17442 (N_17442,N_15119,N_14536);
or U17443 (N_17443,N_14606,N_14237);
and U17444 (N_17444,N_15972,N_14391);
and U17445 (N_17445,N_14661,N_14471);
and U17446 (N_17446,N_14289,N_15917);
xnor U17447 (N_17447,N_14780,N_15225);
and U17448 (N_17448,N_14821,N_14748);
and U17449 (N_17449,N_14801,N_15639);
or U17450 (N_17450,N_14820,N_15803);
and U17451 (N_17451,N_15583,N_15357);
or U17452 (N_17452,N_15429,N_14103);
xor U17453 (N_17453,N_14402,N_15179);
nor U17454 (N_17454,N_14296,N_14808);
nand U17455 (N_17455,N_14650,N_15515);
and U17456 (N_17456,N_15752,N_14787);
or U17457 (N_17457,N_15039,N_14400);
or U17458 (N_17458,N_14526,N_14309);
and U17459 (N_17459,N_15488,N_15042);
nand U17460 (N_17460,N_14526,N_15665);
and U17461 (N_17461,N_14116,N_14618);
and U17462 (N_17462,N_14536,N_14270);
nor U17463 (N_17463,N_14608,N_15880);
nor U17464 (N_17464,N_14024,N_14244);
or U17465 (N_17465,N_14264,N_14382);
nor U17466 (N_17466,N_14325,N_15957);
and U17467 (N_17467,N_14810,N_14492);
or U17468 (N_17468,N_15848,N_15942);
nor U17469 (N_17469,N_14142,N_15904);
nor U17470 (N_17470,N_15155,N_15347);
nor U17471 (N_17471,N_14934,N_14816);
nor U17472 (N_17472,N_15743,N_15407);
or U17473 (N_17473,N_15707,N_15062);
nand U17474 (N_17474,N_15443,N_14479);
and U17475 (N_17475,N_15051,N_15114);
xor U17476 (N_17476,N_14005,N_15106);
nor U17477 (N_17477,N_15119,N_15351);
nand U17478 (N_17478,N_14205,N_14207);
nor U17479 (N_17479,N_15340,N_15611);
xor U17480 (N_17480,N_14643,N_15042);
nor U17481 (N_17481,N_14044,N_14032);
nor U17482 (N_17482,N_15694,N_15659);
and U17483 (N_17483,N_15789,N_15018);
and U17484 (N_17484,N_14668,N_14913);
nor U17485 (N_17485,N_14238,N_14671);
or U17486 (N_17486,N_14113,N_15603);
nor U17487 (N_17487,N_15275,N_14304);
nand U17488 (N_17488,N_15086,N_15707);
nor U17489 (N_17489,N_14563,N_14569);
nand U17490 (N_17490,N_15196,N_15452);
nand U17491 (N_17491,N_14081,N_15456);
or U17492 (N_17492,N_15873,N_14031);
xnor U17493 (N_17493,N_14835,N_14680);
nand U17494 (N_17494,N_15265,N_15626);
nor U17495 (N_17495,N_15963,N_15785);
or U17496 (N_17496,N_14215,N_15862);
nor U17497 (N_17497,N_15843,N_15811);
xor U17498 (N_17498,N_15223,N_15759);
nand U17499 (N_17499,N_14594,N_14172);
xor U17500 (N_17500,N_15108,N_14051);
or U17501 (N_17501,N_14279,N_15670);
xnor U17502 (N_17502,N_14648,N_15612);
xor U17503 (N_17503,N_15709,N_14778);
nand U17504 (N_17504,N_14207,N_14090);
or U17505 (N_17505,N_15270,N_14745);
xor U17506 (N_17506,N_15639,N_14214);
xnor U17507 (N_17507,N_14478,N_15941);
nor U17508 (N_17508,N_14393,N_14387);
nand U17509 (N_17509,N_14456,N_14917);
or U17510 (N_17510,N_15497,N_14600);
and U17511 (N_17511,N_15628,N_14049);
or U17512 (N_17512,N_14877,N_15143);
or U17513 (N_17513,N_14438,N_14022);
nor U17514 (N_17514,N_14508,N_14141);
nand U17515 (N_17515,N_15663,N_15675);
or U17516 (N_17516,N_15091,N_14097);
or U17517 (N_17517,N_15867,N_14837);
or U17518 (N_17518,N_15072,N_15100);
nand U17519 (N_17519,N_14976,N_15416);
nand U17520 (N_17520,N_15036,N_14077);
and U17521 (N_17521,N_15994,N_15039);
nand U17522 (N_17522,N_15700,N_15237);
and U17523 (N_17523,N_14407,N_14018);
or U17524 (N_17524,N_15601,N_15508);
nand U17525 (N_17525,N_15791,N_14331);
nor U17526 (N_17526,N_15389,N_14906);
or U17527 (N_17527,N_15799,N_14998);
nor U17528 (N_17528,N_15700,N_14235);
or U17529 (N_17529,N_14385,N_14735);
nand U17530 (N_17530,N_15647,N_14379);
nand U17531 (N_17531,N_15056,N_15092);
or U17532 (N_17532,N_15997,N_15523);
and U17533 (N_17533,N_15482,N_14905);
nor U17534 (N_17534,N_15182,N_15739);
nand U17535 (N_17535,N_15139,N_15156);
or U17536 (N_17536,N_15714,N_14028);
xor U17537 (N_17537,N_14259,N_15953);
xnor U17538 (N_17538,N_15177,N_14768);
and U17539 (N_17539,N_14815,N_15079);
and U17540 (N_17540,N_14412,N_14481);
nor U17541 (N_17541,N_14463,N_15977);
nand U17542 (N_17542,N_14942,N_15203);
and U17543 (N_17543,N_14496,N_14981);
or U17544 (N_17544,N_15817,N_14442);
or U17545 (N_17545,N_14600,N_14783);
or U17546 (N_17546,N_15255,N_15507);
xor U17547 (N_17547,N_14919,N_15726);
or U17548 (N_17548,N_15246,N_14755);
and U17549 (N_17549,N_15238,N_14413);
xor U17550 (N_17550,N_15889,N_15538);
and U17551 (N_17551,N_14321,N_15598);
and U17552 (N_17552,N_15091,N_15537);
or U17553 (N_17553,N_15773,N_15237);
xor U17554 (N_17554,N_15087,N_14348);
nor U17555 (N_17555,N_15505,N_14930);
and U17556 (N_17556,N_14801,N_14479);
nor U17557 (N_17557,N_14356,N_15582);
nor U17558 (N_17558,N_15559,N_15933);
and U17559 (N_17559,N_15296,N_14027);
xnor U17560 (N_17560,N_14002,N_15192);
nor U17561 (N_17561,N_15507,N_14687);
nand U17562 (N_17562,N_15764,N_15610);
nand U17563 (N_17563,N_15116,N_14293);
nand U17564 (N_17564,N_15746,N_15288);
and U17565 (N_17565,N_15422,N_14525);
nand U17566 (N_17566,N_15462,N_14000);
nand U17567 (N_17567,N_14874,N_14325);
or U17568 (N_17568,N_14211,N_15282);
or U17569 (N_17569,N_14487,N_15973);
and U17570 (N_17570,N_14688,N_14231);
and U17571 (N_17571,N_15807,N_14816);
xor U17572 (N_17572,N_15235,N_14068);
and U17573 (N_17573,N_15447,N_14791);
and U17574 (N_17574,N_15905,N_15653);
nand U17575 (N_17575,N_14246,N_14817);
xor U17576 (N_17576,N_14641,N_15100);
or U17577 (N_17577,N_15645,N_15676);
xor U17578 (N_17578,N_15688,N_14445);
xor U17579 (N_17579,N_14084,N_14428);
and U17580 (N_17580,N_15168,N_14045);
and U17581 (N_17581,N_14112,N_15929);
nor U17582 (N_17582,N_14253,N_14322);
and U17583 (N_17583,N_14214,N_15204);
xnor U17584 (N_17584,N_14743,N_15452);
xnor U17585 (N_17585,N_15890,N_14736);
and U17586 (N_17586,N_15990,N_15342);
nor U17587 (N_17587,N_15798,N_15056);
xnor U17588 (N_17588,N_15667,N_15979);
xor U17589 (N_17589,N_15075,N_14352);
nand U17590 (N_17590,N_15109,N_15924);
nand U17591 (N_17591,N_14971,N_14565);
nand U17592 (N_17592,N_14159,N_14739);
xnor U17593 (N_17593,N_15009,N_14205);
nor U17594 (N_17594,N_15929,N_14337);
nor U17595 (N_17595,N_15832,N_15256);
xnor U17596 (N_17596,N_15636,N_15718);
or U17597 (N_17597,N_14249,N_14020);
and U17598 (N_17598,N_14464,N_15794);
nand U17599 (N_17599,N_15919,N_15817);
nor U17600 (N_17600,N_14791,N_15113);
and U17601 (N_17601,N_15901,N_15702);
nand U17602 (N_17602,N_14712,N_15661);
nand U17603 (N_17603,N_14972,N_14016);
nor U17604 (N_17604,N_15268,N_14130);
or U17605 (N_17605,N_15368,N_14497);
nor U17606 (N_17606,N_14975,N_14548);
or U17607 (N_17607,N_15738,N_15318);
and U17608 (N_17608,N_14483,N_15812);
nand U17609 (N_17609,N_14080,N_15919);
nor U17610 (N_17610,N_14355,N_14559);
nor U17611 (N_17611,N_15953,N_14557);
nor U17612 (N_17612,N_15518,N_14133);
or U17613 (N_17613,N_14763,N_14854);
and U17614 (N_17614,N_14970,N_14570);
and U17615 (N_17615,N_14774,N_14870);
and U17616 (N_17616,N_14691,N_15474);
nand U17617 (N_17617,N_15023,N_15978);
or U17618 (N_17618,N_15494,N_15642);
or U17619 (N_17619,N_15084,N_15078);
and U17620 (N_17620,N_14496,N_15735);
nor U17621 (N_17621,N_15071,N_15582);
xor U17622 (N_17622,N_14114,N_14567);
or U17623 (N_17623,N_14570,N_15426);
xnor U17624 (N_17624,N_15605,N_15244);
or U17625 (N_17625,N_14535,N_15576);
nand U17626 (N_17626,N_14018,N_15771);
nand U17627 (N_17627,N_15085,N_14461);
and U17628 (N_17628,N_14287,N_15592);
nand U17629 (N_17629,N_14802,N_14993);
or U17630 (N_17630,N_14939,N_15542);
and U17631 (N_17631,N_15785,N_15171);
and U17632 (N_17632,N_14398,N_15534);
and U17633 (N_17633,N_14700,N_15508);
nor U17634 (N_17634,N_15512,N_15237);
xnor U17635 (N_17635,N_14372,N_15847);
or U17636 (N_17636,N_14444,N_14901);
xor U17637 (N_17637,N_15953,N_15975);
or U17638 (N_17638,N_15528,N_14496);
or U17639 (N_17639,N_15201,N_15422);
nand U17640 (N_17640,N_14247,N_14169);
and U17641 (N_17641,N_14248,N_14602);
nand U17642 (N_17642,N_14130,N_15428);
or U17643 (N_17643,N_14564,N_14227);
xnor U17644 (N_17644,N_15860,N_14775);
and U17645 (N_17645,N_15243,N_14891);
or U17646 (N_17646,N_14366,N_15940);
and U17647 (N_17647,N_15624,N_15655);
or U17648 (N_17648,N_15225,N_14626);
or U17649 (N_17649,N_14183,N_14630);
nor U17650 (N_17650,N_14323,N_14127);
xor U17651 (N_17651,N_15913,N_14011);
nand U17652 (N_17652,N_14878,N_15219);
or U17653 (N_17653,N_14385,N_14827);
nor U17654 (N_17654,N_14367,N_15501);
nor U17655 (N_17655,N_14178,N_15220);
nor U17656 (N_17656,N_15725,N_15354);
nor U17657 (N_17657,N_15463,N_15883);
and U17658 (N_17658,N_15639,N_15368);
and U17659 (N_17659,N_15727,N_15213);
nor U17660 (N_17660,N_15084,N_14009);
nand U17661 (N_17661,N_14140,N_15921);
xor U17662 (N_17662,N_15431,N_14575);
and U17663 (N_17663,N_14179,N_15758);
or U17664 (N_17664,N_15092,N_15283);
nor U17665 (N_17665,N_14897,N_15780);
or U17666 (N_17666,N_14199,N_15087);
or U17667 (N_17667,N_15336,N_14010);
nor U17668 (N_17668,N_15385,N_15717);
nand U17669 (N_17669,N_15023,N_15459);
and U17670 (N_17670,N_15676,N_14115);
nor U17671 (N_17671,N_14951,N_14931);
nor U17672 (N_17672,N_14573,N_14776);
and U17673 (N_17673,N_15423,N_15951);
or U17674 (N_17674,N_15481,N_15913);
and U17675 (N_17675,N_14296,N_14038);
or U17676 (N_17676,N_14205,N_14148);
and U17677 (N_17677,N_14819,N_15179);
and U17678 (N_17678,N_14183,N_15367);
and U17679 (N_17679,N_15871,N_14123);
nor U17680 (N_17680,N_15024,N_14895);
nand U17681 (N_17681,N_14589,N_15168);
nor U17682 (N_17682,N_15891,N_15210);
nand U17683 (N_17683,N_14277,N_15637);
nor U17684 (N_17684,N_14752,N_15974);
xnor U17685 (N_17685,N_15023,N_14756);
or U17686 (N_17686,N_14318,N_14770);
xor U17687 (N_17687,N_14425,N_14055);
or U17688 (N_17688,N_14535,N_14532);
nand U17689 (N_17689,N_14340,N_14215);
nand U17690 (N_17690,N_14931,N_14902);
and U17691 (N_17691,N_15080,N_14389);
nand U17692 (N_17692,N_14992,N_14658);
or U17693 (N_17693,N_15810,N_14433);
and U17694 (N_17694,N_15912,N_15507);
and U17695 (N_17695,N_15283,N_15629);
nand U17696 (N_17696,N_15848,N_15107);
nand U17697 (N_17697,N_14486,N_14467);
and U17698 (N_17698,N_15031,N_15271);
or U17699 (N_17699,N_15443,N_14001);
and U17700 (N_17700,N_14582,N_14705);
nor U17701 (N_17701,N_15017,N_14838);
xor U17702 (N_17702,N_14700,N_14622);
nand U17703 (N_17703,N_14818,N_14903);
xnor U17704 (N_17704,N_15001,N_14175);
xnor U17705 (N_17705,N_15710,N_14245);
xor U17706 (N_17706,N_14259,N_15527);
or U17707 (N_17707,N_15721,N_15505);
nand U17708 (N_17708,N_14078,N_15946);
nand U17709 (N_17709,N_14275,N_14833);
nor U17710 (N_17710,N_15273,N_14677);
xnor U17711 (N_17711,N_15877,N_14434);
and U17712 (N_17712,N_15591,N_14874);
nor U17713 (N_17713,N_14126,N_15078);
nand U17714 (N_17714,N_14793,N_14676);
and U17715 (N_17715,N_15452,N_14649);
xnor U17716 (N_17716,N_14414,N_14666);
xor U17717 (N_17717,N_14758,N_14777);
or U17718 (N_17718,N_14742,N_14335);
nand U17719 (N_17719,N_15996,N_15751);
or U17720 (N_17720,N_15354,N_14015);
nor U17721 (N_17721,N_14474,N_14685);
xnor U17722 (N_17722,N_15471,N_15801);
nand U17723 (N_17723,N_14454,N_15474);
or U17724 (N_17724,N_15016,N_15494);
xnor U17725 (N_17725,N_15509,N_14193);
nand U17726 (N_17726,N_15556,N_14000);
nand U17727 (N_17727,N_14611,N_15215);
xnor U17728 (N_17728,N_15087,N_14903);
or U17729 (N_17729,N_14114,N_15383);
xnor U17730 (N_17730,N_15036,N_14673);
or U17731 (N_17731,N_15307,N_14043);
nor U17732 (N_17732,N_15759,N_14399);
and U17733 (N_17733,N_15231,N_15458);
and U17734 (N_17734,N_14005,N_15588);
or U17735 (N_17735,N_15643,N_15407);
and U17736 (N_17736,N_15744,N_15937);
and U17737 (N_17737,N_14650,N_14791);
and U17738 (N_17738,N_14687,N_14141);
nor U17739 (N_17739,N_15113,N_15081);
nand U17740 (N_17740,N_15200,N_15383);
xnor U17741 (N_17741,N_14001,N_14428);
nor U17742 (N_17742,N_14431,N_15092);
nand U17743 (N_17743,N_14299,N_14758);
or U17744 (N_17744,N_15379,N_14848);
nor U17745 (N_17745,N_15810,N_15647);
and U17746 (N_17746,N_14314,N_15448);
xor U17747 (N_17747,N_15740,N_15496);
or U17748 (N_17748,N_15154,N_15867);
or U17749 (N_17749,N_14716,N_14071);
xor U17750 (N_17750,N_15943,N_14695);
nor U17751 (N_17751,N_15898,N_15424);
and U17752 (N_17752,N_14746,N_15264);
nor U17753 (N_17753,N_14912,N_15679);
nor U17754 (N_17754,N_15835,N_15461);
and U17755 (N_17755,N_15765,N_15496);
xor U17756 (N_17756,N_15202,N_14338);
nor U17757 (N_17757,N_15009,N_14275);
or U17758 (N_17758,N_15135,N_15738);
and U17759 (N_17759,N_14312,N_15524);
or U17760 (N_17760,N_15254,N_14323);
or U17761 (N_17761,N_15850,N_15641);
or U17762 (N_17762,N_15969,N_14322);
nand U17763 (N_17763,N_15642,N_15847);
or U17764 (N_17764,N_15689,N_14062);
and U17765 (N_17765,N_14406,N_14744);
nor U17766 (N_17766,N_15166,N_15169);
nor U17767 (N_17767,N_15616,N_15220);
or U17768 (N_17768,N_15499,N_14959);
or U17769 (N_17769,N_14972,N_14585);
or U17770 (N_17770,N_14611,N_14339);
nand U17771 (N_17771,N_14155,N_14909);
nor U17772 (N_17772,N_14944,N_15366);
nand U17773 (N_17773,N_14658,N_14104);
xor U17774 (N_17774,N_15932,N_14272);
and U17775 (N_17775,N_14457,N_15466);
nor U17776 (N_17776,N_15483,N_14191);
nor U17777 (N_17777,N_15094,N_15847);
nand U17778 (N_17778,N_15695,N_15115);
xnor U17779 (N_17779,N_15467,N_14928);
nor U17780 (N_17780,N_15858,N_14617);
and U17781 (N_17781,N_14135,N_14208);
nor U17782 (N_17782,N_14777,N_14108);
nand U17783 (N_17783,N_15562,N_15242);
nand U17784 (N_17784,N_15721,N_15768);
nor U17785 (N_17785,N_15809,N_15895);
xnor U17786 (N_17786,N_14449,N_15627);
and U17787 (N_17787,N_14159,N_14955);
nand U17788 (N_17788,N_14548,N_14497);
xor U17789 (N_17789,N_14586,N_15336);
nor U17790 (N_17790,N_15149,N_14533);
xor U17791 (N_17791,N_14930,N_14293);
and U17792 (N_17792,N_14799,N_15100);
nor U17793 (N_17793,N_14946,N_15060);
nand U17794 (N_17794,N_14712,N_15243);
xor U17795 (N_17795,N_15281,N_14451);
nand U17796 (N_17796,N_15309,N_14838);
nor U17797 (N_17797,N_14620,N_15591);
xnor U17798 (N_17798,N_14334,N_15095);
and U17799 (N_17799,N_14750,N_15579);
nor U17800 (N_17800,N_14734,N_14726);
nand U17801 (N_17801,N_14283,N_14620);
xor U17802 (N_17802,N_15523,N_14828);
nand U17803 (N_17803,N_15877,N_14375);
or U17804 (N_17804,N_15347,N_14995);
and U17805 (N_17805,N_15380,N_14595);
nand U17806 (N_17806,N_14167,N_15030);
or U17807 (N_17807,N_14820,N_15067);
nand U17808 (N_17808,N_14574,N_15910);
or U17809 (N_17809,N_14776,N_15090);
nand U17810 (N_17810,N_14125,N_14524);
and U17811 (N_17811,N_15474,N_14257);
xnor U17812 (N_17812,N_14630,N_15721);
and U17813 (N_17813,N_14990,N_15798);
nor U17814 (N_17814,N_15580,N_15807);
nor U17815 (N_17815,N_15689,N_14831);
and U17816 (N_17816,N_14594,N_14318);
and U17817 (N_17817,N_15647,N_14993);
nand U17818 (N_17818,N_15477,N_14793);
xor U17819 (N_17819,N_15555,N_14643);
nor U17820 (N_17820,N_14127,N_14496);
nor U17821 (N_17821,N_15056,N_14560);
or U17822 (N_17822,N_14858,N_14438);
nand U17823 (N_17823,N_14628,N_15077);
nand U17824 (N_17824,N_14176,N_15016);
and U17825 (N_17825,N_14703,N_14821);
and U17826 (N_17826,N_15082,N_14378);
nand U17827 (N_17827,N_14365,N_14221);
or U17828 (N_17828,N_15027,N_14667);
xnor U17829 (N_17829,N_15524,N_14219);
xor U17830 (N_17830,N_15624,N_15373);
nor U17831 (N_17831,N_15555,N_15757);
nand U17832 (N_17832,N_14344,N_15532);
xnor U17833 (N_17833,N_15012,N_15844);
xnor U17834 (N_17834,N_15495,N_14549);
and U17835 (N_17835,N_15768,N_15758);
or U17836 (N_17836,N_15679,N_14659);
and U17837 (N_17837,N_14443,N_15137);
or U17838 (N_17838,N_14186,N_14291);
nand U17839 (N_17839,N_15254,N_14023);
or U17840 (N_17840,N_15544,N_15040);
or U17841 (N_17841,N_15498,N_15126);
and U17842 (N_17842,N_14859,N_14937);
and U17843 (N_17843,N_15018,N_15637);
and U17844 (N_17844,N_15841,N_14809);
nor U17845 (N_17845,N_15342,N_14748);
xor U17846 (N_17846,N_15842,N_15094);
or U17847 (N_17847,N_14365,N_14967);
nand U17848 (N_17848,N_15425,N_14960);
and U17849 (N_17849,N_14935,N_14030);
nand U17850 (N_17850,N_15400,N_14378);
or U17851 (N_17851,N_14726,N_14305);
xnor U17852 (N_17852,N_14184,N_14519);
nand U17853 (N_17853,N_14065,N_14541);
nor U17854 (N_17854,N_14592,N_14134);
nand U17855 (N_17855,N_14656,N_14243);
and U17856 (N_17856,N_14557,N_14055);
or U17857 (N_17857,N_14237,N_15760);
nand U17858 (N_17858,N_14314,N_14425);
and U17859 (N_17859,N_14299,N_15687);
xnor U17860 (N_17860,N_14780,N_14413);
and U17861 (N_17861,N_14798,N_14512);
nor U17862 (N_17862,N_14774,N_14938);
xnor U17863 (N_17863,N_14273,N_15220);
nor U17864 (N_17864,N_15551,N_15039);
or U17865 (N_17865,N_14073,N_15811);
nand U17866 (N_17866,N_14641,N_14381);
or U17867 (N_17867,N_15131,N_15938);
xnor U17868 (N_17868,N_14962,N_14781);
and U17869 (N_17869,N_14492,N_15761);
or U17870 (N_17870,N_15893,N_15788);
nand U17871 (N_17871,N_15882,N_15472);
xor U17872 (N_17872,N_15019,N_14789);
and U17873 (N_17873,N_15802,N_14325);
or U17874 (N_17874,N_14392,N_14411);
and U17875 (N_17875,N_15534,N_14972);
and U17876 (N_17876,N_15681,N_14425);
xor U17877 (N_17877,N_15275,N_15394);
nand U17878 (N_17878,N_14454,N_14573);
nand U17879 (N_17879,N_14340,N_15024);
nor U17880 (N_17880,N_14699,N_15641);
nand U17881 (N_17881,N_14961,N_14798);
and U17882 (N_17882,N_14407,N_15179);
nor U17883 (N_17883,N_14044,N_15589);
nor U17884 (N_17884,N_14375,N_15069);
or U17885 (N_17885,N_15153,N_14958);
nand U17886 (N_17886,N_15073,N_14685);
nor U17887 (N_17887,N_14182,N_15115);
or U17888 (N_17888,N_15991,N_14179);
xor U17889 (N_17889,N_15879,N_15607);
nor U17890 (N_17890,N_14416,N_14905);
and U17891 (N_17891,N_14524,N_15015);
nor U17892 (N_17892,N_14810,N_15596);
xor U17893 (N_17893,N_14719,N_14814);
xnor U17894 (N_17894,N_14279,N_15362);
nand U17895 (N_17895,N_14573,N_14155);
nand U17896 (N_17896,N_15428,N_15083);
nand U17897 (N_17897,N_15700,N_14917);
or U17898 (N_17898,N_15930,N_14691);
and U17899 (N_17899,N_15028,N_14787);
and U17900 (N_17900,N_14157,N_15566);
and U17901 (N_17901,N_14613,N_14705);
nor U17902 (N_17902,N_14999,N_14914);
or U17903 (N_17903,N_14862,N_15714);
nand U17904 (N_17904,N_15507,N_15615);
or U17905 (N_17905,N_15949,N_14231);
xor U17906 (N_17906,N_15795,N_14223);
nand U17907 (N_17907,N_15057,N_15631);
nor U17908 (N_17908,N_15259,N_15848);
nor U17909 (N_17909,N_15789,N_14201);
and U17910 (N_17910,N_14529,N_14035);
nor U17911 (N_17911,N_15214,N_15413);
nand U17912 (N_17912,N_15838,N_15828);
or U17913 (N_17913,N_15422,N_14778);
nor U17914 (N_17914,N_14520,N_14870);
nand U17915 (N_17915,N_14062,N_14654);
nor U17916 (N_17916,N_15790,N_14062);
nor U17917 (N_17917,N_15637,N_14499);
or U17918 (N_17918,N_15728,N_15980);
and U17919 (N_17919,N_14506,N_15894);
or U17920 (N_17920,N_14989,N_15214);
and U17921 (N_17921,N_15668,N_14681);
nand U17922 (N_17922,N_15167,N_14262);
nor U17923 (N_17923,N_14637,N_15404);
nor U17924 (N_17924,N_15019,N_14877);
nor U17925 (N_17925,N_15222,N_15423);
or U17926 (N_17926,N_14753,N_14859);
or U17927 (N_17927,N_15382,N_14560);
nor U17928 (N_17928,N_15520,N_14418);
and U17929 (N_17929,N_14427,N_15645);
and U17930 (N_17930,N_14461,N_14699);
or U17931 (N_17931,N_14551,N_15811);
and U17932 (N_17932,N_15952,N_15102);
nor U17933 (N_17933,N_15458,N_14249);
or U17934 (N_17934,N_14796,N_14061);
xor U17935 (N_17935,N_15563,N_14060);
nand U17936 (N_17936,N_14752,N_14732);
xnor U17937 (N_17937,N_15172,N_14921);
and U17938 (N_17938,N_14649,N_15191);
nor U17939 (N_17939,N_14421,N_14710);
or U17940 (N_17940,N_15299,N_15768);
or U17941 (N_17941,N_14139,N_14448);
nor U17942 (N_17942,N_14745,N_15721);
nor U17943 (N_17943,N_15520,N_14186);
or U17944 (N_17944,N_14489,N_14980);
nand U17945 (N_17945,N_14099,N_15527);
or U17946 (N_17946,N_15650,N_15850);
xnor U17947 (N_17947,N_14339,N_14891);
nor U17948 (N_17948,N_15336,N_14610);
xor U17949 (N_17949,N_14130,N_15010);
nand U17950 (N_17950,N_14079,N_14038);
xnor U17951 (N_17951,N_14515,N_15294);
nand U17952 (N_17952,N_14598,N_15970);
nand U17953 (N_17953,N_14211,N_15762);
nor U17954 (N_17954,N_15150,N_14394);
xor U17955 (N_17955,N_15422,N_14323);
and U17956 (N_17956,N_14263,N_15158);
nor U17957 (N_17957,N_15409,N_14938);
or U17958 (N_17958,N_15539,N_14512);
or U17959 (N_17959,N_15698,N_15669);
xor U17960 (N_17960,N_15427,N_15651);
or U17961 (N_17961,N_15841,N_15471);
and U17962 (N_17962,N_15414,N_14362);
or U17963 (N_17963,N_14901,N_14352);
nor U17964 (N_17964,N_15802,N_14015);
or U17965 (N_17965,N_14732,N_15400);
or U17966 (N_17966,N_14212,N_15821);
xor U17967 (N_17967,N_15612,N_15040);
and U17968 (N_17968,N_15779,N_15897);
or U17969 (N_17969,N_15830,N_15233);
xor U17970 (N_17970,N_14866,N_15548);
nor U17971 (N_17971,N_14696,N_15288);
or U17972 (N_17972,N_15488,N_14792);
nand U17973 (N_17973,N_14618,N_14939);
nor U17974 (N_17974,N_15057,N_15126);
and U17975 (N_17975,N_15909,N_15412);
or U17976 (N_17976,N_15977,N_15043);
xor U17977 (N_17977,N_14669,N_15725);
and U17978 (N_17978,N_14204,N_15812);
xor U17979 (N_17979,N_14716,N_14725);
xor U17980 (N_17980,N_14071,N_14476);
xor U17981 (N_17981,N_15504,N_15522);
or U17982 (N_17982,N_15473,N_15263);
xnor U17983 (N_17983,N_14632,N_14024);
nor U17984 (N_17984,N_15255,N_15817);
nand U17985 (N_17985,N_14905,N_15618);
and U17986 (N_17986,N_14829,N_15415);
and U17987 (N_17987,N_15291,N_14674);
nor U17988 (N_17988,N_15500,N_15842);
nand U17989 (N_17989,N_14123,N_15886);
nand U17990 (N_17990,N_15413,N_14858);
xnor U17991 (N_17991,N_14327,N_15653);
nor U17992 (N_17992,N_14663,N_15056);
nand U17993 (N_17993,N_14017,N_15839);
xor U17994 (N_17994,N_15241,N_14557);
xnor U17995 (N_17995,N_15458,N_14470);
and U17996 (N_17996,N_15670,N_14503);
nand U17997 (N_17997,N_14441,N_15466);
xnor U17998 (N_17998,N_14609,N_14671);
or U17999 (N_17999,N_15683,N_15878);
nand U18000 (N_18000,N_17019,N_16187);
and U18001 (N_18001,N_17076,N_16648);
nor U18002 (N_18002,N_17669,N_16273);
and U18003 (N_18003,N_17363,N_17618);
or U18004 (N_18004,N_17124,N_17601);
nand U18005 (N_18005,N_16325,N_16163);
nand U18006 (N_18006,N_16730,N_17354);
and U18007 (N_18007,N_17734,N_16917);
or U18008 (N_18008,N_17792,N_17255);
nor U18009 (N_18009,N_16921,N_16549);
and U18010 (N_18010,N_16841,N_16109);
xnor U18011 (N_18011,N_16903,N_17395);
nand U18012 (N_18012,N_16586,N_17544);
nand U18013 (N_18013,N_16885,N_16265);
nor U18014 (N_18014,N_16520,N_17310);
xnor U18015 (N_18015,N_17326,N_17700);
or U18016 (N_18016,N_16983,N_17082);
or U18017 (N_18017,N_17041,N_16387);
or U18018 (N_18018,N_17654,N_16287);
nand U18019 (N_18019,N_17085,N_16898);
and U18020 (N_18020,N_17987,N_17693);
nor U18021 (N_18021,N_16042,N_16130);
or U18022 (N_18022,N_17442,N_17362);
nand U18023 (N_18023,N_16366,N_16859);
nand U18024 (N_18024,N_17629,N_16064);
nand U18025 (N_18025,N_16143,N_16598);
and U18026 (N_18026,N_16432,N_16077);
xnor U18027 (N_18027,N_17995,N_17893);
and U18028 (N_18028,N_16112,N_16745);
or U18029 (N_18029,N_16926,N_16892);
xor U18030 (N_18030,N_16846,N_16528);
nor U18031 (N_18031,N_16182,N_16637);
nor U18032 (N_18032,N_16605,N_17619);
nand U18033 (N_18033,N_16963,N_17391);
nor U18034 (N_18034,N_16170,N_16172);
nor U18035 (N_18035,N_17592,N_17635);
or U18036 (N_18036,N_16680,N_17532);
nor U18037 (N_18037,N_17199,N_16041);
xor U18038 (N_18038,N_17923,N_16925);
and U18039 (N_18039,N_16496,N_17279);
or U18040 (N_18040,N_17115,N_16357);
nor U18041 (N_18041,N_16213,N_17841);
and U18042 (N_18042,N_16247,N_17180);
and U18043 (N_18043,N_17133,N_17768);
and U18044 (N_18044,N_17691,N_16495);
xnor U18045 (N_18045,N_16094,N_17811);
xnor U18046 (N_18046,N_17595,N_16578);
xnor U18047 (N_18047,N_17024,N_16322);
nor U18048 (N_18048,N_16568,N_16938);
xnor U18049 (N_18049,N_17212,N_16615);
nor U18050 (N_18050,N_17930,N_16952);
and U18051 (N_18051,N_16764,N_17485);
nand U18052 (N_18052,N_17039,N_16774);
and U18053 (N_18053,N_17806,N_17773);
or U18054 (N_18054,N_16304,N_17189);
xnor U18055 (N_18055,N_16297,N_17671);
nand U18056 (N_18056,N_16812,N_16973);
nand U18057 (N_18057,N_16439,N_16884);
xnor U18058 (N_18058,N_17661,N_16639);
nand U18059 (N_18059,N_16338,N_17822);
or U18060 (N_18060,N_16302,N_16013);
nor U18061 (N_18061,N_17946,N_17584);
and U18062 (N_18062,N_17044,N_16239);
nand U18063 (N_18063,N_17507,N_16089);
nand U18064 (N_18064,N_16236,N_16434);
nor U18065 (N_18065,N_17439,N_17608);
and U18066 (N_18066,N_17373,N_16998);
or U18067 (N_18067,N_17285,N_17665);
or U18068 (N_18068,N_17218,N_17426);
xnor U18069 (N_18069,N_17639,N_16607);
or U18070 (N_18070,N_16240,N_16244);
nor U18071 (N_18071,N_17980,N_17334);
xor U18072 (N_18072,N_17481,N_17720);
or U18073 (N_18073,N_16090,N_17386);
nand U18074 (N_18074,N_16275,N_17451);
and U18075 (N_18075,N_17855,N_16369);
nand U18076 (N_18076,N_16719,N_16497);
and U18077 (N_18077,N_16652,N_16819);
nand U18078 (N_18078,N_16294,N_16144);
and U18079 (N_18079,N_17029,N_17933);
or U18080 (N_18080,N_17003,N_16817);
nand U18081 (N_18081,N_17197,N_17256);
and U18082 (N_18082,N_16487,N_17091);
and U18083 (N_18083,N_17702,N_17936);
and U18084 (N_18084,N_17139,N_16243);
nand U18085 (N_18085,N_17847,N_16115);
and U18086 (N_18086,N_16062,N_17515);
nand U18087 (N_18087,N_17820,N_16823);
xnor U18088 (N_18088,N_17273,N_16779);
or U18089 (N_18089,N_16481,N_17746);
or U18090 (N_18090,N_16479,N_17899);
xnor U18091 (N_18091,N_16268,N_16810);
xor U18092 (N_18092,N_16826,N_16448);
xnor U18093 (N_18093,N_16096,N_16845);
nor U18094 (N_18094,N_17129,N_17593);
and U18095 (N_18095,N_16574,N_17027);
and U18096 (N_18096,N_17898,N_17718);
or U18097 (N_18097,N_17598,N_17166);
or U18098 (N_18098,N_16336,N_16346);
and U18099 (N_18099,N_16451,N_17467);
and U18100 (N_18100,N_17525,N_16321);
or U18101 (N_18101,N_17871,N_16691);
nand U18102 (N_18102,N_17501,N_16811);
and U18103 (N_18103,N_17253,N_16397);
xor U18104 (N_18104,N_17788,N_17782);
nand U18105 (N_18105,N_16491,N_17016);
xnor U18106 (N_18106,N_17339,N_16738);
nand U18107 (N_18107,N_17494,N_17178);
nand U18108 (N_18108,N_16954,N_16512);
and U18109 (N_18109,N_17624,N_16022);
nor U18110 (N_18110,N_17135,N_16999);
xnor U18111 (N_18111,N_17920,N_17512);
and U18112 (N_18112,N_17008,N_17397);
xnor U18113 (N_18113,N_17257,N_16185);
xnor U18114 (N_18114,N_16050,N_16421);
or U18115 (N_18115,N_17906,N_16643);
nand U18116 (N_18116,N_17596,N_17996);
xnor U18117 (N_18117,N_17972,N_17134);
or U18118 (N_18118,N_16499,N_16660);
or U18119 (N_18119,N_17123,N_16360);
xor U18120 (N_18120,N_16933,N_16361);
nand U18121 (N_18121,N_17533,N_17190);
and U18122 (N_18122,N_16616,N_16771);
nand U18123 (N_18123,N_16476,N_17796);
and U18124 (N_18124,N_16267,N_17799);
nand U18125 (N_18125,N_17383,N_17406);
nor U18126 (N_18126,N_16551,N_16891);
nor U18127 (N_18127,N_17644,N_16069);
or U18128 (N_18128,N_16186,N_16003);
or U18129 (N_18129,N_17408,N_17430);
nor U18130 (N_18130,N_16405,N_16266);
nand U18131 (N_18131,N_16638,N_16900);
xor U18132 (N_18132,N_17350,N_17832);
nor U18133 (N_18133,N_16039,N_16987);
nor U18134 (N_18134,N_17433,N_16509);
or U18135 (N_18135,N_16494,N_17240);
or U18136 (N_18136,N_17424,N_17114);
nor U18137 (N_18137,N_17534,N_16228);
xor U18138 (N_18138,N_16735,N_16203);
nor U18139 (N_18139,N_16554,N_16004);
xnor U18140 (N_18140,N_17965,N_17264);
or U18141 (N_18141,N_16274,N_17309);
or U18142 (N_18142,N_16184,N_17713);
or U18143 (N_18143,N_16619,N_16118);
or U18144 (N_18144,N_16312,N_16351);
xor U18145 (N_18145,N_16393,N_16128);
and U18146 (N_18146,N_17777,N_16697);
nor U18147 (N_18147,N_17246,N_16376);
and U18148 (N_18148,N_16441,N_16027);
nand U18149 (N_18149,N_17925,N_16125);
nor U18150 (N_18150,N_16521,N_17859);
xor U18151 (N_18151,N_16688,N_17553);
nand U18152 (N_18152,N_16046,N_17294);
and U18153 (N_18153,N_17931,N_17698);
or U18154 (N_18154,N_16656,N_17018);
xor U18155 (N_18155,N_16733,N_17999);
or U18156 (N_18156,N_16552,N_16453);
nand U18157 (N_18157,N_16693,N_16559);
xor U18158 (N_18158,N_16806,N_17719);
xnor U18159 (N_18159,N_16091,N_17234);
and U18160 (N_18160,N_17293,N_16723);
xor U18161 (N_18161,N_17631,N_16659);
nor U18162 (N_18162,N_17472,N_17656);
and U18163 (N_18163,N_17225,N_16458);
and U18164 (N_18164,N_17186,N_17683);
and U18165 (N_18165,N_17181,N_16550);
and U18166 (N_18166,N_17120,N_16911);
nand U18167 (N_18167,N_17443,N_16024);
xnor U18168 (N_18168,N_17325,N_17261);
and U18169 (N_18169,N_16871,N_17548);
or U18170 (N_18170,N_16284,N_16726);
xor U18171 (N_18171,N_17037,N_16743);
nand U18172 (N_18172,N_17603,N_17591);
or U18173 (N_18173,N_16957,N_17108);
and U18174 (N_18174,N_17319,N_16533);
nor U18175 (N_18175,N_17667,N_16583);
or U18176 (N_18176,N_16160,N_16695);
nor U18177 (N_18177,N_17463,N_17049);
nor U18178 (N_18178,N_17382,N_17723);
xor U18179 (N_18179,N_16435,N_16791);
or U18180 (N_18180,N_17609,N_17174);
nand U18181 (N_18181,N_17538,N_17546);
nor U18182 (N_18182,N_16915,N_16640);
or U18183 (N_18183,N_16058,N_16593);
nor U18184 (N_18184,N_17983,N_16761);
nand U18185 (N_18185,N_17098,N_17853);
and U18186 (N_18186,N_17554,N_17416);
or U18187 (N_18187,N_17708,N_17306);
nand U18188 (N_18188,N_17149,N_17356);
nor U18189 (N_18189,N_17945,N_17826);
xnor U18190 (N_18190,N_17454,N_17405);
and U18191 (N_18191,N_17201,N_17524);
and U18192 (N_18192,N_17537,N_16463);
nor U18193 (N_18193,N_17348,N_17461);
and U18194 (N_18194,N_17072,N_17328);
nor U18195 (N_18195,N_16483,N_17958);
nor U18196 (N_18196,N_17500,N_16100);
xor U18197 (N_18197,N_17140,N_16378);
and U18198 (N_18198,N_16960,N_16288);
nand U18199 (N_18199,N_16994,N_16756);
and U18200 (N_18200,N_16959,N_17685);
nor U18201 (N_18201,N_17797,N_16707);
nor U18202 (N_18202,N_17238,N_17881);
nor U18203 (N_18203,N_16445,N_17298);
or U18204 (N_18204,N_17540,N_17484);
or U18205 (N_18205,N_17521,N_16264);
or U18206 (N_18206,N_17096,N_16352);
xnor U18207 (N_18207,N_17517,N_16675);
xnor U18208 (N_18208,N_17346,N_16888);
nand U18209 (N_18209,N_16147,N_16278);
nor U18210 (N_18210,N_17167,N_17195);
or U18211 (N_18211,N_16606,N_16237);
xnor U18212 (N_18212,N_17531,N_16602);
or U18213 (N_18213,N_17324,N_17938);
xnor U18214 (N_18214,N_17340,N_17728);
nand U18215 (N_18215,N_16698,N_17229);
and U18216 (N_18216,N_16793,N_16402);
or U18217 (N_18217,N_17307,N_16489);
and U18218 (N_18218,N_17497,N_17668);
or U18219 (N_18219,N_16950,N_16847);
xnor U18220 (N_18220,N_17368,N_17790);
xnor U18221 (N_18221,N_17824,N_16073);
and U18222 (N_18222,N_17342,N_16717);
or U18223 (N_18223,N_16327,N_17252);
nor U18224 (N_18224,N_16008,N_16132);
nand U18225 (N_18225,N_17655,N_17445);
nand U18226 (N_18226,N_17737,N_17961);
nand U18227 (N_18227,N_16498,N_16976);
or U18228 (N_18228,N_17349,N_17845);
xnor U18229 (N_18229,N_17403,N_17457);
nand U18230 (N_18230,N_17605,N_17374);
and U18231 (N_18231,N_17427,N_16010);
or U18232 (N_18232,N_17528,N_17684);
or U18233 (N_18233,N_16544,N_17640);
nor U18234 (N_18234,N_16685,N_17156);
nand U18235 (N_18235,N_17176,N_16941);
nor U18236 (N_18236,N_17244,N_17316);
nand U18237 (N_18237,N_16825,N_16256);
nor U18238 (N_18238,N_17370,N_17105);
or U18239 (N_18239,N_16067,N_17510);
nand U18240 (N_18240,N_17557,N_17075);
nor U18241 (N_18241,N_17814,N_16828);
and U18242 (N_18242,N_17750,N_17150);
nand U18243 (N_18243,N_17440,N_16838);
or U18244 (N_18244,N_16540,N_17864);
nor U18245 (N_18245,N_16250,N_16792);
and U18246 (N_18246,N_17318,N_16683);
xor U18247 (N_18247,N_16519,N_17805);
nor U18248 (N_18248,N_17558,N_16958);
nor U18249 (N_18249,N_16923,N_17121);
nand U18250 (N_18250,N_16134,N_17425);
xor U18251 (N_18251,N_16153,N_17565);
or U18252 (N_18252,N_16469,N_16359);
and U18253 (N_18253,N_16875,N_17081);
or U18254 (N_18254,N_17338,N_17935);
and U18255 (N_18255,N_17606,N_16381);
and U18256 (N_18256,N_16565,N_17755);
or U18257 (N_18257,N_16214,N_16603);
and U18258 (N_18258,N_17753,N_17270);
xnor U18259 (N_18259,N_17874,N_16257);
nand U18260 (N_18260,N_17550,N_16610);
nor U18261 (N_18261,N_16157,N_17882);
nor U18262 (N_18262,N_17955,N_17097);
and U18263 (N_18263,N_16080,N_16460);
nand U18264 (N_18264,N_17284,N_16882);
xnor U18265 (N_18265,N_17227,N_16066);
nor U18266 (N_18266,N_16329,N_16618);
nor U18267 (N_18267,N_17131,N_17361);
xor U18268 (N_18268,N_17269,N_17113);
nand U18269 (N_18269,N_16292,N_16662);
xor U18270 (N_18270,N_17359,N_16017);
nor U18271 (N_18271,N_16804,N_16065);
nor U18272 (N_18272,N_17988,N_16422);
nand U18273 (N_18273,N_16687,N_17968);
xnor U18274 (N_18274,N_16150,N_16371);
or U18275 (N_18275,N_16696,N_17569);
or U18276 (N_18276,N_16235,N_17479);
nand U18277 (N_18277,N_17341,N_17645);
or U18278 (N_18278,N_16148,N_17102);
nand U18279 (N_18279,N_16874,N_16864);
nor U18280 (N_18280,N_17202,N_17030);
or U18281 (N_18281,N_16720,N_16117);
and U18282 (N_18282,N_16566,N_17164);
or U18283 (N_18283,N_16047,N_16083);
or U18284 (N_18284,N_16108,N_16258);
nand U18285 (N_18285,N_17917,N_17077);
or U18286 (N_18286,N_16585,N_16000);
nor U18287 (N_18287,N_17421,N_17069);
nand U18288 (N_18288,N_17660,N_16450);
xor U18289 (N_18289,N_17610,N_16625);
and U18290 (N_18290,N_17211,N_16341);
xnor U18291 (N_18291,N_17207,N_17233);
xnor U18292 (N_18292,N_16632,N_16576);
and U18293 (N_18293,N_16036,N_16121);
nor U18294 (N_18294,N_17809,N_17803);
nor U18295 (N_18295,N_17161,N_17262);
or U18296 (N_18296,N_16149,N_16415);
or U18297 (N_18297,N_17873,N_17947);
and U18298 (N_18298,N_16834,N_17158);
nand U18299 (N_18299,N_16881,N_16613);
nor U18300 (N_18300,N_16682,N_17926);
and U18301 (N_18301,N_17948,N_16635);
nand U18302 (N_18302,N_16703,N_16671);
or U18303 (N_18303,N_16527,N_16485);
nand U18304 (N_18304,N_16873,N_16518);
or U18305 (N_18305,N_16617,N_17854);
nor U18306 (N_18306,N_16399,N_16208);
nor U18307 (N_18307,N_16964,N_17870);
xor U18308 (N_18308,N_16135,N_16946);
xnor U18309 (N_18309,N_16714,N_17078);
nand U18310 (N_18310,N_16689,N_16795);
or U18311 (N_18311,N_17783,N_16282);
and U18312 (N_18312,N_16323,N_17110);
or U18313 (N_18313,N_16155,N_17767);
and U18314 (N_18314,N_17617,N_16829);
or U18315 (N_18315,N_16139,N_16525);
nor U18316 (N_18316,N_17800,N_16866);
and U18317 (N_18317,N_16484,N_17748);
xnor U18318 (N_18318,N_17574,N_17944);
or U18319 (N_18319,N_17827,N_16763);
or U18320 (N_18320,N_17612,N_16464);
xor U18321 (N_18321,N_17675,N_16320);
nor U18322 (N_18322,N_17589,N_17613);
xor U18323 (N_18323,N_17887,N_16220);
xnor U18324 (N_18324,N_16443,N_16951);
xnor U18325 (N_18325,N_17924,N_17004);
xnor U18326 (N_18326,N_17290,N_16466);
nand U18327 (N_18327,N_17280,N_17320);
and U18328 (N_18328,N_16389,N_17474);
nor U18329 (N_18329,N_16556,N_17151);
xor U18330 (N_18330,N_17377,N_17986);
nand U18331 (N_18331,N_16663,N_16541);
or U18332 (N_18332,N_17883,N_17641);
nand U18333 (N_18333,N_17456,N_16383);
nor U18334 (N_18334,N_16651,N_17851);
nor U18335 (N_18335,N_17231,N_17122);
nand U18336 (N_18336,N_16230,N_16515);
and U18337 (N_18337,N_16098,N_16391);
or U18338 (N_18338,N_16621,N_17721);
nor U18339 (N_18339,N_17801,N_17664);
nor U18340 (N_18340,N_17804,N_16043);
and U18341 (N_18341,N_17251,N_16277);
and U18342 (N_18342,N_16055,N_16461);
nand U18343 (N_18343,N_17302,N_17894);
and U18344 (N_18344,N_16584,N_16295);
nor U18345 (N_18345,N_16783,N_16867);
nand U18346 (N_18346,N_17050,N_17380);
or U18347 (N_18347,N_17247,N_17304);
nand U18348 (N_18348,N_17242,N_16626);
nand U18349 (N_18349,N_16390,N_16815);
or U18350 (N_18350,N_16020,N_17818);
nand U18351 (N_18351,N_17017,N_16116);
nand U18352 (N_18352,N_17000,N_16305);
nor U18353 (N_18353,N_16537,N_17848);
nor U18354 (N_18354,N_17505,N_17957);
xor U18355 (N_18355,N_16209,N_17715);
nor U18356 (N_18356,N_17886,N_17100);
xnor U18357 (N_18357,N_16251,N_16192);
nor U18358 (N_18358,N_16194,N_16271);
or U18359 (N_18359,N_16049,N_16562);
xor U18360 (N_18360,N_17688,N_16252);
nand U18361 (N_18361,N_17205,N_16326);
and U18362 (N_18362,N_17058,N_16486);
xnor U18363 (N_18363,N_17080,N_17292);
xnor U18364 (N_18364,N_17198,N_16226);
nor U18365 (N_18365,N_16099,N_16981);
or U18366 (N_18366,N_17545,N_16511);
nand U18367 (N_18367,N_16832,N_16260);
nor U18368 (N_18368,N_17740,N_17840);
and U18369 (N_18369,N_16704,N_17448);
and U18370 (N_18370,N_17147,N_17384);
nor U18371 (N_18371,N_16146,N_16927);
nor U18372 (N_18372,N_16212,N_17117);
xnor U18373 (N_18373,N_16942,N_16347);
xnor U18374 (N_18374,N_16409,N_16989);
nor U18375 (N_18375,N_17288,N_16508);
nor U18376 (N_18376,N_16547,N_16961);
xnor U18377 (N_18377,N_17489,N_16009);
nand U18378 (N_18378,N_17055,N_17813);
nor U18379 (N_18379,N_16372,N_16849);
xnor U18380 (N_18380,N_16851,N_16897);
xnor U18381 (N_18381,N_16503,N_16152);
and U18382 (N_18382,N_16993,N_17191);
xnor U18383 (N_18383,N_16506,N_16427);
xor U18384 (N_18384,N_17892,N_16164);
and U18385 (N_18385,N_17332,N_16138);
xor U18386 (N_18386,N_16018,N_16907);
xnor U18387 (N_18387,N_16301,N_16536);
or U18388 (N_18388,N_17934,N_17301);
nand U18389 (N_18389,N_17763,N_17276);
and U18390 (N_18390,N_16308,N_16104);
xor U18391 (N_18391,N_16014,N_17070);
nand U18392 (N_18392,N_16051,N_16910);
xnor U18393 (N_18393,N_16831,N_17283);
nand U18394 (N_18394,N_16535,N_17973);
or U18395 (N_18395,N_16711,N_16200);
and U18396 (N_18396,N_16860,N_16669);
nor U18397 (N_18397,N_16137,N_17842);
nand U18398 (N_18398,N_17975,N_16385);
nor U18399 (N_18399,N_17045,N_16015);
nand U18400 (N_18400,N_16437,N_17436);
and U18401 (N_18401,N_16839,N_16948);
or U18402 (N_18402,N_17404,N_17530);
or U18403 (N_18403,N_17305,N_17071);
xnor U18404 (N_18404,N_16677,N_17789);
xor U18405 (N_18405,N_17682,N_17877);
nor U18406 (N_18406,N_17837,N_17679);
xor U18407 (N_18407,N_17185,N_16340);
and U18408 (N_18408,N_16931,N_16095);
or U18409 (N_18409,N_16289,N_16916);
and U18410 (N_18410,N_17499,N_17297);
nor U18411 (N_18411,N_17496,N_17317);
nand U18412 (N_18412,N_17575,N_17833);
xor U18413 (N_18413,N_17171,N_17602);
nor U18414 (N_18414,N_17209,N_17065);
nor U18415 (N_18415,N_16702,N_16914);
or U18416 (N_18416,N_17323,N_17327);
nor U18417 (N_18417,N_16581,N_17143);
and U18418 (N_18418,N_16580,N_16488);
and U18419 (N_18419,N_16664,N_17520);
nor U18420 (N_18420,N_16367,N_16814);
xor U18421 (N_18421,N_16335,N_17254);
or U18422 (N_18422,N_16668,N_16345);
xor U18423 (N_18423,N_16579,N_17083);
nor U18424 (N_18424,N_17393,N_16079);
xnor U18425 (N_18425,N_17435,N_17633);
and U18426 (N_18426,N_17969,N_16752);
xor U18427 (N_18427,N_17163,N_17838);
and U18428 (N_18428,N_17217,N_16131);
nand U18429 (N_18429,N_17086,N_17519);
and U18430 (N_18430,N_16673,N_16978);
or U18431 (N_18431,N_17476,N_16166);
xor U18432 (N_18432,N_17681,N_16715);
xnor U18433 (N_18433,N_16548,N_16564);
nor U18434 (N_18434,N_16595,N_17148);
xor U18435 (N_18435,N_16224,N_16798);
nor U18436 (N_18436,N_17104,N_17599);
xor U18437 (N_18437,N_17570,N_17492);
and U18438 (N_18438,N_17007,N_16207);
and U18439 (N_18439,N_16456,N_17040);
or U18440 (N_18440,N_16986,N_17588);
and U18441 (N_18441,N_16530,N_16328);
nor U18442 (N_18442,N_17729,N_17092);
nand U18443 (N_18443,N_16765,N_16883);
xor U18444 (N_18444,N_17761,N_16262);
nor U18445 (N_18445,N_17219,N_17277);
nor U18446 (N_18446,N_16922,N_17490);
and U18447 (N_18447,N_17402,N_17895);
and U18448 (N_18448,N_16869,N_17646);
nor U18449 (N_18449,N_17036,N_17032);
xor U18450 (N_18450,N_16173,N_16248);
and U18451 (N_18451,N_17666,N_17245);
xnor U18452 (N_18452,N_17722,N_17726);
nor U18453 (N_18453,N_17849,N_16136);
nand U18454 (N_18454,N_17127,N_16123);
nor U18455 (N_18455,N_16944,N_16056);
nand U18456 (N_18456,N_16588,N_16316);
nand U18457 (N_18457,N_16344,N_16231);
nand U18458 (N_18458,N_17749,N_16740);
xor U18459 (N_18459,N_17088,N_16234);
and U18460 (N_18460,N_17066,N_17056);
nand U18461 (N_18461,N_16781,N_16545);
or U18462 (N_18462,N_16007,N_16854);
nor U18463 (N_18463,N_16113,N_17954);
nand U18464 (N_18464,N_17703,N_16856);
and U18465 (N_18465,N_17031,N_16201);
xnor U18466 (N_18466,N_17539,N_17657);
nand U18467 (N_18467,N_16667,N_17237);
nand U18468 (N_18468,N_16560,N_16021);
or U18469 (N_18469,N_16416,N_16830);
or U18470 (N_18470,N_16889,N_17872);
or U18471 (N_18471,N_17351,N_17784);
nand U18472 (N_18472,N_17409,N_17099);
nor U18473 (N_18473,N_17552,N_17630);
nor U18474 (N_18474,N_17491,N_17213);
nand U18475 (N_18475,N_16026,N_17358);
and U18476 (N_18476,N_17977,N_16582);
nand U18477 (N_18477,N_17367,N_16759);
and U18478 (N_18478,N_17200,N_17677);
or U18479 (N_18479,N_16894,N_17459);
nand U18480 (N_18480,N_17953,N_16967);
or U18481 (N_18481,N_16174,N_16071);
and U18482 (N_18482,N_16293,N_16417);
and U18483 (N_18483,N_16513,N_16087);
and U18484 (N_18484,N_16997,N_17353);
or U18485 (N_18485,N_17910,N_16468);
xor U18486 (N_18486,N_16424,N_16879);
nand U18487 (N_18487,N_17263,N_17733);
nand U18488 (N_18488,N_17559,N_17503);
nand U18489 (N_18489,N_17689,N_16542);
nor U18490 (N_18490,N_17577,N_17678);
nand U18491 (N_18491,N_17336,N_16646);
nand U18492 (N_18492,N_17952,N_16971);
nand U18493 (N_18493,N_17407,N_17586);
or U18494 (N_18494,N_17692,N_17652);
nand U18495 (N_18495,N_16229,N_16124);
or U18496 (N_18496,N_17431,N_17909);
xor U18497 (N_18497,N_16122,N_16082);
xor U18498 (N_18498,N_17420,N_16311);
xnor U18499 (N_18499,N_17312,N_16475);
and U18500 (N_18500,N_16772,N_17429);
nor U18501 (N_18501,N_16741,N_17686);
xnor U18502 (N_18502,N_17146,N_17366);
nand U18503 (N_18503,N_16449,N_16317);
and U18504 (N_18504,N_17398,N_16852);
nor U18505 (N_18505,N_17468,N_16797);
nand U18506 (N_18506,N_17981,N_17829);
xnor U18507 (N_18507,N_16002,N_17059);
xor U18508 (N_18508,N_17412,N_17950);
xor U18509 (N_18509,N_17839,N_17052);
nand U18510 (N_18510,N_16612,N_16404);
xor U18511 (N_18511,N_16102,N_16016);
xor U18512 (N_18512,N_16362,N_17417);
or U18513 (N_18513,N_17504,N_17576);
and U18514 (N_18514,N_17597,N_16040);
nor U18515 (N_18515,N_16053,N_16622);
or U18516 (N_18516,N_17711,N_17649);
nand U18517 (N_18517,N_16219,N_16929);
and U18518 (N_18518,N_16478,N_16589);
nor U18519 (N_18519,N_16844,N_17258);
nand U18520 (N_18520,N_16665,N_16760);
xor U18521 (N_18521,N_17132,N_17203);
xnor U18522 (N_18522,N_17902,N_16045);
nand U18523 (N_18523,N_16023,N_17775);
and U18524 (N_18524,N_16824,N_17175);
and U18525 (N_18525,N_17696,N_16198);
xor U18526 (N_18526,N_16661,N_17875);
xor U18527 (N_18527,N_17418,N_16835);
or U18528 (N_18528,N_17912,N_17759);
and U18529 (N_18529,N_16650,N_16757);
nor U18530 (N_18530,N_16742,N_16330);
or U18531 (N_18531,N_17614,N_17817);
and U18532 (N_18532,N_16353,N_17107);
and U18533 (N_18533,N_17756,N_17278);
or U18534 (N_18534,N_17876,N_17626);
or U18535 (N_18535,N_17498,N_16753);
and U18536 (N_18536,N_16802,N_16517);
nand U18537 (N_18537,N_17793,N_16546);
nor U18538 (N_18538,N_16608,N_17329);
and U18539 (N_18539,N_17757,N_17053);
or U18540 (N_18540,N_16392,N_16725);
xnor U18541 (N_18541,N_17951,N_17441);
and U18542 (N_18542,N_16692,N_17464);
nand U18543 (N_18543,N_17862,N_17101);
nor U18544 (N_18544,N_16523,N_17674);
xor U18545 (N_18545,N_16199,N_17449);
and U18546 (N_18546,N_17850,N_17028);
or U18547 (N_18547,N_16750,N_17964);
xor U18548 (N_18548,N_16674,N_16827);
nor U18549 (N_18549,N_17615,N_17857);
and U18550 (N_18550,N_17808,N_16375);
or U18551 (N_18551,N_17480,N_16238);
xnor U18552 (N_18552,N_16762,N_17248);
nor U18553 (N_18553,N_17073,N_16400);
or U18554 (N_18554,N_17103,N_16842);
xor U18555 (N_18555,N_16744,N_16363);
nor U18556 (N_18556,N_17184,N_16853);
xnor U18557 (N_18557,N_16342,N_16377);
or U18558 (N_18558,N_16423,N_16044);
or U18559 (N_18559,N_16895,N_17160);
nand U18560 (N_18560,N_16038,N_16171);
nand U18561 (N_18561,N_17780,N_16355);
nand U18562 (N_18562,N_17868,N_17567);
or U18563 (N_18563,N_16522,N_16202);
and U18564 (N_18564,N_16930,N_17653);
or U18565 (N_18565,N_16868,N_17054);
nor U18566 (N_18566,N_17482,N_17971);
or U18567 (N_18567,N_17785,N_17982);
nor U18568 (N_18568,N_17963,N_17224);
xor U18569 (N_18569,N_17090,N_16837);
nor U18570 (N_18570,N_17549,N_16388);
and U18571 (N_18571,N_16012,N_16647);
xnor U18572 (N_18572,N_16276,N_16145);
or U18573 (N_18573,N_17168,N_17087);
and U18574 (N_18574,N_17111,N_17828);
nand U18575 (N_18575,N_17993,N_16614);
nor U18576 (N_18576,N_17043,N_17013);
xnor U18577 (N_18577,N_17516,N_17637);
xnor U18578 (N_18578,N_16782,N_17266);
and U18579 (N_18579,N_17513,N_17787);
nand U18580 (N_18580,N_16384,N_17033);
or U18581 (N_18581,N_17568,N_17432);
or U18582 (N_18582,N_16644,N_17536);
nor U18583 (N_18583,N_17916,N_17236);
and U18584 (N_18584,N_16596,N_16374);
nor U18585 (N_18585,N_16822,N_17672);
and U18586 (N_18586,N_17716,N_16031);
or U18587 (N_18587,N_17786,N_16205);
nor U18588 (N_18588,N_16887,N_16939);
nor U18589 (N_18589,N_17385,N_16555);
nand U18590 (N_18590,N_17437,N_16334);
xor U18591 (N_18591,N_17694,N_17770);
and U18592 (N_18592,N_17835,N_17736);
or U18593 (N_18593,N_17911,N_16721);
and U18594 (N_18594,N_16591,N_16800);
nor U18595 (N_18595,N_16074,N_17778);
or U18596 (N_18596,N_17680,N_17315);
xnor U18597 (N_18597,N_16072,N_16553);
and U18598 (N_18598,N_17493,N_16712);
xnor U18599 (N_18599,N_17172,N_17469);
nand U18600 (N_18600,N_16956,N_16701);
and U18601 (N_18601,N_16269,N_16645);
or U18602 (N_18602,N_16979,N_16382);
nand U18603 (N_18603,N_17130,N_17428);
xor U18604 (N_18604,N_16216,N_16075);
and U18605 (N_18605,N_17452,N_17331);
or U18606 (N_18606,N_17620,N_17600);
xnor U18607 (N_18607,N_17542,N_16705);
nand U18608 (N_18608,N_17878,N_16597);
and U18609 (N_18609,N_17976,N_16057);
xnor U18610 (N_18610,N_17856,N_16204);
nor U18611 (N_18611,N_16318,N_17450);
nand U18612 (N_18612,N_16430,N_17564);
nand U18613 (N_18613,N_17866,N_16431);
nand U18614 (N_18614,N_17760,N_17974);
and U18615 (N_18615,N_16206,N_16350);
xor U18616 (N_18616,N_17526,N_16624);
and U18617 (N_18617,N_17012,N_17118);
xnor U18618 (N_18618,N_16246,N_17155);
and U18619 (N_18619,N_16975,N_16679);
or U18620 (N_18620,N_16493,N_16690);
nand U18621 (N_18621,N_16919,N_16354);
nor U18622 (N_18622,N_17064,N_16129);
and U18623 (N_18623,N_17057,N_16601);
and U18624 (N_18624,N_17663,N_17400);
or U18625 (N_18625,N_16855,N_17891);
nor U18626 (N_18626,N_16935,N_17707);
or U18627 (N_18627,N_16748,N_17890);
and U18628 (N_18628,N_16500,N_16840);
or U18629 (N_18629,N_16955,N_16746);
nand U18630 (N_18630,N_16179,N_17628);
xor U18631 (N_18631,N_16168,N_17243);
or U18632 (N_18632,N_16928,N_16773);
or U18633 (N_18633,N_16455,N_17223);
and U18634 (N_18634,N_16514,N_17011);
and U18635 (N_18635,N_17487,N_17555);
and U18636 (N_18636,N_17365,N_17159);
or U18637 (N_18637,N_16642,N_16641);
and U18638 (N_18638,N_17343,N_17594);
or U18639 (N_18639,N_16974,N_16154);
nor U18640 (N_18640,N_16380,N_16370);
nand U18641 (N_18641,N_17810,N_17230);
xor U18642 (N_18642,N_17551,N_17867);
and U18643 (N_18643,N_16306,N_16790);
xor U18644 (N_18644,N_16953,N_17794);
or U18645 (N_18645,N_17392,N_16365);
nand U18646 (N_18646,N_17462,N_16188);
xnor U18647 (N_18647,N_16599,N_16890);
xnor U18648 (N_18648,N_16092,N_17414);
and U18649 (N_18649,N_17622,N_16425);
and U18650 (N_18650,N_16777,N_17998);
and U18651 (N_18651,N_17410,N_16270);
nand U18652 (N_18652,N_16708,N_16462);
xnor U18653 (N_18653,N_17563,N_17025);
nor U18654 (N_18654,N_16161,N_17754);
nor U18655 (N_18655,N_17411,N_17478);
xor U18656 (N_18656,N_17547,N_17769);
xor U18657 (N_18657,N_16303,N_16934);
or U18658 (N_18658,N_16655,N_17241);
or U18659 (N_18659,N_16232,N_16863);
and U18660 (N_18660,N_16905,N_16331);
nor U18661 (N_18661,N_17812,N_17676);
xnor U18662 (N_18662,N_16348,N_17821);
or U18663 (N_18663,N_17903,N_16937);
or U18664 (N_18664,N_16880,N_16259);
xor U18665 (N_18665,N_16029,N_17394);
xor U18666 (N_18666,N_17061,N_16729);
nor U18667 (N_18667,N_16438,N_16429);
nor U18668 (N_18668,N_17112,N_16472);
xnor U18669 (N_18669,N_16796,N_17699);
nand U18670 (N_18670,N_16426,N_17970);
or U18671 (N_18671,N_17738,N_16718);
nand U18672 (N_18672,N_16151,N_17128);
xor U18673 (N_18673,N_17337,N_17281);
xor U18674 (N_18674,N_16706,N_17741);
xnor U18675 (N_18675,N_16918,N_17194);
xnor U18676 (N_18676,N_16980,N_16534);
nor U18677 (N_18677,N_17731,N_17152);
xor U18678 (N_18678,N_16162,N_16368);
and U18679 (N_18679,N_17001,N_17035);
xor U18680 (N_18680,N_17745,N_17956);
or U18681 (N_18681,N_16636,N_16175);
nor U18682 (N_18682,N_17992,N_16623);
xor U18683 (N_18683,N_16356,N_16313);
xor U18684 (N_18684,N_16786,N_16176);
xnor U18685 (N_18685,N_16727,N_17662);
and U18686 (N_18686,N_17376,N_17330);
or U18687 (N_18687,N_16001,N_16751);
and U18688 (N_18688,N_17730,N_16156);
nor U18689 (N_18689,N_16492,N_16653);
xnor U18690 (N_18690,N_17154,N_17239);
or U18691 (N_18691,N_16700,N_16110);
xnor U18692 (N_18692,N_17632,N_17260);
xor U18693 (N_18693,N_16473,N_16211);
and U18694 (N_18694,N_17732,N_17807);
and U18695 (N_18695,N_17006,N_16731);
xor U18696 (N_18696,N_16893,N_16177);
nor U18697 (N_18697,N_17345,N_17735);
and U18698 (N_18698,N_16444,N_16280);
nor U18699 (N_18699,N_17423,N_16529);
nand U18700 (N_18700,N_17005,N_17145);
nand U18701 (N_18701,N_17831,N_17396);
nand U18702 (N_18702,N_16732,N_17888);
xnor U18703 (N_18703,N_17994,N_17182);
or U18704 (N_18704,N_17566,N_16222);
nor U18705 (N_18705,N_17752,N_16904);
nand U18706 (N_18706,N_17966,N_16114);
or U18707 (N_18707,N_16242,N_16710);
nor U18708 (N_18708,N_17523,N_17214);
nor U18709 (N_18709,N_16505,N_16221);
or U18710 (N_18710,N_17021,N_16364);
xor U18711 (N_18711,N_16969,N_17714);
nor U18712 (N_18712,N_16739,N_16410);
nand U18713 (N_18713,N_17289,N_16805);
nor U18714 (N_18714,N_17063,N_16452);
nand U18715 (N_18715,N_16982,N_17216);
or U18716 (N_18716,N_16337,N_17388);
nor U18717 (N_18717,N_16722,N_16803);
and U18718 (N_18718,N_17465,N_16538);
and U18719 (N_18719,N_16414,N_16672);
xnor U18720 (N_18720,N_16459,N_16571);
nor U18721 (N_18721,N_17772,N_17259);
and U18722 (N_18722,N_17271,N_16401);
nand U18723 (N_18723,N_17322,N_17488);
nor U18724 (N_18724,N_17060,N_16482);
nand U18725 (N_18725,N_16977,N_17267);
and U18726 (N_18726,N_16105,N_16754);
xor U18727 (N_18727,N_17583,N_16225);
nor U18728 (N_18728,N_17744,N_17942);
and U18729 (N_18729,N_16159,N_16126);
nand U18730 (N_18730,N_16788,N_16396);
xor U18731 (N_18731,N_16060,N_17705);
or U18732 (N_18732,N_16563,N_16480);
nand U18733 (N_18733,N_16101,N_16857);
nor U18734 (N_18734,N_17473,N_16085);
nand U18735 (N_18735,N_17670,N_16833);
nor U18736 (N_18736,N_16932,N_17094);
xor U18737 (N_18737,N_17372,N_17250);
nor U18738 (N_18738,N_17165,N_16218);
and U18739 (N_18739,N_16217,N_17169);
and U18740 (N_18740,N_17475,N_16630);
nand U18741 (N_18741,N_16436,N_17858);
nand U18742 (N_18742,N_16106,N_16962);
or U18743 (N_18743,N_17509,N_16787);
or U18744 (N_18744,N_17344,N_16985);
nand U18745 (N_18745,N_17908,N_16255);
or U18746 (N_18746,N_16052,N_16816);
nor U18747 (N_18747,N_17659,N_17299);
nand U18748 (N_18748,N_16924,N_17701);
or U18749 (N_18749,N_16501,N_17188);
nand U18750 (N_18750,N_17210,N_16314);
nor U18751 (N_18751,N_17861,N_17477);
xor U18752 (N_18752,N_17357,N_16557);
nand U18753 (N_18753,N_17453,N_17798);
and U18754 (N_18754,N_16249,N_16666);
nor U18755 (N_18755,N_16600,N_16283);
nor U18756 (N_18756,N_17268,N_17949);
or U18757 (N_18757,N_16319,N_17215);
nor U18758 (N_18758,N_17919,N_16920);
and U18759 (N_18759,N_16902,N_17514);
nand U18760 (N_18760,N_16210,N_17296);
or U18761 (N_18761,N_16567,N_17419);
nor U18762 (N_18762,N_17765,N_17997);
and U18763 (N_18763,N_16315,N_16629);
or U18764 (N_18764,N_16848,N_17743);
and U18765 (N_18765,N_16808,N_16133);
and U18766 (N_18766,N_17771,N_16996);
or U18767 (N_18767,N_16285,N_17896);
xor U18768 (N_18768,N_16223,N_16373);
nand U18769 (N_18769,N_16291,N_16227);
nor U18770 (N_18770,N_17047,N_17162);
nor U18771 (N_18771,N_17422,N_17978);
or U18772 (N_18772,N_17604,N_16609);
nand U18773 (N_18773,N_16970,N_17819);
nand U18774 (N_18774,N_17347,N_16477);
or U18775 (N_18775,N_17795,N_17321);
or U18776 (N_18776,N_16780,N_17438);
or U18777 (N_18777,N_16784,N_17647);
nor U18778 (N_18778,N_17204,N_16906);
and U18779 (N_18779,N_17460,N_17314);
xor U18780 (N_18780,N_17458,N_16794);
and U18781 (N_18781,N_17889,N_17308);
nor U18782 (N_18782,N_16778,N_17369);
or U18783 (N_18783,N_16093,N_17371);
and U18784 (N_18784,N_17561,N_16620);
xor U18785 (N_18785,N_16097,N_16411);
and U18786 (N_18786,N_16048,N_16678);
or U18787 (N_18787,N_17010,N_16858);
nand U18788 (N_18788,N_17381,N_16379);
nand U18789 (N_18789,N_17884,N_17506);
and U18790 (N_18790,N_16972,N_17747);
xnor U18791 (N_18791,N_17390,N_17979);
nor U18792 (N_18792,N_17046,N_17193);
or U18793 (N_18793,N_17885,N_17697);
and U18794 (N_18794,N_17495,N_16286);
xnor U18795 (N_18795,N_17560,N_17984);
and U18796 (N_18796,N_16862,N_17658);
nand U18797 (N_18797,N_17543,N_16870);
or U18798 (N_18798,N_17846,N_16940);
and U18799 (N_18799,N_16633,N_17922);
nand U18800 (N_18800,N_17119,N_17571);
xnor U18801 (N_18801,N_17830,N_16912);
nor U18802 (N_18802,N_17355,N_16412);
nand U18803 (N_18803,N_17643,N_16298);
nand U18804 (N_18804,N_16776,N_16775);
and U18805 (N_18805,N_17125,N_16634);
nand U18806 (N_18806,N_16191,N_17634);
nor U18807 (N_18807,N_16699,N_16809);
xor U18808 (N_18808,N_17836,N_17627);
xor U18809 (N_18809,N_16433,N_16573);
or U18810 (N_18810,N_16821,N_16061);
and U18811 (N_18811,N_17068,N_17106);
nand U18812 (N_18812,N_17623,N_16913);
xnor U18813 (N_18813,N_16716,N_16516);
nor U18814 (N_18814,N_16254,N_17153);
nor U18815 (N_18815,N_16836,N_16531);
nand U18816 (N_18816,N_17904,N_17611);
and U18817 (N_18817,N_17825,N_17823);
xnor U18818 (N_18818,N_17642,N_17335);
xnor U18819 (N_18819,N_16245,N_17562);
xnor U18820 (N_18820,N_16178,N_16358);
and U18821 (N_18821,N_16896,N_16196);
nor U18822 (N_18822,N_16769,N_17616);
nor U18823 (N_18823,N_17774,N_16649);
xor U18824 (N_18824,N_17880,N_17142);
nor U18825 (N_18825,N_17042,N_16332);
nand U18826 (N_18826,N_16684,N_16789);
nor U18827 (N_18827,N_16167,N_17579);
and U18828 (N_18828,N_17126,N_16799);
nor U18829 (N_18829,N_16467,N_16694);
nor U18830 (N_18830,N_16005,N_16310);
xnor U18831 (N_18831,N_17915,N_16878);
xor U18832 (N_18832,N_17585,N_17764);
nor U18833 (N_18833,N_16947,N_17196);
or U18834 (N_18834,N_16681,N_16006);
nor U18835 (N_18835,N_16386,N_16657);
or U18836 (N_18836,N_16886,N_16403);
xor U18837 (N_18837,N_16165,N_17816);
nor U18838 (N_18838,N_16734,N_17751);
xor U18839 (N_18839,N_17022,N_17535);
nand U18840 (N_18840,N_17897,N_17651);
nor U18841 (N_18841,N_17650,N_17274);
nand U18842 (N_18842,N_16086,N_17687);
nor U18843 (N_18843,N_16713,N_16577);
xor U18844 (N_18844,N_16558,N_16333);
nand U18845 (N_18845,N_17776,N_17116);
nor U18846 (N_18846,N_16296,N_16054);
or U18847 (N_18847,N_16454,N_17206);
nand U18848 (N_18848,N_16736,N_17907);
xor U18849 (N_18849,N_17352,N_17921);
and U18850 (N_18850,N_16119,N_17444);
nand U18851 (N_18851,N_16526,N_16801);
nand U18852 (N_18852,N_16654,N_16909);
nand U18853 (N_18853,N_17282,N_16766);
nand U18854 (N_18854,N_17742,N_17413);
nor U18855 (N_18855,N_16028,N_16570);
xor U18856 (N_18856,N_16032,N_17625);
xnor U18857 (N_18857,N_17179,N_16030);
xnor U18858 (N_18858,N_16324,N_16190);
or U18859 (N_18859,N_17062,N_16059);
nand U18860 (N_18860,N_16594,N_17590);
and U18861 (N_18861,N_16088,N_16861);
xor U18862 (N_18862,N_16628,N_17300);
and U18863 (N_18863,N_17802,N_16945);
nor U18864 (N_18864,N_16063,N_16447);
xnor U18865 (N_18865,N_16407,N_16899);
xor U18866 (N_18866,N_16876,N_16507);
and U18867 (N_18867,N_17673,N_17844);
nor U18868 (N_18868,N_17067,N_17572);
or U18869 (N_18869,N_17522,N_17962);
nand U18870 (N_18870,N_17378,N_16572);
nor U18871 (N_18871,N_17914,N_16767);
xnor U18872 (N_18872,N_17852,N_16183);
xnor U18873 (N_18873,N_16749,N_17581);
and U18874 (N_18874,N_16299,N_17286);
and U18875 (N_18875,N_17026,N_16502);
or U18876 (N_18876,N_17901,N_16446);
xor U18877 (N_18877,N_17399,N_16984);
nor U18878 (N_18878,N_16686,N_17303);
or U18879 (N_18879,N_16737,N_16428);
xor U18880 (N_18880,N_16877,N_16543);
or U18881 (N_18881,N_17990,N_16968);
xor U18882 (N_18882,N_16193,N_17084);
nand U18883 (N_18883,N_17991,N_16197);
nand U18884 (N_18884,N_16524,N_16709);
or U18885 (N_18885,N_16510,N_16081);
xnor U18886 (N_18886,N_17863,N_16747);
nand U18887 (N_18887,N_16413,N_17222);
and U18888 (N_18888,N_16343,N_17136);
nand U18889 (N_18889,N_17739,N_17228);
and U18890 (N_18890,N_16471,N_17932);
nor U18891 (N_18891,N_17638,N_16195);
nor U18892 (N_18892,N_17287,N_16539);
and U18893 (N_18893,N_16107,N_17941);
nand U18894 (N_18894,N_17959,N_16307);
xor U18895 (N_18895,N_17587,N_17529);
nor U18896 (N_18896,N_17717,N_16033);
or U18897 (N_18897,N_17582,N_17518);
nor U18898 (N_18898,N_17364,N_16785);
nor U18899 (N_18899,N_16770,N_17989);
or U18900 (N_18900,N_17313,N_17815);
and U18901 (N_18901,N_17295,N_16279);
and U18902 (N_18902,N_17527,N_17486);
nand U18903 (N_18903,N_16457,N_16068);
and U18904 (N_18904,N_17725,N_17221);
and U18905 (N_18905,N_17508,N_17177);
nand U18906 (N_18906,N_17208,N_16169);
nand U18907 (N_18907,N_17791,N_17900);
nor U18908 (N_18908,N_17170,N_16418);
nand U18909 (N_18909,N_16019,N_17928);
or U18910 (N_18910,N_17226,N_17913);
xor U18911 (N_18911,N_16281,N_17727);
nor U18912 (N_18912,N_16575,N_17183);
xnor U18913 (N_18913,N_16807,N_16724);
nand U18914 (N_18914,N_16419,N_16408);
nor U18915 (N_18915,N_16590,N_16901);
or U18916 (N_18916,N_17502,N_16949);
nand U18917 (N_18917,N_16532,N_17636);
nand U18918 (N_18918,N_17109,N_17333);
nor U18919 (N_18919,N_16180,N_17265);
nand U18920 (N_18920,N_16035,N_16943);
or U18921 (N_18921,N_17455,N_16398);
xor U18922 (N_18922,N_17573,N_17220);
nor U18923 (N_18923,N_16127,N_16676);
xor U18924 (N_18924,N_16490,N_17275);
and U18925 (N_18925,N_16070,N_17389);
xnor U18926 (N_18926,N_17762,N_16215);
nor U18927 (N_18927,N_16076,N_17192);
and U18928 (N_18928,N_16181,N_17758);
or U18929 (N_18929,N_17141,N_17051);
nor U18930 (N_18930,N_16442,N_17095);
xnor U18931 (N_18931,N_17860,N_16111);
nor U18932 (N_18932,N_16755,N_17985);
and U18933 (N_18933,N_16872,N_17724);
nand U18934 (N_18934,N_16158,N_17009);
xnor U18935 (N_18935,N_17939,N_17918);
nand U18936 (N_18936,N_16611,N_16865);
or U18937 (N_18937,N_16140,N_17093);
xnor U18938 (N_18938,N_17138,N_17695);
or U18939 (N_18939,N_17387,N_17048);
xor U18940 (N_18940,N_16290,N_17447);
or U18941 (N_18941,N_16758,N_16120);
or U18942 (N_18942,N_17879,N_16768);
nand U18943 (N_18943,N_17015,N_17905);
nor U18944 (N_18944,N_16406,N_16728);
nor U18945 (N_18945,N_16272,N_17272);
nor U18946 (N_18946,N_17466,N_17937);
or U18947 (N_18947,N_16995,N_17434);
nand U18948 (N_18948,N_17157,N_17869);
xor U18949 (N_18949,N_17766,N_16820);
or U18950 (N_18950,N_17311,N_17927);
xnor U18951 (N_18951,N_16241,N_17781);
or U18952 (N_18952,N_17023,N_16470);
and U18953 (N_18953,N_17556,N_17929);
or U18954 (N_18954,N_16142,N_16670);
nand U18955 (N_18955,N_17187,N_17541);
xnor U18956 (N_18956,N_17967,N_17843);
and U18957 (N_18957,N_17014,N_16440);
or U18958 (N_18958,N_17706,N_17648);
or U18959 (N_18959,N_17446,N_16037);
nor U18960 (N_18960,N_16465,N_16395);
xor U18961 (N_18961,N_16309,N_16084);
nand U18962 (N_18962,N_17415,N_16253);
nor U18963 (N_18963,N_17483,N_16966);
nand U18964 (N_18964,N_17943,N_16843);
or U18965 (N_18965,N_16349,N_16658);
nor U18966 (N_18966,N_17704,N_16850);
xnor U18967 (N_18967,N_17621,N_17249);
nand U18968 (N_18968,N_16233,N_16394);
and U18969 (N_18969,N_16078,N_16988);
nor U18970 (N_18970,N_16189,N_16561);
nand U18971 (N_18971,N_16936,N_17002);
nand U18972 (N_18972,N_16261,N_17960);
nor U18973 (N_18973,N_17865,N_17580);
and U18974 (N_18974,N_17471,N_16034);
xor U18975 (N_18975,N_16011,N_16592);
xor U18976 (N_18976,N_17038,N_17173);
and U18977 (N_18977,N_17020,N_16991);
nand U18978 (N_18978,N_17235,N_17034);
or U18979 (N_18979,N_16965,N_16103);
xnor U18980 (N_18980,N_16569,N_16025);
xor U18981 (N_18981,N_16604,N_16818);
nor U18982 (N_18982,N_17401,N_16908);
xor U18983 (N_18983,N_17511,N_16420);
nand U18984 (N_18984,N_17379,N_16300);
or U18985 (N_18985,N_17144,N_16504);
nand U18986 (N_18986,N_17232,N_17607);
or U18987 (N_18987,N_16992,N_17137);
xor U18988 (N_18988,N_17360,N_16990);
and U18989 (N_18989,N_17074,N_17690);
nand U18990 (N_18990,N_16587,N_16263);
nand U18991 (N_18991,N_17291,N_16339);
and U18992 (N_18992,N_17578,N_17712);
nor U18993 (N_18993,N_16474,N_16141);
and U18994 (N_18994,N_16627,N_17710);
nand U18995 (N_18995,N_17079,N_17089);
nand U18996 (N_18996,N_17470,N_17940);
or U18997 (N_18997,N_17834,N_16813);
nand U18998 (N_18998,N_17709,N_17779);
or U18999 (N_18999,N_17375,N_16631);
nor U19000 (N_19000,N_17465,N_16196);
or U19001 (N_19001,N_16778,N_17681);
and U19002 (N_19002,N_16689,N_16954);
xor U19003 (N_19003,N_16071,N_17426);
xor U19004 (N_19004,N_16156,N_17153);
nor U19005 (N_19005,N_16282,N_17021);
nand U19006 (N_19006,N_16054,N_17234);
or U19007 (N_19007,N_17340,N_16994);
nand U19008 (N_19008,N_17503,N_17404);
xnor U19009 (N_19009,N_17046,N_16861);
or U19010 (N_19010,N_17224,N_16656);
or U19011 (N_19011,N_17360,N_17561);
xnor U19012 (N_19012,N_16487,N_17736);
xor U19013 (N_19013,N_17864,N_16711);
or U19014 (N_19014,N_17380,N_17804);
and U19015 (N_19015,N_16933,N_17375);
and U19016 (N_19016,N_17159,N_17312);
or U19017 (N_19017,N_17901,N_17543);
nor U19018 (N_19018,N_17693,N_16172);
or U19019 (N_19019,N_16878,N_17814);
or U19020 (N_19020,N_17697,N_16261);
nor U19021 (N_19021,N_16370,N_17534);
and U19022 (N_19022,N_16495,N_16199);
xor U19023 (N_19023,N_16201,N_16025);
nor U19024 (N_19024,N_17533,N_16415);
nor U19025 (N_19025,N_16814,N_16448);
and U19026 (N_19026,N_17252,N_17567);
nor U19027 (N_19027,N_16290,N_17799);
nand U19028 (N_19028,N_17824,N_17609);
nor U19029 (N_19029,N_17095,N_16285);
xnor U19030 (N_19030,N_16021,N_17342);
nor U19031 (N_19031,N_16756,N_17441);
xnor U19032 (N_19032,N_16907,N_17796);
or U19033 (N_19033,N_17239,N_16648);
nand U19034 (N_19034,N_16539,N_16541);
and U19035 (N_19035,N_17532,N_17633);
xnor U19036 (N_19036,N_16906,N_17652);
nand U19037 (N_19037,N_16911,N_16718);
nor U19038 (N_19038,N_16231,N_17633);
xnor U19039 (N_19039,N_17551,N_16554);
xor U19040 (N_19040,N_17128,N_16292);
nor U19041 (N_19041,N_16520,N_16668);
or U19042 (N_19042,N_17670,N_17224);
and U19043 (N_19043,N_17707,N_17442);
or U19044 (N_19044,N_17974,N_16693);
nor U19045 (N_19045,N_16633,N_17952);
and U19046 (N_19046,N_16465,N_17843);
xor U19047 (N_19047,N_16183,N_17203);
or U19048 (N_19048,N_16492,N_17418);
nor U19049 (N_19049,N_17421,N_17658);
xor U19050 (N_19050,N_16021,N_17600);
nor U19051 (N_19051,N_16583,N_16856);
or U19052 (N_19052,N_16921,N_16343);
or U19053 (N_19053,N_16998,N_17010);
or U19054 (N_19054,N_16846,N_16372);
nor U19055 (N_19055,N_16579,N_16268);
xor U19056 (N_19056,N_16311,N_17442);
nor U19057 (N_19057,N_17270,N_16992);
nor U19058 (N_19058,N_17711,N_16511);
nand U19059 (N_19059,N_16466,N_16139);
nor U19060 (N_19060,N_17925,N_16103);
xnor U19061 (N_19061,N_17306,N_16842);
and U19062 (N_19062,N_16116,N_17527);
nand U19063 (N_19063,N_16549,N_17768);
nand U19064 (N_19064,N_17759,N_17469);
or U19065 (N_19065,N_16132,N_17103);
nor U19066 (N_19066,N_16424,N_17909);
or U19067 (N_19067,N_17154,N_17027);
nand U19068 (N_19068,N_16821,N_17126);
nand U19069 (N_19069,N_16808,N_17772);
xnor U19070 (N_19070,N_16705,N_17116);
nor U19071 (N_19071,N_16363,N_17041);
xor U19072 (N_19072,N_16717,N_17290);
nand U19073 (N_19073,N_16435,N_17323);
and U19074 (N_19074,N_16611,N_16006);
nand U19075 (N_19075,N_17084,N_16671);
or U19076 (N_19076,N_16683,N_17651);
nand U19077 (N_19077,N_16037,N_16609);
xnor U19078 (N_19078,N_17417,N_16957);
xnor U19079 (N_19079,N_16169,N_16475);
xnor U19080 (N_19080,N_17754,N_17327);
or U19081 (N_19081,N_17979,N_16551);
and U19082 (N_19082,N_17872,N_17119);
or U19083 (N_19083,N_16993,N_17115);
nor U19084 (N_19084,N_16934,N_17844);
nand U19085 (N_19085,N_16822,N_16346);
nand U19086 (N_19086,N_17265,N_17554);
xor U19087 (N_19087,N_16739,N_17191);
nor U19088 (N_19088,N_16422,N_17583);
or U19089 (N_19089,N_16416,N_16343);
nor U19090 (N_19090,N_16991,N_16581);
nand U19091 (N_19091,N_17064,N_16653);
nor U19092 (N_19092,N_17445,N_16740);
and U19093 (N_19093,N_17099,N_17845);
nand U19094 (N_19094,N_16990,N_17966);
or U19095 (N_19095,N_17873,N_17146);
or U19096 (N_19096,N_16520,N_17115);
and U19097 (N_19097,N_17473,N_16220);
nor U19098 (N_19098,N_17514,N_16730);
nor U19099 (N_19099,N_17208,N_17293);
and U19100 (N_19100,N_16347,N_17476);
or U19101 (N_19101,N_16803,N_17938);
nand U19102 (N_19102,N_17343,N_16234);
nand U19103 (N_19103,N_16814,N_16416);
nor U19104 (N_19104,N_17700,N_17772);
xor U19105 (N_19105,N_16770,N_16822);
xnor U19106 (N_19106,N_16211,N_16465);
nand U19107 (N_19107,N_16216,N_16115);
or U19108 (N_19108,N_16020,N_17848);
and U19109 (N_19109,N_16094,N_16606);
or U19110 (N_19110,N_16137,N_17770);
xnor U19111 (N_19111,N_16605,N_16058);
or U19112 (N_19112,N_17498,N_16156);
and U19113 (N_19113,N_16352,N_16963);
and U19114 (N_19114,N_16530,N_16206);
or U19115 (N_19115,N_17197,N_17486);
nand U19116 (N_19116,N_17355,N_16464);
xnor U19117 (N_19117,N_17615,N_16745);
nand U19118 (N_19118,N_17689,N_16625);
nand U19119 (N_19119,N_17501,N_16165);
xnor U19120 (N_19120,N_16084,N_16617);
nor U19121 (N_19121,N_17593,N_16358);
or U19122 (N_19122,N_17404,N_16465);
and U19123 (N_19123,N_17958,N_17189);
and U19124 (N_19124,N_17134,N_16124);
nand U19125 (N_19125,N_17675,N_17605);
and U19126 (N_19126,N_17524,N_16318);
xor U19127 (N_19127,N_17219,N_17779);
or U19128 (N_19128,N_17525,N_16360);
nor U19129 (N_19129,N_16853,N_17434);
or U19130 (N_19130,N_16025,N_16029);
nand U19131 (N_19131,N_17464,N_17619);
xnor U19132 (N_19132,N_17902,N_16522);
xnor U19133 (N_19133,N_17560,N_17541);
nand U19134 (N_19134,N_16894,N_17254);
xnor U19135 (N_19135,N_17064,N_16627);
and U19136 (N_19136,N_17057,N_16786);
xor U19137 (N_19137,N_16409,N_16594);
xnor U19138 (N_19138,N_16751,N_17319);
and U19139 (N_19139,N_16162,N_16700);
xnor U19140 (N_19140,N_16699,N_16152);
nand U19141 (N_19141,N_17672,N_17341);
nand U19142 (N_19142,N_17870,N_16107);
nor U19143 (N_19143,N_16056,N_16176);
and U19144 (N_19144,N_17878,N_17502);
xnor U19145 (N_19145,N_17954,N_16183);
nand U19146 (N_19146,N_17472,N_17878);
nand U19147 (N_19147,N_17225,N_17233);
or U19148 (N_19148,N_17300,N_17788);
nor U19149 (N_19149,N_17915,N_16102);
xor U19150 (N_19150,N_16665,N_16595);
and U19151 (N_19151,N_16497,N_16823);
and U19152 (N_19152,N_16498,N_17517);
nand U19153 (N_19153,N_17877,N_16563);
nor U19154 (N_19154,N_17236,N_17910);
and U19155 (N_19155,N_17743,N_16502);
xor U19156 (N_19156,N_16413,N_16950);
xnor U19157 (N_19157,N_16051,N_16480);
xnor U19158 (N_19158,N_17229,N_16838);
nor U19159 (N_19159,N_17135,N_16148);
and U19160 (N_19160,N_17539,N_17357);
nand U19161 (N_19161,N_17222,N_16424);
xnor U19162 (N_19162,N_17184,N_17338);
nand U19163 (N_19163,N_17234,N_16486);
or U19164 (N_19164,N_16750,N_17343);
nand U19165 (N_19165,N_16449,N_17307);
nor U19166 (N_19166,N_16210,N_16259);
xor U19167 (N_19167,N_17110,N_17986);
xor U19168 (N_19168,N_17827,N_16432);
nor U19169 (N_19169,N_17462,N_16718);
and U19170 (N_19170,N_16305,N_17891);
or U19171 (N_19171,N_17939,N_17519);
and U19172 (N_19172,N_16466,N_16556);
nand U19173 (N_19173,N_16564,N_17163);
or U19174 (N_19174,N_16160,N_16085);
or U19175 (N_19175,N_17520,N_17134);
or U19176 (N_19176,N_17798,N_16112);
nor U19177 (N_19177,N_16791,N_17988);
nand U19178 (N_19178,N_17561,N_17376);
and U19179 (N_19179,N_17229,N_17363);
or U19180 (N_19180,N_17060,N_16596);
and U19181 (N_19181,N_16055,N_17851);
and U19182 (N_19182,N_17791,N_17065);
nand U19183 (N_19183,N_17048,N_16925);
xnor U19184 (N_19184,N_17654,N_16089);
or U19185 (N_19185,N_17617,N_16590);
nor U19186 (N_19186,N_17228,N_17517);
or U19187 (N_19187,N_17324,N_17232);
nor U19188 (N_19188,N_16126,N_17639);
and U19189 (N_19189,N_17913,N_17772);
xnor U19190 (N_19190,N_17290,N_17779);
or U19191 (N_19191,N_17537,N_17017);
nor U19192 (N_19192,N_17198,N_16337);
nor U19193 (N_19193,N_17246,N_16600);
or U19194 (N_19194,N_17175,N_17763);
and U19195 (N_19195,N_16144,N_16649);
nand U19196 (N_19196,N_16630,N_16661);
or U19197 (N_19197,N_17829,N_17976);
xnor U19198 (N_19198,N_17409,N_17615);
xor U19199 (N_19199,N_16446,N_16777);
nand U19200 (N_19200,N_17255,N_16457);
xnor U19201 (N_19201,N_16193,N_17246);
and U19202 (N_19202,N_16847,N_16639);
nand U19203 (N_19203,N_16806,N_16284);
and U19204 (N_19204,N_17551,N_16321);
or U19205 (N_19205,N_17101,N_17479);
nor U19206 (N_19206,N_17662,N_17000);
xor U19207 (N_19207,N_16384,N_16096);
and U19208 (N_19208,N_16184,N_17047);
xnor U19209 (N_19209,N_17922,N_17422);
nor U19210 (N_19210,N_17851,N_16917);
nor U19211 (N_19211,N_16657,N_17630);
and U19212 (N_19212,N_16418,N_16324);
and U19213 (N_19213,N_17072,N_17149);
nor U19214 (N_19214,N_17491,N_17625);
or U19215 (N_19215,N_16647,N_16620);
and U19216 (N_19216,N_17382,N_17070);
or U19217 (N_19217,N_17114,N_16675);
xnor U19218 (N_19218,N_16476,N_16960);
nor U19219 (N_19219,N_17793,N_17045);
nand U19220 (N_19220,N_17954,N_16032);
and U19221 (N_19221,N_17771,N_17233);
or U19222 (N_19222,N_16012,N_17468);
nand U19223 (N_19223,N_17239,N_16942);
or U19224 (N_19224,N_16415,N_16229);
nand U19225 (N_19225,N_16092,N_17287);
or U19226 (N_19226,N_17918,N_16045);
and U19227 (N_19227,N_16322,N_17363);
nand U19228 (N_19228,N_16289,N_17013);
and U19229 (N_19229,N_16893,N_16287);
xor U19230 (N_19230,N_17897,N_16045);
or U19231 (N_19231,N_16500,N_16772);
nor U19232 (N_19232,N_16868,N_17398);
nor U19233 (N_19233,N_17672,N_17806);
and U19234 (N_19234,N_16640,N_16504);
nor U19235 (N_19235,N_16576,N_16778);
nor U19236 (N_19236,N_16713,N_16482);
nand U19237 (N_19237,N_17989,N_16598);
or U19238 (N_19238,N_17014,N_17195);
and U19239 (N_19239,N_17789,N_16115);
nand U19240 (N_19240,N_16438,N_16178);
nor U19241 (N_19241,N_16982,N_17259);
xor U19242 (N_19242,N_17017,N_17573);
or U19243 (N_19243,N_16870,N_17864);
and U19244 (N_19244,N_16913,N_16975);
or U19245 (N_19245,N_17014,N_16487);
nand U19246 (N_19246,N_17839,N_17879);
and U19247 (N_19247,N_16220,N_17299);
and U19248 (N_19248,N_17476,N_17639);
nand U19249 (N_19249,N_17471,N_16754);
and U19250 (N_19250,N_16085,N_16987);
and U19251 (N_19251,N_17878,N_16660);
and U19252 (N_19252,N_16327,N_16295);
xor U19253 (N_19253,N_16404,N_17752);
nor U19254 (N_19254,N_17317,N_17444);
and U19255 (N_19255,N_16049,N_16426);
nand U19256 (N_19256,N_17926,N_17334);
or U19257 (N_19257,N_16248,N_17978);
nor U19258 (N_19258,N_17907,N_16938);
nand U19259 (N_19259,N_16108,N_17941);
nor U19260 (N_19260,N_17452,N_17741);
and U19261 (N_19261,N_17880,N_17727);
xnor U19262 (N_19262,N_16116,N_17980);
and U19263 (N_19263,N_17545,N_16196);
xor U19264 (N_19264,N_16060,N_16969);
or U19265 (N_19265,N_16260,N_17978);
xor U19266 (N_19266,N_17704,N_16103);
and U19267 (N_19267,N_16928,N_17153);
nand U19268 (N_19268,N_16797,N_17857);
xnor U19269 (N_19269,N_17584,N_16162);
xor U19270 (N_19270,N_16647,N_16252);
xnor U19271 (N_19271,N_17401,N_17905);
nand U19272 (N_19272,N_16386,N_16385);
or U19273 (N_19273,N_16116,N_17687);
nor U19274 (N_19274,N_17975,N_17005);
nor U19275 (N_19275,N_17270,N_17669);
xor U19276 (N_19276,N_17595,N_16171);
and U19277 (N_19277,N_17378,N_16876);
xor U19278 (N_19278,N_17342,N_16829);
and U19279 (N_19279,N_16334,N_17126);
xnor U19280 (N_19280,N_17973,N_16317);
nand U19281 (N_19281,N_17794,N_17143);
or U19282 (N_19282,N_16470,N_17357);
and U19283 (N_19283,N_16246,N_17585);
and U19284 (N_19284,N_17683,N_16470);
and U19285 (N_19285,N_16728,N_17193);
xnor U19286 (N_19286,N_16639,N_16955);
nand U19287 (N_19287,N_16766,N_17067);
and U19288 (N_19288,N_17311,N_17847);
nand U19289 (N_19289,N_16167,N_17657);
or U19290 (N_19290,N_16131,N_17999);
xor U19291 (N_19291,N_16457,N_17033);
or U19292 (N_19292,N_16834,N_17379);
nand U19293 (N_19293,N_16868,N_17244);
xor U19294 (N_19294,N_16768,N_17916);
nand U19295 (N_19295,N_17569,N_16620);
xnor U19296 (N_19296,N_17817,N_17384);
and U19297 (N_19297,N_17976,N_16505);
or U19298 (N_19298,N_17981,N_17430);
nor U19299 (N_19299,N_17778,N_17185);
nand U19300 (N_19300,N_17314,N_16015);
nor U19301 (N_19301,N_16338,N_16801);
nand U19302 (N_19302,N_17711,N_16949);
and U19303 (N_19303,N_16484,N_17680);
nand U19304 (N_19304,N_16848,N_17712);
nor U19305 (N_19305,N_17175,N_16464);
nor U19306 (N_19306,N_16428,N_16469);
nor U19307 (N_19307,N_16671,N_17468);
or U19308 (N_19308,N_17022,N_16566);
xor U19309 (N_19309,N_16587,N_16995);
or U19310 (N_19310,N_16840,N_17981);
xor U19311 (N_19311,N_17229,N_16987);
nor U19312 (N_19312,N_17108,N_16093);
nor U19313 (N_19313,N_17106,N_16643);
nand U19314 (N_19314,N_17385,N_16054);
and U19315 (N_19315,N_16692,N_17740);
nor U19316 (N_19316,N_16799,N_16305);
and U19317 (N_19317,N_16440,N_17424);
or U19318 (N_19318,N_17793,N_17170);
and U19319 (N_19319,N_17396,N_16736);
nand U19320 (N_19320,N_16722,N_17211);
nand U19321 (N_19321,N_16735,N_16690);
xor U19322 (N_19322,N_17303,N_17959);
nor U19323 (N_19323,N_16072,N_16425);
and U19324 (N_19324,N_17121,N_17388);
nand U19325 (N_19325,N_17519,N_16626);
nand U19326 (N_19326,N_16948,N_16473);
nor U19327 (N_19327,N_17880,N_17370);
and U19328 (N_19328,N_17165,N_17517);
and U19329 (N_19329,N_17486,N_16525);
xor U19330 (N_19330,N_17503,N_16643);
nor U19331 (N_19331,N_16218,N_17533);
or U19332 (N_19332,N_16882,N_17054);
or U19333 (N_19333,N_17668,N_17300);
and U19334 (N_19334,N_16963,N_16801);
or U19335 (N_19335,N_17970,N_17684);
xnor U19336 (N_19336,N_16764,N_16760);
and U19337 (N_19337,N_16678,N_16861);
xor U19338 (N_19338,N_17399,N_16417);
nor U19339 (N_19339,N_16712,N_16683);
or U19340 (N_19340,N_17847,N_16825);
or U19341 (N_19341,N_17962,N_16309);
nand U19342 (N_19342,N_16266,N_16997);
nand U19343 (N_19343,N_17585,N_17527);
or U19344 (N_19344,N_16307,N_16124);
and U19345 (N_19345,N_17264,N_16618);
nor U19346 (N_19346,N_16571,N_17046);
xor U19347 (N_19347,N_17113,N_17606);
xor U19348 (N_19348,N_17363,N_17739);
xnor U19349 (N_19349,N_17483,N_16057);
xor U19350 (N_19350,N_17790,N_17578);
and U19351 (N_19351,N_16120,N_17751);
and U19352 (N_19352,N_17564,N_17426);
nand U19353 (N_19353,N_17338,N_17698);
nand U19354 (N_19354,N_17919,N_17166);
and U19355 (N_19355,N_16458,N_16453);
and U19356 (N_19356,N_17988,N_16259);
and U19357 (N_19357,N_16728,N_17255);
nor U19358 (N_19358,N_17593,N_16518);
nand U19359 (N_19359,N_17259,N_17729);
or U19360 (N_19360,N_17469,N_16707);
xnor U19361 (N_19361,N_16844,N_17988);
nand U19362 (N_19362,N_16150,N_17917);
and U19363 (N_19363,N_16458,N_17211);
xor U19364 (N_19364,N_16297,N_16319);
and U19365 (N_19365,N_16726,N_16122);
and U19366 (N_19366,N_17741,N_16730);
and U19367 (N_19367,N_17333,N_17252);
xnor U19368 (N_19368,N_17579,N_16146);
nand U19369 (N_19369,N_17406,N_16212);
xor U19370 (N_19370,N_17490,N_16028);
or U19371 (N_19371,N_16844,N_17140);
and U19372 (N_19372,N_17276,N_16298);
and U19373 (N_19373,N_16078,N_17138);
or U19374 (N_19374,N_16482,N_16505);
nand U19375 (N_19375,N_16508,N_17517);
xnor U19376 (N_19376,N_17241,N_16932);
xnor U19377 (N_19377,N_16875,N_17325);
nand U19378 (N_19378,N_17549,N_16115);
nor U19379 (N_19379,N_16918,N_17741);
nor U19380 (N_19380,N_17905,N_16681);
or U19381 (N_19381,N_16851,N_17054);
nor U19382 (N_19382,N_16196,N_17373);
xor U19383 (N_19383,N_16539,N_17204);
nand U19384 (N_19384,N_17206,N_17106);
and U19385 (N_19385,N_17440,N_16738);
xor U19386 (N_19386,N_16204,N_16595);
and U19387 (N_19387,N_17775,N_17081);
xnor U19388 (N_19388,N_16142,N_17266);
or U19389 (N_19389,N_16832,N_16610);
xnor U19390 (N_19390,N_16043,N_17981);
or U19391 (N_19391,N_17375,N_16820);
or U19392 (N_19392,N_17985,N_17092);
nor U19393 (N_19393,N_17684,N_16914);
or U19394 (N_19394,N_16101,N_16085);
or U19395 (N_19395,N_17136,N_17986);
xnor U19396 (N_19396,N_17596,N_17385);
or U19397 (N_19397,N_17210,N_16865);
nor U19398 (N_19398,N_16898,N_16356);
and U19399 (N_19399,N_16121,N_16128);
nand U19400 (N_19400,N_16816,N_16334);
xor U19401 (N_19401,N_16024,N_16266);
or U19402 (N_19402,N_17479,N_17340);
and U19403 (N_19403,N_16053,N_16716);
nor U19404 (N_19404,N_16595,N_16459);
nand U19405 (N_19405,N_17762,N_17051);
nor U19406 (N_19406,N_16289,N_16419);
and U19407 (N_19407,N_17041,N_16526);
nor U19408 (N_19408,N_16461,N_17136);
nor U19409 (N_19409,N_17362,N_16456);
or U19410 (N_19410,N_17352,N_17847);
nor U19411 (N_19411,N_16898,N_16598);
xor U19412 (N_19412,N_16554,N_17763);
xnor U19413 (N_19413,N_16244,N_17260);
nand U19414 (N_19414,N_16941,N_17403);
nor U19415 (N_19415,N_16613,N_17144);
and U19416 (N_19416,N_17961,N_17690);
nor U19417 (N_19417,N_17473,N_17288);
nand U19418 (N_19418,N_16351,N_16358);
and U19419 (N_19419,N_16688,N_16442);
nand U19420 (N_19420,N_17286,N_17566);
and U19421 (N_19421,N_17385,N_16343);
nand U19422 (N_19422,N_17562,N_16183);
xor U19423 (N_19423,N_17466,N_17994);
or U19424 (N_19424,N_16083,N_17855);
nor U19425 (N_19425,N_16174,N_16318);
and U19426 (N_19426,N_17538,N_16772);
nor U19427 (N_19427,N_17216,N_16752);
and U19428 (N_19428,N_16369,N_17183);
and U19429 (N_19429,N_16978,N_16412);
xnor U19430 (N_19430,N_17824,N_16746);
xor U19431 (N_19431,N_16742,N_17544);
or U19432 (N_19432,N_17982,N_17731);
nor U19433 (N_19433,N_17403,N_16665);
nand U19434 (N_19434,N_17150,N_17367);
xnor U19435 (N_19435,N_16972,N_17885);
nand U19436 (N_19436,N_16096,N_17186);
nor U19437 (N_19437,N_16599,N_17728);
nor U19438 (N_19438,N_17223,N_16286);
nand U19439 (N_19439,N_17750,N_17554);
or U19440 (N_19440,N_16900,N_16159);
xnor U19441 (N_19441,N_16455,N_17366);
and U19442 (N_19442,N_17603,N_17172);
xnor U19443 (N_19443,N_16091,N_17158);
or U19444 (N_19444,N_17534,N_17643);
or U19445 (N_19445,N_17222,N_17056);
and U19446 (N_19446,N_16673,N_16561);
xor U19447 (N_19447,N_17986,N_16449);
or U19448 (N_19448,N_17503,N_17076);
and U19449 (N_19449,N_17973,N_16824);
and U19450 (N_19450,N_16825,N_17942);
nand U19451 (N_19451,N_17054,N_17969);
and U19452 (N_19452,N_16145,N_16319);
nand U19453 (N_19453,N_17880,N_16157);
xor U19454 (N_19454,N_16483,N_17172);
xor U19455 (N_19455,N_17734,N_17571);
nor U19456 (N_19456,N_17872,N_16447);
or U19457 (N_19457,N_17104,N_17589);
nand U19458 (N_19458,N_17502,N_16646);
nand U19459 (N_19459,N_16132,N_17806);
or U19460 (N_19460,N_16790,N_17289);
and U19461 (N_19461,N_16894,N_17641);
xor U19462 (N_19462,N_16554,N_17020);
nand U19463 (N_19463,N_16234,N_17818);
and U19464 (N_19464,N_16036,N_16667);
nand U19465 (N_19465,N_17927,N_16623);
nand U19466 (N_19466,N_16940,N_17991);
nor U19467 (N_19467,N_17602,N_17977);
or U19468 (N_19468,N_16629,N_17396);
nand U19469 (N_19469,N_16015,N_17542);
and U19470 (N_19470,N_16742,N_17569);
nand U19471 (N_19471,N_16001,N_17274);
or U19472 (N_19472,N_16066,N_16129);
and U19473 (N_19473,N_16044,N_17152);
nor U19474 (N_19474,N_17782,N_16067);
nor U19475 (N_19475,N_17934,N_16220);
and U19476 (N_19476,N_16647,N_17447);
or U19477 (N_19477,N_16424,N_17119);
nor U19478 (N_19478,N_17892,N_16147);
nand U19479 (N_19479,N_17743,N_16322);
or U19480 (N_19480,N_17683,N_16947);
nand U19481 (N_19481,N_17620,N_16332);
nor U19482 (N_19482,N_16462,N_17334);
or U19483 (N_19483,N_17005,N_16324);
or U19484 (N_19484,N_17300,N_16093);
xnor U19485 (N_19485,N_17515,N_17393);
and U19486 (N_19486,N_17416,N_16029);
nor U19487 (N_19487,N_17130,N_16069);
nand U19488 (N_19488,N_17860,N_17999);
xnor U19489 (N_19489,N_16715,N_16777);
nand U19490 (N_19490,N_16947,N_17107);
xor U19491 (N_19491,N_17981,N_17183);
nor U19492 (N_19492,N_16733,N_17658);
nand U19493 (N_19493,N_17866,N_16748);
xor U19494 (N_19494,N_17227,N_17889);
xor U19495 (N_19495,N_17983,N_16355);
or U19496 (N_19496,N_16075,N_16610);
nor U19497 (N_19497,N_16713,N_17018);
and U19498 (N_19498,N_16403,N_16844);
nor U19499 (N_19499,N_16448,N_16329);
and U19500 (N_19500,N_16918,N_17372);
nand U19501 (N_19501,N_16791,N_17121);
nor U19502 (N_19502,N_16354,N_17607);
and U19503 (N_19503,N_17778,N_16876);
and U19504 (N_19504,N_17030,N_16520);
nand U19505 (N_19505,N_17677,N_16050);
nor U19506 (N_19506,N_16277,N_16658);
nor U19507 (N_19507,N_16850,N_17562);
nand U19508 (N_19508,N_16168,N_16172);
and U19509 (N_19509,N_16884,N_17428);
xnor U19510 (N_19510,N_17299,N_17226);
xnor U19511 (N_19511,N_16781,N_16114);
xnor U19512 (N_19512,N_17056,N_17177);
xor U19513 (N_19513,N_16029,N_16717);
nor U19514 (N_19514,N_17124,N_17474);
or U19515 (N_19515,N_17345,N_16332);
xnor U19516 (N_19516,N_16875,N_16010);
and U19517 (N_19517,N_16101,N_17220);
or U19518 (N_19518,N_16436,N_16570);
nor U19519 (N_19519,N_17718,N_16904);
xor U19520 (N_19520,N_17284,N_17631);
and U19521 (N_19521,N_17288,N_17914);
xor U19522 (N_19522,N_17337,N_16955);
nand U19523 (N_19523,N_17308,N_16995);
or U19524 (N_19524,N_17442,N_17555);
nor U19525 (N_19525,N_17266,N_17470);
or U19526 (N_19526,N_16165,N_16178);
xnor U19527 (N_19527,N_17120,N_17301);
nand U19528 (N_19528,N_16427,N_16698);
xor U19529 (N_19529,N_17865,N_16643);
nand U19530 (N_19530,N_16513,N_16866);
xnor U19531 (N_19531,N_17613,N_17014);
nand U19532 (N_19532,N_16631,N_17161);
or U19533 (N_19533,N_16980,N_16680);
xnor U19534 (N_19534,N_17755,N_16836);
and U19535 (N_19535,N_17437,N_16205);
nor U19536 (N_19536,N_17043,N_17330);
and U19537 (N_19537,N_17818,N_17276);
nand U19538 (N_19538,N_17643,N_17042);
nor U19539 (N_19539,N_16576,N_16017);
xnor U19540 (N_19540,N_17907,N_17870);
and U19541 (N_19541,N_16124,N_17675);
nand U19542 (N_19542,N_17832,N_17113);
xor U19543 (N_19543,N_16086,N_16595);
nand U19544 (N_19544,N_16588,N_16711);
and U19545 (N_19545,N_17664,N_17315);
and U19546 (N_19546,N_17702,N_16700);
nand U19547 (N_19547,N_17108,N_17635);
xor U19548 (N_19548,N_16748,N_17484);
nand U19549 (N_19549,N_16285,N_16564);
and U19550 (N_19550,N_16907,N_17543);
nand U19551 (N_19551,N_17673,N_16538);
or U19552 (N_19552,N_16393,N_16663);
nor U19553 (N_19553,N_16146,N_17950);
nor U19554 (N_19554,N_17259,N_17483);
nor U19555 (N_19555,N_17052,N_17562);
xor U19556 (N_19556,N_17329,N_16819);
and U19557 (N_19557,N_17550,N_17070);
nand U19558 (N_19558,N_16174,N_16822);
nand U19559 (N_19559,N_17909,N_16383);
or U19560 (N_19560,N_17580,N_17823);
nand U19561 (N_19561,N_16084,N_16880);
nor U19562 (N_19562,N_16927,N_16690);
or U19563 (N_19563,N_17536,N_16001);
or U19564 (N_19564,N_17815,N_16253);
nor U19565 (N_19565,N_17004,N_16208);
nor U19566 (N_19566,N_16226,N_17478);
or U19567 (N_19567,N_16524,N_17606);
nor U19568 (N_19568,N_16424,N_17489);
nand U19569 (N_19569,N_16382,N_17608);
nand U19570 (N_19570,N_16452,N_16466);
or U19571 (N_19571,N_17910,N_17836);
xnor U19572 (N_19572,N_16101,N_16066);
nand U19573 (N_19573,N_17689,N_16549);
nor U19574 (N_19574,N_16939,N_16278);
nand U19575 (N_19575,N_16703,N_17871);
and U19576 (N_19576,N_17341,N_16671);
or U19577 (N_19577,N_17964,N_16260);
or U19578 (N_19578,N_16418,N_17045);
and U19579 (N_19579,N_16474,N_17536);
xor U19580 (N_19580,N_16156,N_17004);
nor U19581 (N_19581,N_17678,N_17822);
or U19582 (N_19582,N_16811,N_17366);
or U19583 (N_19583,N_17895,N_16217);
xnor U19584 (N_19584,N_17389,N_16198);
nor U19585 (N_19585,N_16264,N_16605);
and U19586 (N_19586,N_17018,N_17105);
xor U19587 (N_19587,N_16490,N_16984);
xor U19588 (N_19588,N_16914,N_17820);
or U19589 (N_19589,N_16619,N_16183);
nor U19590 (N_19590,N_17656,N_17021);
nor U19591 (N_19591,N_16788,N_17209);
nand U19592 (N_19592,N_17053,N_17806);
or U19593 (N_19593,N_17698,N_17553);
or U19594 (N_19594,N_17174,N_17417);
or U19595 (N_19595,N_16102,N_16216);
or U19596 (N_19596,N_16534,N_16024);
nor U19597 (N_19597,N_16815,N_16939);
or U19598 (N_19598,N_17387,N_16767);
or U19599 (N_19599,N_16139,N_17052);
xor U19600 (N_19600,N_16837,N_16937);
nand U19601 (N_19601,N_16774,N_16605);
xor U19602 (N_19602,N_16686,N_16729);
nand U19603 (N_19603,N_16434,N_16793);
xor U19604 (N_19604,N_17882,N_16342);
xor U19605 (N_19605,N_16353,N_16446);
nor U19606 (N_19606,N_16764,N_16484);
nor U19607 (N_19607,N_16890,N_17881);
or U19608 (N_19608,N_16722,N_16625);
and U19609 (N_19609,N_16013,N_17630);
and U19610 (N_19610,N_17800,N_17623);
nor U19611 (N_19611,N_17877,N_17760);
and U19612 (N_19612,N_17473,N_17296);
xnor U19613 (N_19613,N_16320,N_17311);
and U19614 (N_19614,N_16831,N_17764);
nand U19615 (N_19615,N_17310,N_17983);
xor U19616 (N_19616,N_16766,N_16591);
or U19617 (N_19617,N_16643,N_17149);
nand U19618 (N_19618,N_17226,N_17772);
and U19619 (N_19619,N_16988,N_17260);
nand U19620 (N_19620,N_16995,N_16996);
nand U19621 (N_19621,N_17152,N_16043);
nor U19622 (N_19622,N_16788,N_17257);
and U19623 (N_19623,N_17273,N_17372);
or U19624 (N_19624,N_17452,N_16226);
nor U19625 (N_19625,N_16504,N_17628);
nand U19626 (N_19626,N_16136,N_17423);
or U19627 (N_19627,N_17872,N_16092);
nand U19628 (N_19628,N_17652,N_16065);
xor U19629 (N_19629,N_16822,N_16898);
nor U19630 (N_19630,N_17028,N_16120);
xnor U19631 (N_19631,N_17445,N_16508);
xnor U19632 (N_19632,N_17518,N_17520);
or U19633 (N_19633,N_17986,N_17195);
nand U19634 (N_19634,N_16805,N_16501);
and U19635 (N_19635,N_16443,N_16996);
nand U19636 (N_19636,N_17737,N_16701);
or U19637 (N_19637,N_16566,N_17609);
xor U19638 (N_19638,N_16350,N_17649);
xnor U19639 (N_19639,N_16991,N_16053);
or U19640 (N_19640,N_16326,N_17384);
xor U19641 (N_19641,N_16479,N_17319);
nor U19642 (N_19642,N_16387,N_16852);
nor U19643 (N_19643,N_17324,N_16017);
and U19644 (N_19644,N_16561,N_17446);
or U19645 (N_19645,N_16137,N_16555);
nor U19646 (N_19646,N_17740,N_16269);
and U19647 (N_19647,N_17119,N_16223);
or U19648 (N_19648,N_16933,N_17452);
and U19649 (N_19649,N_17408,N_16618);
nand U19650 (N_19650,N_17076,N_16140);
or U19651 (N_19651,N_17339,N_17486);
or U19652 (N_19652,N_16843,N_16187);
nor U19653 (N_19653,N_17718,N_16757);
xnor U19654 (N_19654,N_16396,N_17436);
nand U19655 (N_19655,N_17239,N_16861);
and U19656 (N_19656,N_17687,N_16471);
nor U19657 (N_19657,N_16804,N_17749);
nand U19658 (N_19658,N_17173,N_16524);
or U19659 (N_19659,N_16184,N_16322);
xnor U19660 (N_19660,N_17400,N_17825);
and U19661 (N_19661,N_17996,N_17777);
nor U19662 (N_19662,N_17751,N_17583);
xor U19663 (N_19663,N_16912,N_16160);
xor U19664 (N_19664,N_17784,N_16242);
nand U19665 (N_19665,N_16580,N_17841);
nor U19666 (N_19666,N_16842,N_17058);
and U19667 (N_19667,N_16322,N_16881);
nor U19668 (N_19668,N_17955,N_17965);
nand U19669 (N_19669,N_17090,N_16871);
xor U19670 (N_19670,N_17472,N_16015);
xor U19671 (N_19671,N_16665,N_17346);
nand U19672 (N_19672,N_16884,N_17203);
xor U19673 (N_19673,N_16616,N_16392);
nand U19674 (N_19674,N_17571,N_17644);
nor U19675 (N_19675,N_17500,N_17244);
nor U19676 (N_19676,N_17157,N_17944);
nor U19677 (N_19677,N_17791,N_16752);
or U19678 (N_19678,N_17581,N_16552);
xor U19679 (N_19679,N_16035,N_17529);
and U19680 (N_19680,N_16011,N_17095);
nand U19681 (N_19681,N_16472,N_16242);
xnor U19682 (N_19682,N_16583,N_16000);
or U19683 (N_19683,N_17991,N_17435);
and U19684 (N_19684,N_17255,N_17534);
nand U19685 (N_19685,N_16501,N_17107);
nand U19686 (N_19686,N_16690,N_16779);
or U19687 (N_19687,N_16719,N_17766);
xnor U19688 (N_19688,N_16640,N_17507);
xor U19689 (N_19689,N_17791,N_17543);
and U19690 (N_19690,N_16697,N_16570);
nand U19691 (N_19691,N_17581,N_16884);
and U19692 (N_19692,N_17600,N_16246);
nand U19693 (N_19693,N_17880,N_17719);
and U19694 (N_19694,N_16215,N_17204);
nand U19695 (N_19695,N_17873,N_16466);
or U19696 (N_19696,N_17993,N_16925);
nor U19697 (N_19697,N_16471,N_17879);
nor U19698 (N_19698,N_17876,N_16039);
xnor U19699 (N_19699,N_17535,N_16267);
nor U19700 (N_19700,N_16786,N_17088);
xnor U19701 (N_19701,N_16753,N_16229);
nor U19702 (N_19702,N_17749,N_16111);
and U19703 (N_19703,N_17011,N_16316);
or U19704 (N_19704,N_16428,N_16165);
xor U19705 (N_19705,N_16892,N_17607);
nor U19706 (N_19706,N_17322,N_17733);
or U19707 (N_19707,N_17436,N_17594);
and U19708 (N_19708,N_16457,N_16632);
and U19709 (N_19709,N_17504,N_17647);
nor U19710 (N_19710,N_17634,N_16221);
nand U19711 (N_19711,N_16338,N_17623);
nor U19712 (N_19712,N_16658,N_16827);
and U19713 (N_19713,N_17500,N_16012);
nand U19714 (N_19714,N_17007,N_17852);
and U19715 (N_19715,N_16845,N_17655);
or U19716 (N_19716,N_16650,N_17961);
and U19717 (N_19717,N_16467,N_16216);
nand U19718 (N_19718,N_16030,N_17691);
xor U19719 (N_19719,N_16818,N_17556);
xnor U19720 (N_19720,N_16565,N_17671);
nor U19721 (N_19721,N_17100,N_17034);
or U19722 (N_19722,N_16458,N_16424);
xor U19723 (N_19723,N_17013,N_17435);
or U19724 (N_19724,N_16215,N_16448);
xor U19725 (N_19725,N_16413,N_16416);
or U19726 (N_19726,N_16507,N_16626);
nand U19727 (N_19727,N_16076,N_16220);
nand U19728 (N_19728,N_17414,N_17673);
nor U19729 (N_19729,N_17579,N_16845);
or U19730 (N_19730,N_16059,N_17544);
xor U19731 (N_19731,N_16648,N_17951);
nor U19732 (N_19732,N_16156,N_17605);
nand U19733 (N_19733,N_16545,N_17240);
xnor U19734 (N_19734,N_17962,N_16670);
and U19735 (N_19735,N_16890,N_17791);
and U19736 (N_19736,N_17451,N_17878);
nor U19737 (N_19737,N_16565,N_16543);
nand U19738 (N_19738,N_16504,N_17115);
or U19739 (N_19739,N_16374,N_17604);
nand U19740 (N_19740,N_16973,N_16827);
and U19741 (N_19741,N_16347,N_16081);
and U19742 (N_19742,N_16380,N_17936);
or U19743 (N_19743,N_16455,N_16643);
or U19744 (N_19744,N_16821,N_17045);
or U19745 (N_19745,N_16591,N_16390);
xnor U19746 (N_19746,N_17473,N_17709);
or U19747 (N_19747,N_17365,N_16302);
nand U19748 (N_19748,N_17291,N_16246);
or U19749 (N_19749,N_16391,N_16644);
or U19750 (N_19750,N_17321,N_17852);
or U19751 (N_19751,N_16258,N_16737);
and U19752 (N_19752,N_16408,N_16451);
nand U19753 (N_19753,N_16686,N_17553);
nand U19754 (N_19754,N_16519,N_17358);
nor U19755 (N_19755,N_16215,N_17027);
xnor U19756 (N_19756,N_17816,N_16401);
or U19757 (N_19757,N_17401,N_17847);
xnor U19758 (N_19758,N_17272,N_17575);
and U19759 (N_19759,N_17700,N_17351);
xor U19760 (N_19760,N_16920,N_16905);
or U19761 (N_19761,N_16393,N_16207);
nor U19762 (N_19762,N_17791,N_17135);
nand U19763 (N_19763,N_17114,N_17597);
nor U19764 (N_19764,N_16318,N_17515);
nand U19765 (N_19765,N_16798,N_17758);
nand U19766 (N_19766,N_16661,N_17363);
nand U19767 (N_19767,N_16139,N_17759);
xor U19768 (N_19768,N_17448,N_17249);
xor U19769 (N_19769,N_17549,N_17152);
nand U19770 (N_19770,N_16069,N_16293);
nor U19771 (N_19771,N_17845,N_17497);
or U19772 (N_19772,N_17889,N_17239);
xnor U19773 (N_19773,N_16755,N_17264);
or U19774 (N_19774,N_16819,N_17403);
nor U19775 (N_19775,N_16517,N_17591);
and U19776 (N_19776,N_16567,N_16065);
xor U19777 (N_19777,N_17940,N_16386);
or U19778 (N_19778,N_17692,N_17414);
or U19779 (N_19779,N_17236,N_17383);
nand U19780 (N_19780,N_17892,N_16252);
xor U19781 (N_19781,N_16667,N_16356);
and U19782 (N_19782,N_16585,N_16570);
nor U19783 (N_19783,N_16501,N_17801);
nor U19784 (N_19784,N_17159,N_16640);
xor U19785 (N_19785,N_16846,N_17054);
or U19786 (N_19786,N_16579,N_16958);
xnor U19787 (N_19787,N_16396,N_17977);
and U19788 (N_19788,N_16338,N_16071);
xnor U19789 (N_19789,N_16880,N_16236);
or U19790 (N_19790,N_17451,N_16519);
nor U19791 (N_19791,N_16729,N_16397);
nor U19792 (N_19792,N_17161,N_16646);
or U19793 (N_19793,N_17265,N_16836);
and U19794 (N_19794,N_17456,N_17444);
xor U19795 (N_19795,N_17234,N_17167);
nand U19796 (N_19796,N_16188,N_17372);
or U19797 (N_19797,N_17415,N_17540);
xnor U19798 (N_19798,N_17698,N_16938);
xor U19799 (N_19799,N_16159,N_17657);
nor U19800 (N_19800,N_17510,N_17828);
and U19801 (N_19801,N_16168,N_17604);
nor U19802 (N_19802,N_16789,N_17532);
nand U19803 (N_19803,N_17159,N_17095);
or U19804 (N_19804,N_17670,N_17361);
or U19805 (N_19805,N_16344,N_17088);
and U19806 (N_19806,N_17557,N_16024);
nand U19807 (N_19807,N_17141,N_16858);
or U19808 (N_19808,N_16016,N_17009);
and U19809 (N_19809,N_16085,N_16729);
nor U19810 (N_19810,N_16990,N_16883);
or U19811 (N_19811,N_17955,N_16226);
nand U19812 (N_19812,N_16447,N_17395);
nand U19813 (N_19813,N_16940,N_17452);
or U19814 (N_19814,N_16793,N_16247);
or U19815 (N_19815,N_16948,N_16300);
or U19816 (N_19816,N_17562,N_16189);
nor U19817 (N_19817,N_17539,N_16858);
nand U19818 (N_19818,N_16879,N_16903);
nor U19819 (N_19819,N_17739,N_17585);
or U19820 (N_19820,N_16701,N_17918);
and U19821 (N_19821,N_17068,N_16991);
or U19822 (N_19822,N_16272,N_17331);
or U19823 (N_19823,N_16676,N_16632);
or U19824 (N_19824,N_17393,N_16054);
and U19825 (N_19825,N_16409,N_17011);
nor U19826 (N_19826,N_16545,N_16345);
nor U19827 (N_19827,N_17419,N_16555);
nor U19828 (N_19828,N_16429,N_16330);
and U19829 (N_19829,N_17465,N_17890);
xnor U19830 (N_19830,N_17284,N_17157);
and U19831 (N_19831,N_16790,N_16015);
xnor U19832 (N_19832,N_17697,N_17958);
xor U19833 (N_19833,N_17813,N_16112);
nand U19834 (N_19834,N_16134,N_17702);
nand U19835 (N_19835,N_16754,N_17439);
nand U19836 (N_19836,N_17918,N_16881);
xnor U19837 (N_19837,N_16252,N_17120);
xnor U19838 (N_19838,N_16436,N_16120);
xor U19839 (N_19839,N_17104,N_17553);
and U19840 (N_19840,N_16318,N_16443);
or U19841 (N_19841,N_16967,N_17252);
or U19842 (N_19842,N_16349,N_16087);
or U19843 (N_19843,N_17541,N_16603);
xor U19844 (N_19844,N_16612,N_16371);
nand U19845 (N_19845,N_16241,N_16024);
or U19846 (N_19846,N_16771,N_17892);
or U19847 (N_19847,N_16866,N_17706);
nand U19848 (N_19848,N_16577,N_17146);
xnor U19849 (N_19849,N_17045,N_17085);
xor U19850 (N_19850,N_16322,N_17849);
nor U19851 (N_19851,N_17199,N_17466);
xnor U19852 (N_19852,N_17922,N_17217);
or U19853 (N_19853,N_16867,N_17909);
nand U19854 (N_19854,N_16306,N_16196);
and U19855 (N_19855,N_16779,N_17488);
or U19856 (N_19856,N_17420,N_16000);
nand U19857 (N_19857,N_17547,N_16424);
or U19858 (N_19858,N_16068,N_17639);
nor U19859 (N_19859,N_16442,N_17980);
or U19860 (N_19860,N_17591,N_17537);
and U19861 (N_19861,N_17409,N_17108);
nand U19862 (N_19862,N_16876,N_16642);
nor U19863 (N_19863,N_17536,N_16832);
nor U19864 (N_19864,N_17648,N_17345);
and U19865 (N_19865,N_17776,N_16953);
or U19866 (N_19866,N_17245,N_17441);
nor U19867 (N_19867,N_16476,N_16332);
nor U19868 (N_19868,N_16317,N_17476);
nand U19869 (N_19869,N_17623,N_16957);
and U19870 (N_19870,N_17385,N_16944);
nand U19871 (N_19871,N_16087,N_16527);
nand U19872 (N_19872,N_17134,N_17946);
and U19873 (N_19873,N_16891,N_16669);
and U19874 (N_19874,N_16778,N_16548);
xnor U19875 (N_19875,N_16364,N_16422);
or U19876 (N_19876,N_17538,N_17596);
or U19877 (N_19877,N_16071,N_17198);
or U19878 (N_19878,N_17453,N_16194);
nand U19879 (N_19879,N_16286,N_17770);
nand U19880 (N_19880,N_17774,N_17676);
xor U19881 (N_19881,N_17329,N_17451);
or U19882 (N_19882,N_16187,N_16830);
or U19883 (N_19883,N_16566,N_17016);
nand U19884 (N_19884,N_17090,N_17013);
nand U19885 (N_19885,N_16754,N_17905);
or U19886 (N_19886,N_16763,N_16772);
and U19887 (N_19887,N_16618,N_16858);
nand U19888 (N_19888,N_17736,N_16956);
nor U19889 (N_19889,N_16583,N_16569);
xor U19890 (N_19890,N_17242,N_16620);
nand U19891 (N_19891,N_16237,N_16012);
nand U19892 (N_19892,N_16573,N_17139);
nand U19893 (N_19893,N_16954,N_17879);
nand U19894 (N_19894,N_16669,N_16555);
nand U19895 (N_19895,N_17004,N_16908);
or U19896 (N_19896,N_17685,N_17014);
nand U19897 (N_19897,N_16445,N_16416);
nor U19898 (N_19898,N_16329,N_17654);
and U19899 (N_19899,N_17281,N_17221);
and U19900 (N_19900,N_17647,N_16290);
nand U19901 (N_19901,N_17205,N_16100);
or U19902 (N_19902,N_16200,N_17484);
or U19903 (N_19903,N_16025,N_16083);
nand U19904 (N_19904,N_17055,N_16851);
nor U19905 (N_19905,N_17979,N_16958);
xnor U19906 (N_19906,N_17476,N_17307);
nand U19907 (N_19907,N_16991,N_16469);
nor U19908 (N_19908,N_17604,N_16626);
or U19909 (N_19909,N_16530,N_17386);
or U19910 (N_19910,N_16332,N_16613);
or U19911 (N_19911,N_16478,N_17108);
or U19912 (N_19912,N_17405,N_16145);
nand U19913 (N_19913,N_17750,N_17405);
or U19914 (N_19914,N_16375,N_17989);
xnor U19915 (N_19915,N_16835,N_16248);
or U19916 (N_19916,N_16148,N_17970);
and U19917 (N_19917,N_17273,N_17966);
xnor U19918 (N_19918,N_17627,N_16734);
xnor U19919 (N_19919,N_17915,N_17950);
and U19920 (N_19920,N_16419,N_16948);
and U19921 (N_19921,N_17689,N_16961);
nand U19922 (N_19922,N_16100,N_16819);
nand U19923 (N_19923,N_17022,N_17757);
xnor U19924 (N_19924,N_16520,N_17716);
nand U19925 (N_19925,N_17142,N_17094);
xor U19926 (N_19926,N_16507,N_16470);
nor U19927 (N_19927,N_17983,N_16673);
nand U19928 (N_19928,N_17352,N_17720);
and U19929 (N_19929,N_17520,N_16486);
or U19930 (N_19930,N_17973,N_16933);
or U19931 (N_19931,N_16585,N_16463);
xnor U19932 (N_19932,N_17381,N_17284);
nor U19933 (N_19933,N_16307,N_17315);
and U19934 (N_19934,N_16886,N_17534);
or U19935 (N_19935,N_17382,N_17665);
nor U19936 (N_19936,N_16280,N_17519);
nor U19937 (N_19937,N_17905,N_17445);
or U19938 (N_19938,N_16378,N_17983);
xor U19939 (N_19939,N_16537,N_17800);
or U19940 (N_19940,N_17106,N_17759);
nand U19941 (N_19941,N_16444,N_16282);
nor U19942 (N_19942,N_16996,N_17169);
xnor U19943 (N_19943,N_16622,N_17438);
or U19944 (N_19944,N_16763,N_16314);
nor U19945 (N_19945,N_17700,N_16294);
or U19946 (N_19946,N_16182,N_16731);
nand U19947 (N_19947,N_16144,N_16787);
and U19948 (N_19948,N_16967,N_17583);
or U19949 (N_19949,N_17709,N_16560);
or U19950 (N_19950,N_16322,N_16982);
xor U19951 (N_19951,N_17687,N_16605);
xnor U19952 (N_19952,N_16653,N_16881);
xnor U19953 (N_19953,N_17674,N_16075);
nor U19954 (N_19954,N_16910,N_16895);
or U19955 (N_19955,N_16257,N_16471);
nand U19956 (N_19956,N_16447,N_16073);
and U19957 (N_19957,N_16458,N_17640);
or U19958 (N_19958,N_17505,N_16245);
and U19959 (N_19959,N_17918,N_17105);
or U19960 (N_19960,N_16820,N_17541);
and U19961 (N_19961,N_16021,N_17588);
xnor U19962 (N_19962,N_17418,N_16534);
nand U19963 (N_19963,N_16066,N_17962);
nand U19964 (N_19964,N_16069,N_16308);
nor U19965 (N_19965,N_16951,N_17449);
nand U19966 (N_19966,N_16850,N_16507);
nor U19967 (N_19967,N_17733,N_16506);
nand U19968 (N_19968,N_16016,N_16435);
xor U19969 (N_19969,N_16219,N_17255);
and U19970 (N_19970,N_17886,N_16960);
or U19971 (N_19971,N_16044,N_17257);
xor U19972 (N_19972,N_16994,N_17402);
and U19973 (N_19973,N_16575,N_17473);
and U19974 (N_19974,N_17003,N_16150);
nor U19975 (N_19975,N_17368,N_17926);
nor U19976 (N_19976,N_17322,N_16179);
nand U19977 (N_19977,N_16758,N_17774);
nor U19978 (N_19978,N_16621,N_17668);
and U19979 (N_19979,N_16881,N_16950);
or U19980 (N_19980,N_17055,N_16470);
nand U19981 (N_19981,N_17357,N_16426);
nand U19982 (N_19982,N_17709,N_17941);
and U19983 (N_19983,N_17899,N_17444);
nor U19984 (N_19984,N_16176,N_16672);
or U19985 (N_19985,N_16198,N_16098);
xor U19986 (N_19986,N_16789,N_16749);
and U19987 (N_19987,N_17799,N_17414);
xor U19988 (N_19988,N_17649,N_17881);
and U19989 (N_19989,N_16406,N_16994);
nor U19990 (N_19990,N_16735,N_17879);
or U19991 (N_19991,N_17913,N_16401);
xnor U19992 (N_19992,N_17141,N_16957);
nor U19993 (N_19993,N_17809,N_17970);
nor U19994 (N_19994,N_16895,N_17290);
nand U19995 (N_19995,N_16017,N_16700);
nand U19996 (N_19996,N_16978,N_17728);
or U19997 (N_19997,N_16670,N_17232);
or U19998 (N_19998,N_17333,N_16263);
nor U19999 (N_19999,N_16045,N_17692);
xor UO_0 (O_0,N_19449,N_18446);
or UO_1 (O_1,N_19269,N_18009);
or UO_2 (O_2,N_19111,N_19530);
or UO_3 (O_3,N_18260,N_19287);
or UO_4 (O_4,N_18371,N_18325);
nand UO_5 (O_5,N_19288,N_19725);
or UO_6 (O_6,N_19778,N_19254);
and UO_7 (O_7,N_19233,N_18410);
or UO_8 (O_8,N_19826,N_18581);
xor UO_9 (O_9,N_18298,N_18011);
nor UO_10 (O_10,N_18555,N_19391);
xnor UO_11 (O_11,N_18820,N_18074);
nand UO_12 (O_12,N_19546,N_19856);
nor UO_13 (O_13,N_19389,N_18908);
nor UO_14 (O_14,N_19251,N_19790);
nor UO_15 (O_15,N_19944,N_18360);
nor UO_16 (O_16,N_18996,N_18274);
and UO_17 (O_17,N_19306,N_19132);
and UO_18 (O_18,N_18015,N_19216);
nor UO_19 (O_19,N_18923,N_18247);
nor UO_20 (O_20,N_19866,N_18070);
xnor UO_21 (O_21,N_18078,N_18183);
and UO_22 (O_22,N_18541,N_18758);
nor UO_23 (O_23,N_19584,N_19550);
and UO_24 (O_24,N_18327,N_18077);
nor UO_25 (O_25,N_19358,N_19068);
or UO_26 (O_26,N_19548,N_19788);
or UO_27 (O_27,N_18817,N_18320);
or UO_28 (O_28,N_18664,N_19632);
or UO_29 (O_29,N_18357,N_18135);
and UO_30 (O_30,N_18699,N_18189);
nor UO_31 (O_31,N_18290,N_19424);
and UO_32 (O_32,N_18493,N_18337);
xnor UO_33 (O_33,N_18958,N_19884);
and UO_34 (O_34,N_18711,N_18466);
or UO_35 (O_35,N_19119,N_18725);
nand UO_36 (O_36,N_19112,N_19137);
nor UO_37 (O_37,N_18947,N_19334);
or UO_38 (O_38,N_18782,N_18252);
or UO_39 (O_39,N_18429,N_19455);
nor UO_40 (O_40,N_18995,N_18838);
or UO_41 (O_41,N_18791,N_19409);
xnor UO_42 (O_42,N_19145,N_19036);
and UO_43 (O_43,N_19074,N_19158);
or UO_44 (O_44,N_18764,N_19598);
xnor UO_45 (O_45,N_19395,N_18677);
and UO_46 (O_46,N_18729,N_18308);
nand UO_47 (O_47,N_19559,N_19753);
and UO_48 (O_48,N_18738,N_18959);
or UO_49 (O_49,N_19961,N_19760);
nor UO_50 (O_50,N_19766,N_18380);
xor UO_51 (O_51,N_18319,N_19755);
or UO_52 (O_52,N_19918,N_19450);
and UO_53 (O_53,N_19983,N_18673);
xor UO_54 (O_54,N_18229,N_19237);
and UO_55 (O_55,N_18770,N_18355);
xor UO_56 (O_56,N_19714,N_19190);
xnor UO_57 (O_57,N_19321,N_19581);
nand UO_58 (O_58,N_18113,N_19654);
or UO_59 (O_59,N_19602,N_19017);
or UO_60 (O_60,N_19862,N_18747);
and UO_61 (O_61,N_19996,N_18472);
and UO_62 (O_62,N_18259,N_18579);
nor UO_63 (O_63,N_19451,N_18656);
xnor UO_64 (O_64,N_18629,N_19404);
and UO_65 (O_65,N_18519,N_19730);
or UO_66 (O_66,N_19098,N_18220);
nor UO_67 (O_67,N_19255,N_18846);
and UO_68 (O_68,N_18815,N_18151);
nand UO_69 (O_69,N_19023,N_18407);
nor UO_70 (O_70,N_18148,N_18652);
nor UO_71 (O_71,N_18690,N_18640);
xor UO_72 (O_72,N_19894,N_19720);
or UO_73 (O_73,N_19244,N_18241);
or UO_74 (O_74,N_18988,N_19301);
or UO_75 (O_75,N_19200,N_19828);
nand UO_76 (O_76,N_18623,N_18287);
nand UO_77 (O_77,N_19292,N_19590);
xnor UO_78 (O_78,N_19011,N_18695);
xnor UO_79 (O_79,N_19470,N_18864);
nor UO_80 (O_80,N_19136,N_19263);
xnor UO_81 (O_81,N_18423,N_19250);
and UO_82 (O_82,N_18731,N_18847);
nand UO_83 (O_83,N_19049,N_18588);
and UO_84 (O_84,N_18683,N_19796);
xnor UO_85 (O_85,N_19600,N_19012);
or UO_86 (O_86,N_18089,N_19882);
nand UO_87 (O_87,N_18885,N_18515);
xor UO_88 (O_88,N_18524,N_19733);
and UO_89 (O_89,N_19507,N_19718);
nor UO_90 (O_90,N_19296,N_18055);
nand UO_91 (O_91,N_19658,N_18426);
nand UO_92 (O_92,N_19503,N_19184);
nand UO_93 (O_93,N_19523,N_18072);
xnor UO_94 (O_94,N_19784,N_18806);
or UO_95 (O_95,N_19633,N_19312);
and UO_96 (O_96,N_18253,N_19577);
and UO_97 (O_97,N_19278,N_18296);
and UO_98 (O_98,N_19282,N_18457);
or UO_99 (O_99,N_19643,N_18217);
nand UO_100 (O_100,N_18102,N_18739);
nor UO_101 (O_101,N_18542,N_18348);
xnor UO_102 (O_102,N_18293,N_18850);
nand UO_103 (O_103,N_18223,N_19813);
nand UO_104 (O_104,N_18147,N_18053);
xnor UO_105 (O_105,N_18018,N_18076);
xor UO_106 (O_106,N_19138,N_18309);
and UO_107 (O_107,N_18970,N_19483);
or UO_108 (O_108,N_19479,N_18992);
nor UO_109 (O_109,N_19147,N_19408);
and UO_110 (O_110,N_18586,N_19426);
nand UO_111 (O_111,N_19226,N_18757);
nand UO_112 (O_112,N_19497,N_19436);
or UO_113 (O_113,N_18462,N_18924);
and UO_114 (O_114,N_19195,N_18709);
xor UO_115 (O_115,N_18300,N_18152);
or UO_116 (O_116,N_19139,N_19231);
or UO_117 (O_117,N_18932,N_19955);
xor UO_118 (O_118,N_18544,N_19360);
or UO_119 (O_119,N_19751,N_18759);
or UO_120 (O_120,N_18655,N_19325);
xor UO_121 (O_121,N_19780,N_19355);
nand UO_122 (O_122,N_19171,N_18352);
and UO_123 (O_123,N_19401,N_18827);
nor UO_124 (O_124,N_19261,N_18632);
nor UO_125 (O_125,N_19574,N_19934);
nand UO_126 (O_126,N_18546,N_18798);
and UO_127 (O_127,N_18349,N_19242);
xor UO_128 (O_128,N_18278,N_19880);
xor UO_129 (O_129,N_19843,N_19765);
and UO_130 (O_130,N_19326,N_18245);
xnor UO_131 (O_131,N_18843,N_19384);
or UO_132 (O_132,N_19700,N_18029);
nand UO_133 (O_133,N_18963,N_18103);
or UO_134 (O_134,N_19383,N_18477);
nor UO_135 (O_135,N_18935,N_19063);
xor UO_136 (O_136,N_18956,N_18765);
xnor UO_137 (O_137,N_19810,N_19965);
xor UO_138 (O_138,N_19073,N_18143);
nand UO_139 (O_139,N_19474,N_18511);
and UO_140 (O_140,N_18538,N_18284);
or UO_141 (O_141,N_18505,N_19442);
and UO_142 (O_142,N_18039,N_19217);
xor UO_143 (O_143,N_18645,N_19086);
or UO_144 (O_144,N_19797,N_19125);
and UO_145 (O_145,N_18985,N_18498);
nand UO_146 (O_146,N_19427,N_18949);
nor UO_147 (O_147,N_19169,N_18957);
xor UO_148 (O_148,N_19123,N_19560);
or UO_149 (O_149,N_19986,N_19623);
and UO_150 (O_150,N_18481,N_19709);
nand UO_151 (O_151,N_18385,N_18227);
and UO_152 (O_152,N_18574,N_19281);
or UO_153 (O_153,N_18326,N_18510);
nand UO_154 (O_154,N_19743,N_18315);
nand UO_155 (O_155,N_19890,N_18177);
and UO_156 (O_156,N_18350,N_18697);
xor UO_157 (O_157,N_18431,N_19363);
nor UO_158 (O_158,N_19656,N_19435);
nand UO_159 (O_159,N_18718,N_18445);
xor UO_160 (O_160,N_18624,N_19738);
nand UO_161 (O_161,N_18210,N_18618);
and UO_162 (O_162,N_18744,N_19844);
and UO_163 (O_163,N_18473,N_18083);
nor UO_164 (O_164,N_19247,N_19614);
nor UO_165 (O_165,N_18316,N_19886);
and UO_166 (O_166,N_19798,N_18080);
xor UO_167 (O_167,N_18133,N_19518);
and UO_168 (O_168,N_18037,N_19815);
nand UO_169 (O_169,N_18363,N_19445);
or UO_170 (O_170,N_18937,N_19601);
xor UO_171 (O_171,N_19239,N_18318);
or UO_172 (O_172,N_18863,N_19531);
or UO_173 (O_173,N_18277,N_19650);
nand UO_174 (O_174,N_19716,N_18345);
nor UO_175 (O_175,N_18386,N_19877);
nor UO_176 (O_176,N_18688,N_19888);
and UO_177 (O_177,N_19723,N_19500);
or UO_178 (O_178,N_18031,N_19154);
xnor UO_179 (O_179,N_19291,N_18601);
nor UO_180 (O_180,N_19144,N_18006);
or UO_181 (O_181,N_19431,N_18399);
or UO_182 (O_182,N_18328,N_18366);
or UO_183 (O_183,N_18915,N_18035);
and UO_184 (O_184,N_18365,N_19839);
or UO_185 (O_185,N_19127,N_19083);
or UO_186 (O_186,N_18767,N_19998);
and UO_187 (O_187,N_19094,N_18983);
or UO_188 (O_188,N_18897,N_18132);
nor UO_189 (O_189,N_19447,N_19202);
nor UO_190 (O_190,N_18818,N_19690);
xor UO_191 (O_191,N_19003,N_19979);
or UO_192 (O_192,N_18666,N_19108);
nor UO_193 (O_193,N_19628,N_19543);
nor UO_194 (O_194,N_19100,N_18156);
nor UO_195 (O_195,N_19051,N_18643);
or UO_196 (O_196,N_18192,N_18911);
nand UO_197 (O_197,N_18403,N_19759);
or UO_198 (O_198,N_18000,N_19230);
xor UO_199 (O_199,N_18974,N_19113);
or UO_200 (O_200,N_19569,N_18454);
nor UO_201 (O_201,N_19433,N_18107);
and UO_202 (O_202,N_19864,N_18990);
nor UO_203 (O_203,N_18310,N_19679);
xnor UO_204 (O_204,N_18548,N_18794);
nand UO_205 (O_205,N_18166,N_18531);
and UO_206 (O_206,N_19176,N_19423);
and UO_207 (O_207,N_18153,N_18237);
nor UO_208 (O_208,N_19993,N_18880);
and UO_209 (O_209,N_18458,N_19150);
xor UO_210 (O_210,N_19583,N_19077);
and UO_211 (O_211,N_19564,N_19678);
xor UO_212 (O_212,N_19280,N_18727);
nor UO_213 (O_213,N_19731,N_19453);
xor UO_214 (O_214,N_18435,N_18048);
or UO_215 (O_215,N_19624,N_18614);
nor UO_216 (O_216,N_19960,N_18594);
nand UO_217 (O_217,N_18825,N_18225);
xor UO_218 (O_218,N_19914,N_19345);
nor UO_219 (O_219,N_18517,N_19201);
and UO_220 (O_220,N_18194,N_18672);
and UO_221 (O_221,N_19014,N_19713);
or UO_222 (O_222,N_18181,N_19735);
xnor UO_223 (O_223,N_18188,N_19367);
xnor UO_224 (O_224,N_19323,N_19018);
or UO_225 (O_225,N_18002,N_19681);
or UO_226 (O_226,N_19505,N_19495);
xnor UO_227 (O_227,N_18321,N_18495);
nand UO_228 (O_228,N_19517,N_18874);
nand UO_229 (O_229,N_18397,N_18859);
and UO_230 (O_230,N_18788,N_19361);
nand UO_231 (O_231,N_18136,N_18636);
xor UO_232 (O_232,N_18617,N_19277);
xnor UO_233 (O_233,N_18269,N_19131);
nand UO_234 (O_234,N_18370,N_19124);
nand UO_235 (O_235,N_19508,N_18719);
nor UO_236 (O_236,N_18020,N_18175);
nand UO_237 (O_237,N_18250,N_19787);
xor UO_238 (O_238,N_18613,N_19067);
and UO_239 (O_239,N_19210,N_18134);
nor UO_240 (O_240,N_19982,N_18082);
xor UO_241 (O_241,N_18242,N_19529);
xnor UO_242 (O_242,N_19472,N_19331);
and UO_243 (O_243,N_19706,N_18966);
or UO_244 (O_244,N_19480,N_19163);
nand UO_245 (O_245,N_19610,N_19398);
nand UO_246 (O_246,N_19902,N_18249);
xnor UO_247 (O_247,N_18030,N_18761);
nand UO_248 (O_248,N_18584,N_18630);
or UO_249 (O_249,N_18282,N_18648);
xor UO_250 (O_250,N_18131,N_18987);
nor UO_251 (O_251,N_18808,N_18170);
xor UO_252 (O_252,N_19421,N_19207);
and UO_253 (O_253,N_18696,N_18060);
nand UO_254 (O_254,N_19537,N_19005);
xnor UO_255 (O_255,N_19981,N_19392);
nand UO_256 (O_256,N_19803,N_19310);
nand UO_257 (O_257,N_18575,N_18722);
or UO_258 (O_258,N_18221,N_19318);
xor UO_259 (O_259,N_18101,N_18207);
or UO_260 (O_260,N_18989,N_19985);
nand UO_261 (O_261,N_18219,N_18839);
and UO_262 (O_262,N_18805,N_18778);
nor UO_263 (O_263,N_19910,N_18663);
nor UO_264 (O_264,N_19314,N_19061);
xor UO_265 (O_265,N_19465,N_19443);
or UO_266 (O_266,N_18649,N_19037);
and UO_267 (O_267,N_18781,N_18596);
nand UO_268 (O_268,N_19348,N_18377);
and UO_269 (O_269,N_19873,N_18669);
nor UO_270 (O_270,N_18324,N_19079);
nor UO_271 (O_271,N_19043,N_18138);
and UO_272 (O_272,N_18291,N_18639);
nor UO_273 (O_273,N_18085,N_19867);
xor UO_274 (O_274,N_19002,N_19387);
nor UO_275 (O_275,N_19557,N_19140);
nand UO_276 (O_276,N_18023,N_18787);
nand UO_277 (O_277,N_18314,N_18773);
or UO_278 (O_278,N_18341,N_18208);
or UO_279 (O_279,N_18705,N_18566);
nor UO_280 (O_280,N_19305,N_18137);
nand UO_281 (O_281,N_18496,N_18154);
xor UO_282 (O_282,N_18523,N_18396);
and UO_283 (O_283,N_18028,N_18465);
and UO_284 (O_284,N_19736,N_19861);
and UO_285 (O_285,N_19257,N_19177);
and UO_286 (O_286,N_19708,N_19703);
xnor UO_287 (O_287,N_19109,N_18046);
xnor UO_288 (O_288,N_19126,N_18860);
nor UO_289 (O_289,N_18793,N_19309);
and UO_290 (O_290,N_19252,N_18740);
and UO_291 (O_291,N_18530,N_18772);
and UO_292 (O_292,N_19594,N_19904);
xnor UO_293 (O_293,N_19031,N_18003);
xnor UO_294 (O_294,N_19938,N_18200);
nand UO_295 (O_295,N_19354,N_18280);
nor UO_296 (O_296,N_19820,N_18368);
xnor UO_297 (O_297,N_19368,N_19576);
or UO_298 (O_298,N_19419,N_19072);
xor UO_299 (O_299,N_19804,N_18126);
nor UO_300 (O_300,N_18901,N_18164);
xnor UO_301 (O_301,N_19940,N_19382);
nand UO_302 (O_302,N_18275,N_18411);
xnor UO_303 (O_303,N_18312,N_19498);
xor UO_304 (O_304,N_19157,N_19117);
nor UO_305 (O_305,N_19087,N_18338);
nor UO_306 (O_306,N_18886,N_18842);
xnor UO_307 (O_307,N_19726,N_19997);
nor UO_308 (O_308,N_18563,N_18243);
nand UO_309 (O_309,N_19621,N_18564);
or UO_310 (O_310,N_19041,N_19187);
and UO_311 (O_311,N_19189,N_19053);
and UO_312 (O_312,N_18950,N_19829);
or UO_313 (O_313,N_19327,N_19204);
and UO_314 (O_314,N_18329,N_19402);
and UO_315 (O_315,N_19651,N_19511);
or UO_316 (O_316,N_19089,N_19777);
or UO_317 (O_317,N_18230,N_18882);
xnor UO_318 (O_318,N_19212,N_19352);
nor UO_319 (O_319,N_19967,N_19313);
or UO_320 (O_320,N_18942,N_18551);
and UO_321 (O_321,N_19871,N_19710);
and UO_322 (O_322,N_18822,N_19227);
or UO_323 (O_323,N_18255,N_19071);
nor UO_324 (O_324,N_18807,N_18813);
nand UO_325 (O_325,N_19812,N_18344);
nor UO_326 (O_326,N_18869,N_19728);
xor UO_327 (O_327,N_19417,N_18733);
nor UO_328 (O_328,N_19460,N_18169);
or UO_329 (O_329,N_18797,N_19028);
nand UO_330 (O_330,N_18266,N_19040);
nor UO_331 (O_331,N_19928,N_19682);
and UO_332 (O_332,N_19616,N_19478);
xnor UO_333 (O_333,N_18647,N_19711);
nor UO_334 (O_334,N_18065,N_18215);
xnor UO_335 (O_335,N_19283,N_19380);
xor UO_336 (O_336,N_19185,N_19534);
or UO_337 (O_337,N_18257,N_19146);
and UO_338 (O_338,N_18706,N_18038);
or UO_339 (O_339,N_18714,N_19636);
xor UO_340 (O_340,N_18339,N_19842);
nor UO_341 (O_341,N_19851,N_18689);
and UO_342 (O_342,N_18660,N_18894);
and UO_343 (O_343,N_18883,N_19625);
nor UO_344 (O_344,N_19399,N_19205);
nor UO_345 (O_345,N_19547,N_19410);
nand UO_346 (O_346,N_18490,N_19042);
or UO_347 (O_347,N_19865,N_18091);
and UO_348 (O_348,N_19980,N_19764);
xnor UO_349 (O_349,N_18022,N_19400);
xor UO_350 (O_350,N_18111,N_19156);
and UO_351 (O_351,N_18346,N_18703);
xor UO_352 (O_352,N_18354,N_19892);
or UO_353 (O_353,N_18866,N_19987);
or UO_354 (O_354,N_19704,N_19935);
and UO_355 (O_355,N_18340,N_19836);
or UO_356 (O_356,N_18216,N_18067);
nor UO_357 (O_357,N_18606,N_18394);
nor UO_358 (O_358,N_19954,N_18891);
and UO_359 (O_359,N_19162,N_18094);
nand UO_360 (O_360,N_18603,N_18191);
and UO_361 (O_361,N_18066,N_18088);
nand UO_362 (O_362,N_19452,N_18514);
nor UO_363 (O_363,N_19817,N_19415);
and UO_364 (O_364,N_18736,N_19129);
or UO_365 (O_365,N_19622,N_19418);
and UO_366 (O_366,N_19091,N_19270);
nor UO_367 (O_367,N_18383,N_19665);
xnor UO_368 (O_368,N_19193,N_19330);
and UO_369 (O_369,N_18218,N_18910);
nor UO_370 (O_370,N_19732,N_19153);
or UO_371 (O_371,N_19805,N_19082);
nor UO_372 (O_372,N_18299,N_18508);
xnor UO_373 (O_373,N_18425,N_18779);
nor UO_374 (O_374,N_18984,N_19640);
and UO_375 (O_375,N_18125,N_19208);
and UO_376 (O_376,N_18141,N_19487);
xnor UO_377 (O_377,N_19824,N_18941);
xor UO_378 (O_378,N_19223,N_19744);
or UO_379 (O_379,N_18934,N_18019);
nor UO_380 (O_380,N_19613,N_19057);
and UO_381 (O_381,N_19661,N_18206);
nand UO_382 (O_382,N_18059,N_18240);
nand UO_383 (O_383,N_19416,N_18816);
and UO_384 (O_384,N_19775,N_18750);
or UO_385 (O_385,N_18422,N_19976);
nor UO_386 (O_386,N_18185,N_18971);
xor UO_387 (O_387,N_19385,N_18993);
or UO_388 (O_388,N_19350,N_18145);
or UO_389 (O_389,N_19722,N_18627);
or UO_390 (O_390,N_18746,N_18372);
nor UO_391 (O_391,N_18420,N_18605);
xnor UO_392 (O_392,N_19274,N_18232);
nor UO_393 (O_393,N_18917,N_19490);
nand UO_394 (O_394,N_19845,N_19930);
or UO_395 (O_395,N_18121,N_19170);
xnor UO_396 (O_396,N_18187,N_19116);
or UO_397 (O_397,N_18569,N_18359);
or UO_398 (O_398,N_18671,N_18246);
and UO_399 (O_399,N_19906,N_19852);
and UO_400 (O_400,N_19901,N_19816);
nand UO_401 (O_401,N_18186,N_18196);
nand UO_402 (O_402,N_18879,N_19868);
or UO_403 (O_403,N_19933,N_18854);
or UO_404 (O_404,N_18592,N_18506);
xnor UO_405 (O_405,N_19062,N_19923);
and UO_406 (O_406,N_18600,N_18635);
nand UO_407 (O_407,N_19249,N_18682);
or UO_408 (O_408,N_18491,N_18751);
nand UO_409 (O_409,N_19475,N_18093);
or UO_410 (O_410,N_18953,N_18991);
and UO_411 (O_411,N_19376,N_18898);
or UO_412 (O_412,N_18497,N_19821);
nand UO_413 (O_413,N_19526,N_19078);
nor UO_414 (O_414,N_18589,N_18862);
nor UO_415 (O_415,N_19586,N_19235);
nor UO_416 (O_416,N_19060,N_19908);
and UO_417 (O_417,N_18610,N_18155);
nor UO_418 (O_418,N_19687,N_19595);
nor UO_419 (O_419,N_18783,N_18033);
or UO_420 (O_420,N_19454,N_18693);
nor UO_421 (O_421,N_19489,N_19858);
or UO_422 (O_422,N_19631,N_18962);
nand UO_423 (O_423,N_18373,N_18844);
nand UO_424 (O_424,N_18071,N_19811);
nor UO_425 (O_425,N_18471,N_18443);
xor UO_426 (O_426,N_19717,N_18453);
nand UO_427 (O_427,N_18001,N_19224);
nor UO_428 (O_428,N_18470,N_19657);
or UO_429 (O_429,N_19048,N_18870);
nor UO_430 (O_430,N_19397,N_18620);
nand UO_431 (O_431,N_19587,N_18812);
nor UO_432 (O_432,N_19357,N_19152);
nand UO_433 (O_433,N_18478,N_19855);
xnor UO_434 (O_434,N_19022,N_19101);
and UO_435 (O_435,N_18042,N_18374);
and UO_436 (O_436,N_18118,N_19029);
nor UO_437 (O_437,N_18896,N_18149);
nand UO_438 (O_438,N_18073,N_18480);
nor UO_439 (O_439,N_18097,N_18486);
and UO_440 (O_440,N_19192,N_19971);
nand UO_441 (O_441,N_18796,N_18721);
nand UO_442 (O_442,N_18052,N_19374);
nor UO_443 (O_443,N_18233,N_18434);
xnor UO_444 (O_444,N_18356,N_19070);
nor UO_445 (O_445,N_19552,N_19693);
and UO_446 (O_446,N_18641,N_18301);
and UO_447 (O_447,N_19333,N_18529);
nand UO_448 (O_448,N_18754,N_18025);
nand UO_449 (O_449,N_18040,N_19501);
xor UO_450 (O_450,N_19860,N_18675);
or UO_451 (O_451,N_19608,N_18938);
or UO_452 (O_452,N_19461,N_19729);
nor UO_453 (O_453,N_18939,N_19411);
nor UO_454 (O_454,N_19335,N_19106);
nand UO_455 (O_455,N_18205,N_19444);
or UO_456 (O_456,N_19551,N_19630);
nand UO_457 (O_457,N_18388,N_19471);
nand UO_458 (O_458,N_18167,N_18068);
nor UO_459 (O_459,N_18769,N_19970);
nand UO_460 (O_460,N_19521,N_18313);
xor UO_461 (O_461,N_19995,N_18840);
xnor UO_462 (O_462,N_18182,N_18157);
nor UO_463 (O_463,N_19064,N_19853);
or UO_464 (O_464,N_18853,N_19883);
xor UO_465 (O_465,N_18877,N_19258);
or UO_466 (O_466,N_18027,N_18484);
and UO_467 (O_467,N_19915,N_18447);
or UO_468 (O_468,N_19105,N_19248);
xnor UO_469 (O_469,N_19857,N_19545);
or UO_470 (O_470,N_18428,N_19832);
nor UO_471 (O_471,N_18800,N_18317);
nor UO_472 (O_472,N_19683,N_18214);
nand UO_473 (O_473,N_19527,N_18213);
nor UO_474 (O_474,N_19702,N_18527);
and UO_475 (O_475,N_19434,N_19835);
nor UO_476 (O_476,N_18836,N_18903);
or UO_477 (O_477,N_18804,N_19662);
or UO_478 (O_478,N_18451,N_18295);
nand UO_479 (O_479,N_18165,N_18916);
nor UO_480 (O_480,N_18026,N_18464);
xnor UO_481 (O_481,N_19677,N_19808);
nand UO_482 (O_482,N_19615,N_19128);
and UO_483 (O_483,N_18438,N_18092);
nand UO_484 (O_484,N_18568,N_18599);
or UO_485 (O_485,N_19689,N_18271);
and UO_486 (O_486,N_19893,N_18159);
nor UO_487 (O_487,N_18051,N_19834);
xnor UO_488 (O_488,N_19038,N_18235);
and UO_489 (O_489,N_19715,N_19298);
or UO_490 (O_490,N_19294,N_19688);
or UO_491 (O_491,N_19311,N_19180);
and UO_492 (O_492,N_18920,N_18814);
or UO_493 (O_493,N_19055,N_18848);
nor UO_494 (O_494,N_19191,N_19203);
xnor UO_495 (O_495,N_18698,N_19491);
nor UO_496 (O_496,N_18264,N_18565);
nand UO_497 (O_497,N_18406,N_19076);
nand UO_498 (O_498,N_18913,N_19343);
and UO_499 (O_499,N_19114,N_19482);
nand UO_500 (O_500,N_19197,N_19638);
xor UO_501 (O_501,N_19641,N_19155);
xor UO_502 (O_502,N_18774,N_18289);
nor UO_503 (O_503,N_18980,N_19440);
xor UO_504 (O_504,N_19992,N_18681);
and UO_505 (O_505,N_19238,N_18554);
and UO_506 (O_506,N_18732,N_18829);
or UO_507 (O_507,N_18276,N_19562);
nor UO_508 (O_508,N_18461,N_18710);
or UO_509 (O_509,N_19379,N_19373);
or UO_510 (O_510,N_19909,N_19695);
nor UO_511 (O_511,N_19936,N_19182);
and UO_512 (O_512,N_19618,N_18571);
xor UO_513 (O_513,N_19222,N_19611);
xnor UO_514 (O_514,N_18239,N_19634);
xor UO_515 (O_515,N_18590,N_18286);
xor UO_516 (O_516,N_19916,N_18526);
nor UO_517 (O_517,N_19351,N_18268);
and UO_518 (O_518,N_18109,N_18890);
nand UO_519 (O_519,N_18171,N_18168);
nand UO_520 (O_520,N_18528,N_19603);
and UO_521 (O_521,N_19456,N_19667);
or UO_522 (O_522,N_19990,N_19822);
xor UO_523 (O_523,N_18199,N_19302);
or UO_524 (O_524,N_18906,N_18771);
and UO_525 (O_525,N_19299,N_18389);
and UO_526 (O_526,N_18516,N_18922);
nor UO_527 (O_527,N_18621,N_18550);
and UO_528 (O_528,N_19267,N_19556);
and UO_529 (O_529,N_19605,N_19342);
and UO_530 (O_530,N_18504,N_19196);
nor UO_531 (O_531,N_18595,N_19554);
nor UO_532 (O_532,N_18545,N_19568);
nor UO_533 (O_533,N_18408,N_18330);
xor UO_534 (O_534,N_18598,N_19206);
xnor UO_535 (O_535,N_18492,N_18304);
or UO_536 (O_536,N_19308,N_18105);
xnor UO_537 (O_537,N_18198,N_18534);
or UO_538 (O_538,N_18176,N_19831);
or UO_539 (O_539,N_18972,N_19046);
and UO_540 (O_540,N_18212,N_18343);
and UO_541 (O_541,N_19705,N_18888);
or UO_542 (O_542,N_19340,N_19422);
or UO_543 (O_543,N_19540,N_18261);
and UO_544 (O_544,N_18331,N_18743);
or UO_545 (O_545,N_19737,N_18591);
or UO_546 (O_546,N_19653,N_18904);
nor UO_547 (O_547,N_18895,N_18307);
xor UO_548 (O_548,N_19473,N_19900);
nor UO_549 (O_549,N_19359,N_18892);
xnor UO_550 (O_550,N_18998,N_18455);
and UO_551 (O_551,N_18283,N_18401);
nand UO_552 (O_552,N_19807,N_19052);
nand UO_553 (O_553,N_19019,N_18694);
xnor UO_554 (O_554,N_18918,N_19649);
xnor UO_555 (O_555,N_18982,N_19927);
nand UO_556 (O_556,N_19365,N_19265);
nor UO_557 (O_557,N_19289,N_19015);
or UO_558 (O_558,N_19823,N_19209);
nand UO_559 (O_559,N_19830,N_18961);
or UO_560 (O_560,N_19538,N_18726);
nor UO_561 (O_561,N_19951,N_19260);
nand UO_562 (O_562,N_19789,N_18440);
xnor UO_563 (O_563,N_19520,N_19898);
xor UO_564 (O_564,N_18512,N_19448);
or UO_565 (O_565,N_18098,N_19591);
xnor UO_566 (O_566,N_18604,N_18116);
nor UO_567 (O_567,N_18919,N_19942);
or UO_568 (O_568,N_19428,N_19854);
nor UO_569 (O_569,N_18755,N_18079);
nand UO_570 (O_570,N_18108,N_18122);
or UO_571 (O_571,N_18659,N_19167);
nor UO_572 (O_572,N_18433,N_19093);
or UO_573 (O_573,N_18479,N_19872);
nor UO_574 (O_574,N_18358,N_19008);
nor UO_575 (O_575,N_18872,N_19972);
or UO_576 (O_576,N_19840,N_19390);
or UO_577 (O_577,N_18832,N_18900);
or UO_578 (O_578,N_18752,N_18775);
nand UO_579 (O_579,N_18158,N_19774);
nor UO_580 (O_580,N_19887,N_19950);
nand UO_581 (O_581,N_19425,N_19604);
or UO_582 (O_582,N_19194,N_18790);
and UO_583 (O_583,N_18567,N_18871);
nand UO_584 (O_584,N_19370,N_18190);
nor UO_585 (O_585,N_18238,N_18625);
or UO_586 (O_586,N_18997,N_19025);
and UO_587 (O_587,N_19637,N_19499);
and UO_588 (O_588,N_18267,N_18821);
xor UO_589 (O_589,N_18146,N_18851);
and UO_590 (O_590,N_18943,N_18611);
or UO_591 (O_591,N_19420,N_18562);
xnor UO_592 (O_592,N_19000,N_18849);
nor UO_593 (O_593,N_18819,N_19555);
or UO_594 (O_594,N_19437,N_18593);
and UO_595 (O_595,N_19045,N_19246);
xor UO_596 (O_596,N_19462,N_19988);
and UO_597 (O_597,N_18050,N_18008);
nor UO_598 (O_598,N_18704,N_18834);
nor UO_599 (O_599,N_19477,N_18303);
or UO_600 (O_600,N_18734,N_19234);
or UO_601 (O_601,N_19148,N_18557);
or UO_602 (O_602,N_19859,N_19050);
nand UO_603 (O_603,N_18224,N_19758);
xnor UO_604 (O_604,N_18856,N_19782);
xnor UO_605 (O_605,N_18717,N_18075);
nor UO_606 (O_606,N_19570,N_19671);
or UO_607 (O_607,N_18855,N_19572);
and UO_608 (O_608,N_19596,N_19752);
xnor UO_609 (O_609,N_19549,N_18256);
nand UO_610 (O_610,N_19999,N_18114);
xor UO_611 (O_611,N_18297,N_19514);
and UO_612 (O_612,N_19791,N_19949);
and UO_613 (O_613,N_18502,N_19142);
nor UO_614 (O_614,N_19806,N_18905);
or UO_615 (O_615,N_18835,N_18522);
or UO_616 (O_616,N_19745,N_19103);
xor UO_617 (O_617,N_18081,N_18865);
or UO_618 (O_618,N_18150,N_19488);
nor UO_619 (O_619,N_18202,N_18485);
nand UO_620 (O_620,N_18715,N_18533);
nand UO_621 (O_621,N_19885,N_19945);
nor UO_622 (O_622,N_18378,N_18367);
or UO_623 (O_623,N_19741,N_19118);
or UO_624 (O_624,N_18391,N_18826);
nand UO_625 (O_625,N_18811,N_19629);
nand UO_626 (O_626,N_19353,N_18409);
xnor UO_627 (O_627,N_18402,N_18427);
xnor UO_628 (O_628,N_18708,N_18634);
xnor UO_629 (O_629,N_19925,N_18057);
or UO_630 (O_630,N_19635,N_19178);
xor UO_631 (O_631,N_19044,N_19324);
and UO_632 (O_632,N_19863,N_19558);
nand UO_633 (O_633,N_19964,N_19284);
or UO_634 (O_634,N_19328,N_18889);
and UO_635 (O_635,N_18004,N_18204);
and UO_636 (O_636,N_19199,N_18902);
or UO_637 (O_637,N_18069,N_18713);
xnor UO_638 (O_638,N_19393,N_19519);
nor UO_639 (O_639,N_19959,N_19229);
and UO_640 (O_640,N_19802,N_19266);
xnor UO_641 (O_641,N_18142,N_18558);
nor UO_642 (O_642,N_19588,N_18658);
xnor UO_643 (O_643,N_18830,N_19211);
nand UO_644 (O_644,N_19243,N_18556);
xor UO_645 (O_645,N_18288,N_18263);
xnor UO_646 (O_646,N_18967,N_18981);
xor UO_647 (O_647,N_18054,N_19366);
and UO_648 (O_648,N_18270,N_18973);
and UO_649 (O_649,N_18728,N_18748);
and UO_650 (O_650,N_18347,N_19372);
nand UO_651 (O_651,N_19179,N_18535);
or UO_652 (O_652,N_19673,N_19275);
or UO_653 (O_653,N_19219,N_18763);
nor UO_654 (O_654,N_18047,N_19956);
or UO_655 (O_655,N_19020,N_18597);
and UO_656 (O_656,N_19663,N_19617);
or UO_657 (O_657,N_19186,N_18450);
nand UO_658 (O_658,N_19033,N_19347);
nand UO_659 (O_659,N_19580,N_19407);
xnor UO_660 (O_660,N_18376,N_19903);
and UO_661 (O_661,N_18174,N_18948);
nand UO_662 (O_662,N_18691,N_19750);
or UO_663 (O_663,N_19533,N_19719);
xor UO_664 (O_664,N_19001,N_18858);
or UO_665 (O_665,N_18010,N_19652);
nor UO_666 (O_666,N_18127,N_19542);
xor UO_667 (O_667,N_19924,N_18322);
or UO_668 (O_668,N_19528,N_18881);
nor UO_669 (O_669,N_18979,N_18016);
xor UO_670 (O_670,N_18684,N_19770);
nor UO_671 (O_671,N_19297,N_18884);
or UO_672 (O_672,N_19338,N_19484);
nand UO_673 (O_673,N_18430,N_18628);
and UO_674 (O_674,N_19319,N_19414);
or UO_675 (O_675,N_19220,N_18017);
and UO_676 (O_676,N_19848,N_19509);
nand UO_677 (O_677,N_19833,N_19561);
nor UO_678 (O_678,N_18211,N_18977);
xnor UO_679 (O_679,N_19486,N_19563);
nor UO_680 (O_680,N_18927,N_19166);
nor UO_681 (O_681,N_18180,N_19962);
and UO_682 (O_682,N_19021,N_19030);
nor UO_683 (O_683,N_19241,N_19458);
and UO_684 (O_684,N_18852,N_18119);
nand UO_685 (O_685,N_18685,N_19994);
nand UO_686 (O_686,N_19080,N_18474);
or UO_687 (O_687,N_18539,N_18580);
nor UO_688 (O_688,N_19841,N_19337);
nor UO_689 (O_689,N_19875,N_19215);
and UO_690 (O_690,N_19566,N_18762);
xor UO_691 (O_691,N_18400,N_19096);
xnor UO_692 (O_692,N_19403,N_19592);
or UO_693 (O_693,N_19225,N_18930);
xor UO_694 (O_694,N_19304,N_19589);
nand UO_695 (O_695,N_19897,N_19007);
or UO_696 (O_696,N_19320,N_18095);
and UO_697 (O_697,N_18680,N_18679);
nand UO_698 (O_698,N_18612,N_19388);
nor UO_699 (O_699,N_18417,N_18421);
nand UO_700 (O_700,N_19439,N_19779);
nand UO_701 (O_701,N_18489,N_19686);
and UO_702 (O_702,N_18201,N_19213);
or UO_703 (O_703,N_19739,N_19271);
or UO_704 (O_704,N_19920,N_19792);
or UO_705 (O_705,N_19692,N_19691);
xnor UO_706 (O_706,N_18766,N_18064);
and UO_707 (O_707,N_18195,N_19627);
or UO_708 (O_708,N_18323,N_19065);
or UO_709 (O_709,N_19847,N_19099);
xnor UO_710 (O_710,N_19809,N_19870);
nand UO_711 (O_711,N_19740,N_18444);
xor UO_712 (O_712,N_19198,N_19054);
and UO_713 (O_713,N_19571,N_18572);
xnor UO_714 (O_714,N_19502,N_18707);
nand UO_715 (O_715,N_18873,N_19339);
nand UO_716 (O_716,N_19698,N_19075);
nor UO_717 (O_717,N_18405,N_18745);
nor UO_718 (O_718,N_18965,N_18364);
and UO_719 (O_719,N_19609,N_18063);
xor UO_720 (O_720,N_18667,N_19612);
nand UO_721 (O_721,N_19164,N_19757);
or UO_722 (O_722,N_19869,N_18414);
nor UO_723 (O_723,N_18570,N_19092);
and UO_724 (O_724,N_19532,N_19946);
xnor UO_725 (O_725,N_19953,N_19849);
and UO_726 (O_726,N_19272,N_18547);
nor UO_727 (O_727,N_18161,N_19459);
nand UO_728 (O_728,N_19369,N_18553);
and UO_729 (O_729,N_18653,N_19039);
or UO_730 (O_730,N_18756,N_19669);
nand UO_731 (O_731,N_19941,N_19646);
and UO_732 (O_732,N_18390,N_19027);
xnor UO_733 (O_733,N_18720,N_19214);
or UO_734 (O_734,N_18236,N_18032);
nor UO_735 (O_735,N_19772,N_19585);
and UO_736 (O_736,N_19727,N_18665);
or UO_737 (O_737,N_18931,N_18914);
xnor UO_738 (O_738,N_19307,N_18173);
nand UO_739 (O_739,N_18058,N_19290);
or UO_740 (O_740,N_19783,N_19763);
and UO_741 (O_741,N_19102,N_18654);
xor UO_742 (O_742,N_18452,N_19221);
nand UO_743 (O_743,N_19377,N_18899);
nand UO_744 (O_744,N_19536,N_18559);
nor UO_745 (O_745,N_18602,N_19814);
nand UO_746 (O_746,N_19672,N_19929);
xnor UO_747 (O_747,N_19680,N_18500);
or UO_748 (O_748,N_19768,N_18306);
and UO_749 (O_749,N_18503,N_18449);
xnor UO_750 (O_750,N_18012,N_18944);
nor UO_751 (O_751,N_18049,N_19446);
nor UO_752 (O_752,N_19707,N_18144);
nand UO_753 (O_753,N_18946,N_18831);
xor UO_754 (O_754,N_19607,N_19120);
or UO_755 (O_755,N_19838,N_19748);
and UO_756 (O_756,N_18608,N_18104);
nor UO_757 (O_757,N_18090,N_19922);
and UO_758 (O_758,N_18824,N_19273);
and UO_759 (O_759,N_19771,N_19639);
and UO_760 (O_760,N_19597,N_19285);
xnor UO_761 (O_761,N_18940,N_18578);
nand UO_762 (O_762,N_19648,N_18753);
nor UO_763 (O_763,N_19966,N_19026);
nor UO_764 (O_764,N_19825,N_18573);
or UO_765 (O_765,N_18415,N_19218);
and UO_766 (O_766,N_19010,N_19801);
nor UO_767 (O_767,N_18130,N_18723);
or UO_768 (O_768,N_19522,N_19697);
nand UO_769 (O_769,N_18978,N_18668);
xor UO_770 (O_770,N_18928,N_18737);
nand UO_771 (O_771,N_19795,N_19943);
and UO_772 (O_772,N_18110,N_18921);
nand UO_773 (O_773,N_18488,N_19674);
nor UO_774 (O_774,N_18311,N_18441);
and UO_775 (O_775,N_19160,N_19937);
and UO_776 (O_776,N_18416,N_18678);
and UO_777 (O_777,N_18460,N_19781);
and UO_778 (O_778,N_19776,N_18140);
xnor UO_779 (O_779,N_18792,N_18442);
and UO_780 (O_780,N_19485,N_18335);
nand UO_781 (O_781,N_19188,N_18507);
nand UO_782 (O_782,N_19371,N_18945);
nor UO_783 (O_783,N_19899,N_19891);
or UO_784 (O_784,N_18724,N_19183);
or UO_785 (O_785,N_19989,N_18044);
nor UO_786 (O_786,N_19513,N_19315);
nand UO_787 (O_787,N_19510,N_19386);
nor UO_788 (O_788,N_18975,N_19675);
xor UO_789 (O_789,N_18638,N_18115);
nand UO_790 (O_790,N_19264,N_19303);
xor UO_791 (O_791,N_19069,N_18273);
xnor UO_792 (O_792,N_18785,N_19579);
nor UO_793 (O_793,N_18803,N_19626);
and UO_794 (O_794,N_19846,N_19756);
and UO_795 (O_795,N_18867,N_19084);
or UO_796 (O_796,N_18128,N_19913);
nand UO_797 (O_797,N_18518,N_19464);
and UO_798 (O_798,N_18552,N_19912);
xor UO_799 (O_799,N_19056,N_19115);
or UO_800 (O_800,N_18789,N_18459);
or UO_801 (O_801,N_19122,N_19161);
nor UO_802 (O_802,N_19481,N_19541);
nor UO_803 (O_803,N_18014,N_18193);
nand UO_804 (O_804,N_18845,N_19175);
nand UO_805 (O_805,N_18467,N_18285);
nand UO_806 (O_806,N_19141,N_18439);
nor UO_807 (O_807,N_19939,N_18828);
nand UO_808 (O_808,N_18248,N_18837);
and UO_809 (O_809,N_19159,N_18007);
or UO_810 (O_810,N_18404,N_18809);
nand UO_811 (O_811,N_19432,N_18305);
or UO_812 (O_812,N_18609,N_18536);
xnor UO_813 (O_813,N_18876,N_19228);
and UO_814 (O_814,N_19095,N_19104);
or UO_815 (O_815,N_18692,N_19800);
or UO_816 (O_816,N_19767,N_19364);
nand UO_817 (O_817,N_18576,N_19276);
xor UO_818 (O_818,N_18100,N_19975);
nand UO_819 (O_819,N_19647,N_19676);
nand UO_820 (O_820,N_19911,N_19620);
nor UO_821 (O_821,N_18619,N_18036);
nor UO_822 (O_822,N_19958,N_19133);
nor UO_823 (O_823,N_18615,N_19984);
and UO_824 (O_824,N_19493,N_19977);
xnor UO_825 (O_825,N_19085,N_19785);
xor UO_826 (O_826,N_19684,N_18086);
nand UO_827 (O_827,N_19724,N_19878);
nor UO_828 (O_828,N_18222,N_18661);
or UO_829 (O_829,N_18833,N_18432);
or UO_830 (O_830,N_19236,N_18369);
xor UO_831 (O_831,N_19963,N_18361);
xor UO_832 (O_832,N_18179,N_18084);
nand UO_833 (O_833,N_18795,N_19794);
nand UO_834 (O_834,N_18543,N_18540);
nor UO_835 (O_835,N_18332,N_18062);
and UO_836 (O_836,N_19874,N_19168);
and UO_837 (O_837,N_18521,N_18583);
nand UO_838 (O_838,N_19172,N_19827);
xor UO_839 (O_839,N_19837,N_19346);
xnor UO_840 (O_840,N_18735,N_19619);
xnor UO_841 (O_841,N_18265,N_18244);
xnor UO_842 (O_842,N_19819,N_18381);
xor UO_843 (O_843,N_19088,N_19721);
nor UO_844 (O_844,N_18160,N_19553);
nand UO_845 (O_845,N_19492,N_18184);
nand UO_846 (O_846,N_18525,N_19896);
nor UO_847 (O_847,N_19286,N_18178);
xnor UO_848 (O_848,N_19259,N_18272);
xnor UO_849 (O_849,N_19655,N_19664);
and UO_850 (O_850,N_19850,N_19317);
xor UO_851 (O_851,N_18395,N_18482);
nor UO_852 (O_852,N_18336,N_19668);
nor UO_853 (O_853,N_18099,N_19644);
xnor UO_854 (O_854,N_19107,N_19818);
and UO_855 (O_855,N_19336,N_19712);
nor UO_856 (O_856,N_19149,N_18909);
and UO_857 (O_857,N_19256,N_19316);
nor UO_858 (O_858,N_18520,N_19582);
nand UO_859 (O_859,N_18096,N_19926);
and UO_860 (O_860,N_18021,N_18448);
nor UO_861 (O_861,N_18857,N_18139);
and UO_862 (O_862,N_18626,N_18933);
xor UO_863 (O_863,N_18509,N_19525);
nor UO_864 (O_864,N_18976,N_19032);
nor UO_865 (O_865,N_18646,N_18398);
xnor UO_866 (O_866,N_18912,N_18622);
and UO_867 (O_867,N_19699,N_19438);
nor UO_868 (O_868,N_18056,N_18741);
nand UO_869 (O_869,N_18823,N_18760);
xnor UO_870 (O_870,N_19066,N_18642);
nor UO_871 (O_871,N_19441,N_19300);
and UO_872 (O_872,N_19058,N_18585);
or UO_873 (O_873,N_18968,N_19539);
and UO_874 (O_874,N_19991,N_18532);
or UO_875 (O_875,N_18878,N_18986);
and UO_876 (O_876,N_19349,N_18687);
xor UO_877 (O_877,N_19494,N_18670);
or UO_878 (O_878,N_18469,N_18162);
nor UO_879 (O_879,N_18375,N_18952);
and UO_880 (O_880,N_18334,N_18024);
nand UO_881 (O_881,N_19932,N_19024);
and UO_882 (O_882,N_18582,N_19413);
nand UO_883 (O_883,N_18875,N_19279);
nand UO_884 (O_884,N_19362,N_18701);
xor UO_885 (O_885,N_19378,N_18925);
nor UO_886 (O_886,N_19134,N_18254);
nand UO_887 (O_887,N_19516,N_19957);
nor UO_888 (O_888,N_18362,N_19515);
and UO_889 (O_889,N_19948,N_18549);
xor UO_890 (O_890,N_18437,N_19973);
nor UO_891 (O_891,N_18700,N_18112);
nand UO_892 (O_892,N_18587,N_18294);
xor UO_893 (O_893,N_19429,N_19394);
or UO_894 (O_894,N_18712,N_19694);
or UO_895 (O_895,N_18468,N_19165);
and UO_896 (O_896,N_19754,N_19905);
xor UO_897 (O_897,N_19969,N_19332);
nand UO_898 (O_898,N_18716,N_19047);
xor UO_899 (O_899,N_18456,N_19666);
and UO_900 (O_900,N_19907,N_18413);
and UO_901 (O_901,N_18333,N_18351);
and UO_902 (O_902,N_18768,N_19978);
and UO_903 (O_903,N_18633,N_19761);
xnor UO_904 (O_904,N_18251,N_19573);
and UO_905 (O_905,N_19430,N_18120);
and UO_906 (O_906,N_19535,N_19463);
xor UO_907 (O_907,N_18637,N_18964);
xnor UO_908 (O_908,N_18907,N_18676);
xor UO_909 (O_909,N_18499,N_19881);
and UO_910 (O_910,N_18129,N_19457);
nand UO_911 (O_911,N_19685,N_19174);
or UO_912 (O_912,N_19467,N_18117);
nand UO_913 (O_913,N_19262,N_18045);
and UO_914 (O_914,N_19606,N_18926);
or UO_915 (O_915,N_18262,N_19013);
or UO_916 (O_916,N_18537,N_19341);
and UO_917 (O_917,N_18893,N_19356);
xor UO_918 (O_918,N_19295,N_18041);
or UO_919 (O_919,N_19034,N_19059);
or UO_920 (O_920,N_18234,N_18353);
nor UO_921 (O_921,N_18861,N_18342);
xor UO_922 (O_922,N_18674,N_19701);
nor UO_923 (O_923,N_19097,N_18419);
or UO_924 (O_924,N_19496,N_19660);
nand UO_925 (O_925,N_19375,N_18424);
or UO_926 (O_926,N_19524,N_18487);
and UO_927 (O_927,N_18969,N_18802);
nor UO_928 (O_928,N_19181,N_19110);
or UO_929 (O_929,N_19268,N_18801);
and UO_930 (O_930,N_18501,N_18631);
and UO_931 (O_931,N_18475,N_18686);
nand UO_932 (O_932,N_18197,N_19917);
xnor UO_933 (O_933,N_18034,N_18644);
nor UO_934 (O_934,N_19466,N_18799);
and UO_935 (O_935,N_19344,N_19130);
nor UO_936 (O_936,N_18258,N_18936);
and UO_937 (O_937,N_18463,N_18087);
or UO_938 (O_938,N_18954,N_18005);
and UO_939 (O_939,N_19506,N_18841);
and UO_940 (O_940,N_19921,N_18387);
nor UO_941 (O_941,N_18412,N_18616);
nand UO_942 (O_942,N_18887,N_19412);
xnor UO_943 (O_943,N_19565,N_19895);
nor UO_944 (O_944,N_19879,N_19143);
and UO_945 (O_945,N_19405,N_19512);
and UO_946 (O_946,N_18784,N_19322);
and UO_947 (O_947,N_18279,N_19016);
or UO_948 (O_948,N_19135,N_18476);
nor UO_949 (O_949,N_18203,N_19245);
and UO_950 (O_950,N_18123,N_19876);
xnor UO_951 (O_951,N_18393,N_18061);
nor UO_952 (O_952,N_19469,N_18780);
nor UO_953 (O_953,N_19746,N_19293);
or UO_954 (O_954,N_19974,N_18384);
nor UO_955 (O_955,N_19642,N_18951);
or UO_956 (O_956,N_19081,N_19659);
and UO_957 (O_957,N_18955,N_18777);
and UO_958 (O_958,N_18868,N_19747);
and UO_959 (O_959,N_19578,N_19952);
nand UO_960 (O_960,N_18702,N_18650);
and UO_961 (O_961,N_19599,N_18810);
nor UO_962 (O_962,N_19799,N_19329);
xnor UO_963 (O_963,N_18302,N_19769);
nand UO_964 (O_964,N_19009,N_18776);
or UO_965 (O_965,N_19749,N_19006);
or UO_966 (O_966,N_19696,N_18960);
and UO_967 (O_967,N_19773,N_18043);
nor UO_968 (O_968,N_18013,N_18209);
xor UO_969 (O_969,N_18786,N_18382);
nand UO_970 (O_970,N_18577,N_19240);
and UO_971 (O_971,N_19575,N_18994);
or UO_972 (O_972,N_18749,N_18172);
nand UO_973 (O_973,N_19035,N_19931);
or UO_974 (O_974,N_19786,N_19670);
or UO_975 (O_975,N_19734,N_18379);
or UO_976 (O_976,N_19253,N_18231);
xor UO_977 (O_977,N_19476,N_19947);
nand UO_978 (O_978,N_19504,N_19173);
nor UO_979 (O_979,N_18651,N_18742);
and UO_980 (O_980,N_18929,N_18124);
and UO_981 (O_981,N_18281,N_18226);
or UO_982 (O_982,N_18730,N_18561);
nand UO_983 (O_983,N_18999,N_19121);
nand UO_984 (O_984,N_18607,N_19151);
and UO_985 (O_985,N_18513,N_19468);
nor UO_986 (O_986,N_18106,N_19381);
nand UO_987 (O_987,N_19090,N_19889);
nor UO_988 (O_988,N_18483,N_19793);
xor UO_989 (O_989,N_18163,N_18560);
nand UO_990 (O_990,N_18436,N_19593);
or UO_991 (O_991,N_18228,N_18494);
xor UO_992 (O_992,N_18662,N_19742);
or UO_993 (O_993,N_19232,N_18657);
and UO_994 (O_994,N_19645,N_19762);
or UO_995 (O_995,N_19406,N_18292);
nand UO_996 (O_996,N_18392,N_18418);
xnor UO_997 (O_997,N_19919,N_19396);
xnor UO_998 (O_998,N_19004,N_19968);
nand UO_999 (O_999,N_19567,N_19544);
and UO_1000 (O_1000,N_19769,N_18739);
or UO_1001 (O_1001,N_18669,N_19016);
xnor UO_1002 (O_1002,N_18785,N_19672);
xnor UO_1003 (O_1003,N_19333,N_19038);
nand UO_1004 (O_1004,N_18021,N_19786);
nand UO_1005 (O_1005,N_18103,N_19190);
nor UO_1006 (O_1006,N_18545,N_19451);
xor UO_1007 (O_1007,N_19481,N_19759);
nand UO_1008 (O_1008,N_19226,N_19954);
or UO_1009 (O_1009,N_18783,N_18018);
nor UO_1010 (O_1010,N_18205,N_18406);
nor UO_1011 (O_1011,N_19981,N_19772);
nand UO_1012 (O_1012,N_19161,N_18640);
nor UO_1013 (O_1013,N_18540,N_18027);
and UO_1014 (O_1014,N_19803,N_18131);
xnor UO_1015 (O_1015,N_18122,N_19801);
nor UO_1016 (O_1016,N_19431,N_18315);
and UO_1017 (O_1017,N_19092,N_19691);
or UO_1018 (O_1018,N_19068,N_19864);
and UO_1019 (O_1019,N_18657,N_19827);
nand UO_1020 (O_1020,N_18406,N_19037);
xor UO_1021 (O_1021,N_18597,N_18240);
and UO_1022 (O_1022,N_18472,N_19556);
nor UO_1023 (O_1023,N_18671,N_18691);
nand UO_1024 (O_1024,N_19262,N_19038);
or UO_1025 (O_1025,N_18608,N_18473);
nand UO_1026 (O_1026,N_19143,N_19162);
and UO_1027 (O_1027,N_18978,N_18580);
and UO_1028 (O_1028,N_19286,N_18823);
xnor UO_1029 (O_1029,N_18086,N_19770);
xnor UO_1030 (O_1030,N_18258,N_19467);
nand UO_1031 (O_1031,N_19982,N_19815);
nand UO_1032 (O_1032,N_19334,N_18350);
nor UO_1033 (O_1033,N_18043,N_19445);
nor UO_1034 (O_1034,N_19081,N_18942);
and UO_1035 (O_1035,N_18949,N_19971);
nor UO_1036 (O_1036,N_18712,N_18231);
nor UO_1037 (O_1037,N_18851,N_18015);
nor UO_1038 (O_1038,N_18024,N_19936);
nor UO_1039 (O_1039,N_19021,N_18900);
nand UO_1040 (O_1040,N_18180,N_18359);
or UO_1041 (O_1041,N_19086,N_19034);
nand UO_1042 (O_1042,N_19479,N_19826);
or UO_1043 (O_1043,N_19045,N_18637);
and UO_1044 (O_1044,N_19832,N_19304);
nor UO_1045 (O_1045,N_18828,N_18930);
nor UO_1046 (O_1046,N_18702,N_18112);
and UO_1047 (O_1047,N_18496,N_18931);
nor UO_1048 (O_1048,N_19145,N_19104);
or UO_1049 (O_1049,N_19054,N_19191);
and UO_1050 (O_1050,N_19326,N_18188);
and UO_1051 (O_1051,N_18625,N_19360);
or UO_1052 (O_1052,N_19068,N_19239);
or UO_1053 (O_1053,N_18657,N_19944);
and UO_1054 (O_1054,N_18977,N_19906);
or UO_1055 (O_1055,N_19263,N_18532);
nor UO_1056 (O_1056,N_18655,N_19521);
nand UO_1057 (O_1057,N_19559,N_18247);
and UO_1058 (O_1058,N_19669,N_19399);
and UO_1059 (O_1059,N_19387,N_18776);
nand UO_1060 (O_1060,N_18668,N_18349);
and UO_1061 (O_1061,N_18442,N_19435);
nand UO_1062 (O_1062,N_18192,N_18072);
xnor UO_1063 (O_1063,N_18808,N_19550);
nor UO_1064 (O_1064,N_19414,N_18603);
nand UO_1065 (O_1065,N_18685,N_18995);
xnor UO_1066 (O_1066,N_19680,N_19506);
and UO_1067 (O_1067,N_18418,N_19716);
or UO_1068 (O_1068,N_19145,N_18543);
nand UO_1069 (O_1069,N_18266,N_19382);
nand UO_1070 (O_1070,N_19299,N_19741);
nor UO_1071 (O_1071,N_19197,N_19517);
nand UO_1072 (O_1072,N_18831,N_19111);
or UO_1073 (O_1073,N_18392,N_19889);
or UO_1074 (O_1074,N_18611,N_18227);
xnor UO_1075 (O_1075,N_18011,N_18813);
and UO_1076 (O_1076,N_19171,N_19918);
nand UO_1077 (O_1077,N_19068,N_18934);
xnor UO_1078 (O_1078,N_18143,N_19031);
and UO_1079 (O_1079,N_19605,N_18025);
or UO_1080 (O_1080,N_19231,N_18625);
xnor UO_1081 (O_1081,N_18734,N_19123);
or UO_1082 (O_1082,N_18269,N_18191);
or UO_1083 (O_1083,N_19009,N_18463);
and UO_1084 (O_1084,N_18450,N_18155);
and UO_1085 (O_1085,N_19084,N_18923);
or UO_1086 (O_1086,N_19500,N_18207);
nor UO_1087 (O_1087,N_19467,N_18975);
and UO_1088 (O_1088,N_19388,N_18850);
xor UO_1089 (O_1089,N_18261,N_18651);
nor UO_1090 (O_1090,N_18956,N_18676);
or UO_1091 (O_1091,N_19558,N_19644);
nand UO_1092 (O_1092,N_19683,N_19596);
and UO_1093 (O_1093,N_18074,N_19085);
nor UO_1094 (O_1094,N_19374,N_19528);
xor UO_1095 (O_1095,N_18781,N_18458);
nor UO_1096 (O_1096,N_19166,N_19046);
nand UO_1097 (O_1097,N_19360,N_18863);
nor UO_1098 (O_1098,N_18074,N_18457);
xnor UO_1099 (O_1099,N_19343,N_18206);
nor UO_1100 (O_1100,N_18317,N_18627);
nand UO_1101 (O_1101,N_19589,N_18250);
nand UO_1102 (O_1102,N_18213,N_19236);
xnor UO_1103 (O_1103,N_18385,N_19053);
or UO_1104 (O_1104,N_18657,N_18851);
or UO_1105 (O_1105,N_18878,N_18893);
xnor UO_1106 (O_1106,N_18106,N_19832);
and UO_1107 (O_1107,N_18884,N_18238);
xnor UO_1108 (O_1108,N_19298,N_19697);
nor UO_1109 (O_1109,N_19022,N_19883);
and UO_1110 (O_1110,N_19722,N_18278);
or UO_1111 (O_1111,N_19564,N_19975);
nand UO_1112 (O_1112,N_18679,N_18616);
xor UO_1113 (O_1113,N_18511,N_18791);
nor UO_1114 (O_1114,N_18073,N_18174);
xor UO_1115 (O_1115,N_18072,N_18915);
and UO_1116 (O_1116,N_18076,N_18337);
and UO_1117 (O_1117,N_19253,N_19430);
nor UO_1118 (O_1118,N_18693,N_18042);
and UO_1119 (O_1119,N_19713,N_18442);
and UO_1120 (O_1120,N_18385,N_18204);
nand UO_1121 (O_1121,N_18128,N_18154);
xor UO_1122 (O_1122,N_19953,N_18591);
or UO_1123 (O_1123,N_18772,N_18822);
nor UO_1124 (O_1124,N_18103,N_18617);
nor UO_1125 (O_1125,N_18290,N_18779);
nand UO_1126 (O_1126,N_18174,N_18129);
and UO_1127 (O_1127,N_19963,N_18822);
xnor UO_1128 (O_1128,N_19921,N_18385);
xor UO_1129 (O_1129,N_18063,N_19614);
xnor UO_1130 (O_1130,N_18125,N_18420);
nor UO_1131 (O_1131,N_18448,N_18275);
and UO_1132 (O_1132,N_19372,N_18097);
nor UO_1133 (O_1133,N_19985,N_18307);
and UO_1134 (O_1134,N_18232,N_19086);
or UO_1135 (O_1135,N_19004,N_19428);
xnor UO_1136 (O_1136,N_19482,N_19631);
or UO_1137 (O_1137,N_19456,N_18807);
xor UO_1138 (O_1138,N_18975,N_19482);
or UO_1139 (O_1139,N_19638,N_19061);
nand UO_1140 (O_1140,N_19586,N_18303);
xor UO_1141 (O_1141,N_19440,N_19945);
and UO_1142 (O_1142,N_18911,N_18295);
and UO_1143 (O_1143,N_18233,N_18347);
nor UO_1144 (O_1144,N_18164,N_19472);
xnor UO_1145 (O_1145,N_19898,N_19707);
or UO_1146 (O_1146,N_19443,N_19864);
or UO_1147 (O_1147,N_19085,N_18019);
nor UO_1148 (O_1148,N_18449,N_18712);
and UO_1149 (O_1149,N_18445,N_18687);
and UO_1150 (O_1150,N_18861,N_18437);
or UO_1151 (O_1151,N_18795,N_19284);
xor UO_1152 (O_1152,N_18101,N_18515);
nor UO_1153 (O_1153,N_18213,N_19132);
xnor UO_1154 (O_1154,N_19427,N_19748);
xor UO_1155 (O_1155,N_19355,N_19842);
or UO_1156 (O_1156,N_18248,N_19014);
nand UO_1157 (O_1157,N_18049,N_19489);
and UO_1158 (O_1158,N_19878,N_19222);
or UO_1159 (O_1159,N_18017,N_18297);
nor UO_1160 (O_1160,N_19601,N_19317);
or UO_1161 (O_1161,N_19845,N_19079);
or UO_1162 (O_1162,N_19904,N_19477);
nand UO_1163 (O_1163,N_19844,N_18677);
xnor UO_1164 (O_1164,N_18195,N_19897);
xnor UO_1165 (O_1165,N_19838,N_18191);
nand UO_1166 (O_1166,N_18269,N_19544);
nand UO_1167 (O_1167,N_19200,N_18109);
and UO_1168 (O_1168,N_19063,N_18473);
nand UO_1169 (O_1169,N_18692,N_19751);
nor UO_1170 (O_1170,N_18854,N_19066);
xnor UO_1171 (O_1171,N_19869,N_18251);
xor UO_1172 (O_1172,N_18722,N_19457);
and UO_1173 (O_1173,N_18958,N_18831);
and UO_1174 (O_1174,N_18186,N_19458);
or UO_1175 (O_1175,N_18138,N_19162);
nor UO_1176 (O_1176,N_19179,N_18548);
or UO_1177 (O_1177,N_18841,N_18176);
nand UO_1178 (O_1178,N_18080,N_19228);
nand UO_1179 (O_1179,N_18114,N_18677);
nor UO_1180 (O_1180,N_18203,N_18317);
xnor UO_1181 (O_1181,N_18411,N_18217);
nand UO_1182 (O_1182,N_18710,N_18171);
nor UO_1183 (O_1183,N_19957,N_19724);
nor UO_1184 (O_1184,N_18310,N_19125);
or UO_1185 (O_1185,N_18278,N_18826);
nor UO_1186 (O_1186,N_18919,N_19910);
and UO_1187 (O_1187,N_18816,N_18215);
xor UO_1188 (O_1188,N_18916,N_18637);
and UO_1189 (O_1189,N_19985,N_18539);
xnor UO_1190 (O_1190,N_18891,N_18574);
nand UO_1191 (O_1191,N_18928,N_18337);
nand UO_1192 (O_1192,N_19741,N_18900);
or UO_1193 (O_1193,N_19290,N_18312);
nand UO_1194 (O_1194,N_19515,N_19353);
nand UO_1195 (O_1195,N_18363,N_19748);
or UO_1196 (O_1196,N_19771,N_18730);
or UO_1197 (O_1197,N_19734,N_18242);
or UO_1198 (O_1198,N_18559,N_19596);
and UO_1199 (O_1199,N_18120,N_19811);
and UO_1200 (O_1200,N_18913,N_19260);
nand UO_1201 (O_1201,N_18298,N_19000);
nor UO_1202 (O_1202,N_19029,N_19301);
or UO_1203 (O_1203,N_18452,N_19501);
or UO_1204 (O_1204,N_19910,N_18035);
or UO_1205 (O_1205,N_18172,N_19966);
or UO_1206 (O_1206,N_18416,N_19736);
and UO_1207 (O_1207,N_18368,N_19774);
xor UO_1208 (O_1208,N_19942,N_19177);
and UO_1209 (O_1209,N_18942,N_19139);
and UO_1210 (O_1210,N_19927,N_19320);
or UO_1211 (O_1211,N_18970,N_18165);
nor UO_1212 (O_1212,N_19124,N_18161);
and UO_1213 (O_1213,N_19552,N_18014);
nor UO_1214 (O_1214,N_19722,N_19310);
nor UO_1215 (O_1215,N_19914,N_18483);
or UO_1216 (O_1216,N_19638,N_18657);
nand UO_1217 (O_1217,N_19725,N_18216);
and UO_1218 (O_1218,N_18451,N_19042);
or UO_1219 (O_1219,N_19831,N_18355);
nor UO_1220 (O_1220,N_19940,N_19182);
or UO_1221 (O_1221,N_18901,N_19909);
or UO_1222 (O_1222,N_19750,N_19988);
xor UO_1223 (O_1223,N_18007,N_19039);
or UO_1224 (O_1224,N_19992,N_18421);
nand UO_1225 (O_1225,N_18578,N_19369);
nor UO_1226 (O_1226,N_19451,N_19812);
nor UO_1227 (O_1227,N_18050,N_19549);
xor UO_1228 (O_1228,N_19012,N_18724);
nand UO_1229 (O_1229,N_18907,N_18115);
or UO_1230 (O_1230,N_18544,N_18934);
nor UO_1231 (O_1231,N_18443,N_18733);
nand UO_1232 (O_1232,N_18039,N_19195);
nor UO_1233 (O_1233,N_18937,N_19556);
xor UO_1234 (O_1234,N_18844,N_18338);
xor UO_1235 (O_1235,N_18649,N_19533);
nand UO_1236 (O_1236,N_18276,N_18018);
or UO_1237 (O_1237,N_18940,N_19509);
nor UO_1238 (O_1238,N_19721,N_19702);
xnor UO_1239 (O_1239,N_19800,N_18917);
or UO_1240 (O_1240,N_19665,N_18879);
or UO_1241 (O_1241,N_19183,N_19692);
xor UO_1242 (O_1242,N_18176,N_18007);
nor UO_1243 (O_1243,N_19430,N_19674);
and UO_1244 (O_1244,N_18943,N_19902);
xor UO_1245 (O_1245,N_18558,N_18186);
nand UO_1246 (O_1246,N_18675,N_18964);
and UO_1247 (O_1247,N_18656,N_19048);
nand UO_1248 (O_1248,N_19505,N_18528);
or UO_1249 (O_1249,N_18152,N_19867);
nand UO_1250 (O_1250,N_19328,N_19146);
xor UO_1251 (O_1251,N_18773,N_19014);
nand UO_1252 (O_1252,N_18987,N_19839);
nor UO_1253 (O_1253,N_18843,N_19116);
or UO_1254 (O_1254,N_19284,N_18444);
nand UO_1255 (O_1255,N_18616,N_18411);
nor UO_1256 (O_1256,N_19791,N_18020);
xnor UO_1257 (O_1257,N_18929,N_19619);
xnor UO_1258 (O_1258,N_19245,N_18184);
and UO_1259 (O_1259,N_19374,N_18634);
xor UO_1260 (O_1260,N_19041,N_19381);
xnor UO_1261 (O_1261,N_19260,N_19006);
xor UO_1262 (O_1262,N_18634,N_19476);
nand UO_1263 (O_1263,N_19605,N_18411);
xor UO_1264 (O_1264,N_18401,N_19891);
xnor UO_1265 (O_1265,N_19049,N_19411);
or UO_1266 (O_1266,N_18199,N_18329);
nor UO_1267 (O_1267,N_19833,N_19381);
xor UO_1268 (O_1268,N_18439,N_19219);
and UO_1269 (O_1269,N_19957,N_19308);
nand UO_1270 (O_1270,N_19043,N_19391);
nor UO_1271 (O_1271,N_18266,N_18475);
nor UO_1272 (O_1272,N_19805,N_18686);
or UO_1273 (O_1273,N_18310,N_18671);
nor UO_1274 (O_1274,N_18229,N_19486);
nand UO_1275 (O_1275,N_18802,N_19724);
or UO_1276 (O_1276,N_19419,N_18389);
xor UO_1277 (O_1277,N_18541,N_18530);
or UO_1278 (O_1278,N_19604,N_18168);
or UO_1279 (O_1279,N_19420,N_19668);
and UO_1280 (O_1280,N_19403,N_18608);
xor UO_1281 (O_1281,N_18413,N_18793);
xnor UO_1282 (O_1282,N_18053,N_19768);
and UO_1283 (O_1283,N_19397,N_18010);
nand UO_1284 (O_1284,N_19646,N_18935);
nor UO_1285 (O_1285,N_19810,N_18503);
and UO_1286 (O_1286,N_19169,N_18041);
and UO_1287 (O_1287,N_18855,N_18258);
or UO_1288 (O_1288,N_19083,N_19398);
nor UO_1289 (O_1289,N_19270,N_18558);
or UO_1290 (O_1290,N_19162,N_18824);
nand UO_1291 (O_1291,N_19166,N_19590);
and UO_1292 (O_1292,N_19998,N_18320);
nor UO_1293 (O_1293,N_19343,N_19676);
and UO_1294 (O_1294,N_18522,N_19050);
and UO_1295 (O_1295,N_19368,N_19419);
or UO_1296 (O_1296,N_18541,N_18088);
xnor UO_1297 (O_1297,N_19143,N_18533);
and UO_1298 (O_1298,N_18483,N_18348);
or UO_1299 (O_1299,N_19565,N_19265);
or UO_1300 (O_1300,N_18122,N_19962);
and UO_1301 (O_1301,N_18488,N_19372);
xnor UO_1302 (O_1302,N_18552,N_18794);
nand UO_1303 (O_1303,N_18116,N_19564);
nor UO_1304 (O_1304,N_18022,N_18811);
nand UO_1305 (O_1305,N_19193,N_19133);
nand UO_1306 (O_1306,N_19271,N_19673);
xor UO_1307 (O_1307,N_18988,N_19738);
and UO_1308 (O_1308,N_18943,N_18981);
nor UO_1309 (O_1309,N_19159,N_18403);
nor UO_1310 (O_1310,N_18495,N_18712);
nor UO_1311 (O_1311,N_19975,N_18143);
or UO_1312 (O_1312,N_19813,N_19046);
xor UO_1313 (O_1313,N_19649,N_19612);
and UO_1314 (O_1314,N_19297,N_18740);
or UO_1315 (O_1315,N_18589,N_18323);
or UO_1316 (O_1316,N_18484,N_19507);
and UO_1317 (O_1317,N_18317,N_19733);
or UO_1318 (O_1318,N_18644,N_19115);
nor UO_1319 (O_1319,N_18034,N_18470);
nor UO_1320 (O_1320,N_18915,N_18687);
xor UO_1321 (O_1321,N_19654,N_19148);
and UO_1322 (O_1322,N_19011,N_18013);
or UO_1323 (O_1323,N_19618,N_18429);
and UO_1324 (O_1324,N_19379,N_18426);
or UO_1325 (O_1325,N_19358,N_18398);
and UO_1326 (O_1326,N_18611,N_19988);
or UO_1327 (O_1327,N_18635,N_18024);
and UO_1328 (O_1328,N_19553,N_18814);
and UO_1329 (O_1329,N_19953,N_18488);
and UO_1330 (O_1330,N_19124,N_18910);
nand UO_1331 (O_1331,N_18005,N_18948);
nand UO_1332 (O_1332,N_18262,N_18048);
nor UO_1333 (O_1333,N_18273,N_18219);
nor UO_1334 (O_1334,N_18944,N_18905);
and UO_1335 (O_1335,N_19319,N_18880);
or UO_1336 (O_1336,N_19292,N_18776);
and UO_1337 (O_1337,N_18291,N_18505);
and UO_1338 (O_1338,N_19810,N_19790);
nand UO_1339 (O_1339,N_19496,N_18411);
nor UO_1340 (O_1340,N_18335,N_18205);
xor UO_1341 (O_1341,N_19764,N_18118);
and UO_1342 (O_1342,N_18675,N_19296);
nor UO_1343 (O_1343,N_18907,N_18543);
nand UO_1344 (O_1344,N_19577,N_18905);
xnor UO_1345 (O_1345,N_18435,N_18957);
or UO_1346 (O_1346,N_18214,N_18611);
xnor UO_1347 (O_1347,N_19417,N_19908);
and UO_1348 (O_1348,N_18204,N_18132);
nand UO_1349 (O_1349,N_19151,N_19535);
nor UO_1350 (O_1350,N_19814,N_18307);
and UO_1351 (O_1351,N_19115,N_18757);
or UO_1352 (O_1352,N_19360,N_19461);
nor UO_1353 (O_1353,N_18093,N_19158);
or UO_1354 (O_1354,N_18597,N_19589);
or UO_1355 (O_1355,N_19221,N_19175);
and UO_1356 (O_1356,N_19687,N_18418);
nand UO_1357 (O_1357,N_18571,N_19589);
and UO_1358 (O_1358,N_19506,N_18378);
and UO_1359 (O_1359,N_19387,N_18657);
and UO_1360 (O_1360,N_18819,N_18323);
nand UO_1361 (O_1361,N_18001,N_18536);
or UO_1362 (O_1362,N_19776,N_18002);
nand UO_1363 (O_1363,N_19007,N_18561);
xnor UO_1364 (O_1364,N_19495,N_18684);
nor UO_1365 (O_1365,N_19440,N_19206);
nor UO_1366 (O_1366,N_19833,N_18935);
nand UO_1367 (O_1367,N_19325,N_18593);
xnor UO_1368 (O_1368,N_19308,N_19295);
and UO_1369 (O_1369,N_18771,N_19959);
and UO_1370 (O_1370,N_19411,N_18235);
xnor UO_1371 (O_1371,N_19930,N_19394);
nand UO_1372 (O_1372,N_18628,N_19118);
and UO_1373 (O_1373,N_19216,N_19137);
and UO_1374 (O_1374,N_19968,N_18865);
or UO_1375 (O_1375,N_19835,N_18116);
and UO_1376 (O_1376,N_18722,N_19132);
nand UO_1377 (O_1377,N_18653,N_18785);
and UO_1378 (O_1378,N_19174,N_19418);
and UO_1379 (O_1379,N_18035,N_18154);
nand UO_1380 (O_1380,N_18571,N_18926);
nand UO_1381 (O_1381,N_18991,N_19816);
xnor UO_1382 (O_1382,N_18434,N_19822);
xnor UO_1383 (O_1383,N_19735,N_18922);
nor UO_1384 (O_1384,N_19669,N_19704);
xnor UO_1385 (O_1385,N_19857,N_19185);
or UO_1386 (O_1386,N_18476,N_18641);
xnor UO_1387 (O_1387,N_19322,N_19394);
xnor UO_1388 (O_1388,N_18956,N_18284);
xor UO_1389 (O_1389,N_19986,N_19688);
xnor UO_1390 (O_1390,N_18729,N_19475);
nor UO_1391 (O_1391,N_18050,N_19591);
or UO_1392 (O_1392,N_18918,N_19752);
xor UO_1393 (O_1393,N_19763,N_18624);
xor UO_1394 (O_1394,N_19372,N_19417);
nand UO_1395 (O_1395,N_18758,N_18089);
or UO_1396 (O_1396,N_18520,N_19480);
nand UO_1397 (O_1397,N_18785,N_18602);
xnor UO_1398 (O_1398,N_19652,N_18267);
or UO_1399 (O_1399,N_19078,N_18733);
xor UO_1400 (O_1400,N_18182,N_19883);
xor UO_1401 (O_1401,N_19827,N_19807);
and UO_1402 (O_1402,N_18812,N_19043);
or UO_1403 (O_1403,N_18419,N_19162);
and UO_1404 (O_1404,N_19627,N_18417);
xor UO_1405 (O_1405,N_19031,N_19140);
nand UO_1406 (O_1406,N_18686,N_18029);
or UO_1407 (O_1407,N_19347,N_19756);
or UO_1408 (O_1408,N_19073,N_18972);
nand UO_1409 (O_1409,N_18390,N_18675);
nand UO_1410 (O_1410,N_18176,N_18498);
or UO_1411 (O_1411,N_19974,N_18723);
nor UO_1412 (O_1412,N_18172,N_19570);
and UO_1413 (O_1413,N_18336,N_19256);
or UO_1414 (O_1414,N_19710,N_19719);
xor UO_1415 (O_1415,N_19558,N_18274);
nor UO_1416 (O_1416,N_18176,N_19918);
and UO_1417 (O_1417,N_19242,N_18235);
or UO_1418 (O_1418,N_18960,N_18294);
or UO_1419 (O_1419,N_19727,N_19068);
or UO_1420 (O_1420,N_18954,N_18856);
xnor UO_1421 (O_1421,N_19989,N_18381);
nand UO_1422 (O_1422,N_19051,N_18717);
nor UO_1423 (O_1423,N_19169,N_19657);
or UO_1424 (O_1424,N_19701,N_19083);
or UO_1425 (O_1425,N_18322,N_19057);
nand UO_1426 (O_1426,N_18437,N_18600);
nand UO_1427 (O_1427,N_19450,N_18974);
nand UO_1428 (O_1428,N_19931,N_19767);
and UO_1429 (O_1429,N_19539,N_18116);
xor UO_1430 (O_1430,N_19991,N_18924);
and UO_1431 (O_1431,N_18248,N_19069);
nor UO_1432 (O_1432,N_18162,N_19080);
nand UO_1433 (O_1433,N_18434,N_19891);
nor UO_1434 (O_1434,N_19428,N_18310);
or UO_1435 (O_1435,N_19175,N_18626);
or UO_1436 (O_1436,N_19502,N_18090);
xor UO_1437 (O_1437,N_19693,N_19179);
or UO_1438 (O_1438,N_19984,N_19879);
and UO_1439 (O_1439,N_19075,N_19529);
nor UO_1440 (O_1440,N_19482,N_19818);
nor UO_1441 (O_1441,N_19885,N_18082);
or UO_1442 (O_1442,N_19668,N_18570);
nand UO_1443 (O_1443,N_18064,N_18835);
nand UO_1444 (O_1444,N_19630,N_18516);
or UO_1445 (O_1445,N_18657,N_19104);
xnor UO_1446 (O_1446,N_19924,N_18057);
xnor UO_1447 (O_1447,N_19332,N_18388);
xnor UO_1448 (O_1448,N_19643,N_18919);
or UO_1449 (O_1449,N_19723,N_18349);
or UO_1450 (O_1450,N_18529,N_18419);
or UO_1451 (O_1451,N_18275,N_19719);
nor UO_1452 (O_1452,N_19980,N_18486);
and UO_1453 (O_1453,N_19171,N_19184);
nor UO_1454 (O_1454,N_19664,N_18181);
nand UO_1455 (O_1455,N_19887,N_19743);
or UO_1456 (O_1456,N_19230,N_18772);
nor UO_1457 (O_1457,N_19324,N_18297);
nand UO_1458 (O_1458,N_18509,N_18984);
nand UO_1459 (O_1459,N_18170,N_18369);
and UO_1460 (O_1460,N_19233,N_18322);
nand UO_1461 (O_1461,N_18503,N_18678);
and UO_1462 (O_1462,N_18307,N_18489);
nor UO_1463 (O_1463,N_18722,N_19114);
nor UO_1464 (O_1464,N_18409,N_18750);
xor UO_1465 (O_1465,N_19805,N_18490);
and UO_1466 (O_1466,N_18467,N_19145);
xor UO_1467 (O_1467,N_18034,N_18025);
nor UO_1468 (O_1468,N_19398,N_18057);
and UO_1469 (O_1469,N_19821,N_19680);
and UO_1470 (O_1470,N_19090,N_19016);
nor UO_1471 (O_1471,N_19207,N_18808);
nand UO_1472 (O_1472,N_18057,N_19505);
and UO_1473 (O_1473,N_19873,N_18655);
nor UO_1474 (O_1474,N_19006,N_19897);
nor UO_1475 (O_1475,N_18254,N_19962);
or UO_1476 (O_1476,N_18190,N_18742);
and UO_1477 (O_1477,N_18465,N_19075);
nand UO_1478 (O_1478,N_19054,N_19845);
xnor UO_1479 (O_1479,N_18732,N_19731);
or UO_1480 (O_1480,N_19377,N_19028);
or UO_1481 (O_1481,N_19479,N_18786);
nand UO_1482 (O_1482,N_18598,N_19658);
or UO_1483 (O_1483,N_19791,N_19495);
nand UO_1484 (O_1484,N_19594,N_19764);
xor UO_1485 (O_1485,N_19979,N_18063);
xnor UO_1486 (O_1486,N_18273,N_19469);
nor UO_1487 (O_1487,N_18716,N_19762);
xnor UO_1488 (O_1488,N_18269,N_19188);
xnor UO_1489 (O_1489,N_18165,N_18418);
nand UO_1490 (O_1490,N_19730,N_19712);
xor UO_1491 (O_1491,N_18888,N_19265);
nor UO_1492 (O_1492,N_18259,N_19267);
nand UO_1493 (O_1493,N_18375,N_18149);
xnor UO_1494 (O_1494,N_19065,N_18361);
and UO_1495 (O_1495,N_18164,N_19648);
xnor UO_1496 (O_1496,N_19541,N_18544);
nand UO_1497 (O_1497,N_19523,N_18213);
nor UO_1498 (O_1498,N_19643,N_19340);
nand UO_1499 (O_1499,N_18588,N_18131);
and UO_1500 (O_1500,N_18168,N_19362);
nor UO_1501 (O_1501,N_18309,N_19054);
nor UO_1502 (O_1502,N_18823,N_19005);
xor UO_1503 (O_1503,N_19127,N_19908);
nand UO_1504 (O_1504,N_19131,N_18592);
and UO_1505 (O_1505,N_18581,N_18106);
and UO_1506 (O_1506,N_19170,N_18532);
nor UO_1507 (O_1507,N_18637,N_18471);
and UO_1508 (O_1508,N_19461,N_19087);
nand UO_1509 (O_1509,N_19230,N_19700);
or UO_1510 (O_1510,N_18209,N_18695);
or UO_1511 (O_1511,N_18322,N_18317);
xor UO_1512 (O_1512,N_18713,N_18621);
nor UO_1513 (O_1513,N_19825,N_19211);
nor UO_1514 (O_1514,N_18110,N_18400);
nor UO_1515 (O_1515,N_19073,N_18364);
nand UO_1516 (O_1516,N_19197,N_19199);
xor UO_1517 (O_1517,N_19949,N_19755);
and UO_1518 (O_1518,N_18766,N_19237);
nor UO_1519 (O_1519,N_19967,N_18908);
and UO_1520 (O_1520,N_18652,N_18414);
and UO_1521 (O_1521,N_18652,N_19695);
and UO_1522 (O_1522,N_19730,N_18674);
or UO_1523 (O_1523,N_19511,N_19721);
nand UO_1524 (O_1524,N_18304,N_18769);
and UO_1525 (O_1525,N_18002,N_19638);
nand UO_1526 (O_1526,N_18791,N_19427);
nand UO_1527 (O_1527,N_19107,N_19147);
nor UO_1528 (O_1528,N_19681,N_19785);
or UO_1529 (O_1529,N_19372,N_19444);
nand UO_1530 (O_1530,N_18050,N_18299);
and UO_1531 (O_1531,N_19775,N_18472);
or UO_1532 (O_1532,N_19842,N_18966);
nor UO_1533 (O_1533,N_19881,N_18028);
xnor UO_1534 (O_1534,N_19547,N_19842);
or UO_1535 (O_1535,N_19714,N_18577);
nand UO_1536 (O_1536,N_19604,N_18214);
nor UO_1537 (O_1537,N_18593,N_19356);
xnor UO_1538 (O_1538,N_18864,N_18190);
xor UO_1539 (O_1539,N_18099,N_19135);
nand UO_1540 (O_1540,N_19616,N_19667);
nor UO_1541 (O_1541,N_19691,N_18059);
or UO_1542 (O_1542,N_19759,N_18251);
nand UO_1543 (O_1543,N_18336,N_18274);
xor UO_1544 (O_1544,N_19030,N_19001);
nand UO_1545 (O_1545,N_18841,N_19187);
nand UO_1546 (O_1546,N_18668,N_19674);
nand UO_1547 (O_1547,N_18931,N_19750);
xnor UO_1548 (O_1548,N_19508,N_18606);
xnor UO_1549 (O_1549,N_18863,N_19388);
and UO_1550 (O_1550,N_18581,N_19485);
nor UO_1551 (O_1551,N_18128,N_18216);
or UO_1552 (O_1552,N_18609,N_19672);
nor UO_1553 (O_1553,N_19002,N_19523);
and UO_1554 (O_1554,N_19732,N_19976);
xnor UO_1555 (O_1555,N_18223,N_19050);
and UO_1556 (O_1556,N_18466,N_18366);
nand UO_1557 (O_1557,N_19812,N_19861);
nor UO_1558 (O_1558,N_18686,N_19769);
nor UO_1559 (O_1559,N_18634,N_18063);
nand UO_1560 (O_1560,N_19858,N_18429);
nor UO_1561 (O_1561,N_18848,N_19160);
and UO_1562 (O_1562,N_18878,N_19202);
and UO_1563 (O_1563,N_18473,N_18894);
xor UO_1564 (O_1564,N_19500,N_19039);
nor UO_1565 (O_1565,N_18669,N_19229);
xnor UO_1566 (O_1566,N_18510,N_19632);
and UO_1567 (O_1567,N_19186,N_18904);
or UO_1568 (O_1568,N_19984,N_18148);
and UO_1569 (O_1569,N_19412,N_18342);
xnor UO_1570 (O_1570,N_18054,N_19377);
nor UO_1571 (O_1571,N_19095,N_19996);
nand UO_1572 (O_1572,N_19321,N_19370);
or UO_1573 (O_1573,N_18157,N_18073);
and UO_1574 (O_1574,N_18140,N_19126);
xnor UO_1575 (O_1575,N_19666,N_19178);
and UO_1576 (O_1576,N_18516,N_19223);
or UO_1577 (O_1577,N_19921,N_18435);
nor UO_1578 (O_1578,N_19029,N_19947);
and UO_1579 (O_1579,N_18468,N_18150);
or UO_1580 (O_1580,N_18551,N_19628);
xnor UO_1581 (O_1581,N_19182,N_18711);
nor UO_1582 (O_1582,N_19676,N_19172);
xnor UO_1583 (O_1583,N_18924,N_19685);
or UO_1584 (O_1584,N_18576,N_18277);
xnor UO_1585 (O_1585,N_19907,N_19243);
xnor UO_1586 (O_1586,N_18521,N_19168);
xor UO_1587 (O_1587,N_19336,N_19154);
nand UO_1588 (O_1588,N_18548,N_19686);
nor UO_1589 (O_1589,N_19472,N_18567);
nor UO_1590 (O_1590,N_19905,N_18923);
and UO_1591 (O_1591,N_18902,N_19606);
nor UO_1592 (O_1592,N_19784,N_19754);
nor UO_1593 (O_1593,N_19815,N_18238);
and UO_1594 (O_1594,N_19586,N_18594);
nand UO_1595 (O_1595,N_18224,N_18219);
nor UO_1596 (O_1596,N_18216,N_18303);
and UO_1597 (O_1597,N_19783,N_18461);
nand UO_1598 (O_1598,N_19072,N_19905);
nor UO_1599 (O_1599,N_18973,N_18741);
or UO_1600 (O_1600,N_18296,N_19476);
or UO_1601 (O_1601,N_19866,N_19517);
nor UO_1602 (O_1602,N_19554,N_19804);
nor UO_1603 (O_1603,N_18970,N_18236);
or UO_1604 (O_1604,N_19717,N_19600);
nor UO_1605 (O_1605,N_19648,N_18566);
nand UO_1606 (O_1606,N_19896,N_18773);
and UO_1607 (O_1607,N_18397,N_18112);
or UO_1608 (O_1608,N_19210,N_18416);
nand UO_1609 (O_1609,N_18498,N_18018);
nand UO_1610 (O_1610,N_18410,N_18883);
or UO_1611 (O_1611,N_19642,N_19172);
nand UO_1612 (O_1612,N_18086,N_18825);
or UO_1613 (O_1613,N_19866,N_19037);
or UO_1614 (O_1614,N_18057,N_18095);
nand UO_1615 (O_1615,N_19114,N_18115);
and UO_1616 (O_1616,N_18395,N_18759);
or UO_1617 (O_1617,N_19382,N_19635);
and UO_1618 (O_1618,N_18274,N_19544);
nor UO_1619 (O_1619,N_19661,N_18120);
xnor UO_1620 (O_1620,N_19624,N_18698);
nor UO_1621 (O_1621,N_19944,N_19340);
nor UO_1622 (O_1622,N_18790,N_19211);
or UO_1623 (O_1623,N_19923,N_18507);
or UO_1624 (O_1624,N_18548,N_18763);
and UO_1625 (O_1625,N_18906,N_18140);
nor UO_1626 (O_1626,N_19176,N_19471);
or UO_1627 (O_1627,N_19496,N_19407);
nor UO_1628 (O_1628,N_19116,N_19939);
nor UO_1629 (O_1629,N_19193,N_19104);
or UO_1630 (O_1630,N_19711,N_18952);
nor UO_1631 (O_1631,N_19609,N_18580);
nor UO_1632 (O_1632,N_19886,N_18064);
or UO_1633 (O_1633,N_19867,N_19592);
or UO_1634 (O_1634,N_19121,N_19574);
xnor UO_1635 (O_1635,N_19244,N_19285);
nand UO_1636 (O_1636,N_19662,N_19774);
or UO_1637 (O_1637,N_19591,N_18866);
nor UO_1638 (O_1638,N_19091,N_18223);
or UO_1639 (O_1639,N_18647,N_19844);
or UO_1640 (O_1640,N_18477,N_18966);
xnor UO_1641 (O_1641,N_19029,N_18468);
nor UO_1642 (O_1642,N_19602,N_19717);
nor UO_1643 (O_1643,N_19249,N_19786);
xnor UO_1644 (O_1644,N_19421,N_18810);
nand UO_1645 (O_1645,N_18774,N_18172);
or UO_1646 (O_1646,N_18750,N_19374);
nand UO_1647 (O_1647,N_19221,N_18114);
nand UO_1648 (O_1648,N_19970,N_19159);
nand UO_1649 (O_1649,N_19459,N_18392);
nand UO_1650 (O_1650,N_18593,N_19544);
nor UO_1651 (O_1651,N_19992,N_19331);
nor UO_1652 (O_1652,N_18471,N_18957);
xnor UO_1653 (O_1653,N_19100,N_19451);
nand UO_1654 (O_1654,N_18755,N_19685);
nor UO_1655 (O_1655,N_19858,N_19133);
nor UO_1656 (O_1656,N_19491,N_18008);
xor UO_1657 (O_1657,N_19527,N_19705);
or UO_1658 (O_1658,N_18143,N_18476);
xnor UO_1659 (O_1659,N_19338,N_19723);
or UO_1660 (O_1660,N_18375,N_19284);
nand UO_1661 (O_1661,N_19822,N_19251);
xor UO_1662 (O_1662,N_19321,N_18359);
and UO_1663 (O_1663,N_18438,N_19511);
xnor UO_1664 (O_1664,N_18043,N_18545);
nor UO_1665 (O_1665,N_18825,N_18113);
nand UO_1666 (O_1666,N_19312,N_18601);
nor UO_1667 (O_1667,N_19596,N_18824);
xor UO_1668 (O_1668,N_19218,N_19628);
xor UO_1669 (O_1669,N_18900,N_18124);
xnor UO_1670 (O_1670,N_18647,N_18418);
nand UO_1671 (O_1671,N_19414,N_19336);
xor UO_1672 (O_1672,N_19660,N_18641);
nand UO_1673 (O_1673,N_19955,N_19938);
and UO_1674 (O_1674,N_19663,N_18081);
nor UO_1675 (O_1675,N_19169,N_19147);
and UO_1676 (O_1676,N_18756,N_19255);
xor UO_1677 (O_1677,N_19469,N_19905);
xnor UO_1678 (O_1678,N_19864,N_18733);
nand UO_1679 (O_1679,N_19164,N_18228);
nor UO_1680 (O_1680,N_18420,N_19316);
nor UO_1681 (O_1681,N_18717,N_18203);
and UO_1682 (O_1682,N_18366,N_18977);
or UO_1683 (O_1683,N_19153,N_18249);
and UO_1684 (O_1684,N_18746,N_19460);
xor UO_1685 (O_1685,N_18869,N_18054);
nor UO_1686 (O_1686,N_18641,N_19411);
nand UO_1687 (O_1687,N_18614,N_19356);
or UO_1688 (O_1688,N_18965,N_19863);
and UO_1689 (O_1689,N_18549,N_19232);
and UO_1690 (O_1690,N_18623,N_19182);
and UO_1691 (O_1691,N_18044,N_18992);
and UO_1692 (O_1692,N_18720,N_18283);
nor UO_1693 (O_1693,N_18947,N_18779);
or UO_1694 (O_1694,N_19502,N_19622);
nand UO_1695 (O_1695,N_18699,N_19134);
or UO_1696 (O_1696,N_18267,N_19871);
nor UO_1697 (O_1697,N_18056,N_18486);
and UO_1698 (O_1698,N_18497,N_19159);
or UO_1699 (O_1699,N_18679,N_18530);
nand UO_1700 (O_1700,N_19437,N_18016);
nor UO_1701 (O_1701,N_18606,N_18765);
or UO_1702 (O_1702,N_18426,N_18348);
or UO_1703 (O_1703,N_18343,N_19863);
nand UO_1704 (O_1704,N_18235,N_18892);
nand UO_1705 (O_1705,N_18731,N_18630);
nor UO_1706 (O_1706,N_19027,N_18083);
nor UO_1707 (O_1707,N_18415,N_18701);
nor UO_1708 (O_1708,N_18960,N_19902);
or UO_1709 (O_1709,N_18519,N_18660);
nand UO_1710 (O_1710,N_18417,N_18506);
nor UO_1711 (O_1711,N_19097,N_18314);
xnor UO_1712 (O_1712,N_18691,N_19800);
nor UO_1713 (O_1713,N_18047,N_18940);
nor UO_1714 (O_1714,N_19275,N_19378);
nand UO_1715 (O_1715,N_18793,N_19570);
nand UO_1716 (O_1716,N_19914,N_18602);
xnor UO_1717 (O_1717,N_19137,N_19478);
and UO_1718 (O_1718,N_19058,N_19351);
nor UO_1719 (O_1719,N_19347,N_19064);
xor UO_1720 (O_1720,N_19321,N_18237);
nor UO_1721 (O_1721,N_18107,N_19593);
or UO_1722 (O_1722,N_19468,N_18818);
and UO_1723 (O_1723,N_19695,N_19659);
xor UO_1724 (O_1724,N_18083,N_18591);
or UO_1725 (O_1725,N_18203,N_19426);
and UO_1726 (O_1726,N_18157,N_18192);
or UO_1727 (O_1727,N_19390,N_19384);
nand UO_1728 (O_1728,N_18967,N_19339);
xor UO_1729 (O_1729,N_18054,N_19634);
nor UO_1730 (O_1730,N_18821,N_19982);
nor UO_1731 (O_1731,N_19140,N_19239);
and UO_1732 (O_1732,N_19115,N_18236);
and UO_1733 (O_1733,N_18570,N_18538);
and UO_1734 (O_1734,N_19513,N_18094);
and UO_1735 (O_1735,N_19037,N_18691);
or UO_1736 (O_1736,N_18371,N_18198);
or UO_1737 (O_1737,N_19174,N_19623);
nor UO_1738 (O_1738,N_18626,N_18166);
xor UO_1739 (O_1739,N_18728,N_19002);
xor UO_1740 (O_1740,N_19968,N_19012);
and UO_1741 (O_1741,N_19832,N_18254);
xnor UO_1742 (O_1742,N_18178,N_19497);
and UO_1743 (O_1743,N_18648,N_18244);
nand UO_1744 (O_1744,N_18414,N_18323);
nor UO_1745 (O_1745,N_18869,N_18344);
xor UO_1746 (O_1746,N_18165,N_19205);
or UO_1747 (O_1747,N_19030,N_19669);
and UO_1748 (O_1748,N_19461,N_19343);
and UO_1749 (O_1749,N_19896,N_18763);
nor UO_1750 (O_1750,N_19479,N_19898);
nor UO_1751 (O_1751,N_19430,N_19038);
or UO_1752 (O_1752,N_18292,N_18811);
and UO_1753 (O_1753,N_19321,N_19414);
nor UO_1754 (O_1754,N_19517,N_18962);
nand UO_1755 (O_1755,N_18419,N_19884);
nor UO_1756 (O_1756,N_19840,N_18098);
and UO_1757 (O_1757,N_19259,N_19866);
or UO_1758 (O_1758,N_19348,N_18897);
nor UO_1759 (O_1759,N_18382,N_18839);
nor UO_1760 (O_1760,N_19986,N_19930);
nand UO_1761 (O_1761,N_19954,N_18253);
or UO_1762 (O_1762,N_18692,N_18431);
or UO_1763 (O_1763,N_19207,N_18309);
xnor UO_1764 (O_1764,N_19421,N_19551);
nor UO_1765 (O_1765,N_18474,N_18608);
xnor UO_1766 (O_1766,N_19312,N_18377);
nand UO_1767 (O_1767,N_19210,N_19479);
nand UO_1768 (O_1768,N_18846,N_18129);
nor UO_1769 (O_1769,N_19582,N_19099);
nor UO_1770 (O_1770,N_18858,N_19380);
and UO_1771 (O_1771,N_18106,N_19297);
xnor UO_1772 (O_1772,N_19559,N_19631);
nor UO_1773 (O_1773,N_18673,N_19902);
nand UO_1774 (O_1774,N_19684,N_18910);
xor UO_1775 (O_1775,N_19863,N_19590);
or UO_1776 (O_1776,N_18108,N_19618);
nand UO_1777 (O_1777,N_18646,N_18864);
and UO_1778 (O_1778,N_18726,N_19595);
nor UO_1779 (O_1779,N_18091,N_18984);
and UO_1780 (O_1780,N_19053,N_18536);
and UO_1781 (O_1781,N_18505,N_19420);
nor UO_1782 (O_1782,N_19502,N_18249);
nor UO_1783 (O_1783,N_19103,N_19340);
xor UO_1784 (O_1784,N_19482,N_18886);
xnor UO_1785 (O_1785,N_18559,N_19487);
nand UO_1786 (O_1786,N_19789,N_19590);
xor UO_1787 (O_1787,N_19362,N_18452);
nand UO_1788 (O_1788,N_18012,N_18007);
xor UO_1789 (O_1789,N_19868,N_19372);
or UO_1790 (O_1790,N_18833,N_18177);
nand UO_1791 (O_1791,N_19593,N_18245);
nand UO_1792 (O_1792,N_19027,N_19374);
nand UO_1793 (O_1793,N_19124,N_18690);
and UO_1794 (O_1794,N_18431,N_18990);
or UO_1795 (O_1795,N_19139,N_18838);
nor UO_1796 (O_1796,N_19054,N_19816);
and UO_1797 (O_1797,N_18049,N_19215);
nor UO_1798 (O_1798,N_19143,N_19547);
nand UO_1799 (O_1799,N_18757,N_18742);
and UO_1800 (O_1800,N_18584,N_19064);
xnor UO_1801 (O_1801,N_18479,N_19661);
and UO_1802 (O_1802,N_18821,N_18670);
and UO_1803 (O_1803,N_19567,N_18125);
or UO_1804 (O_1804,N_19736,N_19170);
nand UO_1805 (O_1805,N_18852,N_18645);
xor UO_1806 (O_1806,N_18674,N_18945);
and UO_1807 (O_1807,N_19174,N_19170);
or UO_1808 (O_1808,N_18885,N_18091);
xor UO_1809 (O_1809,N_18774,N_18402);
nand UO_1810 (O_1810,N_19425,N_18587);
xor UO_1811 (O_1811,N_18798,N_18265);
nand UO_1812 (O_1812,N_18967,N_19474);
nor UO_1813 (O_1813,N_19115,N_19276);
or UO_1814 (O_1814,N_18343,N_19760);
and UO_1815 (O_1815,N_19812,N_19053);
xnor UO_1816 (O_1816,N_19161,N_19649);
xnor UO_1817 (O_1817,N_18231,N_19020);
and UO_1818 (O_1818,N_18888,N_19759);
nor UO_1819 (O_1819,N_18369,N_18090);
xnor UO_1820 (O_1820,N_19840,N_18521);
nor UO_1821 (O_1821,N_18979,N_19798);
nor UO_1822 (O_1822,N_19623,N_19419);
and UO_1823 (O_1823,N_18311,N_18461);
nor UO_1824 (O_1824,N_18752,N_19467);
nor UO_1825 (O_1825,N_19205,N_19470);
and UO_1826 (O_1826,N_18556,N_19354);
or UO_1827 (O_1827,N_19626,N_18206);
or UO_1828 (O_1828,N_19695,N_19734);
or UO_1829 (O_1829,N_18843,N_18937);
or UO_1830 (O_1830,N_18191,N_19633);
xnor UO_1831 (O_1831,N_19031,N_18985);
nor UO_1832 (O_1832,N_18865,N_18980);
and UO_1833 (O_1833,N_19187,N_19073);
xor UO_1834 (O_1834,N_19929,N_18901);
xnor UO_1835 (O_1835,N_19793,N_18650);
nand UO_1836 (O_1836,N_18212,N_18049);
nor UO_1837 (O_1837,N_19857,N_19034);
and UO_1838 (O_1838,N_18406,N_19906);
nand UO_1839 (O_1839,N_18588,N_19931);
nor UO_1840 (O_1840,N_19649,N_19459);
nand UO_1841 (O_1841,N_18580,N_18453);
or UO_1842 (O_1842,N_18185,N_18130);
nor UO_1843 (O_1843,N_19085,N_18463);
or UO_1844 (O_1844,N_19616,N_19864);
and UO_1845 (O_1845,N_19015,N_19093);
nor UO_1846 (O_1846,N_19188,N_18355);
nor UO_1847 (O_1847,N_19481,N_19273);
and UO_1848 (O_1848,N_19198,N_18463);
xnor UO_1849 (O_1849,N_19446,N_18386);
or UO_1850 (O_1850,N_19551,N_18059);
xnor UO_1851 (O_1851,N_18318,N_19465);
or UO_1852 (O_1852,N_18541,N_19554);
or UO_1853 (O_1853,N_19065,N_18237);
nand UO_1854 (O_1854,N_18565,N_18353);
and UO_1855 (O_1855,N_18760,N_18078);
and UO_1856 (O_1856,N_19923,N_18202);
and UO_1857 (O_1857,N_19199,N_18475);
nand UO_1858 (O_1858,N_18090,N_19261);
or UO_1859 (O_1859,N_18589,N_19906);
or UO_1860 (O_1860,N_19383,N_18942);
nand UO_1861 (O_1861,N_19375,N_19366);
and UO_1862 (O_1862,N_18385,N_19938);
nand UO_1863 (O_1863,N_18420,N_19837);
nand UO_1864 (O_1864,N_19689,N_19084);
or UO_1865 (O_1865,N_19296,N_19028);
xnor UO_1866 (O_1866,N_18458,N_19347);
nor UO_1867 (O_1867,N_19759,N_18902);
and UO_1868 (O_1868,N_18604,N_19049);
nand UO_1869 (O_1869,N_18464,N_18188);
xor UO_1870 (O_1870,N_18482,N_19371);
nand UO_1871 (O_1871,N_18537,N_18920);
or UO_1872 (O_1872,N_19344,N_18451);
nor UO_1873 (O_1873,N_18139,N_18415);
or UO_1874 (O_1874,N_18614,N_18157);
and UO_1875 (O_1875,N_18983,N_19158);
and UO_1876 (O_1876,N_19988,N_18351);
xor UO_1877 (O_1877,N_18402,N_19433);
and UO_1878 (O_1878,N_18859,N_19648);
nand UO_1879 (O_1879,N_18101,N_19725);
nor UO_1880 (O_1880,N_19365,N_19890);
nand UO_1881 (O_1881,N_18697,N_18827);
nand UO_1882 (O_1882,N_19370,N_18555);
nand UO_1883 (O_1883,N_18600,N_19059);
nand UO_1884 (O_1884,N_19353,N_18214);
nand UO_1885 (O_1885,N_18114,N_19907);
nor UO_1886 (O_1886,N_19942,N_19381);
and UO_1887 (O_1887,N_19794,N_19073);
nand UO_1888 (O_1888,N_19464,N_18572);
and UO_1889 (O_1889,N_18577,N_18052);
and UO_1890 (O_1890,N_18680,N_19361);
xor UO_1891 (O_1891,N_18511,N_18800);
xor UO_1892 (O_1892,N_18524,N_19638);
xor UO_1893 (O_1893,N_19030,N_18347);
xor UO_1894 (O_1894,N_19543,N_19449);
or UO_1895 (O_1895,N_19216,N_19036);
and UO_1896 (O_1896,N_18960,N_19122);
and UO_1897 (O_1897,N_18066,N_18140);
nand UO_1898 (O_1898,N_18439,N_18475);
xnor UO_1899 (O_1899,N_19089,N_19337);
or UO_1900 (O_1900,N_18432,N_18845);
or UO_1901 (O_1901,N_18257,N_19546);
and UO_1902 (O_1902,N_18931,N_19194);
or UO_1903 (O_1903,N_19763,N_19657);
nor UO_1904 (O_1904,N_18169,N_19494);
nor UO_1905 (O_1905,N_18629,N_18992);
nor UO_1906 (O_1906,N_19367,N_18365);
nor UO_1907 (O_1907,N_19701,N_19723);
or UO_1908 (O_1908,N_19532,N_18111);
nand UO_1909 (O_1909,N_18607,N_18913);
nor UO_1910 (O_1910,N_19796,N_18171);
nor UO_1911 (O_1911,N_18733,N_19087);
or UO_1912 (O_1912,N_18387,N_18573);
nand UO_1913 (O_1913,N_19638,N_19852);
nor UO_1914 (O_1914,N_19737,N_18853);
nor UO_1915 (O_1915,N_18588,N_18877);
xor UO_1916 (O_1916,N_19618,N_19691);
or UO_1917 (O_1917,N_18045,N_18334);
nor UO_1918 (O_1918,N_19662,N_18655);
or UO_1919 (O_1919,N_19369,N_19653);
and UO_1920 (O_1920,N_18998,N_19176);
or UO_1921 (O_1921,N_18548,N_18908);
or UO_1922 (O_1922,N_19963,N_19858);
and UO_1923 (O_1923,N_18106,N_19722);
nand UO_1924 (O_1924,N_19052,N_19992);
xnor UO_1925 (O_1925,N_19611,N_18463);
xor UO_1926 (O_1926,N_18903,N_19442);
and UO_1927 (O_1927,N_18816,N_18077);
nor UO_1928 (O_1928,N_18793,N_19023);
nor UO_1929 (O_1929,N_18190,N_19496);
and UO_1930 (O_1930,N_19578,N_18029);
nor UO_1931 (O_1931,N_18399,N_19998);
nand UO_1932 (O_1932,N_18393,N_18908);
and UO_1933 (O_1933,N_19932,N_18318);
and UO_1934 (O_1934,N_18921,N_18537);
nor UO_1935 (O_1935,N_19346,N_18642);
nor UO_1936 (O_1936,N_18934,N_19292);
or UO_1937 (O_1937,N_18795,N_19259);
xor UO_1938 (O_1938,N_19905,N_19883);
and UO_1939 (O_1939,N_19661,N_18546);
nand UO_1940 (O_1940,N_18608,N_19366);
xor UO_1941 (O_1941,N_19566,N_19747);
nor UO_1942 (O_1942,N_19698,N_19370);
or UO_1943 (O_1943,N_19993,N_18626);
nor UO_1944 (O_1944,N_18976,N_19726);
nand UO_1945 (O_1945,N_18851,N_19478);
or UO_1946 (O_1946,N_19225,N_19925);
or UO_1947 (O_1947,N_19506,N_19786);
nor UO_1948 (O_1948,N_18080,N_19611);
nor UO_1949 (O_1949,N_18943,N_18710);
and UO_1950 (O_1950,N_19760,N_18897);
and UO_1951 (O_1951,N_19573,N_18279);
and UO_1952 (O_1952,N_19738,N_18850);
nor UO_1953 (O_1953,N_19295,N_19050);
nor UO_1954 (O_1954,N_18195,N_18897);
xor UO_1955 (O_1955,N_19322,N_18533);
nor UO_1956 (O_1956,N_18006,N_18962);
nand UO_1957 (O_1957,N_19523,N_19408);
nand UO_1958 (O_1958,N_18715,N_18049);
or UO_1959 (O_1959,N_18073,N_19251);
or UO_1960 (O_1960,N_19835,N_18068);
nor UO_1961 (O_1961,N_19963,N_18225);
or UO_1962 (O_1962,N_19263,N_19488);
and UO_1963 (O_1963,N_19816,N_19977);
or UO_1964 (O_1964,N_18054,N_18597);
xnor UO_1965 (O_1965,N_18241,N_19732);
nor UO_1966 (O_1966,N_18814,N_18423);
or UO_1967 (O_1967,N_19073,N_19290);
nor UO_1968 (O_1968,N_18423,N_19445);
nor UO_1969 (O_1969,N_19374,N_19618);
or UO_1970 (O_1970,N_18154,N_19735);
xnor UO_1971 (O_1971,N_18393,N_18511);
xor UO_1972 (O_1972,N_18343,N_19102);
nand UO_1973 (O_1973,N_19013,N_18344);
nor UO_1974 (O_1974,N_18495,N_18316);
or UO_1975 (O_1975,N_19878,N_19688);
nor UO_1976 (O_1976,N_19608,N_18759);
nor UO_1977 (O_1977,N_19478,N_19047);
nor UO_1978 (O_1978,N_18530,N_18956);
xnor UO_1979 (O_1979,N_18894,N_19888);
or UO_1980 (O_1980,N_19119,N_18318);
nand UO_1981 (O_1981,N_18695,N_18583);
xor UO_1982 (O_1982,N_18136,N_19335);
and UO_1983 (O_1983,N_19962,N_19163);
or UO_1984 (O_1984,N_18251,N_19330);
nand UO_1985 (O_1985,N_19255,N_18806);
nor UO_1986 (O_1986,N_19258,N_18505);
xnor UO_1987 (O_1987,N_19236,N_18317);
nor UO_1988 (O_1988,N_18111,N_19590);
nand UO_1989 (O_1989,N_18671,N_18321);
nor UO_1990 (O_1990,N_18488,N_19292);
nor UO_1991 (O_1991,N_19283,N_18152);
nand UO_1992 (O_1992,N_19512,N_19655);
nand UO_1993 (O_1993,N_19533,N_18970);
xnor UO_1994 (O_1994,N_18168,N_18495);
and UO_1995 (O_1995,N_19188,N_18895);
xor UO_1996 (O_1996,N_18358,N_18632);
and UO_1997 (O_1997,N_18900,N_18398);
nor UO_1998 (O_1998,N_18302,N_18751);
and UO_1999 (O_1999,N_19403,N_19796);
nor UO_2000 (O_2000,N_19156,N_19768);
or UO_2001 (O_2001,N_19485,N_19565);
and UO_2002 (O_2002,N_19269,N_19656);
and UO_2003 (O_2003,N_19427,N_18047);
xnor UO_2004 (O_2004,N_19913,N_18047);
and UO_2005 (O_2005,N_18648,N_19354);
xnor UO_2006 (O_2006,N_19765,N_19196);
xor UO_2007 (O_2007,N_19639,N_19551);
nor UO_2008 (O_2008,N_19141,N_18332);
nor UO_2009 (O_2009,N_18194,N_19489);
xor UO_2010 (O_2010,N_18083,N_19832);
nand UO_2011 (O_2011,N_19272,N_19012);
nand UO_2012 (O_2012,N_18257,N_19523);
nor UO_2013 (O_2013,N_18355,N_18210);
or UO_2014 (O_2014,N_18759,N_18117);
nor UO_2015 (O_2015,N_19242,N_18179);
nor UO_2016 (O_2016,N_19569,N_19882);
nor UO_2017 (O_2017,N_19175,N_18924);
nor UO_2018 (O_2018,N_18441,N_19594);
xor UO_2019 (O_2019,N_18690,N_18172);
nor UO_2020 (O_2020,N_18851,N_19147);
nor UO_2021 (O_2021,N_18265,N_18841);
nor UO_2022 (O_2022,N_18757,N_19558);
nor UO_2023 (O_2023,N_18145,N_19112);
nor UO_2024 (O_2024,N_18327,N_19277);
xnor UO_2025 (O_2025,N_18607,N_18550);
nor UO_2026 (O_2026,N_18075,N_19643);
xor UO_2027 (O_2027,N_19308,N_19259);
nand UO_2028 (O_2028,N_19028,N_19355);
nor UO_2029 (O_2029,N_18337,N_18214);
nand UO_2030 (O_2030,N_18898,N_19280);
nand UO_2031 (O_2031,N_19945,N_19286);
xor UO_2032 (O_2032,N_18431,N_19427);
nor UO_2033 (O_2033,N_18352,N_18222);
and UO_2034 (O_2034,N_18702,N_19701);
nor UO_2035 (O_2035,N_18254,N_19859);
and UO_2036 (O_2036,N_18541,N_18291);
or UO_2037 (O_2037,N_19929,N_18823);
nand UO_2038 (O_2038,N_18149,N_18238);
or UO_2039 (O_2039,N_19383,N_18775);
nor UO_2040 (O_2040,N_18091,N_19148);
or UO_2041 (O_2041,N_18172,N_18189);
and UO_2042 (O_2042,N_18260,N_18893);
xnor UO_2043 (O_2043,N_18970,N_18281);
and UO_2044 (O_2044,N_19344,N_18698);
and UO_2045 (O_2045,N_18464,N_18347);
nand UO_2046 (O_2046,N_18180,N_19822);
or UO_2047 (O_2047,N_18328,N_19943);
or UO_2048 (O_2048,N_19740,N_19846);
xor UO_2049 (O_2049,N_18464,N_18499);
nand UO_2050 (O_2050,N_19557,N_19039);
xor UO_2051 (O_2051,N_19399,N_19238);
nor UO_2052 (O_2052,N_18236,N_19590);
xor UO_2053 (O_2053,N_19319,N_19747);
and UO_2054 (O_2054,N_19956,N_19305);
nand UO_2055 (O_2055,N_18949,N_18894);
nand UO_2056 (O_2056,N_19996,N_19673);
nor UO_2057 (O_2057,N_18135,N_19933);
nand UO_2058 (O_2058,N_19049,N_18555);
nand UO_2059 (O_2059,N_18576,N_19438);
or UO_2060 (O_2060,N_19007,N_18932);
xnor UO_2061 (O_2061,N_18951,N_19091);
or UO_2062 (O_2062,N_19489,N_19734);
nor UO_2063 (O_2063,N_18812,N_19423);
nand UO_2064 (O_2064,N_18322,N_19372);
nor UO_2065 (O_2065,N_19071,N_19044);
xor UO_2066 (O_2066,N_19966,N_19954);
xnor UO_2067 (O_2067,N_18759,N_19414);
nand UO_2068 (O_2068,N_18777,N_19550);
xnor UO_2069 (O_2069,N_19699,N_18668);
nand UO_2070 (O_2070,N_19061,N_18234);
nor UO_2071 (O_2071,N_19126,N_19630);
xnor UO_2072 (O_2072,N_19636,N_18479);
nor UO_2073 (O_2073,N_19245,N_19147);
or UO_2074 (O_2074,N_18960,N_19498);
or UO_2075 (O_2075,N_19027,N_18323);
xor UO_2076 (O_2076,N_18868,N_19920);
nor UO_2077 (O_2077,N_19129,N_18868);
nor UO_2078 (O_2078,N_18363,N_18547);
xor UO_2079 (O_2079,N_19080,N_19256);
nand UO_2080 (O_2080,N_19743,N_19971);
nor UO_2081 (O_2081,N_19345,N_19197);
nand UO_2082 (O_2082,N_18964,N_19430);
nand UO_2083 (O_2083,N_19732,N_18613);
nor UO_2084 (O_2084,N_19331,N_19224);
or UO_2085 (O_2085,N_19091,N_18106);
or UO_2086 (O_2086,N_18065,N_18129);
or UO_2087 (O_2087,N_19122,N_19379);
or UO_2088 (O_2088,N_18149,N_18983);
or UO_2089 (O_2089,N_18902,N_18533);
nand UO_2090 (O_2090,N_19597,N_19797);
or UO_2091 (O_2091,N_18993,N_19563);
and UO_2092 (O_2092,N_19624,N_19714);
nor UO_2093 (O_2093,N_18801,N_19450);
nand UO_2094 (O_2094,N_18182,N_18643);
or UO_2095 (O_2095,N_18115,N_19752);
and UO_2096 (O_2096,N_19207,N_18361);
nand UO_2097 (O_2097,N_19292,N_19325);
or UO_2098 (O_2098,N_19383,N_19148);
and UO_2099 (O_2099,N_19205,N_19615);
and UO_2100 (O_2100,N_19711,N_18701);
nand UO_2101 (O_2101,N_19221,N_19028);
xor UO_2102 (O_2102,N_19262,N_18512);
and UO_2103 (O_2103,N_19205,N_18721);
or UO_2104 (O_2104,N_18630,N_18032);
nand UO_2105 (O_2105,N_19589,N_19352);
nand UO_2106 (O_2106,N_19637,N_18307);
or UO_2107 (O_2107,N_19121,N_19840);
nand UO_2108 (O_2108,N_18423,N_18445);
or UO_2109 (O_2109,N_19777,N_19491);
nor UO_2110 (O_2110,N_18768,N_18104);
and UO_2111 (O_2111,N_19602,N_18690);
nand UO_2112 (O_2112,N_18935,N_18923);
or UO_2113 (O_2113,N_18781,N_18186);
and UO_2114 (O_2114,N_18303,N_18254);
or UO_2115 (O_2115,N_18308,N_18319);
nor UO_2116 (O_2116,N_18771,N_19816);
and UO_2117 (O_2117,N_19207,N_18682);
nor UO_2118 (O_2118,N_19857,N_19498);
nor UO_2119 (O_2119,N_19344,N_18909);
nor UO_2120 (O_2120,N_18811,N_19525);
xor UO_2121 (O_2121,N_19400,N_19519);
nand UO_2122 (O_2122,N_19705,N_18000);
and UO_2123 (O_2123,N_18085,N_18301);
nand UO_2124 (O_2124,N_18569,N_19628);
nor UO_2125 (O_2125,N_19177,N_18762);
nand UO_2126 (O_2126,N_19841,N_18835);
nor UO_2127 (O_2127,N_18701,N_19976);
or UO_2128 (O_2128,N_19312,N_19202);
nand UO_2129 (O_2129,N_19954,N_18020);
xnor UO_2130 (O_2130,N_18134,N_19700);
and UO_2131 (O_2131,N_18344,N_18520);
nand UO_2132 (O_2132,N_18237,N_18874);
nor UO_2133 (O_2133,N_18539,N_18327);
nand UO_2134 (O_2134,N_19085,N_18558);
xor UO_2135 (O_2135,N_19228,N_19769);
or UO_2136 (O_2136,N_19581,N_19658);
nand UO_2137 (O_2137,N_19094,N_18882);
nand UO_2138 (O_2138,N_19415,N_18647);
and UO_2139 (O_2139,N_18594,N_19812);
and UO_2140 (O_2140,N_19925,N_18520);
nand UO_2141 (O_2141,N_19812,N_18845);
and UO_2142 (O_2142,N_19346,N_18697);
and UO_2143 (O_2143,N_19556,N_19597);
nor UO_2144 (O_2144,N_19755,N_18963);
or UO_2145 (O_2145,N_18430,N_19897);
nand UO_2146 (O_2146,N_18082,N_18188);
nand UO_2147 (O_2147,N_18228,N_19101);
and UO_2148 (O_2148,N_19277,N_19750);
xor UO_2149 (O_2149,N_18924,N_19393);
nand UO_2150 (O_2150,N_19021,N_19207);
xnor UO_2151 (O_2151,N_18994,N_19771);
nand UO_2152 (O_2152,N_18301,N_18600);
or UO_2153 (O_2153,N_18446,N_18019);
nand UO_2154 (O_2154,N_18646,N_19590);
nand UO_2155 (O_2155,N_19093,N_19867);
nor UO_2156 (O_2156,N_18642,N_18767);
nand UO_2157 (O_2157,N_18638,N_18121);
xnor UO_2158 (O_2158,N_19648,N_18721);
nand UO_2159 (O_2159,N_18385,N_18178);
or UO_2160 (O_2160,N_19776,N_19437);
nand UO_2161 (O_2161,N_18975,N_18184);
nor UO_2162 (O_2162,N_19650,N_18719);
xor UO_2163 (O_2163,N_19915,N_18123);
or UO_2164 (O_2164,N_19921,N_19900);
nand UO_2165 (O_2165,N_18484,N_19680);
and UO_2166 (O_2166,N_18909,N_18062);
nor UO_2167 (O_2167,N_18648,N_19301);
or UO_2168 (O_2168,N_18139,N_19222);
nor UO_2169 (O_2169,N_19149,N_19492);
nand UO_2170 (O_2170,N_18772,N_18358);
xnor UO_2171 (O_2171,N_19639,N_18593);
or UO_2172 (O_2172,N_19510,N_19515);
and UO_2173 (O_2173,N_19577,N_19385);
nor UO_2174 (O_2174,N_18053,N_18102);
nand UO_2175 (O_2175,N_19544,N_19041);
nand UO_2176 (O_2176,N_19302,N_18552);
xnor UO_2177 (O_2177,N_19690,N_19931);
nand UO_2178 (O_2178,N_18585,N_18044);
or UO_2179 (O_2179,N_19284,N_18428);
and UO_2180 (O_2180,N_19880,N_18863);
xor UO_2181 (O_2181,N_19273,N_18372);
xnor UO_2182 (O_2182,N_19534,N_18034);
xnor UO_2183 (O_2183,N_18220,N_19955);
and UO_2184 (O_2184,N_18937,N_19073);
xor UO_2185 (O_2185,N_18572,N_19511);
and UO_2186 (O_2186,N_19793,N_19983);
or UO_2187 (O_2187,N_19903,N_19271);
and UO_2188 (O_2188,N_19253,N_18490);
nor UO_2189 (O_2189,N_18279,N_19901);
or UO_2190 (O_2190,N_19156,N_19999);
and UO_2191 (O_2191,N_19448,N_18075);
nand UO_2192 (O_2192,N_19554,N_19767);
and UO_2193 (O_2193,N_19317,N_19922);
or UO_2194 (O_2194,N_19787,N_18056);
nor UO_2195 (O_2195,N_18350,N_18931);
or UO_2196 (O_2196,N_18363,N_18952);
and UO_2197 (O_2197,N_19553,N_18276);
and UO_2198 (O_2198,N_18724,N_19271);
nor UO_2199 (O_2199,N_18896,N_18325);
nand UO_2200 (O_2200,N_18295,N_19375);
xnor UO_2201 (O_2201,N_18370,N_18573);
nand UO_2202 (O_2202,N_18086,N_18768);
xnor UO_2203 (O_2203,N_19385,N_19699);
xor UO_2204 (O_2204,N_19390,N_18095);
or UO_2205 (O_2205,N_18667,N_18975);
nor UO_2206 (O_2206,N_19185,N_18745);
or UO_2207 (O_2207,N_18797,N_18814);
nor UO_2208 (O_2208,N_19191,N_18303);
or UO_2209 (O_2209,N_18654,N_19571);
nor UO_2210 (O_2210,N_18892,N_19263);
nor UO_2211 (O_2211,N_18178,N_19467);
and UO_2212 (O_2212,N_18189,N_18477);
nand UO_2213 (O_2213,N_19351,N_19260);
and UO_2214 (O_2214,N_19383,N_18538);
and UO_2215 (O_2215,N_18394,N_19689);
or UO_2216 (O_2216,N_19699,N_18714);
nand UO_2217 (O_2217,N_19959,N_19633);
nand UO_2218 (O_2218,N_19584,N_19165);
or UO_2219 (O_2219,N_18925,N_18200);
xnor UO_2220 (O_2220,N_18776,N_18807);
nand UO_2221 (O_2221,N_18992,N_18644);
nand UO_2222 (O_2222,N_18371,N_19532);
nand UO_2223 (O_2223,N_18752,N_18730);
or UO_2224 (O_2224,N_19299,N_18513);
nor UO_2225 (O_2225,N_19833,N_18699);
or UO_2226 (O_2226,N_18606,N_18813);
or UO_2227 (O_2227,N_18118,N_19180);
or UO_2228 (O_2228,N_19261,N_19343);
xor UO_2229 (O_2229,N_19054,N_18512);
or UO_2230 (O_2230,N_19121,N_18182);
nor UO_2231 (O_2231,N_19752,N_19623);
xnor UO_2232 (O_2232,N_19290,N_19706);
xnor UO_2233 (O_2233,N_18719,N_18858);
nand UO_2234 (O_2234,N_19730,N_19142);
or UO_2235 (O_2235,N_18221,N_19749);
and UO_2236 (O_2236,N_19431,N_18428);
or UO_2237 (O_2237,N_18870,N_19829);
nand UO_2238 (O_2238,N_18809,N_18364);
xor UO_2239 (O_2239,N_18095,N_18529);
xnor UO_2240 (O_2240,N_19290,N_19770);
or UO_2241 (O_2241,N_18972,N_19091);
nor UO_2242 (O_2242,N_18096,N_19791);
nand UO_2243 (O_2243,N_19648,N_19607);
and UO_2244 (O_2244,N_19750,N_19881);
nand UO_2245 (O_2245,N_19261,N_19158);
nand UO_2246 (O_2246,N_18532,N_18072);
or UO_2247 (O_2247,N_19222,N_18802);
and UO_2248 (O_2248,N_19926,N_18641);
or UO_2249 (O_2249,N_18914,N_19557);
nor UO_2250 (O_2250,N_18949,N_18563);
nor UO_2251 (O_2251,N_19698,N_19912);
nand UO_2252 (O_2252,N_18198,N_19495);
nor UO_2253 (O_2253,N_19399,N_18382);
nand UO_2254 (O_2254,N_18609,N_19677);
or UO_2255 (O_2255,N_18032,N_19370);
or UO_2256 (O_2256,N_18271,N_18210);
or UO_2257 (O_2257,N_18161,N_18151);
nor UO_2258 (O_2258,N_18474,N_19047);
xor UO_2259 (O_2259,N_19888,N_19343);
xor UO_2260 (O_2260,N_18465,N_19486);
nand UO_2261 (O_2261,N_18198,N_19148);
or UO_2262 (O_2262,N_19536,N_18976);
xnor UO_2263 (O_2263,N_19300,N_19916);
and UO_2264 (O_2264,N_18053,N_19281);
and UO_2265 (O_2265,N_18807,N_18651);
nor UO_2266 (O_2266,N_18509,N_19062);
nand UO_2267 (O_2267,N_18879,N_19424);
or UO_2268 (O_2268,N_18109,N_18427);
nand UO_2269 (O_2269,N_18243,N_19106);
or UO_2270 (O_2270,N_19077,N_18348);
nand UO_2271 (O_2271,N_19923,N_18162);
nor UO_2272 (O_2272,N_19798,N_19492);
nor UO_2273 (O_2273,N_18479,N_19875);
or UO_2274 (O_2274,N_19060,N_18716);
nor UO_2275 (O_2275,N_18680,N_18832);
nand UO_2276 (O_2276,N_19965,N_19361);
nand UO_2277 (O_2277,N_19096,N_18530);
nand UO_2278 (O_2278,N_18789,N_19609);
xnor UO_2279 (O_2279,N_18818,N_19271);
xnor UO_2280 (O_2280,N_19514,N_19448);
nor UO_2281 (O_2281,N_19018,N_19477);
and UO_2282 (O_2282,N_19517,N_18798);
xnor UO_2283 (O_2283,N_19835,N_18133);
and UO_2284 (O_2284,N_18661,N_18070);
xor UO_2285 (O_2285,N_19364,N_18352);
xor UO_2286 (O_2286,N_18404,N_18160);
and UO_2287 (O_2287,N_19923,N_19307);
and UO_2288 (O_2288,N_19790,N_18011);
xor UO_2289 (O_2289,N_18534,N_18888);
xnor UO_2290 (O_2290,N_18537,N_18268);
xnor UO_2291 (O_2291,N_18017,N_19183);
nor UO_2292 (O_2292,N_19129,N_18804);
or UO_2293 (O_2293,N_18860,N_18468);
or UO_2294 (O_2294,N_18796,N_19914);
xnor UO_2295 (O_2295,N_18506,N_19721);
and UO_2296 (O_2296,N_19317,N_19731);
nand UO_2297 (O_2297,N_19469,N_18688);
nand UO_2298 (O_2298,N_18296,N_18437);
nor UO_2299 (O_2299,N_18885,N_18198);
nor UO_2300 (O_2300,N_18661,N_18532);
nor UO_2301 (O_2301,N_18051,N_19300);
nand UO_2302 (O_2302,N_18416,N_19782);
and UO_2303 (O_2303,N_19666,N_18572);
nand UO_2304 (O_2304,N_18597,N_19708);
or UO_2305 (O_2305,N_18890,N_19112);
nor UO_2306 (O_2306,N_18316,N_19934);
and UO_2307 (O_2307,N_18153,N_19714);
nor UO_2308 (O_2308,N_19185,N_18831);
or UO_2309 (O_2309,N_19396,N_18607);
nor UO_2310 (O_2310,N_19969,N_19079);
and UO_2311 (O_2311,N_19395,N_18693);
nand UO_2312 (O_2312,N_19239,N_19668);
nand UO_2313 (O_2313,N_19817,N_19584);
or UO_2314 (O_2314,N_19854,N_19762);
xnor UO_2315 (O_2315,N_18758,N_18225);
and UO_2316 (O_2316,N_18078,N_18129);
xor UO_2317 (O_2317,N_18386,N_18291);
xnor UO_2318 (O_2318,N_19125,N_18343);
or UO_2319 (O_2319,N_18062,N_19208);
nand UO_2320 (O_2320,N_19195,N_18474);
nor UO_2321 (O_2321,N_18206,N_19261);
or UO_2322 (O_2322,N_18144,N_19299);
or UO_2323 (O_2323,N_18925,N_18288);
or UO_2324 (O_2324,N_19627,N_18357);
nor UO_2325 (O_2325,N_18228,N_18790);
nor UO_2326 (O_2326,N_18650,N_18425);
and UO_2327 (O_2327,N_19973,N_18431);
nand UO_2328 (O_2328,N_19205,N_19329);
nand UO_2329 (O_2329,N_19328,N_19366);
nor UO_2330 (O_2330,N_19533,N_18387);
nor UO_2331 (O_2331,N_18539,N_19186);
nor UO_2332 (O_2332,N_18783,N_18935);
nand UO_2333 (O_2333,N_18989,N_19692);
or UO_2334 (O_2334,N_18469,N_18632);
or UO_2335 (O_2335,N_19977,N_19005);
or UO_2336 (O_2336,N_19269,N_19923);
xor UO_2337 (O_2337,N_19326,N_18267);
nor UO_2338 (O_2338,N_19294,N_19749);
or UO_2339 (O_2339,N_19040,N_19314);
or UO_2340 (O_2340,N_18098,N_19342);
and UO_2341 (O_2341,N_18318,N_18320);
nor UO_2342 (O_2342,N_18462,N_19390);
xnor UO_2343 (O_2343,N_19140,N_18320);
or UO_2344 (O_2344,N_19978,N_18401);
nor UO_2345 (O_2345,N_18991,N_18867);
or UO_2346 (O_2346,N_19384,N_19512);
xor UO_2347 (O_2347,N_19589,N_19940);
nor UO_2348 (O_2348,N_19274,N_18792);
nor UO_2349 (O_2349,N_18890,N_19687);
nand UO_2350 (O_2350,N_19547,N_18379);
and UO_2351 (O_2351,N_18840,N_19875);
nor UO_2352 (O_2352,N_18037,N_19993);
nor UO_2353 (O_2353,N_19546,N_18436);
nor UO_2354 (O_2354,N_18411,N_19843);
and UO_2355 (O_2355,N_19565,N_18833);
nand UO_2356 (O_2356,N_18080,N_18136);
nand UO_2357 (O_2357,N_19539,N_19406);
xor UO_2358 (O_2358,N_19252,N_19984);
nor UO_2359 (O_2359,N_18074,N_18730);
xor UO_2360 (O_2360,N_19775,N_19856);
and UO_2361 (O_2361,N_19666,N_18462);
xor UO_2362 (O_2362,N_19845,N_19444);
nand UO_2363 (O_2363,N_18968,N_18599);
nand UO_2364 (O_2364,N_19840,N_19423);
and UO_2365 (O_2365,N_19694,N_18673);
nand UO_2366 (O_2366,N_18030,N_19675);
or UO_2367 (O_2367,N_18480,N_19560);
nand UO_2368 (O_2368,N_19511,N_18005);
nand UO_2369 (O_2369,N_18637,N_18377);
xnor UO_2370 (O_2370,N_19597,N_18691);
nor UO_2371 (O_2371,N_19542,N_18664);
nand UO_2372 (O_2372,N_18453,N_19212);
nor UO_2373 (O_2373,N_19177,N_19853);
and UO_2374 (O_2374,N_18649,N_18542);
nor UO_2375 (O_2375,N_19218,N_18911);
xnor UO_2376 (O_2376,N_18906,N_19440);
nor UO_2377 (O_2377,N_19773,N_18966);
nand UO_2378 (O_2378,N_19698,N_18191);
or UO_2379 (O_2379,N_18871,N_18191);
nand UO_2380 (O_2380,N_19493,N_18945);
nor UO_2381 (O_2381,N_18760,N_18312);
xor UO_2382 (O_2382,N_18524,N_18960);
nand UO_2383 (O_2383,N_18434,N_18778);
nand UO_2384 (O_2384,N_18594,N_19291);
and UO_2385 (O_2385,N_19912,N_18229);
or UO_2386 (O_2386,N_18595,N_19677);
or UO_2387 (O_2387,N_18748,N_18493);
xnor UO_2388 (O_2388,N_19773,N_18536);
or UO_2389 (O_2389,N_18478,N_19315);
nand UO_2390 (O_2390,N_18720,N_19094);
nand UO_2391 (O_2391,N_18245,N_18967);
and UO_2392 (O_2392,N_18453,N_19533);
nand UO_2393 (O_2393,N_18412,N_18191);
nor UO_2394 (O_2394,N_19261,N_18624);
nor UO_2395 (O_2395,N_18171,N_19897);
and UO_2396 (O_2396,N_18777,N_18362);
xor UO_2397 (O_2397,N_18007,N_18827);
nand UO_2398 (O_2398,N_19326,N_19809);
or UO_2399 (O_2399,N_19392,N_19670);
xnor UO_2400 (O_2400,N_19270,N_19677);
or UO_2401 (O_2401,N_19093,N_18691);
nor UO_2402 (O_2402,N_18734,N_19175);
nand UO_2403 (O_2403,N_18906,N_19449);
or UO_2404 (O_2404,N_19899,N_18309);
or UO_2405 (O_2405,N_18066,N_18567);
or UO_2406 (O_2406,N_19372,N_19357);
nor UO_2407 (O_2407,N_18840,N_18229);
nand UO_2408 (O_2408,N_18105,N_19906);
and UO_2409 (O_2409,N_19389,N_19706);
nand UO_2410 (O_2410,N_19822,N_19130);
and UO_2411 (O_2411,N_19839,N_19076);
nand UO_2412 (O_2412,N_18074,N_18128);
xor UO_2413 (O_2413,N_19079,N_19131);
and UO_2414 (O_2414,N_19818,N_19497);
or UO_2415 (O_2415,N_19674,N_19853);
nand UO_2416 (O_2416,N_19605,N_19577);
xnor UO_2417 (O_2417,N_19050,N_19617);
xor UO_2418 (O_2418,N_19307,N_19304);
nand UO_2419 (O_2419,N_18755,N_18752);
and UO_2420 (O_2420,N_19267,N_18570);
xnor UO_2421 (O_2421,N_18278,N_18373);
or UO_2422 (O_2422,N_19779,N_18708);
xnor UO_2423 (O_2423,N_19592,N_19212);
xnor UO_2424 (O_2424,N_18592,N_19493);
nor UO_2425 (O_2425,N_19294,N_19001);
or UO_2426 (O_2426,N_19136,N_19015);
xor UO_2427 (O_2427,N_18914,N_18887);
xnor UO_2428 (O_2428,N_18176,N_19433);
or UO_2429 (O_2429,N_19788,N_19772);
and UO_2430 (O_2430,N_19512,N_18364);
nand UO_2431 (O_2431,N_19258,N_19949);
xor UO_2432 (O_2432,N_19691,N_18318);
xor UO_2433 (O_2433,N_18712,N_19168);
or UO_2434 (O_2434,N_19403,N_18834);
or UO_2435 (O_2435,N_18731,N_18840);
nand UO_2436 (O_2436,N_19604,N_19247);
and UO_2437 (O_2437,N_19822,N_19273);
or UO_2438 (O_2438,N_19709,N_18563);
nor UO_2439 (O_2439,N_18064,N_19444);
nor UO_2440 (O_2440,N_19372,N_18354);
nand UO_2441 (O_2441,N_19737,N_19422);
and UO_2442 (O_2442,N_19219,N_18714);
nand UO_2443 (O_2443,N_19528,N_18681);
nor UO_2444 (O_2444,N_19058,N_18763);
nand UO_2445 (O_2445,N_18688,N_18547);
xnor UO_2446 (O_2446,N_19143,N_19651);
or UO_2447 (O_2447,N_19998,N_19766);
xnor UO_2448 (O_2448,N_19289,N_18719);
xnor UO_2449 (O_2449,N_18034,N_19791);
xor UO_2450 (O_2450,N_18101,N_19739);
xor UO_2451 (O_2451,N_19409,N_18705);
xor UO_2452 (O_2452,N_19693,N_18332);
nand UO_2453 (O_2453,N_18518,N_18562);
nor UO_2454 (O_2454,N_19686,N_18451);
xor UO_2455 (O_2455,N_19705,N_18933);
or UO_2456 (O_2456,N_19264,N_18749);
or UO_2457 (O_2457,N_18430,N_19137);
nor UO_2458 (O_2458,N_19592,N_19870);
or UO_2459 (O_2459,N_18001,N_18483);
nand UO_2460 (O_2460,N_18649,N_18363);
or UO_2461 (O_2461,N_19294,N_19100);
xnor UO_2462 (O_2462,N_18158,N_18299);
and UO_2463 (O_2463,N_18008,N_18571);
nor UO_2464 (O_2464,N_19412,N_19592);
or UO_2465 (O_2465,N_18272,N_19416);
or UO_2466 (O_2466,N_18687,N_18352);
nor UO_2467 (O_2467,N_18055,N_19138);
xor UO_2468 (O_2468,N_19171,N_18767);
xnor UO_2469 (O_2469,N_19861,N_18912);
nor UO_2470 (O_2470,N_18675,N_18548);
or UO_2471 (O_2471,N_18357,N_18086);
or UO_2472 (O_2472,N_19113,N_18331);
nand UO_2473 (O_2473,N_18003,N_19300);
nand UO_2474 (O_2474,N_18525,N_19531);
and UO_2475 (O_2475,N_19941,N_18076);
or UO_2476 (O_2476,N_18147,N_18162);
nor UO_2477 (O_2477,N_19264,N_19103);
or UO_2478 (O_2478,N_19726,N_19058);
and UO_2479 (O_2479,N_18677,N_18484);
or UO_2480 (O_2480,N_18135,N_19663);
nor UO_2481 (O_2481,N_18260,N_19967);
or UO_2482 (O_2482,N_18129,N_19133);
and UO_2483 (O_2483,N_18077,N_18378);
xor UO_2484 (O_2484,N_18742,N_18895);
nor UO_2485 (O_2485,N_19693,N_19470);
nand UO_2486 (O_2486,N_18246,N_19286);
or UO_2487 (O_2487,N_19821,N_18148);
nand UO_2488 (O_2488,N_19151,N_18786);
nand UO_2489 (O_2489,N_18810,N_19692);
xnor UO_2490 (O_2490,N_18080,N_19497);
nor UO_2491 (O_2491,N_19162,N_18912);
xor UO_2492 (O_2492,N_19662,N_19036);
or UO_2493 (O_2493,N_19789,N_19717);
nor UO_2494 (O_2494,N_19781,N_19179);
xnor UO_2495 (O_2495,N_18414,N_19084);
or UO_2496 (O_2496,N_18802,N_18457);
nand UO_2497 (O_2497,N_19933,N_19453);
nand UO_2498 (O_2498,N_19910,N_18664);
xnor UO_2499 (O_2499,N_19248,N_18473);
endmodule