module basic_1000_10000_1500_4_levels_1xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nand U0 (N_0,In_323,In_398);
nor U1 (N_1,In_988,In_5);
or U2 (N_2,In_577,In_886);
and U3 (N_3,In_592,In_86);
and U4 (N_4,In_287,In_943);
and U5 (N_5,In_362,In_769);
nor U6 (N_6,In_735,In_609);
nor U7 (N_7,In_834,In_783);
nand U8 (N_8,In_320,In_620);
and U9 (N_9,In_542,In_188);
or U10 (N_10,In_97,In_861);
nand U11 (N_11,In_129,In_731);
and U12 (N_12,In_556,In_419);
or U13 (N_13,In_139,In_972);
nand U14 (N_14,In_543,In_640);
and U15 (N_15,In_215,In_779);
xor U16 (N_16,In_402,In_102);
and U17 (N_17,In_406,In_273);
nor U18 (N_18,In_767,In_182);
and U19 (N_19,In_270,In_278);
and U20 (N_20,In_817,In_751);
nor U21 (N_21,In_246,In_255);
nor U22 (N_22,In_967,In_969);
nor U23 (N_23,In_551,In_451);
nand U24 (N_24,In_448,In_656);
or U25 (N_25,In_688,In_281);
nor U26 (N_26,In_984,In_253);
or U27 (N_27,In_891,In_890);
and U28 (N_28,In_898,In_839);
nor U29 (N_29,In_385,In_47);
nor U30 (N_30,In_96,In_144);
and U31 (N_31,In_141,In_899);
nand U32 (N_32,In_78,In_279);
and U33 (N_33,In_858,In_316);
nor U34 (N_34,In_616,In_617);
and U35 (N_35,In_780,In_503);
and U36 (N_36,In_558,In_622);
nor U37 (N_37,In_582,In_999);
and U38 (N_38,In_480,In_122);
or U39 (N_39,In_686,In_781);
nor U40 (N_40,In_876,In_401);
nand U41 (N_41,In_677,In_304);
nand U42 (N_42,In_681,In_927);
nand U43 (N_43,In_707,In_505);
nor U44 (N_44,In_206,In_605);
or U45 (N_45,In_303,In_319);
nor U46 (N_46,In_459,In_321);
nor U47 (N_47,In_113,In_164);
or U48 (N_48,In_661,In_272);
nand U49 (N_49,In_74,In_189);
nand U50 (N_50,In_805,In_752);
nand U51 (N_51,In_108,In_691);
nand U52 (N_52,In_655,In_233);
or U53 (N_53,In_914,In_717);
and U54 (N_54,In_554,In_470);
and U55 (N_55,In_387,In_361);
nand U56 (N_56,In_719,In_975);
nor U57 (N_57,In_147,In_513);
or U58 (N_58,In_338,In_920);
nand U59 (N_59,In_589,In_520);
nand U60 (N_60,In_350,In_776);
and U61 (N_61,In_159,In_302);
nor U62 (N_62,In_822,In_185);
nand U63 (N_63,In_283,In_940);
nand U64 (N_64,In_375,In_814);
nand U65 (N_65,In_366,In_262);
nand U66 (N_66,In_658,In_296);
nand U67 (N_67,In_700,In_669);
nand U68 (N_68,In_985,In_696);
and U69 (N_69,In_705,In_389);
and U70 (N_70,In_538,In_312);
and U71 (N_71,In_862,In_412);
nor U72 (N_72,In_176,In_469);
nand U73 (N_73,In_257,In_787);
nand U74 (N_74,In_693,In_137);
nor U75 (N_75,In_720,In_405);
and U76 (N_76,In_439,In_824);
and U77 (N_77,In_210,In_831);
or U78 (N_78,In_25,In_732);
and U79 (N_79,In_778,In_794);
and U80 (N_80,In_784,In_836);
nand U81 (N_81,In_235,In_23);
nand U82 (N_82,In_963,In_68);
and U83 (N_83,In_928,In_414);
nor U84 (N_84,In_652,In_601);
nand U85 (N_85,In_293,In_827);
and U86 (N_86,In_841,In_659);
and U87 (N_87,In_379,In_529);
nor U88 (N_88,In_21,In_197);
nand U89 (N_89,In_62,In_76);
or U90 (N_90,In_248,In_26);
or U91 (N_91,In_344,In_602);
or U92 (N_92,In_804,In_260);
nor U93 (N_93,In_367,In_567);
or U94 (N_94,In_675,In_333);
nand U95 (N_95,In_431,In_692);
and U96 (N_96,In_650,In_703);
nand U97 (N_97,In_646,In_351);
nor U98 (N_98,In_791,In_777);
xnor U99 (N_99,In_764,In_536);
nor U100 (N_100,In_423,In_219);
and U101 (N_101,In_107,In_501);
nor U102 (N_102,In_427,In_966);
and U103 (N_103,In_167,In_29);
or U104 (N_104,In_932,In_917);
nor U105 (N_105,In_729,In_924);
nor U106 (N_106,In_586,In_530);
or U107 (N_107,In_823,In_328);
and U108 (N_108,In_936,In_918);
and U109 (N_109,In_873,In_741);
nor U110 (N_110,In_606,In_343);
or U111 (N_111,In_865,In_156);
nand U112 (N_112,In_90,In_243);
nand U113 (N_113,In_926,In_34);
or U114 (N_114,In_464,In_285);
or U115 (N_115,In_789,In_193);
and U116 (N_116,In_992,In_826);
nand U117 (N_117,In_610,In_575);
nand U118 (N_118,In_6,In_840);
or U119 (N_119,In_736,In_438);
nor U120 (N_120,In_178,In_458);
nand U121 (N_121,In_810,In_629);
nand U122 (N_122,In_523,In_549);
xor U123 (N_123,In_88,In_493);
nand U124 (N_124,In_757,In_980);
nor U125 (N_125,In_689,In_157);
nand U126 (N_126,In_591,In_919);
nor U127 (N_127,In_382,In_734);
or U128 (N_128,In_508,In_221);
nand U129 (N_129,In_968,In_702);
nand U130 (N_130,In_54,In_801);
or U131 (N_131,In_881,In_290);
or U132 (N_132,In_668,In_504);
or U133 (N_133,In_939,In_550);
and U134 (N_134,In_1,In_642);
and U135 (N_135,In_748,In_138);
nand U136 (N_136,In_247,In_695);
nand U137 (N_137,In_733,In_258);
or U138 (N_138,In_747,In_983);
nand U139 (N_139,In_244,In_329);
or U140 (N_140,In_368,In_394);
or U141 (N_141,In_45,In_982);
nand U142 (N_142,In_690,In_771);
and U143 (N_143,In_165,In_978);
nor U144 (N_144,In_938,In_208);
or U145 (N_145,In_421,In_973);
or U146 (N_146,In_745,In_326);
nand U147 (N_147,In_65,In_224);
and U148 (N_148,In_654,In_715);
and U149 (N_149,In_704,In_190);
nand U150 (N_150,In_388,In_832);
and U151 (N_151,In_179,In_666);
and U152 (N_152,In_670,In_657);
and U153 (N_153,In_802,In_191);
or U154 (N_154,In_103,In_130);
nand U155 (N_155,In_433,In_492);
nor U156 (N_156,In_941,In_685);
or U157 (N_157,In_237,In_502);
nand U158 (N_158,In_168,In_590);
nand U159 (N_159,In_819,In_879);
or U160 (N_160,In_58,In_949);
xnor U161 (N_161,In_796,In_81);
or U162 (N_162,In_317,In_560);
or U163 (N_163,In_626,In_430);
nor U164 (N_164,In_486,In_718);
nand U165 (N_165,In_305,In_454);
xor U166 (N_166,In_466,In_204);
nor U167 (N_167,In_73,In_393);
or U168 (N_168,In_599,In_94);
or U169 (N_169,In_331,In_568);
or U170 (N_170,In_516,In_99);
or U171 (N_171,In_183,In_298);
or U172 (N_172,In_825,In_623);
nor U173 (N_173,In_953,In_479);
nand U174 (N_174,In_201,In_628);
nor U175 (N_175,In_739,In_607);
nand U176 (N_176,In_223,In_7);
or U177 (N_177,In_209,In_476);
nand U178 (N_178,In_674,In_227);
nand U179 (N_179,In_291,In_14);
or U180 (N_180,In_484,In_989);
or U181 (N_181,In_61,In_32);
nand U182 (N_182,In_821,In_300);
nor U183 (N_183,In_284,In_813);
nor U184 (N_184,In_267,In_820);
or U185 (N_185,In_254,In_756);
or U186 (N_186,In_797,In_318);
nor U187 (N_187,In_85,In_104);
nor U188 (N_188,In_684,In_462);
and U189 (N_189,In_613,In_136);
nor U190 (N_190,In_962,In_251);
nor U191 (N_191,In_403,In_916);
nand U192 (N_192,In_954,In_649);
nor U193 (N_193,In_994,In_709);
nand U194 (N_194,In_539,In_935);
nor U195 (N_195,In_811,In_816);
nand U196 (N_196,In_497,In_866);
nand U197 (N_197,In_915,In_860);
or U198 (N_198,In_410,In_473);
and U199 (N_199,In_180,In_19);
nand U200 (N_200,In_990,In_611);
or U201 (N_201,In_614,In_250);
or U202 (N_202,In_397,In_175);
nor U203 (N_203,In_639,In_63);
nand U204 (N_204,In_425,In_378);
nor U205 (N_205,In_441,In_728);
or U206 (N_206,In_0,In_697);
and U207 (N_207,In_564,In_521);
and U208 (N_208,In_971,In_905);
or U209 (N_209,In_212,In_460);
xnor U210 (N_210,In_222,In_913);
nor U211 (N_211,In_488,In_581);
or U212 (N_212,In_349,In_481);
and U213 (N_213,In_597,In_958);
xor U214 (N_214,In_286,In_311);
nor U215 (N_215,In_461,In_447);
and U216 (N_216,In_584,In_566);
and U217 (N_217,In_146,In_637);
nor U218 (N_218,In_143,In_651);
nand U219 (N_219,In_337,In_2);
and U220 (N_220,In_773,In_901);
and U221 (N_221,In_496,In_517);
and U222 (N_222,In_772,In_280);
nand U223 (N_223,In_569,In_548);
and U224 (N_224,In_765,In_242);
or U225 (N_225,In_509,In_452);
or U226 (N_226,In_274,In_422);
or U227 (N_227,In_843,In_432);
nand U228 (N_228,In_960,In_396);
and U229 (N_229,In_562,In_721);
or U230 (N_230,In_116,In_112);
nor U231 (N_231,In_526,In_544);
nand U232 (N_232,In_815,In_489);
or U233 (N_233,In_155,In_522);
and U234 (N_234,In_869,In_580);
and U235 (N_235,In_140,In_578);
nand U236 (N_236,In_987,In_663);
nor U237 (N_237,In_51,In_877);
nor U238 (N_238,In_514,In_234);
nand U239 (N_239,In_959,In_648);
and U240 (N_240,In_341,In_373);
or U241 (N_241,In_231,In_854);
nor U242 (N_242,In_946,In_912);
and U243 (N_243,In_332,In_166);
and U244 (N_244,In_31,In_956);
or U245 (N_245,In_33,In_534);
and U246 (N_246,In_67,In_12);
and U247 (N_247,In_662,In_131);
and U248 (N_248,In_878,In_744);
nand U249 (N_249,In_892,In_216);
or U250 (N_250,In_803,In_428);
and U251 (N_251,In_603,In_339);
and U252 (N_252,In_485,In_135);
nand U253 (N_253,In_371,In_335);
and U254 (N_254,In_618,In_519);
or U255 (N_255,In_105,In_615);
or U256 (N_256,In_173,In_181);
and U257 (N_257,In_923,In_118);
and U258 (N_258,In_738,In_408);
nand U259 (N_259,In_314,In_903);
nand U260 (N_260,In_199,In_565);
and U261 (N_261,In_202,In_245);
and U262 (N_262,In_882,In_383);
and U263 (N_263,In_906,In_585);
and U264 (N_264,In_524,In_844);
or U265 (N_265,In_798,In_330);
nand U266 (N_266,In_357,In_295);
xnor U267 (N_267,In_993,In_859);
or U268 (N_268,In_334,In_698);
or U269 (N_269,In_354,In_760);
nand U270 (N_270,In_997,In_996);
and U271 (N_271,In_856,In_4);
nor U272 (N_272,In_55,In_874);
and U273 (N_273,In_345,In_894);
and U274 (N_274,In_535,In_482);
nand U275 (N_275,In_364,In_92);
and U276 (N_276,In_644,In_265);
or U277 (N_277,In_353,In_845);
nor U278 (N_278,In_145,In_604);
or U279 (N_279,In_490,In_456);
and U280 (N_280,In_790,In_16);
nor U281 (N_281,In_676,In_848);
and U282 (N_282,In_352,In_424);
and U283 (N_283,In_301,In_386);
and U284 (N_284,In_249,In_214);
or U285 (N_285,In_277,In_200);
and U286 (N_286,In_647,In_977);
and U287 (N_287,In_171,In_902);
and U288 (N_288,In_818,In_380);
or U289 (N_289,In_151,In_714);
nand U290 (N_290,In_125,In_974);
nand U291 (N_291,In_170,In_477);
nor U292 (N_292,In_163,In_627);
nor U293 (N_293,In_785,In_995);
nor U294 (N_294,In_788,In_115);
and U295 (N_295,In_36,In_437);
nand U296 (N_296,In_268,In_225);
nand U297 (N_297,In_392,In_89);
nand U298 (N_298,In_643,In_863);
or U299 (N_299,In_263,In_411);
and U300 (N_300,In_8,In_327);
or U301 (N_301,In_404,In_358);
nand U302 (N_302,In_724,In_399);
or U303 (N_303,In_109,In_533);
nor U304 (N_304,In_18,In_236);
nor U305 (N_305,In_812,In_619);
nor U306 (N_306,In_981,In_429);
and U307 (N_307,In_722,In_857);
nand U308 (N_308,In_294,In_893);
and U309 (N_309,In_871,In_495);
or U310 (N_310,In_415,In_678);
nand U311 (N_311,In_758,In_537);
nor U312 (N_312,In_518,In_56);
nor U313 (N_313,In_727,In_596);
nor U314 (N_314,In_541,In_100);
or U315 (N_315,In_395,In_557);
and U316 (N_316,In_483,In_52);
nor U317 (N_317,In_576,In_699);
nor U318 (N_318,In_908,In_570);
and U319 (N_319,In_413,In_515);
or U320 (N_320,In_712,In_474);
and U321 (N_321,In_683,In_774);
and U322 (N_322,In_252,In_309);
or U323 (N_323,In_842,In_838);
and U324 (N_324,In_49,In_187);
nand U325 (N_325,In_75,In_443);
nor U326 (N_326,In_71,In_241);
and U327 (N_327,In_883,In_407);
nor U328 (N_328,In_846,In_297);
xor U329 (N_329,In_500,In_494);
nand U330 (N_330,In_746,In_851);
or U331 (N_331,In_952,In_673);
nor U332 (N_332,In_239,In_847);
nand U333 (N_333,In_763,In_348);
nand U334 (N_334,In_929,In_192);
xor U335 (N_335,In_240,In_306);
and U336 (N_336,In_3,In_540);
or U337 (N_337,In_121,In_900);
nand U338 (N_338,In_340,In_48);
or U339 (N_339,In_28,In_740);
nand U340 (N_340,In_755,In_148);
nor U341 (N_341,In_964,In_679);
or U342 (N_342,In_895,In_664);
nor U343 (N_343,In_372,In_743);
nand U344 (N_344,In_446,In_829);
nand U345 (N_345,In_608,In_95);
and U346 (N_346,In_682,In_853);
or U347 (N_347,In_359,In_587);
or U348 (N_348,In_633,In_849);
or U349 (N_349,In_934,In_672);
or U350 (N_350,In_313,In_83);
nor U351 (N_351,In_128,In_991);
nor U352 (N_352,In_194,In_630);
and U353 (N_353,In_979,In_119);
nand U354 (N_354,In_635,In_24);
nor U355 (N_355,In_976,In_792);
nor U356 (N_356,In_87,In_44);
and U357 (N_357,In_716,In_855);
nor U358 (N_358,In_594,In_416);
or U359 (N_359,In_324,In_299);
nand U360 (N_360,In_117,In_336);
or U361 (N_361,In_806,In_282);
xnor U362 (N_362,In_573,In_571);
or U363 (N_363,In_711,In_742);
or U364 (N_364,In_725,In_226);
and U365 (N_365,In_218,In_275);
nor U366 (N_366,In_833,In_381);
nand U367 (N_367,In_561,In_835);
nor U368 (N_368,In_713,In_922);
nor U369 (N_369,In_64,In_205);
nor U370 (N_370,In_641,In_98);
nor U371 (N_371,In_754,In_525);
and U372 (N_372,In_17,In_292);
nand U373 (N_373,In_203,In_793);
or U374 (N_374,In_213,In_123);
and U375 (N_375,In_376,In_708);
and U376 (N_376,In_911,In_434);
or U377 (N_377,In_872,In_101);
nor U378 (N_378,In_595,In_868);
or U379 (N_379,In_445,In_761);
nand U380 (N_380,In_307,In_355);
or U381 (N_381,In_435,In_921);
nor U382 (N_382,In_468,In_638);
or U383 (N_383,In_775,In_888);
nand U384 (N_384,In_471,In_261);
and U385 (N_385,In_198,In_77);
nand U386 (N_386,In_256,In_726);
nand U387 (N_387,In_807,In_782);
and U388 (N_388,In_84,In_134);
nor U389 (N_389,In_632,In_232);
nand U390 (N_390,In_162,In_950);
nand U391 (N_391,In_79,In_126);
nor U392 (N_392,In_120,In_152);
or U393 (N_393,In_910,In_114);
nand U394 (N_394,In_887,In_830);
nand U395 (N_395,In_217,In_467);
or U396 (N_396,In_532,In_799);
and U397 (N_397,In_370,In_510);
or U398 (N_398,In_37,In_27);
and U399 (N_399,In_694,In_93);
nand U400 (N_400,In_211,In_947);
and U401 (N_401,In_172,In_528);
nor U402 (N_402,In_264,In_390);
nor U403 (N_403,In_965,In_885);
and U404 (N_404,In_491,In_653);
and U405 (N_405,In_444,In_706);
and U406 (N_406,In_583,In_15);
nor U407 (N_407,In_82,In_961);
or U408 (N_408,In_195,In_259);
and U409 (N_409,In_72,In_749);
or U410 (N_410,In_50,In_955);
or U411 (N_411,In_600,In_322);
nor U412 (N_412,In_527,In_625);
nand U413 (N_413,In_455,In_356);
or U414 (N_414,In_110,In_342);
and U415 (N_415,In_70,In_153);
nor U416 (N_416,In_436,In_759);
nand U417 (N_417,In_38,In_230);
nor U418 (N_418,In_942,In_269);
nand U419 (N_419,In_636,In_420);
and U420 (N_420,In_10,In_154);
and U421 (N_421,In_150,In_409);
or U422 (N_422,In_475,In_347);
nand U423 (N_423,In_453,In_426);
or U424 (N_424,In_660,In_160);
nand U425 (N_425,In_907,In_91);
and U426 (N_426,In_680,In_465);
and U427 (N_427,In_808,In_60);
and U428 (N_428,In_365,In_933);
nor U429 (N_429,In_572,In_391);
or U430 (N_430,In_800,In_127);
nor U431 (N_431,In_850,In_621);
nand U432 (N_432,In_369,In_80);
and U433 (N_433,In_238,In_864);
and U434 (N_434,In_795,In_889);
and U435 (N_435,In_870,In_310);
and U436 (N_436,In_43,In_579);
nor U437 (N_437,In_867,In_184);
nand U438 (N_438,In_762,In_400);
nor U439 (N_439,In_487,In_266);
nand U440 (N_440,In_809,In_645);
or U441 (N_441,In_512,In_897);
nor U442 (N_442,In_308,In_612);
nand U443 (N_443,In_545,In_884);
nand U444 (N_444,In_418,In_142);
nor U445 (N_445,In_970,In_315);
or U446 (N_446,In_132,In_40);
nand U447 (N_447,In_289,In_106);
nand U448 (N_448,In_472,In_149);
nand U449 (N_449,In_9,In_687);
and U450 (N_450,In_768,In_770);
nor U451 (N_451,In_701,In_229);
or U452 (N_452,In_730,In_417);
and U453 (N_453,In_440,In_925);
or U454 (N_454,In_753,In_133);
and U455 (N_455,In_559,In_880);
nor U456 (N_456,In_384,In_111);
nand U457 (N_457,In_547,In_174);
or U458 (N_458,In_377,In_931);
nand U459 (N_459,In_463,In_998);
nor U460 (N_460,In_325,In_66);
nand U461 (N_461,In_220,In_634);
nor U462 (N_462,In_531,In_41);
nand U463 (N_463,In_948,In_786);
and U464 (N_464,In_896,In_13);
nand U465 (N_465,In_750,In_507);
and U466 (N_466,In_161,In_563);
nor U467 (N_467,In_723,In_186);
nor U468 (N_468,In_546,In_671);
nand U469 (N_469,In_937,In_42);
or U470 (N_470,In_957,In_574);
and U471 (N_471,In_930,In_598);
nand U472 (N_472,In_498,In_631);
nor U473 (N_473,In_442,In_20);
or U474 (N_474,In_506,In_499);
nand U475 (N_475,In_553,In_35);
nand U476 (N_476,In_588,In_710);
and U477 (N_477,In_986,In_449);
xor U478 (N_478,In_457,In_22);
or U479 (N_479,In_363,In_69);
nor U480 (N_480,In_30,In_904);
and U481 (N_481,In_511,In_228);
and U482 (N_482,In_478,In_593);
or U483 (N_483,In_59,In_39);
nand U484 (N_484,In_945,In_450);
and U485 (N_485,In_169,In_552);
nand U486 (N_486,In_667,In_124);
and U487 (N_487,In_46,In_276);
nor U488 (N_488,In_875,In_737);
and U489 (N_489,In_207,In_346);
nand U490 (N_490,In_57,In_909);
nand U491 (N_491,In_360,In_944);
or U492 (N_492,In_177,In_288);
nor U493 (N_493,In_624,In_951);
or U494 (N_494,In_852,In_196);
or U495 (N_495,In_53,In_665);
nand U496 (N_496,In_374,In_766);
and U497 (N_497,In_828,In_271);
and U498 (N_498,In_158,In_11);
nand U499 (N_499,In_555,In_837);
nor U500 (N_500,In_251,In_159);
or U501 (N_501,In_333,In_516);
nand U502 (N_502,In_926,In_703);
nand U503 (N_503,In_297,In_499);
nor U504 (N_504,In_461,In_730);
nand U505 (N_505,In_924,In_985);
and U506 (N_506,In_223,In_982);
nand U507 (N_507,In_116,In_144);
nor U508 (N_508,In_716,In_199);
nor U509 (N_509,In_93,In_607);
nor U510 (N_510,In_919,In_832);
nor U511 (N_511,In_234,In_331);
or U512 (N_512,In_850,In_359);
nand U513 (N_513,In_813,In_285);
nor U514 (N_514,In_769,In_265);
nand U515 (N_515,In_738,In_494);
nand U516 (N_516,In_996,In_910);
nand U517 (N_517,In_594,In_312);
or U518 (N_518,In_107,In_95);
or U519 (N_519,In_133,In_946);
and U520 (N_520,In_686,In_637);
and U521 (N_521,In_623,In_454);
nand U522 (N_522,In_954,In_938);
and U523 (N_523,In_983,In_584);
and U524 (N_524,In_710,In_592);
nor U525 (N_525,In_792,In_35);
or U526 (N_526,In_960,In_253);
nor U527 (N_527,In_646,In_761);
nand U528 (N_528,In_419,In_646);
nand U529 (N_529,In_720,In_363);
nand U530 (N_530,In_647,In_771);
and U531 (N_531,In_199,In_182);
and U532 (N_532,In_895,In_870);
and U533 (N_533,In_206,In_169);
and U534 (N_534,In_640,In_191);
and U535 (N_535,In_811,In_883);
nor U536 (N_536,In_166,In_543);
nor U537 (N_537,In_782,In_350);
and U538 (N_538,In_169,In_73);
and U539 (N_539,In_541,In_552);
and U540 (N_540,In_967,In_232);
and U541 (N_541,In_881,In_694);
nor U542 (N_542,In_223,In_297);
nand U543 (N_543,In_516,In_421);
nand U544 (N_544,In_180,In_188);
or U545 (N_545,In_839,In_694);
or U546 (N_546,In_657,In_912);
nor U547 (N_547,In_284,In_927);
and U548 (N_548,In_617,In_149);
and U549 (N_549,In_365,In_767);
or U550 (N_550,In_56,In_111);
nand U551 (N_551,In_942,In_319);
nand U552 (N_552,In_123,In_53);
nor U553 (N_553,In_34,In_311);
and U554 (N_554,In_184,In_570);
nor U555 (N_555,In_914,In_972);
and U556 (N_556,In_104,In_818);
or U557 (N_557,In_38,In_741);
nand U558 (N_558,In_830,In_714);
or U559 (N_559,In_360,In_841);
and U560 (N_560,In_402,In_969);
nand U561 (N_561,In_407,In_352);
nand U562 (N_562,In_689,In_382);
nor U563 (N_563,In_748,In_511);
or U564 (N_564,In_327,In_301);
and U565 (N_565,In_271,In_640);
nand U566 (N_566,In_742,In_581);
or U567 (N_567,In_452,In_996);
or U568 (N_568,In_592,In_948);
nor U569 (N_569,In_509,In_374);
nor U570 (N_570,In_254,In_666);
nor U571 (N_571,In_337,In_909);
nor U572 (N_572,In_803,In_960);
nand U573 (N_573,In_159,In_643);
and U574 (N_574,In_33,In_651);
or U575 (N_575,In_55,In_243);
and U576 (N_576,In_787,In_266);
and U577 (N_577,In_709,In_342);
nand U578 (N_578,In_377,In_360);
nor U579 (N_579,In_492,In_278);
and U580 (N_580,In_614,In_437);
nor U581 (N_581,In_359,In_390);
and U582 (N_582,In_838,In_465);
nand U583 (N_583,In_432,In_235);
xor U584 (N_584,In_864,In_279);
nand U585 (N_585,In_684,In_797);
nand U586 (N_586,In_438,In_333);
and U587 (N_587,In_730,In_989);
nor U588 (N_588,In_638,In_499);
nor U589 (N_589,In_803,In_104);
or U590 (N_590,In_971,In_74);
nor U591 (N_591,In_498,In_995);
nand U592 (N_592,In_118,In_320);
nand U593 (N_593,In_660,In_410);
or U594 (N_594,In_47,In_892);
nand U595 (N_595,In_784,In_991);
or U596 (N_596,In_348,In_737);
nand U597 (N_597,In_785,In_934);
nor U598 (N_598,In_287,In_848);
or U599 (N_599,In_187,In_634);
and U600 (N_600,In_512,In_167);
nor U601 (N_601,In_52,In_949);
or U602 (N_602,In_511,In_731);
nand U603 (N_603,In_801,In_690);
or U604 (N_604,In_537,In_218);
and U605 (N_605,In_802,In_819);
nand U606 (N_606,In_204,In_279);
nand U607 (N_607,In_126,In_469);
or U608 (N_608,In_968,In_363);
or U609 (N_609,In_929,In_507);
and U610 (N_610,In_69,In_308);
nor U611 (N_611,In_956,In_305);
nand U612 (N_612,In_309,In_941);
and U613 (N_613,In_704,In_756);
and U614 (N_614,In_824,In_534);
or U615 (N_615,In_822,In_79);
nor U616 (N_616,In_33,In_171);
xor U617 (N_617,In_103,In_77);
or U618 (N_618,In_905,In_694);
or U619 (N_619,In_102,In_300);
and U620 (N_620,In_652,In_231);
nor U621 (N_621,In_765,In_376);
nor U622 (N_622,In_314,In_590);
nor U623 (N_623,In_628,In_743);
nand U624 (N_624,In_578,In_274);
and U625 (N_625,In_354,In_360);
nor U626 (N_626,In_449,In_946);
and U627 (N_627,In_692,In_819);
nor U628 (N_628,In_992,In_572);
nor U629 (N_629,In_909,In_310);
nor U630 (N_630,In_50,In_579);
nand U631 (N_631,In_660,In_827);
nor U632 (N_632,In_257,In_357);
or U633 (N_633,In_731,In_476);
nand U634 (N_634,In_661,In_866);
or U635 (N_635,In_804,In_389);
or U636 (N_636,In_539,In_60);
or U637 (N_637,In_162,In_960);
or U638 (N_638,In_564,In_835);
nor U639 (N_639,In_81,In_591);
and U640 (N_640,In_432,In_784);
nand U641 (N_641,In_544,In_460);
or U642 (N_642,In_855,In_913);
nor U643 (N_643,In_321,In_1);
nand U644 (N_644,In_531,In_418);
nor U645 (N_645,In_229,In_718);
nand U646 (N_646,In_930,In_905);
and U647 (N_647,In_906,In_655);
or U648 (N_648,In_745,In_146);
nor U649 (N_649,In_534,In_357);
nand U650 (N_650,In_645,In_245);
nand U651 (N_651,In_286,In_321);
nand U652 (N_652,In_195,In_524);
and U653 (N_653,In_708,In_609);
and U654 (N_654,In_676,In_744);
nand U655 (N_655,In_776,In_665);
nand U656 (N_656,In_305,In_378);
nand U657 (N_657,In_365,In_299);
or U658 (N_658,In_874,In_313);
or U659 (N_659,In_982,In_730);
and U660 (N_660,In_621,In_10);
or U661 (N_661,In_929,In_985);
or U662 (N_662,In_78,In_224);
nor U663 (N_663,In_56,In_938);
or U664 (N_664,In_261,In_795);
or U665 (N_665,In_902,In_220);
and U666 (N_666,In_376,In_579);
nor U667 (N_667,In_765,In_936);
or U668 (N_668,In_60,In_923);
nor U669 (N_669,In_281,In_272);
nand U670 (N_670,In_491,In_304);
nor U671 (N_671,In_713,In_174);
and U672 (N_672,In_396,In_733);
and U673 (N_673,In_726,In_849);
nor U674 (N_674,In_225,In_143);
and U675 (N_675,In_195,In_858);
and U676 (N_676,In_710,In_272);
nor U677 (N_677,In_769,In_363);
and U678 (N_678,In_664,In_879);
nand U679 (N_679,In_858,In_45);
or U680 (N_680,In_443,In_989);
and U681 (N_681,In_325,In_734);
nor U682 (N_682,In_997,In_646);
and U683 (N_683,In_17,In_111);
and U684 (N_684,In_861,In_370);
nor U685 (N_685,In_14,In_672);
and U686 (N_686,In_599,In_26);
nor U687 (N_687,In_530,In_171);
nor U688 (N_688,In_631,In_533);
nand U689 (N_689,In_972,In_639);
nor U690 (N_690,In_282,In_458);
nor U691 (N_691,In_954,In_377);
or U692 (N_692,In_395,In_531);
nor U693 (N_693,In_783,In_265);
nand U694 (N_694,In_983,In_353);
or U695 (N_695,In_101,In_623);
or U696 (N_696,In_687,In_371);
nor U697 (N_697,In_857,In_507);
or U698 (N_698,In_151,In_775);
and U699 (N_699,In_691,In_789);
nor U700 (N_700,In_777,In_42);
and U701 (N_701,In_575,In_671);
and U702 (N_702,In_838,In_258);
or U703 (N_703,In_145,In_556);
or U704 (N_704,In_255,In_459);
or U705 (N_705,In_344,In_65);
nand U706 (N_706,In_827,In_519);
nor U707 (N_707,In_31,In_435);
nor U708 (N_708,In_739,In_672);
or U709 (N_709,In_211,In_763);
and U710 (N_710,In_286,In_791);
nor U711 (N_711,In_538,In_316);
nor U712 (N_712,In_233,In_789);
nor U713 (N_713,In_779,In_716);
nor U714 (N_714,In_576,In_849);
and U715 (N_715,In_156,In_365);
and U716 (N_716,In_105,In_586);
or U717 (N_717,In_153,In_750);
and U718 (N_718,In_605,In_805);
or U719 (N_719,In_380,In_544);
and U720 (N_720,In_497,In_444);
and U721 (N_721,In_961,In_260);
nand U722 (N_722,In_545,In_704);
nand U723 (N_723,In_826,In_428);
and U724 (N_724,In_379,In_879);
and U725 (N_725,In_761,In_199);
nor U726 (N_726,In_754,In_349);
nor U727 (N_727,In_939,In_420);
and U728 (N_728,In_615,In_837);
or U729 (N_729,In_204,In_514);
and U730 (N_730,In_496,In_633);
and U731 (N_731,In_506,In_565);
nor U732 (N_732,In_582,In_937);
nor U733 (N_733,In_851,In_410);
and U734 (N_734,In_429,In_556);
nor U735 (N_735,In_96,In_463);
or U736 (N_736,In_305,In_968);
or U737 (N_737,In_322,In_75);
or U738 (N_738,In_545,In_342);
and U739 (N_739,In_58,In_48);
and U740 (N_740,In_767,In_179);
nand U741 (N_741,In_773,In_555);
or U742 (N_742,In_752,In_145);
and U743 (N_743,In_353,In_267);
nand U744 (N_744,In_459,In_472);
and U745 (N_745,In_827,In_381);
nand U746 (N_746,In_855,In_45);
and U747 (N_747,In_793,In_34);
nor U748 (N_748,In_948,In_792);
nand U749 (N_749,In_116,In_367);
and U750 (N_750,In_288,In_374);
and U751 (N_751,In_891,In_518);
nor U752 (N_752,In_266,In_809);
nand U753 (N_753,In_156,In_782);
and U754 (N_754,In_925,In_729);
or U755 (N_755,In_475,In_90);
or U756 (N_756,In_922,In_665);
and U757 (N_757,In_485,In_274);
xnor U758 (N_758,In_567,In_550);
nand U759 (N_759,In_127,In_721);
nand U760 (N_760,In_258,In_37);
or U761 (N_761,In_327,In_926);
nor U762 (N_762,In_199,In_542);
nor U763 (N_763,In_206,In_894);
and U764 (N_764,In_814,In_408);
or U765 (N_765,In_748,In_49);
nor U766 (N_766,In_619,In_805);
or U767 (N_767,In_3,In_36);
or U768 (N_768,In_399,In_600);
xor U769 (N_769,In_57,In_552);
nand U770 (N_770,In_917,In_870);
and U771 (N_771,In_283,In_218);
and U772 (N_772,In_581,In_995);
nor U773 (N_773,In_171,In_775);
or U774 (N_774,In_163,In_21);
and U775 (N_775,In_441,In_679);
and U776 (N_776,In_260,In_330);
nand U777 (N_777,In_596,In_427);
nand U778 (N_778,In_779,In_704);
nor U779 (N_779,In_817,In_966);
nand U780 (N_780,In_649,In_651);
nor U781 (N_781,In_594,In_507);
and U782 (N_782,In_108,In_939);
or U783 (N_783,In_176,In_173);
nor U784 (N_784,In_200,In_971);
or U785 (N_785,In_47,In_519);
nand U786 (N_786,In_35,In_195);
nand U787 (N_787,In_605,In_792);
and U788 (N_788,In_6,In_558);
nand U789 (N_789,In_666,In_37);
nand U790 (N_790,In_653,In_80);
nand U791 (N_791,In_934,In_783);
nand U792 (N_792,In_315,In_527);
and U793 (N_793,In_571,In_459);
or U794 (N_794,In_775,In_208);
nand U795 (N_795,In_631,In_662);
or U796 (N_796,In_385,In_500);
nor U797 (N_797,In_49,In_878);
nor U798 (N_798,In_857,In_435);
or U799 (N_799,In_465,In_295);
xor U800 (N_800,In_846,In_649);
nand U801 (N_801,In_654,In_596);
or U802 (N_802,In_496,In_42);
nor U803 (N_803,In_182,In_679);
or U804 (N_804,In_287,In_695);
nand U805 (N_805,In_293,In_775);
nor U806 (N_806,In_566,In_469);
or U807 (N_807,In_7,In_22);
or U808 (N_808,In_53,In_867);
nand U809 (N_809,In_285,In_956);
and U810 (N_810,In_266,In_642);
or U811 (N_811,In_29,In_536);
and U812 (N_812,In_739,In_975);
nand U813 (N_813,In_198,In_838);
nand U814 (N_814,In_871,In_9);
and U815 (N_815,In_943,In_19);
nand U816 (N_816,In_733,In_966);
nand U817 (N_817,In_644,In_710);
xor U818 (N_818,In_755,In_646);
or U819 (N_819,In_101,In_72);
nand U820 (N_820,In_66,In_138);
and U821 (N_821,In_852,In_587);
nor U822 (N_822,In_897,In_539);
or U823 (N_823,In_909,In_287);
and U824 (N_824,In_162,In_315);
nand U825 (N_825,In_88,In_181);
nor U826 (N_826,In_273,In_390);
or U827 (N_827,In_467,In_594);
nor U828 (N_828,In_398,In_244);
nor U829 (N_829,In_932,In_625);
nand U830 (N_830,In_318,In_993);
and U831 (N_831,In_124,In_473);
nand U832 (N_832,In_955,In_846);
nor U833 (N_833,In_445,In_195);
nor U834 (N_834,In_788,In_328);
nand U835 (N_835,In_8,In_390);
nand U836 (N_836,In_769,In_160);
nor U837 (N_837,In_871,In_419);
nand U838 (N_838,In_296,In_33);
nor U839 (N_839,In_538,In_423);
and U840 (N_840,In_122,In_762);
nor U841 (N_841,In_530,In_798);
nand U842 (N_842,In_125,In_257);
or U843 (N_843,In_603,In_541);
xor U844 (N_844,In_320,In_314);
and U845 (N_845,In_412,In_645);
nand U846 (N_846,In_712,In_709);
or U847 (N_847,In_669,In_743);
and U848 (N_848,In_502,In_893);
or U849 (N_849,In_489,In_635);
or U850 (N_850,In_460,In_702);
and U851 (N_851,In_121,In_910);
nor U852 (N_852,In_706,In_879);
nand U853 (N_853,In_948,In_563);
nand U854 (N_854,In_828,In_514);
nand U855 (N_855,In_274,In_923);
nor U856 (N_856,In_849,In_905);
and U857 (N_857,In_362,In_316);
nor U858 (N_858,In_789,In_34);
and U859 (N_859,In_62,In_603);
or U860 (N_860,In_126,In_184);
or U861 (N_861,In_153,In_315);
or U862 (N_862,In_922,In_81);
and U863 (N_863,In_71,In_332);
and U864 (N_864,In_940,In_373);
or U865 (N_865,In_472,In_950);
nand U866 (N_866,In_260,In_721);
nand U867 (N_867,In_468,In_699);
nor U868 (N_868,In_643,In_191);
and U869 (N_869,In_172,In_289);
and U870 (N_870,In_887,In_771);
or U871 (N_871,In_946,In_922);
and U872 (N_872,In_248,In_710);
and U873 (N_873,In_883,In_765);
and U874 (N_874,In_467,In_244);
or U875 (N_875,In_166,In_865);
and U876 (N_876,In_784,In_207);
or U877 (N_877,In_198,In_188);
nand U878 (N_878,In_742,In_321);
and U879 (N_879,In_610,In_45);
nor U880 (N_880,In_146,In_206);
or U881 (N_881,In_985,In_317);
nand U882 (N_882,In_381,In_318);
nand U883 (N_883,In_239,In_882);
nand U884 (N_884,In_350,In_195);
xnor U885 (N_885,In_794,In_306);
and U886 (N_886,In_180,In_586);
nor U887 (N_887,In_423,In_665);
and U888 (N_888,In_711,In_378);
or U889 (N_889,In_893,In_398);
or U890 (N_890,In_408,In_892);
nor U891 (N_891,In_252,In_666);
nor U892 (N_892,In_921,In_150);
nand U893 (N_893,In_563,In_391);
or U894 (N_894,In_817,In_727);
and U895 (N_895,In_167,In_111);
and U896 (N_896,In_487,In_544);
or U897 (N_897,In_415,In_187);
or U898 (N_898,In_805,In_670);
nor U899 (N_899,In_567,In_767);
nor U900 (N_900,In_318,In_199);
and U901 (N_901,In_473,In_161);
nor U902 (N_902,In_42,In_389);
nor U903 (N_903,In_33,In_786);
and U904 (N_904,In_813,In_291);
or U905 (N_905,In_97,In_390);
or U906 (N_906,In_591,In_183);
nor U907 (N_907,In_737,In_503);
nor U908 (N_908,In_294,In_122);
nor U909 (N_909,In_62,In_725);
and U910 (N_910,In_995,In_306);
nand U911 (N_911,In_518,In_339);
and U912 (N_912,In_703,In_450);
nor U913 (N_913,In_168,In_959);
and U914 (N_914,In_443,In_981);
nand U915 (N_915,In_818,In_381);
nand U916 (N_916,In_478,In_5);
or U917 (N_917,In_918,In_845);
or U918 (N_918,In_536,In_477);
or U919 (N_919,In_133,In_403);
xnor U920 (N_920,In_916,In_513);
and U921 (N_921,In_757,In_31);
nand U922 (N_922,In_167,In_804);
nand U923 (N_923,In_209,In_859);
or U924 (N_924,In_973,In_180);
nor U925 (N_925,In_514,In_850);
xnor U926 (N_926,In_397,In_781);
and U927 (N_927,In_909,In_582);
and U928 (N_928,In_584,In_875);
nand U929 (N_929,In_694,In_980);
nor U930 (N_930,In_593,In_136);
nand U931 (N_931,In_81,In_336);
and U932 (N_932,In_506,In_302);
nand U933 (N_933,In_126,In_187);
and U934 (N_934,In_176,In_590);
nor U935 (N_935,In_499,In_892);
or U936 (N_936,In_962,In_330);
or U937 (N_937,In_693,In_789);
and U938 (N_938,In_61,In_797);
nand U939 (N_939,In_204,In_209);
or U940 (N_940,In_785,In_713);
nor U941 (N_941,In_485,In_708);
nand U942 (N_942,In_231,In_364);
and U943 (N_943,In_524,In_527);
or U944 (N_944,In_520,In_438);
and U945 (N_945,In_765,In_654);
and U946 (N_946,In_38,In_142);
nor U947 (N_947,In_487,In_751);
nor U948 (N_948,In_600,In_17);
and U949 (N_949,In_266,In_212);
and U950 (N_950,In_252,In_651);
and U951 (N_951,In_468,In_819);
nand U952 (N_952,In_397,In_34);
nand U953 (N_953,In_449,In_67);
nor U954 (N_954,In_605,In_878);
or U955 (N_955,In_181,In_499);
and U956 (N_956,In_625,In_729);
nor U957 (N_957,In_788,In_815);
nand U958 (N_958,In_420,In_934);
nor U959 (N_959,In_796,In_664);
nand U960 (N_960,In_539,In_943);
nand U961 (N_961,In_827,In_377);
or U962 (N_962,In_251,In_493);
nand U963 (N_963,In_574,In_650);
or U964 (N_964,In_165,In_907);
nor U965 (N_965,In_704,In_270);
and U966 (N_966,In_21,In_645);
nor U967 (N_967,In_57,In_464);
nand U968 (N_968,In_388,In_855);
nand U969 (N_969,In_454,In_763);
nor U970 (N_970,In_790,In_40);
and U971 (N_971,In_943,In_824);
and U972 (N_972,In_361,In_314);
nor U973 (N_973,In_767,In_896);
and U974 (N_974,In_123,In_202);
or U975 (N_975,In_575,In_582);
and U976 (N_976,In_495,In_258);
nor U977 (N_977,In_19,In_685);
nand U978 (N_978,In_702,In_144);
and U979 (N_979,In_211,In_876);
nand U980 (N_980,In_721,In_219);
or U981 (N_981,In_778,In_416);
or U982 (N_982,In_651,In_486);
or U983 (N_983,In_911,In_622);
or U984 (N_984,In_248,In_247);
nand U985 (N_985,In_842,In_583);
nor U986 (N_986,In_99,In_374);
nand U987 (N_987,In_269,In_216);
nor U988 (N_988,In_94,In_485);
nor U989 (N_989,In_620,In_542);
or U990 (N_990,In_569,In_502);
nand U991 (N_991,In_243,In_697);
and U992 (N_992,In_871,In_320);
or U993 (N_993,In_571,In_575);
nor U994 (N_994,In_460,In_248);
or U995 (N_995,In_796,In_918);
nand U996 (N_996,In_850,In_336);
nor U997 (N_997,In_520,In_585);
nor U998 (N_998,In_347,In_756);
or U999 (N_999,In_144,In_411);
nor U1000 (N_1000,In_66,In_215);
xnor U1001 (N_1001,In_874,In_559);
and U1002 (N_1002,In_960,In_535);
and U1003 (N_1003,In_355,In_58);
nand U1004 (N_1004,In_10,In_941);
or U1005 (N_1005,In_577,In_576);
nor U1006 (N_1006,In_111,In_465);
and U1007 (N_1007,In_233,In_40);
or U1008 (N_1008,In_767,In_788);
nor U1009 (N_1009,In_910,In_643);
nor U1010 (N_1010,In_139,In_981);
or U1011 (N_1011,In_389,In_882);
nor U1012 (N_1012,In_441,In_228);
nor U1013 (N_1013,In_852,In_384);
and U1014 (N_1014,In_902,In_6);
or U1015 (N_1015,In_246,In_71);
nand U1016 (N_1016,In_798,In_115);
nand U1017 (N_1017,In_41,In_645);
nor U1018 (N_1018,In_627,In_77);
nand U1019 (N_1019,In_618,In_806);
or U1020 (N_1020,In_511,In_225);
nand U1021 (N_1021,In_706,In_33);
nand U1022 (N_1022,In_600,In_529);
nor U1023 (N_1023,In_668,In_7);
or U1024 (N_1024,In_168,In_69);
and U1025 (N_1025,In_414,In_264);
or U1026 (N_1026,In_259,In_698);
or U1027 (N_1027,In_762,In_511);
nor U1028 (N_1028,In_887,In_979);
and U1029 (N_1029,In_42,In_88);
and U1030 (N_1030,In_344,In_77);
nand U1031 (N_1031,In_212,In_37);
and U1032 (N_1032,In_508,In_192);
nand U1033 (N_1033,In_301,In_542);
and U1034 (N_1034,In_992,In_633);
nand U1035 (N_1035,In_458,In_832);
and U1036 (N_1036,In_853,In_942);
and U1037 (N_1037,In_71,In_437);
nor U1038 (N_1038,In_576,In_63);
nor U1039 (N_1039,In_416,In_925);
and U1040 (N_1040,In_731,In_146);
nand U1041 (N_1041,In_630,In_675);
nand U1042 (N_1042,In_274,In_659);
xor U1043 (N_1043,In_928,In_778);
nand U1044 (N_1044,In_979,In_501);
nand U1045 (N_1045,In_206,In_393);
nand U1046 (N_1046,In_255,In_760);
nand U1047 (N_1047,In_791,In_423);
or U1048 (N_1048,In_837,In_795);
or U1049 (N_1049,In_100,In_865);
and U1050 (N_1050,In_386,In_928);
nor U1051 (N_1051,In_68,In_13);
nand U1052 (N_1052,In_982,In_660);
and U1053 (N_1053,In_861,In_355);
nand U1054 (N_1054,In_397,In_980);
or U1055 (N_1055,In_34,In_22);
nor U1056 (N_1056,In_49,In_241);
or U1057 (N_1057,In_511,In_833);
nand U1058 (N_1058,In_683,In_356);
and U1059 (N_1059,In_418,In_55);
and U1060 (N_1060,In_954,In_67);
or U1061 (N_1061,In_594,In_352);
and U1062 (N_1062,In_476,In_321);
and U1063 (N_1063,In_702,In_563);
nor U1064 (N_1064,In_874,In_572);
or U1065 (N_1065,In_511,In_573);
nor U1066 (N_1066,In_905,In_550);
nor U1067 (N_1067,In_279,In_663);
nor U1068 (N_1068,In_359,In_51);
or U1069 (N_1069,In_936,In_426);
and U1070 (N_1070,In_124,In_314);
and U1071 (N_1071,In_719,In_814);
nand U1072 (N_1072,In_162,In_753);
nand U1073 (N_1073,In_427,In_282);
nor U1074 (N_1074,In_847,In_105);
or U1075 (N_1075,In_478,In_524);
and U1076 (N_1076,In_345,In_410);
nor U1077 (N_1077,In_519,In_884);
or U1078 (N_1078,In_593,In_106);
nor U1079 (N_1079,In_212,In_354);
nand U1080 (N_1080,In_436,In_703);
nand U1081 (N_1081,In_440,In_601);
or U1082 (N_1082,In_806,In_237);
nor U1083 (N_1083,In_390,In_537);
and U1084 (N_1084,In_451,In_585);
nand U1085 (N_1085,In_241,In_338);
or U1086 (N_1086,In_221,In_46);
and U1087 (N_1087,In_514,In_879);
or U1088 (N_1088,In_884,In_254);
and U1089 (N_1089,In_205,In_865);
or U1090 (N_1090,In_576,In_917);
and U1091 (N_1091,In_967,In_342);
or U1092 (N_1092,In_28,In_578);
and U1093 (N_1093,In_555,In_200);
and U1094 (N_1094,In_909,In_602);
nand U1095 (N_1095,In_402,In_258);
nand U1096 (N_1096,In_496,In_316);
nor U1097 (N_1097,In_318,In_932);
and U1098 (N_1098,In_953,In_413);
or U1099 (N_1099,In_832,In_790);
or U1100 (N_1100,In_754,In_311);
or U1101 (N_1101,In_236,In_172);
nand U1102 (N_1102,In_637,In_533);
nand U1103 (N_1103,In_266,In_12);
xnor U1104 (N_1104,In_511,In_468);
or U1105 (N_1105,In_9,In_986);
nand U1106 (N_1106,In_464,In_644);
and U1107 (N_1107,In_840,In_299);
nor U1108 (N_1108,In_905,In_525);
or U1109 (N_1109,In_952,In_132);
and U1110 (N_1110,In_690,In_121);
or U1111 (N_1111,In_316,In_419);
nor U1112 (N_1112,In_945,In_692);
or U1113 (N_1113,In_536,In_969);
and U1114 (N_1114,In_691,In_126);
nand U1115 (N_1115,In_935,In_981);
nand U1116 (N_1116,In_717,In_340);
nor U1117 (N_1117,In_936,In_793);
nor U1118 (N_1118,In_877,In_98);
or U1119 (N_1119,In_868,In_189);
nor U1120 (N_1120,In_712,In_797);
and U1121 (N_1121,In_974,In_556);
nand U1122 (N_1122,In_423,In_994);
and U1123 (N_1123,In_180,In_450);
xnor U1124 (N_1124,In_677,In_676);
nor U1125 (N_1125,In_683,In_889);
nand U1126 (N_1126,In_678,In_449);
and U1127 (N_1127,In_144,In_543);
nor U1128 (N_1128,In_573,In_154);
nand U1129 (N_1129,In_91,In_932);
nand U1130 (N_1130,In_166,In_626);
and U1131 (N_1131,In_765,In_97);
nand U1132 (N_1132,In_589,In_873);
or U1133 (N_1133,In_133,In_929);
xor U1134 (N_1134,In_748,In_296);
nand U1135 (N_1135,In_525,In_668);
nor U1136 (N_1136,In_300,In_439);
or U1137 (N_1137,In_452,In_747);
nor U1138 (N_1138,In_917,In_46);
nand U1139 (N_1139,In_173,In_43);
nand U1140 (N_1140,In_928,In_154);
nor U1141 (N_1141,In_475,In_587);
nor U1142 (N_1142,In_11,In_206);
and U1143 (N_1143,In_5,In_207);
and U1144 (N_1144,In_176,In_546);
and U1145 (N_1145,In_575,In_859);
nor U1146 (N_1146,In_418,In_101);
nand U1147 (N_1147,In_828,In_157);
and U1148 (N_1148,In_986,In_698);
or U1149 (N_1149,In_376,In_153);
or U1150 (N_1150,In_194,In_403);
nand U1151 (N_1151,In_17,In_105);
nand U1152 (N_1152,In_355,In_394);
nor U1153 (N_1153,In_307,In_207);
or U1154 (N_1154,In_663,In_860);
nand U1155 (N_1155,In_794,In_307);
or U1156 (N_1156,In_182,In_560);
and U1157 (N_1157,In_477,In_874);
or U1158 (N_1158,In_231,In_141);
and U1159 (N_1159,In_677,In_709);
and U1160 (N_1160,In_401,In_348);
and U1161 (N_1161,In_198,In_815);
nor U1162 (N_1162,In_829,In_344);
nor U1163 (N_1163,In_872,In_822);
and U1164 (N_1164,In_508,In_77);
nand U1165 (N_1165,In_908,In_306);
nor U1166 (N_1166,In_822,In_217);
nor U1167 (N_1167,In_647,In_873);
and U1168 (N_1168,In_894,In_358);
or U1169 (N_1169,In_430,In_631);
and U1170 (N_1170,In_392,In_571);
or U1171 (N_1171,In_127,In_558);
nor U1172 (N_1172,In_832,In_99);
nand U1173 (N_1173,In_466,In_51);
or U1174 (N_1174,In_201,In_352);
nor U1175 (N_1175,In_511,In_323);
nand U1176 (N_1176,In_935,In_380);
nand U1177 (N_1177,In_201,In_978);
and U1178 (N_1178,In_270,In_342);
and U1179 (N_1179,In_70,In_713);
and U1180 (N_1180,In_768,In_481);
and U1181 (N_1181,In_287,In_649);
and U1182 (N_1182,In_269,In_564);
nand U1183 (N_1183,In_752,In_826);
nand U1184 (N_1184,In_932,In_718);
or U1185 (N_1185,In_779,In_46);
or U1186 (N_1186,In_490,In_696);
nor U1187 (N_1187,In_488,In_875);
nand U1188 (N_1188,In_784,In_390);
and U1189 (N_1189,In_976,In_466);
and U1190 (N_1190,In_362,In_356);
nor U1191 (N_1191,In_488,In_67);
or U1192 (N_1192,In_962,In_927);
and U1193 (N_1193,In_385,In_59);
nor U1194 (N_1194,In_795,In_416);
and U1195 (N_1195,In_453,In_656);
or U1196 (N_1196,In_47,In_348);
nor U1197 (N_1197,In_246,In_754);
and U1198 (N_1198,In_321,In_549);
and U1199 (N_1199,In_980,In_235);
nand U1200 (N_1200,In_413,In_32);
and U1201 (N_1201,In_184,In_810);
and U1202 (N_1202,In_320,In_697);
or U1203 (N_1203,In_431,In_483);
nor U1204 (N_1204,In_90,In_747);
or U1205 (N_1205,In_589,In_295);
or U1206 (N_1206,In_865,In_619);
nand U1207 (N_1207,In_267,In_897);
and U1208 (N_1208,In_188,In_377);
nand U1209 (N_1209,In_887,In_445);
nor U1210 (N_1210,In_749,In_439);
nor U1211 (N_1211,In_73,In_307);
and U1212 (N_1212,In_100,In_796);
or U1213 (N_1213,In_734,In_175);
nand U1214 (N_1214,In_650,In_602);
or U1215 (N_1215,In_721,In_903);
nor U1216 (N_1216,In_497,In_787);
nand U1217 (N_1217,In_366,In_352);
nand U1218 (N_1218,In_49,In_67);
nor U1219 (N_1219,In_347,In_334);
nor U1220 (N_1220,In_454,In_446);
and U1221 (N_1221,In_431,In_557);
nand U1222 (N_1222,In_641,In_246);
and U1223 (N_1223,In_588,In_69);
and U1224 (N_1224,In_681,In_986);
and U1225 (N_1225,In_233,In_613);
and U1226 (N_1226,In_471,In_662);
nor U1227 (N_1227,In_549,In_884);
or U1228 (N_1228,In_858,In_740);
nor U1229 (N_1229,In_55,In_863);
nand U1230 (N_1230,In_444,In_325);
and U1231 (N_1231,In_756,In_96);
nor U1232 (N_1232,In_702,In_404);
nor U1233 (N_1233,In_443,In_940);
xnor U1234 (N_1234,In_898,In_515);
or U1235 (N_1235,In_76,In_80);
and U1236 (N_1236,In_724,In_957);
nand U1237 (N_1237,In_830,In_927);
and U1238 (N_1238,In_785,In_119);
nor U1239 (N_1239,In_66,In_686);
nor U1240 (N_1240,In_790,In_767);
or U1241 (N_1241,In_699,In_916);
or U1242 (N_1242,In_522,In_935);
nor U1243 (N_1243,In_320,In_574);
nand U1244 (N_1244,In_428,In_582);
or U1245 (N_1245,In_683,In_611);
and U1246 (N_1246,In_14,In_568);
nand U1247 (N_1247,In_740,In_976);
nor U1248 (N_1248,In_8,In_34);
nor U1249 (N_1249,In_567,In_978);
nor U1250 (N_1250,In_758,In_670);
and U1251 (N_1251,In_115,In_313);
or U1252 (N_1252,In_750,In_249);
or U1253 (N_1253,In_802,In_504);
nand U1254 (N_1254,In_141,In_788);
and U1255 (N_1255,In_5,In_558);
and U1256 (N_1256,In_888,In_906);
or U1257 (N_1257,In_441,In_283);
nand U1258 (N_1258,In_908,In_15);
and U1259 (N_1259,In_196,In_748);
and U1260 (N_1260,In_599,In_981);
nand U1261 (N_1261,In_187,In_827);
nand U1262 (N_1262,In_790,In_462);
or U1263 (N_1263,In_607,In_60);
nand U1264 (N_1264,In_546,In_250);
or U1265 (N_1265,In_492,In_364);
nand U1266 (N_1266,In_950,In_957);
nand U1267 (N_1267,In_891,In_585);
or U1268 (N_1268,In_329,In_754);
nand U1269 (N_1269,In_139,In_186);
nor U1270 (N_1270,In_60,In_574);
and U1271 (N_1271,In_185,In_622);
nor U1272 (N_1272,In_767,In_433);
nand U1273 (N_1273,In_171,In_946);
and U1274 (N_1274,In_219,In_661);
or U1275 (N_1275,In_590,In_290);
nor U1276 (N_1276,In_493,In_786);
and U1277 (N_1277,In_146,In_249);
nor U1278 (N_1278,In_726,In_587);
nor U1279 (N_1279,In_336,In_156);
or U1280 (N_1280,In_703,In_880);
or U1281 (N_1281,In_793,In_822);
or U1282 (N_1282,In_722,In_335);
nand U1283 (N_1283,In_940,In_378);
or U1284 (N_1284,In_135,In_487);
nand U1285 (N_1285,In_716,In_46);
nor U1286 (N_1286,In_990,In_382);
and U1287 (N_1287,In_588,In_97);
or U1288 (N_1288,In_632,In_656);
nand U1289 (N_1289,In_182,In_264);
and U1290 (N_1290,In_230,In_35);
or U1291 (N_1291,In_679,In_653);
nor U1292 (N_1292,In_880,In_983);
or U1293 (N_1293,In_707,In_969);
nor U1294 (N_1294,In_567,In_903);
nor U1295 (N_1295,In_91,In_627);
xnor U1296 (N_1296,In_108,In_892);
or U1297 (N_1297,In_942,In_321);
nand U1298 (N_1298,In_316,In_688);
nand U1299 (N_1299,In_980,In_940);
nor U1300 (N_1300,In_306,In_225);
or U1301 (N_1301,In_698,In_853);
or U1302 (N_1302,In_776,In_278);
nand U1303 (N_1303,In_321,In_355);
or U1304 (N_1304,In_203,In_864);
nand U1305 (N_1305,In_886,In_16);
nor U1306 (N_1306,In_467,In_887);
nor U1307 (N_1307,In_173,In_5);
or U1308 (N_1308,In_366,In_571);
or U1309 (N_1309,In_402,In_857);
and U1310 (N_1310,In_65,In_30);
xor U1311 (N_1311,In_496,In_826);
nand U1312 (N_1312,In_738,In_79);
or U1313 (N_1313,In_557,In_76);
or U1314 (N_1314,In_940,In_798);
nand U1315 (N_1315,In_437,In_740);
and U1316 (N_1316,In_942,In_177);
nor U1317 (N_1317,In_126,In_799);
and U1318 (N_1318,In_27,In_167);
nor U1319 (N_1319,In_187,In_149);
nand U1320 (N_1320,In_389,In_542);
and U1321 (N_1321,In_560,In_584);
or U1322 (N_1322,In_829,In_21);
nor U1323 (N_1323,In_202,In_346);
and U1324 (N_1324,In_174,In_143);
nor U1325 (N_1325,In_171,In_494);
and U1326 (N_1326,In_894,In_59);
and U1327 (N_1327,In_257,In_855);
or U1328 (N_1328,In_596,In_750);
and U1329 (N_1329,In_962,In_24);
xor U1330 (N_1330,In_21,In_750);
and U1331 (N_1331,In_265,In_347);
and U1332 (N_1332,In_603,In_24);
or U1333 (N_1333,In_537,In_653);
or U1334 (N_1334,In_466,In_298);
and U1335 (N_1335,In_262,In_161);
nor U1336 (N_1336,In_81,In_114);
or U1337 (N_1337,In_957,In_836);
nor U1338 (N_1338,In_330,In_46);
nand U1339 (N_1339,In_706,In_598);
nand U1340 (N_1340,In_896,In_310);
and U1341 (N_1341,In_869,In_690);
or U1342 (N_1342,In_775,In_809);
and U1343 (N_1343,In_52,In_64);
nor U1344 (N_1344,In_663,In_64);
or U1345 (N_1345,In_862,In_982);
nor U1346 (N_1346,In_618,In_782);
nand U1347 (N_1347,In_75,In_311);
and U1348 (N_1348,In_385,In_193);
and U1349 (N_1349,In_963,In_15);
or U1350 (N_1350,In_250,In_720);
nor U1351 (N_1351,In_647,In_889);
nor U1352 (N_1352,In_259,In_810);
nor U1353 (N_1353,In_545,In_973);
or U1354 (N_1354,In_97,In_675);
nor U1355 (N_1355,In_365,In_255);
or U1356 (N_1356,In_717,In_237);
nand U1357 (N_1357,In_990,In_549);
nand U1358 (N_1358,In_236,In_360);
or U1359 (N_1359,In_146,In_903);
and U1360 (N_1360,In_190,In_218);
nor U1361 (N_1361,In_761,In_652);
or U1362 (N_1362,In_66,In_850);
nor U1363 (N_1363,In_421,In_56);
and U1364 (N_1364,In_262,In_432);
or U1365 (N_1365,In_229,In_569);
nor U1366 (N_1366,In_732,In_735);
or U1367 (N_1367,In_587,In_546);
or U1368 (N_1368,In_191,In_219);
nand U1369 (N_1369,In_274,In_310);
nand U1370 (N_1370,In_940,In_35);
nand U1371 (N_1371,In_914,In_374);
nand U1372 (N_1372,In_851,In_186);
or U1373 (N_1373,In_813,In_596);
or U1374 (N_1374,In_828,In_830);
nor U1375 (N_1375,In_573,In_976);
and U1376 (N_1376,In_160,In_223);
or U1377 (N_1377,In_345,In_8);
nand U1378 (N_1378,In_24,In_687);
nand U1379 (N_1379,In_387,In_976);
and U1380 (N_1380,In_73,In_171);
and U1381 (N_1381,In_375,In_462);
nor U1382 (N_1382,In_721,In_336);
or U1383 (N_1383,In_83,In_8);
and U1384 (N_1384,In_653,In_210);
nor U1385 (N_1385,In_261,In_404);
nor U1386 (N_1386,In_798,In_153);
or U1387 (N_1387,In_663,In_82);
nand U1388 (N_1388,In_752,In_56);
nor U1389 (N_1389,In_682,In_794);
nor U1390 (N_1390,In_370,In_745);
and U1391 (N_1391,In_415,In_493);
nand U1392 (N_1392,In_161,In_630);
or U1393 (N_1393,In_577,In_794);
and U1394 (N_1394,In_757,In_452);
nor U1395 (N_1395,In_103,In_571);
nand U1396 (N_1396,In_882,In_829);
nor U1397 (N_1397,In_706,In_452);
nand U1398 (N_1398,In_896,In_924);
or U1399 (N_1399,In_237,In_384);
nor U1400 (N_1400,In_836,In_281);
nand U1401 (N_1401,In_703,In_863);
nor U1402 (N_1402,In_30,In_943);
and U1403 (N_1403,In_775,In_359);
nand U1404 (N_1404,In_625,In_167);
or U1405 (N_1405,In_481,In_568);
or U1406 (N_1406,In_356,In_784);
nor U1407 (N_1407,In_908,In_206);
nand U1408 (N_1408,In_975,In_870);
nand U1409 (N_1409,In_610,In_296);
xor U1410 (N_1410,In_798,In_685);
and U1411 (N_1411,In_882,In_839);
or U1412 (N_1412,In_822,In_778);
or U1413 (N_1413,In_534,In_293);
and U1414 (N_1414,In_676,In_810);
nor U1415 (N_1415,In_374,In_136);
or U1416 (N_1416,In_672,In_239);
or U1417 (N_1417,In_418,In_725);
and U1418 (N_1418,In_70,In_285);
nor U1419 (N_1419,In_274,In_939);
nor U1420 (N_1420,In_503,In_252);
nand U1421 (N_1421,In_579,In_219);
and U1422 (N_1422,In_795,In_158);
or U1423 (N_1423,In_204,In_750);
nand U1424 (N_1424,In_393,In_96);
nor U1425 (N_1425,In_574,In_267);
or U1426 (N_1426,In_136,In_341);
or U1427 (N_1427,In_582,In_723);
nand U1428 (N_1428,In_470,In_999);
xnor U1429 (N_1429,In_972,In_82);
and U1430 (N_1430,In_160,In_355);
and U1431 (N_1431,In_426,In_90);
and U1432 (N_1432,In_99,In_997);
or U1433 (N_1433,In_251,In_57);
or U1434 (N_1434,In_613,In_481);
nand U1435 (N_1435,In_986,In_767);
or U1436 (N_1436,In_833,In_221);
nand U1437 (N_1437,In_895,In_364);
nor U1438 (N_1438,In_84,In_710);
or U1439 (N_1439,In_762,In_771);
and U1440 (N_1440,In_131,In_409);
nand U1441 (N_1441,In_201,In_9);
nor U1442 (N_1442,In_535,In_621);
and U1443 (N_1443,In_345,In_120);
or U1444 (N_1444,In_388,In_577);
xor U1445 (N_1445,In_793,In_188);
or U1446 (N_1446,In_460,In_137);
and U1447 (N_1447,In_131,In_271);
and U1448 (N_1448,In_956,In_327);
and U1449 (N_1449,In_604,In_971);
and U1450 (N_1450,In_624,In_543);
or U1451 (N_1451,In_979,In_819);
nor U1452 (N_1452,In_305,In_490);
or U1453 (N_1453,In_989,In_206);
or U1454 (N_1454,In_74,In_875);
or U1455 (N_1455,In_172,In_347);
nand U1456 (N_1456,In_138,In_901);
and U1457 (N_1457,In_983,In_807);
and U1458 (N_1458,In_472,In_178);
and U1459 (N_1459,In_982,In_767);
nand U1460 (N_1460,In_987,In_208);
nor U1461 (N_1461,In_321,In_198);
or U1462 (N_1462,In_826,In_469);
and U1463 (N_1463,In_759,In_573);
nand U1464 (N_1464,In_889,In_698);
and U1465 (N_1465,In_960,In_407);
nor U1466 (N_1466,In_353,In_923);
nand U1467 (N_1467,In_647,In_162);
nor U1468 (N_1468,In_547,In_655);
or U1469 (N_1469,In_276,In_821);
nand U1470 (N_1470,In_949,In_196);
and U1471 (N_1471,In_126,In_835);
and U1472 (N_1472,In_46,In_5);
and U1473 (N_1473,In_956,In_973);
or U1474 (N_1474,In_570,In_445);
nor U1475 (N_1475,In_33,In_950);
xor U1476 (N_1476,In_393,In_741);
nor U1477 (N_1477,In_238,In_994);
nor U1478 (N_1478,In_142,In_790);
or U1479 (N_1479,In_236,In_600);
and U1480 (N_1480,In_607,In_367);
and U1481 (N_1481,In_897,In_407);
nor U1482 (N_1482,In_286,In_482);
nand U1483 (N_1483,In_930,In_245);
or U1484 (N_1484,In_660,In_546);
nand U1485 (N_1485,In_565,In_723);
nor U1486 (N_1486,In_65,In_761);
nand U1487 (N_1487,In_456,In_652);
nand U1488 (N_1488,In_295,In_738);
nand U1489 (N_1489,In_227,In_163);
nand U1490 (N_1490,In_159,In_759);
and U1491 (N_1491,In_533,In_144);
or U1492 (N_1492,In_209,In_332);
or U1493 (N_1493,In_650,In_99);
nand U1494 (N_1494,In_780,In_847);
nand U1495 (N_1495,In_544,In_343);
or U1496 (N_1496,In_481,In_124);
nand U1497 (N_1497,In_256,In_909);
or U1498 (N_1498,In_337,In_718);
nor U1499 (N_1499,In_516,In_597);
nand U1500 (N_1500,In_346,In_165);
nor U1501 (N_1501,In_492,In_267);
nor U1502 (N_1502,In_487,In_570);
and U1503 (N_1503,In_500,In_347);
nor U1504 (N_1504,In_916,In_36);
nand U1505 (N_1505,In_310,In_857);
nand U1506 (N_1506,In_636,In_785);
or U1507 (N_1507,In_742,In_947);
and U1508 (N_1508,In_457,In_81);
nand U1509 (N_1509,In_929,In_13);
and U1510 (N_1510,In_440,In_467);
nand U1511 (N_1511,In_567,In_998);
and U1512 (N_1512,In_109,In_210);
or U1513 (N_1513,In_986,In_464);
and U1514 (N_1514,In_49,In_421);
nor U1515 (N_1515,In_598,In_288);
nor U1516 (N_1516,In_616,In_11);
or U1517 (N_1517,In_621,In_230);
or U1518 (N_1518,In_500,In_473);
or U1519 (N_1519,In_683,In_811);
or U1520 (N_1520,In_294,In_240);
or U1521 (N_1521,In_613,In_238);
nor U1522 (N_1522,In_764,In_838);
and U1523 (N_1523,In_910,In_638);
and U1524 (N_1524,In_467,In_830);
nor U1525 (N_1525,In_265,In_283);
and U1526 (N_1526,In_242,In_743);
nor U1527 (N_1527,In_894,In_263);
and U1528 (N_1528,In_963,In_50);
nand U1529 (N_1529,In_331,In_797);
nor U1530 (N_1530,In_33,In_247);
and U1531 (N_1531,In_836,In_982);
or U1532 (N_1532,In_101,In_388);
nand U1533 (N_1533,In_731,In_843);
nor U1534 (N_1534,In_41,In_399);
nor U1535 (N_1535,In_493,In_662);
nand U1536 (N_1536,In_363,In_381);
nand U1537 (N_1537,In_297,In_486);
and U1538 (N_1538,In_927,In_674);
nor U1539 (N_1539,In_882,In_128);
and U1540 (N_1540,In_559,In_901);
nand U1541 (N_1541,In_398,In_817);
or U1542 (N_1542,In_179,In_619);
or U1543 (N_1543,In_857,In_237);
nor U1544 (N_1544,In_119,In_658);
or U1545 (N_1545,In_279,In_638);
nor U1546 (N_1546,In_879,In_257);
and U1547 (N_1547,In_841,In_885);
or U1548 (N_1548,In_893,In_577);
and U1549 (N_1549,In_990,In_710);
nand U1550 (N_1550,In_649,In_235);
nand U1551 (N_1551,In_787,In_157);
nand U1552 (N_1552,In_230,In_266);
nor U1553 (N_1553,In_483,In_279);
nand U1554 (N_1554,In_79,In_25);
or U1555 (N_1555,In_904,In_283);
nand U1556 (N_1556,In_868,In_584);
nand U1557 (N_1557,In_618,In_838);
nand U1558 (N_1558,In_926,In_930);
nand U1559 (N_1559,In_679,In_176);
or U1560 (N_1560,In_4,In_422);
and U1561 (N_1561,In_496,In_878);
and U1562 (N_1562,In_848,In_366);
and U1563 (N_1563,In_284,In_228);
or U1564 (N_1564,In_413,In_321);
or U1565 (N_1565,In_665,In_520);
nor U1566 (N_1566,In_724,In_434);
or U1567 (N_1567,In_684,In_564);
and U1568 (N_1568,In_846,In_798);
and U1569 (N_1569,In_602,In_162);
and U1570 (N_1570,In_664,In_229);
and U1571 (N_1571,In_743,In_579);
nor U1572 (N_1572,In_210,In_145);
or U1573 (N_1573,In_606,In_412);
nand U1574 (N_1574,In_899,In_956);
and U1575 (N_1575,In_934,In_444);
or U1576 (N_1576,In_696,In_232);
nand U1577 (N_1577,In_882,In_518);
and U1578 (N_1578,In_602,In_464);
nor U1579 (N_1579,In_937,In_105);
and U1580 (N_1580,In_931,In_476);
nor U1581 (N_1581,In_320,In_802);
nor U1582 (N_1582,In_971,In_683);
nor U1583 (N_1583,In_585,In_985);
and U1584 (N_1584,In_164,In_575);
nand U1585 (N_1585,In_291,In_387);
nor U1586 (N_1586,In_471,In_720);
and U1587 (N_1587,In_614,In_937);
nand U1588 (N_1588,In_877,In_706);
and U1589 (N_1589,In_73,In_551);
or U1590 (N_1590,In_413,In_199);
nand U1591 (N_1591,In_627,In_690);
nand U1592 (N_1592,In_962,In_392);
or U1593 (N_1593,In_316,In_410);
or U1594 (N_1594,In_756,In_785);
nand U1595 (N_1595,In_523,In_241);
or U1596 (N_1596,In_441,In_314);
nand U1597 (N_1597,In_276,In_397);
and U1598 (N_1598,In_770,In_862);
nor U1599 (N_1599,In_288,In_71);
or U1600 (N_1600,In_963,In_11);
nand U1601 (N_1601,In_400,In_925);
and U1602 (N_1602,In_656,In_644);
and U1603 (N_1603,In_815,In_773);
or U1604 (N_1604,In_918,In_590);
nand U1605 (N_1605,In_570,In_706);
and U1606 (N_1606,In_807,In_702);
nand U1607 (N_1607,In_648,In_330);
nand U1608 (N_1608,In_960,In_356);
nor U1609 (N_1609,In_39,In_470);
or U1610 (N_1610,In_783,In_619);
nand U1611 (N_1611,In_589,In_75);
nand U1612 (N_1612,In_261,In_131);
nand U1613 (N_1613,In_214,In_165);
or U1614 (N_1614,In_302,In_457);
and U1615 (N_1615,In_446,In_67);
and U1616 (N_1616,In_290,In_963);
nor U1617 (N_1617,In_567,In_108);
nand U1618 (N_1618,In_337,In_122);
nand U1619 (N_1619,In_966,In_636);
and U1620 (N_1620,In_774,In_732);
nor U1621 (N_1621,In_988,In_966);
or U1622 (N_1622,In_693,In_726);
nor U1623 (N_1623,In_919,In_691);
or U1624 (N_1624,In_760,In_175);
and U1625 (N_1625,In_547,In_196);
nand U1626 (N_1626,In_216,In_601);
and U1627 (N_1627,In_851,In_273);
nor U1628 (N_1628,In_105,In_468);
nor U1629 (N_1629,In_97,In_25);
nand U1630 (N_1630,In_660,In_642);
or U1631 (N_1631,In_836,In_505);
nor U1632 (N_1632,In_679,In_907);
nor U1633 (N_1633,In_862,In_370);
and U1634 (N_1634,In_163,In_664);
nor U1635 (N_1635,In_419,In_227);
nand U1636 (N_1636,In_561,In_666);
or U1637 (N_1637,In_542,In_396);
nand U1638 (N_1638,In_470,In_41);
or U1639 (N_1639,In_280,In_76);
and U1640 (N_1640,In_273,In_211);
and U1641 (N_1641,In_440,In_316);
or U1642 (N_1642,In_339,In_245);
and U1643 (N_1643,In_774,In_633);
nor U1644 (N_1644,In_9,In_768);
nand U1645 (N_1645,In_929,In_27);
and U1646 (N_1646,In_143,In_879);
nor U1647 (N_1647,In_986,In_799);
and U1648 (N_1648,In_897,In_831);
xor U1649 (N_1649,In_505,In_740);
nand U1650 (N_1650,In_721,In_194);
nand U1651 (N_1651,In_485,In_589);
nor U1652 (N_1652,In_604,In_876);
nor U1653 (N_1653,In_772,In_216);
nor U1654 (N_1654,In_591,In_719);
nor U1655 (N_1655,In_280,In_363);
and U1656 (N_1656,In_837,In_895);
and U1657 (N_1657,In_992,In_430);
nand U1658 (N_1658,In_264,In_835);
and U1659 (N_1659,In_963,In_873);
or U1660 (N_1660,In_208,In_773);
nor U1661 (N_1661,In_438,In_799);
nand U1662 (N_1662,In_914,In_607);
nand U1663 (N_1663,In_676,In_594);
xnor U1664 (N_1664,In_622,In_75);
or U1665 (N_1665,In_165,In_567);
nor U1666 (N_1666,In_446,In_153);
or U1667 (N_1667,In_321,In_924);
nor U1668 (N_1668,In_326,In_177);
or U1669 (N_1669,In_170,In_722);
and U1670 (N_1670,In_473,In_876);
nand U1671 (N_1671,In_718,In_941);
or U1672 (N_1672,In_850,In_666);
xor U1673 (N_1673,In_871,In_47);
or U1674 (N_1674,In_125,In_645);
or U1675 (N_1675,In_573,In_170);
and U1676 (N_1676,In_504,In_336);
nor U1677 (N_1677,In_261,In_522);
nor U1678 (N_1678,In_487,In_796);
or U1679 (N_1679,In_135,In_352);
nor U1680 (N_1680,In_312,In_194);
or U1681 (N_1681,In_3,In_183);
xnor U1682 (N_1682,In_205,In_334);
and U1683 (N_1683,In_724,In_394);
nor U1684 (N_1684,In_288,In_937);
nand U1685 (N_1685,In_434,In_455);
or U1686 (N_1686,In_721,In_641);
or U1687 (N_1687,In_709,In_215);
and U1688 (N_1688,In_249,In_72);
and U1689 (N_1689,In_755,In_40);
nand U1690 (N_1690,In_804,In_428);
nor U1691 (N_1691,In_147,In_602);
nor U1692 (N_1692,In_57,In_349);
nand U1693 (N_1693,In_829,In_159);
nand U1694 (N_1694,In_993,In_15);
nor U1695 (N_1695,In_691,In_850);
nor U1696 (N_1696,In_746,In_846);
nand U1697 (N_1697,In_435,In_600);
or U1698 (N_1698,In_370,In_569);
and U1699 (N_1699,In_143,In_52);
nand U1700 (N_1700,In_331,In_615);
nor U1701 (N_1701,In_136,In_102);
nand U1702 (N_1702,In_139,In_932);
nand U1703 (N_1703,In_607,In_104);
or U1704 (N_1704,In_588,In_795);
nor U1705 (N_1705,In_11,In_584);
and U1706 (N_1706,In_565,In_862);
or U1707 (N_1707,In_181,In_288);
nand U1708 (N_1708,In_584,In_622);
and U1709 (N_1709,In_759,In_264);
or U1710 (N_1710,In_507,In_401);
and U1711 (N_1711,In_161,In_467);
nor U1712 (N_1712,In_761,In_671);
or U1713 (N_1713,In_186,In_902);
nand U1714 (N_1714,In_733,In_72);
nand U1715 (N_1715,In_768,In_91);
and U1716 (N_1716,In_356,In_498);
nand U1717 (N_1717,In_410,In_757);
nand U1718 (N_1718,In_432,In_369);
nor U1719 (N_1719,In_529,In_51);
nor U1720 (N_1720,In_24,In_392);
nand U1721 (N_1721,In_145,In_823);
nor U1722 (N_1722,In_271,In_742);
or U1723 (N_1723,In_42,In_888);
or U1724 (N_1724,In_621,In_181);
or U1725 (N_1725,In_731,In_99);
and U1726 (N_1726,In_859,In_729);
or U1727 (N_1727,In_660,In_188);
nand U1728 (N_1728,In_676,In_311);
and U1729 (N_1729,In_329,In_402);
nor U1730 (N_1730,In_268,In_840);
nand U1731 (N_1731,In_769,In_691);
nor U1732 (N_1732,In_433,In_224);
nor U1733 (N_1733,In_817,In_977);
nor U1734 (N_1734,In_337,In_371);
nor U1735 (N_1735,In_93,In_154);
nor U1736 (N_1736,In_75,In_867);
nor U1737 (N_1737,In_816,In_996);
nand U1738 (N_1738,In_545,In_955);
nor U1739 (N_1739,In_661,In_892);
and U1740 (N_1740,In_465,In_369);
and U1741 (N_1741,In_529,In_665);
or U1742 (N_1742,In_112,In_447);
nand U1743 (N_1743,In_946,In_288);
and U1744 (N_1744,In_206,In_42);
or U1745 (N_1745,In_77,In_606);
or U1746 (N_1746,In_756,In_988);
or U1747 (N_1747,In_31,In_385);
nor U1748 (N_1748,In_182,In_822);
or U1749 (N_1749,In_106,In_217);
or U1750 (N_1750,In_128,In_28);
nand U1751 (N_1751,In_914,In_526);
nand U1752 (N_1752,In_607,In_249);
nor U1753 (N_1753,In_863,In_751);
and U1754 (N_1754,In_426,In_165);
and U1755 (N_1755,In_44,In_674);
nand U1756 (N_1756,In_285,In_1);
and U1757 (N_1757,In_978,In_823);
nand U1758 (N_1758,In_339,In_497);
nor U1759 (N_1759,In_755,In_861);
and U1760 (N_1760,In_373,In_498);
and U1761 (N_1761,In_962,In_403);
nor U1762 (N_1762,In_679,In_738);
nor U1763 (N_1763,In_451,In_12);
nand U1764 (N_1764,In_699,In_706);
nor U1765 (N_1765,In_857,In_447);
and U1766 (N_1766,In_789,In_767);
nand U1767 (N_1767,In_972,In_730);
or U1768 (N_1768,In_420,In_964);
nand U1769 (N_1769,In_55,In_278);
or U1770 (N_1770,In_582,In_861);
or U1771 (N_1771,In_328,In_536);
nor U1772 (N_1772,In_806,In_309);
or U1773 (N_1773,In_449,In_111);
nor U1774 (N_1774,In_896,In_776);
nor U1775 (N_1775,In_564,In_429);
and U1776 (N_1776,In_320,In_674);
and U1777 (N_1777,In_336,In_787);
and U1778 (N_1778,In_666,In_621);
nand U1779 (N_1779,In_253,In_884);
nor U1780 (N_1780,In_331,In_495);
and U1781 (N_1781,In_167,In_885);
nand U1782 (N_1782,In_515,In_427);
nand U1783 (N_1783,In_312,In_133);
nor U1784 (N_1784,In_777,In_137);
and U1785 (N_1785,In_802,In_106);
and U1786 (N_1786,In_527,In_38);
or U1787 (N_1787,In_456,In_784);
or U1788 (N_1788,In_891,In_702);
and U1789 (N_1789,In_860,In_208);
and U1790 (N_1790,In_816,In_824);
and U1791 (N_1791,In_780,In_954);
or U1792 (N_1792,In_408,In_102);
and U1793 (N_1793,In_360,In_755);
xnor U1794 (N_1794,In_46,In_150);
or U1795 (N_1795,In_75,In_620);
and U1796 (N_1796,In_20,In_619);
nand U1797 (N_1797,In_868,In_767);
nor U1798 (N_1798,In_9,In_742);
and U1799 (N_1799,In_451,In_362);
nor U1800 (N_1800,In_864,In_914);
nor U1801 (N_1801,In_452,In_398);
nand U1802 (N_1802,In_235,In_146);
or U1803 (N_1803,In_593,In_434);
nor U1804 (N_1804,In_62,In_93);
and U1805 (N_1805,In_444,In_850);
or U1806 (N_1806,In_397,In_910);
nand U1807 (N_1807,In_91,In_949);
nor U1808 (N_1808,In_344,In_46);
and U1809 (N_1809,In_589,In_468);
nand U1810 (N_1810,In_542,In_442);
nor U1811 (N_1811,In_974,In_792);
nand U1812 (N_1812,In_203,In_0);
or U1813 (N_1813,In_427,In_415);
or U1814 (N_1814,In_737,In_35);
nand U1815 (N_1815,In_179,In_183);
and U1816 (N_1816,In_957,In_441);
nor U1817 (N_1817,In_35,In_593);
and U1818 (N_1818,In_770,In_369);
nor U1819 (N_1819,In_268,In_393);
nand U1820 (N_1820,In_105,In_426);
nand U1821 (N_1821,In_402,In_134);
nor U1822 (N_1822,In_656,In_711);
or U1823 (N_1823,In_238,In_1);
and U1824 (N_1824,In_51,In_181);
and U1825 (N_1825,In_303,In_335);
or U1826 (N_1826,In_615,In_16);
and U1827 (N_1827,In_47,In_612);
nor U1828 (N_1828,In_626,In_446);
nand U1829 (N_1829,In_753,In_415);
nor U1830 (N_1830,In_308,In_871);
and U1831 (N_1831,In_226,In_160);
or U1832 (N_1832,In_734,In_968);
nor U1833 (N_1833,In_923,In_829);
nand U1834 (N_1834,In_583,In_939);
and U1835 (N_1835,In_417,In_220);
and U1836 (N_1836,In_389,In_106);
and U1837 (N_1837,In_722,In_791);
nand U1838 (N_1838,In_201,In_898);
or U1839 (N_1839,In_512,In_658);
nand U1840 (N_1840,In_365,In_443);
nand U1841 (N_1841,In_750,In_630);
nor U1842 (N_1842,In_566,In_287);
or U1843 (N_1843,In_117,In_770);
nor U1844 (N_1844,In_385,In_362);
xnor U1845 (N_1845,In_888,In_264);
nor U1846 (N_1846,In_342,In_477);
nor U1847 (N_1847,In_723,In_941);
and U1848 (N_1848,In_274,In_39);
and U1849 (N_1849,In_30,In_451);
nor U1850 (N_1850,In_221,In_175);
or U1851 (N_1851,In_930,In_755);
nor U1852 (N_1852,In_648,In_596);
and U1853 (N_1853,In_707,In_797);
nand U1854 (N_1854,In_13,In_604);
nor U1855 (N_1855,In_398,In_824);
nand U1856 (N_1856,In_497,In_879);
nor U1857 (N_1857,In_18,In_20);
nand U1858 (N_1858,In_187,In_279);
nand U1859 (N_1859,In_794,In_915);
nand U1860 (N_1860,In_708,In_373);
nand U1861 (N_1861,In_400,In_287);
and U1862 (N_1862,In_423,In_868);
nand U1863 (N_1863,In_78,In_18);
nand U1864 (N_1864,In_305,In_965);
and U1865 (N_1865,In_258,In_696);
nor U1866 (N_1866,In_822,In_874);
and U1867 (N_1867,In_903,In_565);
or U1868 (N_1868,In_958,In_700);
and U1869 (N_1869,In_15,In_468);
nor U1870 (N_1870,In_591,In_961);
and U1871 (N_1871,In_477,In_997);
nand U1872 (N_1872,In_471,In_629);
or U1873 (N_1873,In_608,In_912);
nand U1874 (N_1874,In_489,In_811);
nor U1875 (N_1875,In_358,In_415);
nor U1876 (N_1876,In_122,In_825);
nand U1877 (N_1877,In_346,In_32);
nand U1878 (N_1878,In_657,In_451);
nand U1879 (N_1879,In_448,In_729);
nor U1880 (N_1880,In_6,In_256);
nor U1881 (N_1881,In_521,In_33);
or U1882 (N_1882,In_99,In_744);
and U1883 (N_1883,In_522,In_223);
nand U1884 (N_1884,In_984,In_950);
and U1885 (N_1885,In_797,In_358);
or U1886 (N_1886,In_941,In_31);
or U1887 (N_1887,In_124,In_792);
nand U1888 (N_1888,In_30,In_768);
and U1889 (N_1889,In_166,In_95);
and U1890 (N_1890,In_952,In_499);
and U1891 (N_1891,In_390,In_96);
nand U1892 (N_1892,In_459,In_670);
nor U1893 (N_1893,In_575,In_289);
or U1894 (N_1894,In_579,In_747);
and U1895 (N_1895,In_984,In_488);
and U1896 (N_1896,In_301,In_340);
and U1897 (N_1897,In_431,In_600);
and U1898 (N_1898,In_929,In_251);
and U1899 (N_1899,In_925,In_714);
nor U1900 (N_1900,In_833,In_754);
or U1901 (N_1901,In_8,In_1);
nor U1902 (N_1902,In_933,In_538);
nor U1903 (N_1903,In_711,In_653);
and U1904 (N_1904,In_615,In_866);
nor U1905 (N_1905,In_87,In_533);
or U1906 (N_1906,In_309,In_136);
or U1907 (N_1907,In_589,In_884);
nor U1908 (N_1908,In_72,In_125);
nor U1909 (N_1909,In_16,In_963);
and U1910 (N_1910,In_570,In_115);
nand U1911 (N_1911,In_817,In_70);
nand U1912 (N_1912,In_891,In_165);
nor U1913 (N_1913,In_811,In_814);
and U1914 (N_1914,In_531,In_818);
nor U1915 (N_1915,In_306,In_663);
nand U1916 (N_1916,In_660,In_343);
and U1917 (N_1917,In_628,In_386);
nand U1918 (N_1918,In_732,In_813);
and U1919 (N_1919,In_98,In_924);
nor U1920 (N_1920,In_337,In_24);
nor U1921 (N_1921,In_866,In_191);
nor U1922 (N_1922,In_371,In_243);
nor U1923 (N_1923,In_52,In_471);
nor U1924 (N_1924,In_208,In_296);
and U1925 (N_1925,In_209,In_435);
or U1926 (N_1926,In_535,In_294);
and U1927 (N_1927,In_877,In_474);
or U1928 (N_1928,In_756,In_34);
and U1929 (N_1929,In_21,In_419);
and U1930 (N_1930,In_246,In_127);
and U1931 (N_1931,In_645,In_642);
nand U1932 (N_1932,In_431,In_247);
or U1933 (N_1933,In_981,In_6);
nor U1934 (N_1934,In_360,In_640);
and U1935 (N_1935,In_647,In_140);
and U1936 (N_1936,In_80,In_904);
or U1937 (N_1937,In_67,In_715);
and U1938 (N_1938,In_752,In_848);
nor U1939 (N_1939,In_669,In_864);
nand U1940 (N_1940,In_15,In_876);
or U1941 (N_1941,In_139,In_862);
and U1942 (N_1942,In_208,In_152);
nand U1943 (N_1943,In_954,In_454);
or U1944 (N_1944,In_657,In_542);
or U1945 (N_1945,In_539,In_198);
and U1946 (N_1946,In_10,In_767);
nor U1947 (N_1947,In_651,In_717);
and U1948 (N_1948,In_233,In_798);
nand U1949 (N_1949,In_989,In_655);
and U1950 (N_1950,In_106,In_12);
nor U1951 (N_1951,In_891,In_313);
nand U1952 (N_1952,In_417,In_77);
or U1953 (N_1953,In_294,In_940);
nand U1954 (N_1954,In_999,In_895);
or U1955 (N_1955,In_312,In_137);
nand U1956 (N_1956,In_982,In_724);
or U1957 (N_1957,In_377,In_991);
nor U1958 (N_1958,In_373,In_684);
and U1959 (N_1959,In_667,In_51);
and U1960 (N_1960,In_943,In_0);
and U1961 (N_1961,In_50,In_798);
and U1962 (N_1962,In_407,In_888);
or U1963 (N_1963,In_737,In_411);
or U1964 (N_1964,In_332,In_555);
nand U1965 (N_1965,In_942,In_41);
or U1966 (N_1966,In_865,In_162);
or U1967 (N_1967,In_161,In_203);
and U1968 (N_1968,In_877,In_393);
nor U1969 (N_1969,In_67,In_735);
nand U1970 (N_1970,In_151,In_551);
nor U1971 (N_1971,In_296,In_21);
and U1972 (N_1972,In_547,In_621);
and U1973 (N_1973,In_340,In_764);
and U1974 (N_1974,In_242,In_154);
nor U1975 (N_1975,In_963,In_60);
or U1976 (N_1976,In_789,In_299);
or U1977 (N_1977,In_570,In_196);
and U1978 (N_1978,In_949,In_455);
and U1979 (N_1979,In_943,In_127);
and U1980 (N_1980,In_666,In_849);
or U1981 (N_1981,In_348,In_492);
nand U1982 (N_1982,In_550,In_734);
or U1983 (N_1983,In_231,In_856);
nor U1984 (N_1984,In_927,In_479);
or U1985 (N_1985,In_980,In_730);
or U1986 (N_1986,In_355,In_493);
and U1987 (N_1987,In_459,In_973);
and U1988 (N_1988,In_10,In_412);
or U1989 (N_1989,In_946,In_167);
nor U1990 (N_1990,In_960,In_793);
and U1991 (N_1991,In_615,In_374);
nand U1992 (N_1992,In_952,In_753);
nor U1993 (N_1993,In_338,In_34);
nand U1994 (N_1994,In_160,In_649);
nor U1995 (N_1995,In_428,In_700);
nor U1996 (N_1996,In_876,In_271);
nor U1997 (N_1997,In_646,In_141);
nand U1998 (N_1998,In_455,In_888);
or U1999 (N_1999,In_561,In_475);
nand U2000 (N_2000,In_955,In_851);
nand U2001 (N_2001,In_616,In_92);
nand U2002 (N_2002,In_335,In_492);
nor U2003 (N_2003,In_808,In_811);
and U2004 (N_2004,In_284,In_349);
nand U2005 (N_2005,In_937,In_598);
nand U2006 (N_2006,In_95,In_454);
or U2007 (N_2007,In_548,In_5);
nand U2008 (N_2008,In_742,In_300);
nand U2009 (N_2009,In_905,In_658);
and U2010 (N_2010,In_248,In_195);
or U2011 (N_2011,In_822,In_808);
nor U2012 (N_2012,In_955,In_190);
or U2013 (N_2013,In_138,In_773);
or U2014 (N_2014,In_344,In_927);
or U2015 (N_2015,In_792,In_598);
nand U2016 (N_2016,In_40,In_382);
nand U2017 (N_2017,In_277,In_19);
or U2018 (N_2018,In_714,In_881);
or U2019 (N_2019,In_892,In_933);
nor U2020 (N_2020,In_477,In_221);
or U2021 (N_2021,In_115,In_941);
or U2022 (N_2022,In_65,In_987);
or U2023 (N_2023,In_992,In_982);
nand U2024 (N_2024,In_922,In_19);
nand U2025 (N_2025,In_163,In_976);
and U2026 (N_2026,In_660,In_857);
nand U2027 (N_2027,In_159,In_372);
and U2028 (N_2028,In_549,In_915);
xnor U2029 (N_2029,In_428,In_895);
and U2030 (N_2030,In_614,In_914);
nor U2031 (N_2031,In_800,In_555);
and U2032 (N_2032,In_305,In_580);
or U2033 (N_2033,In_140,In_307);
nand U2034 (N_2034,In_113,In_709);
and U2035 (N_2035,In_66,In_837);
nor U2036 (N_2036,In_145,In_939);
nand U2037 (N_2037,In_876,In_559);
or U2038 (N_2038,In_944,In_372);
nor U2039 (N_2039,In_369,In_938);
and U2040 (N_2040,In_318,In_185);
or U2041 (N_2041,In_378,In_481);
and U2042 (N_2042,In_815,In_86);
or U2043 (N_2043,In_110,In_269);
and U2044 (N_2044,In_827,In_755);
or U2045 (N_2045,In_704,In_525);
or U2046 (N_2046,In_194,In_365);
nor U2047 (N_2047,In_747,In_895);
nand U2048 (N_2048,In_340,In_291);
nor U2049 (N_2049,In_347,In_476);
nand U2050 (N_2050,In_747,In_701);
nor U2051 (N_2051,In_143,In_252);
nand U2052 (N_2052,In_217,In_348);
nor U2053 (N_2053,In_41,In_391);
and U2054 (N_2054,In_26,In_629);
and U2055 (N_2055,In_867,In_99);
or U2056 (N_2056,In_719,In_830);
nand U2057 (N_2057,In_799,In_994);
or U2058 (N_2058,In_905,In_733);
or U2059 (N_2059,In_2,In_196);
nor U2060 (N_2060,In_129,In_87);
or U2061 (N_2061,In_515,In_528);
nor U2062 (N_2062,In_670,In_928);
and U2063 (N_2063,In_453,In_564);
or U2064 (N_2064,In_910,In_915);
nor U2065 (N_2065,In_20,In_33);
and U2066 (N_2066,In_744,In_109);
nand U2067 (N_2067,In_346,In_64);
nor U2068 (N_2068,In_250,In_834);
nor U2069 (N_2069,In_53,In_788);
nand U2070 (N_2070,In_860,In_837);
nand U2071 (N_2071,In_847,In_606);
or U2072 (N_2072,In_102,In_92);
or U2073 (N_2073,In_515,In_940);
and U2074 (N_2074,In_65,In_856);
or U2075 (N_2075,In_661,In_18);
nor U2076 (N_2076,In_540,In_232);
nor U2077 (N_2077,In_266,In_332);
and U2078 (N_2078,In_981,In_223);
and U2079 (N_2079,In_327,In_791);
nor U2080 (N_2080,In_62,In_260);
or U2081 (N_2081,In_625,In_637);
and U2082 (N_2082,In_117,In_815);
nor U2083 (N_2083,In_53,In_214);
and U2084 (N_2084,In_170,In_696);
nor U2085 (N_2085,In_361,In_590);
and U2086 (N_2086,In_495,In_328);
and U2087 (N_2087,In_519,In_869);
nor U2088 (N_2088,In_754,In_188);
or U2089 (N_2089,In_83,In_749);
and U2090 (N_2090,In_389,In_576);
nor U2091 (N_2091,In_880,In_823);
and U2092 (N_2092,In_47,In_778);
or U2093 (N_2093,In_339,In_921);
and U2094 (N_2094,In_428,In_730);
nand U2095 (N_2095,In_643,In_683);
nand U2096 (N_2096,In_246,In_215);
nor U2097 (N_2097,In_324,In_457);
nand U2098 (N_2098,In_353,In_238);
nand U2099 (N_2099,In_270,In_473);
nor U2100 (N_2100,In_671,In_760);
nor U2101 (N_2101,In_847,In_916);
and U2102 (N_2102,In_870,In_623);
nor U2103 (N_2103,In_542,In_835);
and U2104 (N_2104,In_358,In_532);
or U2105 (N_2105,In_117,In_173);
or U2106 (N_2106,In_30,In_465);
nand U2107 (N_2107,In_726,In_160);
or U2108 (N_2108,In_798,In_910);
nand U2109 (N_2109,In_435,In_291);
nand U2110 (N_2110,In_72,In_560);
or U2111 (N_2111,In_380,In_454);
nand U2112 (N_2112,In_795,In_398);
or U2113 (N_2113,In_382,In_118);
nand U2114 (N_2114,In_507,In_224);
and U2115 (N_2115,In_243,In_8);
or U2116 (N_2116,In_758,In_818);
and U2117 (N_2117,In_241,In_309);
and U2118 (N_2118,In_244,In_554);
or U2119 (N_2119,In_501,In_90);
or U2120 (N_2120,In_152,In_965);
nand U2121 (N_2121,In_49,In_549);
or U2122 (N_2122,In_258,In_974);
or U2123 (N_2123,In_138,In_839);
and U2124 (N_2124,In_634,In_143);
nand U2125 (N_2125,In_435,In_431);
nor U2126 (N_2126,In_251,In_454);
or U2127 (N_2127,In_647,In_583);
or U2128 (N_2128,In_823,In_547);
nand U2129 (N_2129,In_559,In_611);
nand U2130 (N_2130,In_920,In_312);
and U2131 (N_2131,In_67,In_864);
or U2132 (N_2132,In_688,In_705);
nand U2133 (N_2133,In_879,In_468);
and U2134 (N_2134,In_107,In_935);
and U2135 (N_2135,In_361,In_193);
and U2136 (N_2136,In_916,In_88);
nand U2137 (N_2137,In_455,In_693);
or U2138 (N_2138,In_360,In_468);
and U2139 (N_2139,In_162,In_972);
or U2140 (N_2140,In_260,In_794);
and U2141 (N_2141,In_957,In_584);
nand U2142 (N_2142,In_612,In_244);
nand U2143 (N_2143,In_867,In_35);
and U2144 (N_2144,In_639,In_638);
nand U2145 (N_2145,In_182,In_585);
and U2146 (N_2146,In_327,In_922);
nor U2147 (N_2147,In_896,In_930);
or U2148 (N_2148,In_485,In_228);
nor U2149 (N_2149,In_345,In_227);
or U2150 (N_2150,In_198,In_766);
and U2151 (N_2151,In_683,In_6);
nand U2152 (N_2152,In_380,In_968);
or U2153 (N_2153,In_599,In_557);
nand U2154 (N_2154,In_273,In_152);
and U2155 (N_2155,In_654,In_73);
and U2156 (N_2156,In_409,In_711);
and U2157 (N_2157,In_513,In_365);
or U2158 (N_2158,In_591,In_281);
xor U2159 (N_2159,In_483,In_636);
nand U2160 (N_2160,In_135,In_305);
or U2161 (N_2161,In_815,In_6);
or U2162 (N_2162,In_786,In_140);
nand U2163 (N_2163,In_323,In_715);
and U2164 (N_2164,In_960,In_467);
or U2165 (N_2165,In_788,In_997);
nor U2166 (N_2166,In_308,In_974);
nor U2167 (N_2167,In_443,In_620);
xor U2168 (N_2168,In_215,In_350);
and U2169 (N_2169,In_618,In_249);
nor U2170 (N_2170,In_691,In_870);
nand U2171 (N_2171,In_597,In_87);
nor U2172 (N_2172,In_194,In_736);
nand U2173 (N_2173,In_318,In_937);
or U2174 (N_2174,In_912,In_880);
or U2175 (N_2175,In_814,In_26);
or U2176 (N_2176,In_567,In_78);
and U2177 (N_2177,In_158,In_758);
or U2178 (N_2178,In_891,In_236);
nand U2179 (N_2179,In_402,In_363);
or U2180 (N_2180,In_286,In_55);
and U2181 (N_2181,In_529,In_416);
nand U2182 (N_2182,In_986,In_258);
nor U2183 (N_2183,In_363,In_110);
nor U2184 (N_2184,In_147,In_510);
nand U2185 (N_2185,In_494,In_485);
and U2186 (N_2186,In_917,In_779);
nand U2187 (N_2187,In_945,In_368);
nor U2188 (N_2188,In_895,In_557);
and U2189 (N_2189,In_932,In_344);
and U2190 (N_2190,In_303,In_391);
nand U2191 (N_2191,In_21,In_60);
and U2192 (N_2192,In_492,In_818);
or U2193 (N_2193,In_612,In_594);
nand U2194 (N_2194,In_640,In_876);
nand U2195 (N_2195,In_877,In_804);
nand U2196 (N_2196,In_691,In_241);
and U2197 (N_2197,In_248,In_382);
nor U2198 (N_2198,In_949,In_870);
nand U2199 (N_2199,In_66,In_475);
and U2200 (N_2200,In_982,In_233);
or U2201 (N_2201,In_195,In_238);
nor U2202 (N_2202,In_628,In_53);
or U2203 (N_2203,In_621,In_485);
or U2204 (N_2204,In_556,In_120);
and U2205 (N_2205,In_936,In_995);
or U2206 (N_2206,In_628,In_147);
or U2207 (N_2207,In_164,In_933);
and U2208 (N_2208,In_179,In_962);
nand U2209 (N_2209,In_918,In_41);
and U2210 (N_2210,In_859,In_501);
nand U2211 (N_2211,In_747,In_421);
and U2212 (N_2212,In_373,In_119);
and U2213 (N_2213,In_157,In_733);
nand U2214 (N_2214,In_687,In_636);
or U2215 (N_2215,In_80,In_157);
nand U2216 (N_2216,In_452,In_296);
xor U2217 (N_2217,In_36,In_348);
nand U2218 (N_2218,In_639,In_118);
and U2219 (N_2219,In_963,In_858);
nand U2220 (N_2220,In_783,In_456);
or U2221 (N_2221,In_684,In_410);
or U2222 (N_2222,In_579,In_460);
nor U2223 (N_2223,In_247,In_198);
nand U2224 (N_2224,In_460,In_664);
nand U2225 (N_2225,In_623,In_467);
or U2226 (N_2226,In_306,In_23);
or U2227 (N_2227,In_94,In_697);
or U2228 (N_2228,In_135,In_108);
nor U2229 (N_2229,In_345,In_40);
and U2230 (N_2230,In_496,In_676);
nor U2231 (N_2231,In_3,In_515);
nand U2232 (N_2232,In_649,In_558);
and U2233 (N_2233,In_79,In_255);
nand U2234 (N_2234,In_272,In_201);
nand U2235 (N_2235,In_440,In_785);
and U2236 (N_2236,In_752,In_7);
and U2237 (N_2237,In_10,In_228);
and U2238 (N_2238,In_26,In_800);
nand U2239 (N_2239,In_836,In_423);
or U2240 (N_2240,In_208,In_11);
or U2241 (N_2241,In_232,In_947);
nor U2242 (N_2242,In_474,In_399);
and U2243 (N_2243,In_686,In_880);
nor U2244 (N_2244,In_673,In_905);
nand U2245 (N_2245,In_613,In_65);
nand U2246 (N_2246,In_974,In_868);
and U2247 (N_2247,In_738,In_490);
and U2248 (N_2248,In_668,In_777);
xor U2249 (N_2249,In_617,In_205);
and U2250 (N_2250,In_301,In_111);
nor U2251 (N_2251,In_438,In_82);
nor U2252 (N_2252,In_345,In_616);
and U2253 (N_2253,In_953,In_830);
nand U2254 (N_2254,In_388,In_831);
and U2255 (N_2255,In_741,In_608);
nor U2256 (N_2256,In_589,In_304);
nand U2257 (N_2257,In_103,In_69);
nand U2258 (N_2258,In_40,In_918);
and U2259 (N_2259,In_219,In_348);
nand U2260 (N_2260,In_112,In_569);
and U2261 (N_2261,In_24,In_273);
nand U2262 (N_2262,In_827,In_390);
or U2263 (N_2263,In_561,In_807);
nor U2264 (N_2264,In_906,In_731);
or U2265 (N_2265,In_27,In_49);
and U2266 (N_2266,In_490,In_832);
and U2267 (N_2267,In_596,In_46);
or U2268 (N_2268,In_119,In_456);
or U2269 (N_2269,In_280,In_931);
nand U2270 (N_2270,In_854,In_872);
and U2271 (N_2271,In_249,In_866);
nor U2272 (N_2272,In_358,In_646);
and U2273 (N_2273,In_466,In_936);
and U2274 (N_2274,In_515,In_452);
nor U2275 (N_2275,In_925,In_337);
or U2276 (N_2276,In_209,In_3);
and U2277 (N_2277,In_955,In_606);
or U2278 (N_2278,In_736,In_264);
and U2279 (N_2279,In_416,In_609);
nand U2280 (N_2280,In_297,In_25);
or U2281 (N_2281,In_755,In_142);
nand U2282 (N_2282,In_345,In_839);
nor U2283 (N_2283,In_418,In_466);
or U2284 (N_2284,In_610,In_564);
or U2285 (N_2285,In_209,In_877);
nor U2286 (N_2286,In_879,In_300);
and U2287 (N_2287,In_747,In_184);
and U2288 (N_2288,In_129,In_213);
nand U2289 (N_2289,In_433,In_827);
nor U2290 (N_2290,In_607,In_524);
or U2291 (N_2291,In_497,In_482);
or U2292 (N_2292,In_954,In_916);
nor U2293 (N_2293,In_610,In_409);
and U2294 (N_2294,In_397,In_394);
or U2295 (N_2295,In_623,In_654);
nand U2296 (N_2296,In_282,In_246);
nand U2297 (N_2297,In_115,In_958);
nand U2298 (N_2298,In_907,In_313);
nand U2299 (N_2299,In_317,In_780);
and U2300 (N_2300,In_755,In_909);
nand U2301 (N_2301,In_700,In_480);
nand U2302 (N_2302,In_146,In_66);
nand U2303 (N_2303,In_367,In_127);
and U2304 (N_2304,In_653,In_72);
nand U2305 (N_2305,In_505,In_266);
or U2306 (N_2306,In_974,In_366);
nand U2307 (N_2307,In_656,In_998);
nor U2308 (N_2308,In_441,In_695);
nand U2309 (N_2309,In_790,In_812);
nand U2310 (N_2310,In_472,In_527);
nand U2311 (N_2311,In_346,In_647);
or U2312 (N_2312,In_957,In_928);
or U2313 (N_2313,In_55,In_351);
nor U2314 (N_2314,In_821,In_982);
or U2315 (N_2315,In_184,In_140);
nand U2316 (N_2316,In_362,In_44);
or U2317 (N_2317,In_656,In_205);
nand U2318 (N_2318,In_796,In_679);
nand U2319 (N_2319,In_648,In_769);
nor U2320 (N_2320,In_356,In_374);
nand U2321 (N_2321,In_300,In_924);
or U2322 (N_2322,In_702,In_440);
and U2323 (N_2323,In_117,In_176);
nor U2324 (N_2324,In_266,In_549);
nand U2325 (N_2325,In_547,In_757);
nand U2326 (N_2326,In_398,In_160);
nor U2327 (N_2327,In_736,In_946);
or U2328 (N_2328,In_743,In_713);
nand U2329 (N_2329,In_714,In_746);
nor U2330 (N_2330,In_770,In_798);
and U2331 (N_2331,In_867,In_332);
and U2332 (N_2332,In_473,In_597);
nor U2333 (N_2333,In_73,In_931);
or U2334 (N_2334,In_519,In_678);
nand U2335 (N_2335,In_308,In_328);
nor U2336 (N_2336,In_896,In_838);
and U2337 (N_2337,In_531,In_57);
and U2338 (N_2338,In_530,In_622);
and U2339 (N_2339,In_386,In_869);
nand U2340 (N_2340,In_58,In_675);
nor U2341 (N_2341,In_496,In_883);
and U2342 (N_2342,In_717,In_864);
or U2343 (N_2343,In_538,In_753);
and U2344 (N_2344,In_569,In_642);
and U2345 (N_2345,In_212,In_153);
nand U2346 (N_2346,In_876,In_504);
and U2347 (N_2347,In_108,In_775);
nand U2348 (N_2348,In_380,In_691);
or U2349 (N_2349,In_779,In_656);
and U2350 (N_2350,In_22,In_94);
nand U2351 (N_2351,In_465,In_476);
nor U2352 (N_2352,In_180,In_706);
nand U2353 (N_2353,In_314,In_363);
nor U2354 (N_2354,In_737,In_847);
and U2355 (N_2355,In_309,In_910);
and U2356 (N_2356,In_105,In_964);
nand U2357 (N_2357,In_82,In_695);
nor U2358 (N_2358,In_867,In_630);
nand U2359 (N_2359,In_530,In_294);
and U2360 (N_2360,In_199,In_740);
nor U2361 (N_2361,In_794,In_797);
nor U2362 (N_2362,In_548,In_696);
and U2363 (N_2363,In_608,In_551);
xor U2364 (N_2364,In_408,In_776);
nand U2365 (N_2365,In_642,In_502);
nand U2366 (N_2366,In_763,In_120);
nor U2367 (N_2367,In_46,In_480);
nor U2368 (N_2368,In_847,In_679);
or U2369 (N_2369,In_729,In_456);
nand U2370 (N_2370,In_891,In_125);
or U2371 (N_2371,In_460,In_211);
and U2372 (N_2372,In_582,In_731);
and U2373 (N_2373,In_599,In_451);
nand U2374 (N_2374,In_422,In_234);
and U2375 (N_2375,In_287,In_464);
and U2376 (N_2376,In_939,In_711);
or U2377 (N_2377,In_728,In_352);
nor U2378 (N_2378,In_932,In_73);
and U2379 (N_2379,In_367,In_94);
nor U2380 (N_2380,In_389,In_679);
nand U2381 (N_2381,In_108,In_680);
nor U2382 (N_2382,In_318,In_798);
nor U2383 (N_2383,In_337,In_602);
and U2384 (N_2384,In_972,In_116);
and U2385 (N_2385,In_612,In_530);
nor U2386 (N_2386,In_533,In_89);
nor U2387 (N_2387,In_228,In_828);
nand U2388 (N_2388,In_679,In_474);
nor U2389 (N_2389,In_344,In_880);
nor U2390 (N_2390,In_389,In_772);
or U2391 (N_2391,In_919,In_881);
or U2392 (N_2392,In_664,In_104);
nand U2393 (N_2393,In_842,In_737);
nand U2394 (N_2394,In_534,In_693);
nand U2395 (N_2395,In_289,In_648);
and U2396 (N_2396,In_514,In_326);
nand U2397 (N_2397,In_892,In_472);
and U2398 (N_2398,In_1,In_264);
nand U2399 (N_2399,In_393,In_243);
nand U2400 (N_2400,In_487,In_230);
nand U2401 (N_2401,In_645,In_286);
or U2402 (N_2402,In_841,In_242);
and U2403 (N_2403,In_527,In_329);
and U2404 (N_2404,In_662,In_32);
xor U2405 (N_2405,In_581,In_734);
nor U2406 (N_2406,In_155,In_809);
or U2407 (N_2407,In_218,In_416);
nor U2408 (N_2408,In_856,In_31);
and U2409 (N_2409,In_779,In_815);
and U2410 (N_2410,In_82,In_130);
nor U2411 (N_2411,In_653,In_785);
and U2412 (N_2412,In_659,In_669);
or U2413 (N_2413,In_348,In_334);
or U2414 (N_2414,In_408,In_351);
and U2415 (N_2415,In_8,In_898);
nand U2416 (N_2416,In_57,In_580);
nand U2417 (N_2417,In_591,In_631);
or U2418 (N_2418,In_593,In_937);
and U2419 (N_2419,In_577,In_317);
nor U2420 (N_2420,In_135,In_296);
and U2421 (N_2421,In_504,In_78);
or U2422 (N_2422,In_508,In_484);
nor U2423 (N_2423,In_905,In_300);
nand U2424 (N_2424,In_598,In_765);
or U2425 (N_2425,In_883,In_497);
and U2426 (N_2426,In_742,In_489);
or U2427 (N_2427,In_215,In_958);
nand U2428 (N_2428,In_337,In_135);
or U2429 (N_2429,In_576,In_95);
or U2430 (N_2430,In_59,In_340);
nand U2431 (N_2431,In_556,In_226);
nand U2432 (N_2432,In_923,In_795);
nand U2433 (N_2433,In_486,In_91);
nor U2434 (N_2434,In_742,In_36);
or U2435 (N_2435,In_624,In_782);
or U2436 (N_2436,In_916,In_156);
nor U2437 (N_2437,In_872,In_27);
xor U2438 (N_2438,In_676,In_517);
nand U2439 (N_2439,In_412,In_749);
nor U2440 (N_2440,In_339,In_153);
nor U2441 (N_2441,In_516,In_182);
and U2442 (N_2442,In_823,In_932);
nor U2443 (N_2443,In_482,In_388);
and U2444 (N_2444,In_463,In_517);
or U2445 (N_2445,In_657,In_817);
and U2446 (N_2446,In_435,In_494);
nand U2447 (N_2447,In_449,In_972);
and U2448 (N_2448,In_299,In_876);
nor U2449 (N_2449,In_958,In_512);
or U2450 (N_2450,In_7,In_36);
and U2451 (N_2451,In_232,In_504);
nor U2452 (N_2452,In_740,In_533);
and U2453 (N_2453,In_640,In_468);
nor U2454 (N_2454,In_637,In_626);
nor U2455 (N_2455,In_858,In_63);
or U2456 (N_2456,In_646,In_472);
nor U2457 (N_2457,In_855,In_333);
nor U2458 (N_2458,In_242,In_382);
nand U2459 (N_2459,In_942,In_608);
or U2460 (N_2460,In_698,In_720);
nor U2461 (N_2461,In_897,In_550);
nand U2462 (N_2462,In_998,In_469);
nand U2463 (N_2463,In_187,In_935);
nor U2464 (N_2464,In_742,In_456);
and U2465 (N_2465,In_368,In_61);
or U2466 (N_2466,In_954,In_203);
nor U2467 (N_2467,In_673,In_208);
nor U2468 (N_2468,In_22,In_904);
nand U2469 (N_2469,In_361,In_519);
nor U2470 (N_2470,In_720,In_463);
nor U2471 (N_2471,In_347,In_813);
and U2472 (N_2472,In_366,In_329);
or U2473 (N_2473,In_542,In_440);
and U2474 (N_2474,In_766,In_147);
nor U2475 (N_2475,In_279,In_399);
or U2476 (N_2476,In_960,In_434);
or U2477 (N_2477,In_54,In_767);
and U2478 (N_2478,In_43,In_63);
nand U2479 (N_2479,In_102,In_293);
and U2480 (N_2480,In_925,In_109);
or U2481 (N_2481,In_377,In_660);
nand U2482 (N_2482,In_918,In_38);
or U2483 (N_2483,In_972,In_518);
and U2484 (N_2484,In_775,In_805);
and U2485 (N_2485,In_446,In_331);
nor U2486 (N_2486,In_905,In_774);
nor U2487 (N_2487,In_328,In_341);
or U2488 (N_2488,In_696,In_395);
nand U2489 (N_2489,In_805,In_234);
or U2490 (N_2490,In_19,In_24);
or U2491 (N_2491,In_650,In_867);
nand U2492 (N_2492,In_80,In_952);
nand U2493 (N_2493,In_419,In_910);
nor U2494 (N_2494,In_108,In_144);
and U2495 (N_2495,In_271,In_934);
nand U2496 (N_2496,In_549,In_827);
or U2497 (N_2497,In_348,In_319);
nand U2498 (N_2498,In_332,In_214);
and U2499 (N_2499,In_687,In_922);
nor U2500 (N_2500,N_1139,N_611);
and U2501 (N_2501,N_2077,N_1676);
or U2502 (N_2502,N_559,N_1921);
xnor U2503 (N_2503,N_1286,N_2326);
nor U2504 (N_2504,N_1000,N_1154);
and U2505 (N_2505,N_405,N_2108);
nand U2506 (N_2506,N_1791,N_1652);
nand U2507 (N_2507,N_1929,N_667);
nor U2508 (N_2508,N_22,N_1101);
and U2509 (N_2509,N_52,N_2418);
nand U2510 (N_2510,N_1495,N_2286);
and U2511 (N_2511,N_2278,N_1811);
and U2512 (N_2512,N_929,N_679);
and U2513 (N_2513,N_2293,N_2364);
and U2514 (N_2514,N_1850,N_486);
and U2515 (N_2515,N_1093,N_2339);
or U2516 (N_2516,N_102,N_169);
nor U2517 (N_2517,N_422,N_1043);
nand U2518 (N_2518,N_469,N_355);
nor U2519 (N_2519,N_1035,N_222);
nand U2520 (N_2520,N_1959,N_189);
and U2521 (N_2521,N_1982,N_1031);
and U2522 (N_2522,N_1648,N_2375);
or U2523 (N_2523,N_696,N_1974);
xor U2524 (N_2524,N_2014,N_959);
nor U2525 (N_2525,N_2123,N_2304);
and U2526 (N_2526,N_92,N_1052);
nand U2527 (N_2527,N_1072,N_481);
and U2528 (N_2528,N_2086,N_1186);
nand U2529 (N_2529,N_556,N_121);
or U2530 (N_2530,N_376,N_60);
nor U2531 (N_2531,N_836,N_1868);
and U2532 (N_2532,N_810,N_1143);
and U2533 (N_2533,N_1026,N_726);
nand U2534 (N_2534,N_1119,N_879);
nand U2535 (N_2535,N_1025,N_2346);
or U2536 (N_2536,N_1034,N_110);
nand U2537 (N_2537,N_2206,N_203);
xor U2538 (N_2538,N_843,N_2218);
nor U2539 (N_2539,N_1231,N_821);
and U2540 (N_2540,N_1613,N_517);
nand U2541 (N_2541,N_971,N_2456);
nor U2542 (N_2542,N_2315,N_419);
and U2543 (N_2543,N_1349,N_2076);
nor U2544 (N_2544,N_744,N_673);
or U2545 (N_2545,N_501,N_2004);
nand U2546 (N_2546,N_15,N_255);
or U2547 (N_2547,N_46,N_1115);
or U2548 (N_2548,N_2089,N_1279);
or U2549 (N_2549,N_1109,N_2342);
nand U2550 (N_2550,N_1305,N_2193);
nand U2551 (N_2551,N_721,N_2397);
and U2552 (N_2552,N_1928,N_2032);
and U2553 (N_2553,N_2092,N_107);
nand U2554 (N_2554,N_860,N_916);
nand U2555 (N_2555,N_2462,N_1416);
or U2556 (N_2556,N_2121,N_973);
nor U2557 (N_2557,N_2327,N_300);
nor U2558 (N_2558,N_322,N_2195);
nand U2559 (N_2559,N_1065,N_1189);
and U2560 (N_2560,N_72,N_1359);
nand U2561 (N_2561,N_2067,N_812);
nand U2562 (N_2562,N_2330,N_990);
and U2563 (N_2563,N_566,N_2290);
and U2564 (N_2564,N_1311,N_941);
nand U2565 (N_2565,N_174,N_263);
nand U2566 (N_2566,N_2492,N_1370);
nand U2567 (N_2567,N_2249,N_1250);
or U2568 (N_2568,N_2196,N_2384);
and U2569 (N_2569,N_1263,N_934);
nand U2570 (N_2570,N_880,N_1494);
xnor U2571 (N_2571,N_506,N_1967);
nor U2572 (N_2572,N_2259,N_1661);
nand U2573 (N_2573,N_1782,N_1222);
and U2574 (N_2574,N_514,N_428);
and U2575 (N_2575,N_887,N_1457);
nand U2576 (N_2576,N_1419,N_1369);
and U2577 (N_2577,N_807,N_1789);
or U2578 (N_2578,N_440,N_1134);
or U2579 (N_2579,N_652,N_551);
nand U2580 (N_2580,N_485,N_1546);
and U2581 (N_2581,N_2372,N_2228);
nor U2582 (N_2582,N_573,N_1893);
or U2583 (N_2583,N_2145,N_988);
nor U2584 (N_2584,N_1217,N_206);
and U2585 (N_2585,N_1267,N_281);
or U2586 (N_2586,N_228,N_105);
nor U2587 (N_2587,N_2210,N_961);
and U2588 (N_2588,N_438,N_1597);
or U2589 (N_2589,N_581,N_1469);
or U2590 (N_2590,N_1174,N_1671);
nand U2591 (N_2591,N_1049,N_1752);
nand U2592 (N_2592,N_2055,N_369);
or U2593 (N_2593,N_1294,N_678);
nor U2594 (N_2594,N_1287,N_2002);
and U2595 (N_2595,N_177,N_2325);
or U2596 (N_2596,N_693,N_444);
and U2597 (N_2597,N_1721,N_301);
nand U2598 (N_2598,N_1654,N_1593);
or U2599 (N_2599,N_2017,N_1491);
nand U2600 (N_2600,N_317,N_636);
and U2601 (N_2601,N_1407,N_2157);
nand U2602 (N_2602,N_1431,N_982);
nor U2603 (N_2603,N_2178,N_85);
nor U2604 (N_2604,N_286,N_1525);
and U2605 (N_2605,N_185,N_1187);
or U2606 (N_2606,N_705,N_1575);
nor U2607 (N_2607,N_1796,N_615);
or U2608 (N_2608,N_260,N_2306);
and U2609 (N_2609,N_1740,N_2042);
and U2610 (N_2610,N_670,N_2485);
or U2611 (N_2611,N_2066,N_1596);
nor U2612 (N_2612,N_1883,N_1071);
nor U2613 (N_2613,N_2053,N_2080);
nand U2614 (N_2614,N_2352,N_1836);
nand U2615 (N_2615,N_125,N_1650);
nand U2616 (N_2616,N_1995,N_394);
and U2617 (N_2617,N_2147,N_681);
and U2618 (N_2618,N_1411,N_1427);
or U2619 (N_2619,N_2497,N_2318);
nand U2620 (N_2620,N_1647,N_1140);
and U2621 (N_2621,N_1367,N_710);
or U2622 (N_2622,N_1934,N_1832);
and U2623 (N_2623,N_802,N_1114);
and U2624 (N_2624,N_1335,N_1122);
nor U2625 (N_2625,N_1601,N_229);
nor U2626 (N_2626,N_822,N_717);
nand U2627 (N_2627,N_2487,N_1182);
and U2628 (N_2628,N_1218,N_2159);
and U2629 (N_2629,N_1646,N_1441);
nand U2630 (N_2630,N_868,N_1913);
xnor U2631 (N_2631,N_1986,N_69);
and U2632 (N_2632,N_2000,N_1410);
and U2633 (N_2633,N_799,N_427);
and U2634 (N_2634,N_1015,N_980);
and U2635 (N_2635,N_2096,N_830);
xor U2636 (N_2636,N_599,N_280);
or U2637 (N_2637,N_1787,N_1903);
nand U2638 (N_2638,N_126,N_1687);
and U2639 (N_2639,N_176,N_160);
or U2640 (N_2640,N_2124,N_743);
and U2641 (N_2641,N_460,N_2133);
nand U2642 (N_2642,N_230,N_2253);
or U2643 (N_2643,N_509,N_1664);
nand U2644 (N_2644,N_2209,N_99);
and U2645 (N_2645,N_781,N_2496);
and U2646 (N_2646,N_252,N_544);
nor U2647 (N_2647,N_77,N_2394);
nor U2648 (N_2648,N_132,N_2482);
xor U2649 (N_2649,N_1033,N_1138);
nor U2650 (N_2650,N_1537,N_128);
nand U2651 (N_2651,N_2439,N_742);
and U2652 (N_2652,N_1141,N_59);
and U2653 (N_2653,N_1777,N_1608);
nor U2654 (N_2654,N_1091,N_1164);
nor U2655 (N_2655,N_1800,N_1726);
or U2656 (N_2656,N_2460,N_212);
or U2657 (N_2657,N_97,N_1429);
nand U2658 (N_2658,N_1761,N_1762);
and U2659 (N_2659,N_1188,N_1508);
nor U2660 (N_2660,N_1935,N_313);
nand U2661 (N_2661,N_170,N_1943);
nor U2662 (N_2662,N_1492,N_2069);
or U2663 (N_2663,N_1145,N_2098);
nand U2664 (N_2664,N_454,N_1798);
nand U2665 (N_2665,N_2440,N_2225);
or U2666 (N_2666,N_1313,N_2243);
or U2667 (N_2667,N_2234,N_832);
nand U2668 (N_2668,N_841,N_2113);
nand U2669 (N_2669,N_1044,N_1497);
nor U2670 (N_2670,N_138,N_666);
nand U2671 (N_2671,N_1024,N_596);
or U2672 (N_2672,N_1634,N_2045);
nor U2673 (N_2673,N_1715,N_2305);
and U2674 (N_2674,N_1064,N_1042);
nand U2675 (N_2675,N_1340,N_870);
nor U2676 (N_2676,N_1858,N_2361);
or U2677 (N_2677,N_217,N_757);
and U2678 (N_2678,N_2090,N_1068);
nor U2679 (N_2679,N_351,N_1204);
nor U2680 (N_2680,N_299,N_2411);
nor U2681 (N_2681,N_463,N_958);
nor U2682 (N_2682,N_2469,N_274);
nor U2683 (N_2683,N_2382,N_541);
nand U2684 (N_2684,N_18,N_1892);
and U2685 (N_2685,N_42,N_1297);
nand U2686 (N_2686,N_2363,N_642);
nor U2687 (N_2687,N_1422,N_619);
and U2688 (N_2688,N_1701,N_88);
nor U2689 (N_2689,N_1126,N_1523);
nand U2690 (N_2690,N_87,N_2144);
or U2691 (N_2691,N_976,N_1315);
or U2692 (N_2692,N_1406,N_998);
nand U2693 (N_2693,N_1922,N_1957);
nand U2694 (N_2694,N_11,N_29);
and U2695 (N_2695,N_1307,N_633);
nand U2696 (N_2696,N_828,N_1048);
or U2697 (N_2697,N_901,N_1057);
nor U2698 (N_2698,N_760,N_1301);
nor U2699 (N_2699,N_1628,N_1554);
and U2700 (N_2700,N_2205,N_2186);
and U2701 (N_2701,N_1309,N_1919);
or U2702 (N_2702,N_395,N_1861);
and U2703 (N_2703,N_1496,N_2387);
and U2704 (N_2704,N_312,N_1124);
nand U2705 (N_2705,N_159,N_1388);
or U2706 (N_2706,N_1036,N_25);
or U2707 (N_2707,N_1321,N_50);
nand U2708 (N_2708,N_1442,N_964);
nor U2709 (N_2709,N_1285,N_656);
or U2710 (N_2710,N_1172,N_186);
and U2711 (N_2711,N_133,N_1585);
nand U2712 (N_2712,N_716,N_1978);
nand U2713 (N_2713,N_2283,N_644);
and U2714 (N_2714,N_967,N_1105);
and U2715 (N_2715,N_68,N_1481);
nor U2716 (N_2716,N_104,N_1066);
nand U2717 (N_2717,N_1353,N_302);
nand U2718 (N_2718,N_946,N_856);
or U2719 (N_2719,N_1606,N_279);
and U2720 (N_2720,N_2356,N_2480);
nor U2721 (N_2721,N_2208,N_2321);
nor U2722 (N_2722,N_2065,N_1845);
nor U2723 (N_2723,N_2493,N_1260);
or U2724 (N_2724,N_324,N_1907);
or U2725 (N_2725,N_1630,N_1629);
or U2726 (N_2726,N_1021,N_466);
nor U2727 (N_2727,N_411,N_1941);
or U2728 (N_2728,N_724,N_753);
nand U2729 (N_2729,N_381,N_1955);
nand U2730 (N_2730,N_2282,N_917);
nor U2731 (N_2731,N_2192,N_1149);
and U2732 (N_2732,N_984,N_1853);
or U2733 (N_2733,N_2110,N_2250);
and U2734 (N_2734,N_1830,N_1135);
nor U2735 (N_2735,N_477,N_198);
nand U2736 (N_2736,N_926,N_494);
and U2737 (N_2737,N_2051,N_1703);
nor U2738 (N_2738,N_1567,N_920);
or U2739 (N_2739,N_1932,N_2162);
and U2740 (N_2740,N_1743,N_2132);
and U2741 (N_2741,N_801,N_2189);
and U2742 (N_2742,N_2454,N_819);
or U2743 (N_2743,N_2434,N_348);
or U2744 (N_2744,N_1750,N_1272);
or U2745 (N_2745,N_2166,N_2430);
or U2746 (N_2746,N_2248,N_855);
or U2747 (N_2747,N_1656,N_284);
xor U2748 (N_2748,N_1001,N_2498);
or U2749 (N_2749,N_928,N_1700);
nand U2750 (N_2750,N_730,N_2095);
nand U2751 (N_2751,N_831,N_1591);
and U2752 (N_2752,N_144,N_344);
nor U2753 (N_2753,N_145,N_40);
xnor U2754 (N_2754,N_650,N_790);
or U2755 (N_2755,N_2395,N_2422);
nor U2756 (N_2756,N_776,N_1478);
or U2757 (N_2757,N_1960,N_334);
or U2758 (N_2758,N_1560,N_2393);
and U2759 (N_2759,N_1851,N_937);
nor U2760 (N_2760,N_1289,N_1350);
nor U2761 (N_2761,N_1237,N_1310);
xnor U2762 (N_2762,N_242,N_1563);
nor U2763 (N_2763,N_413,N_1151);
nand U2764 (N_2764,N_1163,N_1631);
nand U2765 (N_2765,N_1856,N_2255);
nand U2766 (N_2766,N_2258,N_1724);
nand U2767 (N_2767,N_1773,N_1007);
or U2768 (N_2768,N_960,N_881);
or U2769 (N_2769,N_1621,N_180);
and U2770 (N_2770,N_2217,N_453);
and U2771 (N_2771,N_588,N_2235);
and U2772 (N_2772,N_1709,N_752);
or U2773 (N_2773,N_357,N_1480);
xor U2774 (N_2774,N_649,N_2345);
nand U2775 (N_2775,N_1067,N_375);
or U2776 (N_2776,N_2115,N_2219);
and U2777 (N_2777,N_2062,N_1860);
or U2778 (N_2778,N_979,N_2221);
nand U2779 (N_2779,N_1998,N_362);
nand U2780 (N_2780,N_2368,N_291);
nand U2781 (N_2781,N_1840,N_1873);
and U2782 (N_2782,N_335,N_2336);
or U2783 (N_2783,N_2379,N_1206);
nand U2784 (N_2784,N_241,N_2030);
and U2785 (N_2785,N_2262,N_1888);
nor U2786 (N_2786,N_808,N_2371);
nor U2787 (N_2787,N_844,N_1805);
nor U2788 (N_2788,N_2458,N_1938);
xnor U2789 (N_2789,N_1233,N_646);
and U2790 (N_2790,N_780,N_1516);
or U2791 (N_2791,N_864,N_1622);
and U2792 (N_2792,N_1396,N_519);
nand U2793 (N_2793,N_202,N_1637);
and U2794 (N_2794,N_755,N_2489);
or U2795 (N_2795,N_1522,N_1341);
nand U2796 (N_2796,N_2486,N_641);
or U2797 (N_2797,N_311,N_793);
nor U2798 (N_2798,N_2229,N_1318);
nand U2799 (N_2799,N_1268,N_316);
nor U2800 (N_2800,N_1747,N_306);
and U2801 (N_2801,N_1612,N_482);
nor U2802 (N_2802,N_2310,N_797);
nand U2803 (N_2803,N_545,N_648);
and U2804 (N_2804,N_2285,N_285);
or U2805 (N_2805,N_476,N_2349);
nand U2806 (N_2806,N_788,N_1061);
or U2807 (N_2807,N_2129,N_238);
and U2808 (N_2808,N_2187,N_1574);
and U2809 (N_2809,N_10,N_1925);
or U2810 (N_2810,N_2347,N_1870);
or U2811 (N_2811,N_402,N_707);
or U2812 (N_2812,N_2294,N_1060);
or U2813 (N_2813,N_1504,N_912);
and U2814 (N_2814,N_806,N_1463);
nor U2815 (N_2815,N_379,N_507);
and U2816 (N_2816,N_1299,N_1990);
nand U2817 (N_2817,N_2022,N_607);
nor U2818 (N_2818,N_1714,N_834);
nand U2819 (N_2819,N_669,N_91);
nand U2820 (N_2820,N_1110,N_1981);
nand U2821 (N_2821,N_643,N_1550);
or U2822 (N_2822,N_2275,N_248);
or U2823 (N_2823,N_249,N_1519);
nor U2824 (N_2824,N_722,N_1937);
and U2825 (N_2825,N_2391,N_1282);
and U2826 (N_2826,N_2260,N_1618);
nand U2827 (N_2827,N_1723,N_268);
and U2828 (N_2828,N_2455,N_1930);
xor U2829 (N_2829,N_784,N_554);
and U2830 (N_2830,N_2023,N_626);
nand U2831 (N_2831,N_835,N_2010);
nand U2832 (N_2832,N_1449,N_2024);
and U2833 (N_2833,N_1768,N_2466);
and U2834 (N_2834,N_2064,N_2463);
nand U2835 (N_2835,N_1243,N_2451);
and U2836 (N_2836,N_1423,N_2152);
nor U2837 (N_2837,N_449,N_1090);
and U2838 (N_2838,N_2146,N_2385);
or U2839 (N_2839,N_1733,N_731);
nand U2840 (N_2840,N_421,N_1939);
or U2841 (N_2841,N_1357,N_2274);
or U2842 (N_2842,N_1694,N_1384);
or U2843 (N_2843,N_2019,N_14);
nor U2844 (N_2844,N_325,N_2331);
nor U2845 (N_2845,N_1663,N_1566);
nand U2846 (N_2846,N_1765,N_41);
and U2847 (N_2847,N_1440,N_533);
nor U2848 (N_2848,N_927,N_711);
nand U2849 (N_2849,N_385,N_1707);
or U2850 (N_2850,N_245,N_1588);
and U2851 (N_2851,N_188,N_106);
nand U2852 (N_2852,N_617,N_898);
nand U2853 (N_2853,N_272,N_1535);
and U2854 (N_2854,N_567,N_1843);
or U2855 (N_2855,N_1728,N_1878);
or U2856 (N_2856,N_829,N_1354);
or U2857 (N_2857,N_2029,N_137);
or U2858 (N_2858,N_497,N_1404);
or U2859 (N_2859,N_161,N_388);
and U2860 (N_2860,N_127,N_1215);
and U2861 (N_2861,N_558,N_1711);
and U2862 (N_2862,N_2426,N_1437);
or U2863 (N_2863,N_356,N_179);
nor U2864 (N_2864,N_1326,N_1316);
nor U2865 (N_2865,N_384,N_900);
nor U2866 (N_2866,N_1680,N_1727);
nor U2867 (N_2867,N_1436,N_1632);
nor U2868 (N_2868,N_604,N_515);
nand U2869 (N_2869,N_546,N_1118);
nor U2870 (N_2870,N_1541,N_972);
nor U2871 (N_2871,N_103,N_1261);
nand U2872 (N_2872,N_1039,N_459);
and U2873 (N_2873,N_2329,N_1660);
nor U2874 (N_2874,N_602,N_2226);
nand U2875 (N_2875,N_2158,N_783);
or U2876 (N_2876,N_2403,N_932);
nor U2877 (N_2877,N_450,N_1275);
and U2878 (N_2878,N_2081,N_2165);
nand U2879 (N_2879,N_2273,N_205);
nor U2880 (N_2880,N_2443,N_863);
and U2881 (N_2881,N_2168,N_761);
and U2882 (N_2882,N_1842,N_1414);
nand U2883 (N_2883,N_1202,N_1512);
or U2884 (N_2884,N_1100,N_913);
and U2885 (N_2885,N_845,N_2070);
or U2886 (N_2886,N_2340,N_1337);
nand U2887 (N_2887,N_2276,N_942);
or U2888 (N_2888,N_234,N_1710);
or U2889 (N_2889,N_2164,N_2314);
and U2890 (N_2890,N_1692,N_1984);
nand U2891 (N_2891,N_847,N_2016);
nand U2892 (N_2892,N_1940,N_814);
nor U2893 (N_2893,N_1116,N_2223);
nor U2894 (N_2894,N_1882,N_1584);
or U2895 (N_2895,N_1230,N_309);
and U2896 (N_2896,N_2204,N_1155);
or U2897 (N_2897,N_2130,N_1371);
and U2898 (N_2898,N_593,N_434);
nor U2899 (N_2899,N_310,N_1586);
and U2900 (N_2900,N_1417,N_2453);
or U2901 (N_2901,N_1615,N_474);
nand U2902 (N_2902,N_1214,N_1327);
and U2903 (N_2903,N_2377,N_1605);
nor U2904 (N_2904,N_952,N_2362);
xnor U2905 (N_2905,N_2406,N_1815);
or U2906 (N_2906,N_1078,N_739);
and U2907 (N_2907,N_1019,N_1885);
nor U2908 (N_2908,N_1177,N_141);
nor U2909 (N_2909,N_2118,N_473);
and U2910 (N_2910,N_1844,N_2200);
nand U2911 (N_2911,N_2061,N_452);
nor U2912 (N_2912,N_1308,N_1557);
and U2913 (N_2913,N_1399,N_713);
and U2914 (N_2914,N_516,N_1665);
nor U2915 (N_2915,N_1686,N_2107);
nor U2916 (N_2916,N_2236,N_1894);
or U2917 (N_2917,N_258,N_603);
and U2918 (N_2918,N_1533,N_622);
and U2919 (N_2919,N_1526,N_795);
nor U2920 (N_2920,N_1636,N_684);
or U2921 (N_2921,N_1089,N_1659);
nand U2922 (N_2922,N_1344,N_904);
or U2923 (N_2923,N_433,N_2308);
nand U2924 (N_2924,N_813,N_1846);
and U2925 (N_2925,N_2307,N_872);
and U2926 (N_2926,N_2049,N_1424);
or U2927 (N_2927,N_1833,N_425);
and U2928 (N_2928,N_1292,N_664);
or U2929 (N_2929,N_1381,N_1642);
nor U2930 (N_2930,N_2074,N_1010);
or U2931 (N_2931,N_383,N_233);
and U2932 (N_2932,N_674,N_1295);
nand U2933 (N_2933,N_45,N_512);
nor U2934 (N_2934,N_1054,N_1988);
or U2935 (N_2935,N_1531,N_1510);
and U2936 (N_2936,N_475,N_1806);
or U2937 (N_2937,N_1573,N_2039);
nand U2938 (N_2938,N_1320,N_2323);
nand U2939 (N_2939,N_1073,N_1786);
or U2940 (N_2940,N_2142,N_254);
or U2941 (N_2941,N_572,N_995);
nand U2942 (N_2942,N_1253,N_2150);
nor U2943 (N_2943,N_1319,N_2190);
and U2944 (N_2944,N_1259,N_680);
or U2945 (N_2945,N_2091,N_1587);
or U2946 (N_2946,N_38,N_216);
nor U2947 (N_2947,N_314,N_271);
nand U2948 (N_2948,N_1972,N_1120);
nand U2949 (N_2949,N_727,N_108);
nor U2950 (N_2950,N_1390,N_756);
or U2951 (N_2951,N_1975,N_56);
or U2952 (N_2952,N_530,N_800);
nor U2953 (N_2953,N_70,N_253);
nand U2954 (N_2954,N_2112,N_247);
nor U2955 (N_2955,N_909,N_577);
nor U2956 (N_2956,N_82,N_1799);
nor U2957 (N_2957,N_115,N_2043);
and U2958 (N_2958,N_1997,N_1592);
nand U2959 (N_2959,N_2141,N_297);
and U2960 (N_2960,N_214,N_2483);
nor U2961 (N_2961,N_2139,N_1132);
and U2962 (N_2962,N_1343,N_367);
nor U2963 (N_2963,N_1070,N_2052);
nand U2964 (N_2964,N_1616,N_1183);
nor U2965 (N_2965,N_548,N_2438);
and U2966 (N_2966,N_1831,N_1047);
or U2967 (N_2967,N_1809,N_1581);
nor U2968 (N_2968,N_955,N_1949);
and U2969 (N_2969,N_1756,N_719);
nand U2970 (N_2970,N_1037,N_1336);
nor U2971 (N_2971,N_2338,N_1966);
and U2972 (N_2972,N_223,N_598);
nand U2973 (N_2973,N_1241,N_1763);
and U2974 (N_2974,N_1524,N_2244);
and U2975 (N_2975,N_439,N_275);
nand U2976 (N_2976,N_237,N_1857);
and U2977 (N_2977,N_1046,N_2003);
or U2978 (N_2978,N_2311,N_1559);
or U2979 (N_2979,N_1102,N_308);
nor U2980 (N_2980,N_227,N_2058);
nand U2981 (N_2981,N_2419,N_889);
nor U2982 (N_2982,N_627,N_677);
or U2983 (N_2983,N_2215,N_358);
nand U2984 (N_2984,N_798,N_2399);
nand U2985 (N_2985,N_1705,N_1590);
nand U2986 (N_2986,N_1178,N_590);
nor U2987 (N_2987,N_49,N_1617);
or U2988 (N_2988,N_470,N_2442);
or U2989 (N_2989,N_1804,N_584);
and U2990 (N_2990,N_1079,N_2271);
nand U2991 (N_2991,N_374,N_1987);
nand U2992 (N_2992,N_827,N_747);
nor U2993 (N_2993,N_580,N_1041);
nand U2994 (N_2994,N_2,N_1216);
and U2995 (N_2995,N_1964,N_158);
and U2996 (N_2996,N_2001,N_542);
nor U2997 (N_2997,N_1103,N_1273);
or U2998 (N_2998,N_98,N_1780);
or U2999 (N_2999,N_1438,N_815);
nor U3000 (N_3000,N_1002,N_436);
and U3001 (N_3001,N_2474,N_44);
nand U3002 (N_3002,N_163,N_733);
or U3003 (N_3003,N_2170,N_741);
nor U3004 (N_3004,N_1127,N_999);
and U3005 (N_3005,N_859,N_147);
and U3006 (N_3006,N_277,N_592);
nand U3007 (N_3007,N_1142,N_329);
nor U3008 (N_3008,N_526,N_991);
nor U3009 (N_3009,N_172,N_1144);
or U3010 (N_3010,N_414,N_1509);
nor U3011 (N_3011,N_1754,N_1755);
nand U3012 (N_3012,N_1439,N_1028);
nor U3013 (N_3013,N_574,N_1130);
or U3014 (N_3014,N_1099,N_1589);
and U3015 (N_3015,N_1402,N_771);
and U3016 (N_3016,N_640,N_754);
nand U3017 (N_3017,N_1758,N_304);
and U3018 (N_3018,N_2180,N_1389);
nand U3019 (N_3019,N_2301,N_1245);
and U3020 (N_3020,N_2446,N_465);
or U3021 (N_3021,N_1225,N_616);
nor U3022 (N_3022,N_1985,N_2357);
nor U3023 (N_3023,N_1415,N_489);
or U3024 (N_3024,N_511,N_1916);
or U3025 (N_3025,N_9,N_1459);
nor U3026 (N_3026,N_521,N_625);
nand U3027 (N_3027,N_890,N_1822);
nand U3028 (N_3028,N_1785,N_171);
nand U3029 (N_3029,N_2034,N_360);
and U3030 (N_3030,N_232,N_155);
or U3031 (N_3031,N_373,N_430);
nor U3032 (N_3032,N_2179,N_1810);
nor U3033 (N_3033,N_1201,N_1625);
nand U3034 (N_3034,N_1500,N_2490);
nand U3035 (N_3035,N_759,N_488);
nand U3036 (N_3036,N_2026,N_1108);
and U3037 (N_3037,N_173,N_1266);
or U3038 (N_3038,N_2174,N_921);
xor U3039 (N_3039,N_1848,N_219);
nand U3040 (N_3040,N_2280,N_215);
nor U3041 (N_3041,N_1433,N_493);
and U3042 (N_3042,N_1718,N_1970);
and U3043 (N_3043,N_1244,N_2432);
and U3044 (N_3044,N_340,N_1197);
nand U3045 (N_3045,N_181,N_153);
nor U3046 (N_3046,N_490,N_936);
nor U3047 (N_3047,N_2299,N_867);
and U3048 (N_3048,N_79,N_1129);
and U3049 (N_3049,N_1083,N_1479);
and U3050 (N_3050,N_1869,N_67);
nand U3051 (N_3051,N_492,N_1450);
or U3052 (N_3052,N_1651,N_1018);
or U3053 (N_3053,N_1540,N_398);
and U3054 (N_3054,N_1377,N_1672);
nand U3055 (N_3055,N_2104,N_939);
and U3056 (N_3056,N_1871,N_1195);
or U3057 (N_3057,N_287,N_957);
nand U3058 (N_3058,N_2435,N_2005);
nor U3059 (N_3059,N_694,N_1558);
nand U3060 (N_3060,N_1051,N_495);
nor U3061 (N_3061,N_1505,N_2351);
and U3062 (N_3062,N_539,N_849);
nand U3063 (N_3063,N_1849,N_1136);
or U3064 (N_3064,N_2279,N_532);
xnor U3065 (N_3065,N_1173,N_1322);
nand U3066 (N_3066,N_894,N_2400);
or U3067 (N_3067,N_2428,N_907);
and U3068 (N_3068,N_2102,N_266);
or U3069 (N_3069,N_2128,N_969);
nor U3070 (N_3070,N_480,N_2436);
nor U3071 (N_3071,N_1466,N_1859);
nand U3072 (N_3072,N_565,N_371);
and U3073 (N_3073,N_1801,N_168);
nor U3074 (N_3074,N_458,N_1578);
or U3075 (N_3075,N_536,N_662);
nand U3076 (N_3076,N_2136,N_2122);
nor U3077 (N_3077,N_579,N_1600);
nor U3078 (N_3078,N_165,N_1838);
nor U3079 (N_3079,N_1689,N_122);
nand U3080 (N_3080,N_632,N_140);
nand U3081 (N_3081,N_1973,N_2185);
nor U3082 (N_3082,N_1994,N_35);
nand U3083 (N_3083,N_143,N_1738);
nand U3084 (N_3084,N_1876,N_1556);
or U3085 (N_3085,N_1852,N_902);
nor U3086 (N_3086,N_639,N_978);
or U3087 (N_3087,N_1482,N_1161);
nand U3088 (N_3088,N_471,N_209);
and U3089 (N_3089,N_2257,N_763);
nand U3090 (N_3090,N_2407,N_1221);
xnor U3091 (N_3091,N_1329,N_142);
nand U3092 (N_3092,N_2389,N_1148);
or U3093 (N_3093,N_989,N_853);
nor U3094 (N_3094,N_528,N_318);
and U3095 (N_3095,N_1212,N_750);
nor U3096 (N_3096,N_804,N_396);
or U3097 (N_3097,N_1640,N_1426);
or U3098 (N_3098,N_1168,N_1082);
nand U3099 (N_3099,N_748,N_1739);
nor U3100 (N_3100,N_191,N_1317);
nor U3101 (N_3101,N_187,N_956);
nand U3102 (N_3102,N_23,N_1477);
nor U3103 (N_3103,N_1264,N_1004);
nor U3104 (N_3104,N_562,N_1977);
nand U3105 (N_3105,N_1382,N_100);
nand U3106 (N_3106,N_1699,N_337);
nor U3107 (N_3107,N_723,N_861);
nor U3108 (N_3108,N_1513,N_2127);
or U3109 (N_3109,N_1468,N_663);
or U3110 (N_3110,N_1641,N_688);
and U3111 (N_3111,N_1199,N_2059);
or U3112 (N_3112,N_2231,N_1391);
nand U3113 (N_3113,N_1125,N_930);
nor U3114 (N_3114,N_20,N_2175);
nor U3115 (N_3115,N_996,N_702);
nor U3116 (N_3116,N_1794,N_17);
nor U3117 (N_3117,N_791,N_2203);
and U3118 (N_3118,N_184,N_1901);
or U3119 (N_3119,N_1834,N_403);
and U3120 (N_3120,N_659,N_1395);
nand U3121 (N_3121,N_57,N_354);
or U3122 (N_3122,N_1770,N_897);
nand U3123 (N_3123,N_1053,N_1824);
and U3124 (N_3124,N_1874,N_2383);
and U3125 (N_3125,N_2008,N_151);
or U3126 (N_3126,N_1887,N_1555);
nor U3127 (N_3127,N_2367,N_211);
nor U3128 (N_3128,N_2060,N_1484);
nand U3129 (N_3129,N_871,N_257);
or U3130 (N_3130,N_1895,N_605);
nor U3131 (N_3131,N_657,N_1249);
nand U3132 (N_3132,N_1029,N_1485);
nand U3133 (N_3133,N_2335,N_51);
or U3134 (N_3134,N_2046,N_2036);
or U3135 (N_3135,N_1570,N_1160);
and U3136 (N_3136,N_89,N_1989);
nor U3137 (N_3137,N_1198,N_1069);
nand U3138 (N_3138,N_668,N_483);
or U3139 (N_3139,N_692,N_1633);
nor U3140 (N_3140,N_326,N_363);
or U3141 (N_3141,N_148,N_2025);
and U3142 (N_3142,N_676,N_2020);
or U3143 (N_3143,N_869,N_840);
or U3144 (N_3144,N_2073,N_2343);
nor U3145 (N_3145,N_838,N_415);
nor U3146 (N_3146,N_1400,N_613);
or U3147 (N_3147,N_1247,N_2267);
and U3148 (N_3148,N_2057,N_349);
nor U3149 (N_3149,N_1814,N_130);
or U3150 (N_3150,N_1331,N_409);
nor U3151 (N_3151,N_2298,N_1022);
nor U3152 (N_3152,N_2097,N_1062);
nand U3153 (N_3153,N_1507,N_854);
nor U3154 (N_3154,N_1312,N_1226);
or U3155 (N_3155,N_1936,N_1175);
or U3156 (N_3156,N_1889,N_850);
or U3157 (N_3157,N_950,N_903);
nand U3158 (N_3158,N_1050,N_1708);
and U3159 (N_3159,N_36,N_412);
nor U3160 (N_3160,N_1674,N_83);
or U3161 (N_3161,N_1345,N_74);
nor U3162 (N_3162,N_706,N_1228);
or U3163 (N_3163,N_377,N_895);
or U3164 (N_3164,N_2083,N_1807);
or U3165 (N_3165,N_261,N_635);
nor U3166 (N_3166,N_387,N_442);
nor U3167 (N_3167,N_1368,N_1194);
and U3168 (N_3168,N_1854,N_1094);
nand U3169 (N_3169,N_1948,N_392);
or U3170 (N_3170,N_1950,N_1448);
nand U3171 (N_3171,N_332,N_614);
or U3172 (N_3172,N_2100,N_732);
nor U3173 (N_3173,N_352,N_1983);
nand U3174 (N_3174,N_282,N_1639);
nand U3175 (N_3175,N_905,N_661);
or U3176 (N_3176,N_30,N_728);
nand U3177 (N_3177,N_769,N_1224);
or U3178 (N_3178,N_2354,N_3);
or U3179 (N_3179,N_1428,N_1915);
or U3180 (N_3180,N_2360,N_1162);
nor U3181 (N_3181,N_2319,N_472);
nor U3182 (N_3182,N_298,N_2181);
or U3183 (N_3183,N_196,N_61);
or U3184 (N_3184,N_1363,N_2182);
or U3185 (N_3185,N_368,N_1460);
nor U3186 (N_3186,N_114,N_518);
or U3187 (N_3187,N_1432,N_685);
nor U3188 (N_3188,N_923,N_1819);
or U3189 (N_3189,N_1339,N_66);
or U3190 (N_3190,N_865,N_975);
and U3191 (N_3191,N_2072,N_2194);
nand U3192 (N_3192,N_1547,N_1527);
or U3193 (N_3193,N_523,N_1920);
or U3194 (N_3194,N_729,N_1536);
nor U3195 (N_3195,N_774,N_1398);
and U3196 (N_3196,N_970,N_1355);
and U3197 (N_3197,N_1751,N_1553);
nor U3198 (N_3198,N_1795,N_1802);
nor U3199 (N_3199,N_2353,N_120);
nor U3200 (N_3200,N_908,N_305);
or U3201 (N_3201,N_461,N_1486);
and U3202 (N_3202,N_350,N_1776);
nor U3203 (N_3203,N_1569,N_2452);
and U3204 (N_3204,N_2447,N_448);
nand U3205 (N_3205,N_687,N_924);
nor U3206 (N_3206,N_455,N_1684);
or U3207 (N_3207,N_820,N_2071);
or U3208 (N_3208,N_1487,N_1521);
or U3209 (N_3209,N_178,N_119);
or U3210 (N_3210,N_204,N_1465);
or U3211 (N_3211,N_164,N_1734);
or U3212 (N_3212,N_1284,N_235);
and U3213 (N_3213,N_71,N_1475);
and U3214 (N_3214,N_167,N_197);
or U3215 (N_3215,N_2103,N_117);
nand U3216 (N_3216,N_1619,N_500);
or U3217 (N_3217,N_1330,N_1991);
or U3218 (N_3218,N_2094,N_1157);
nor U3219 (N_3219,N_583,N_1467);
nand U3220 (N_3220,N_2358,N_1270);
nand U3221 (N_3221,N_1627,N_1678);
nor U3222 (N_3222,N_224,N_1111);
or U3223 (N_3223,N_818,N_527);
and U3224 (N_3224,N_2241,N_2084);
nor U3225 (N_3225,N_262,N_1302);
nor U3226 (N_3226,N_1488,N_977);
nand U3227 (N_3227,N_608,N_1325);
nand U3228 (N_3228,N_2481,N_2240);
and U3229 (N_3229,N_862,N_2207);
or U3230 (N_3230,N_1693,N_944);
nand U3231 (N_3231,N_1107,N_1013);
nand U3232 (N_3232,N_372,N_239);
nor U3233 (N_3233,N_2048,N_504);
or U3234 (N_3234,N_131,N_1385);
or U3235 (N_3235,N_2370,N_1274);
and U3236 (N_3236,N_606,N_112);
nand U3237 (N_3237,N_2188,N_1595);
nor U3238 (N_3238,N_2238,N_1);
nand U3239 (N_3239,N_885,N_2264);
or U3240 (N_3240,N_1180,N_2461);
or U3241 (N_3241,N_1005,N_2263);
and U3242 (N_3242,N_1645,N_782);
or U3243 (N_3243,N_1897,N_2239);
nand U3244 (N_3244,N_2459,N_424);
and U3245 (N_3245,N_81,N_1695);
nand U3246 (N_3246,N_962,N_1087);
nand U3247 (N_3247,N_2355,N_296);
or U3248 (N_3248,N_531,N_1232);
or U3249 (N_3249,N_1203,N_540);
nor U3250 (N_3250,N_1112,N_839);
or U3251 (N_3251,N_1670,N_2465);
nand U3252 (N_3252,N_824,N_1435);
and U3253 (N_3253,N_1918,N_1303);
or U3254 (N_3254,N_1683,N_193);
or U3255 (N_3255,N_1564,N_1511);
and U3256 (N_3256,N_1405,N_1020);
or U3257 (N_3257,N_1610,N_464);
and U3258 (N_3258,N_1011,N_883);
or U3259 (N_3259,N_162,N_2341);
or U3260 (N_3260,N_1200,N_1582);
nor U3261 (N_3261,N_1702,N_2126);
nor U3262 (N_3262,N_1835,N_1378);
or U3263 (N_3263,N_1529,N_346);
and U3264 (N_3264,N_382,N_1153);
nor U3265 (N_3265,N_2153,N_2012);
nor U3266 (N_3266,N_37,N_1278);
nand U3267 (N_3267,N_1254,N_529);
nor U3268 (N_3268,N_2376,N_1375);
nand U3269 (N_3269,N_2151,N_2499);
and U3270 (N_3270,N_365,N_1745);
nor U3271 (N_3271,N_1604,N_1867);
nor U3272 (N_3272,N_1741,N_479);
nand U3273 (N_3273,N_891,N_1820);
nand U3274 (N_3274,N_1818,N_1032);
nand U3275 (N_3275,N_6,N_1379);
and U3276 (N_3276,N_1992,N_1905);
and U3277 (N_3277,N_1746,N_816);
or U3278 (N_3278,N_2479,N_1544);
or U3279 (N_3279,N_1227,N_2167);
or U3280 (N_3280,N_1655,N_906);
nor U3281 (N_3281,N_637,N_1624);
or U3282 (N_3282,N_2457,N_1373);
nand U3283 (N_3283,N_595,N_675);
or U3284 (N_3284,N_1150,N_1548);
nor U3285 (N_3285,N_378,N_875);
nand U3286 (N_3286,N_1501,N_1165);
or U3287 (N_3287,N_1192,N_2256);
and U3288 (N_3288,N_157,N_293);
and U3289 (N_3289,N_1271,N_1193);
nor U3290 (N_3290,N_2031,N_503);
and U3291 (N_3291,N_1418,N_1826);
nand U3292 (N_3292,N_111,N_925);
nor U3293 (N_3293,N_1839,N_1008);
nand U3294 (N_3294,N_1443,N_2047);
or U3295 (N_3295,N_1999,N_393);
and U3296 (N_3296,N_43,N_968);
nor U3297 (N_3297,N_520,N_2494);
or U3298 (N_3298,N_1729,N_766);
nand U3299 (N_3299,N_951,N_1012);
or U3300 (N_3300,N_628,N_462);
nand U3301 (N_3301,N_1685,N_2119);
nor U3302 (N_3302,N_1403,N_873);
nand U3303 (N_3303,N_2313,N_1506);
and U3304 (N_3304,N_264,N_498);
or U3305 (N_3305,N_2429,N_2148);
and U3306 (N_3306,N_2410,N_445);
and U3307 (N_3307,N_589,N_1499);
and U3308 (N_3308,N_510,N_1352);
or U3309 (N_3309,N_416,N_342);
or U3310 (N_3310,N_823,N_2224);
nor U3311 (N_3311,N_534,N_256);
or U3312 (N_3312,N_1808,N_1931);
nand U3313 (N_3313,N_1236,N_1866);
or U3314 (N_3314,N_1210,N_250);
nor U3315 (N_3315,N_1760,N_899);
and U3316 (N_3316,N_1517,N_672);
nand U3317 (N_3317,N_1953,N_2245);
or U3318 (N_3318,N_361,N_1383);
and U3319 (N_3319,N_2491,N_1532);
nand U3320 (N_3320,N_953,N_825);
or U3321 (N_3321,N_1968,N_1277);
and U3322 (N_3322,N_708,N_2199);
or U3323 (N_3323,N_1328,N_1131);
and U3324 (N_3324,N_124,N_80);
and U3325 (N_3325,N_1291,N_1886);
nor U3326 (N_3326,N_2011,N_2470);
nand U3327 (N_3327,N_1300,N_734);
nand U3328 (N_3328,N_2448,N_93);
nor U3329 (N_3329,N_1735,N_1864);
or U3330 (N_3330,N_1716,N_243);
nor U3331 (N_3331,N_1908,N_1862);
and U3332 (N_3332,N_1393,N_65);
nor U3333 (N_3333,N_1265,N_1324);
nand U3334 (N_3334,N_1626,N_1397);
or U3335 (N_3335,N_1171,N_2495);
nor U3336 (N_3336,N_2177,N_1579);
nand U3337 (N_3337,N_2213,N_2233);
nor U3338 (N_3338,N_1963,N_370);
xor U3339 (N_3339,N_555,N_2033);
nand U3340 (N_3340,N_981,N_1784);
nor U3341 (N_3341,N_682,N_1081);
or U3342 (N_3342,N_2365,N_1583);
nand U3343 (N_3343,N_1817,N_1577);
nor U3344 (N_3344,N_2050,N_918);
and U3345 (N_3345,N_1248,N_1290);
or U3346 (N_3346,N_772,N_2252);
or U3347 (N_3347,N_2437,N_39);
or U3348 (N_3348,N_2296,N_837);
and U3349 (N_3349,N_265,N_1338);
or U3350 (N_3350,N_218,N_803);
and U3351 (N_3351,N_134,N_720);
and U3352 (N_3352,N_1779,N_16);
nor U3353 (N_3353,N_1394,N_745);
or U3354 (N_3354,N_1003,N_947);
or U3355 (N_3355,N_64,N_195);
nor U3356 (N_3356,N_429,N_612);
and U3357 (N_3357,N_276,N_1965);
or U3358 (N_3358,N_910,N_207);
nor U3359 (N_3359,N_1713,N_484);
nor U3360 (N_3360,N_691,N_1598);
nor U3361 (N_3361,N_2131,N_2216);
or U3362 (N_3362,N_331,N_1911);
or U3363 (N_3363,N_1446,N_2471);
nor U3364 (N_3364,N_397,N_192);
nor U3365 (N_3365,N_149,N_1958);
and U3366 (N_3366,N_1976,N_945);
and U3367 (N_3367,N_1704,N_933);
nand U3368 (N_3368,N_892,N_1599);
nand U3369 (N_3369,N_2106,N_292);
nand U3370 (N_3370,N_1293,N_502);
and U3371 (N_3371,N_884,N_2220);
nand U3372 (N_3372,N_1865,N_1812);
and U3373 (N_3373,N_333,N_221);
xnor U3374 (N_3374,N_2197,N_1257);
or U3375 (N_3375,N_1445,N_2468);
nor U3376 (N_3376,N_1543,N_156);
nand U3377 (N_3377,N_601,N_1179);
nand U3378 (N_3378,N_740,N_1551);
or U3379 (N_3379,N_456,N_767);
or U3380 (N_3380,N_1387,N_1996);
and U3381 (N_3381,N_1847,N_686);
or U3382 (N_3382,N_846,N_983);
nand U3383 (N_3383,N_714,N_336);
nor U3384 (N_3384,N_2289,N_2173);
nand U3385 (N_3385,N_12,N_1912);
or U3386 (N_3386,N_594,N_655);
nand U3387 (N_3387,N_1884,N_2201);
nand U3388 (N_3388,N_1611,N_1927);
and U3389 (N_3389,N_1900,N_1281);
and U3390 (N_3390,N_447,N_785);
nor U3391 (N_3391,N_1304,N_2063);
nor U3392 (N_3392,N_2085,N_1169);
nand U3393 (N_3393,N_621,N_2078);
nor U3394 (N_3394,N_404,N_2309);
nand U3395 (N_3395,N_1483,N_1667);
and U3396 (N_3396,N_1803,N_2114);
and U3397 (N_3397,N_1891,N_787);
nor U3398 (N_3398,N_2251,N_2392);
and U3399 (N_3399,N_1781,N_407);
or U3400 (N_3400,N_1753,N_591);
or U3401 (N_3401,N_886,N_2038);
or U3402 (N_3402,N_90,N_410);
and U3403 (N_3403,N_338,N_1841);
or U3404 (N_3404,N_1190,N_123);
and U3405 (N_3405,N_32,N_2450);
nand U3406 (N_3406,N_2154,N_1821);
nand U3407 (N_3407,N_1969,N_1095);
nand U3408 (N_3408,N_789,N_1732);
or U3409 (N_3409,N_1898,N_2013);
nand U3410 (N_3410,N_2472,N_660);
and U3411 (N_3411,N_1828,N_671);
or U3412 (N_3412,N_366,N_319);
nor U3413 (N_3413,N_1717,N_1334);
and U3414 (N_3414,N_893,N_1766);
and U3415 (N_3415,N_2445,N_1666);
or U3416 (N_3416,N_432,N_1176);
and U3417 (N_3417,N_1620,N_1923);
or U3418 (N_3418,N_1945,N_2246);
and U3419 (N_3419,N_1520,N_796);
and U3420 (N_3420,N_2369,N_778);
xnor U3421 (N_3421,N_2035,N_634);
and U3422 (N_3422,N_1476,N_709);
nor U3423 (N_3423,N_2302,N_2155);
or U3424 (N_3424,N_1152,N_2320);
or U3425 (N_3425,N_2421,N_1653);
or U3426 (N_3426,N_2134,N_697);
or U3427 (N_3427,N_200,N_21);
nand U3428 (N_3428,N_4,N_852);
nand U3429 (N_3429,N_624,N_2261);
or U3430 (N_3430,N_704,N_1691);
or U3431 (N_3431,N_1872,N_1323);
nand U3432 (N_3432,N_1133,N_2427);
nand U3433 (N_3433,N_896,N_2191);
nor U3434 (N_3434,N_773,N_1058);
xnor U3435 (N_3435,N_1890,N_631);
and U3436 (N_3436,N_1823,N_1879);
or U3437 (N_3437,N_1366,N_1649);
or U3438 (N_3438,N_2202,N_1951);
nor U3439 (N_3439,N_2350,N_1239);
nand U3440 (N_3440,N_1643,N_2444);
and U3441 (N_3441,N_1764,N_1023);
nor U3442 (N_3442,N_1877,N_1454);
and U3443 (N_3443,N_443,N_505);
nand U3444 (N_3444,N_2328,N_689);
and U3445 (N_3445,N_525,N_1742);
nor U3446 (N_3446,N_109,N_2449);
nand U3447 (N_3447,N_811,N_1502);
and U3448 (N_3448,N_1545,N_339);
nand U3449 (N_3449,N_1092,N_1542);
nor U3450 (N_3450,N_343,N_210);
and U3451 (N_3451,N_154,N_1944);
nand U3452 (N_3452,N_2161,N_746);
or U3453 (N_3453,N_328,N_1528);
and U3454 (N_3454,N_1346,N_1342);
nor U3455 (N_3455,N_1009,N_95);
xnor U3456 (N_3456,N_63,N_1515);
or U3457 (N_3457,N_2237,N_1376);
nand U3458 (N_3458,N_1471,N_1561);
nand U3459 (N_3459,N_2254,N_78);
nand U3460 (N_3460,N_866,N_1235);
nor U3461 (N_3461,N_53,N_2087);
or U3462 (N_3462,N_587,N_1675);
nand U3463 (N_3463,N_341,N_288);
or U3464 (N_3464,N_940,N_386);
nand U3465 (N_3465,N_2270,N_2284);
nand U3466 (N_3466,N_321,N_576);
nand U3467 (N_3467,N_922,N_1306);
nor U3468 (N_3468,N_877,N_1783);
or U3469 (N_3469,N_1147,N_1113);
or U3470 (N_3470,N_1993,N_231);
nand U3471 (N_3471,N_1493,N_2374);
nor U3472 (N_3472,N_451,N_764);
nand U3473 (N_3473,N_347,N_1123);
nor U3474 (N_3474,N_2041,N_2018);
or U3475 (N_3475,N_1696,N_943);
nor U3476 (N_3476,N_236,N_543);
and U3477 (N_3477,N_987,N_73);
nand U3478 (N_3478,N_1088,N_1332);
nor U3479 (N_3479,N_2317,N_353);
nand U3480 (N_3480,N_183,N_1775);
nand U3481 (N_3481,N_658,N_2475);
nor U3482 (N_3482,N_1961,N_2378);
and U3483 (N_3483,N_1191,N_1117);
and U3484 (N_3484,N_1906,N_1238);
nor U3485 (N_3485,N_1720,N_1562);
and U3486 (N_3486,N_468,N_2088);
or U3487 (N_3487,N_552,N_775);
and U3488 (N_3488,N_568,N_623);
and U3489 (N_3489,N_1690,N_1462);
or U3490 (N_3490,N_1262,N_2417);
nand U3491 (N_3491,N_270,N_2156);
and U3492 (N_3492,N_805,N_2303);
and U3493 (N_3493,N_2227,N_1952);
nand U3494 (N_3494,N_1256,N_878);
nand U3495 (N_3495,N_1825,N_1211);
or U3496 (N_3496,N_1444,N_1788);
and U3497 (N_3497,N_914,N_75);
or U3498 (N_3498,N_1863,N_2291);
nand U3499 (N_3499,N_575,N_101);
nand U3500 (N_3500,N_1607,N_963);
and U3501 (N_3501,N_765,N_758);
or U3502 (N_3502,N_136,N_1793);
and U3503 (N_3503,N_2172,N_2093);
nor U3504 (N_3504,N_1769,N_1926);
or U3505 (N_3505,N_2402,N_1408);
nor U3506 (N_3506,N_273,N_1706);
nor U3507 (N_3507,N_2405,N_600);
and U3508 (N_3508,N_1016,N_1933);
or U3509 (N_3509,N_1181,N_2322);
nand U3510 (N_3510,N_2082,N_1464);
nand U3511 (N_3511,N_1096,N_965);
nand U3512 (N_3512,N_690,N_1255);
and U3513 (N_3513,N_327,N_1409);
and U3514 (N_3514,N_2348,N_1246);
and U3515 (N_3515,N_330,N_1458);
or U3516 (N_3516,N_610,N_858);
nand U3517 (N_3517,N_2359,N_208);
nor U3518 (N_3518,N_563,N_2431);
nand U3519 (N_3519,N_618,N_320);
and U3520 (N_3520,N_1534,N_2316);
or U3521 (N_3521,N_700,N_2425);
or U3522 (N_3522,N_513,N_560);
nor U3523 (N_3523,N_2344,N_1962);
nor U3524 (N_3524,N_129,N_1434);
or U3525 (N_3525,N_794,N_1669);
or U3526 (N_3526,N_1196,N_2232);
or U3527 (N_3527,N_1855,N_1063);
and U3528 (N_3528,N_166,N_1372);
or U3529 (N_3529,N_1452,N_1979);
and U3530 (N_3530,N_2415,N_2478);
nand U3531 (N_3531,N_779,N_2212);
xnor U3532 (N_3532,N_1077,N_997);
and U3533 (N_3533,N_2398,N_1121);
nor U3534 (N_3534,N_1472,N_874);
and U3535 (N_3535,N_1412,N_1565);
and U3536 (N_3536,N_182,N_725);
xor U3537 (N_3537,N_1137,N_1682);
and U3538 (N_3538,N_1351,N_919);
nand U3539 (N_3539,N_1461,N_550);
and U3540 (N_3540,N_54,N_882);
nor U3541 (N_3541,N_1075,N_1875);
or U3542 (N_3542,N_1744,N_1571);
nor U3543 (N_3543,N_2312,N_406);
and U3544 (N_3544,N_647,N_2075);
and U3545 (N_3545,N_715,N_2079);
nand U3546 (N_3546,N_86,N_1731);
and U3547 (N_3547,N_2366,N_1772);
nor U3548 (N_3548,N_522,N_1374);
or U3549 (N_3549,N_94,N_1455);
or U3550 (N_3550,N_2222,N_7);
or U3551 (N_3551,N_2007,N_315);
or U3552 (N_3552,N_283,N_399);
or U3553 (N_3553,N_1014,N_994);
or U3554 (N_3554,N_1473,N_571);
or U3555 (N_3555,N_524,N_294);
and U3556 (N_3556,N_55,N_401);
nor U3557 (N_3557,N_1314,N_1401);
nor U3558 (N_3558,N_2021,N_390);
nor U3559 (N_3559,N_1364,N_2176);
nand U3560 (N_3560,N_1602,N_1076);
nor U3561 (N_3561,N_2413,N_1638);
and U3562 (N_3562,N_1910,N_699);
nor U3563 (N_3563,N_2281,N_954);
and U3564 (N_3564,N_2169,N_1697);
nand U3565 (N_3565,N_1917,N_2117);
and U3566 (N_3566,N_2101,N_2420);
nor U3567 (N_3567,N_1954,N_570);
and U3568 (N_3568,N_2380,N_2211);
or U3569 (N_3569,N_2272,N_1017);
nor U3570 (N_3570,N_948,N_2412);
nand U3571 (N_3571,N_2230,N_1722);
nand U3572 (N_3572,N_1430,N_2441);
nor U3573 (N_3573,N_1358,N_1219);
nand U3574 (N_3574,N_1576,N_736);
and U3575 (N_3575,N_84,N_762);
or U3576 (N_3576,N_848,N_1609);
and U3577 (N_3577,N_1594,N_1156);
and U3578 (N_3578,N_408,N_851);
nand U3579 (N_3579,N_2300,N_240);
nor U3580 (N_3580,N_194,N_1159);
nor U3581 (N_3581,N_1829,N_1208);
or U3582 (N_3582,N_1045,N_307);
nor U3583 (N_3583,N_2099,N_1474);
or U3584 (N_3584,N_1668,N_1881);
nor U3585 (N_3585,N_2044,N_2324);
or U3586 (N_3586,N_1538,N_2381);
nand U3587 (N_3587,N_695,N_2140);
nand U3588 (N_3588,N_1421,N_2337);
or U3589 (N_3589,N_1234,N_2137);
nor U3590 (N_3590,N_630,N_1790);
nand U3591 (N_3591,N_698,N_1361);
nand U3592 (N_3592,N_1006,N_2333);
and U3593 (N_3593,N_364,N_1658);
and U3594 (N_3594,N_557,N_1209);
and U3595 (N_3595,N_701,N_28);
nand U3596 (N_3596,N_653,N_547);
nor U3597 (N_3597,N_2242,N_888);
nor U3598 (N_3598,N_2125,N_417);
nand U3599 (N_3599,N_1712,N_423);
and U3600 (N_3600,N_986,N_0);
and U3601 (N_3601,N_569,N_1185);
nor U3602 (N_3602,N_2295,N_792);
or U3603 (N_3603,N_665,N_1909);
nand U3604 (N_3604,N_2467,N_2266);
or U3605 (N_3605,N_278,N_1767);
nor U3606 (N_3606,N_564,N_992);
and U3607 (N_3607,N_139,N_1056);
nor U3608 (N_3608,N_1251,N_735);
nand U3609 (N_3609,N_1942,N_295);
nor U3610 (N_3610,N_2297,N_1080);
and U3611 (N_3611,N_538,N_1679);
and U3612 (N_3612,N_1098,N_467);
or U3613 (N_3613,N_2287,N_1748);
and U3614 (N_3614,N_47,N_251);
nand U3615 (N_3615,N_8,N_586);
and U3616 (N_3616,N_62,N_1220);
or U3617 (N_3617,N_1420,N_620);
nand U3618 (N_3618,N_535,N_1899);
or U3619 (N_3619,N_391,N_1749);
and U3620 (N_3620,N_1880,N_1205);
nand U3621 (N_3621,N_2473,N_2163);
and U3622 (N_3622,N_437,N_1549);
and U3623 (N_3623,N_496,N_2386);
nand U3624 (N_3624,N_1106,N_2149);
or U3625 (N_3625,N_1298,N_1447);
and U3626 (N_3626,N_1413,N_27);
and U3627 (N_3627,N_1456,N_2265);
nand U3628 (N_3628,N_712,N_2292);
nor U3629 (N_3629,N_2056,N_966);
nor U3630 (N_3630,N_2247,N_1681);
nand U3631 (N_3631,N_749,N_116);
nand U3632 (N_3632,N_1837,N_1348);
nor U3633 (N_3633,N_703,N_1518);
or U3634 (N_3634,N_76,N_561);
nand U3635 (N_3635,N_2477,N_1603);
or U3636 (N_3636,N_2138,N_2054);
or U3637 (N_3637,N_226,N_2416);
nand U3638 (N_3638,N_553,N_2269);
or U3639 (N_3639,N_578,N_1392);
or U3640 (N_3640,N_225,N_1827);
nor U3641 (N_3641,N_597,N_34);
nand U3642 (N_3642,N_2277,N_2484);
or U3643 (N_3643,N_1086,N_2268);
nand U3644 (N_3644,N_2408,N_1771);
or U3645 (N_3645,N_1280,N_738);
nand U3646 (N_3646,N_2068,N_1688);
and U3647 (N_3647,N_857,N_2424);
or U3648 (N_3648,N_508,N_2388);
and U3649 (N_3649,N_1184,N_96);
or U3650 (N_3650,N_426,N_2396);
nor U3651 (N_3651,N_380,N_1386);
xnor U3652 (N_3652,N_2409,N_1539);
and U3653 (N_3653,N_1737,N_2040);
and U3654 (N_3654,N_33,N_1166);
or U3655 (N_3655,N_199,N_1269);
or U3656 (N_3656,N_446,N_303);
nand U3657 (N_3657,N_420,N_1223);
or U3658 (N_3658,N_718,N_1074);
nand U3659 (N_3659,N_1170,N_1971);
nor U3660 (N_3660,N_2105,N_1283);
nand U3661 (N_3661,N_935,N_842);
and U3662 (N_3662,N_1774,N_58);
and U3663 (N_3663,N_220,N_2171);
nand U3664 (N_3664,N_1296,N_777);
and U3665 (N_3665,N_1902,N_2332);
nor U3666 (N_3666,N_435,N_1229);
or U3667 (N_3667,N_246,N_645);
or U3668 (N_3668,N_1657,N_638);
or U3669 (N_3669,N_1719,N_1425);
nor U3670 (N_3670,N_1085,N_2037);
and U3671 (N_3671,N_2111,N_2184);
nand U3672 (N_3672,N_1797,N_1167);
nand U3673 (N_3673,N_267,N_135);
nand U3674 (N_3674,N_2414,N_876);
nand U3675 (N_3675,N_190,N_1453);
and U3676 (N_3676,N_118,N_549);
nor U3677 (N_3677,N_269,N_938);
nand U3678 (N_3678,N_2373,N_1027);
nand U3679 (N_3679,N_259,N_1380);
and U3680 (N_3680,N_1038,N_1498);
nor U3681 (N_3681,N_1242,N_817);
and U3682 (N_3682,N_2109,N_770);
or U3683 (N_3683,N_1514,N_1030);
nor U3684 (N_3684,N_2488,N_1736);
or U3685 (N_3685,N_400,N_24);
or U3686 (N_3686,N_809,N_737);
or U3687 (N_3687,N_244,N_1530);
and U3688 (N_3688,N_1104,N_418);
xnor U3689 (N_3689,N_2404,N_949);
and U3690 (N_3690,N_1207,N_1059);
nor U3691 (N_3691,N_826,N_915);
nor U3692 (N_3692,N_323,N_1347);
nand U3693 (N_3693,N_201,N_786);
nand U3694 (N_3694,N_609,N_290);
nor U3695 (N_3695,N_113,N_1252);
and U3696 (N_3696,N_654,N_457);
or U3697 (N_3697,N_651,N_582);
or U3698 (N_3698,N_1128,N_2120);
xor U3699 (N_3699,N_629,N_1698);
nand U3700 (N_3700,N_1623,N_1362);
nand U3701 (N_3701,N_146,N_1759);
or U3702 (N_3702,N_345,N_1333);
and U3703 (N_3703,N_2116,N_31);
or U3704 (N_3704,N_1673,N_1816);
nor U3705 (N_3705,N_1097,N_2464);
nand U3706 (N_3706,N_768,N_1490);
nor U3707 (N_3707,N_585,N_1956);
nand U3708 (N_3708,N_1896,N_1503);
nor U3709 (N_3709,N_19,N_1040);
nor U3710 (N_3710,N_1792,N_441);
and U3711 (N_3711,N_152,N_2027);
and U3712 (N_3712,N_1213,N_289);
and U3713 (N_3713,N_1240,N_1276);
and U3714 (N_3714,N_48,N_2135);
and U3715 (N_3715,N_2183,N_5);
nand U3716 (N_3716,N_175,N_213);
and U3717 (N_3717,N_974,N_1356);
nor U3718 (N_3718,N_1365,N_1258);
nor U3719 (N_3719,N_1677,N_1158);
nor U3720 (N_3720,N_1552,N_683);
or U3721 (N_3721,N_1055,N_2334);
and U3722 (N_3722,N_1084,N_1580);
and U3723 (N_3723,N_2390,N_1904);
and U3724 (N_3724,N_478,N_1914);
and U3725 (N_3725,N_2015,N_1288);
and U3726 (N_3726,N_487,N_1568);
and U3727 (N_3727,N_2476,N_1778);
nor U3728 (N_3728,N_1360,N_2433);
nand U3729 (N_3729,N_2006,N_2028);
nand U3730 (N_3730,N_499,N_491);
nand U3731 (N_3731,N_1924,N_1489);
and U3732 (N_3732,N_431,N_2009);
or U3733 (N_3733,N_1662,N_1813);
nand U3734 (N_3734,N_26,N_13);
nand U3735 (N_3735,N_833,N_1614);
and U3736 (N_3736,N_1730,N_1725);
nor U3737 (N_3737,N_2401,N_911);
and U3738 (N_3738,N_2143,N_2198);
nand U3739 (N_3739,N_985,N_1644);
or U3740 (N_3740,N_1757,N_1635);
or U3741 (N_3741,N_1146,N_1451);
and U3742 (N_3742,N_1946,N_1980);
and U3743 (N_3743,N_150,N_2288);
and U3744 (N_3744,N_1947,N_2160);
or U3745 (N_3745,N_1572,N_993);
nand U3746 (N_3746,N_359,N_931);
nand U3747 (N_3747,N_2214,N_751);
or U3748 (N_3748,N_2423,N_1470);
and U3749 (N_3749,N_389,N_537);
or U3750 (N_3750,N_2414,N_1725);
and U3751 (N_3751,N_798,N_2374);
and U3752 (N_3752,N_26,N_1305);
nand U3753 (N_3753,N_1366,N_824);
nand U3754 (N_3754,N_105,N_200);
and U3755 (N_3755,N_90,N_965);
or U3756 (N_3756,N_631,N_2034);
and U3757 (N_3757,N_1719,N_192);
and U3758 (N_3758,N_2348,N_912);
nand U3759 (N_3759,N_248,N_364);
and U3760 (N_3760,N_2291,N_48);
nand U3761 (N_3761,N_548,N_928);
nor U3762 (N_3762,N_2465,N_1606);
or U3763 (N_3763,N_1360,N_1015);
nand U3764 (N_3764,N_1274,N_2460);
nor U3765 (N_3765,N_2067,N_1850);
nor U3766 (N_3766,N_1335,N_453);
nor U3767 (N_3767,N_6,N_444);
and U3768 (N_3768,N_79,N_2316);
and U3769 (N_3769,N_1882,N_187);
nor U3770 (N_3770,N_1445,N_2064);
or U3771 (N_3771,N_2356,N_1633);
nand U3772 (N_3772,N_1585,N_297);
and U3773 (N_3773,N_761,N_1008);
and U3774 (N_3774,N_1524,N_236);
nor U3775 (N_3775,N_42,N_361);
and U3776 (N_3776,N_1515,N_2387);
nor U3777 (N_3777,N_1196,N_1202);
or U3778 (N_3778,N_1616,N_300);
nand U3779 (N_3779,N_2071,N_317);
and U3780 (N_3780,N_1401,N_1932);
or U3781 (N_3781,N_491,N_1515);
nor U3782 (N_3782,N_634,N_1805);
and U3783 (N_3783,N_983,N_1132);
nor U3784 (N_3784,N_22,N_1553);
or U3785 (N_3785,N_1183,N_950);
nor U3786 (N_3786,N_1739,N_49);
or U3787 (N_3787,N_742,N_2276);
nand U3788 (N_3788,N_1435,N_505);
xnor U3789 (N_3789,N_1851,N_824);
nand U3790 (N_3790,N_1717,N_559);
nor U3791 (N_3791,N_206,N_1715);
and U3792 (N_3792,N_189,N_1450);
or U3793 (N_3793,N_1785,N_398);
and U3794 (N_3794,N_1542,N_1216);
nor U3795 (N_3795,N_1257,N_2155);
and U3796 (N_3796,N_302,N_1304);
and U3797 (N_3797,N_2448,N_2120);
or U3798 (N_3798,N_2255,N_1546);
and U3799 (N_3799,N_792,N_879);
nor U3800 (N_3800,N_3,N_576);
nor U3801 (N_3801,N_260,N_1209);
and U3802 (N_3802,N_490,N_442);
and U3803 (N_3803,N_1845,N_170);
nor U3804 (N_3804,N_147,N_1853);
nor U3805 (N_3805,N_575,N_757);
or U3806 (N_3806,N_1988,N_1061);
nand U3807 (N_3807,N_2200,N_2323);
nand U3808 (N_3808,N_1014,N_1055);
nand U3809 (N_3809,N_1779,N_786);
nand U3810 (N_3810,N_21,N_421);
or U3811 (N_3811,N_1925,N_1316);
and U3812 (N_3812,N_359,N_508);
nor U3813 (N_3813,N_101,N_1675);
or U3814 (N_3814,N_892,N_2306);
nand U3815 (N_3815,N_439,N_445);
and U3816 (N_3816,N_1555,N_1979);
nand U3817 (N_3817,N_1203,N_758);
and U3818 (N_3818,N_1730,N_258);
and U3819 (N_3819,N_2462,N_2299);
or U3820 (N_3820,N_264,N_783);
or U3821 (N_3821,N_848,N_1917);
nor U3822 (N_3822,N_1245,N_627);
nand U3823 (N_3823,N_1535,N_1065);
nand U3824 (N_3824,N_1857,N_426);
and U3825 (N_3825,N_2024,N_1750);
and U3826 (N_3826,N_2365,N_257);
or U3827 (N_3827,N_1564,N_185);
nor U3828 (N_3828,N_1559,N_2122);
and U3829 (N_3829,N_1819,N_299);
or U3830 (N_3830,N_1905,N_451);
or U3831 (N_3831,N_1433,N_371);
nor U3832 (N_3832,N_2180,N_1356);
nor U3833 (N_3833,N_865,N_1157);
nor U3834 (N_3834,N_1830,N_2410);
or U3835 (N_3835,N_892,N_877);
and U3836 (N_3836,N_176,N_2002);
nor U3837 (N_3837,N_355,N_2258);
and U3838 (N_3838,N_1377,N_2140);
nand U3839 (N_3839,N_1983,N_299);
nand U3840 (N_3840,N_2300,N_2216);
nand U3841 (N_3841,N_1175,N_311);
nand U3842 (N_3842,N_665,N_1251);
and U3843 (N_3843,N_2135,N_1997);
nor U3844 (N_3844,N_2155,N_1206);
nor U3845 (N_3845,N_84,N_473);
nand U3846 (N_3846,N_1560,N_1376);
nor U3847 (N_3847,N_1992,N_705);
or U3848 (N_3848,N_1555,N_1191);
nand U3849 (N_3849,N_527,N_687);
nand U3850 (N_3850,N_2256,N_656);
or U3851 (N_3851,N_1849,N_1551);
nor U3852 (N_3852,N_415,N_641);
and U3853 (N_3853,N_13,N_1721);
or U3854 (N_3854,N_209,N_666);
nor U3855 (N_3855,N_1886,N_1132);
nor U3856 (N_3856,N_399,N_1335);
nor U3857 (N_3857,N_404,N_58);
nand U3858 (N_3858,N_327,N_2093);
nand U3859 (N_3859,N_1090,N_377);
or U3860 (N_3860,N_799,N_1719);
or U3861 (N_3861,N_2486,N_409);
nand U3862 (N_3862,N_1440,N_2412);
or U3863 (N_3863,N_650,N_683);
nor U3864 (N_3864,N_1441,N_1139);
nand U3865 (N_3865,N_2038,N_1008);
nor U3866 (N_3866,N_1005,N_518);
or U3867 (N_3867,N_1193,N_200);
nor U3868 (N_3868,N_1235,N_277);
nor U3869 (N_3869,N_2385,N_605);
nand U3870 (N_3870,N_1624,N_180);
nand U3871 (N_3871,N_955,N_1180);
nand U3872 (N_3872,N_1190,N_300);
or U3873 (N_3873,N_2010,N_74);
nand U3874 (N_3874,N_107,N_126);
nor U3875 (N_3875,N_621,N_1133);
nor U3876 (N_3876,N_916,N_1121);
or U3877 (N_3877,N_1728,N_1209);
nand U3878 (N_3878,N_840,N_2486);
and U3879 (N_3879,N_607,N_2027);
nand U3880 (N_3880,N_635,N_2358);
nand U3881 (N_3881,N_662,N_1774);
or U3882 (N_3882,N_1001,N_133);
nor U3883 (N_3883,N_117,N_713);
nor U3884 (N_3884,N_563,N_1754);
and U3885 (N_3885,N_2339,N_213);
nand U3886 (N_3886,N_110,N_1546);
and U3887 (N_3887,N_2054,N_887);
nor U3888 (N_3888,N_900,N_1445);
or U3889 (N_3889,N_1277,N_2355);
nand U3890 (N_3890,N_507,N_2357);
or U3891 (N_3891,N_78,N_2238);
or U3892 (N_3892,N_1560,N_1182);
nor U3893 (N_3893,N_1692,N_1095);
nor U3894 (N_3894,N_988,N_1956);
nand U3895 (N_3895,N_1317,N_1063);
and U3896 (N_3896,N_1798,N_881);
nand U3897 (N_3897,N_634,N_1014);
nor U3898 (N_3898,N_1488,N_2269);
and U3899 (N_3899,N_460,N_717);
or U3900 (N_3900,N_2457,N_101);
or U3901 (N_3901,N_1374,N_609);
nand U3902 (N_3902,N_255,N_2083);
and U3903 (N_3903,N_440,N_363);
nor U3904 (N_3904,N_422,N_83);
and U3905 (N_3905,N_915,N_1855);
nor U3906 (N_3906,N_1526,N_90);
and U3907 (N_3907,N_1640,N_1169);
and U3908 (N_3908,N_1926,N_201);
and U3909 (N_3909,N_248,N_1401);
nand U3910 (N_3910,N_1891,N_2391);
and U3911 (N_3911,N_266,N_109);
and U3912 (N_3912,N_743,N_767);
nand U3913 (N_3913,N_1554,N_2301);
nor U3914 (N_3914,N_686,N_2205);
nand U3915 (N_3915,N_506,N_736);
or U3916 (N_3916,N_2219,N_1299);
nor U3917 (N_3917,N_1414,N_1295);
or U3918 (N_3918,N_1104,N_726);
or U3919 (N_3919,N_204,N_1443);
nor U3920 (N_3920,N_466,N_1587);
and U3921 (N_3921,N_355,N_685);
nand U3922 (N_3922,N_557,N_2029);
nand U3923 (N_3923,N_693,N_1908);
or U3924 (N_3924,N_207,N_896);
nand U3925 (N_3925,N_1114,N_1012);
nor U3926 (N_3926,N_716,N_2395);
nor U3927 (N_3927,N_2181,N_758);
and U3928 (N_3928,N_2140,N_908);
nor U3929 (N_3929,N_495,N_915);
nor U3930 (N_3930,N_2112,N_1425);
or U3931 (N_3931,N_1703,N_351);
or U3932 (N_3932,N_755,N_2052);
or U3933 (N_3933,N_1787,N_61);
and U3934 (N_3934,N_908,N_80);
nand U3935 (N_3935,N_531,N_2090);
and U3936 (N_3936,N_978,N_1277);
nand U3937 (N_3937,N_860,N_1784);
nor U3938 (N_3938,N_1766,N_347);
nor U3939 (N_3939,N_905,N_636);
nand U3940 (N_3940,N_94,N_1503);
nand U3941 (N_3941,N_875,N_1998);
nand U3942 (N_3942,N_1523,N_1936);
nor U3943 (N_3943,N_1428,N_11);
and U3944 (N_3944,N_1706,N_1648);
and U3945 (N_3945,N_1431,N_1669);
nand U3946 (N_3946,N_911,N_1390);
nor U3947 (N_3947,N_0,N_1363);
or U3948 (N_3948,N_1665,N_2350);
or U3949 (N_3949,N_1423,N_1654);
nand U3950 (N_3950,N_1514,N_305);
or U3951 (N_3951,N_2188,N_110);
or U3952 (N_3952,N_199,N_1078);
nor U3953 (N_3953,N_1355,N_592);
nand U3954 (N_3954,N_2200,N_1786);
nand U3955 (N_3955,N_951,N_198);
nand U3956 (N_3956,N_1355,N_537);
and U3957 (N_3957,N_1484,N_1449);
and U3958 (N_3958,N_2182,N_16);
nor U3959 (N_3959,N_2027,N_834);
and U3960 (N_3960,N_1129,N_2240);
and U3961 (N_3961,N_1243,N_1817);
and U3962 (N_3962,N_1617,N_1018);
nor U3963 (N_3963,N_201,N_1715);
and U3964 (N_3964,N_580,N_1439);
nand U3965 (N_3965,N_1574,N_310);
xor U3966 (N_3966,N_1943,N_147);
nand U3967 (N_3967,N_227,N_557);
nor U3968 (N_3968,N_219,N_2284);
nand U3969 (N_3969,N_381,N_671);
nor U3970 (N_3970,N_1963,N_2388);
xor U3971 (N_3971,N_2289,N_775);
nand U3972 (N_3972,N_1279,N_1204);
xnor U3973 (N_3973,N_361,N_1613);
or U3974 (N_3974,N_1015,N_1650);
or U3975 (N_3975,N_603,N_2410);
or U3976 (N_3976,N_1559,N_625);
or U3977 (N_3977,N_1803,N_1703);
nand U3978 (N_3978,N_42,N_1582);
and U3979 (N_3979,N_649,N_1914);
nor U3980 (N_3980,N_1597,N_1226);
or U3981 (N_3981,N_756,N_1267);
nor U3982 (N_3982,N_216,N_2209);
and U3983 (N_3983,N_1534,N_1778);
and U3984 (N_3984,N_441,N_1030);
nor U3985 (N_3985,N_2427,N_597);
nand U3986 (N_3986,N_1050,N_228);
xor U3987 (N_3987,N_715,N_1352);
xor U3988 (N_3988,N_1564,N_2408);
nand U3989 (N_3989,N_1468,N_361);
nor U3990 (N_3990,N_1121,N_1066);
nand U3991 (N_3991,N_2127,N_1662);
nand U3992 (N_3992,N_1213,N_2405);
nor U3993 (N_3993,N_38,N_2077);
and U3994 (N_3994,N_1584,N_1956);
or U3995 (N_3995,N_2172,N_90);
and U3996 (N_3996,N_2300,N_837);
and U3997 (N_3997,N_1663,N_2211);
and U3998 (N_3998,N_1265,N_1912);
and U3999 (N_3999,N_34,N_1937);
nor U4000 (N_4000,N_850,N_923);
nand U4001 (N_4001,N_2271,N_578);
or U4002 (N_4002,N_825,N_2215);
and U4003 (N_4003,N_2310,N_2007);
nand U4004 (N_4004,N_1857,N_1428);
or U4005 (N_4005,N_2363,N_1879);
nor U4006 (N_4006,N_2461,N_73);
or U4007 (N_4007,N_93,N_2107);
nand U4008 (N_4008,N_431,N_209);
and U4009 (N_4009,N_45,N_2181);
or U4010 (N_4010,N_669,N_1861);
or U4011 (N_4011,N_109,N_2352);
nand U4012 (N_4012,N_1228,N_1087);
or U4013 (N_4013,N_130,N_1282);
and U4014 (N_4014,N_72,N_815);
and U4015 (N_4015,N_1131,N_218);
nor U4016 (N_4016,N_397,N_2207);
nand U4017 (N_4017,N_79,N_1323);
or U4018 (N_4018,N_356,N_1456);
and U4019 (N_4019,N_1539,N_396);
nand U4020 (N_4020,N_1081,N_2071);
nand U4021 (N_4021,N_1131,N_1748);
nor U4022 (N_4022,N_345,N_53);
nand U4023 (N_4023,N_1630,N_1786);
and U4024 (N_4024,N_2177,N_1031);
and U4025 (N_4025,N_79,N_350);
or U4026 (N_4026,N_1803,N_1708);
nand U4027 (N_4027,N_1997,N_1009);
or U4028 (N_4028,N_2326,N_396);
nand U4029 (N_4029,N_1989,N_514);
nand U4030 (N_4030,N_540,N_1427);
and U4031 (N_4031,N_1173,N_1468);
or U4032 (N_4032,N_1576,N_580);
and U4033 (N_4033,N_1080,N_1350);
and U4034 (N_4034,N_750,N_30);
nand U4035 (N_4035,N_2437,N_1114);
nand U4036 (N_4036,N_397,N_1611);
or U4037 (N_4037,N_2408,N_2295);
nand U4038 (N_4038,N_2480,N_589);
nor U4039 (N_4039,N_608,N_1526);
nand U4040 (N_4040,N_794,N_1766);
and U4041 (N_4041,N_606,N_2055);
xnor U4042 (N_4042,N_951,N_1534);
nor U4043 (N_4043,N_2411,N_1482);
nor U4044 (N_4044,N_2294,N_1949);
or U4045 (N_4045,N_1178,N_1508);
nor U4046 (N_4046,N_273,N_721);
and U4047 (N_4047,N_2241,N_2006);
and U4048 (N_4048,N_1065,N_1194);
and U4049 (N_4049,N_1863,N_961);
and U4050 (N_4050,N_256,N_187);
nand U4051 (N_4051,N_358,N_704);
nand U4052 (N_4052,N_1570,N_1455);
and U4053 (N_4053,N_2025,N_379);
nand U4054 (N_4054,N_1214,N_2319);
and U4055 (N_4055,N_358,N_130);
nor U4056 (N_4056,N_408,N_1149);
nor U4057 (N_4057,N_2401,N_1301);
nand U4058 (N_4058,N_742,N_365);
nor U4059 (N_4059,N_1908,N_1170);
and U4060 (N_4060,N_140,N_1704);
or U4061 (N_4061,N_1244,N_2405);
or U4062 (N_4062,N_2196,N_2181);
and U4063 (N_4063,N_748,N_74);
nand U4064 (N_4064,N_1184,N_2382);
and U4065 (N_4065,N_989,N_1697);
or U4066 (N_4066,N_204,N_809);
xor U4067 (N_4067,N_358,N_993);
and U4068 (N_4068,N_2193,N_2496);
or U4069 (N_4069,N_244,N_1436);
nand U4070 (N_4070,N_45,N_1196);
or U4071 (N_4071,N_1087,N_133);
or U4072 (N_4072,N_46,N_885);
nand U4073 (N_4073,N_897,N_2063);
nor U4074 (N_4074,N_99,N_1595);
or U4075 (N_4075,N_2450,N_1208);
nand U4076 (N_4076,N_853,N_654);
nand U4077 (N_4077,N_608,N_97);
or U4078 (N_4078,N_977,N_1631);
or U4079 (N_4079,N_1242,N_731);
or U4080 (N_4080,N_474,N_2108);
and U4081 (N_4081,N_842,N_110);
nand U4082 (N_4082,N_1614,N_1431);
and U4083 (N_4083,N_1355,N_1282);
and U4084 (N_4084,N_1769,N_100);
nor U4085 (N_4085,N_724,N_1186);
and U4086 (N_4086,N_1634,N_1519);
or U4087 (N_4087,N_689,N_1724);
nand U4088 (N_4088,N_1946,N_689);
and U4089 (N_4089,N_2319,N_1538);
nor U4090 (N_4090,N_2165,N_1937);
nor U4091 (N_4091,N_2203,N_1193);
or U4092 (N_4092,N_230,N_0);
or U4093 (N_4093,N_1282,N_2176);
and U4094 (N_4094,N_409,N_1335);
nand U4095 (N_4095,N_900,N_1537);
or U4096 (N_4096,N_2073,N_778);
or U4097 (N_4097,N_1231,N_1730);
nor U4098 (N_4098,N_2240,N_1320);
nand U4099 (N_4099,N_874,N_1938);
and U4100 (N_4100,N_1883,N_452);
and U4101 (N_4101,N_1313,N_1183);
nor U4102 (N_4102,N_2334,N_987);
nand U4103 (N_4103,N_868,N_19);
nand U4104 (N_4104,N_717,N_13);
and U4105 (N_4105,N_1612,N_93);
nand U4106 (N_4106,N_1284,N_1773);
and U4107 (N_4107,N_690,N_1780);
and U4108 (N_4108,N_402,N_1901);
nand U4109 (N_4109,N_1098,N_1076);
or U4110 (N_4110,N_856,N_1977);
nand U4111 (N_4111,N_444,N_841);
nor U4112 (N_4112,N_1114,N_2278);
or U4113 (N_4113,N_1668,N_1671);
and U4114 (N_4114,N_2263,N_1274);
and U4115 (N_4115,N_81,N_1330);
nor U4116 (N_4116,N_83,N_712);
nor U4117 (N_4117,N_823,N_1759);
nand U4118 (N_4118,N_314,N_1041);
and U4119 (N_4119,N_2225,N_2295);
nand U4120 (N_4120,N_877,N_1246);
and U4121 (N_4121,N_140,N_0);
or U4122 (N_4122,N_113,N_1466);
and U4123 (N_4123,N_2135,N_658);
or U4124 (N_4124,N_2132,N_1028);
or U4125 (N_4125,N_457,N_1777);
and U4126 (N_4126,N_575,N_176);
or U4127 (N_4127,N_1273,N_1601);
and U4128 (N_4128,N_60,N_185);
or U4129 (N_4129,N_810,N_39);
or U4130 (N_4130,N_1667,N_1071);
or U4131 (N_4131,N_174,N_1044);
and U4132 (N_4132,N_935,N_1043);
nand U4133 (N_4133,N_1983,N_1156);
or U4134 (N_4134,N_2019,N_1637);
and U4135 (N_4135,N_1378,N_1011);
nand U4136 (N_4136,N_600,N_1444);
and U4137 (N_4137,N_527,N_1335);
nand U4138 (N_4138,N_1363,N_2230);
nor U4139 (N_4139,N_1759,N_664);
nand U4140 (N_4140,N_242,N_532);
and U4141 (N_4141,N_1880,N_1440);
nor U4142 (N_4142,N_1124,N_1833);
nor U4143 (N_4143,N_1169,N_1586);
nand U4144 (N_4144,N_246,N_347);
nor U4145 (N_4145,N_451,N_2129);
nor U4146 (N_4146,N_1991,N_937);
and U4147 (N_4147,N_184,N_1318);
or U4148 (N_4148,N_861,N_574);
nor U4149 (N_4149,N_1773,N_466);
nand U4150 (N_4150,N_1639,N_1225);
or U4151 (N_4151,N_40,N_1307);
and U4152 (N_4152,N_416,N_435);
nand U4153 (N_4153,N_603,N_1676);
and U4154 (N_4154,N_1710,N_2372);
xnor U4155 (N_4155,N_175,N_1581);
nor U4156 (N_4156,N_2041,N_1401);
or U4157 (N_4157,N_1653,N_2329);
nand U4158 (N_4158,N_2485,N_876);
and U4159 (N_4159,N_835,N_434);
nor U4160 (N_4160,N_2465,N_2309);
nand U4161 (N_4161,N_698,N_684);
nor U4162 (N_4162,N_1255,N_596);
nand U4163 (N_4163,N_32,N_711);
nand U4164 (N_4164,N_1693,N_2391);
and U4165 (N_4165,N_2069,N_1954);
nor U4166 (N_4166,N_1001,N_2337);
nand U4167 (N_4167,N_83,N_1027);
or U4168 (N_4168,N_696,N_863);
and U4169 (N_4169,N_2309,N_640);
nor U4170 (N_4170,N_1524,N_437);
nor U4171 (N_4171,N_546,N_1757);
nand U4172 (N_4172,N_1278,N_554);
xor U4173 (N_4173,N_1319,N_1810);
nor U4174 (N_4174,N_2097,N_181);
nand U4175 (N_4175,N_1045,N_454);
or U4176 (N_4176,N_275,N_304);
and U4177 (N_4177,N_1989,N_422);
nand U4178 (N_4178,N_1620,N_306);
and U4179 (N_4179,N_2426,N_407);
and U4180 (N_4180,N_2019,N_1052);
or U4181 (N_4181,N_1330,N_2001);
and U4182 (N_4182,N_850,N_2495);
nand U4183 (N_4183,N_1689,N_1913);
nand U4184 (N_4184,N_647,N_2394);
nand U4185 (N_4185,N_707,N_804);
xor U4186 (N_4186,N_695,N_79);
and U4187 (N_4187,N_268,N_485);
or U4188 (N_4188,N_1524,N_36);
or U4189 (N_4189,N_164,N_523);
nor U4190 (N_4190,N_507,N_444);
and U4191 (N_4191,N_1653,N_648);
and U4192 (N_4192,N_3,N_373);
or U4193 (N_4193,N_225,N_969);
nor U4194 (N_4194,N_908,N_2259);
or U4195 (N_4195,N_623,N_2027);
nand U4196 (N_4196,N_1141,N_325);
and U4197 (N_4197,N_596,N_503);
nor U4198 (N_4198,N_1712,N_1355);
nor U4199 (N_4199,N_1282,N_1601);
and U4200 (N_4200,N_891,N_1141);
nand U4201 (N_4201,N_630,N_758);
nor U4202 (N_4202,N_643,N_62);
or U4203 (N_4203,N_507,N_944);
or U4204 (N_4204,N_204,N_997);
xor U4205 (N_4205,N_2069,N_1775);
and U4206 (N_4206,N_1443,N_758);
or U4207 (N_4207,N_2017,N_2210);
or U4208 (N_4208,N_284,N_1843);
nand U4209 (N_4209,N_703,N_1218);
or U4210 (N_4210,N_2114,N_324);
nor U4211 (N_4211,N_378,N_1528);
nor U4212 (N_4212,N_1308,N_1655);
nor U4213 (N_4213,N_2377,N_1104);
or U4214 (N_4214,N_1926,N_1032);
nand U4215 (N_4215,N_236,N_1385);
nand U4216 (N_4216,N_1086,N_600);
nor U4217 (N_4217,N_1874,N_1962);
or U4218 (N_4218,N_1530,N_1220);
and U4219 (N_4219,N_2076,N_2116);
and U4220 (N_4220,N_150,N_1639);
or U4221 (N_4221,N_203,N_2031);
nand U4222 (N_4222,N_884,N_1224);
nor U4223 (N_4223,N_1479,N_121);
nand U4224 (N_4224,N_2077,N_774);
and U4225 (N_4225,N_319,N_865);
nand U4226 (N_4226,N_238,N_1435);
and U4227 (N_4227,N_1414,N_1662);
nor U4228 (N_4228,N_2336,N_1157);
or U4229 (N_4229,N_1614,N_2412);
nand U4230 (N_4230,N_1850,N_143);
and U4231 (N_4231,N_683,N_2308);
nor U4232 (N_4232,N_2092,N_1527);
or U4233 (N_4233,N_1733,N_1562);
and U4234 (N_4234,N_529,N_721);
or U4235 (N_4235,N_1225,N_819);
and U4236 (N_4236,N_839,N_2082);
nor U4237 (N_4237,N_796,N_1373);
nand U4238 (N_4238,N_1708,N_2495);
nor U4239 (N_4239,N_2350,N_1537);
and U4240 (N_4240,N_2242,N_390);
nand U4241 (N_4241,N_556,N_73);
nand U4242 (N_4242,N_1698,N_1560);
nor U4243 (N_4243,N_601,N_1020);
nand U4244 (N_4244,N_962,N_752);
and U4245 (N_4245,N_2210,N_95);
or U4246 (N_4246,N_1354,N_936);
and U4247 (N_4247,N_1859,N_2124);
or U4248 (N_4248,N_2040,N_598);
or U4249 (N_4249,N_719,N_1699);
nor U4250 (N_4250,N_1466,N_1933);
and U4251 (N_4251,N_200,N_875);
or U4252 (N_4252,N_1076,N_2244);
nand U4253 (N_4253,N_721,N_454);
or U4254 (N_4254,N_638,N_1533);
and U4255 (N_4255,N_2280,N_2260);
or U4256 (N_4256,N_444,N_2197);
and U4257 (N_4257,N_1466,N_2305);
nor U4258 (N_4258,N_1242,N_215);
or U4259 (N_4259,N_1606,N_2041);
or U4260 (N_4260,N_1578,N_2304);
nor U4261 (N_4261,N_2255,N_1903);
and U4262 (N_4262,N_1431,N_749);
or U4263 (N_4263,N_1620,N_1533);
or U4264 (N_4264,N_1740,N_1319);
nor U4265 (N_4265,N_1506,N_1488);
nor U4266 (N_4266,N_1512,N_2446);
or U4267 (N_4267,N_1269,N_491);
and U4268 (N_4268,N_1066,N_1667);
nor U4269 (N_4269,N_248,N_1372);
nor U4270 (N_4270,N_2494,N_2334);
and U4271 (N_4271,N_980,N_409);
nor U4272 (N_4272,N_1801,N_2094);
nor U4273 (N_4273,N_1428,N_1513);
and U4274 (N_4274,N_68,N_2005);
and U4275 (N_4275,N_133,N_861);
or U4276 (N_4276,N_2060,N_1712);
and U4277 (N_4277,N_1572,N_672);
and U4278 (N_4278,N_2408,N_98);
or U4279 (N_4279,N_2353,N_1015);
or U4280 (N_4280,N_2336,N_360);
or U4281 (N_4281,N_2371,N_1926);
nor U4282 (N_4282,N_88,N_436);
nand U4283 (N_4283,N_1748,N_1248);
nor U4284 (N_4284,N_795,N_997);
nor U4285 (N_4285,N_703,N_1422);
and U4286 (N_4286,N_1837,N_250);
and U4287 (N_4287,N_2099,N_963);
and U4288 (N_4288,N_564,N_2039);
nor U4289 (N_4289,N_56,N_810);
nand U4290 (N_4290,N_916,N_258);
nand U4291 (N_4291,N_1340,N_407);
or U4292 (N_4292,N_1472,N_693);
or U4293 (N_4293,N_653,N_1677);
and U4294 (N_4294,N_886,N_2259);
nand U4295 (N_4295,N_2436,N_1776);
nand U4296 (N_4296,N_2358,N_1900);
nor U4297 (N_4297,N_1237,N_2060);
or U4298 (N_4298,N_1942,N_1803);
nand U4299 (N_4299,N_2002,N_1796);
nor U4300 (N_4300,N_265,N_1634);
or U4301 (N_4301,N_2156,N_156);
nor U4302 (N_4302,N_1459,N_779);
and U4303 (N_4303,N_2187,N_1806);
nand U4304 (N_4304,N_1338,N_1712);
nand U4305 (N_4305,N_1112,N_711);
and U4306 (N_4306,N_1590,N_1187);
nor U4307 (N_4307,N_1767,N_885);
xnor U4308 (N_4308,N_1760,N_402);
and U4309 (N_4309,N_2405,N_2020);
or U4310 (N_4310,N_1255,N_617);
or U4311 (N_4311,N_2412,N_1817);
nand U4312 (N_4312,N_1626,N_84);
nand U4313 (N_4313,N_113,N_1682);
or U4314 (N_4314,N_820,N_438);
and U4315 (N_4315,N_316,N_1530);
or U4316 (N_4316,N_942,N_1871);
nor U4317 (N_4317,N_2280,N_1371);
and U4318 (N_4318,N_861,N_1526);
nor U4319 (N_4319,N_1495,N_1443);
or U4320 (N_4320,N_1291,N_1862);
nand U4321 (N_4321,N_1986,N_559);
nor U4322 (N_4322,N_107,N_392);
or U4323 (N_4323,N_1692,N_177);
or U4324 (N_4324,N_364,N_1364);
nand U4325 (N_4325,N_570,N_2416);
and U4326 (N_4326,N_598,N_909);
and U4327 (N_4327,N_1800,N_1115);
and U4328 (N_4328,N_1485,N_382);
nor U4329 (N_4329,N_1534,N_2202);
or U4330 (N_4330,N_916,N_1942);
or U4331 (N_4331,N_1336,N_1613);
and U4332 (N_4332,N_1989,N_276);
nand U4333 (N_4333,N_1077,N_2112);
nand U4334 (N_4334,N_1365,N_2020);
and U4335 (N_4335,N_363,N_1848);
and U4336 (N_4336,N_2465,N_345);
or U4337 (N_4337,N_441,N_2284);
nor U4338 (N_4338,N_1518,N_204);
nor U4339 (N_4339,N_1481,N_147);
and U4340 (N_4340,N_1877,N_1503);
xnor U4341 (N_4341,N_1661,N_1233);
nand U4342 (N_4342,N_2352,N_2155);
nand U4343 (N_4343,N_496,N_314);
or U4344 (N_4344,N_51,N_2133);
nand U4345 (N_4345,N_893,N_360);
nor U4346 (N_4346,N_1580,N_2459);
or U4347 (N_4347,N_809,N_1623);
and U4348 (N_4348,N_1196,N_501);
and U4349 (N_4349,N_642,N_43);
or U4350 (N_4350,N_1087,N_2429);
nor U4351 (N_4351,N_2293,N_1410);
nor U4352 (N_4352,N_872,N_855);
and U4353 (N_4353,N_1483,N_742);
or U4354 (N_4354,N_1448,N_218);
or U4355 (N_4355,N_1100,N_1385);
nand U4356 (N_4356,N_2459,N_2225);
xnor U4357 (N_4357,N_532,N_2196);
nand U4358 (N_4358,N_2363,N_682);
nor U4359 (N_4359,N_784,N_1741);
nor U4360 (N_4360,N_1601,N_89);
nor U4361 (N_4361,N_2297,N_1289);
nand U4362 (N_4362,N_201,N_227);
and U4363 (N_4363,N_2470,N_1801);
or U4364 (N_4364,N_1375,N_2274);
nor U4365 (N_4365,N_1748,N_2405);
or U4366 (N_4366,N_2162,N_1805);
and U4367 (N_4367,N_106,N_1318);
nand U4368 (N_4368,N_930,N_1758);
nor U4369 (N_4369,N_1429,N_1489);
nand U4370 (N_4370,N_758,N_2080);
or U4371 (N_4371,N_297,N_372);
nor U4372 (N_4372,N_1839,N_1981);
nor U4373 (N_4373,N_1480,N_741);
nand U4374 (N_4374,N_673,N_1334);
nor U4375 (N_4375,N_428,N_1453);
nor U4376 (N_4376,N_206,N_1997);
and U4377 (N_4377,N_1810,N_1297);
and U4378 (N_4378,N_2188,N_1863);
and U4379 (N_4379,N_2390,N_19);
nor U4380 (N_4380,N_1116,N_2323);
nand U4381 (N_4381,N_2498,N_1769);
nand U4382 (N_4382,N_126,N_1359);
or U4383 (N_4383,N_582,N_1173);
or U4384 (N_4384,N_190,N_2041);
nor U4385 (N_4385,N_2037,N_1459);
or U4386 (N_4386,N_2459,N_2024);
or U4387 (N_4387,N_1931,N_1439);
nand U4388 (N_4388,N_2163,N_1858);
or U4389 (N_4389,N_1056,N_1777);
nor U4390 (N_4390,N_1896,N_2290);
and U4391 (N_4391,N_2315,N_2004);
nand U4392 (N_4392,N_2413,N_1504);
nand U4393 (N_4393,N_365,N_20);
nor U4394 (N_4394,N_2491,N_228);
and U4395 (N_4395,N_1920,N_250);
and U4396 (N_4396,N_382,N_2314);
nor U4397 (N_4397,N_2388,N_2417);
or U4398 (N_4398,N_2388,N_1902);
nand U4399 (N_4399,N_45,N_2385);
and U4400 (N_4400,N_396,N_627);
or U4401 (N_4401,N_379,N_2270);
or U4402 (N_4402,N_995,N_1265);
and U4403 (N_4403,N_776,N_742);
nand U4404 (N_4404,N_1523,N_1383);
nor U4405 (N_4405,N_2387,N_2315);
and U4406 (N_4406,N_2241,N_2350);
or U4407 (N_4407,N_2115,N_787);
or U4408 (N_4408,N_1528,N_1115);
nand U4409 (N_4409,N_162,N_540);
nor U4410 (N_4410,N_325,N_2215);
and U4411 (N_4411,N_1562,N_1369);
or U4412 (N_4412,N_1916,N_983);
nand U4413 (N_4413,N_214,N_1863);
nor U4414 (N_4414,N_2403,N_2118);
and U4415 (N_4415,N_1533,N_1341);
or U4416 (N_4416,N_2263,N_506);
nand U4417 (N_4417,N_1600,N_208);
nor U4418 (N_4418,N_1286,N_397);
or U4419 (N_4419,N_2481,N_603);
or U4420 (N_4420,N_1008,N_1085);
nor U4421 (N_4421,N_1528,N_1847);
or U4422 (N_4422,N_1719,N_490);
and U4423 (N_4423,N_1230,N_1);
or U4424 (N_4424,N_2098,N_2466);
and U4425 (N_4425,N_2300,N_1976);
nand U4426 (N_4426,N_110,N_220);
nor U4427 (N_4427,N_2028,N_936);
nor U4428 (N_4428,N_2103,N_2251);
or U4429 (N_4429,N_692,N_2360);
and U4430 (N_4430,N_1282,N_990);
or U4431 (N_4431,N_303,N_1188);
or U4432 (N_4432,N_700,N_613);
nor U4433 (N_4433,N_2088,N_1931);
and U4434 (N_4434,N_885,N_1092);
or U4435 (N_4435,N_1453,N_93);
and U4436 (N_4436,N_2206,N_1450);
nand U4437 (N_4437,N_2219,N_70);
nor U4438 (N_4438,N_1566,N_2289);
or U4439 (N_4439,N_247,N_31);
or U4440 (N_4440,N_1785,N_2093);
and U4441 (N_4441,N_520,N_1296);
nand U4442 (N_4442,N_1265,N_2153);
and U4443 (N_4443,N_1399,N_949);
or U4444 (N_4444,N_2248,N_451);
or U4445 (N_4445,N_1726,N_912);
nand U4446 (N_4446,N_215,N_1714);
nor U4447 (N_4447,N_635,N_231);
nand U4448 (N_4448,N_1970,N_204);
and U4449 (N_4449,N_2203,N_2090);
nand U4450 (N_4450,N_717,N_1682);
or U4451 (N_4451,N_1927,N_1698);
nor U4452 (N_4452,N_280,N_772);
nand U4453 (N_4453,N_235,N_132);
and U4454 (N_4454,N_407,N_1835);
and U4455 (N_4455,N_1687,N_1454);
and U4456 (N_4456,N_92,N_1213);
or U4457 (N_4457,N_831,N_268);
nor U4458 (N_4458,N_2493,N_212);
and U4459 (N_4459,N_428,N_411);
or U4460 (N_4460,N_1823,N_81);
or U4461 (N_4461,N_1870,N_1282);
and U4462 (N_4462,N_795,N_2399);
xnor U4463 (N_4463,N_1415,N_2030);
nor U4464 (N_4464,N_611,N_2200);
and U4465 (N_4465,N_1510,N_450);
nand U4466 (N_4466,N_1127,N_1717);
and U4467 (N_4467,N_2085,N_1969);
and U4468 (N_4468,N_1331,N_1068);
nor U4469 (N_4469,N_73,N_1705);
and U4470 (N_4470,N_714,N_1810);
nand U4471 (N_4471,N_2410,N_2460);
nor U4472 (N_4472,N_1772,N_1506);
or U4473 (N_4473,N_364,N_1962);
or U4474 (N_4474,N_1805,N_1275);
or U4475 (N_4475,N_2294,N_1909);
and U4476 (N_4476,N_1646,N_1219);
or U4477 (N_4477,N_2027,N_1573);
or U4478 (N_4478,N_2166,N_37);
nand U4479 (N_4479,N_73,N_897);
and U4480 (N_4480,N_465,N_453);
and U4481 (N_4481,N_454,N_786);
nor U4482 (N_4482,N_1496,N_733);
nor U4483 (N_4483,N_787,N_1475);
and U4484 (N_4484,N_875,N_2381);
nand U4485 (N_4485,N_584,N_124);
and U4486 (N_4486,N_661,N_1042);
and U4487 (N_4487,N_1321,N_1169);
or U4488 (N_4488,N_802,N_480);
and U4489 (N_4489,N_1496,N_567);
nand U4490 (N_4490,N_1418,N_1099);
or U4491 (N_4491,N_58,N_1402);
or U4492 (N_4492,N_1357,N_1147);
and U4493 (N_4493,N_805,N_1756);
nand U4494 (N_4494,N_856,N_532);
nand U4495 (N_4495,N_1877,N_1886);
or U4496 (N_4496,N_208,N_2128);
nor U4497 (N_4497,N_0,N_180);
and U4498 (N_4498,N_1685,N_477);
nor U4499 (N_4499,N_67,N_2255);
nand U4500 (N_4500,N_684,N_1946);
nand U4501 (N_4501,N_44,N_1405);
nand U4502 (N_4502,N_2022,N_2073);
and U4503 (N_4503,N_1861,N_208);
or U4504 (N_4504,N_2051,N_284);
or U4505 (N_4505,N_1598,N_1042);
nand U4506 (N_4506,N_2300,N_2047);
nand U4507 (N_4507,N_1654,N_776);
nor U4508 (N_4508,N_170,N_693);
nor U4509 (N_4509,N_1418,N_309);
nand U4510 (N_4510,N_1914,N_1335);
xor U4511 (N_4511,N_1471,N_1601);
nand U4512 (N_4512,N_973,N_34);
xnor U4513 (N_4513,N_2433,N_1938);
nor U4514 (N_4514,N_773,N_1126);
nor U4515 (N_4515,N_983,N_1211);
or U4516 (N_4516,N_1307,N_672);
nand U4517 (N_4517,N_1574,N_2430);
nand U4518 (N_4518,N_1714,N_1797);
nand U4519 (N_4519,N_1160,N_1903);
nor U4520 (N_4520,N_395,N_2311);
and U4521 (N_4521,N_1956,N_1197);
or U4522 (N_4522,N_2393,N_292);
nor U4523 (N_4523,N_882,N_1264);
nor U4524 (N_4524,N_1134,N_1430);
or U4525 (N_4525,N_259,N_908);
or U4526 (N_4526,N_996,N_1844);
or U4527 (N_4527,N_558,N_1140);
and U4528 (N_4528,N_2001,N_501);
or U4529 (N_4529,N_168,N_2027);
nor U4530 (N_4530,N_468,N_2187);
nor U4531 (N_4531,N_1548,N_970);
or U4532 (N_4532,N_1638,N_2279);
nand U4533 (N_4533,N_794,N_2250);
or U4534 (N_4534,N_152,N_1385);
or U4535 (N_4535,N_1065,N_2379);
or U4536 (N_4536,N_2059,N_759);
and U4537 (N_4537,N_453,N_1156);
nand U4538 (N_4538,N_927,N_2373);
nor U4539 (N_4539,N_492,N_1019);
or U4540 (N_4540,N_494,N_874);
nand U4541 (N_4541,N_2373,N_777);
nand U4542 (N_4542,N_527,N_931);
or U4543 (N_4543,N_1820,N_371);
nor U4544 (N_4544,N_2470,N_184);
and U4545 (N_4545,N_1043,N_1992);
or U4546 (N_4546,N_107,N_947);
nand U4547 (N_4547,N_222,N_2272);
and U4548 (N_4548,N_685,N_1583);
and U4549 (N_4549,N_440,N_1193);
or U4550 (N_4550,N_587,N_2362);
nand U4551 (N_4551,N_2297,N_936);
or U4552 (N_4552,N_683,N_1240);
nand U4553 (N_4553,N_1203,N_1031);
nand U4554 (N_4554,N_1971,N_1333);
nand U4555 (N_4555,N_689,N_624);
nor U4556 (N_4556,N_125,N_1507);
nor U4557 (N_4557,N_1046,N_1525);
and U4558 (N_4558,N_2218,N_190);
or U4559 (N_4559,N_1239,N_1086);
or U4560 (N_4560,N_237,N_900);
and U4561 (N_4561,N_269,N_2294);
nand U4562 (N_4562,N_43,N_1199);
or U4563 (N_4563,N_68,N_192);
nand U4564 (N_4564,N_2123,N_992);
nor U4565 (N_4565,N_1239,N_2305);
or U4566 (N_4566,N_990,N_2308);
or U4567 (N_4567,N_1120,N_2415);
and U4568 (N_4568,N_436,N_905);
nand U4569 (N_4569,N_514,N_1413);
or U4570 (N_4570,N_745,N_2111);
or U4571 (N_4571,N_2311,N_1860);
nor U4572 (N_4572,N_1872,N_62);
nand U4573 (N_4573,N_181,N_173);
nand U4574 (N_4574,N_194,N_2410);
nand U4575 (N_4575,N_34,N_951);
or U4576 (N_4576,N_325,N_62);
nand U4577 (N_4577,N_1215,N_235);
or U4578 (N_4578,N_2060,N_738);
and U4579 (N_4579,N_2299,N_1242);
nand U4580 (N_4580,N_323,N_1518);
nor U4581 (N_4581,N_398,N_754);
nor U4582 (N_4582,N_1194,N_1369);
nor U4583 (N_4583,N_531,N_299);
or U4584 (N_4584,N_484,N_203);
or U4585 (N_4585,N_1416,N_563);
nand U4586 (N_4586,N_790,N_1480);
or U4587 (N_4587,N_2033,N_2290);
or U4588 (N_4588,N_618,N_652);
or U4589 (N_4589,N_2056,N_1880);
nand U4590 (N_4590,N_2431,N_2216);
or U4591 (N_4591,N_1378,N_1630);
or U4592 (N_4592,N_1924,N_2107);
nand U4593 (N_4593,N_2399,N_468);
nor U4594 (N_4594,N_2166,N_1931);
and U4595 (N_4595,N_307,N_214);
and U4596 (N_4596,N_1245,N_1223);
xor U4597 (N_4597,N_555,N_1612);
nand U4598 (N_4598,N_1939,N_1260);
or U4599 (N_4599,N_180,N_2008);
nor U4600 (N_4600,N_1073,N_1800);
and U4601 (N_4601,N_2059,N_1550);
nor U4602 (N_4602,N_441,N_858);
nor U4603 (N_4603,N_305,N_2278);
and U4604 (N_4604,N_2052,N_954);
nand U4605 (N_4605,N_2143,N_1831);
and U4606 (N_4606,N_1441,N_1291);
nor U4607 (N_4607,N_2170,N_569);
or U4608 (N_4608,N_2228,N_2107);
nand U4609 (N_4609,N_1733,N_1182);
and U4610 (N_4610,N_296,N_26);
nand U4611 (N_4611,N_1539,N_453);
and U4612 (N_4612,N_771,N_1997);
nand U4613 (N_4613,N_24,N_2394);
or U4614 (N_4614,N_1404,N_653);
nand U4615 (N_4615,N_2011,N_1642);
nand U4616 (N_4616,N_1739,N_767);
nand U4617 (N_4617,N_1590,N_1662);
or U4618 (N_4618,N_1110,N_22);
or U4619 (N_4619,N_717,N_485);
or U4620 (N_4620,N_1627,N_704);
or U4621 (N_4621,N_1055,N_430);
nor U4622 (N_4622,N_294,N_1859);
or U4623 (N_4623,N_1968,N_1784);
nor U4624 (N_4624,N_1126,N_1650);
xor U4625 (N_4625,N_1738,N_1394);
nor U4626 (N_4626,N_1354,N_680);
and U4627 (N_4627,N_2362,N_1296);
nor U4628 (N_4628,N_62,N_1620);
nor U4629 (N_4629,N_83,N_2318);
nand U4630 (N_4630,N_2291,N_1623);
or U4631 (N_4631,N_1842,N_2007);
and U4632 (N_4632,N_2377,N_1406);
and U4633 (N_4633,N_1081,N_958);
nor U4634 (N_4634,N_579,N_2218);
or U4635 (N_4635,N_2233,N_1966);
nor U4636 (N_4636,N_1502,N_531);
or U4637 (N_4637,N_1387,N_823);
nand U4638 (N_4638,N_1180,N_2481);
nand U4639 (N_4639,N_1049,N_325);
or U4640 (N_4640,N_1019,N_1630);
nand U4641 (N_4641,N_169,N_425);
or U4642 (N_4642,N_1192,N_1317);
nor U4643 (N_4643,N_2394,N_1064);
nor U4644 (N_4644,N_1860,N_1296);
nand U4645 (N_4645,N_2002,N_1423);
nand U4646 (N_4646,N_1436,N_1717);
nor U4647 (N_4647,N_1815,N_2454);
nand U4648 (N_4648,N_1236,N_1999);
nor U4649 (N_4649,N_103,N_1814);
and U4650 (N_4650,N_1417,N_1810);
or U4651 (N_4651,N_1364,N_799);
or U4652 (N_4652,N_868,N_1295);
or U4653 (N_4653,N_346,N_2381);
and U4654 (N_4654,N_1393,N_981);
and U4655 (N_4655,N_1488,N_827);
or U4656 (N_4656,N_1869,N_1984);
and U4657 (N_4657,N_166,N_561);
and U4658 (N_4658,N_2132,N_1244);
and U4659 (N_4659,N_1710,N_1808);
nand U4660 (N_4660,N_2146,N_279);
nand U4661 (N_4661,N_1604,N_2349);
nand U4662 (N_4662,N_1849,N_1126);
nand U4663 (N_4663,N_882,N_1713);
nand U4664 (N_4664,N_1895,N_1084);
or U4665 (N_4665,N_1432,N_1522);
or U4666 (N_4666,N_1024,N_2333);
nand U4667 (N_4667,N_303,N_509);
nor U4668 (N_4668,N_1784,N_384);
nor U4669 (N_4669,N_2464,N_1009);
nand U4670 (N_4670,N_2097,N_1478);
nand U4671 (N_4671,N_1778,N_584);
or U4672 (N_4672,N_2264,N_1424);
and U4673 (N_4673,N_554,N_742);
nor U4674 (N_4674,N_2456,N_2445);
nor U4675 (N_4675,N_185,N_2396);
nor U4676 (N_4676,N_916,N_893);
and U4677 (N_4677,N_1253,N_933);
nor U4678 (N_4678,N_2466,N_1375);
nor U4679 (N_4679,N_1615,N_2180);
and U4680 (N_4680,N_1023,N_443);
or U4681 (N_4681,N_2380,N_1752);
nand U4682 (N_4682,N_1298,N_1653);
nand U4683 (N_4683,N_1040,N_1015);
or U4684 (N_4684,N_683,N_1416);
nor U4685 (N_4685,N_63,N_158);
nand U4686 (N_4686,N_2462,N_1688);
nor U4687 (N_4687,N_1628,N_2129);
nand U4688 (N_4688,N_499,N_736);
and U4689 (N_4689,N_1327,N_2347);
or U4690 (N_4690,N_751,N_1717);
nand U4691 (N_4691,N_721,N_903);
and U4692 (N_4692,N_307,N_1251);
nand U4693 (N_4693,N_1855,N_2267);
nand U4694 (N_4694,N_2033,N_2231);
or U4695 (N_4695,N_404,N_2209);
and U4696 (N_4696,N_547,N_735);
and U4697 (N_4697,N_190,N_1655);
xor U4698 (N_4698,N_1519,N_646);
nor U4699 (N_4699,N_2144,N_672);
nand U4700 (N_4700,N_1891,N_2250);
and U4701 (N_4701,N_1785,N_1842);
or U4702 (N_4702,N_1056,N_1554);
nand U4703 (N_4703,N_666,N_1239);
nand U4704 (N_4704,N_1121,N_605);
and U4705 (N_4705,N_1543,N_401);
nand U4706 (N_4706,N_1767,N_1895);
nand U4707 (N_4707,N_1121,N_322);
or U4708 (N_4708,N_45,N_2053);
nand U4709 (N_4709,N_2084,N_58);
nand U4710 (N_4710,N_1743,N_801);
nand U4711 (N_4711,N_76,N_1133);
nor U4712 (N_4712,N_154,N_1711);
or U4713 (N_4713,N_1066,N_1819);
nand U4714 (N_4714,N_718,N_336);
nor U4715 (N_4715,N_191,N_2200);
nor U4716 (N_4716,N_417,N_1180);
or U4717 (N_4717,N_1084,N_389);
nor U4718 (N_4718,N_418,N_1618);
nand U4719 (N_4719,N_587,N_1723);
nand U4720 (N_4720,N_1825,N_2072);
nor U4721 (N_4721,N_721,N_199);
or U4722 (N_4722,N_1973,N_2211);
nand U4723 (N_4723,N_1738,N_866);
or U4724 (N_4724,N_2412,N_1367);
and U4725 (N_4725,N_2436,N_2068);
nand U4726 (N_4726,N_2133,N_2257);
and U4727 (N_4727,N_2123,N_381);
nand U4728 (N_4728,N_2426,N_2095);
or U4729 (N_4729,N_500,N_2479);
and U4730 (N_4730,N_1237,N_488);
nand U4731 (N_4731,N_542,N_1500);
nor U4732 (N_4732,N_579,N_1341);
or U4733 (N_4733,N_594,N_510);
nand U4734 (N_4734,N_1455,N_1888);
nand U4735 (N_4735,N_896,N_2003);
and U4736 (N_4736,N_187,N_1550);
and U4737 (N_4737,N_407,N_171);
and U4738 (N_4738,N_2021,N_542);
and U4739 (N_4739,N_620,N_2065);
nor U4740 (N_4740,N_899,N_1399);
nor U4741 (N_4741,N_1728,N_1182);
nand U4742 (N_4742,N_1188,N_1839);
or U4743 (N_4743,N_722,N_2370);
nor U4744 (N_4744,N_2268,N_1771);
or U4745 (N_4745,N_1752,N_1024);
nor U4746 (N_4746,N_1438,N_253);
or U4747 (N_4747,N_1239,N_632);
nor U4748 (N_4748,N_939,N_911);
or U4749 (N_4749,N_53,N_2083);
nor U4750 (N_4750,N_1767,N_113);
or U4751 (N_4751,N_2491,N_2108);
and U4752 (N_4752,N_2241,N_1750);
nand U4753 (N_4753,N_2169,N_236);
and U4754 (N_4754,N_477,N_1020);
or U4755 (N_4755,N_518,N_1586);
or U4756 (N_4756,N_1302,N_936);
nand U4757 (N_4757,N_1594,N_2472);
and U4758 (N_4758,N_2113,N_106);
nor U4759 (N_4759,N_1564,N_237);
xnor U4760 (N_4760,N_432,N_1592);
nand U4761 (N_4761,N_2169,N_816);
or U4762 (N_4762,N_1654,N_831);
nand U4763 (N_4763,N_1856,N_1483);
nand U4764 (N_4764,N_2169,N_1914);
nor U4765 (N_4765,N_1375,N_1577);
and U4766 (N_4766,N_315,N_41);
nor U4767 (N_4767,N_654,N_2252);
or U4768 (N_4768,N_697,N_1772);
xnor U4769 (N_4769,N_533,N_1989);
nand U4770 (N_4770,N_1069,N_294);
nor U4771 (N_4771,N_1808,N_382);
nand U4772 (N_4772,N_612,N_652);
and U4773 (N_4773,N_1256,N_1074);
nand U4774 (N_4774,N_2105,N_207);
and U4775 (N_4775,N_1343,N_837);
nor U4776 (N_4776,N_1751,N_2293);
and U4777 (N_4777,N_2178,N_1001);
nand U4778 (N_4778,N_1109,N_2445);
nand U4779 (N_4779,N_161,N_2405);
and U4780 (N_4780,N_2492,N_2340);
or U4781 (N_4781,N_1715,N_1363);
nand U4782 (N_4782,N_1539,N_756);
nor U4783 (N_4783,N_1175,N_2306);
nand U4784 (N_4784,N_1536,N_1286);
nor U4785 (N_4785,N_10,N_2307);
nand U4786 (N_4786,N_390,N_1820);
nor U4787 (N_4787,N_2493,N_1216);
nor U4788 (N_4788,N_1990,N_1639);
or U4789 (N_4789,N_1287,N_2147);
and U4790 (N_4790,N_168,N_941);
nand U4791 (N_4791,N_501,N_1042);
and U4792 (N_4792,N_1090,N_2205);
nand U4793 (N_4793,N_1269,N_628);
or U4794 (N_4794,N_1208,N_1121);
or U4795 (N_4795,N_303,N_1425);
nor U4796 (N_4796,N_1232,N_547);
nor U4797 (N_4797,N_694,N_196);
xor U4798 (N_4798,N_731,N_1017);
or U4799 (N_4799,N_1283,N_1418);
or U4800 (N_4800,N_2128,N_197);
nand U4801 (N_4801,N_759,N_937);
nor U4802 (N_4802,N_2294,N_885);
or U4803 (N_4803,N_256,N_1003);
or U4804 (N_4804,N_1770,N_1567);
nor U4805 (N_4805,N_436,N_2345);
nand U4806 (N_4806,N_1741,N_1080);
and U4807 (N_4807,N_44,N_2472);
nand U4808 (N_4808,N_697,N_358);
nand U4809 (N_4809,N_475,N_347);
nor U4810 (N_4810,N_988,N_2259);
nand U4811 (N_4811,N_1992,N_1111);
nand U4812 (N_4812,N_348,N_1199);
and U4813 (N_4813,N_1305,N_2127);
nor U4814 (N_4814,N_1886,N_1066);
nand U4815 (N_4815,N_372,N_1865);
or U4816 (N_4816,N_1237,N_1434);
nor U4817 (N_4817,N_1246,N_695);
xor U4818 (N_4818,N_722,N_1677);
nor U4819 (N_4819,N_436,N_517);
nor U4820 (N_4820,N_1446,N_2313);
and U4821 (N_4821,N_205,N_1379);
or U4822 (N_4822,N_1366,N_757);
and U4823 (N_4823,N_1491,N_1670);
nor U4824 (N_4824,N_53,N_1612);
nor U4825 (N_4825,N_2101,N_2405);
nor U4826 (N_4826,N_1844,N_961);
nand U4827 (N_4827,N_872,N_2003);
or U4828 (N_4828,N_515,N_433);
nor U4829 (N_4829,N_1554,N_1072);
nand U4830 (N_4830,N_2217,N_461);
nand U4831 (N_4831,N_1927,N_520);
and U4832 (N_4832,N_2347,N_1444);
and U4833 (N_4833,N_1045,N_1372);
and U4834 (N_4834,N_706,N_106);
nand U4835 (N_4835,N_1048,N_1206);
or U4836 (N_4836,N_1858,N_1135);
nand U4837 (N_4837,N_2465,N_2380);
or U4838 (N_4838,N_956,N_2293);
or U4839 (N_4839,N_1079,N_1608);
or U4840 (N_4840,N_1506,N_1640);
and U4841 (N_4841,N_2217,N_2312);
and U4842 (N_4842,N_347,N_2075);
nand U4843 (N_4843,N_651,N_2222);
nor U4844 (N_4844,N_691,N_164);
or U4845 (N_4845,N_1329,N_1670);
nand U4846 (N_4846,N_1069,N_1334);
nand U4847 (N_4847,N_112,N_1683);
and U4848 (N_4848,N_1523,N_2);
and U4849 (N_4849,N_1126,N_1134);
or U4850 (N_4850,N_2294,N_1160);
nor U4851 (N_4851,N_2487,N_1680);
and U4852 (N_4852,N_2492,N_2213);
or U4853 (N_4853,N_1346,N_67);
or U4854 (N_4854,N_1472,N_700);
or U4855 (N_4855,N_1831,N_230);
nand U4856 (N_4856,N_1019,N_1218);
or U4857 (N_4857,N_1563,N_2117);
nand U4858 (N_4858,N_1444,N_1373);
xor U4859 (N_4859,N_1361,N_342);
or U4860 (N_4860,N_683,N_302);
and U4861 (N_4861,N_1820,N_1909);
nor U4862 (N_4862,N_1733,N_1653);
nor U4863 (N_4863,N_548,N_2470);
and U4864 (N_4864,N_359,N_1964);
or U4865 (N_4865,N_1271,N_1099);
nor U4866 (N_4866,N_1654,N_346);
nor U4867 (N_4867,N_143,N_1943);
or U4868 (N_4868,N_2427,N_1056);
nor U4869 (N_4869,N_960,N_1069);
nand U4870 (N_4870,N_1599,N_1359);
nor U4871 (N_4871,N_61,N_2071);
nor U4872 (N_4872,N_103,N_340);
nor U4873 (N_4873,N_72,N_1469);
nand U4874 (N_4874,N_640,N_1763);
or U4875 (N_4875,N_1758,N_1491);
nor U4876 (N_4876,N_1860,N_1496);
or U4877 (N_4877,N_872,N_1059);
nand U4878 (N_4878,N_1709,N_396);
or U4879 (N_4879,N_1642,N_601);
and U4880 (N_4880,N_711,N_634);
xor U4881 (N_4881,N_249,N_483);
and U4882 (N_4882,N_162,N_300);
nand U4883 (N_4883,N_184,N_1279);
nand U4884 (N_4884,N_2187,N_1199);
or U4885 (N_4885,N_531,N_2163);
nand U4886 (N_4886,N_593,N_2028);
or U4887 (N_4887,N_1820,N_1120);
or U4888 (N_4888,N_239,N_1265);
nor U4889 (N_4889,N_650,N_2201);
or U4890 (N_4890,N_2167,N_1471);
nand U4891 (N_4891,N_1339,N_211);
or U4892 (N_4892,N_514,N_438);
nand U4893 (N_4893,N_1124,N_1804);
nand U4894 (N_4894,N_1295,N_825);
nand U4895 (N_4895,N_1378,N_1796);
nand U4896 (N_4896,N_897,N_672);
and U4897 (N_4897,N_2214,N_115);
nand U4898 (N_4898,N_569,N_1181);
or U4899 (N_4899,N_1996,N_920);
or U4900 (N_4900,N_659,N_272);
or U4901 (N_4901,N_820,N_19);
and U4902 (N_4902,N_1481,N_1756);
or U4903 (N_4903,N_2217,N_1983);
or U4904 (N_4904,N_83,N_250);
or U4905 (N_4905,N_1083,N_96);
and U4906 (N_4906,N_966,N_2351);
nor U4907 (N_4907,N_1063,N_627);
and U4908 (N_4908,N_823,N_2463);
or U4909 (N_4909,N_493,N_123);
or U4910 (N_4910,N_1150,N_177);
nand U4911 (N_4911,N_463,N_546);
and U4912 (N_4912,N_2254,N_1399);
nand U4913 (N_4913,N_320,N_2013);
nand U4914 (N_4914,N_741,N_2053);
nand U4915 (N_4915,N_1157,N_2273);
or U4916 (N_4916,N_2426,N_300);
or U4917 (N_4917,N_1999,N_1376);
and U4918 (N_4918,N_737,N_2010);
and U4919 (N_4919,N_91,N_1);
nand U4920 (N_4920,N_411,N_25);
nor U4921 (N_4921,N_596,N_484);
nor U4922 (N_4922,N_1960,N_1726);
and U4923 (N_4923,N_2063,N_2323);
and U4924 (N_4924,N_235,N_1835);
nor U4925 (N_4925,N_768,N_1284);
nor U4926 (N_4926,N_1711,N_2059);
nand U4927 (N_4927,N_2020,N_874);
and U4928 (N_4928,N_1123,N_704);
nand U4929 (N_4929,N_697,N_1636);
and U4930 (N_4930,N_1202,N_797);
nand U4931 (N_4931,N_2483,N_1030);
and U4932 (N_4932,N_630,N_2333);
nor U4933 (N_4933,N_2379,N_2030);
nor U4934 (N_4934,N_1537,N_2216);
or U4935 (N_4935,N_1920,N_1959);
or U4936 (N_4936,N_1086,N_847);
nor U4937 (N_4937,N_806,N_2210);
nand U4938 (N_4938,N_1679,N_1377);
nor U4939 (N_4939,N_294,N_1691);
nand U4940 (N_4940,N_2026,N_826);
and U4941 (N_4941,N_16,N_277);
nand U4942 (N_4942,N_727,N_712);
and U4943 (N_4943,N_728,N_1817);
nor U4944 (N_4944,N_2196,N_889);
and U4945 (N_4945,N_595,N_1777);
nor U4946 (N_4946,N_1886,N_740);
and U4947 (N_4947,N_554,N_1588);
or U4948 (N_4948,N_1369,N_119);
nand U4949 (N_4949,N_1161,N_158);
and U4950 (N_4950,N_1047,N_1271);
nand U4951 (N_4951,N_702,N_1024);
nand U4952 (N_4952,N_1372,N_667);
nand U4953 (N_4953,N_500,N_805);
and U4954 (N_4954,N_1824,N_836);
nand U4955 (N_4955,N_850,N_1006);
or U4956 (N_4956,N_1885,N_1435);
or U4957 (N_4957,N_2120,N_1538);
and U4958 (N_4958,N_905,N_1169);
nor U4959 (N_4959,N_826,N_1341);
nor U4960 (N_4960,N_255,N_2301);
or U4961 (N_4961,N_2114,N_490);
and U4962 (N_4962,N_1980,N_29);
nor U4963 (N_4963,N_839,N_1468);
nand U4964 (N_4964,N_1083,N_602);
or U4965 (N_4965,N_279,N_909);
xor U4966 (N_4966,N_2317,N_1290);
nor U4967 (N_4967,N_549,N_2487);
nand U4968 (N_4968,N_1787,N_590);
or U4969 (N_4969,N_2022,N_762);
and U4970 (N_4970,N_1141,N_37);
nor U4971 (N_4971,N_1968,N_2048);
and U4972 (N_4972,N_2047,N_65);
nor U4973 (N_4973,N_1205,N_853);
and U4974 (N_4974,N_338,N_960);
and U4975 (N_4975,N_547,N_641);
or U4976 (N_4976,N_1116,N_1085);
and U4977 (N_4977,N_1033,N_2082);
or U4978 (N_4978,N_2010,N_1001);
and U4979 (N_4979,N_1153,N_2067);
nand U4980 (N_4980,N_675,N_416);
and U4981 (N_4981,N_344,N_1425);
and U4982 (N_4982,N_1093,N_1249);
and U4983 (N_4983,N_561,N_2492);
nor U4984 (N_4984,N_354,N_1017);
nor U4985 (N_4985,N_2478,N_1825);
or U4986 (N_4986,N_1695,N_1340);
or U4987 (N_4987,N_1074,N_1241);
or U4988 (N_4988,N_234,N_279);
nand U4989 (N_4989,N_1786,N_1151);
or U4990 (N_4990,N_2095,N_286);
nand U4991 (N_4991,N_951,N_217);
and U4992 (N_4992,N_1538,N_93);
or U4993 (N_4993,N_963,N_1992);
and U4994 (N_4994,N_2267,N_1066);
nand U4995 (N_4995,N_458,N_701);
nand U4996 (N_4996,N_2061,N_1520);
and U4997 (N_4997,N_298,N_1164);
and U4998 (N_4998,N_1933,N_1352);
nand U4999 (N_4999,N_916,N_2433);
nor U5000 (N_5000,N_2502,N_4851);
or U5001 (N_5001,N_4212,N_4073);
and U5002 (N_5002,N_3758,N_2725);
nand U5003 (N_5003,N_3637,N_3396);
and U5004 (N_5004,N_4028,N_3827);
nand U5005 (N_5005,N_3529,N_4251);
nand U5006 (N_5006,N_2604,N_3669);
nand U5007 (N_5007,N_3777,N_3711);
and U5008 (N_5008,N_3653,N_3883);
and U5009 (N_5009,N_3083,N_4164);
nor U5010 (N_5010,N_3671,N_3029);
or U5011 (N_5011,N_4126,N_2510);
nor U5012 (N_5012,N_4962,N_2576);
nand U5013 (N_5013,N_4849,N_3231);
and U5014 (N_5014,N_2799,N_3884);
and U5015 (N_5015,N_3489,N_2930);
nor U5016 (N_5016,N_4972,N_3795);
or U5017 (N_5017,N_4238,N_2951);
and U5018 (N_5018,N_3522,N_4348);
nand U5019 (N_5019,N_3076,N_3215);
nand U5020 (N_5020,N_3324,N_3689);
and U5021 (N_5021,N_4135,N_3280);
or U5022 (N_5022,N_3276,N_4436);
or U5023 (N_5023,N_3935,N_3882);
xor U5024 (N_5024,N_3577,N_4969);
and U5025 (N_5025,N_4020,N_3414);
nand U5026 (N_5026,N_3038,N_4258);
nand U5027 (N_5027,N_4506,N_4247);
or U5028 (N_5028,N_2997,N_3063);
and U5029 (N_5029,N_4374,N_2609);
nor U5030 (N_5030,N_3971,N_3184);
or U5031 (N_5031,N_2505,N_4694);
nor U5032 (N_5032,N_3298,N_2732);
nor U5033 (N_5033,N_3739,N_4669);
and U5034 (N_5034,N_4572,N_3846);
nor U5035 (N_5035,N_3997,N_3850);
nor U5036 (N_5036,N_2612,N_2824);
nor U5037 (N_5037,N_3956,N_4958);
nand U5038 (N_5038,N_4625,N_4954);
and U5039 (N_5039,N_3273,N_4319);
nand U5040 (N_5040,N_3514,N_4553);
nand U5041 (N_5041,N_4057,N_4529);
nor U5042 (N_5042,N_4875,N_3830);
nor U5043 (N_5043,N_4353,N_3047);
nand U5044 (N_5044,N_3111,N_4573);
nand U5045 (N_5045,N_4086,N_4205);
or U5046 (N_5046,N_4216,N_2896);
and U5047 (N_5047,N_2961,N_4167);
nand U5048 (N_5048,N_3761,N_4383);
and U5049 (N_5049,N_3246,N_4062);
nor U5050 (N_5050,N_4345,N_4880);
nand U5051 (N_5051,N_2787,N_3542);
or U5052 (N_5052,N_3188,N_3318);
nand U5053 (N_5053,N_4366,N_2808);
nor U5054 (N_5054,N_3286,N_3892);
nand U5055 (N_5055,N_3574,N_4037);
and U5056 (N_5056,N_2971,N_4809);
nand U5057 (N_5057,N_2722,N_4194);
and U5058 (N_5058,N_4059,N_3960);
and U5059 (N_5059,N_3364,N_3617);
or U5060 (N_5060,N_3311,N_2914);
or U5061 (N_5061,N_3948,N_4261);
and U5062 (N_5062,N_4523,N_2897);
nand U5063 (N_5063,N_2624,N_4598);
and U5064 (N_5064,N_4481,N_4600);
or U5065 (N_5065,N_2641,N_3566);
or U5066 (N_5066,N_3423,N_4977);
and U5067 (N_5067,N_3167,N_4584);
and U5068 (N_5068,N_2689,N_2955);
nand U5069 (N_5069,N_4489,N_4505);
and U5070 (N_5070,N_4510,N_3419);
or U5071 (N_5071,N_3260,N_4555);
or U5072 (N_5072,N_2585,N_3752);
or U5073 (N_5073,N_3282,N_3572);
or U5074 (N_5074,N_3141,N_3980);
or U5075 (N_5075,N_3170,N_4372);
or U5076 (N_5076,N_4437,N_4661);
nor U5077 (N_5077,N_4776,N_4961);
or U5078 (N_5078,N_3274,N_3564);
nor U5079 (N_5079,N_3943,N_4341);
nand U5080 (N_5080,N_2775,N_4796);
or U5081 (N_5081,N_3779,N_4960);
nor U5082 (N_5082,N_4400,N_3261);
nor U5083 (N_5083,N_3908,N_4351);
nor U5084 (N_5084,N_4861,N_3180);
nor U5085 (N_5085,N_3493,N_2654);
or U5086 (N_5086,N_4690,N_2621);
and U5087 (N_5087,N_2786,N_4454);
and U5088 (N_5088,N_3648,N_2942);
nand U5089 (N_5089,N_4778,N_3057);
or U5090 (N_5090,N_4340,N_2635);
nor U5091 (N_5091,N_2707,N_4603);
or U5092 (N_5092,N_3148,N_2773);
or U5093 (N_5093,N_4065,N_3426);
nand U5094 (N_5094,N_3309,N_4482);
or U5095 (N_5095,N_2927,N_4906);
and U5096 (N_5096,N_3343,N_3152);
or U5097 (N_5097,N_2593,N_4492);
nor U5098 (N_5098,N_4330,N_3270);
nand U5099 (N_5099,N_2757,N_2628);
nor U5100 (N_5100,N_4200,N_3305);
nor U5101 (N_5101,N_3291,N_3622);
or U5102 (N_5102,N_2868,N_4871);
nand U5103 (N_5103,N_4434,N_3374);
nor U5104 (N_5104,N_4180,N_3645);
nand U5105 (N_5105,N_2727,N_3510);
or U5106 (N_5106,N_3536,N_2771);
or U5107 (N_5107,N_2573,N_3046);
nor U5108 (N_5108,N_3609,N_4371);
or U5109 (N_5109,N_4605,N_4166);
and U5110 (N_5110,N_2873,N_4344);
or U5111 (N_5111,N_3546,N_4987);
or U5112 (N_5112,N_4772,N_2848);
nand U5113 (N_5113,N_3904,N_3495);
nand U5114 (N_5114,N_2895,N_3719);
or U5115 (N_5115,N_2846,N_2575);
nand U5116 (N_5116,N_3920,N_3154);
or U5117 (N_5117,N_2945,N_4115);
and U5118 (N_5118,N_3941,N_4269);
and U5119 (N_5119,N_4663,N_2683);
nand U5120 (N_5120,N_3857,N_3266);
and U5121 (N_5121,N_4445,N_4373);
and U5122 (N_5122,N_4362,N_4633);
and U5123 (N_5123,N_3762,N_4550);
or U5124 (N_5124,N_4222,N_4827);
nand U5125 (N_5125,N_3936,N_4939);
and U5126 (N_5126,N_2640,N_3604);
or U5127 (N_5127,N_4545,N_3297);
nand U5128 (N_5128,N_2687,N_2948);
nand U5129 (N_5129,N_4936,N_4350);
nand U5130 (N_5130,N_4485,N_4302);
nand U5131 (N_5131,N_3796,N_2867);
nor U5132 (N_5132,N_4324,N_2507);
and U5133 (N_5133,N_2923,N_4855);
nor U5134 (N_5134,N_3547,N_3443);
nor U5135 (N_5135,N_2605,N_4478);
and U5136 (N_5136,N_3627,N_3717);
and U5137 (N_5137,N_4322,N_2835);
nand U5138 (N_5138,N_3558,N_2663);
and U5139 (N_5139,N_3050,N_3766);
or U5140 (N_5140,N_4512,N_4068);
or U5141 (N_5141,N_4380,N_2550);
and U5142 (N_5142,N_4092,N_3650);
xor U5143 (N_5143,N_4777,N_2639);
or U5144 (N_5144,N_2847,N_4432);
or U5145 (N_5145,N_2552,N_2764);
and U5146 (N_5146,N_2519,N_3649);
or U5147 (N_5147,N_2840,N_4081);
and U5148 (N_5148,N_4655,N_3416);
and U5149 (N_5149,N_3596,N_3737);
or U5150 (N_5150,N_4027,N_4475);
or U5151 (N_5151,N_3687,N_4365);
and U5152 (N_5152,N_4786,N_3177);
or U5153 (N_5153,N_4779,N_2857);
nand U5154 (N_5154,N_3683,N_4812);
nor U5155 (N_5155,N_3285,N_3483);
and U5156 (N_5156,N_3565,N_4336);
nor U5157 (N_5157,N_3688,N_3078);
nor U5158 (N_5158,N_3149,N_4137);
xor U5159 (N_5159,N_4014,N_3675);
and U5160 (N_5160,N_4920,N_4199);
nand U5161 (N_5161,N_2828,N_4108);
nand U5162 (N_5162,N_2884,N_3087);
nand U5163 (N_5163,N_4176,N_3020);
and U5164 (N_5164,N_4997,N_4986);
and U5165 (N_5165,N_3178,N_4943);
nor U5166 (N_5166,N_4173,N_4246);
and U5167 (N_5167,N_3644,N_4206);
and U5168 (N_5168,N_4533,N_2827);
nor U5169 (N_5169,N_3800,N_4589);
nor U5170 (N_5170,N_4797,N_4240);
nand U5171 (N_5171,N_4901,N_3983);
and U5172 (N_5172,N_2563,N_3191);
and U5173 (N_5173,N_3162,N_3219);
and U5174 (N_5174,N_3608,N_4160);
and U5175 (N_5175,N_4941,N_2819);
nand U5176 (N_5176,N_2843,N_4386);
and U5177 (N_5177,N_2655,N_4892);
and U5178 (N_5178,N_2728,N_4189);
nand U5179 (N_5179,N_2622,N_2752);
or U5180 (N_5180,N_3958,N_4641);
and U5181 (N_5181,N_4472,N_4213);
or U5182 (N_5182,N_2511,N_4318);
nor U5183 (N_5183,N_3080,N_3887);
and U5184 (N_5184,N_4817,N_3898);
nand U5185 (N_5185,N_2924,N_4711);
or U5186 (N_5186,N_2937,N_4984);
nand U5187 (N_5187,N_3321,N_2623);
nor U5188 (N_5188,N_2570,N_4171);
and U5189 (N_5189,N_4254,N_2525);
or U5190 (N_5190,N_4680,N_4747);
nand U5191 (N_5191,N_4542,N_2803);
or U5192 (N_5192,N_4539,N_3094);
or U5193 (N_5193,N_2934,N_3700);
nand U5194 (N_5194,N_4606,N_3938);
and U5195 (N_5195,N_3233,N_2599);
and U5196 (N_5196,N_2932,N_4498);
nor U5197 (N_5197,N_3332,N_4963);
and U5198 (N_5198,N_3756,N_4384);
nor U5199 (N_5199,N_3702,N_2922);
or U5200 (N_5200,N_3832,N_4563);
nor U5201 (N_5201,N_4967,N_4684);
or U5202 (N_5202,N_3890,N_2796);
or U5203 (N_5203,N_4844,N_3728);
and U5204 (N_5204,N_2761,N_3699);
and U5205 (N_5205,N_3831,N_3151);
or U5206 (N_5206,N_4905,N_4700);
and U5207 (N_5207,N_3862,N_3275);
and U5208 (N_5208,N_4976,N_2671);
or U5209 (N_5209,N_3137,N_4032);
nor U5210 (N_5210,N_4295,N_4034);
and U5211 (N_5211,N_2712,N_2996);
nand U5212 (N_5212,N_4487,N_2870);
xor U5213 (N_5213,N_3866,N_4921);
nand U5214 (N_5214,N_2931,N_4930);
nor U5215 (N_5215,N_4713,N_3239);
or U5216 (N_5216,N_4628,N_3126);
nor U5217 (N_5217,N_4927,N_3032);
nor U5218 (N_5218,N_3742,N_2984);
or U5219 (N_5219,N_3924,N_3491);
and U5220 (N_5220,N_4576,N_3272);
and U5221 (N_5221,N_2957,N_2925);
nand U5222 (N_5222,N_4204,N_2856);
nor U5223 (N_5223,N_4703,N_3549);
nand U5224 (N_5224,N_3281,N_4128);
nor U5225 (N_5225,N_2851,N_3401);
or U5226 (N_5226,N_3150,N_4058);
nand U5227 (N_5227,N_2561,N_3433);
nor U5228 (N_5228,N_3183,N_2916);
and U5229 (N_5229,N_3654,N_4428);
nor U5230 (N_5230,N_2619,N_3475);
or U5231 (N_5231,N_2672,N_2657);
and U5232 (N_5232,N_4673,N_4076);
nor U5233 (N_5233,N_4677,N_3330);
and U5234 (N_5234,N_3110,N_3302);
nand U5235 (N_5235,N_3996,N_3216);
xnor U5236 (N_5236,N_4187,N_4968);
nor U5237 (N_5237,N_4267,N_3505);
or U5238 (N_5238,N_3048,N_4040);
and U5239 (N_5239,N_4352,N_3258);
nor U5240 (N_5240,N_2795,N_4337);
nand U5241 (N_5241,N_3528,N_2545);
and U5242 (N_5242,N_4736,N_4734);
or U5243 (N_5243,N_2814,N_2523);
nand U5244 (N_5244,N_2664,N_3068);
or U5245 (N_5245,N_3293,N_2594);
nor U5246 (N_5246,N_4015,N_2969);
nor U5247 (N_5247,N_2962,N_4234);
or U5248 (N_5248,N_2766,N_4273);
or U5249 (N_5249,N_2705,N_3470);
nor U5250 (N_5250,N_4647,N_4847);
and U5251 (N_5251,N_3678,N_3553);
nand U5252 (N_5252,N_4789,N_2928);
nor U5253 (N_5253,N_3469,N_3860);
or U5254 (N_5254,N_3791,N_3060);
nand U5255 (N_5255,N_2558,N_4398);
nor U5256 (N_5256,N_4536,N_4785);
and U5257 (N_5257,N_4253,N_4250);
xnor U5258 (N_5258,N_3847,N_3434);
and U5259 (N_5259,N_4169,N_4157);
or U5260 (N_5260,N_3835,N_3658);
and U5261 (N_5261,N_3679,N_3561);
nor U5262 (N_5262,N_4334,N_3121);
nor U5263 (N_5263,N_4893,N_4136);
and U5264 (N_5264,N_2580,N_2972);
nand U5265 (N_5265,N_3142,N_4170);
or U5266 (N_5266,N_2739,N_4668);
nor U5267 (N_5267,N_4966,N_2888);
and U5268 (N_5268,N_4834,N_4784);
or U5269 (N_5269,N_3037,N_2529);
nand U5270 (N_5270,N_4538,N_2515);
nand U5271 (N_5271,N_2721,N_3236);
or U5272 (N_5272,N_4911,N_2941);
nor U5273 (N_5273,N_4638,N_3515);
or U5274 (N_5274,N_3441,N_4575);
nand U5275 (N_5275,N_2645,N_4473);
nor U5276 (N_5276,N_3328,N_3462);
and U5277 (N_5277,N_3389,N_2581);
or U5278 (N_5278,N_2681,N_2564);
nand U5279 (N_5279,N_3550,N_4887);
nor U5280 (N_5280,N_4501,N_3498);
or U5281 (N_5281,N_3303,N_4816);
and U5282 (N_5282,N_2789,N_4802);
nand U5283 (N_5283,N_3573,N_3362);
or U5284 (N_5284,N_3575,N_2993);
xnor U5285 (N_5285,N_2596,N_4728);
or U5286 (N_5286,N_2533,N_3271);
nor U5287 (N_5287,N_3845,N_4026);
or U5288 (N_5288,N_3946,N_3125);
nor U5289 (N_5289,N_4069,N_3715);
and U5290 (N_5290,N_3605,N_2544);
and U5291 (N_5291,N_2565,N_4708);
nor U5292 (N_5292,N_2853,N_2811);
nor U5293 (N_5293,N_3815,N_2894);
or U5294 (N_5294,N_4821,N_4678);
nor U5295 (N_5295,N_3801,N_4780);
nor U5296 (N_5296,N_4265,N_4613);
and U5297 (N_5297,N_3339,N_4029);
and U5298 (N_5298,N_2949,N_4056);
and U5299 (N_5299,N_2528,N_4163);
and U5300 (N_5300,N_4612,N_4944);
and U5301 (N_5301,N_2709,N_3349);
nor U5302 (N_5302,N_3400,N_3289);
or U5303 (N_5303,N_4903,N_4094);
nor U5304 (N_5304,N_3894,N_3072);
or U5305 (N_5305,N_2652,N_3576);
nand U5306 (N_5306,N_3316,N_3221);
or U5307 (N_5307,N_2666,N_4074);
xnor U5308 (N_5308,N_2807,N_4438);
nor U5309 (N_5309,N_4975,N_4839);
and U5310 (N_5310,N_3198,N_3753);
nor U5311 (N_5311,N_3770,N_3583);
nor U5312 (N_5312,N_2661,N_3869);
nor U5313 (N_5313,N_4477,N_4325);
nor U5314 (N_5314,N_4154,N_4774);
and U5315 (N_5315,N_4971,N_2555);
and U5316 (N_5316,N_3432,N_3371);
or U5317 (N_5317,N_2889,N_4608);
xnor U5318 (N_5318,N_3283,N_4009);
and U5319 (N_5319,N_4574,N_4629);
nand U5320 (N_5320,N_4635,N_3732);
and U5321 (N_5321,N_4743,N_4441);
or U5322 (N_5322,N_3868,N_3212);
nor U5323 (N_5323,N_2823,N_4982);
nor U5324 (N_5324,N_3383,N_2559);
or U5325 (N_5325,N_3825,N_4965);
nor U5326 (N_5326,N_4357,N_4278);
or U5327 (N_5327,N_3359,N_3952);
nand U5328 (N_5328,N_4460,N_4964);
or U5329 (N_5329,N_4660,N_3234);
nand U5330 (N_5330,N_3993,N_4063);
and U5331 (N_5331,N_4041,N_3899);
and U5332 (N_5332,N_4075,N_3747);
nor U5333 (N_5333,N_3407,N_3836);
and U5334 (N_5334,N_4403,N_3773);
nand U5335 (N_5335,N_4299,N_4153);
nand U5336 (N_5336,N_3481,N_3524);
or U5337 (N_5337,N_4787,N_2861);
nor U5338 (N_5338,N_3457,N_3660);
and U5339 (N_5339,N_4649,N_4271);
nand U5340 (N_5340,N_3409,N_3730);
and U5341 (N_5341,N_4053,N_4355);
and U5342 (N_5342,N_3533,N_4951);
or U5343 (N_5343,N_3012,N_4804);
nor U5344 (N_5344,N_4172,N_2735);
nor U5345 (N_5345,N_4450,N_4885);
nor U5346 (N_5346,N_4509,N_4272);
and U5347 (N_5347,N_3064,N_3992);
or U5348 (N_5348,N_4395,N_2917);
and U5349 (N_5349,N_4599,N_2584);
nor U5350 (N_5350,N_4994,N_4084);
nor U5351 (N_5351,N_3257,N_3799);
or U5352 (N_5352,N_4266,N_3634);
and U5353 (N_5353,N_2751,N_3933);
nor U5354 (N_5354,N_4888,N_3740);
nand U5355 (N_5355,N_3543,N_3300);
nor U5356 (N_5356,N_3519,N_2610);
nand U5357 (N_5357,N_3697,N_4717);
or U5358 (N_5358,N_3696,N_3394);
nor U5359 (N_5359,N_3054,N_2591);
nor U5360 (N_5360,N_2920,N_4497);
or U5361 (N_5361,N_3059,N_4733);
nor U5362 (N_5362,N_2973,N_3393);
and U5363 (N_5363,N_4055,N_3814);
or U5364 (N_5364,N_4739,N_4359);
nor U5365 (N_5365,N_2947,N_3361);
nor U5366 (N_5366,N_3181,N_3222);
or U5367 (N_5367,N_3749,N_3010);
nand U5368 (N_5368,N_3703,N_3278);
nor U5369 (N_5369,N_2913,N_3245);
nor U5370 (N_5370,N_3351,N_3379);
or U5371 (N_5371,N_2818,N_3584);
nand U5372 (N_5372,N_4064,N_3372);
nor U5373 (N_5373,N_2720,N_2734);
nand U5374 (N_5374,N_2694,N_4465);
or U5375 (N_5375,N_4106,N_4183);
nand U5376 (N_5376,N_4766,N_3325);
nor U5377 (N_5377,N_4597,N_2836);
or U5378 (N_5378,N_3138,N_3007);
and U5379 (N_5379,N_4518,N_4195);
or U5380 (N_5380,N_4702,N_3987);
and U5381 (N_5381,N_3218,N_2643);
nand U5382 (N_5382,N_3085,N_3895);
and U5383 (N_5383,N_3725,N_4347);
or U5384 (N_5384,N_2697,N_2765);
or U5385 (N_5385,N_3461,N_3193);
and U5386 (N_5386,N_4731,N_3968);
nand U5387 (N_5387,N_3733,N_3849);
and U5388 (N_5388,N_4645,N_3859);
nor U5389 (N_5389,N_3552,N_4242);
nand U5390 (N_5390,N_4186,N_4174);
and U5391 (N_5391,N_4534,N_4051);
nand U5392 (N_5392,N_2631,N_4914);
and U5393 (N_5393,N_4863,N_4294);
nand U5394 (N_5394,N_2620,N_2503);
or U5395 (N_5395,N_3976,N_2710);
xnor U5396 (N_5396,N_4202,N_3502);
nand U5397 (N_5397,N_2755,N_3521);
nor U5398 (N_5398,N_3492,N_3002);
nor U5399 (N_5399,N_3207,N_4754);
nor U5400 (N_5400,N_2770,N_3243);
or U5401 (N_5401,N_3705,N_3066);
nor U5402 (N_5402,N_4358,N_2571);
and U5403 (N_5403,N_2560,N_2959);
or U5404 (N_5404,N_4184,N_4751);
nor U5405 (N_5405,N_4502,N_2702);
nor U5406 (N_5406,N_2826,N_4822);
nor U5407 (N_5407,N_4177,N_3822);
nor U5408 (N_5408,N_4474,N_2668);
and U5409 (N_5409,N_4626,N_4704);
or U5410 (N_5410,N_4850,N_3579);
and U5411 (N_5411,N_3865,N_3140);
nor U5412 (N_5412,N_4577,N_4671);
nand U5413 (N_5413,N_4531,N_3472);
nor U5414 (N_5414,N_4689,N_4031);
nand U5415 (N_5415,N_3413,N_4017);
or U5416 (N_5416,N_2574,N_3560);
or U5417 (N_5417,N_4223,N_4910);
nor U5418 (N_5418,N_3967,N_4289);
or U5419 (N_5419,N_4527,N_3269);
or U5420 (N_5420,N_2965,N_3312);
nor U5421 (N_5421,N_3919,N_2915);
and U5422 (N_5422,N_3395,N_2714);
or U5423 (N_5423,N_4333,N_4002);
or U5424 (N_5424,N_3019,N_4721);
and U5425 (N_5425,N_4952,N_3252);
nor U5426 (N_5426,N_4624,N_4602);
nand U5427 (N_5427,N_2750,N_3099);
and U5428 (N_5428,N_3594,N_4561);
nand U5429 (N_5429,N_4453,N_4042);
and U5430 (N_5430,N_3721,N_2603);
nand U5431 (N_5431,N_2967,N_4884);
or U5432 (N_5432,N_3681,N_3652);
nor U5433 (N_5433,N_3331,N_3011);
nand U5434 (N_5434,N_3656,N_3663);
nand U5435 (N_5435,N_2670,N_4162);
nor U5436 (N_5436,N_2842,N_4416);
or U5437 (N_5437,N_3834,N_3345);
or U5438 (N_5438,N_2821,N_2893);
and U5439 (N_5439,N_3338,N_4879);
and U5440 (N_5440,N_4862,N_4898);
and U5441 (N_5441,N_4521,N_3179);
or U5442 (N_5442,N_4687,N_3763);
and U5443 (N_5443,N_3440,N_3000);
nor U5444 (N_5444,N_2817,N_4520);
nor U5445 (N_5445,N_4118,N_3506);
nor U5446 (N_5446,N_4415,N_4946);
and U5447 (N_5447,N_3417,N_2582);
nor U5448 (N_5448,N_3449,N_2514);
or U5449 (N_5449,N_3714,N_4131);
and U5450 (N_5450,N_3620,N_2758);
and U5451 (N_5451,N_4500,N_2810);
nand U5452 (N_5452,N_4124,N_2557);
nand U5453 (N_5453,N_4396,N_3436);
nand U5454 (N_5454,N_2798,N_2911);
and U5455 (N_5455,N_4329,N_3488);
nand U5456 (N_5456,N_3296,N_3885);
or U5457 (N_5457,N_3455,N_2832);
and U5458 (N_5458,N_4864,N_3033);
nand U5459 (N_5459,N_4653,N_2679);
nor U5460 (N_5460,N_3691,N_4760);
nor U5461 (N_5461,N_3826,N_2686);
or U5462 (N_5462,N_3001,N_4564);
and U5463 (N_5463,N_3267,N_2538);
nor U5464 (N_5464,N_2611,N_3718);
nor U5465 (N_5465,N_4368,N_3597);
nor U5466 (N_5466,N_3357,N_3105);
or U5467 (N_5467,N_3411,N_4443);
or U5468 (N_5468,N_4099,N_3378);
nand U5469 (N_5469,N_4551,N_3464);
nand U5470 (N_5470,N_2608,N_3384);
or U5471 (N_5471,N_2968,N_4596);
and U5472 (N_5472,N_3035,N_3334);
or U5473 (N_5473,N_4306,N_2699);
nor U5474 (N_5474,N_3381,N_3006);
nand U5475 (N_5475,N_2740,N_3963);
nand U5476 (N_5476,N_2617,N_4248);
or U5477 (N_5477,N_2567,N_2837);
nor U5478 (N_5478,N_3373,N_4039);
and U5479 (N_5479,N_2845,N_4815);
nand U5480 (N_5480,N_4196,N_3599);
nand U5481 (N_5481,N_3544,N_2695);
nor U5482 (N_5482,N_2590,N_4670);
nor U5483 (N_5483,N_2938,N_4339);
nand U5484 (N_5484,N_2776,N_4096);
nand U5485 (N_5485,N_3520,N_4013);
nand U5486 (N_5486,N_3166,N_2820);
nor U5487 (N_5487,N_3202,N_2601);
or U5488 (N_5488,N_3160,N_3451);
xnor U5489 (N_5489,N_4088,N_4953);
xnor U5490 (N_5490,N_4631,N_4033);
or U5491 (N_5491,N_3129,N_4852);
and U5492 (N_5492,N_3672,N_3102);
and U5493 (N_5493,N_3415,N_2543);
nand U5494 (N_5494,N_2852,N_4567);
nor U5495 (N_5495,N_3499,N_4219);
nand U5496 (N_5496,N_3144,N_3726);
nor U5497 (N_5497,N_3255,N_4256);
nor U5498 (N_5498,N_2586,N_2688);
and U5499 (N_5499,N_3387,N_4741);
nand U5500 (N_5500,N_4493,N_2809);
or U5501 (N_5501,N_4654,N_2659);
or U5502 (N_5502,N_2780,N_2833);
nand U5503 (N_5503,N_4105,N_4899);
nand U5504 (N_5504,N_4259,N_4858);
and U5505 (N_5505,N_4637,N_4209);
nor U5506 (N_5506,N_3944,N_4840);
or U5507 (N_5507,N_4705,N_4364);
and U5508 (N_5508,N_4024,N_2691);
nand U5509 (N_5509,N_3227,N_3055);
and U5510 (N_5510,N_4882,N_4021);
nand U5511 (N_5511,N_3176,N_3844);
xnor U5512 (N_5512,N_4729,N_2900);
and U5513 (N_5513,N_3810,N_3548);
or U5514 (N_5514,N_3902,N_2901);
nor U5515 (N_5515,N_3984,N_4197);
and U5516 (N_5516,N_2849,N_4912);
or U5517 (N_5517,N_4354,N_3244);
and U5518 (N_5518,N_4314,N_3329);
nand U5519 (N_5519,N_3682,N_4119);
nand U5520 (N_5520,N_4825,N_3045);
nand U5521 (N_5521,N_3635,N_2904);
nand U5522 (N_5522,N_4201,N_3657);
or U5523 (N_5523,N_3232,N_2551);
nand U5524 (N_5524,N_2879,N_4270);
nand U5525 (N_5525,N_2899,N_4349);
nor U5526 (N_5526,N_4807,N_3685);
nor U5527 (N_5527,N_2975,N_3235);
and U5528 (N_5528,N_3662,N_4439);
nand U5529 (N_5529,N_2642,N_2815);
nand U5530 (N_5530,N_3525,N_3341);
or U5531 (N_5531,N_3568,N_3397);
or U5532 (N_5532,N_4883,N_4495);
and U5533 (N_5533,N_4735,N_3256);
or U5534 (N_5534,N_3042,N_2531);
nand U5535 (N_5535,N_3893,N_3768);
and U5536 (N_5536,N_4208,N_3427);
or U5537 (N_5537,N_4408,N_3173);
and U5538 (N_5538,N_2746,N_3342);
nand U5539 (N_5539,N_4499,N_2793);
nand U5540 (N_5540,N_4685,N_2978);
and U5541 (N_5541,N_3623,N_3442);
nand U5542 (N_5542,N_2921,N_3881);
nor U5543 (N_5543,N_4085,N_2804);
or U5544 (N_5544,N_4681,N_4742);
or U5545 (N_5545,N_3614,N_2535);
nor U5546 (N_5546,N_2625,N_3124);
and U5547 (N_5547,N_3823,N_4107);
or U5548 (N_5548,N_4066,N_2602);
and U5549 (N_5549,N_4005,N_4665);
or U5550 (N_5550,N_3643,N_3053);
nor U5551 (N_5551,N_3886,N_3391);
and U5552 (N_5552,N_4091,N_4405);
or U5553 (N_5553,N_3399,N_4988);
and U5554 (N_5554,N_2998,N_2935);
nand U5555 (N_5555,N_3949,N_4297);
nand U5556 (N_5556,N_4980,N_4591);
nand U5557 (N_5557,N_4651,N_2943);
nor U5558 (N_5558,N_2813,N_4989);
or U5559 (N_5559,N_4854,N_3545);
nand U5560 (N_5560,N_4469,N_4090);
and U5561 (N_5561,N_4528,N_3953);
and U5562 (N_5562,N_4227,N_4928);
or U5563 (N_5563,N_3858,N_4312);
or U5564 (N_5564,N_4132,N_2522);
or U5565 (N_5565,N_3158,N_2577);
and U5566 (N_5566,N_3490,N_3588);
or U5567 (N_5567,N_3313,N_3735);
or U5568 (N_5568,N_3213,N_2977);
or U5569 (N_5569,N_3238,N_3587);
and U5570 (N_5570,N_3074,N_3631);
or U5571 (N_5571,N_3913,N_4973);
nand U5572 (N_5572,N_3677,N_2785);
nand U5573 (N_5573,N_4841,N_4356);
nand U5574 (N_5574,N_3217,N_2919);
and U5575 (N_5575,N_3804,N_3808);
nor U5576 (N_5576,N_3497,N_3081);
and U5577 (N_5577,N_4215,N_3592);
and U5578 (N_5578,N_3931,N_4483);
nand U5579 (N_5579,N_3199,N_4819);
nor U5580 (N_5580,N_3798,N_4182);
nor U5581 (N_5581,N_4471,N_2887);
nand U5582 (N_5582,N_3909,N_3724);
and U5583 (N_5583,N_3722,N_3406);
and U5584 (N_5584,N_3673,N_3168);
and U5585 (N_5585,N_4225,N_4627);
or U5586 (N_5586,N_2976,N_3315);
nor U5587 (N_5587,N_3790,N_4583);
or U5588 (N_5588,N_4701,N_2876);
and U5589 (N_5589,N_4621,N_4006);
nand U5590 (N_5590,N_4578,N_3789);
or U5591 (N_5591,N_4956,N_4748);
or U5592 (N_5592,N_3242,N_2742);
xor U5593 (N_5593,N_3069,N_2954);
and U5594 (N_5594,N_4548,N_2700);
nor U5595 (N_5595,N_3708,N_3727);
and U5596 (N_5596,N_3674,N_4857);
and U5597 (N_5597,N_3551,N_4793);
nand U5598 (N_5598,N_2595,N_4950);
nand U5599 (N_5599,N_4646,N_4752);
nor U5600 (N_5600,N_4249,N_3995);
nor U5601 (N_5601,N_3240,N_4363);
or U5602 (N_5602,N_3517,N_4399);
and U5603 (N_5603,N_2706,N_4038);
or U5604 (N_5604,N_2918,N_4672);
or U5605 (N_5605,N_3333,N_3308);
and U5606 (N_5606,N_3842,N_3051);
and U5607 (N_5607,N_4837,N_2877);
and U5608 (N_5608,N_4869,N_2791);
nand U5609 (N_5609,N_4061,N_4934);
and U5610 (N_5610,N_3230,N_2539);
and U5611 (N_5611,N_4342,N_3065);
nand U5612 (N_5612,N_4803,N_3377);
nand U5613 (N_5613,N_2569,N_4425);
nor U5614 (N_5614,N_2805,N_4769);
or U5615 (N_5615,N_4103,N_3156);
nor U5616 (N_5616,N_4012,N_2546);
and U5617 (N_5617,N_4008,N_3248);
or U5618 (N_5618,N_3277,N_3082);
or U5619 (N_5619,N_3422,N_4394);
and U5620 (N_5620,N_2980,N_3437);
nand U5621 (N_5621,N_4764,N_3593);
or U5622 (N_5622,N_2907,N_3005);
nor U5623 (N_5623,N_2606,N_2794);
and U5624 (N_5624,N_2933,N_3290);
nor U5625 (N_5625,N_4810,N_3581);
nor U5626 (N_5626,N_3974,N_3878);
nand U5627 (N_5627,N_3966,N_4594);
nor U5628 (N_5628,N_2890,N_3916);
nor U5629 (N_5629,N_3431,N_3874);
or U5630 (N_5630,N_3172,N_4916);
or U5631 (N_5631,N_4799,N_3091);
nand U5632 (N_5632,N_4097,N_4146);
or U5633 (N_5633,N_3210,N_4759);
and U5634 (N_5634,N_4604,N_2730);
or U5635 (N_5635,N_4507,N_2777);
nand U5636 (N_5636,N_3049,N_4666);
nor U5637 (N_5637,N_3265,N_3205);
nand U5638 (N_5638,N_3910,N_3382);
nand U5639 (N_5639,N_2747,N_3326);
nand U5640 (N_5640,N_3153,N_4464);
and U5641 (N_5641,N_3964,N_3320);
or U5642 (N_5642,N_4141,N_4149);
nand U5643 (N_5643,N_2982,N_4444);
xnor U5644 (N_5644,N_4902,N_4046);
or U5645 (N_5645,N_3294,N_3096);
nand U5646 (N_5646,N_2638,N_3116);
nand U5647 (N_5647,N_4379,N_4470);
or U5648 (N_5648,N_4252,N_3390);
and U5649 (N_5649,N_3136,N_2862);
nor U5650 (N_5650,N_3448,N_4393);
nor U5651 (N_5651,N_3961,N_4725);
and U5652 (N_5652,N_4795,N_4722);
and U5653 (N_5653,N_2527,N_4652);
nor U5654 (N_5654,N_4719,N_2698);
or U5655 (N_5655,N_2858,N_3420);
and U5656 (N_5656,N_2629,N_2745);
and U5657 (N_5657,N_3071,N_2613);
nand U5658 (N_5658,N_4838,N_4264);
or U5659 (N_5659,N_4650,N_3709);
and U5660 (N_5660,N_2537,N_3465);
and U5661 (N_5661,N_3973,N_2504);
nor U5662 (N_5662,N_2753,N_3562);
nand U5663 (N_5663,N_3911,N_3571);
nand U5664 (N_5664,N_2825,N_4782);
nand U5665 (N_5665,N_2940,N_4552);
and U5666 (N_5666,N_3023,N_3322);
and U5667 (N_5667,N_3704,N_4410);
nand U5668 (N_5668,N_3208,N_4853);
nor U5669 (N_5669,N_3196,N_4848);
nor U5670 (N_5670,N_4095,N_4139);
and U5671 (N_5671,N_4925,N_4011);
nand U5672 (N_5672,N_3556,N_3806);
and U5673 (N_5673,N_4544,N_4480);
and U5674 (N_5674,N_3058,N_2637);
nand U5675 (N_5675,N_3220,N_4143);
and U5676 (N_5676,N_3224,N_3358);
nor U5677 (N_5677,N_3595,N_4369);
nor U5678 (N_5678,N_2532,N_2762);
or U5679 (N_5679,N_4897,N_3459);
nand U5680 (N_5680,N_3538,N_2756);
nand U5681 (N_5681,N_3680,N_4909);
or U5682 (N_5682,N_2607,N_3606);
or U5683 (N_5683,N_4442,N_4116);
and U5684 (N_5684,N_4757,N_4211);
nand U5685 (N_5685,N_3185,N_2829);
or U5686 (N_5686,N_4190,N_4104);
nor U5687 (N_5687,N_3421,N_3907);
nor U5688 (N_5688,N_3636,N_4224);
nand U5689 (N_5689,N_3089,N_4656);
and U5690 (N_5690,N_3092,N_2738);
and U5691 (N_5691,N_2675,N_4262);
nor U5692 (N_5692,N_3356,N_4089);
nand U5693 (N_5693,N_3375,N_3120);
or U5694 (N_5694,N_3776,N_2806);
nor U5695 (N_5695,N_4346,N_3788);
nor U5696 (N_5696,N_4231,N_3017);
nand U5697 (N_5697,N_4933,N_3811);
nand U5698 (N_5698,N_3978,N_4123);
nand U5699 (N_5699,N_4152,N_2910);
or U5700 (N_5700,N_4998,N_3641);
nand U5701 (N_5701,N_4235,N_4244);
and U5702 (N_5702,N_3783,N_4377);
nand U5703 (N_5703,N_3578,N_3603);
nand U5704 (N_5704,N_2860,N_3077);
nand U5705 (N_5705,N_2981,N_4657);
nor U5706 (N_5706,N_2906,N_4315);
or U5707 (N_5707,N_4054,N_4018);
nor U5708 (N_5708,N_4727,N_3405);
nand U5709 (N_5709,N_3539,N_4800);
nor U5710 (N_5710,N_4381,N_3661);
nand U5711 (N_5711,N_3292,N_3600);
nor U5712 (N_5712,N_3353,N_4640);
or U5713 (N_5713,N_3534,N_4504);
or U5714 (N_5714,N_4999,N_3438);
or U5715 (N_5715,N_2630,N_3474);
nand U5716 (N_5716,N_3851,N_4991);
and U5717 (N_5717,N_2600,N_4724);
or U5718 (N_5718,N_3853,N_2649);
nor U5719 (N_5719,N_4462,N_4370);
or U5720 (N_5720,N_4592,N_4726);
nor U5721 (N_5721,N_3601,N_4826);
or U5722 (N_5722,N_4891,N_2778);
or U5723 (N_5723,N_3194,N_4609);
nand U5724 (N_5724,N_3873,N_2784);
nand U5725 (N_5725,N_3738,N_2542);
and U5726 (N_5726,N_4387,N_3824);
or U5727 (N_5727,N_3446,N_4035);
nor U5728 (N_5728,N_4161,N_4047);
nor U5729 (N_5729,N_4755,N_3555);
and U5730 (N_5730,N_2875,N_4148);
and U5731 (N_5731,N_4113,N_2703);
nor U5732 (N_5732,N_3692,N_2572);
or U5733 (N_5733,N_4908,N_2839);
or U5734 (N_5734,N_4808,N_4435);
or U5735 (N_5735,N_4562,N_4706);
nor U5736 (N_5736,N_2995,N_2724);
nand U5737 (N_5737,N_3344,N_4236);
nor U5738 (N_5738,N_2614,N_2729);
or U5739 (N_5739,N_3301,N_3921);
nand U5740 (N_5740,N_3896,N_4214);
or U5741 (N_5741,N_3569,N_2749);
nor U5742 (N_5742,N_4310,N_3965);
and U5743 (N_5743,N_4404,N_4737);
nor U5744 (N_5744,N_4375,N_3912);
or U5745 (N_5745,N_3314,N_3781);
or U5746 (N_5746,N_4636,N_2963);
or U5747 (N_5747,N_4221,N_4634);
or U5748 (N_5748,N_4412,N_4083);
nor U5749 (N_5749,N_4308,N_4601);
nand U5750 (N_5750,N_4378,N_2711);
nor U5751 (N_5751,N_3024,N_4229);
and U5752 (N_5752,N_3695,N_2736);
nand U5753 (N_5753,N_2974,N_4526);
nor U5754 (N_5754,N_2983,N_4767);
nor U5755 (N_5755,N_4109,N_2549);
or U5756 (N_5756,N_3778,N_3192);
nand U5757 (N_5757,N_3062,N_4642);
nor U5758 (N_5758,N_4805,N_3701);
or U5759 (N_5759,N_4422,N_3570);
or U5760 (N_5760,N_4874,N_3211);
or U5761 (N_5761,N_3430,N_3485);
nor U5762 (N_5762,N_3473,N_3951);
or U5763 (N_5763,N_3145,N_3977);
nor U5764 (N_5764,N_4753,N_2953);
nor U5765 (N_5765,N_3945,N_4343);
nand U5766 (N_5766,N_4121,N_3200);
or U5767 (N_5767,N_3241,N_2838);
or U5768 (N_5768,N_3251,N_2863);
nand U5769 (N_5769,N_3513,N_3425);
nand U5770 (N_5770,N_4112,N_4712);
and U5771 (N_5771,N_2944,N_3424);
nand U5772 (N_5772,N_3182,N_3676);
and U5773 (N_5773,N_3003,N_4765);
nor U5774 (N_5774,N_4761,N_3134);
nor U5775 (N_5775,N_4077,N_3368);
or U5776 (N_5776,N_3540,N_4549);
nand U5777 (N_5777,N_4309,N_3249);
nor U5778 (N_5778,N_2597,N_3729);
nor U5779 (N_5779,N_4079,N_4618);
nand U5780 (N_5780,N_4648,N_4098);
nand U5781 (N_5781,N_2871,N_3888);
or U5782 (N_5782,N_3745,N_4746);
or U5783 (N_5783,N_3487,N_3877);
or U5784 (N_5784,N_3990,N_2966);
and U5785 (N_5785,N_4050,N_3337);
and U5786 (N_5786,N_4587,N_3365);
nor U5787 (N_5787,N_2992,N_3288);
nor U5788 (N_5788,N_4830,N_3640);
nor U5789 (N_5789,N_2540,N_3454);
and U5790 (N_5790,N_3501,N_2656);
and U5791 (N_5791,N_3484,N_4317);
nor U5792 (N_5792,N_4593,N_4894);
or U5793 (N_5793,N_3186,N_3712);
nor U5794 (N_5794,N_2731,N_2693);
and U5795 (N_5795,N_4268,N_3030);
nor U5796 (N_5796,N_4750,N_4643);
and U5797 (N_5797,N_3975,N_2874);
and U5798 (N_5798,N_4992,N_3914);
nor U5799 (N_5799,N_4191,N_4915);
or U5800 (N_5800,N_4740,N_2760);
or U5801 (N_5801,N_2513,N_4134);
nand U5802 (N_5802,N_3757,N_3444);
nand U5803 (N_5803,N_3061,N_3716);
nand U5804 (N_5804,N_2859,N_3901);
nand U5805 (N_5805,N_4300,N_3508);
nand U5806 (N_5806,N_4220,N_3115);
and U5807 (N_5807,N_3854,N_3629);
nand U5808 (N_5808,N_4285,N_4100);
or U5809 (N_5809,N_4175,N_4938);
or U5810 (N_5810,N_3197,N_3633);
nor U5811 (N_5811,N_2556,N_4421);
nor U5812 (N_5812,N_2822,N_4376);
nand U5813 (N_5813,N_4479,N_3848);
nand U5814 (N_5814,N_2589,N_4449);
or U5815 (N_5815,N_4316,N_2660);
nor U5816 (N_5816,N_3229,N_3025);
or U5817 (N_5817,N_4516,N_3782);
nor U5818 (N_5818,N_3348,N_3582);
nand U5819 (N_5819,N_3875,N_4659);
and U5820 (N_5820,N_4237,N_4566);
nand U5821 (N_5821,N_3335,N_3095);
or U5822 (N_5822,N_4207,N_4768);
or U5823 (N_5823,N_4114,N_2898);
and U5824 (N_5824,N_2526,N_4232);
nand U5825 (N_5825,N_3073,N_4335);
or U5826 (N_5826,N_3428,N_3664);
nor U5827 (N_5827,N_3041,N_2754);
nor U5828 (N_5828,N_2598,N_3360);
or U5829 (N_5829,N_4843,N_3855);
nor U5830 (N_5830,N_4801,N_3467);
or U5831 (N_5831,N_3404,N_4525);
or U5832 (N_5832,N_4291,N_2797);
and U5833 (N_5833,N_4494,N_3867);
nand U5834 (N_5834,N_3070,N_3056);
or U5835 (N_5835,N_3106,N_4243);
and U5836 (N_5836,N_2518,N_2627);
and U5837 (N_5837,N_3925,N_3793);
nand U5838 (N_5838,N_3897,N_4983);
and U5839 (N_5839,N_3471,N_2989);
nand U5840 (N_5840,N_3693,N_4560);
or U5841 (N_5841,N_4679,N_4284);
or U5842 (N_5842,N_3304,N_4682);
nor U5843 (N_5843,N_3263,N_4392);
or U5844 (N_5844,N_4693,N_2684);
or U5845 (N_5845,N_2986,N_4707);
or U5846 (N_5846,N_4792,N_3927);
and U5847 (N_5847,N_3163,N_3370);
nand U5848 (N_5848,N_3838,N_4277);
or U5849 (N_5849,N_3340,N_4845);
and U5850 (N_5850,N_3731,N_3554);
or U5851 (N_5851,N_2674,N_4274);
and U5852 (N_5852,N_2772,N_3780);
or U5853 (N_5853,N_2816,N_2650);
xor U5854 (N_5854,N_2704,N_4762);
or U5855 (N_5855,N_3805,N_3253);
nand U5856 (N_5856,N_2790,N_3619);
and U5857 (N_5857,N_2583,N_3223);
nor U5858 (N_5858,N_4102,N_3585);
xnor U5859 (N_5859,N_4569,N_3027);
xnor U5860 (N_5860,N_2676,N_3478);
or U5861 (N_5861,N_3468,N_2719);
nand U5862 (N_5862,N_3999,N_3647);
nor U5863 (N_5863,N_4524,N_4674);
nor U5864 (N_5864,N_3410,N_4699);
and U5865 (N_5865,N_3755,N_4067);
and U5866 (N_5866,N_3034,N_3098);
or U5867 (N_5867,N_3347,N_3127);
or U5868 (N_5868,N_3818,N_2912);
and U5869 (N_5869,N_4217,N_4491);
or U5870 (N_5870,N_4889,N_4241);
or U5871 (N_5871,N_3785,N_2716);
or U5872 (N_5872,N_4010,N_4181);
nor U5873 (N_5873,N_3580,N_4431);
nand U5874 (N_5874,N_3100,N_4686);
nand U5875 (N_5875,N_3247,N_4697);
or U5876 (N_5876,N_3103,N_3479);
nand U5877 (N_5877,N_2994,N_3355);
or U5878 (N_5878,N_3171,N_3612);
and U5879 (N_5879,N_3090,N_3526);
nand U5880 (N_5880,N_2500,N_4283);
nor U5881 (N_5881,N_3429,N_4280);
nand U5882 (N_5882,N_4049,N_3760);
and U5883 (N_5883,N_2883,N_3744);
or U5884 (N_5884,N_3932,N_4959);
and U5885 (N_5885,N_4303,N_4078);
nand U5886 (N_5886,N_3214,N_4457);
or U5887 (N_5887,N_4541,N_2759);
and U5888 (N_5888,N_3503,N_4831);
nand U5889 (N_5889,N_3668,N_2866);
nand U5890 (N_5890,N_3969,N_4919);
and U5891 (N_5891,N_4866,N_3988);
nand U5892 (N_5892,N_2579,N_4382);
nor U5893 (N_5893,N_4043,N_4922);
or U5894 (N_5894,N_2678,N_2929);
nand U5895 (N_5895,N_3418,N_3929);
and U5896 (N_5896,N_4846,N_2717);
nor U5897 (N_5897,N_2854,N_4305);
nor U5898 (N_5898,N_4588,N_2960);
nand U5899 (N_5899,N_4179,N_2715);
nand U5900 (N_5900,N_3204,N_2767);
nor U5901 (N_5901,N_4995,N_4935);
and U5902 (N_5902,N_3559,N_3187);
xnor U5903 (N_5903,N_4947,N_4949);
xnor U5904 (N_5904,N_3477,N_3323);
or U5905 (N_5905,N_4287,N_4448);
nor U5906 (N_5906,N_4007,N_3135);
and U5907 (N_5907,N_4331,N_3480);
nand U5908 (N_5908,N_4630,N_2885);
and U5909 (N_5909,N_4151,N_2632);
and U5910 (N_5910,N_3306,N_3746);
and U5911 (N_5911,N_3456,N_4579);
and U5912 (N_5912,N_3117,N_4486);
nor U5913 (N_5913,N_4585,N_2909);
or U5914 (N_5914,N_4615,N_3044);
or U5915 (N_5915,N_3146,N_4036);
nor U5916 (N_5916,N_4878,N_4420);
nand U5917 (N_5917,N_2516,N_4446);
and U5918 (N_5918,N_4865,N_3937);
nor U5919 (N_5919,N_3870,N_3748);
and U5920 (N_5920,N_4133,N_4929);
and U5921 (N_5921,N_4048,N_2677);
or U5922 (N_5922,N_4515,N_4896);
nand U5923 (N_5923,N_3535,N_4508);
nor U5924 (N_5924,N_4868,N_3839);
or U5925 (N_5925,N_3075,N_3947);
nor U5926 (N_5926,N_4876,N_3922);
and U5927 (N_5927,N_4923,N_3307);
or U5928 (N_5928,N_3802,N_4535);
nor U5929 (N_5929,N_2743,N_4978);
or U5930 (N_5930,N_4093,N_3774);
nand U5931 (N_5931,N_4872,N_4496);
or U5932 (N_5932,N_2653,N_4419);
nand U5933 (N_5933,N_4060,N_3021);
nor U5934 (N_5934,N_4781,N_4447);
nand U5935 (N_5935,N_4142,N_2774);
and U5936 (N_5936,N_4913,N_4022);
or U5937 (N_5937,N_3787,N_3392);
or U5938 (N_5938,N_2781,N_3482);
nand U5939 (N_5939,N_4720,N_4532);
and U5940 (N_5940,N_3625,N_4019);
and U5941 (N_5941,N_3310,N_4313);
nor U5942 (N_5942,N_4835,N_3346);
or U5943 (N_5943,N_2985,N_2763);
or U5944 (N_5944,N_3453,N_3250);
and U5945 (N_5945,N_4924,N_3816);
or U5946 (N_5946,N_2708,N_3014);
nand U5947 (N_5947,N_3226,N_4813);
nand U5948 (N_5948,N_3206,N_3108);
nor U5949 (N_5949,N_4178,N_3646);
nor U5950 (N_5950,N_3710,N_4979);
and U5951 (N_5951,N_3743,N_4696);
nand U5952 (N_5952,N_4540,N_3317);
or U5953 (N_5953,N_3630,N_4168);
or U5954 (N_5954,N_3403,N_4957);
and U5955 (N_5955,N_3797,N_4818);
nor U5956 (N_5956,N_3228,N_3764);
nor U5957 (N_5957,N_4467,N_2718);
nand U5958 (N_5958,N_2667,N_3486);
xnor U5959 (N_5959,N_4522,N_3741);
nor U5960 (N_5960,N_4756,N_3284);
or U5961 (N_5961,N_2713,N_4981);
or U5962 (N_5962,N_3621,N_3903);
and U5963 (N_5963,N_4001,N_3626);
nor U5964 (N_5964,N_2788,N_3563);
and U5965 (N_5965,N_3591,N_3819);
nor U5966 (N_5966,N_4292,N_3567);
and U5967 (N_5967,N_3713,N_2812);
nand U5968 (N_5968,N_3189,N_4080);
nor U5969 (N_5969,N_3079,N_3209);
and U5970 (N_5970,N_4537,N_2521);
nand U5971 (N_5971,N_2646,N_3439);
nand U5972 (N_5972,N_4311,N_2530);
nand U5973 (N_5973,N_3928,N_4937);
and U5974 (N_5974,N_3557,N_4715);
or U5975 (N_5975,N_3507,N_4758);
and U5976 (N_5976,N_3016,N_4870);
and U5977 (N_5977,N_3161,N_4619);
or U5978 (N_5978,N_4255,N_3013);
or U5979 (N_5979,N_3934,N_4293);
nor U5980 (N_5980,N_3336,N_4558);
or U5981 (N_5981,N_3861,N_4198);
nor U5982 (N_5982,N_3628,N_2566);
or U5983 (N_5983,N_3511,N_3452);
or U5984 (N_5984,N_3254,N_4931);
or U5985 (N_5985,N_3642,N_3130);
or U5986 (N_5986,N_3101,N_2651);
and U5987 (N_5987,N_3723,N_2903);
nand U5988 (N_5988,N_3841,N_4463);
nand U5989 (N_5989,N_3624,N_4833);
and U5990 (N_5990,N_3939,N_2669);
or U5991 (N_5991,N_4320,N_4245);
nor U5992 (N_5992,N_2869,N_3537);
nor U5993 (N_5993,N_4867,N_3460);
nand U5994 (N_5994,N_4907,N_3767);
or U5995 (N_5995,N_3666,N_4145);
or U5996 (N_5996,N_4771,N_3119);
and U5997 (N_5997,N_4859,N_4468);
nor U5998 (N_5998,N_3979,N_3039);
or U5999 (N_5999,N_4586,N_3807);
and U6000 (N_6000,N_3616,N_2636);
nand U6001 (N_6001,N_3067,N_4530);
nor U6002 (N_6002,N_4140,N_3107);
nand U6003 (N_6003,N_2902,N_3036);
or U6004 (N_6004,N_3821,N_3157);
and U6005 (N_6005,N_3155,N_4144);
nor U6006 (N_6006,N_4045,N_2541);
nor U6007 (N_6007,N_4582,N_4138);
or U6008 (N_6008,N_2644,N_4714);
and U6009 (N_6009,N_3295,N_2723);
nor U6010 (N_6010,N_2844,N_3786);
nor U6011 (N_6011,N_4890,N_2506);
nand U6012 (N_6012,N_4000,N_3651);
or U6013 (N_6013,N_4275,N_4610);
nand U6014 (N_6014,N_3532,N_3915);
and U6015 (N_6015,N_2782,N_2647);
nor U6016 (N_6016,N_2685,N_4732);
nor U6017 (N_6017,N_4770,N_3784);
nand U6018 (N_6018,N_2633,N_3917);
nor U6019 (N_6019,N_2648,N_4547);
nor U6020 (N_6020,N_3523,N_3775);
and U6021 (N_6021,N_3287,N_4565);
and U6022 (N_6022,N_3516,N_3803);
and U6023 (N_6023,N_3813,N_4406);
nor U6024 (N_6024,N_4709,N_4461);
or U6025 (N_6025,N_3792,N_3496);
or U6026 (N_6026,N_3930,N_4571);
or U6027 (N_6027,N_2520,N_4127);
nand U6028 (N_6028,N_2886,N_4985);
nand U6029 (N_6029,N_4484,N_2878);
nand U6030 (N_6030,N_4557,N_3639);
nor U6031 (N_6031,N_3445,N_3905);
and U6032 (N_6032,N_2665,N_4745);
or U6033 (N_6033,N_2801,N_2536);
nor U6034 (N_6034,N_2950,N_4823);
and U6035 (N_6035,N_2626,N_4970);
or U6036 (N_6036,N_4307,N_2880);
nor U6037 (N_6037,N_4580,N_3026);
nand U6038 (N_6038,N_3607,N_4413);
nor U6039 (N_6039,N_3500,N_3950);
nor U6040 (N_6040,N_3113,N_3852);
and U6041 (N_6041,N_3531,N_3970);
nor U6042 (N_6042,N_4718,N_3165);
and U6043 (N_6043,N_2882,N_3772);
nand U6044 (N_6044,N_4829,N_2864);
nor U6045 (N_6045,N_4147,N_4433);
nor U6046 (N_6046,N_4125,N_2501);
and U6047 (N_6047,N_4842,N_4820);
nand U6048 (N_6048,N_2547,N_4791);
and U6049 (N_6049,N_4620,N_2905);
or U6050 (N_6050,N_2939,N_3589);
or U6051 (N_6051,N_2956,N_4476);
nand U6052 (N_6052,N_3843,N_4623);
or U6053 (N_6053,N_4418,N_4110);
and U6054 (N_6054,N_3225,N_3203);
and U6055 (N_6055,N_2970,N_2508);
and U6056 (N_6056,N_3942,N_2658);
nor U6057 (N_6057,N_3765,N_2800);
nor U6058 (N_6058,N_2680,N_3985);
nor U6059 (N_6059,N_2512,N_2592);
or U6060 (N_6060,N_3367,N_4794);
or U6061 (N_6061,N_3615,N_4856);
and U6062 (N_6062,N_4798,N_4773);
or U6063 (N_6063,N_4451,N_4321);
nand U6064 (N_6064,N_3632,N_3398);
or U6065 (N_6065,N_4662,N_3957);
nand U6066 (N_6066,N_4644,N_3618);
nand U6067 (N_6067,N_4326,N_4738);
and U6068 (N_6068,N_2999,N_4716);
and U6069 (N_6069,N_4632,N_3143);
nor U6070 (N_6070,N_4581,N_4877);
nor U6071 (N_6071,N_3655,N_4044);
nor U6072 (N_6072,N_3476,N_3043);
or U6073 (N_6073,N_3955,N_3366);
nand U6074 (N_6074,N_3694,N_3872);
nand U6075 (N_6075,N_3093,N_4230);
nand U6076 (N_6076,N_4543,N_4570);
nand U6077 (N_6077,N_2692,N_3435);
and U6078 (N_6078,N_4193,N_4554);
nand U6079 (N_6079,N_3837,N_4417);
or U6080 (N_6080,N_2634,N_4886);
or U6081 (N_6081,N_2554,N_4188);
nor U6082 (N_6082,N_4904,N_4401);
nor U6083 (N_6083,N_2524,N_3771);
nand U6084 (N_6084,N_4429,N_3879);
or U6085 (N_6085,N_4452,N_2726);
nand U6086 (N_6086,N_3817,N_2733);
or U6087 (N_6087,N_4744,N_4932);
or U6088 (N_6088,N_3380,N_4590);
and U6089 (N_6089,N_3994,N_4459);
and U6090 (N_6090,N_4723,N_4257);
or U6091 (N_6091,N_4203,N_3118);
or U6092 (N_6092,N_3131,N_2979);
and U6093 (N_6093,N_2802,N_4233);
nand U6094 (N_6094,N_4301,N_4411);
nand U6095 (N_6095,N_4860,N_4948);
or U6096 (N_6096,N_3104,N_2578);
nand U6097 (N_6097,N_3750,N_3820);
nand U6098 (N_6098,N_2779,N_4407);
and U6099 (N_6099,N_3940,N_4282);
or U6100 (N_6100,N_4873,N_3530);
or U6101 (N_6101,N_4490,N_4622);
and U6102 (N_6102,N_3864,N_4281);
nand U6103 (N_6103,N_3923,N_2926);
and U6104 (N_6104,N_4806,N_3684);
and U6105 (N_6105,N_4290,N_2990);
and U6106 (N_6106,N_4228,N_4811);
nand U6107 (N_6107,N_2892,N_4117);
and U6108 (N_6108,N_4430,N_3707);
and U6109 (N_6109,N_3769,N_4511);
or U6110 (N_6110,N_3164,N_4304);
nand U6111 (N_6111,N_2891,N_2748);
nand U6112 (N_6112,N_3891,N_2991);
and U6113 (N_6113,N_3918,N_4323);
nor U6114 (N_6114,N_4122,N_4101);
and U6115 (N_6115,N_3327,N_3386);
and U6116 (N_6116,N_4917,N_2701);
or U6117 (N_6117,N_4616,N_4071);
or U6118 (N_6118,N_4676,N_3829);
nand U6119 (N_6119,N_3686,N_2744);
nor U6120 (N_6120,N_4832,N_4052);
nor U6121 (N_6121,N_3354,N_3363);
and U6122 (N_6122,N_4286,N_3665);
nand U6123 (N_6123,N_4710,N_3009);
and U6124 (N_6124,N_2769,N_3751);
and U6125 (N_6125,N_4218,N_2737);
nand U6126 (N_6126,N_4611,N_4990);
nand U6127 (N_6127,N_4226,N_2588);
and U6128 (N_6128,N_3112,N_3369);
and U6129 (N_6129,N_4458,N_4288);
nor U6130 (N_6130,N_4881,N_3638);
and U6131 (N_6131,N_3900,N_4695);
or U6132 (N_6132,N_3754,N_2881);
or U6133 (N_6133,N_4488,N_4129);
nor U6134 (N_6134,N_2696,N_2662);
or U6135 (N_6135,N_4260,N_3986);
or U6136 (N_6136,N_4814,N_3876);
and U6137 (N_6137,N_4639,N_3706);
or U6138 (N_6138,N_3463,N_3086);
and U6139 (N_6139,N_4828,N_4926);
or U6140 (N_6140,N_3698,N_3175);
or U6141 (N_6141,N_2618,N_3159);
nor U6142 (N_6142,N_2946,N_3264);
or U6143 (N_6143,N_3794,N_4595);
and U6144 (N_6144,N_3319,N_3122);
nor U6145 (N_6145,N_4082,N_3959);
and U6146 (N_6146,N_3613,N_4298);
and U6147 (N_6147,N_4023,N_4568);
and U6148 (N_6148,N_4456,N_4332);
nand U6149 (N_6149,N_3504,N_3962);
nand U6150 (N_6150,N_4296,N_4130);
nand U6151 (N_6151,N_4388,N_4030);
or U6152 (N_6152,N_3088,N_3018);
and U6153 (N_6153,N_4514,N_3518);
and U6154 (N_6154,N_4185,N_3926);
and U6155 (N_6155,N_3734,N_3954);
and U6156 (N_6156,N_3114,N_2616);
and U6157 (N_6157,N_3812,N_4159);
nor U6158 (N_6158,N_4955,N_4426);
and U6159 (N_6159,N_3123,N_2792);
nor U6160 (N_6160,N_2783,N_2587);
nand U6161 (N_6161,N_3402,N_2865);
or U6162 (N_6162,N_3412,N_3259);
or U6163 (N_6163,N_4614,N_2534);
nor U6164 (N_6164,N_4895,N_2958);
or U6165 (N_6165,N_4158,N_3352);
and U6166 (N_6166,N_3736,N_4556);
or U6167 (N_6167,N_4996,N_3139);
nand U6168 (N_6168,N_4775,N_3376);
nor U6169 (N_6169,N_4276,N_3856);
and U6170 (N_6170,N_4279,N_3880);
nor U6171 (N_6171,N_3527,N_4918);
nand U6172 (N_6172,N_3262,N_3299);
or U6173 (N_6173,N_4409,N_4414);
and U6174 (N_6174,N_3004,N_3408);
nand U6175 (N_6175,N_4824,N_4503);
and U6176 (N_6176,N_3833,N_4698);
and U6177 (N_6177,N_2841,N_2690);
nand U6178 (N_6178,N_4360,N_4790);
nor U6179 (N_6179,N_4327,N_3097);
nand U6180 (N_6180,N_4210,N_4942);
and U6181 (N_6181,N_4427,N_4155);
xnor U6182 (N_6182,N_4423,N_2568);
and U6183 (N_6183,N_4940,N_3981);
or U6184 (N_6184,N_3982,N_3190);
nor U6185 (N_6185,N_3809,N_3450);
and U6186 (N_6186,N_2673,N_3015);
and U6187 (N_6187,N_4607,N_4239);
and U6188 (N_6188,N_3128,N_3586);
nor U6189 (N_6189,N_4730,N_4688);
nand U6190 (N_6190,N_2509,N_2548);
or U6191 (N_6191,N_4367,N_3031);
or U6192 (N_6192,N_2517,N_3388);
nor U6193 (N_6193,N_2553,N_2936);
nand U6194 (N_6194,N_4070,N_3659);
nor U6195 (N_6195,N_4559,N_3201);
xor U6196 (N_6196,N_3906,N_3195);
nand U6197 (N_6197,N_4397,N_4391);
nor U6198 (N_6198,N_4111,N_3494);
and U6199 (N_6199,N_3871,N_3279);
or U6200 (N_6200,N_3602,N_3889);
or U6201 (N_6201,N_4004,N_4900);
nor U6202 (N_6202,N_4945,N_2830);
nor U6203 (N_6203,N_4455,N_4424);
and U6204 (N_6204,N_3458,N_3998);
and U6205 (N_6205,N_3512,N_3132);
nand U6206 (N_6206,N_3466,N_3541);
nand U6207 (N_6207,N_2952,N_3147);
or U6208 (N_6208,N_3040,N_4338);
nand U6209 (N_6209,N_2562,N_2768);
or U6210 (N_6210,N_3133,N_2988);
or U6211 (N_6211,N_3610,N_3989);
nand U6212 (N_6212,N_4749,N_3840);
xnor U6213 (N_6213,N_2855,N_3169);
nand U6214 (N_6214,N_2615,N_3972);
or U6215 (N_6215,N_4517,N_3991);
nand U6216 (N_6216,N_3670,N_4087);
xor U6217 (N_6217,N_4763,N_4667);
nand U6218 (N_6218,N_4519,N_4664);
or U6219 (N_6219,N_2831,N_4675);
nand U6220 (N_6220,N_3052,N_3720);
and U6221 (N_6221,N_4263,N_4385);
or U6222 (N_6222,N_3590,N_4683);
nand U6223 (N_6223,N_4389,N_4150);
and U6224 (N_6224,N_3008,N_2850);
nand U6225 (N_6225,N_4192,N_4993);
nor U6226 (N_6226,N_2964,N_3598);
xor U6227 (N_6227,N_4658,N_2834);
or U6228 (N_6228,N_4440,N_3828);
or U6229 (N_6229,N_4466,N_3350);
and U6230 (N_6230,N_3447,N_3174);
or U6231 (N_6231,N_3509,N_4003);
or U6232 (N_6232,N_4120,N_4836);
and U6233 (N_6233,N_3109,N_3237);
and U6234 (N_6234,N_2872,N_2908);
and U6235 (N_6235,N_4328,N_4513);
nand U6236 (N_6236,N_2741,N_4974);
nor U6237 (N_6237,N_4692,N_4788);
or U6238 (N_6238,N_4402,N_3611);
or U6239 (N_6239,N_3690,N_4546);
or U6240 (N_6240,N_4390,N_2682);
nor U6241 (N_6241,N_4361,N_4025);
or U6242 (N_6242,N_4165,N_3268);
nand U6243 (N_6243,N_4016,N_3667);
nor U6244 (N_6244,N_3028,N_3863);
and U6245 (N_6245,N_4617,N_3759);
or U6246 (N_6246,N_4783,N_3385);
nor U6247 (N_6247,N_3084,N_4072);
or U6248 (N_6248,N_3022,N_2987);
or U6249 (N_6249,N_4691,N_4156);
and U6250 (N_6250,N_3995,N_2654);
or U6251 (N_6251,N_3119,N_4838);
and U6252 (N_6252,N_3916,N_3442);
or U6253 (N_6253,N_2985,N_2851);
nand U6254 (N_6254,N_3844,N_3987);
or U6255 (N_6255,N_4123,N_3779);
or U6256 (N_6256,N_3448,N_3872);
or U6257 (N_6257,N_4849,N_3701);
or U6258 (N_6258,N_2636,N_3199);
nor U6259 (N_6259,N_4973,N_2544);
and U6260 (N_6260,N_4314,N_3175);
nand U6261 (N_6261,N_4224,N_3238);
and U6262 (N_6262,N_4583,N_4448);
nand U6263 (N_6263,N_4366,N_3243);
nand U6264 (N_6264,N_3832,N_2681);
and U6265 (N_6265,N_3024,N_2713);
and U6266 (N_6266,N_4178,N_4365);
or U6267 (N_6267,N_3433,N_3958);
nor U6268 (N_6268,N_3116,N_3717);
or U6269 (N_6269,N_4078,N_3066);
or U6270 (N_6270,N_2872,N_3807);
nor U6271 (N_6271,N_3099,N_3230);
and U6272 (N_6272,N_4165,N_3770);
nor U6273 (N_6273,N_2813,N_3834);
and U6274 (N_6274,N_4268,N_3414);
nand U6275 (N_6275,N_3205,N_3739);
nor U6276 (N_6276,N_2832,N_3902);
or U6277 (N_6277,N_2717,N_4579);
and U6278 (N_6278,N_3230,N_3892);
nor U6279 (N_6279,N_2510,N_3965);
or U6280 (N_6280,N_3987,N_2520);
nor U6281 (N_6281,N_2750,N_2860);
and U6282 (N_6282,N_2967,N_4422);
or U6283 (N_6283,N_3304,N_4409);
nor U6284 (N_6284,N_3255,N_3902);
nor U6285 (N_6285,N_2635,N_4396);
nand U6286 (N_6286,N_4513,N_3937);
or U6287 (N_6287,N_4953,N_4598);
or U6288 (N_6288,N_4471,N_2628);
or U6289 (N_6289,N_3315,N_3439);
nand U6290 (N_6290,N_2631,N_4247);
nor U6291 (N_6291,N_2569,N_3006);
and U6292 (N_6292,N_4792,N_2939);
nor U6293 (N_6293,N_2828,N_4310);
and U6294 (N_6294,N_4045,N_3612);
and U6295 (N_6295,N_4939,N_2962);
or U6296 (N_6296,N_3354,N_4331);
and U6297 (N_6297,N_4547,N_3299);
nor U6298 (N_6298,N_2844,N_4539);
nor U6299 (N_6299,N_2514,N_2976);
or U6300 (N_6300,N_4904,N_3587);
or U6301 (N_6301,N_2865,N_4629);
or U6302 (N_6302,N_4979,N_2883);
nor U6303 (N_6303,N_2664,N_4924);
and U6304 (N_6304,N_4928,N_3908);
nor U6305 (N_6305,N_4047,N_3423);
and U6306 (N_6306,N_3467,N_3505);
and U6307 (N_6307,N_3037,N_2926);
nand U6308 (N_6308,N_3870,N_4634);
nor U6309 (N_6309,N_4770,N_3685);
nand U6310 (N_6310,N_3095,N_3085);
nand U6311 (N_6311,N_2701,N_3693);
xnor U6312 (N_6312,N_3823,N_4092);
and U6313 (N_6313,N_3613,N_3163);
or U6314 (N_6314,N_2850,N_2806);
nand U6315 (N_6315,N_2569,N_3631);
nand U6316 (N_6316,N_3280,N_4285);
nand U6317 (N_6317,N_4177,N_4625);
or U6318 (N_6318,N_3000,N_3742);
nor U6319 (N_6319,N_3617,N_4283);
and U6320 (N_6320,N_3958,N_2601);
nand U6321 (N_6321,N_2797,N_2509);
nand U6322 (N_6322,N_4951,N_3352);
and U6323 (N_6323,N_3091,N_4542);
and U6324 (N_6324,N_4239,N_3151);
nand U6325 (N_6325,N_4734,N_3152);
nor U6326 (N_6326,N_4999,N_3255);
nor U6327 (N_6327,N_4776,N_2636);
or U6328 (N_6328,N_4974,N_4695);
nor U6329 (N_6329,N_3013,N_3856);
or U6330 (N_6330,N_4545,N_3628);
or U6331 (N_6331,N_3860,N_3610);
or U6332 (N_6332,N_4914,N_2975);
and U6333 (N_6333,N_2993,N_2701);
nand U6334 (N_6334,N_4183,N_4725);
and U6335 (N_6335,N_2851,N_4115);
or U6336 (N_6336,N_4830,N_3991);
nand U6337 (N_6337,N_2640,N_4578);
nand U6338 (N_6338,N_2767,N_3171);
or U6339 (N_6339,N_3051,N_4716);
and U6340 (N_6340,N_4955,N_4887);
nand U6341 (N_6341,N_2747,N_3565);
nor U6342 (N_6342,N_4913,N_4776);
and U6343 (N_6343,N_4870,N_3882);
nand U6344 (N_6344,N_3360,N_3646);
nor U6345 (N_6345,N_3091,N_4987);
and U6346 (N_6346,N_3216,N_4975);
and U6347 (N_6347,N_2832,N_4377);
or U6348 (N_6348,N_4918,N_4401);
nor U6349 (N_6349,N_4998,N_2694);
nand U6350 (N_6350,N_3968,N_3806);
nand U6351 (N_6351,N_4963,N_4796);
and U6352 (N_6352,N_2878,N_4816);
xnor U6353 (N_6353,N_3383,N_3832);
nand U6354 (N_6354,N_4701,N_3280);
or U6355 (N_6355,N_3491,N_4541);
nor U6356 (N_6356,N_4055,N_3122);
xnor U6357 (N_6357,N_2566,N_3258);
or U6358 (N_6358,N_3451,N_3382);
nor U6359 (N_6359,N_4368,N_3549);
or U6360 (N_6360,N_4004,N_4937);
or U6361 (N_6361,N_2820,N_3098);
or U6362 (N_6362,N_4533,N_4206);
nor U6363 (N_6363,N_2802,N_3007);
nand U6364 (N_6364,N_2985,N_4910);
or U6365 (N_6365,N_3503,N_4581);
or U6366 (N_6366,N_3667,N_2837);
nor U6367 (N_6367,N_3850,N_2882);
nand U6368 (N_6368,N_4659,N_4330);
nor U6369 (N_6369,N_3177,N_3872);
nand U6370 (N_6370,N_2712,N_3409);
and U6371 (N_6371,N_3209,N_2681);
and U6372 (N_6372,N_2773,N_3260);
nor U6373 (N_6373,N_4827,N_2569);
nand U6374 (N_6374,N_3331,N_2786);
nand U6375 (N_6375,N_3541,N_3662);
nor U6376 (N_6376,N_4341,N_2836);
or U6377 (N_6377,N_4573,N_4261);
and U6378 (N_6378,N_4977,N_2926);
nand U6379 (N_6379,N_4092,N_3982);
or U6380 (N_6380,N_4175,N_2567);
nor U6381 (N_6381,N_2930,N_4549);
nand U6382 (N_6382,N_3649,N_4406);
or U6383 (N_6383,N_2579,N_3252);
nand U6384 (N_6384,N_2562,N_3036);
and U6385 (N_6385,N_3617,N_4902);
nand U6386 (N_6386,N_4337,N_4762);
nor U6387 (N_6387,N_2605,N_3415);
nor U6388 (N_6388,N_2649,N_2647);
nor U6389 (N_6389,N_3284,N_2776);
or U6390 (N_6390,N_3904,N_4507);
nor U6391 (N_6391,N_2908,N_2775);
nor U6392 (N_6392,N_3964,N_4789);
nor U6393 (N_6393,N_3177,N_4558);
and U6394 (N_6394,N_3650,N_4178);
nand U6395 (N_6395,N_3711,N_2522);
or U6396 (N_6396,N_4382,N_3204);
nor U6397 (N_6397,N_2847,N_3908);
or U6398 (N_6398,N_4088,N_3050);
nand U6399 (N_6399,N_3947,N_2537);
and U6400 (N_6400,N_3302,N_4685);
nor U6401 (N_6401,N_4378,N_4341);
or U6402 (N_6402,N_3224,N_2922);
and U6403 (N_6403,N_3041,N_4406);
or U6404 (N_6404,N_4873,N_3351);
nand U6405 (N_6405,N_3677,N_4853);
nor U6406 (N_6406,N_3499,N_4556);
nand U6407 (N_6407,N_3124,N_4013);
and U6408 (N_6408,N_4764,N_4845);
or U6409 (N_6409,N_2662,N_4082);
nand U6410 (N_6410,N_4215,N_3999);
or U6411 (N_6411,N_3618,N_4906);
and U6412 (N_6412,N_4093,N_2597);
nand U6413 (N_6413,N_2627,N_4263);
or U6414 (N_6414,N_4683,N_4337);
or U6415 (N_6415,N_2803,N_2628);
and U6416 (N_6416,N_3659,N_4402);
or U6417 (N_6417,N_2923,N_2568);
or U6418 (N_6418,N_3220,N_3828);
and U6419 (N_6419,N_4941,N_4475);
nand U6420 (N_6420,N_3286,N_3370);
nor U6421 (N_6421,N_4900,N_3673);
and U6422 (N_6422,N_4772,N_2736);
and U6423 (N_6423,N_4235,N_4811);
nand U6424 (N_6424,N_4535,N_2940);
nor U6425 (N_6425,N_3581,N_2732);
or U6426 (N_6426,N_3812,N_3263);
or U6427 (N_6427,N_4285,N_3927);
or U6428 (N_6428,N_4980,N_3834);
or U6429 (N_6429,N_3580,N_3924);
nor U6430 (N_6430,N_4619,N_4936);
nand U6431 (N_6431,N_4067,N_3123);
nand U6432 (N_6432,N_4570,N_4568);
or U6433 (N_6433,N_4361,N_3281);
or U6434 (N_6434,N_2777,N_4729);
or U6435 (N_6435,N_4456,N_4943);
nand U6436 (N_6436,N_3711,N_3005);
or U6437 (N_6437,N_4486,N_3316);
or U6438 (N_6438,N_2949,N_3639);
or U6439 (N_6439,N_2780,N_4501);
or U6440 (N_6440,N_2616,N_4826);
or U6441 (N_6441,N_3417,N_4158);
xnor U6442 (N_6442,N_2680,N_2666);
nor U6443 (N_6443,N_4685,N_3474);
and U6444 (N_6444,N_4243,N_4417);
nand U6445 (N_6445,N_2993,N_3525);
or U6446 (N_6446,N_3787,N_4069);
and U6447 (N_6447,N_4054,N_4852);
nand U6448 (N_6448,N_3057,N_2771);
nand U6449 (N_6449,N_2701,N_3874);
nand U6450 (N_6450,N_2956,N_3168);
nand U6451 (N_6451,N_3453,N_3468);
nand U6452 (N_6452,N_4374,N_3370);
nor U6453 (N_6453,N_4783,N_3639);
nor U6454 (N_6454,N_2522,N_3645);
nand U6455 (N_6455,N_2893,N_2770);
and U6456 (N_6456,N_3035,N_4552);
nor U6457 (N_6457,N_4805,N_3713);
nand U6458 (N_6458,N_4992,N_2797);
nor U6459 (N_6459,N_2656,N_4604);
or U6460 (N_6460,N_2643,N_2727);
nand U6461 (N_6461,N_4696,N_3964);
and U6462 (N_6462,N_2810,N_4865);
nor U6463 (N_6463,N_3516,N_3302);
or U6464 (N_6464,N_2516,N_4003);
or U6465 (N_6465,N_2755,N_2789);
and U6466 (N_6466,N_4354,N_3938);
or U6467 (N_6467,N_3335,N_4695);
or U6468 (N_6468,N_2569,N_3900);
and U6469 (N_6469,N_4100,N_3787);
and U6470 (N_6470,N_2791,N_2765);
or U6471 (N_6471,N_3192,N_3873);
nand U6472 (N_6472,N_4268,N_2503);
or U6473 (N_6473,N_4652,N_2977);
or U6474 (N_6474,N_3033,N_3976);
or U6475 (N_6475,N_4596,N_3470);
nand U6476 (N_6476,N_3201,N_3568);
or U6477 (N_6477,N_3881,N_4707);
nor U6478 (N_6478,N_3993,N_3435);
and U6479 (N_6479,N_3144,N_3471);
nand U6480 (N_6480,N_3452,N_4146);
nor U6481 (N_6481,N_4577,N_4495);
nor U6482 (N_6482,N_4343,N_3068);
or U6483 (N_6483,N_3094,N_3102);
or U6484 (N_6484,N_4656,N_3183);
or U6485 (N_6485,N_2792,N_3232);
or U6486 (N_6486,N_4008,N_4065);
nand U6487 (N_6487,N_4302,N_3672);
nand U6488 (N_6488,N_3592,N_2620);
and U6489 (N_6489,N_4770,N_3800);
nor U6490 (N_6490,N_3611,N_4141);
and U6491 (N_6491,N_4625,N_2728);
nand U6492 (N_6492,N_2670,N_3845);
nand U6493 (N_6493,N_4273,N_3440);
nand U6494 (N_6494,N_4016,N_4953);
or U6495 (N_6495,N_3582,N_4878);
or U6496 (N_6496,N_3304,N_4449);
nand U6497 (N_6497,N_4274,N_2992);
nand U6498 (N_6498,N_4240,N_4412);
nor U6499 (N_6499,N_4557,N_4076);
nand U6500 (N_6500,N_2730,N_2804);
or U6501 (N_6501,N_4810,N_3834);
and U6502 (N_6502,N_4362,N_2683);
nor U6503 (N_6503,N_2709,N_3713);
nor U6504 (N_6504,N_4004,N_4164);
and U6505 (N_6505,N_3244,N_3813);
and U6506 (N_6506,N_4943,N_2691);
nand U6507 (N_6507,N_2618,N_2989);
nor U6508 (N_6508,N_3833,N_3159);
or U6509 (N_6509,N_4048,N_3741);
or U6510 (N_6510,N_2629,N_4902);
and U6511 (N_6511,N_4001,N_4209);
and U6512 (N_6512,N_3033,N_3691);
or U6513 (N_6513,N_4977,N_4858);
and U6514 (N_6514,N_4550,N_3472);
and U6515 (N_6515,N_4310,N_3370);
and U6516 (N_6516,N_2548,N_2939);
or U6517 (N_6517,N_4962,N_3173);
nand U6518 (N_6518,N_3812,N_4830);
or U6519 (N_6519,N_2592,N_4279);
or U6520 (N_6520,N_4594,N_2516);
or U6521 (N_6521,N_3941,N_2597);
nand U6522 (N_6522,N_4551,N_4419);
or U6523 (N_6523,N_4395,N_4694);
nor U6524 (N_6524,N_2572,N_3141);
nand U6525 (N_6525,N_3810,N_4988);
nand U6526 (N_6526,N_4171,N_3505);
or U6527 (N_6527,N_2638,N_4365);
nand U6528 (N_6528,N_3690,N_4856);
and U6529 (N_6529,N_3439,N_3736);
nor U6530 (N_6530,N_3528,N_3403);
or U6531 (N_6531,N_4933,N_4497);
or U6532 (N_6532,N_3837,N_4773);
nor U6533 (N_6533,N_4679,N_3093);
or U6534 (N_6534,N_4260,N_4566);
nor U6535 (N_6535,N_4164,N_2865);
or U6536 (N_6536,N_4011,N_4800);
nor U6537 (N_6537,N_4733,N_4800);
nor U6538 (N_6538,N_4896,N_4554);
nand U6539 (N_6539,N_4105,N_2516);
or U6540 (N_6540,N_3506,N_3576);
or U6541 (N_6541,N_2865,N_3429);
and U6542 (N_6542,N_2755,N_4351);
and U6543 (N_6543,N_2744,N_4559);
nand U6544 (N_6544,N_4051,N_3617);
nor U6545 (N_6545,N_3188,N_4154);
nor U6546 (N_6546,N_3380,N_4132);
nor U6547 (N_6547,N_4462,N_3796);
nor U6548 (N_6548,N_4416,N_3146);
nor U6549 (N_6549,N_3097,N_2522);
or U6550 (N_6550,N_4061,N_4037);
nor U6551 (N_6551,N_3676,N_3048);
or U6552 (N_6552,N_4128,N_3617);
nor U6553 (N_6553,N_3335,N_3265);
nand U6554 (N_6554,N_2767,N_2780);
or U6555 (N_6555,N_2930,N_3211);
and U6556 (N_6556,N_3791,N_4041);
or U6557 (N_6557,N_3056,N_4555);
nor U6558 (N_6558,N_4571,N_3657);
nand U6559 (N_6559,N_3221,N_4126);
nor U6560 (N_6560,N_2741,N_3566);
xor U6561 (N_6561,N_4045,N_4083);
nand U6562 (N_6562,N_4692,N_3988);
or U6563 (N_6563,N_4453,N_3418);
or U6564 (N_6564,N_3839,N_3771);
and U6565 (N_6565,N_3783,N_4974);
and U6566 (N_6566,N_3555,N_3839);
nor U6567 (N_6567,N_3530,N_4293);
nor U6568 (N_6568,N_3959,N_4817);
or U6569 (N_6569,N_2739,N_3465);
nor U6570 (N_6570,N_4708,N_3806);
nand U6571 (N_6571,N_3717,N_4807);
nor U6572 (N_6572,N_4398,N_3341);
nand U6573 (N_6573,N_3757,N_3655);
nor U6574 (N_6574,N_4640,N_3541);
nand U6575 (N_6575,N_2758,N_2663);
and U6576 (N_6576,N_3370,N_4601);
nand U6577 (N_6577,N_4725,N_4086);
nand U6578 (N_6578,N_4059,N_4853);
or U6579 (N_6579,N_3986,N_4378);
nor U6580 (N_6580,N_4934,N_2574);
and U6581 (N_6581,N_2886,N_3451);
or U6582 (N_6582,N_2683,N_3283);
and U6583 (N_6583,N_3991,N_4903);
or U6584 (N_6584,N_3000,N_3524);
nand U6585 (N_6585,N_4026,N_4297);
or U6586 (N_6586,N_3390,N_4318);
and U6587 (N_6587,N_3339,N_4253);
nor U6588 (N_6588,N_3407,N_2995);
nand U6589 (N_6589,N_4079,N_3474);
or U6590 (N_6590,N_4265,N_4238);
and U6591 (N_6591,N_2511,N_3879);
nor U6592 (N_6592,N_3254,N_3548);
and U6593 (N_6593,N_4498,N_2588);
nand U6594 (N_6594,N_3774,N_3238);
or U6595 (N_6595,N_3077,N_3900);
or U6596 (N_6596,N_3263,N_3655);
or U6597 (N_6597,N_4339,N_2801);
and U6598 (N_6598,N_4160,N_3716);
or U6599 (N_6599,N_4765,N_4338);
or U6600 (N_6600,N_4048,N_4257);
nand U6601 (N_6601,N_3662,N_3503);
or U6602 (N_6602,N_3109,N_3999);
and U6603 (N_6603,N_3022,N_4412);
xor U6604 (N_6604,N_2661,N_4158);
nor U6605 (N_6605,N_3640,N_3351);
nor U6606 (N_6606,N_4223,N_4690);
nor U6607 (N_6607,N_4346,N_4083);
nor U6608 (N_6608,N_4555,N_3169);
nor U6609 (N_6609,N_4476,N_3353);
or U6610 (N_6610,N_4198,N_4345);
and U6611 (N_6611,N_4564,N_3111);
and U6612 (N_6612,N_4062,N_2729);
or U6613 (N_6613,N_4676,N_3087);
nand U6614 (N_6614,N_3160,N_2861);
or U6615 (N_6615,N_3063,N_2714);
nand U6616 (N_6616,N_2890,N_4585);
and U6617 (N_6617,N_3446,N_2889);
nand U6618 (N_6618,N_2850,N_3309);
nor U6619 (N_6619,N_4833,N_3557);
and U6620 (N_6620,N_2661,N_4392);
nor U6621 (N_6621,N_2846,N_3033);
nor U6622 (N_6622,N_2778,N_4767);
nor U6623 (N_6623,N_4392,N_2971);
nand U6624 (N_6624,N_3650,N_4968);
nor U6625 (N_6625,N_2570,N_3826);
nand U6626 (N_6626,N_4482,N_3053);
and U6627 (N_6627,N_4836,N_3873);
nand U6628 (N_6628,N_3199,N_3147);
and U6629 (N_6629,N_4164,N_4105);
and U6630 (N_6630,N_3851,N_4694);
or U6631 (N_6631,N_4415,N_3574);
and U6632 (N_6632,N_3326,N_2881);
or U6633 (N_6633,N_4405,N_2568);
nor U6634 (N_6634,N_4957,N_4959);
nor U6635 (N_6635,N_4637,N_4246);
nand U6636 (N_6636,N_4848,N_3589);
and U6637 (N_6637,N_2528,N_4160);
nand U6638 (N_6638,N_3150,N_3032);
nand U6639 (N_6639,N_4196,N_3371);
or U6640 (N_6640,N_3558,N_2587);
and U6641 (N_6641,N_3490,N_4118);
nor U6642 (N_6642,N_4913,N_4448);
nand U6643 (N_6643,N_4120,N_3749);
nor U6644 (N_6644,N_4612,N_2810);
or U6645 (N_6645,N_4080,N_4415);
nor U6646 (N_6646,N_3327,N_4877);
nand U6647 (N_6647,N_4683,N_2671);
nand U6648 (N_6648,N_4908,N_4242);
nand U6649 (N_6649,N_4387,N_3620);
nor U6650 (N_6650,N_4272,N_4810);
or U6651 (N_6651,N_3753,N_4053);
and U6652 (N_6652,N_2856,N_2535);
nand U6653 (N_6653,N_3469,N_3530);
nand U6654 (N_6654,N_4853,N_4516);
nand U6655 (N_6655,N_2602,N_3911);
nor U6656 (N_6656,N_4317,N_4818);
or U6657 (N_6657,N_4931,N_4161);
nand U6658 (N_6658,N_4378,N_2749);
and U6659 (N_6659,N_4136,N_3943);
or U6660 (N_6660,N_3733,N_3234);
nor U6661 (N_6661,N_4647,N_3871);
and U6662 (N_6662,N_3168,N_3514);
nand U6663 (N_6663,N_4160,N_3746);
nor U6664 (N_6664,N_4418,N_4032);
or U6665 (N_6665,N_3707,N_4620);
or U6666 (N_6666,N_3530,N_4964);
nor U6667 (N_6667,N_3518,N_4425);
nand U6668 (N_6668,N_4031,N_4535);
nand U6669 (N_6669,N_4574,N_4219);
or U6670 (N_6670,N_4266,N_4624);
nand U6671 (N_6671,N_3694,N_2504);
nor U6672 (N_6672,N_4261,N_4788);
nand U6673 (N_6673,N_3975,N_2696);
nand U6674 (N_6674,N_4631,N_3632);
and U6675 (N_6675,N_3730,N_4635);
nand U6676 (N_6676,N_4289,N_4248);
nand U6677 (N_6677,N_4816,N_4802);
nor U6678 (N_6678,N_2882,N_3550);
and U6679 (N_6679,N_3362,N_4983);
and U6680 (N_6680,N_4774,N_3903);
and U6681 (N_6681,N_4124,N_3187);
and U6682 (N_6682,N_4390,N_2750);
nor U6683 (N_6683,N_3177,N_4273);
and U6684 (N_6684,N_4645,N_2723);
nor U6685 (N_6685,N_2552,N_4822);
nand U6686 (N_6686,N_4823,N_3146);
nand U6687 (N_6687,N_3306,N_3266);
and U6688 (N_6688,N_4383,N_4491);
nor U6689 (N_6689,N_4349,N_3890);
or U6690 (N_6690,N_4774,N_3890);
nor U6691 (N_6691,N_3044,N_3983);
and U6692 (N_6692,N_3042,N_3060);
and U6693 (N_6693,N_2722,N_4041);
and U6694 (N_6694,N_4822,N_2607);
nor U6695 (N_6695,N_4856,N_3792);
and U6696 (N_6696,N_2549,N_4787);
nand U6697 (N_6697,N_3684,N_4408);
nor U6698 (N_6698,N_4756,N_3106);
or U6699 (N_6699,N_3951,N_3030);
nand U6700 (N_6700,N_3984,N_3791);
and U6701 (N_6701,N_3106,N_3542);
or U6702 (N_6702,N_4688,N_4475);
and U6703 (N_6703,N_4604,N_2757);
nor U6704 (N_6704,N_2605,N_3520);
or U6705 (N_6705,N_4819,N_2849);
nor U6706 (N_6706,N_3459,N_3397);
nor U6707 (N_6707,N_4277,N_4317);
nor U6708 (N_6708,N_3985,N_2537);
nand U6709 (N_6709,N_4936,N_4798);
and U6710 (N_6710,N_2646,N_4377);
nor U6711 (N_6711,N_3383,N_3174);
nand U6712 (N_6712,N_3652,N_4624);
or U6713 (N_6713,N_4112,N_4878);
nor U6714 (N_6714,N_2564,N_4505);
or U6715 (N_6715,N_3463,N_2616);
and U6716 (N_6716,N_4169,N_2579);
or U6717 (N_6717,N_4228,N_4026);
or U6718 (N_6718,N_2991,N_2588);
or U6719 (N_6719,N_4079,N_4446);
or U6720 (N_6720,N_3904,N_4743);
or U6721 (N_6721,N_3167,N_3584);
nand U6722 (N_6722,N_3331,N_4788);
and U6723 (N_6723,N_3953,N_3493);
nor U6724 (N_6724,N_3607,N_2604);
and U6725 (N_6725,N_4781,N_2626);
or U6726 (N_6726,N_4463,N_3312);
or U6727 (N_6727,N_3127,N_4865);
nand U6728 (N_6728,N_3437,N_2714);
nand U6729 (N_6729,N_4826,N_2556);
nand U6730 (N_6730,N_4029,N_4697);
nand U6731 (N_6731,N_4320,N_2537);
and U6732 (N_6732,N_3682,N_4304);
nand U6733 (N_6733,N_4876,N_2689);
and U6734 (N_6734,N_3008,N_2958);
nand U6735 (N_6735,N_3617,N_4348);
and U6736 (N_6736,N_3838,N_3514);
nor U6737 (N_6737,N_3860,N_3566);
nand U6738 (N_6738,N_3591,N_4866);
xor U6739 (N_6739,N_3659,N_4392);
nand U6740 (N_6740,N_3286,N_3004);
nand U6741 (N_6741,N_3763,N_2904);
and U6742 (N_6742,N_4779,N_4507);
or U6743 (N_6743,N_4753,N_3236);
or U6744 (N_6744,N_3179,N_2773);
nor U6745 (N_6745,N_3527,N_2639);
and U6746 (N_6746,N_4464,N_2815);
nand U6747 (N_6747,N_3280,N_3810);
nor U6748 (N_6748,N_2760,N_4228);
nand U6749 (N_6749,N_3993,N_4689);
nor U6750 (N_6750,N_3058,N_3348);
or U6751 (N_6751,N_3958,N_4959);
and U6752 (N_6752,N_4283,N_4842);
nand U6753 (N_6753,N_3713,N_4282);
nand U6754 (N_6754,N_4484,N_3959);
nand U6755 (N_6755,N_4279,N_4570);
nand U6756 (N_6756,N_4797,N_4908);
and U6757 (N_6757,N_2686,N_3487);
and U6758 (N_6758,N_2828,N_4907);
and U6759 (N_6759,N_3448,N_4189);
nand U6760 (N_6760,N_4093,N_2973);
nand U6761 (N_6761,N_2987,N_3796);
nand U6762 (N_6762,N_4558,N_3375);
nor U6763 (N_6763,N_2871,N_2815);
nor U6764 (N_6764,N_2715,N_2663);
and U6765 (N_6765,N_3417,N_3603);
and U6766 (N_6766,N_3136,N_4642);
or U6767 (N_6767,N_4262,N_2644);
nor U6768 (N_6768,N_2882,N_4685);
and U6769 (N_6769,N_3862,N_4074);
and U6770 (N_6770,N_4998,N_2857);
nor U6771 (N_6771,N_3557,N_3996);
nor U6772 (N_6772,N_4287,N_4696);
nor U6773 (N_6773,N_4744,N_4795);
or U6774 (N_6774,N_2534,N_4456);
nand U6775 (N_6775,N_3929,N_3499);
or U6776 (N_6776,N_3306,N_4195);
and U6777 (N_6777,N_4485,N_2921);
or U6778 (N_6778,N_3454,N_4656);
or U6779 (N_6779,N_3298,N_4719);
or U6780 (N_6780,N_3339,N_2834);
nand U6781 (N_6781,N_4950,N_2916);
and U6782 (N_6782,N_2547,N_4456);
or U6783 (N_6783,N_4746,N_4015);
nand U6784 (N_6784,N_2671,N_3246);
nand U6785 (N_6785,N_3516,N_4205);
nor U6786 (N_6786,N_3279,N_3134);
nand U6787 (N_6787,N_2760,N_3048);
nor U6788 (N_6788,N_3076,N_4330);
nand U6789 (N_6789,N_3228,N_3125);
and U6790 (N_6790,N_3326,N_3661);
and U6791 (N_6791,N_2747,N_3756);
and U6792 (N_6792,N_2795,N_4016);
or U6793 (N_6793,N_4898,N_3688);
or U6794 (N_6794,N_2605,N_2687);
nor U6795 (N_6795,N_3705,N_3972);
and U6796 (N_6796,N_3471,N_3502);
or U6797 (N_6797,N_3388,N_3679);
and U6798 (N_6798,N_2826,N_4965);
or U6799 (N_6799,N_3457,N_4404);
or U6800 (N_6800,N_3344,N_3729);
nand U6801 (N_6801,N_3372,N_3565);
and U6802 (N_6802,N_4627,N_4292);
nor U6803 (N_6803,N_3415,N_3474);
or U6804 (N_6804,N_3041,N_2542);
and U6805 (N_6805,N_2725,N_4580);
and U6806 (N_6806,N_4291,N_4586);
or U6807 (N_6807,N_3602,N_4978);
and U6808 (N_6808,N_4064,N_2571);
or U6809 (N_6809,N_2849,N_3562);
nor U6810 (N_6810,N_3009,N_2712);
nand U6811 (N_6811,N_4719,N_2673);
nor U6812 (N_6812,N_4888,N_3205);
nor U6813 (N_6813,N_4809,N_4804);
nand U6814 (N_6814,N_4085,N_4415);
nor U6815 (N_6815,N_3357,N_4361);
or U6816 (N_6816,N_4374,N_3789);
nor U6817 (N_6817,N_3816,N_3849);
nand U6818 (N_6818,N_2572,N_3890);
or U6819 (N_6819,N_4166,N_2551);
or U6820 (N_6820,N_4501,N_4619);
nand U6821 (N_6821,N_4666,N_3672);
nor U6822 (N_6822,N_2728,N_4388);
or U6823 (N_6823,N_4961,N_3284);
and U6824 (N_6824,N_3364,N_4308);
nor U6825 (N_6825,N_2513,N_3144);
nand U6826 (N_6826,N_3629,N_4617);
nand U6827 (N_6827,N_3766,N_3000);
or U6828 (N_6828,N_3938,N_2759);
nor U6829 (N_6829,N_2770,N_4511);
nor U6830 (N_6830,N_3086,N_4515);
nor U6831 (N_6831,N_3622,N_2789);
xnor U6832 (N_6832,N_4337,N_4423);
nor U6833 (N_6833,N_4333,N_4139);
or U6834 (N_6834,N_3490,N_4325);
and U6835 (N_6835,N_3551,N_3603);
and U6836 (N_6836,N_4204,N_4648);
or U6837 (N_6837,N_4121,N_3146);
nand U6838 (N_6838,N_4625,N_4477);
nand U6839 (N_6839,N_3243,N_2548);
nand U6840 (N_6840,N_4457,N_4489);
and U6841 (N_6841,N_3255,N_3249);
nor U6842 (N_6842,N_3985,N_4546);
nand U6843 (N_6843,N_2873,N_3917);
and U6844 (N_6844,N_3792,N_2703);
nor U6845 (N_6845,N_3836,N_4513);
or U6846 (N_6846,N_4941,N_4437);
nor U6847 (N_6847,N_4480,N_2570);
nand U6848 (N_6848,N_3471,N_3364);
nand U6849 (N_6849,N_2675,N_3545);
nand U6850 (N_6850,N_4278,N_4593);
nand U6851 (N_6851,N_3494,N_4215);
or U6852 (N_6852,N_3270,N_3851);
or U6853 (N_6853,N_4216,N_3020);
and U6854 (N_6854,N_2973,N_4811);
and U6855 (N_6855,N_2747,N_4423);
and U6856 (N_6856,N_4844,N_4432);
or U6857 (N_6857,N_3367,N_3210);
nand U6858 (N_6858,N_3381,N_4186);
and U6859 (N_6859,N_2838,N_3153);
nor U6860 (N_6860,N_3095,N_3614);
or U6861 (N_6861,N_3807,N_4942);
nand U6862 (N_6862,N_4258,N_3740);
nand U6863 (N_6863,N_2804,N_2936);
nand U6864 (N_6864,N_4179,N_4045);
nand U6865 (N_6865,N_2859,N_2721);
nor U6866 (N_6866,N_2588,N_4275);
or U6867 (N_6867,N_2511,N_3269);
and U6868 (N_6868,N_4681,N_3681);
or U6869 (N_6869,N_2527,N_4248);
nand U6870 (N_6870,N_4154,N_4524);
or U6871 (N_6871,N_3735,N_3622);
or U6872 (N_6872,N_2870,N_4353);
nand U6873 (N_6873,N_2508,N_4669);
nand U6874 (N_6874,N_2957,N_4273);
and U6875 (N_6875,N_3984,N_2862);
nor U6876 (N_6876,N_4079,N_4336);
or U6877 (N_6877,N_4712,N_4777);
nor U6878 (N_6878,N_4212,N_4588);
nand U6879 (N_6879,N_4561,N_4626);
nand U6880 (N_6880,N_3250,N_2961);
nand U6881 (N_6881,N_4874,N_4038);
nand U6882 (N_6882,N_4888,N_3584);
nor U6883 (N_6883,N_4521,N_3454);
nor U6884 (N_6884,N_4631,N_3901);
and U6885 (N_6885,N_4408,N_3668);
nor U6886 (N_6886,N_4964,N_4157);
or U6887 (N_6887,N_3306,N_3316);
or U6888 (N_6888,N_3026,N_3666);
nand U6889 (N_6889,N_3721,N_2774);
nand U6890 (N_6890,N_2728,N_2960);
and U6891 (N_6891,N_2825,N_3268);
and U6892 (N_6892,N_2644,N_3940);
and U6893 (N_6893,N_4592,N_3741);
and U6894 (N_6894,N_3275,N_3626);
nor U6895 (N_6895,N_4887,N_3775);
or U6896 (N_6896,N_3771,N_4423);
nand U6897 (N_6897,N_4597,N_2576);
or U6898 (N_6898,N_2787,N_4971);
or U6899 (N_6899,N_4524,N_3775);
and U6900 (N_6900,N_4076,N_3774);
nor U6901 (N_6901,N_3216,N_4392);
nand U6902 (N_6902,N_4001,N_3304);
nand U6903 (N_6903,N_3848,N_2711);
nand U6904 (N_6904,N_4843,N_4550);
and U6905 (N_6905,N_2564,N_3384);
and U6906 (N_6906,N_2879,N_2858);
or U6907 (N_6907,N_4947,N_2690);
nand U6908 (N_6908,N_4920,N_3338);
and U6909 (N_6909,N_4631,N_4804);
or U6910 (N_6910,N_3009,N_4888);
or U6911 (N_6911,N_3117,N_3330);
nor U6912 (N_6912,N_3244,N_2802);
and U6913 (N_6913,N_4518,N_4156);
or U6914 (N_6914,N_4882,N_3403);
or U6915 (N_6915,N_2918,N_4711);
and U6916 (N_6916,N_2605,N_3050);
or U6917 (N_6917,N_3097,N_2519);
and U6918 (N_6918,N_3435,N_2826);
or U6919 (N_6919,N_4067,N_4806);
nand U6920 (N_6920,N_4062,N_2503);
or U6921 (N_6921,N_4480,N_2615);
nor U6922 (N_6922,N_2626,N_3056);
nand U6923 (N_6923,N_2789,N_2561);
or U6924 (N_6924,N_4180,N_4259);
nand U6925 (N_6925,N_3038,N_4513);
nor U6926 (N_6926,N_4080,N_4648);
and U6927 (N_6927,N_3625,N_4825);
and U6928 (N_6928,N_3777,N_4252);
nor U6929 (N_6929,N_4666,N_3381);
and U6930 (N_6930,N_3570,N_4904);
nand U6931 (N_6931,N_4290,N_4783);
or U6932 (N_6932,N_4618,N_4714);
or U6933 (N_6933,N_2901,N_3780);
nor U6934 (N_6934,N_3870,N_2788);
and U6935 (N_6935,N_4224,N_4331);
xor U6936 (N_6936,N_4294,N_4065);
and U6937 (N_6937,N_3412,N_4389);
nand U6938 (N_6938,N_2659,N_4459);
nand U6939 (N_6939,N_4880,N_3054);
and U6940 (N_6940,N_3982,N_3585);
or U6941 (N_6941,N_2671,N_4850);
and U6942 (N_6942,N_4546,N_4710);
nor U6943 (N_6943,N_3632,N_2818);
xor U6944 (N_6944,N_4691,N_2835);
and U6945 (N_6945,N_4894,N_4827);
nor U6946 (N_6946,N_4046,N_3410);
nand U6947 (N_6947,N_3710,N_2840);
or U6948 (N_6948,N_2911,N_3588);
nor U6949 (N_6949,N_3618,N_4040);
or U6950 (N_6950,N_4838,N_3658);
or U6951 (N_6951,N_3935,N_2995);
and U6952 (N_6952,N_2621,N_3456);
nor U6953 (N_6953,N_2520,N_4041);
nor U6954 (N_6954,N_2651,N_4397);
nor U6955 (N_6955,N_3649,N_2671);
or U6956 (N_6956,N_4181,N_3315);
nand U6957 (N_6957,N_3618,N_4219);
and U6958 (N_6958,N_4588,N_3992);
nor U6959 (N_6959,N_4492,N_3380);
nand U6960 (N_6960,N_4539,N_4378);
and U6961 (N_6961,N_3563,N_2805);
nand U6962 (N_6962,N_2715,N_2738);
or U6963 (N_6963,N_2972,N_3770);
nor U6964 (N_6964,N_3936,N_3212);
and U6965 (N_6965,N_4724,N_4574);
nand U6966 (N_6966,N_3657,N_3535);
nor U6967 (N_6967,N_4720,N_4234);
or U6968 (N_6968,N_3298,N_4929);
nand U6969 (N_6969,N_3887,N_4821);
and U6970 (N_6970,N_2704,N_4421);
or U6971 (N_6971,N_3029,N_2514);
and U6972 (N_6972,N_4204,N_4112);
nor U6973 (N_6973,N_2699,N_3975);
or U6974 (N_6974,N_3731,N_2633);
nor U6975 (N_6975,N_4672,N_3588);
nor U6976 (N_6976,N_4700,N_2826);
or U6977 (N_6977,N_3233,N_3000);
or U6978 (N_6978,N_2963,N_3864);
and U6979 (N_6979,N_2644,N_4503);
xnor U6980 (N_6980,N_3378,N_4805);
nor U6981 (N_6981,N_3213,N_4593);
or U6982 (N_6982,N_3427,N_4780);
or U6983 (N_6983,N_3334,N_2713);
nor U6984 (N_6984,N_4924,N_4646);
nor U6985 (N_6985,N_4840,N_4043);
nor U6986 (N_6986,N_3915,N_3501);
nor U6987 (N_6987,N_4682,N_3466);
nor U6988 (N_6988,N_4307,N_2998);
or U6989 (N_6989,N_4567,N_3337);
or U6990 (N_6990,N_4774,N_4276);
nand U6991 (N_6991,N_2930,N_4507);
and U6992 (N_6992,N_4134,N_3652);
nor U6993 (N_6993,N_3811,N_4443);
or U6994 (N_6994,N_2740,N_3162);
and U6995 (N_6995,N_4010,N_3703);
nor U6996 (N_6996,N_3846,N_4557);
nor U6997 (N_6997,N_4179,N_2876);
and U6998 (N_6998,N_4811,N_2954);
nor U6999 (N_6999,N_3817,N_2660);
or U7000 (N_7000,N_4783,N_4793);
or U7001 (N_7001,N_4208,N_4882);
nor U7002 (N_7002,N_3829,N_4153);
nand U7003 (N_7003,N_4938,N_2840);
nor U7004 (N_7004,N_4983,N_3237);
and U7005 (N_7005,N_4373,N_2565);
nand U7006 (N_7006,N_4897,N_3910);
or U7007 (N_7007,N_4458,N_4850);
or U7008 (N_7008,N_4425,N_4941);
xor U7009 (N_7009,N_4077,N_2885);
or U7010 (N_7010,N_3437,N_3776);
or U7011 (N_7011,N_3393,N_3864);
and U7012 (N_7012,N_2771,N_3761);
or U7013 (N_7013,N_3101,N_4367);
nand U7014 (N_7014,N_3606,N_3264);
nor U7015 (N_7015,N_4362,N_3046);
or U7016 (N_7016,N_3744,N_2574);
nor U7017 (N_7017,N_2922,N_2741);
or U7018 (N_7018,N_2865,N_3565);
nand U7019 (N_7019,N_4364,N_4955);
and U7020 (N_7020,N_4081,N_3783);
and U7021 (N_7021,N_3458,N_3501);
nor U7022 (N_7022,N_4993,N_4627);
and U7023 (N_7023,N_4635,N_4935);
nand U7024 (N_7024,N_3667,N_2521);
and U7025 (N_7025,N_3897,N_3819);
or U7026 (N_7026,N_3069,N_3421);
nor U7027 (N_7027,N_3253,N_2800);
and U7028 (N_7028,N_2850,N_3916);
nor U7029 (N_7029,N_3177,N_3063);
or U7030 (N_7030,N_3974,N_4469);
and U7031 (N_7031,N_3048,N_3042);
nor U7032 (N_7032,N_2642,N_3068);
nor U7033 (N_7033,N_3857,N_4636);
and U7034 (N_7034,N_3855,N_3262);
or U7035 (N_7035,N_4862,N_3187);
nor U7036 (N_7036,N_3971,N_3896);
or U7037 (N_7037,N_4887,N_4291);
nor U7038 (N_7038,N_4648,N_2952);
and U7039 (N_7039,N_4210,N_3242);
nand U7040 (N_7040,N_4197,N_2770);
or U7041 (N_7041,N_2664,N_2621);
nor U7042 (N_7042,N_3434,N_3945);
and U7043 (N_7043,N_4895,N_3261);
nor U7044 (N_7044,N_2661,N_4280);
and U7045 (N_7045,N_4657,N_3248);
nor U7046 (N_7046,N_3780,N_3791);
nor U7047 (N_7047,N_3267,N_3355);
nand U7048 (N_7048,N_3835,N_3017);
nor U7049 (N_7049,N_4016,N_2932);
and U7050 (N_7050,N_4486,N_4922);
or U7051 (N_7051,N_2786,N_3087);
nand U7052 (N_7052,N_3405,N_3570);
nand U7053 (N_7053,N_4143,N_3537);
and U7054 (N_7054,N_3630,N_3571);
nor U7055 (N_7055,N_3177,N_4724);
and U7056 (N_7056,N_3028,N_3007);
nand U7057 (N_7057,N_2612,N_3656);
and U7058 (N_7058,N_3865,N_3918);
or U7059 (N_7059,N_3787,N_4568);
nor U7060 (N_7060,N_3996,N_3158);
nor U7061 (N_7061,N_2733,N_4558);
or U7062 (N_7062,N_3344,N_4069);
nand U7063 (N_7063,N_3819,N_2762);
and U7064 (N_7064,N_3501,N_3103);
or U7065 (N_7065,N_4879,N_4429);
nor U7066 (N_7066,N_4524,N_3601);
nand U7067 (N_7067,N_4407,N_3324);
or U7068 (N_7068,N_3944,N_2753);
and U7069 (N_7069,N_4913,N_4105);
or U7070 (N_7070,N_2974,N_3242);
or U7071 (N_7071,N_4028,N_3414);
and U7072 (N_7072,N_4136,N_3988);
or U7073 (N_7073,N_4381,N_4640);
and U7074 (N_7074,N_2718,N_3753);
nand U7075 (N_7075,N_3401,N_4751);
nor U7076 (N_7076,N_4963,N_2898);
and U7077 (N_7077,N_4361,N_4848);
nor U7078 (N_7078,N_2877,N_4762);
or U7079 (N_7079,N_2784,N_4969);
and U7080 (N_7080,N_4149,N_4546);
and U7081 (N_7081,N_3704,N_4183);
and U7082 (N_7082,N_2703,N_3438);
nand U7083 (N_7083,N_4451,N_3909);
nand U7084 (N_7084,N_3784,N_4146);
or U7085 (N_7085,N_4375,N_2618);
nand U7086 (N_7086,N_4097,N_3940);
nand U7087 (N_7087,N_4387,N_2586);
or U7088 (N_7088,N_4388,N_3369);
and U7089 (N_7089,N_4210,N_3193);
nand U7090 (N_7090,N_4192,N_4757);
and U7091 (N_7091,N_2695,N_3962);
nand U7092 (N_7092,N_3038,N_4072);
or U7093 (N_7093,N_4285,N_2993);
nor U7094 (N_7094,N_4307,N_3011);
nor U7095 (N_7095,N_4855,N_4747);
nand U7096 (N_7096,N_4574,N_4457);
or U7097 (N_7097,N_4861,N_4044);
or U7098 (N_7098,N_2916,N_4705);
nand U7099 (N_7099,N_3713,N_4929);
or U7100 (N_7100,N_3182,N_3223);
or U7101 (N_7101,N_4956,N_4442);
or U7102 (N_7102,N_4160,N_4028);
or U7103 (N_7103,N_2938,N_3391);
or U7104 (N_7104,N_3790,N_3924);
nand U7105 (N_7105,N_4172,N_3896);
nor U7106 (N_7106,N_3433,N_3018);
or U7107 (N_7107,N_4767,N_3511);
or U7108 (N_7108,N_2671,N_4864);
or U7109 (N_7109,N_2701,N_3416);
nand U7110 (N_7110,N_3326,N_3590);
nand U7111 (N_7111,N_3236,N_3096);
nand U7112 (N_7112,N_3904,N_4948);
or U7113 (N_7113,N_2802,N_4537);
and U7114 (N_7114,N_4221,N_4731);
nand U7115 (N_7115,N_4354,N_4568);
and U7116 (N_7116,N_2814,N_4739);
or U7117 (N_7117,N_4204,N_4793);
or U7118 (N_7118,N_3285,N_2997);
nand U7119 (N_7119,N_4327,N_2605);
nor U7120 (N_7120,N_2950,N_2856);
or U7121 (N_7121,N_3183,N_4708);
or U7122 (N_7122,N_2548,N_3423);
or U7123 (N_7123,N_4699,N_2881);
nor U7124 (N_7124,N_2511,N_2897);
and U7125 (N_7125,N_2554,N_3362);
and U7126 (N_7126,N_4727,N_3349);
nor U7127 (N_7127,N_4194,N_4270);
nand U7128 (N_7128,N_3853,N_4382);
nand U7129 (N_7129,N_3448,N_4619);
xor U7130 (N_7130,N_3908,N_3108);
nor U7131 (N_7131,N_3216,N_4342);
nor U7132 (N_7132,N_4726,N_4073);
nand U7133 (N_7133,N_4209,N_4433);
or U7134 (N_7134,N_3101,N_4835);
nand U7135 (N_7135,N_4349,N_4570);
and U7136 (N_7136,N_4942,N_3680);
and U7137 (N_7137,N_4095,N_3659);
nand U7138 (N_7138,N_3769,N_3852);
nor U7139 (N_7139,N_3836,N_4931);
and U7140 (N_7140,N_3346,N_4203);
nor U7141 (N_7141,N_3998,N_4560);
or U7142 (N_7142,N_3093,N_4956);
nor U7143 (N_7143,N_4341,N_3111);
and U7144 (N_7144,N_4376,N_4087);
nor U7145 (N_7145,N_3860,N_2716);
or U7146 (N_7146,N_2743,N_4053);
nand U7147 (N_7147,N_3839,N_3406);
nor U7148 (N_7148,N_2594,N_3011);
and U7149 (N_7149,N_4315,N_3047);
nor U7150 (N_7150,N_3990,N_4165);
nand U7151 (N_7151,N_4326,N_3124);
and U7152 (N_7152,N_4191,N_3720);
and U7153 (N_7153,N_3615,N_3939);
nand U7154 (N_7154,N_4264,N_4752);
nand U7155 (N_7155,N_3081,N_4614);
and U7156 (N_7156,N_3752,N_4058);
and U7157 (N_7157,N_3839,N_3904);
nor U7158 (N_7158,N_4138,N_4106);
nor U7159 (N_7159,N_2636,N_3593);
or U7160 (N_7160,N_3741,N_3631);
nor U7161 (N_7161,N_3525,N_4960);
or U7162 (N_7162,N_4092,N_3897);
and U7163 (N_7163,N_4193,N_4225);
or U7164 (N_7164,N_4675,N_4799);
nor U7165 (N_7165,N_3736,N_4053);
nor U7166 (N_7166,N_3286,N_4265);
nand U7167 (N_7167,N_3212,N_3825);
nand U7168 (N_7168,N_4492,N_2982);
nor U7169 (N_7169,N_4147,N_3023);
nand U7170 (N_7170,N_4493,N_4559);
nand U7171 (N_7171,N_3605,N_3280);
nand U7172 (N_7172,N_4883,N_4463);
nor U7173 (N_7173,N_4464,N_3155);
nor U7174 (N_7174,N_3508,N_4681);
or U7175 (N_7175,N_4415,N_3078);
or U7176 (N_7176,N_3105,N_4431);
or U7177 (N_7177,N_3615,N_3252);
and U7178 (N_7178,N_3798,N_2925);
nand U7179 (N_7179,N_3512,N_4787);
and U7180 (N_7180,N_4765,N_3385);
nor U7181 (N_7181,N_3342,N_4491);
nor U7182 (N_7182,N_3663,N_3465);
nor U7183 (N_7183,N_2891,N_3088);
and U7184 (N_7184,N_4996,N_3525);
nand U7185 (N_7185,N_3582,N_4954);
xnor U7186 (N_7186,N_4267,N_4037);
nand U7187 (N_7187,N_3319,N_2993);
and U7188 (N_7188,N_3584,N_4028);
nand U7189 (N_7189,N_3594,N_3554);
nor U7190 (N_7190,N_2563,N_4714);
and U7191 (N_7191,N_2565,N_2875);
nand U7192 (N_7192,N_3876,N_2951);
nand U7193 (N_7193,N_4541,N_4575);
nand U7194 (N_7194,N_4567,N_4574);
or U7195 (N_7195,N_4296,N_4432);
nand U7196 (N_7196,N_3414,N_2717);
nand U7197 (N_7197,N_3257,N_3325);
nand U7198 (N_7198,N_4263,N_4481);
or U7199 (N_7199,N_4687,N_4039);
and U7200 (N_7200,N_4473,N_4289);
nor U7201 (N_7201,N_2589,N_2505);
or U7202 (N_7202,N_3267,N_4517);
and U7203 (N_7203,N_3041,N_4084);
nand U7204 (N_7204,N_4332,N_3674);
or U7205 (N_7205,N_4848,N_3307);
nand U7206 (N_7206,N_4065,N_4620);
nor U7207 (N_7207,N_3925,N_2539);
or U7208 (N_7208,N_2983,N_2896);
or U7209 (N_7209,N_2807,N_3917);
nand U7210 (N_7210,N_3457,N_3931);
and U7211 (N_7211,N_2574,N_2864);
or U7212 (N_7212,N_3727,N_3509);
or U7213 (N_7213,N_4820,N_4133);
and U7214 (N_7214,N_4091,N_3781);
nand U7215 (N_7215,N_3640,N_2899);
nand U7216 (N_7216,N_3903,N_4030);
and U7217 (N_7217,N_3112,N_2522);
and U7218 (N_7218,N_4034,N_4384);
and U7219 (N_7219,N_2604,N_4749);
or U7220 (N_7220,N_3557,N_3697);
nand U7221 (N_7221,N_2937,N_4897);
or U7222 (N_7222,N_2625,N_2831);
xnor U7223 (N_7223,N_4615,N_2651);
nor U7224 (N_7224,N_3975,N_3231);
and U7225 (N_7225,N_4947,N_3831);
and U7226 (N_7226,N_4827,N_2739);
nand U7227 (N_7227,N_3875,N_3675);
nor U7228 (N_7228,N_3033,N_4588);
nand U7229 (N_7229,N_4523,N_2728);
or U7230 (N_7230,N_3458,N_3706);
and U7231 (N_7231,N_2575,N_4395);
nor U7232 (N_7232,N_4694,N_4184);
xor U7233 (N_7233,N_4232,N_3141);
and U7234 (N_7234,N_4056,N_4329);
nand U7235 (N_7235,N_3568,N_3944);
nor U7236 (N_7236,N_3934,N_3477);
or U7237 (N_7237,N_2720,N_2984);
nor U7238 (N_7238,N_3675,N_3404);
nor U7239 (N_7239,N_4285,N_2686);
nor U7240 (N_7240,N_2872,N_3183);
or U7241 (N_7241,N_3901,N_2888);
nand U7242 (N_7242,N_4795,N_2937);
or U7243 (N_7243,N_4921,N_3720);
and U7244 (N_7244,N_3146,N_2991);
and U7245 (N_7245,N_3137,N_4763);
or U7246 (N_7246,N_3052,N_3615);
nor U7247 (N_7247,N_3337,N_4946);
and U7248 (N_7248,N_2568,N_4749);
nor U7249 (N_7249,N_3217,N_4211);
or U7250 (N_7250,N_4381,N_4067);
xnor U7251 (N_7251,N_4305,N_4033);
or U7252 (N_7252,N_3657,N_4086);
nand U7253 (N_7253,N_4589,N_4917);
and U7254 (N_7254,N_3175,N_2746);
or U7255 (N_7255,N_3995,N_4656);
or U7256 (N_7256,N_2711,N_3380);
nor U7257 (N_7257,N_2746,N_3786);
and U7258 (N_7258,N_4215,N_3584);
and U7259 (N_7259,N_4156,N_2904);
nor U7260 (N_7260,N_2661,N_3576);
nand U7261 (N_7261,N_3921,N_2811);
or U7262 (N_7262,N_4680,N_4183);
nor U7263 (N_7263,N_2585,N_3724);
and U7264 (N_7264,N_3738,N_3172);
and U7265 (N_7265,N_4580,N_3542);
nand U7266 (N_7266,N_2681,N_4709);
and U7267 (N_7267,N_4724,N_4688);
nor U7268 (N_7268,N_2713,N_3987);
or U7269 (N_7269,N_4229,N_3063);
nor U7270 (N_7270,N_3089,N_3809);
nand U7271 (N_7271,N_3220,N_4237);
nor U7272 (N_7272,N_2760,N_2666);
and U7273 (N_7273,N_4044,N_3280);
and U7274 (N_7274,N_4309,N_3377);
or U7275 (N_7275,N_4312,N_4661);
nand U7276 (N_7276,N_3399,N_2729);
nor U7277 (N_7277,N_3525,N_2726);
nand U7278 (N_7278,N_4831,N_3920);
or U7279 (N_7279,N_3411,N_3508);
and U7280 (N_7280,N_4745,N_3974);
nand U7281 (N_7281,N_4606,N_4307);
nor U7282 (N_7282,N_3187,N_3942);
xnor U7283 (N_7283,N_4843,N_3399);
and U7284 (N_7284,N_4518,N_3893);
or U7285 (N_7285,N_4360,N_2735);
nand U7286 (N_7286,N_3258,N_3060);
nor U7287 (N_7287,N_4558,N_4007);
and U7288 (N_7288,N_4182,N_2716);
nand U7289 (N_7289,N_3613,N_2719);
and U7290 (N_7290,N_3830,N_3560);
nand U7291 (N_7291,N_3541,N_4574);
and U7292 (N_7292,N_3585,N_3507);
nor U7293 (N_7293,N_4966,N_2911);
nand U7294 (N_7294,N_4008,N_3394);
and U7295 (N_7295,N_2697,N_2645);
and U7296 (N_7296,N_4339,N_3870);
nand U7297 (N_7297,N_3419,N_2777);
and U7298 (N_7298,N_4007,N_4651);
and U7299 (N_7299,N_4929,N_4515);
or U7300 (N_7300,N_3328,N_4126);
or U7301 (N_7301,N_3974,N_4530);
nand U7302 (N_7302,N_3552,N_3650);
or U7303 (N_7303,N_3179,N_3743);
nand U7304 (N_7304,N_3594,N_4796);
or U7305 (N_7305,N_2822,N_3261);
nor U7306 (N_7306,N_2851,N_4767);
and U7307 (N_7307,N_3874,N_4287);
and U7308 (N_7308,N_3302,N_3767);
nor U7309 (N_7309,N_3315,N_3934);
nand U7310 (N_7310,N_3248,N_4833);
nand U7311 (N_7311,N_2713,N_4083);
and U7312 (N_7312,N_3814,N_3907);
and U7313 (N_7313,N_3633,N_4755);
or U7314 (N_7314,N_2561,N_4746);
and U7315 (N_7315,N_3033,N_4737);
nor U7316 (N_7316,N_2635,N_2551);
nor U7317 (N_7317,N_4775,N_3466);
and U7318 (N_7318,N_2776,N_3895);
or U7319 (N_7319,N_3092,N_3473);
nand U7320 (N_7320,N_4451,N_4631);
nand U7321 (N_7321,N_4451,N_4464);
and U7322 (N_7322,N_3588,N_3215);
or U7323 (N_7323,N_4164,N_3057);
or U7324 (N_7324,N_3230,N_2621);
or U7325 (N_7325,N_4926,N_2517);
or U7326 (N_7326,N_4577,N_2758);
or U7327 (N_7327,N_4886,N_4295);
and U7328 (N_7328,N_4585,N_2910);
and U7329 (N_7329,N_3960,N_3033);
nand U7330 (N_7330,N_4808,N_2652);
nor U7331 (N_7331,N_3792,N_4134);
or U7332 (N_7332,N_2808,N_3795);
nor U7333 (N_7333,N_4393,N_3849);
and U7334 (N_7334,N_4065,N_4551);
nor U7335 (N_7335,N_2792,N_4401);
or U7336 (N_7336,N_3444,N_2637);
and U7337 (N_7337,N_2794,N_3080);
nor U7338 (N_7338,N_3234,N_3474);
nand U7339 (N_7339,N_4730,N_4433);
or U7340 (N_7340,N_3841,N_3703);
nor U7341 (N_7341,N_3316,N_4097);
nor U7342 (N_7342,N_3816,N_3059);
nor U7343 (N_7343,N_4028,N_4667);
and U7344 (N_7344,N_3873,N_3900);
or U7345 (N_7345,N_4814,N_2880);
and U7346 (N_7346,N_4529,N_4007);
and U7347 (N_7347,N_2967,N_3769);
and U7348 (N_7348,N_2796,N_3611);
and U7349 (N_7349,N_4407,N_3234);
nor U7350 (N_7350,N_4459,N_4904);
and U7351 (N_7351,N_2883,N_4817);
nand U7352 (N_7352,N_2699,N_4112);
nor U7353 (N_7353,N_3713,N_3991);
or U7354 (N_7354,N_2860,N_3898);
and U7355 (N_7355,N_4623,N_3496);
or U7356 (N_7356,N_2927,N_4657);
nor U7357 (N_7357,N_2568,N_3361);
or U7358 (N_7358,N_2726,N_4374);
nor U7359 (N_7359,N_4443,N_4731);
xor U7360 (N_7360,N_2782,N_3211);
nor U7361 (N_7361,N_4771,N_2974);
or U7362 (N_7362,N_4297,N_4275);
or U7363 (N_7363,N_4444,N_2810);
nand U7364 (N_7364,N_2953,N_4793);
nor U7365 (N_7365,N_3139,N_3149);
and U7366 (N_7366,N_3933,N_4785);
and U7367 (N_7367,N_2552,N_3297);
nand U7368 (N_7368,N_4773,N_2633);
or U7369 (N_7369,N_3845,N_4473);
nand U7370 (N_7370,N_4886,N_4597);
nand U7371 (N_7371,N_3161,N_3798);
or U7372 (N_7372,N_4427,N_4541);
nor U7373 (N_7373,N_4882,N_3990);
or U7374 (N_7374,N_3055,N_4676);
or U7375 (N_7375,N_3981,N_3327);
nand U7376 (N_7376,N_3473,N_3024);
and U7377 (N_7377,N_3958,N_4646);
nand U7378 (N_7378,N_2614,N_4120);
and U7379 (N_7379,N_4352,N_2679);
nor U7380 (N_7380,N_4971,N_3397);
and U7381 (N_7381,N_3275,N_4094);
and U7382 (N_7382,N_3689,N_3380);
nand U7383 (N_7383,N_4657,N_3369);
nor U7384 (N_7384,N_3002,N_4628);
nor U7385 (N_7385,N_3894,N_2700);
or U7386 (N_7386,N_3916,N_4087);
nand U7387 (N_7387,N_4665,N_2738);
nor U7388 (N_7388,N_2863,N_3719);
and U7389 (N_7389,N_3671,N_3146);
nand U7390 (N_7390,N_4029,N_4316);
and U7391 (N_7391,N_4513,N_2787);
and U7392 (N_7392,N_3519,N_3457);
or U7393 (N_7393,N_2631,N_2976);
nand U7394 (N_7394,N_3425,N_3593);
nand U7395 (N_7395,N_4214,N_4824);
nor U7396 (N_7396,N_4564,N_2566);
and U7397 (N_7397,N_2920,N_3657);
and U7398 (N_7398,N_4545,N_3209);
nand U7399 (N_7399,N_2803,N_3363);
nor U7400 (N_7400,N_3993,N_2744);
and U7401 (N_7401,N_3091,N_3006);
or U7402 (N_7402,N_3984,N_4001);
or U7403 (N_7403,N_3479,N_3577);
or U7404 (N_7404,N_2671,N_4869);
or U7405 (N_7405,N_3495,N_3976);
or U7406 (N_7406,N_4626,N_2786);
and U7407 (N_7407,N_3291,N_3404);
nand U7408 (N_7408,N_2850,N_3180);
nand U7409 (N_7409,N_2878,N_3055);
or U7410 (N_7410,N_2708,N_2560);
nand U7411 (N_7411,N_4798,N_3775);
and U7412 (N_7412,N_4400,N_3457);
nand U7413 (N_7413,N_2764,N_4053);
or U7414 (N_7414,N_2554,N_4867);
or U7415 (N_7415,N_4290,N_4033);
or U7416 (N_7416,N_3609,N_3848);
or U7417 (N_7417,N_3379,N_2596);
and U7418 (N_7418,N_4355,N_2851);
nor U7419 (N_7419,N_4208,N_2604);
and U7420 (N_7420,N_3672,N_2982);
or U7421 (N_7421,N_3581,N_4997);
and U7422 (N_7422,N_3127,N_2767);
and U7423 (N_7423,N_3577,N_3247);
nand U7424 (N_7424,N_3196,N_2703);
nor U7425 (N_7425,N_4645,N_4754);
nand U7426 (N_7426,N_4949,N_3622);
nand U7427 (N_7427,N_3976,N_4493);
and U7428 (N_7428,N_4042,N_2558);
or U7429 (N_7429,N_3364,N_3580);
and U7430 (N_7430,N_2600,N_3545);
nand U7431 (N_7431,N_3686,N_4779);
or U7432 (N_7432,N_4932,N_4553);
nor U7433 (N_7433,N_3617,N_4675);
and U7434 (N_7434,N_3711,N_3250);
or U7435 (N_7435,N_4697,N_3192);
and U7436 (N_7436,N_3924,N_3761);
and U7437 (N_7437,N_4419,N_3639);
or U7438 (N_7438,N_4037,N_4597);
and U7439 (N_7439,N_3190,N_4645);
and U7440 (N_7440,N_3147,N_4839);
or U7441 (N_7441,N_2835,N_2911);
nor U7442 (N_7442,N_4612,N_3094);
and U7443 (N_7443,N_2529,N_2766);
or U7444 (N_7444,N_2991,N_2940);
nor U7445 (N_7445,N_3117,N_2813);
nor U7446 (N_7446,N_3164,N_4747);
or U7447 (N_7447,N_3424,N_4099);
nand U7448 (N_7448,N_4310,N_3287);
or U7449 (N_7449,N_4341,N_4452);
nand U7450 (N_7450,N_4522,N_4341);
nand U7451 (N_7451,N_4759,N_2576);
and U7452 (N_7452,N_4816,N_2514);
or U7453 (N_7453,N_3347,N_4863);
and U7454 (N_7454,N_4093,N_4978);
xor U7455 (N_7455,N_4983,N_4004);
nand U7456 (N_7456,N_4220,N_3709);
and U7457 (N_7457,N_3789,N_4462);
or U7458 (N_7458,N_4341,N_3854);
or U7459 (N_7459,N_3550,N_3725);
nor U7460 (N_7460,N_2907,N_4343);
xnor U7461 (N_7461,N_2793,N_4087);
or U7462 (N_7462,N_2689,N_2839);
nor U7463 (N_7463,N_3201,N_3458);
nor U7464 (N_7464,N_4984,N_4952);
and U7465 (N_7465,N_3953,N_3449);
nor U7466 (N_7466,N_4779,N_3620);
or U7467 (N_7467,N_3231,N_4595);
nor U7468 (N_7468,N_2515,N_3248);
or U7469 (N_7469,N_3785,N_4399);
nand U7470 (N_7470,N_3964,N_4463);
nand U7471 (N_7471,N_4801,N_3734);
nand U7472 (N_7472,N_4006,N_3940);
or U7473 (N_7473,N_4266,N_4227);
nor U7474 (N_7474,N_3901,N_3960);
nor U7475 (N_7475,N_4852,N_3879);
nor U7476 (N_7476,N_4128,N_3177);
nor U7477 (N_7477,N_3233,N_3812);
and U7478 (N_7478,N_4094,N_3281);
nor U7479 (N_7479,N_3553,N_4058);
nor U7480 (N_7480,N_4484,N_4094);
nand U7481 (N_7481,N_3257,N_2637);
or U7482 (N_7482,N_3975,N_2534);
or U7483 (N_7483,N_4261,N_3352);
and U7484 (N_7484,N_3550,N_4448);
or U7485 (N_7485,N_3926,N_4537);
nand U7486 (N_7486,N_4089,N_3148);
nand U7487 (N_7487,N_4890,N_4442);
or U7488 (N_7488,N_4212,N_3162);
nor U7489 (N_7489,N_4612,N_4687);
nor U7490 (N_7490,N_4359,N_4706);
and U7491 (N_7491,N_4677,N_3953);
or U7492 (N_7492,N_4085,N_4437);
nor U7493 (N_7493,N_2673,N_4991);
and U7494 (N_7494,N_4029,N_4962);
nand U7495 (N_7495,N_2589,N_3160);
nand U7496 (N_7496,N_2681,N_4153);
nor U7497 (N_7497,N_3697,N_4061);
nor U7498 (N_7498,N_3238,N_4169);
nand U7499 (N_7499,N_3922,N_3128);
and U7500 (N_7500,N_5298,N_5187);
nor U7501 (N_7501,N_6223,N_5361);
and U7502 (N_7502,N_6300,N_5348);
and U7503 (N_7503,N_6461,N_5838);
and U7504 (N_7504,N_6032,N_5626);
nor U7505 (N_7505,N_6417,N_6192);
and U7506 (N_7506,N_6506,N_6212);
and U7507 (N_7507,N_7403,N_6985);
nor U7508 (N_7508,N_5953,N_7209);
nor U7509 (N_7509,N_5273,N_7174);
or U7510 (N_7510,N_5146,N_5745);
and U7511 (N_7511,N_6130,N_5400);
nor U7512 (N_7512,N_6099,N_7217);
nor U7513 (N_7513,N_6518,N_7289);
or U7514 (N_7514,N_6471,N_5657);
nor U7515 (N_7515,N_7142,N_6284);
and U7516 (N_7516,N_5384,N_5342);
or U7517 (N_7517,N_6356,N_6537);
nor U7518 (N_7518,N_7083,N_7230);
nor U7519 (N_7519,N_5917,N_7367);
nor U7520 (N_7520,N_5019,N_6475);
and U7521 (N_7521,N_5508,N_5649);
and U7522 (N_7522,N_5924,N_7244);
nand U7523 (N_7523,N_5392,N_6462);
and U7524 (N_7524,N_5863,N_5344);
nand U7525 (N_7525,N_5164,N_6813);
nor U7526 (N_7526,N_5589,N_6433);
or U7527 (N_7527,N_5394,N_6538);
or U7528 (N_7528,N_5159,N_5484);
nand U7529 (N_7529,N_5189,N_5637);
nor U7530 (N_7530,N_6432,N_5223);
or U7531 (N_7531,N_7489,N_6159);
nor U7532 (N_7532,N_6112,N_6310);
nor U7533 (N_7533,N_6986,N_7307);
and U7534 (N_7534,N_6663,N_7498);
or U7535 (N_7535,N_7013,N_6407);
nor U7536 (N_7536,N_5270,N_5612);
or U7537 (N_7537,N_6157,N_6258);
nor U7538 (N_7538,N_6085,N_6783);
nand U7539 (N_7539,N_7363,N_5524);
nor U7540 (N_7540,N_6853,N_6153);
nor U7541 (N_7541,N_6716,N_5870);
nand U7542 (N_7542,N_7253,N_5422);
and U7543 (N_7543,N_6001,N_5582);
or U7544 (N_7544,N_6394,N_6785);
and U7545 (N_7545,N_5389,N_5831);
or U7546 (N_7546,N_7195,N_5122);
nand U7547 (N_7547,N_6147,N_5026);
nor U7548 (N_7548,N_5502,N_5190);
or U7549 (N_7549,N_7308,N_5480);
nor U7550 (N_7550,N_6060,N_6763);
or U7551 (N_7551,N_5575,N_6013);
or U7552 (N_7552,N_7491,N_5212);
and U7553 (N_7553,N_5101,N_5677);
and U7554 (N_7554,N_6167,N_5903);
or U7555 (N_7555,N_6599,N_6464);
and U7556 (N_7556,N_6844,N_6372);
nand U7557 (N_7557,N_6224,N_5089);
nand U7558 (N_7558,N_6245,N_6272);
nor U7559 (N_7559,N_6875,N_6023);
nor U7560 (N_7560,N_6609,N_7279);
or U7561 (N_7561,N_6279,N_7214);
and U7562 (N_7562,N_6103,N_5888);
nor U7563 (N_7563,N_6846,N_5535);
and U7564 (N_7564,N_5143,N_6689);
nor U7565 (N_7565,N_5209,N_7292);
or U7566 (N_7566,N_7300,N_5703);
nor U7567 (N_7567,N_5965,N_6122);
and U7568 (N_7568,N_6132,N_6522);
and U7569 (N_7569,N_5641,N_5009);
nand U7570 (N_7570,N_6244,N_6362);
nand U7571 (N_7571,N_7290,N_5331);
or U7572 (N_7572,N_6751,N_5606);
nor U7573 (N_7573,N_7486,N_5285);
and U7574 (N_7574,N_5198,N_5148);
or U7575 (N_7575,N_5109,N_6139);
nand U7576 (N_7576,N_5036,N_7313);
or U7577 (N_7577,N_7444,N_5142);
and U7578 (N_7578,N_6250,N_5256);
and U7579 (N_7579,N_5015,N_5245);
nand U7580 (N_7580,N_5987,N_5121);
or U7581 (N_7581,N_5224,N_6830);
nand U7582 (N_7582,N_6927,N_5861);
or U7583 (N_7583,N_7454,N_6347);
or U7584 (N_7584,N_5216,N_5437);
nor U7585 (N_7585,N_5634,N_6893);
nor U7586 (N_7586,N_5200,N_5260);
and U7587 (N_7587,N_6852,N_6177);
nand U7588 (N_7588,N_7457,N_7228);
nor U7589 (N_7589,N_5062,N_7275);
nor U7590 (N_7590,N_5961,N_5787);
nor U7591 (N_7591,N_6924,N_6113);
or U7592 (N_7592,N_7051,N_6694);
or U7593 (N_7593,N_5719,N_6942);
or U7594 (N_7594,N_5968,N_6227);
and U7595 (N_7595,N_7069,N_5429);
and U7596 (N_7596,N_7438,N_7483);
or U7597 (N_7597,N_6596,N_6827);
or U7598 (N_7598,N_5774,N_6190);
and U7599 (N_7599,N_7286,N_5459);
xnor U7600 (N_7600,N_6009,N_7476);
or U7601 (N_7601,N_6217,N_6042);
or U7602 (N_7602,N_5059,N_6088);
and U7603 (N_7603,N_7001,N_6717);
or U7604 (N_7604,N_5057,N_6275);
or U7605 (N_7605,N_5470,N_6077);
nand U7606 (N_7606,N_5145,N_6724);
nor U7607 (N_7607,N_7448,N_5016);
and U7608 (N_7608,N_6532,N_5333);
nor U7609 (N_7609,N_5230,N_6326);
nand U7610 (N_7610,N_5586,N_5613);
nor U7611 (N_7611,N_5085,N_6990);
nand U7612 (N_7612,N_7162,N_6068);
nor U7613 (N_7613,N_6184,N_5744);
and U7614 (N_7614,N_7196,N_5050);
nor U7615 (N_7615,N_7095,N_7257);
and U7616 (N_7616,N_5826,N_5288);
nor U7617 (N_7617,N_5199,N_7254);
or U7618 (N_7618,N_5287,N_6090);
or U7619 (N_7619,N_5785,N_5386);
nand U7620 (N_7620,N_6735,N_6592);
and U7621 (N_7621,N_7382,N_7059);
and U7622 (N_7622,N_7299,N_5832);
nor U7623 (N_7623,N_5654,N_7144);
and U7624 (N_7624,N_6114,N_7213);
and U7625 (N_7625,N_5934,N_6624);
nor U7626 (N_7626,N_6011,N_6989);
or U7627 (N_7627,N_7391,N_5042);
and U7628 (N_7628,N_6238,N_5413);
nand U7629 (N_7629,N_5184,N_6470);
nor U7630 (N_7630,N_5952,N_5229);
nand U7631 (N_7631,N_6836,N_6381);
and U7632 (N_7632,N_7317,N_5000);
and U7633 (N_7633,N_6151,N_6405);
nor U7634 (N_7634,N_6080,N_6962);
or U7635 (N_7635,N_6949,N_5607);
and U7636 (N_7636,N_6947,N_6648);
and U7637 (N_7637,N_6704,N_5995);
nor U7638 (N_7638,N_6858,N_6298);
and U7639 (N_7639,N_7028,N_5897);
or U7640 (N_7640,N_7376,N_5060);
nor U7641 (N_7641,N_6792,N_6322);
and U7642 (N_7642,N_6698,N_6692);
nor U7643 (N_7643,N_5500,N_5098);
and U7644 (N_7644,N_5091,N_5969);
or U7645 (N_7645,N_5963,N_6329);
nand U7646 (N_7646,N_6303,N_5249);
nand U7647 (N_7647,N_5672,N_5879);
nor U7648 (N_7648,N_5100,N_5168);
nor U7649 (N_7649,N_5329,N_5355);
nand U7650 (N_7650,N_7060,N_6014);
and U7651 (N_7651,N_5241,N_6096);
nor U7652 (N_7652,N_5882,N_6387);
or U7653 (N_7653,N_5381,N_6026);
nand U7654 (N_7654,N_6973,N_6677);
nand U7655 (N_7655,N_6832,N_6831);
or U7656 (N_7656,N_6268,N_6450);
nor U7657 (N_7657,N_5681,N_7251);
nor U7658 (N_7658,N_5156,N_5173);
and U7659 (N_7659,N_6489,N_6350);
nand U7660 (N_7660,N_7291,N_6739);
nand U7661 (N_7661,N_5950,N_5372);
nand U7662 (N_7662,N_6640,N_7232);
and U7663 (N_7663,N_7461,N_5578);
nand U7664 (N_7664,N_7080,N_7357);
and U7665 (N_7665,N_7185,N_7139);
nor U7666 (N_7666,N_5306,N_6436);
xnor U7667 (N_7667,N_6109,N_6550);
nor U7668 (N_7668,N_5728,N_5957);
nor U7669 (N_7669,N_7480,N_6528);
nor U7670 (N_7670,N_7406,N_5892);
and U7671 (N_7671,N_6938,N_5583);
nand U7672 (N_7672,N_5880,N_6286);
nand U7673 (N_7673,N_7356,N_6176);
and U7674 (N_7674,N_5814,N_6590);
or U7675 (N_7675,N_6168,N_6043);
nor U7676 (N_7676,N_6871,N_5345);
nand U7677 (N_7677,N_6507,N_5635);
or U7678 (N_7678,N_5175,N_5850);
nand U7679 (N_7679,N_6841,N_6004);
and U7680 (N_7680,N_7204,N_5176);
or U7681 (N_7681,N_6806,N_6292);
and U7682 (N_7682,N_5061,N_6261);
and U7683 (N_7683,N_6822,N_6969);
nor U7684 (N_7684,N_5802,N_7346);
nor U7685 (N_7685,N_7085,N_5558);
xor U7686 (N_7686,N_5662,N_7425);
nand U7687 (N_7687,N_5149,N_7163);
nor U7688 (N_7688,N_6800,N_7442);
nor U7689 (N_7689,N_7038,N_5399);
nand U7690 (N_7690,N_5781,N_6788);
nand U7691 (N_7691,N_7122,N_5035);
xor U7692 (N_7692,N_5926,N_5485);
nor U7693 (N_7693,N_6944,N_5736);
or U7694 (N_7694,N_6236,N_5325);
nor U7695 (N_7695,N_6161,N_7485);
nor U7696 (N_7696,N_5792,N_5281);
and U7697 (N_7697,N_5691,N_5408);
nand U7698 (N_7698,N_6263,N_7295);
nand U7699 (N_7699,N_6600,N_5999);
nor U7700 (N_7700,N_6709,N_7034);
or U7701 (N_7701,N_5630,N_5130);
or U7702 (N_7702,N_6733,N_6943);
nand U7703 (N_7703,N_7337,N_5871);
nand U7704 (N_7704,N_5817,N_6373);
and U7705 (N_7705,N_6655,N_7110);
and U7706 (N_7706,N_5570,N_5152);
and U7707 (N_7707,N_6102,N_7200);
and U7708 (N_7708,N_6910,N_5320);
or U7709 (N_7709,N_5810,N_7130);
or U7710 (N_7710,N_7258,N_7184);
nand U7711 (N_7711,N_6481,N_6512);
nand U7712 (N_7712,N_6406,N_5929);
and U7713 (N_7713,N_6578,N_6273);
or U7714 (N_7714,N_6583,N_6234);
or U7715 (N_7715,N_6000,N_5797);
nor U7716 (N_7716,N_7137,N_5935);
nor U7717 (N_7717,N_5137,N_7424);
and U7718 (N_7718,N_5805,N_5076);
or U7719 (N_7719,N_5599,N_6547);
nand U7720 (N_7720,N_5279,N_5192);
nand U7721 (N_7721,N_7261,N_6597);
nor U7722 (N_7722,N_7041,N_5705);
or U7723 (N_7723,N_5778,N_6270);
nand U7724 (N_7724,N_6045,N_6657);
nand U7725 (N_7725,N_7183,N_5180);
nand U7726 (N_7726,N_6131,N_6777);
nand U7727 (N_7727,N_7349,N_5460);
nor U7728 (N_7728,N_7125,N_5232);
and U7729 (N_7729,N_6363,N_5701);
nand U7730 (N_7730,N_5752,N_5017);
and U7731 (N_7731,N_5486,N_6423);
and U7732 (N_7732,N_5310,N_5828);
nand U7733 (N_7733,N_6584,N_5576);
nor U7734 (N_7734,N_5794,N_5954);
or U7735 (N_7735,N_5020,N_6497);
nor U7736 (N_7736,N_6683,N_5509);
and U7737 (N_7737,N_5825,N_6357);
and U7738 (N_7738,N_6977,N_7000);
or U7739 (N_7739,N_6517,N_5960);
or U7740 (N_7740,N_5990,N_6937);
and U7741 (N_7741,N_5088,N_7282);
and U7742 (N_7742,N_5025,N_5276);
nand U7743 (N_7743,N_5131,N_7381);
nor U7744 (N_7744,N_5956,N_6815);
nor U7745 (N_7745,N_6883,N_5154);
or U7746 (N_7746,N_6759,N_6178);
and U7747 (N_7747,N_7365,N_5418);
nor U7748 (N_7748,N_5447,N_5491);
or U7749 (N_7749,N_5056,N_7255);
and U7750 (N_7750,N_6616,N_6757);
nor U7751 (N_7751,N_5003,N_6542);
nand U7752 (N_7752,N_6679,N_7098);
nor U7753 (N_7753,N_6642,N_6029);
or U7754 (N_7754,N_6035,N_6498);
xor U7755 (N_7755,N_5448,N_5660);
nand U7756 (N_7756,N_6867,N_5067);
nor U7757 (N_7757,N_6331,N_7373);
and U7758 (N_7758,N_5193,N_6059);
nor U7759 (N_7759,N_6401,N_6220);
nand U7760 (N_7760,N_5018,N_5445);
and U7761 (N_7761,N_6144,N_6825);
nand U7762 (N_7762,N_7383,N_6368);
nor U7763 (N_7763,N_6074,N_5207);
nand U7764 (N_7764,N_6249,N_5989);
or U7765 (N_7765,N_5678,N_6732);
nand U7766 (N_7766,N_6050,N_5138);
nor U7767 (N_7767,N_6315,N_6037);
nor U7768 (N_7768,N_5114,N_6749);
nor U7769 (N_7769,N_7327,N_6824);
and U7770 (N_7770,N_7118,N_5706);
or U7771 (N_7771,N_5166,N_5770);
xnor U7772 (N_7772,N_5103,N_5258);
and U7773 (N_7773,N_5412,N_5697);
nor U7774 (N_7774,N_7149,N_7108);
nor U7775 (N_7775,N_5640,N_6545);
and U7776 (N_7776,N_5527,N_6755);
nor U7777 (N_7777,N_7063,N_5219);
and U7778 (N_7778,N_6057,N_6115);
nor U7779 (N_7779,N_7435,N_7193);
nand U7780 (N_7780,N_6402,N_5682);
and U7781 (N_7781,N_5151,N_7322);
nor U7782 (N_7782,N_7011,N_5605);
nand U7783 (N_7783,N_5365,N_6848);
nor U7784 (N_7784,N_6997,N_7090);
or U7785 (N_7785,N_5405,N_5014);
nor U7786 (N_7786,N_5253,N_6073);
or U7787 (N_7787,N_6288,N_7102);
and U7788 (N_7788,N_6586,N_7301);
and U7789 (N_7789,N_5684,N_6750);
and U7790 (N_7790,N_7015,N_6995);
nor U7791 (N_7791,N_5799,N_7452);
and U7792 (N_7792,N_5272,N_6179);
xor U7793 (N_7793,N_5543,N_7283);
or U7794 (N_7794,N_5217,N_5622);
nor U7795 (N_7795,N_6772,N_6964);
or U7796 (N_7796,N_7328,N_5519);
or U7797 (N_7797,N_5139,N_5760);
or U7798 (N_7798,N_6793,N_6604);
nand U7799 (N_7799,N_6202,N_5598);
nor U7800 (N_7800,N_6911,N_6465);
nand U7801 (N_7801,N_6081,N_5443);
or U7802 (N_7802,N_7210,N_5722);
nand U7803 (N_7803,N_6649,N_6318);
nor U7804 (N_7804,N_7086,N_7023);
or U7805 (N_7805,N_5611,N_5140);
and U7806 (N_7806,N_6079,N_7114);
and U7807 (N_7807,N_6511,N_5473);
and U7808 (N_7808,N_6203,N_5743);
nor U7809 (N_7809,N_5402,N_5242);
nand U7810 (N_7810,N_5304,N_5767);
or U7811 (N_7811,N_7306,N_7248);
or U7812 (N_7812,N_5980,N_7032);
nor U7813 (N_7813,N_5975,N_7407);
or U7814 (N_7814,N_7293,N_7459);
nor U7815 (N_7815,N_5120,N_7351);
or U7816 (N_7816,N_5388,N_6534);
nor U7817 (N_7817,N_5510,N_6125);
nor U7818 (N_7818,N_6602,N_5280);
and U7819 (N_7819,N_6370,N_6909);
nand U7820 (N_7820,N_7467,N_6890);
nand U7821 (N_7821,N_5531,N_7026);
or U7822 (N_7822,N_7402,N_6908);
nand U7823 (N_7823,N_7004,N_5488);
nor U7824 (N_7824,N_7329,N_5074);
nand U7825 (N_7825,N_5360,N_7386);
nor U7826 (N_7826,N_6260,N_5983);
and U7827 (N_7827,N_5449,N_6941);
nor U7828 (N_7828,N_6865,N_5548);
nand U7829 (N_7829,N_5552,N_6054);
and U7830 (N_7830,N_6784,N_5064);
or U7831 (N_7831,N_7224,N_7115);
or U7832 (N_7832,N_6525,N_7318);
nor U7833 (N_7833,N_5727,N_5340);
or U7834 (N_7834,N_7159,N_5514);
and U7835 (N_7835,N_7408,N_5133);
nand U7836 (N_7836,N_7256,N_5228);
and U7837 (N_7837,N_5628,N_6371);
or U7838 (N_7838,N_6154,N_5704);
nand U7839 (N_7839,N_7138,N_5659);
and U7840 (N_7840,N_6209,N_5358);
and U7841 (N_7841,N_6119,N_5013);
nand U7842 (N_7842,N_7212,N_5186);
and U7843 (N_7843,N_7339,N_5962);
nor U7844 (N_7844,N_5761,N_7487);
and U7845 (N_7845,N_6175,N_6415);
nor U7846 (N_7846,N_5909,N_6888);
nand U7847 (N_7847,N_6299,N_6691);
nand U7848 (N_7848,N_5873,N_6838);
or U7849 (N_7849,N_7288,N_6182);
nand U7850 (N_7850,N_5658,N_7428);
nor U7851 (N_7851,N_5444,N_7462);
nor U7852 (N_7852,N_5900,N_5645);
nand U7853 (N_7853,N_6505,N_5927);
and U7854 (N_7854,N_7127,N_7415);
or U7855 (N_7855,N_6309,N_6862);
nor U7856 (N_7856,N_7113,N_5991);
and U7857 (N_7857,N_5574,N_5542);
nor U7858 (N_7858,N_6252,N_5433);
nor U7859 (N_7859,N_6451,N_5113);
nor U7860 (N_7860,N_6928,N_7397);
or U7861 (N_7861,N_5762,N_5820);
or U7862 (N_7862,N_6959,N_6398);
and U7863 (N_7863,N_5024,N_5604);
nor U7864 (N_7864,N_5308,N_7150);
and U7865 (N_7865,N_5438,N_6826);
or U7866 (N_7866,N_6473,N_7395);
or U7867 (N_7867,N_6064,N_7325);
and U7868 (N_7868,N_5419,N_7404);
or U7869 (N_7869,N_5373,N_5442);
and U7870 (N_7870,N_5674,N_5467);
and U7871 (N_7871,N_5522,N_7222);
xnor U7872 (N_7872,N_5461,N_6764);
and U7873 (N_7873,N_5702,N_6795);
nand U7874 (N_7874,N_7167,N_5239);
nor U7875 (N_7875,N_6774,N_6193);
xnor U7876 (N_7876,N_7284,N_5231);
nor U7877 (N_7877,N_6851,N_7020);
nor U7878 (N_7878,N_6934,N_7236);
nor U7879 (N_7879,N_6767,N_6577);
or U7880 (N_7880,N_5819,N_5849);
nand U7881 (N_7881,N_6442,N_5925);
or U7882 (N_7882,N_6926,N_5277);
nand U7883 (N_7883,N_5978,N_6998);
and U7884 (N_7884,N_7259,N_6880);
nor U7885 (N_7885,N_5809,N_7104);
or U7886 (N_7886,N_7111,N_6539);
nor U7887 (N_7887,N_6896,N_6654);
nor U7888 (N_7888,N_5343,N_5410);
nor U7889 (N_7889,N_6221,N_5299);
nand U7890 (N_7890,N_6726,N_5503);
nor U7891 (N_7891,N_5047,N_5922);
nand U7892 (N_7892,N_5994,N_7350);
nand U7893 (N_7893,N_7057,N_5763);
nor U7894 (N_7894,N_6705,N_5561);
or U7895 (N_7895,N_7450,N_5933);
nand U7896 (N_7896,N_6520,N_7268);
or U7897 (N_7897,N_5182,N_6095);
nand U7898 (N_7898,N_7099,N_6290);
nor U7899 (N_7899,N_7420,N_6920);
nand U7900 (N_7900,N_5789,N_5165);
nor U7901 (N_7901,N_5895,N_6982);
nand U7902 (N_7902,N_5685,N_5301);
nand U7903 (N_7903,N_5597,N_7134);
nand U7904 (N_7904,N_6984,N_6681);
nor U7905 (N_7905,N_6579,N_7199);
and U7906 (N_7906,N_5893,N_7394);
and U7907 (N_7907,N_6199,N_6603);
xnor U7908 (N_7908,N_6409,N_5843);
and U7909 (N_7909,N_5158,N_5981);
xor U7910 (N_7910,N_6819,N_6488);
and U7911 (N_7911,N_5387,N_5337);
nand U7912 (N_7912,N_6485,N_6173);
or U7913 (N_7913,N_5498,N_7310);
or U7914 (N_7914,N_5568,N_6866);
nand U7915 (N_7915,N_6058,N_6805);
nand U7916 (N_7916,N_6963,N_6491);
nand U7917 (N_7917,N_5124,N_6695);
nand U7918 (N_7918,N_5539,N_5615);
nand U7919 (N_7919,N_5305,N_5840);
and U7920 (N_7920,N_7148,N_6570);
nand U7921 (N_7921,N_7237,N_7492);
and U7922 (N_7922,N_6965,N_7338);
and U7923 (N_7923,N_5516,N_5087);
or U7924 (N_7924,N_6894,N_7323);
and U7925 (N_7925,N_6548,N_5716);
and U7926 (N_7926,N_6480,N_5243);
or U7927 (N_7927,N_6094,N_6515);
nor U7928 (N_7928,N_7445,N_6993);
nor U7929 (N_7929,N_6879,N_5772);
or U7930 (N_7930,N_6658,N_6226);
nand U7931 (N_7931,N_6946,N_6146);
nand U7932 (N_7932,N_6974,N_5110);
or U7933 (N_7933,N_5069,N_5608);
and U7934 (N_7934,N_5732,N_7008);
or U7935 (N_7935,N_5311,N_6377);
and U7936 (N_7936,N_6535,N_7100);
and U7937 (N_7937,N_5376,N_5711);
nand U7938 (N_7938,N_5816,N_5601);
and U7939 (N_7939,N_6421,N_6206);
or U7940 (N_7940,N_6917,N_6747);
and U7941 (N_7941,N_6593,N_6412);
and U7942 (N_7942,N_5153,N_5073);
nor U7943 (N_7943,N_6328,N_6834);
and U7944 (N_7944,N_6799,N_5247);
nand U7945 (N_7945,N_5887,N_5350);
nand U7946 (N_7946,N_7436,N_6435);
and U7947 (N_7947,N_6162,N_5593);
or U7948 (N_7948,N_5815,N_6664);
or U7949 (N_7949,N_7493,N_6697);
nand U7950 (N_7950,N_5300,N_7046);
or U7951 (N_7951,N_6495,N_7164);
or U7952 (N_7952,N_6383,N_6424);
nor U7953 (N_7953,N_5890,N_6960);
and U7954 (N_7954,N_5054,N_7387);
and U7955 (N_7955,N_5590,N_5618);
and U7956 (N_7956,N_6563,N_5097);
nand U7957 (N_7957,N_6891,N_7264);
or U7958 (N_7958,N_5665,N_6386);
nand U7959 (N_7959,N_7319,N_5906);
nor U7960 (N_7960,N_7481,N_7128);
nand U7961 (N_7961,N_6595,N_5988);
and U7962 (N_7962,N_6902,N_6195);
or U7963 (N_7963,N_6644,N_5855);
and U7964 (N_7964,N_6546,N_5913);
and U7965 (N_7965,N_5844,N_7215);
nor U7966 (N_7966,N_5157,N_6174);
and U7967 (N_7967,N_7355,N_5713);
nor U7968 (N_7968,N_5274,N_6181);
and U7969 (N_7969,N_7112,N_5915);
and U7970 (N_7970,N_5268,N_6140);
nor U7971 (N_7971,N_5937,N_6790);
nand U7972 (N_7972,N_6676,N_6005);
and U7973 (N_7973,N_6957,N_6359);
or U7974 (N_7974,N_5172,N_6900);
nor U7975 (N_7975,N_5380,N_7414);
or U7976 (N_7976,N_5595,N_6361);
xnor U7977 (N_7977,N_6991,N_6884);
and U7978 (N_7978,N_7281,N_5235);
or U7979 (N_7979,N_6466,N_5334);
nand U7980 (N_7980,N_7432,N_6607);
nand U7981 (N_7981,N_5709,N_5072);
nand U7982 (N_7982,N_5790,N_5477);
nor U7983 (N_7983,N_5943,N_5338);
nand U7984 (N_7984,N_7263,N_6794);
or U7985 (N_7985,N_6670,N_6551);
or U7986 (N_7986,N_7097,N_6628);
nor U7987 (N_7987,N_7182,N_6802);
and U7988 (N_7988,N_6881,N_5250);
and U7989 (N_7989,N_5594,N_5872);
or U7990 (N_7990,N_5163,N_7044);
nand U7991 (N_7991,N_6098,N_6183);
nor U7992 (N_7992,N_7439,N_6897);
and U7993 (N_7993,N_7398,N_6007);
and U7994 (N_7994,N_5517,N_6445);
nand U7995 (N_7995,N_6929,N_6630);
or U7996 (N_7996,N_5734,N_6594);
nor U7997 (N_7997,N_5958,N_7119);
nor U7998 (N_7998,N_6612,N_6892);
nand U7999 (N_7999,N_5951,N_5775);
xnor U8000 (N_8000,N_6425,N_5862);
and U8001 (N_8001,N_6561,N_6868);
and U8002 (N_8002,N_5330,N_6017);
or U8003 (N_8003,N_6110,N_5255);
or U8004 (N_8004,N_5768,N_6588);
and U8005 (N_8005,N_6492,N_6186);
and U8006 (N_8006,N_7426,N_6791);
nor U8007 (N_8007,N_5518,N_6730);
or U8008 (N_8008,N_7364,N_6048);
nand U8009 (N_8009,N_7273,N_6271);
and U8010 (N_8010,N_5833,N_5251);
nand U8011 (N_8011,N_7027,N_6571);
or U8012 (N_8012,N_5667,N_6727);
and U8013 (N_8013,N_5784,N_6744);
and U8014 (N_8014,N_6194,N_5827);
nor U8015 (N_8015,N_7405,N_5868);
nand U8016 (N_8016,N_5108,N_5857);
nor U8017 (N_8017,N_5044,N_6156);
nand U8018 (N_8018,N_7075,N_7335);
and U8019 (N_8019,N_5504,N_5474);
nor U8020 (N_8020,N_7226,N_6128);
or U8021 (N_8021,N_6378,N_5742);
and U8022 (N_8022,N_6864,N_5170);
and U8023 (N_8023,N_7393,N_5286);
nor U8024 (N_8024,N_6901,N_6930);
or U8025 (N_8025,N_6044,N_6842);
and U8026 (N_8026,N_5490,N_5417);
or U8027 (N_8027,N_6687,N_5039);
and U8028 (N_8028,N_5907,N_6876);
or U8029 (N_8029,N_6527,N_7190);
nand U8030 (N_8030,N_6420,N_7121);
nor U8031 (N_8031,N_5748,N_5396);
nor U8032 (N_8032,N_5824,N_7475);
nand U8033 (N_8033,N_5401,N_6487);
nand U8034 (N_8034,N_5497,N_6948);
nand U8035 (N_8035,N_6496,N_5562);
and U8036 (N_8036,N_7088,N_7479);
nor U8037 (N_8037,N_6283,N_5254);
and U8038 (N_8038,N_6467,N_6105);
or U8039 (N_8039,N_5803,N_7434);
nand U8040 (N_8040,N_5115,N_6444);
and U8041 (N_8041,N_5646,N_6479);
or U8042 (N_8042,N_6311,N_6089);
or U8043 (N_8043,N_5240,N_7176);
nor U8044 (N_8044,N_6118,N_6873);
or U8045 (N_8045,N_5007,N_6335);
or U8046 (N_8046,N_6773,N_7456);
or U8047 (N_8047,N_5123,N_5012);
nand U8048 (N_8048,N_5971,N_7082);
nand U8049 (N_8049,N_5898,N_6418);
and U8050 (N_8050,N_7068,N_7396);
and U8051 (N_8051,N_5379,N_5712);
and U8052 (N_8052,N_5984,N_6615);
nand U8053 (N_8053,N_5786,N_7309);
nor U8054 (N_8054,N_7274,N_7441);
and U8055 (N_8055,N_5908,N_5349);
nor U8056 (N_8056,N_5236,N_6621);
nor U8057 (N_8057,N_6027,N_6287);
nand U8058 (N_8058,N_5839,N_7126);
or U8059 (N_8059,N_6731,N_6531);
or U8060 (N_8060,N_6680,N_7388);
nand U8061 (N_8061,N_6189,N_6093);
nand U8062 (N_8062,N_7460,N_5663);
nand U8063 (N_8063,N_5798,N_6191);
or U8064 (N_8064,N_6274,N_6443);
nand U8065 (N_8065,N_6632,N_6150);
and U8066 (N_8066,N_6385,N_6978);
or U8067 (N_8067,N_5940,N_5125);
and U8068 (N_8068,N_5904,N_7429);
nand U8069 (N_8069,N_5936,N_5021);
nand U8070 (N_8070,N_7240,N_5619);
xnor U8071 (N_8071,N_6276,N_6669);
nand U8072 (N_8072,N_7401,N_5222);
or U8073 (N_8073,N_5836,N_6766);
and U8074 (N_8074,N_6623,N_6919);
or U8075 (N_8075,N_5415,N_6307);
or U8076 (N_8076,N_7353,N_7269);
or U8077 (N_8077,N_6459,N_5031);
nor U8078 (N_8078,N_6979,N_6721);
and U8079 (N_8079,N_6030,N_5409);
nand U8080 (N_8080,N_5686,N_7380);
or U8081 (N_8081,N_7427,N_6219);
nand U8082 (N_8082,N_6549,N_6337);
nor U8083 (N_8083,N_6533,N_5023);
or U8084 (N_8084,N_6672,N_7490);
nor U8085 (N_8085,N_6754,N_7247);
xnor U8086 (N_8086,N_6682,N_5695);
or U8087 (N_8087,N_5878,N_7206);
and U8088 (N_8088,N_6024,N_5391);
nor U8089 (N_8089,N_6706,N_6771);
nor U8090 (N_8090,N_6907,N_5501);
nand U8091 (N_8091,N_7390,N_7449);
nand U8092 (N_8092,N_5269,N_6338);
or U8093 (N_8093,N_5352,N_6810);
nor U8094 (N_8094,N_6660,N_6051);
nand U8095 (N_8095,N_7002,N_6295);
and U8096 (N_8096,N_7389,N_5202);
and U8097 (N_8097,N_6646,N_6003);
and U8098 (N_8098,N_5041,N_7155);
nand U8099 (N_8099,N_6400,N_6699);
or U8100 (N_8100,N_6392,N_6502);
nand U8101 (N_8101,N_5278,N_6877);
nand U8102 (N_8102,N_5759,N_6343);
or U8103 (N_8103,N_6839,N_6513);
nor U8104 (N_8104,N_5483,N_5733);
nand U8105 (N_8105,N_6541,N_5029);
and U8106 (N_8106,N_6396,N_6861);
nor U8107 (N_8107,N_6071,N_6722);
and U8108 (N_8108,N_7463,N_5591);
nand U8109 (N_8109,N_5214,N_7135);
and U8110 (N_8110,N_6185,N_5773);
or U8111 (N_8111,N_7267,N_6454);
and U8112 (N_8112,N_6849,N_5132);
nor U8113 (N_8113,N_5129,N_6887);
nand U8114 (N_8114,N_6840,N_6980);
nor U8115 (N_8115,N_6812,N_5213);
and U8116 (N_8116,N_6782,N_5791);
or U8117 (N_8117,N_6562,N_6124);
nand U8118 (N_8118,N_5911,N_5555);
nand U8119 (N_8119,N_5084,N_6745);
and U8120 (N_8120,N_6560,N_6215);
and U8121 (N_8121,N_5096,N_6951);
nand U8122 (N_8122,N_5972,N_6031);
nor U8123 (N_8123,N_5196,N_5435);
and U8124 (N_8124,N_6133,N_5580);
nand U8125 (N_8125,N_7421,N_6711);
nor U8126 (N_8126,N_7285,N_6707);
nor U8127 (N_8127,N_5475,N_5996);
nand U8128 (N_8128,N_5296,N_5382);
and U8129 (N_8129,N_5928,N_5234);
nor U8130 (N_8130,N_6775,N_7470);
nand U8131 (N_8131,N_5617,N_5867);
and U8132 (N_8132,N_7070,N_7092);
and U8133 (N_8133,N_5549,N_7227);
nor U8134 (N_8134,N_6399,N_6789);
nand U8135 (N_8135,N_5661,N_6477);
and U8136 (N_8136,N_5749,N_5424);
nor U8137 (N_8137,N_6483,N_7326);
nor U8138 (N_8138,N_6746,N_7482);
nand U8139 (N_8139,N_7181,N_6353);
and U8140 (N_8140,N_5807,N_6101);
nand U8141 (N_8141,N_5398,N_6762);
and U8142 (N_8142,N_6668,N_7036);
nor U8143 (N_8143,N_6823,N_5049);
or U8144 (N_8144,N_5896,N_5885);
nor U8145 (N_8145,N_7123,N_5289);
nand U8146 (N_8146,N_6061,N_5631);
or U8147 (N_8147,N_5624,N_6581);
or U8148 (N_8148,N_5694,N_6237);
and U8149 (N_8149,N_5411,N_6104);
or U8150 (N_8150,N_5188,N_6117);
nor U8151 (N_8151,N_5623,N_7205);
and U8152 (N_8152,N_5055,N_7446);
nor U8153 (N_8153,N_7362,N_6559);
or U8154 (N_8154,N_6554,N_6437);
and U8155 (N_8155,N_5451,N_5581);
nor U8156 (N_8156,N_5347,N_6282);
nor U8157 (N_8157,N_5506,N_6885);
nor U8158 (N_8158,N_7071,N_6164);
and U8159 (N_8159,N_6346,N_5739);
and U8160 (N_8160,N_5525,N_6845);
or U8161 (N_8161,N_6524,N_5428);
nor U8162 (N_8162,N_5077,N_5226);
or U8163 (N_8163,N_6006,N_6278);
nand U8164 (N_8164,N_7058,N_7370);
or U8165 (N_8165,N_5197,N_7278);
and U8166 (N_8166,N_5587,N_5420);
nor U8167 (N_8167,N_6262,N_6931);
nor U8168 (N_8168,N_7189,N_6187);
nand U8169 (N_8169,N_5530,N_6675);
nand U8170 (N_8170,N_5700,N_5886);
and U8171 (N_8171,N_5363,N_6494);
and U8172 (N_8172,N_5446,N_5004);
nor U8173 (N_8173,N_7161,N_5540);
nor U8174 (N_8174,N_5144,N_7302);
nand U8175 (N_8175,N_7474,N_5741);
and U8176 (N_8176,N_6500,N_7087);
nor U8177 (N_8177,N_7187,N_5853);
and U8178 (N_8178,N_6345,N_5737);
or U8179 (N_8179,N_7025,N_5656);
nand U8180 (N_8180,N_5823,N_6700);
and U8181 (N_8181,N_7084,N_5829);
nand U8182 (N_8182,N_5690,N_5588);
and U8183 (N_8183,N_5006,N_5793);
or U8184 (N_8184,N_6521,N_6376);
or U8185 (N_8185,N_7280,N_6056);
or U8186 (N_8186,N_6918,N_5547);
nor U8187 (N_8187,N_7072,N_6086);
or U8188 (N_8188,N_7208,N_6458);
nand U8189 (N_8189,N_6662,N_7488);
nand U8190 (N_8190,N_5837,N_5068);
nand U8191 (N_8191,N_6837,N_7296);
and U8192 (N_8192,N_5750,N_5046);
and U8193 (N_8193,N_5974,N_6201);
nor U8194 (N_8194,N_5452,N_5735);
and U8195 (N_8195,N_7294,N_5206);
nand U8196 (N_8196,N_6499,N_5112);
and U8197 (N_8197,N_5430,N_6574);
and U8198 (N_8198,N_5944,N_5456);
or U8199 (N_8199,N_7241,N_6765);
nor U8200 (N_8200,N_7342,N_6312);
nor U8201 (N_8201,N_5689,N_7374);
and U8202 (N_8202,N_5939,N_5638);
or U8203 (N_8203,N_7341,N_6576);
nor U8204 (N_8204,N_5118,N_5265);
nand U8205 (N_8205,N_5246,N_5910);
and U8206 (N_8206,N_6556,N_5830);
nor U8207 (N_8207,N_6304,N_6084);
nand U8208 (N_8208,N_6501,N_7340);
nor U8209 (N_8209,N_6302,N_5367);
and U8210 (N_8210,N_5463,N_7216);
and U8211 (N_8211,N_6364,N_6116);
nor U8212 (N_8212,N_6427,N_5406);
or U8213 (N_8213,N_5921,N_6126);
and U8214 (N_8214,N_7096,N_5579);
nand U8215 (N_8215,N_5353,N_5462);
nand U8216 (N_8216,N_5941,N_6656);
nor U8217 (N_8217,N_7430,N_5967);
nand U8218 (N_8218,N_6267,N_5455);
and U8219 (N_8219,N_7064,N_7437);
or U8220 (N_8220,N_5800,N_6653);
nor U8221 (N_8221,N_6169,N_5377);
xnor U8222 (N_8222,N_6787,N_5813);
or U8223 (N_8223,N_6152,N_7178);
and U8224 (N_8224,N_5692,N_5544);
and U8225 (N_8225,N_7133,N_7277);
nor U8226 (N_8226,N_5889,N_5754);
nor U8227 (N_8227,N_7332,N_6587);
nand U8228 (N_8228,N_6197,N_7012);
or U8229 (N_8229,N_6976,N_6336);
nand U8230 (N_8230,N_5905,N_5859);
nand U8231 (N_8231,N_7156,N_6685);
and U8232 (N_8232,N_6818,N_6761);
nor U8233 (N_8233,N_6915,N_5920);
or U8234 (N_8234,N_6627,N_6365);
xor U8235 (N_8235,N_5315,N_5718);
nand U8236 (N_8236,N_7368,N_5292);
and U8237 (N_8237,N_5439,N_5512);
nor U8238 (N_8238,N_5043,N_5339);
or U8239 (N_8239,N_5676,N_6036);
xnor U8240 (N_8240,N_7170,N_5765);
nor U8241 (N_8241,N_5195,N_6817);
nand U8242 (N_8242,N_6083,N_5466);
nand U8243 (N_8243,N_7179,N_5284);
and U8244 (N_8244,N_6414,N_5717);
or U8245 (N_8245,N_6253,N_6204);
nor U8246 (N_8246,N_7168,N_6966);
nor U8247 (N_8247,N_6393,N_6333);
and U8248 (N_8248,N_6572,N_7496);
or U8249 (N_8249,N_7233,N_6305);
nand U8250 (N_8250,N_6213,N_7022);
and U8251 (N_8251,N_6352,N_5141);
or U8252 (N_8252,N_7375,N_5806);
and U8253 (N_8253,N_6072,N_6354);
or U8254 (N_8254,N_6898,N_6319);
nor U8255 (N_8255,N_6504,N_6940);
nor U8256 (N_8256,N_6629,N_6171);
nor U8257 (N_8257,N_6493,N_7315);
nand U8258 (N_8258,N_6904,N_7378);
nor U8259 (N_8259,N_5191,N_7103);
or U8260 (N_8260,N_5529,N_6033);
nor U8261 (N_8261,N_5629,N_6430);
nor U8262 (N_8262,N_5584,N_5573);
nand U8263 (N_8263,N_5171,N_6342);
and U8264 (N_8264,N_6696,N_6797);
and U8265 (N_8265,N_7466,N_6803);
and U8266 (N_8266,N_5845,N_5550);
nor U8267 (N_8267,N_6486,N_5541);
or U8268 (N_8268,N_7067,N_6330);
nor U8269 (N_8269,N_5453,N_6905);
and U8270 (N_8270,N_6291,N_5696);
nand U8271 (N_8271,N_7120,N_6684);
nand U8272 (N_8272,N_6617,N_5282);
nand U8273 (N_8273,N_7089,N_5513);
nand U8274 (N_8274,N_5632,N_6638);
and U8275 (N_8275,N_6082,N_5938);
and U8276 (N_8276,N_5851,N_6419);
nand U8277 (N_8277,N_7400,N_5652);
nor U8278 (N_8278,N_7078,N_5707);
and U8279 (N_8279,N_6611,N_5045);
nor U8280 (N_8280,N_7007,N_5683);
nor U8281 (N_8281,N_6734,N_6468);
or U8282 (N_8282,N_5650,N_5078);
or U8283 (N_8283,N_5714,N_6686);
or U8284 (N_8284,N_7107,N_6476);
nand U8285 (N_8285,N_7146,N_5693);
and U8286 (N_8286,N_5738,N_5492);
or U8287 (N_8287,N_5603,N_5478);
and U8288 (N_8288,N_5614,N_6994);
or U8289 (N_8289,N_7129,N_5178);
and U8290 (N_8290,N_6526,N_7354);
or U8291 (N_8291,N_5699,N_5847);
and U8292 (N_8292,N_6403,N_5842);
nor U8293 (N_8293,N_7473,N_6440);
or U8294 (N_8294,N_5854,N_5383);
nor U8295 (N_8295,N_7203,N_5093);
and U8296 (N_8296,N_6906,N_5708);
and U8297 (N_8297,N_5639,N_6566);
or U8298 (N_8298,N_5982,N_5092);
and U8299 (N_8299,N_6610,N_5876);
nand U8300 (N_8300,N_6736,N_6134);
or U8301 (N_8301,N_5852,N_7419);
nor U8302 (N_8302,N_7218,N_5881);
or U8303 (N_8303,N_6958,N_5440);
nand U8304 (N_8304,N_6097,N_5675);
or U8305 (N_8305,N_6301,N_5846);
nand U8306 (N_8306,N_5416,N_6141);
nand U8307 (N_8307,N_5357,N_5993);
nor U8308 (N_8308,N_6637,N_5651);
or U8309 (N_8309,N_6557,N_5390);
and U8310 (N_8310,N_6544,N_7469);
nor U8311 (N_8311,N_6369,N_7198);
and U8312 (N_8312,N_6568,N_7186);
nor U8313 (N_8313,N_5818,N_6780);
and U8314 (N_8314,N_6041,N_6246);
nand U8315 (N_8315,N_5499,N_5776);
or U8316 (N_8316,N_6208,N_5065);
and U8317 (N_8317,N_5894,N_7211);
nor U8318 (N_8318,N_6975,N_7330);
nand U8319 (N_8319,N_6950,N_7109);
or U8320 (N_8320,N_6207,N_6809);
nand U8321 (N_8321,N_6285,N_5877);
nor U8322 (N_8322,N_7039,N_5883);
nor U8323 (N_8323,N_5481,N_6970);
nand U8324 (N_8324,N_6297,N_6855);
nor U8325 (N_8325,N_6382,N_6100);
xor U8326 (N_8326,N_7417,N_5600);
and U8327 (N_8327,N_6843,N_5094);
nand U8328 (N_8328,N_7079,N_6779);
nand U8329 (N_8329,N_6608,N_7177);
and U8330 (N_8330,N_5111,N_5811);
nor U8331 (N_8331,N_5538,N_5668);
nor U8332 (N_8332,N_7316,N_5318);
nand U8333 (N_8333,N_5423,N_6434);
and U8334 (N_8334,N_6142,N_6585);
nand U8335 (N_8335,N_5309,N_5621);
nand U8336 (N_8336,N_6921,N_6108);
or U8337 (N_8337,N_5899,N_5271);
or U8338 (N_8338,N_5551,N_6135);
nor U8339 (N_8339,N_6710,N_5328);
and U8340 (N_8340,N_7220,N_6070);
or U8341 (N_8341,N_5884,N_5966);
and U8342 (N_8342,N_5181,N_6770);
nor U8343 (N_8343,N_6856,N_5297);
and U8344 (N_8344,N_5127,N_6650);
nor U8345 (N_8345,N_6022,N_5169);
and U8346 (N_8346,N_5666,N_5167);
nor U8347 (N_8347,N_6247,N_6619);
or U8348 (N_8348,N_6280,N_5082);
or U8349 (N_8349,N_7276,N_6137);
nor U8350 (N_8350,N_6019,N_6040);
and U8351 (N_8351,N_5515,N_6416);
nand U8352 (N_8352,N_6796,N_7239);
nand U8353 (N_8353,N_6723,N_6895);
nand U8354 (N_8354,N_7160,N_7249);
and U8355 (N_8355,N_6643,N_5482);
or U8356 (N_8356,N_7250,N_6257);
and U8357 (N_8357,N_5644,N_7270);
nor U8358 (N_8358,N_6673,N_5536);
nand U8359 (N_8359,N_5721,N_6768);
nor U8360 (N_8360,N_5404,N_5174);
nand U8361 (N_8361,N_5362,N_6214);
or U8362 (N_8362,N_7003,N_6391);
and U8363 (N_8363,N_7431,N_7260);
nor U8364 (N_8364,N_5546,N_7238);
nand U8365 (N_8365,N_6075,N_6039);
nor U8366 (N_8366,N_5079,N_5266);
nand U8367 (N_8367,N_6021,N_7451);
nor U8368 (N_8368,N_6665,N_6380);
nor U8369 (N_8369,N_6446,N_5053);
and U8370 (N_8370,N_7029,N_6543);
nor U8371 (N_8371,N_6332,N_5556);
nor U8372 (N_8372,N_7091,N_5371);
nand U8373 (N_8373,N_5801,N_6988);
or U8374 (N_8374,N_5945,N_6847);
nand U8375 (N_8375,N_6472,N_7031);
nor U8376 (N_8376,N_6953,N_5070);
nand U8377 (N_8377,N_6455,N_5432);
nor U8378 (N_8378,N_7478,N_6170);
and U8379 (N_8379,N_6645,N_7194);
and U8380 (N_8380,N_6457,N_5295);
or U8381 (N_8381,N_5673,N_6854);
nor U8382 (N_8382,N_5620,N_6218);
or U8383 (N_8383,N_6613,N_6091);
or U8384 (N_8384,N_7191,N_5627);
nand U8385 (N_8385,N_5051,N_5569);
nor U8386 (N_8386,N_7157,N_5081);
nand U8387 (N_8387,N_5351,N_5533);
and U8388 (N_8388,N_7494,N_6625);
and U8389 (N_8389,N_5002,N_7336);
nor U8390 (N_8390,N_5680,N_7219);
nand U8391 (N_8391,N_5783,N_7359);
nor U8392 (N_8392,N_5291,N_5307);
nand U8393 (N_8393,N_6552,N_7049);
nand U8394 (N_8394,N_6225,N_6622);
and U8395 (N_8395,N_7005,N_7344);
nor U8396 (N_8396,N_6870,N_5566);
nor U8397 (N_8397,N_5425,N_5080);
nor U8398 (N_8398,N_5869,N_6955);
nor U8399 (N_8399,N_6087,N_6752);
or U8400 (N_8400,N_6138,N_6661);
nor U8401 (N_8401,N_5755,N_6720);
and U8402 (N_8402,N_5471,N_6321);
nand U8403 (N_8403,N_5724,N_7053);
and U8404 (N_8404,N_7343,N_7272);
or U8405 (N_8405,N_6390,N_5321);
or U8406 (N_8406,N_5162,N_6351);
and U8407 (N_8407,N_6923,N_5633);
nor U8408 (N_8408,N_5048,N_6828);
and U8409 (N_8409,N_5998,N_6123);
nand U8410 (N_8410,N_5126,N_6020);
and U8411 (N_8411,N_6760,N_6703);
nor U8412 (N_8412,N_5804,N_6066);
or U8413 (N_8413,N_6536,N_5395);
or U8414 (N_8414,N_5860,N_5161);
and U8415 (N_8415,N_5808,N_6636);
nand U8416 (N_8416,N_5426,N_5314);
nor U8417 (N_8417,N_6659,N_5986);
or U8418 (N_8418,N_6740,N_5902);
and U8419 (N_8419,N_6255,N_5720);
or U8420 (N_8420,N_6882,N_5571);
and U8421 (N_8421,N_7447,N_5848);
and U8422 (N_8422,N_5316,N_6148);
nor U8423 (N_8423,N_7246,N_5227);
nand U8424 (N_8424,N_6018,N_5746);
nand U8425 (N_8425,N_5324,N_7464);
nor U8426 (N_8426,N_5083,N_5027);
nand U8427 (N_8427,N_6620,N_5918);
nor U8428 (N_8428,N_6254,N_7030);
and U8429 (N_8429,N_5211,N_6453);
nor U8430 (N_8430,N_5779,N_7132);
nor U8431 (N_8431,N_5313,N_6508);
and U8432 (N_8432,N_5959,N_7413);
or U8433 (N_8433,N_7320,N_6708);
and U8434 (N_8434,N_5259,N_6163);
and U8435 (N_8435,N_5931,N_7037);
nand U8436 (N_8436,N_5821,N_7472);
and U8437 (N_8437,N_5261,N_5653);
nand U8438 (N_8438,N_7314,N_6053);
xor U8439 (N_8439,N_7019,N_6047);
or U8440 (N_8440,N_5034,N_5102);
nand U8441 (N_8441,N_7171,N_5526);
nand U8442 (N_8442,N_6639,N_6067);
and U8443 (N_8443,N_5397,N_5670);
and U8444 (N_8444,N_7379,N_6863);
nor U8445 (N_8445,N_6062,N_7334);
and U8446 (N_8446,N_7043,N_5058);
nand U8447 (N_8447,N_5010,N_6914);
nand U8448 (N_8448,N_6753,N_5366);
nand U8449 (N_8449,N_5625,N_7093);
or U8450 (N_8450,N_6323,N_5185);
or U8451 (N_8451,N_6565,N_6939);
nand U8452 (N_8452,N_6719,N_5688);
and U8453 (N_8453,N_6737,N_5710);
or U8454 (N_8454,N_6626,N_6235);
and U8455 (N_8455,N_7312,N_5687);
nand U8456 (N_8456,N_5128,N_6635);
nor U8457 (N_8457,N_6936,N_5507);
nand U8458 (N_8458,N_6388,N_6413);
and U8459 (N_8459,N_7017,N_5864);
and U8460 (N_8460,N_6582,N_7305);
and U8461 (N_8461,N_7297,N_6344);
or U8462 (N_8462,N_6999,N_5563);
nand U8463 (N_8463,N_7201,N_5464);
nand U8464 (N_8464,N_7151,N_6046);
or U8465 (N_8465,N_7484,N_6725);
nand U8466 (N_8466,N_5075,N_6422);
nand U8467 (N_8467,N_6598,N_5450);
and U8468 (N_8468,N_6474,N_7369);
or U8469 (N_8469,N_5183,N_5275);
nor U8470 (N_8470,N_6981,N_5891);
nand U8471 (N_8471,N_7409,N_6426);
or U8472 (N_8472,N_7468,N_7033);
or U8473 (N_8473,N_6010,N_6002);
and U8474 (N_8474,N_5257,N_6605);
or U8475 (N_8475,N_6200,N_6742);
nor U8476 (N_8476,N_7066,N_7040);
and U8477 (N_8477,N_7303,N_5215);
or U8478 (N_8478,N_6555,N_5370);
nor U8479 (N_8479,N_6149,N_6972);
nand U8480 (N_8480,N_7311,N_6769);
and U8481 (N_8481,N_6448,N_5769);
nand U8482 (N_8482,N_5441,N_6339);
or U8483 (N_8483,N_5494,N_5973);
or U8484 (N_8484,N_7077,N_6878);
and U8485 (N_8485,N_7153,N_5469);
and U8486 (N_8486,N_5205,N_6166);
and U8487 (N_8487,N_6961,N_6269);
and U8488 (N_8488,N_6293,N_6389);
nand U8489 (N_8489,N_5731,N_7392);
nand U8490 (N_8490,N_7165,N_6614);
nor U8491 (N_8491,N_7197,N_6715);
nand U8492 (N_8492,N_6463,N_5369);
or U8493 (N_8493,N_6289,N_5642);
nor U8494 (N_8494,N_6833,N_6143);
and U8495 (N_8495,N_6316,N_7056);
nand U8496 (N_8496,N_7124,N_7265);
or U8497 (N_8497,N_6452,N_5949);
or U8498 (N_8498,N_6052,N_6441);
and U8499 (N_8499,N_5655,N_7173);
nor U8500 (N_8500,N_6180,N_5495);
nand U8501 (N_8501,N_5523,N_5210);
and U8502 (N_8502,N_7234,N_6530);
nor U8503 (N_8503,N_6449,N_5698);
and U8504 (N_8504,N_6807,N_6428);
and U8505 (N_8505,N_5454,N_7423);
or U8506 (N_8506,N_6801,N_5303);
nand U8507 (N_8507,N_6367,N_5616);
and U8508 (N_8508,N_5496,N_6633);
and U8509 (N_8509,N_6509,N_5312);
and U8510 (N_8510,N_6820,N_6729);
and U8511 (N_8511,N_7458,N_5782);
or U8512 (N_8512,N_7048,N_6155);
or U8513 (N_8513,N_5923,N_6860);
or U8514 (N_8514,N_6925,N_7042);
nand U8515 (N_8515,N_5086,N_5248);
and U8516 (N_8516,N_6529,N_6952);
and U8517 (N_8517,N_5095,N_5874);
and U8518 (N_8518,N_5465,N_5997);
nand U8519 (N_8519,N_6242,N_7105);
nor U8520 (N_8520,N_6484,N_6968);
nor U8521 (N_8521,N_6690,N_6404);
nor U8522 (N_8522,N_5865,N_6313);
nand U8523 (N_8523,N_5458,N_5294);
and U8524 (N_8524,N_6265,N_6165);
nor U8525 (N_8525,N_5747,N_6034);
or U8526 (N_8526,N_6160,N_5263);
or U8527 (N_8527,N_6678,N_5493);
nor U8528 (N_8528,N_6591,N_5796);
and U8529 (N_8529,N_5585,N_6334);
nand U8530 (N_8530,N_5434,N_6349);
nor U8531 (N_8531,N_7094,N_6666);
nand U8532 (N_8532,N_5160,N_7131);
and U8533 (N_8533,N_7180,N_6798);
or U8534 (N_8534,N_5757,N_6835);
or U8535 (N_8535,N_7321,N_5751);
nor U8536 (N_8536,N_6216,N_6375);
nand U8537 (N_8537,N_5643,N_6553);
and U8538 (N_8538,N_7188,N_6055);
or U8539 (N_8539,N_6231,N_5336);
nand U8540 (N_8540,N_5812,N_6360);
or U8541 (N_8541,N_5221,N_5955);
and U8542 (N_8542,N_7054,N_6922);
nor U8543 (N_8543,N_5822,N_6049);
or U8544 (N_8544,N_5119,N_6564);
xor U8545 (N_8545,N_5327,N_6618);
nand U8546 (N_8546,N_6016,N_6850);
nor U8547 (N_8547,N_7235,N_7147);
and U8548 (N_8548,N_7221,N_6967);
nand U8549 (N_8549,N_6514,N_7081);
and U8550 (N_8550,N_6038,N_6395);
or U8551 (N_8551,N_6569,N_6078);
nor U8552 (N_8552,N_7073,N_7009);
nand U8553 (N_8553,N_7231,N_6111);
nor U8554 (N_8554,N_6756,N_7116);
xnor U8555 (N_8555,N_5135,N_5237);
or U8556 (N_8556,N_6012,N_5553);
nor U8557 (N_8557,N_7145,N_5033);
and U8558 (N_8558,N_7453,N_5385);
and U8559 (N_8559,N_5293,N_6232);
nand U8560 (N_8560,N_7495,N_6702);
and U8561 (N_8561,N_5596,N_6983);
nand U8562 (N_8562,N_5323,N_6857);
nor U8563 (N_8563,N_6308,N_6634);
nor U8564 (N_8564,N_7050,N_6741);
nor U8565 (N_8565,N_5730,N_6366);
nor U8566 (N_8566,N_5179,N_5052);
nor U8567 (N_8567,N_7384,N_7440);
nand U8568 (N_8568,N_5393,N_7166);
and U8569 (N_8569,N_5028,N_5560);
and U8570 (N_8570,N_5368,N_6874);
or U8571 (N_8571,N_6903,N_6397);
and U8572 (N_8572,N_6172,N_6431);
and U8573 (N_8573,N_7443,N_6196);
and U8574 (N_8574,N_6728,N_5788);
nand U8575 (N_8575,N_6814,N_6243);
and U8576 (N_8576,N_5715,N_6992);
or U8577 (N_8577,N_7399,N_5610);
or U8578 (N_8578,N_5946,N_5795);
nor U8579 (N_8579,N_7245,N_6743);
or U8580 (N_8580,N_5545,N_6341);
or U8581 (N_8581,N_6478,N_6912);
and U8582 (N_8582,N_5262,N_5866);
nor U8583 (N_8583,N_7154,N_5283);
nor U8584 (N_8584,N_6859,N_6516);
nand U8585 (N_8585,N_7497,N_7035);
and U8586 (N_8586,N_6136,N_6069);
nor U8587 (N_8587,N_6671,N_6935);
and U8588 (N_8588,N_5671,N_5729);
nand U8589 (N_8589,N_7418,N_7499);
or U8590 (N_8590,N_5326,N_5723);
nand U8591 (N_8591,N_7422,N_5479);
and U8592 (N_8592,N_6933,N_6913);
and U8593 (N_8593,N_7106,N_6573);
and U8594 (N_8594,N_5225,N_5346);
or U8595 (N_8595,N_5489,N_6460);
and U8596 (N_8596,N_7385,N_5505);
or U8597 (N_8597,N_6411,N_7333);
nor U8598 (N_8598,N_6256,N_5134);
and U8599 (N_8599,N_6786,N_5038);
or U8600 (N_8600,N_5534,N_6314);
or U8601 (N_8601,N_7465,N_6688);
and U8602 (N_8602,N_7477,N_7158);
or U8603 (N_8603,N_6439,N_6158);
nand U8604 (N_8604,N_6306,N_5011);
and U8605 (N_8605,N_6127,N_5914);
nor U8606 (N_8606,N_5468,N_7010);
nand U8607 (N_8607,N_5992,N_7410);
nand U8608 (N_8608,N_5136,N_5609);
or U8609 (N_8609,N_7331,N_5001);
or U8610 (N_8610,N_5008,N_7024);
or U8611 (N_8611,N_5520,N_5040);
nor U8612 (N_8612,N_6374,N_5740);
nand U8613 (N_8613,N_5554,N_6092);
nor U8614 (N_8614,N_7018,N_5341);
and U8615 (N_8615,N_6358,N_6259);
nor U8616 (N_8616,N_6490,N_5238);
nand U8617 (N_8617,N_6996,N_6889);
and U8618 (N_8618,N_7298,N_6589);
and U8619 (N_8619,N_6355,N_5977);
and U8620 (N_8620,N_7348,N_5037);
nor U8621 (N_8621,N_5106,N_5766);
or U8622 (N_8622,N_7136,N_5107);
or U8623 (N_8623,N_5532,N_7175);
and U8624 (N_8624,N_5771,N_5022);
and U8625 (N_8625,N_5764,N_5194);
and U8626 (N_8626,N_6748,N_5099);
nand U8627 (N_8627,N_5948,N_7324);
and U8628 (N_8628,N_6228,N_5090);
or U8629 (N_8629,N_5218,N_5725);
nor U8630 (N_8630,N_5147,N_6233);
and U8631 (N_8631,N_5564,N_7061);
and U8632 (N_8632,N_5835,N_6558);
nor U8633 (N_8633,N_6956,N_5375);
or U8634 (N_8634,N_6384,N_7371);
or U8635 (N_8635,N_6230,N_6651);
nor U8636 (N_8636,N_5317,N_5875);
nor U8637 (N_8637,N_5414,N_6869);
or U8638 (N_8638,N_7062,N_7360);
nor U8639 (N_8639,N_6808,N_5220);
nor U8640 (N_8640,N_5602,N_5572);
xnor U8641 (N_8641,N_7345,N_5264);
or U8642 (N_8642,N_6266,N_5577);
nor U8643 (N_8643,N_5105,N_7052);
nor U8644 (N_8644,N_6188,N_7377);
nand U8645 (N_8645,N_5150,N_5753);
nor U8646 (N_8646,N_7242,N_7143);
nor U8647 (N_8647,N_5919,N_5421);
nand U8648 (N_8648,N_5155,N_6469);
nand U8649 (N_8649,N_5364,N_6647);
and U8650 (N_8650,N_6106,N_5901);
or U8651 (N_8651,N_5319,N_5528);
or U8652 (N_8652,N_6693,N_5970);
nand U8653 (N_8653,N_6379,N_6025);
nor U8654 (N_8654,N_5780,N_6281);
or U8655 (N_8655,N_5104,N_5916);
nor U8656 (N_8656,N_7412,N_7347);
or U8657 (N_8657,N_6324,N_6945);
or U8658 (N_8658,N_5359,N_5354);
or U8659 (N_8659,N_5244,N_5431);
and U8660 (N_8660,N_5252,N_5356);
nand U8661 (N_8661,N_5567,N_5117);
nor U8662 (N_8662,N_6821,N_6718);
nand U8663 (N_8663,N_7352,N_7411);
nor U8664 (N_8664,N_6205,N_5066);
or U8665 (N_8665,N_7207,N_7229);
or U8666 (N_8666,N_5267,N_5664);
nand U8667 (N_8667,N_5378,N_5290);
nand U8668 (N_8668,N_5302,N_6899);
nor U8669 (N_8669,N_7223,N_5592);
nor U8670 (N_8670,N_7117,N_6758);
and U8671 (N_8671,N_6456,N_5964);
or U8672 (N_8672,N_5436,N_6804);
or U8673 (N_8673,N_7065,N_5116);
nor U8674 (N_8674,N_5511,N_6606);
or U8675 (N_8675,N_6107,N_5487);
and U8676 (N_8676,N_5756,N_5476);
nor U8677 (N_8677,N_5071,N_7372);
nor U8678 (N_8678,N_6240,N_6712);
or U8679 (N_8679,N_7045,N_6631);
and U8680 (N_8680,N_6713,N_6229);
nor U8681 (N_8681,N_5758,N_6248);
xnor U8682 (N_8682,N_5726,N_6674);
or U8683 (N_8683,N_6251,N_6028);
and U8684 (N_8684,N_5942,N_6738);
or U8685 (N_8685,N_5335,N_6410);
nor U8686 (N_8686,N_6340,N_5233);
or U8687 (N_8687,N_6886,N_7055);
and U8688 (N_8688,N_6145,N_6120);
nand U8689 (N_8689,N_6641,N_6916);
nor U8690 (N_8690,N_6438,N_6872);
or U8691 (N_8691,N_6222,N_5537);
or U8692 (N_8692,N_5472,N_7101);
nor U8693 (N_8693,N_5565,N_6510);
and U8694 (N_8694,N_5208,N_6327);
nor U8695 (N_8695,N_6076,N_5559);
or U8696 (N_8696,N_6540,N_7047);
xnor U8697 (N_8697,N_5374,N_7006);
and U8698 (N_8698,N_7304,N_6778);
or U8699 (N_8699,N_6264,N_6519);
or U8700 (N_8700,N_6523,N_7366);
and U8701 (N_8701,N_7141,N_5427);
and U8702 (N_8702,N_5858,N_6129);
nand U8703 (N_8703,N_6829,N_5930);
and U8704 (N_8704,N_5201,N_6816);
nand U8705 (N_8705,N_6210,N_7152);
nand U8706 (N_8706,N_6652,N_5403);
or U8707 (N_8707,N_7262,N_6482);
nand U8708 (N_8708,N_6987,N_5979);
or U8709 (N_8709,N_6065,N_7416);
nand U8710 (N_8710,N_6811,N_6198);
nand U8711 (N_8711,N_5322,N_7192);
nor U8712 (N_8712,N_5063,N_7225);
xor U8713 (N_8713,N_7266,N_7021);
nor U8714 (N_8714,N_5985,N_7202);
nor U8715 (N_8715,N_7172,N_5005);
nand U8716 (N_8716,N_5856,N_7287);
nand U8717 (N_8717,N_7140,N_7252);
and U8718 (N_8718,N_6781,N_7471);
and U8719 (N_8719,N_5203,N_6447);
nor U8720 (N_8720,N_5177,N_6008);
and U8721 (N_8721,N_6325,N_6317);
or U8722 (N_8722,N_6296,N_5636);
nor U8723 (N_8723,N_5457,N_6320);
nor U8724 (N_8724,N_5669,N_6954);
nor U8725 (N_8725,N_7076,N_6429);
nor U8726 (N_8726,N_7271,N_6241);
or U8727 (N_8727,N_6776,N_5647);
or U8728 (N_8728,N_5648,N_6015);
and U8729 (N_8729,N_5521,N_7433);
and U8730 (N_8730,N_5976,N_5557);
nand U8731 (N_8731,N_5777,N_6294);
nor U8732 (N_8732,N_5947,N_7016);
nor U8733 (N_8733,N_6601,N_6121);
and U8734 (N_8734,N_5407,N_6239);
nor U8735 (N_8735,N_6575,N_6932);
nor U8736 (N_8736,N_6277,N_6211);
nor U8737 (N_8737,N_5032,N_5030);
and U8738 (N_8738,N_5932,N_6408);
and U8739 (N_8739,N_7243,N_6503);
nor U8740 (N_8740,N_7455,N_7361);
nand U8741 (N_8741,N_6714,N_6971);
or U8742 (N_8742,N_6348,N_6667);
nand U8743 (N_8743,N_5841,N_7014);
and U8744 (N_8744,N_6701,N_6567);
or U8745 (N_8745,N_5834,N_7358);
nand U8746 (N_8746,N_5912,N_7169);
nor U8747 (N_8747,N_6063,N_7074);
nand U8748 (N_8748,N_6580,N_5204);
and U8749 (N_8749,N_5679,N_5332);
and U8750 (N_8750,N_5229,N_6392);
nor U8751 (N_8751,N_6024,N_5742);
nor U8752 (N_8752,N_6336,N_5646);
nand U8753 (N_8753,N_6947,N_6816);
and U8754 (N_8754,N_5912,N_6574);
nor U8755 (N_8755,N_7117,N_6911);
nand U8756 (N_8756,N_6647,N_6350);
and U8757 (N_8757,N_5963,N_5056);
and U8758 (N_8758,N_5330,N_5253);
nand U8759 (N_8759,N_6139,N_7277);
or U8760 (N_8760,N_5807,N_5926);
and U8761 (N_8761,N_6692,N_6741);
and U8762 (N_8762,N_6948,N_5840);
nand U8763 (N_8763,N_6693,N_6643);
and U8764 (N_8764,N_6662,N_6583);
nor U8765 (N_8765,N_6192,N_5901);
nand U8766 (N_8766,N_6159,N_6368);
xor U8767 (N_8767,N_7129,N_5934);
nand U8768 (N_8768,N_6918,N_6285);
or U8769 (N_8769,N_6503,N_5407);
nor U8770 (N_8770,N_6657,N_5558);
and U8771 (N_8771,N_6090,N_6837);
nand U8772 (N_8772,N_5517,N_5322);
and U8773 (N_8773,N_6571,N_6999);
and U8774 (N_8774,N_5139,N_5193);
nand U8775 (N_8775,N_7435,N_7461);
nor U8776 (N_8776,N_5295,N_7121);
nor U8777 (N_8777,N_5917,N_5303);
nor U8778 (N_8778,N_5235,N_6685);
and U8779 (N_8779,N_5156,N_5263);
and U8780 (N_8780,N_6886,N_6687);
or U8781 (N_8781,N_6974,N_5750);
nor U8782 (N_8782,N_7190,N_6331);
nor U8783 (N_8783,N_7019,N_5320);
or U8784 (N_8784,N_6571,N_6247);
nor U8785 (N_8785,N_5781,N_5136);
nand U8786 (N_8786,N_6928,N_7281);
or U8787 (N_8787,N_6695,N_5995);
or U8788 (N_8788,N_5441,N_5849);
nand U8789 (N_8789,N_6901,N_6244);
nor U8790 (N_8790,N_6341,N_7239);
or U8791 (N_8791,N_5690,N_6301);
nand U8792 (N_8792,N_5018,N_5127);
and U8793 (N_8793,N_6113,N_5177);
nor U8794 (N_8794,N_5654,N_7406);
nand U8795 (N_8795,N_6158,N_6942);
nor U8796 (N_8796,N_5034,N_5186);
or U8797 (N_8797,N_6226,N_6134);
nor U8798 (N_8798,N_5210,N_5311);
or U8799 (N_8799,N_6098,N_5397);
or U8800 (N_8800,N_6033,N_6505);
or U8801 (N_8801,N_6900,N_6882);
nand U8802 (N_8802,N_7405,N_5956);
nor U8803 (N_8803,N_7073,N_6939);
nor U8804 (N_8804,N_6093,N_5332);
or U8805 (N_8805,N_5381,N_6687);
or U8806 (N_8806,N_7304,N_5265);
nor U8807 (N_8807,N_5756,N_6954);
nand U8808 (N_8808,N_5279,N_7345);
nor U8809 (N_8809,N_6410,N_5886);
nor U8810 (N_8810,N_5119,N_6727);
nor U8811 (N_8811,N_5990,N_5235);
nand U8812 (N_8812,N_5234,N_6244);
nand U8813 (N_8813,N_6632,N_5248);
nor U8814 (N_8814,N_7421,N_5498);
xnor U8815 (N_8815,N_7490,N_5152);
and U8816 (N_8816,N_6837,N_5347);
and U8817 (N_8817,N_5082,N_5834);
nand U8818 (N_8818,N_6759,N_5806);
nor U8819 (N_8819,N_6157,N_6947);
nand U8820 (N_8820,N_5876,N_7252);
nand U8821 (N_8821,N_5125,N_7255);
or U8822 (N_8822,N_5353,N_7250);
and U8823 (N_8823,N_6556,N_5255);
and U8824 (N_8824,N_5808,N_6534);
nand U8825 (N_8825,N_7217,N_5156);
or U8826 (N_8826,N_6462,N_5144);
or U8827 (N_8827,N_6569,N_7378);
or U8828 (N_8828,N_5793,N_6649);
or U8829 (N_8829,N_7085,N_6861);
and U8830 (N_8830,N_5847,N_7186);
nand U8831 (N_8831,N_5625,N_7193);
nor U8832 (N_8832,N_5538,N_6514);
xor U8833 (N_8833,N_6979,N_6653);
nor U8834 (N_8834,N_7434,N_5512);
nor U8835 (N_8835,N_6294,N_6242);
nand U8836 (N_8836,N_5350,N_5355);
nor U8837 (N_8837,N_5318,N_7385);
and U8838 (N_8838,N_7385,N_5498);
nand U8839 (N_8839,N_5224,N_5194);
or U8840 (N_8840,N_6872,N_6786);
nand U8841 (N_8841,N_5239,N_6828);
nor U8842 (N_8842,N_7343,N_6656);
nand U8843 (N_8843,N_6462,N_5345);
nand U8844 (N_8844,N_5356,N_5560);
nand U8845 (N_8845,N_7376,N_6031);
nand U8846 (N_8846,N_7400,N_6257);
nand U8847 (N_8847,N_7112,N_5459);
nand U8848 (N_8848,N_5852,N_7466);
nor U8849 (N_8849,N_6511,N_6398);
nor U8850 (N_8850,N_7334,N_6065);
nand U8851 (N_8851,N_5194,N_5372);
nor U8852 (N_8852,N_5579,N_7172);
nor U8853 (N_8853,N_6314,N_6405);
nor U8854 (N_8854,N_6081,N_7166);
and U8855 (N_8855,N_7343,N_7242);
nor U8856 (N_8856,N_5847,N_7276);
and U8857 (N_8857,N_6537,N_7200);
or U8858 (N_8858,N_7417,N_6040);
or U8859 (N_8859,N_5086,N_7455);
nor U8860 (N_8860,N_7080,N_6671);
or U8861 (N_8861,N_6875,N_6686);
nor U8862 (N_8862,N_6414,N_6598);
nor U8863 (N_8863,N_6619,N_6071);
nand U8864 (N_8864,N_5768,N_6845);
and U8865 (N_8865,N_6585,N_5464);
nand U8866 (N_8866,N_7498,N_6462);
or U8867 (N_8867,N_6993,N_7390);
or U8868 (N_8868,N_5878,N_6236);
nor U8869 (N_8869,N_6323,N_5493);
or U8870 (N_8870,N_7281,N_7451);
and U8871 (N_8871,N_6840,N_6345);
and U8872 (N_8872,N_6013,N_6611);
or U8873 (N_8873,N_6455,N_5923);
nand U8874 (N_8874,N_5913,N_7456);
or U8875 (N_8875,N_7019,N_6838);
nand U8876 (N_8876,N_5950,N_5750);
and U8877 (N_8877,N_5481,N_6354);
nand U8878 (N_8878,N_6937,N_5638);
nand U8879 (N_8879,N_7311,N_5297);
or U8880 (N_8880,N_6674,N_6699);
and U8881 (N_8881,N_6907,N_6804);
and U8882 (N_8882,N_5145,N_7281);
and U8883 (N_8883,N_6508,N_5335);
or U8884 (N_8884,N_5716,N_6892);
nand U8885 (N_8885,N_6754,N_5688);
and U8886 (N_8886,N_6375,N_7369);
or U8887 (N_8887,N_7100,N_6388);
or U8888 (N_8888,N_5466,N_7487);
nor U8889 (N_8889,N_5845,N_6185);
or U8890 (N_8890,N_5144,N_6764);
nor U8891 (N_8891,N_6258,N_6163);
and U8892 (N_8892,N_6016,N_5868);
or U8893 (N_8893,N_6012,N_6224);
or U8894 (N_8894,N_5969,N_6710);
or U8895 (N_8895,N_6862,N_7451);
or U8896 (N_8896,N_7437,N_5318);
nand U8897 (N_8897,N_5769,N_6533);
and U8898 (N_8898,N_6512,N_6542);
nor U8899 (N_8899,N_6273,N_6760);
nor U8900 (N_8900,N_7317,N_7446);
nor U8901 (N_8901,N_6634,N_6652);
or U8902 (N_8902,N_7456,N_6408);
nor U8903 (N_8903,N_6213,N_6313);
or U8904 (N_8904,N_5071,N_6132);
or U8905 (N_8905,N_6494,N_6678);
nand U8906 (N_8906,N_6195,N_7239);
or U8907 (N_8907,N_5544,N_5972);
nor U8908 (N_8908,N_5745,N_7230);
and U8909 (N_8909,N_6220,N_5124);
and U8910 (N_8910,N_5759,N_6774);
nor U8911 (N_8911,N_5626,N_5072);
and U8912 (N_8912,N_5829,N_5721);
nand U8913 (N_8913,N_6358,N_7067);
or U8914 (N_8914,N_5809,N_5884);
and U8915 (N_8915,N_5357,N_6423);
and U8916 (N_8916,N_6403,N_5095);
and U8917 (N_8917,N_6407,N_5064);
or U8918 (N_8918,N_5915,N_6086);
nor U8919 (N_8919,N_6409,N_6699);
nand U8920 (N_8920,N_6572,N_5862);
or U8921 (N_8921,N_7485,N_6619);
and U8922 (N_8922,N_5385,N_5063);
or U8923 (N_8923,N_5838,N_6775);
or U8924 (N_8924,N_5686,N_7266);
or U8925 (N_8925,N_5577,N_6879);
nand U8926 (N_8926,N_7036,N_6798);
nor U8927 (N_8927,N_6552,N_7273);
nor U8928 (N_8928,N_5234,N_6959);
and U8929 (N_8929,N_7453,N_5937);
or U8930 (N_8930,N_7432,N_6600);
or U8931 (N_8931,N_6540,N_5066);
nand U8932 (N_8932,N_5916,N_6995);
nor U8933 (N_8933,N_7463,N_5139);
or U8934 (N_8934,N_6575,N_6402);
and U8935 (N_8935,N_5748,N_5259);
nor U8936 (N_8936,N_5528,N_5175);
nor U8937 (N_8937,N_5733,N_7172);
or U8938 (N_8938,N_5801,N_6996);
and U8939 (N_8939,N_5280,N_5000);
and U8940 (N_8940,N_7296,N_5811);
nand U8941 (N_8941,N_5071,N_6910);
or U8942 (N_8942,N_7131,N_6365);
and U8943 (N_8943,N_6629,N_6063);
or U8944 (N_8944,N_5616,N_6021);
or U8945 (N_8945,N_6513,N_6469);
nor U8946 (N_8946,N_6581,N_5552);
or U8947 (N_8947,N_5258,N_6725);
nand U8948 (N_8948,N_5726,N_7321);
nand U8949 (N_8949,N_6354,N_6160);
or U8950 (N_8950,N_6173,N_6750);
nor U8951 (N_8951,N_5279,N_7116);
or U8952 (N_8952,N_7256,N_6165);
or U8953 (N_8953,N_6127,N_6672);
nor U8954 (N_8954,N_6647,N_6479);
and U8955 (N_8955,N_5473,N_6413);
nor U8956 (N_8956,N_7020,N_6071);
and U8957 (N_8957,N_6658,N_5451);
and U8958 (N_8958,N_7479,N_7104);
nor U8959 (N_8959,N_5571,N_5330);
and U8960 (N_8960,N_7490,N_6904);
nand U8961 (N_8961,N_6672,N_5497);
xor U8962 (N_8962,N_6543,N_7232);
nand U8963 (N_8963,N_7154,N_5902);
nor U8964 (N_8964,N_6518,N_6094);
or U8965 (N_8965,N_5374,N_5781);
nor U8966 (N_8966,N_7466,N_7483);
or U8967 (N_8967,N_6486,N_6658);
or U8968 (N_8968,N_7031,N_5599);
xnor U8969 (N_8969,N_5463,N_5362);
nor U8970 (N_8970,N_6585,N_5309);
or U8971 (N_8971,N_5395,N_6500);
or U8972 (N_8972,N_5854,N_6061);
nand U8973 (N_8973,N_6140,N_5974);
and U8974 (N_8974,N_6856,N_6042);
nor U8975 (N_8975,N_6917,N_6368);
and U8976 (N_8976,N_6824,N_5568);
or U8977 (N_8977,N_6992,N_5872);
nor U8978 (N_8978,N_6509,N_6836);
or U8979 (N_8979,N_6747,N_5514);
and U8980 (N_8980,N_5816,N_5108);
nand U8981 (N_8981,N_7059,N_6753);
nand U8982 (N_8982,N_7489,N_6014);
nand U8983 (N_8983,N_5926,N_6677);
nand U8984 (N_8984,N_7035,N_6531);
nand U8985 (N_8985,N_6112,N_6395);
or U8986 (N_8986,N_6615,N_6485);
nand U8987 (N_8987,N_6787,N_6951);
or U8988 (N_8988,N_7267,N_5681);
nor U8989 (N_8989,N_6647,N_6919);
nand U8990 (N_8990,N_6607,N_5102);
nand U8991 (N_8991,N_5101,N_6708);
nand U8992 (N_8992,N_5308,N_6210);
and U8993 (N_8993,N_6052,N_6129);
or U8994 (N_8994,N_5549,N_6509);
or U8995 (N_8995,N_5198,N_5694);
nor U8996 (N_8996,N_5799,N_6193);
nand U8997 (N_8997,N_7276,N_6228);
and U8998 (N_8998,N_6895,N_5550);
and U8999 (N_8999,N_5046,N_7058);
nand U9000 (N_9000,N_5986,N_6810);
nand U9001 (N_9001,N_6683,N_7476);
nand U9002 (N_9002,N_5119,N_6029);
nand U9003 (N_9003,N_5835,N_6950);
nand U9004 (N_9004,N_6991,N_6735);
nand U9005 (N_9005,N_5765,N_6492);
nor U9006 (N_9006,N_5744,N_6145);
nor U9007 (N_9007,N_6428,N_6706);
or U9008 (N_9008,N_5255,N_6516);
nor U9009 (N_9009,N_6419,N_6405);
or U9010 (N_9010,N_5377,N_6733);
or U9011 (N_9011,N_7035,N_6560);
nand U9012 (N_9012,N_5104,N_5747);
or U9013 (N_9013,N_5262,N_6826);
or U9014 (N_9014,N_6461,N_6789);
and U9015 (N_9015,N_6256,N_6781);
and U9016 (N_9016,N_7424,N_7312);
nor U9017 (N_9017,N_5680,N_5703);
or U9018 (N_9018,N_6506,N_6554);
nand U9019 (N_9019,N_6957,N_7318);
nor U9020 (N_9020,N_5393,N_6979);
nor U9021 (N_9021,N_5827,N_6258);
or U9022 (N_9022,N_6360,N_5935);
nand U9023 (N_9023,N_6865,N_5202);
and U9024 (N_9024,N_6171,N_6659);
nand U9025 (N_9025,N_5698,N_6192);
and U9026 (N_9026,N_6696,N_7423);
and U9027 (N_9027,N_6585,N_7065);
and U9028 (N_9028,N_5070,N_6173);
xor U9029 (N_9029,N_5063,N_6252);
nand U9030 (N_9030,N_7083,N_5225);
or U9031 (N_9031,N_6383,N_7382);
or U9032 (N_9032,N_6814,N_7299);
and U9033 (N_9033,N_5666,N_5522);
nor U9034 (N_9034,N_5381,N_5646);
and U9035 (N_9035,N_7237,N_6672);
or U9036 (N_9036,N_5701,N_5941);
nor U9037 (N_9037,N_6272,N_5700);
nor U9038 (N_9038,N_6494,N_6076);
and U9039 (N_9039,N_7431,N_6662);
and U9040 (N_9040,N_5357,N_5237);
nor U9041 (N_9041,N_7051,N_5486);
or U9042 (N_9042,N_6774,N_5529);
nor U9043 (N_9043,N_5491,N_7474);
nor U9044 (N_9044,N_5602,N_6821);
nand U9045 (N_9045,N_5100,N_6496);
or U9046 (N_9046,N_5677,N_7119);
and U9047 (N_9047,N_5131,N_5450);
and U9048 (N_9048,N_5355,N_7418);
and U9049 (N_9049,N_6267,N_7495);
or U9050 (N_9050,N_7396,N_5546);
nor U9051 (N_9051,N_6681,N_6826);
and U9052 (N_9052,N_7251,N_5245);
or U9053 (N_9053,N_7427,N_5759);
nor U9054 (N_9054,N_5902,N_5064);
nand U9055 (N_9055,N_5591,N_6675);
nand U9056 (N_9056,N_6018,N_5083);
nand U9057 (N_9057,N_7228,N_6250);
nand U9058 (N_9058,N_6079,N_6597);
and U9059 (N_9059,N_7162,N_7001);
nand U9060 (N_9060,N_5678,N_5057);
nand U9061 (N_9061,N_5116,N_6935);
xnor U9062 (N_9062,N_5093,N_5478);
nor U9063 (N_9063,N_5759,N_6443);
and U9064 (N_9064,N_6271,N_6989);
nand U9065 (N_9065,N_6254,N_5902);
nand U9066 (N_9066,N_5761,N_6126);
or U9067 (N_9067,N_7450,N_6714);
nor U9068 (N_9068,N_6250,N_5959);
and U9069 (N_9069,N_6599,N_7160);
or U9070 (N_9070,N_6730,N_7184);
and U9071 (N_9071,N_5609,N_5110);
or U9072 (N_9072,N_5879,N_7293);
and U9073 (N_9073,N_6941,N_7351);
nand U9074 (N_9074,N_5161,N_6265);
nor U9075 (N_9075,N_5240,N_6542);
and U9076 (N_9076,N_5818,N_7123);
or U9077 (N_9077,N_6261,N_5831);
nor U9078 (N_9078,N_5779,N_7072);
nand U9079 (N_9079,N_6076,N_6737);
nor U9080 (N_9080,N_5470,N_7327);
and U9081 (N_9081,N_5370,N_6441);
or U9082 (N_9082,N_5075,N_6585);
nor U9083 (N_9083,N_5554,N_5638);
or U9084 (N_9084,N_5777,N_5310);
or U9085 (N_9085,N_5515,N_5637);
and U9086 (N_9086,N_5623,N_5233);
nor U9087 (N_9087,N_7210,N_5547);
or U9088 (N_9088,N_6931,N_5922);
or U9089 (N_9089,N_7247,N_5459);
nand U9090 (N_9090,N_5682,N_6998);
nor U9091 (N_9091,N_7414,N_5336);
nor U9092 (N_9092,N_5367,N_5296);
or U9093 (N_9093,N_6223,N_5225);
nor U9094 (N_9094,N_7464,N_7153);
nand U9095 (N_9095,N_6266,N_5856);
nor U9096 (N_9096,N_6954,N_5521);
or U9097 (N_9097,N_7488,N_6436);
or U9098 (N_9098,N_5866,N_6786);
or U9099 (N_9099,N_6537,N_5369);
nand U9100 (N_9100,N_6214,N_7269);
or U9101 (N_9101,N_7303,N_6399);
nor U9102 (N_9102,N_6478,N_5439);
nor U9103 (N_9103,N_6594,N_5286);
nand U9104 (N_9104,N_5961,N_7055);
nor U9105 (N_9105,N_5684,N_6020);
nand U9106 (N_9106,N_6109,N_6342);
nor U9107 (N_9107,N_5970,N_5587);
nand U9108 (N_9108,N_6718,N_6052);
and U9109 (N_9109,N_5133,N_6171);
or U9110 (N_9110,N_6071,N_5869);
and U9111 (N_9111,N_5232,N_5043);
and U9112 (N_9112,N_7243,N_6414);
nand U9113 (N_9113,N_7285,N_5198);
or U9114 (N_9114,N_6842,N_5350);
nand U9115 (N_9115,N_5186,N_6058);
nand U9116 (N_9116,N_6502,N_5405);
or U9117 (N_9117,N_5059,N_5776);
or U9118 (N_9118,N_5472,N_7068);
nand U9119 (N_9119,N_6569,N_6223);
xnor U9120 (N_9120,N_5243,N_6350);
and U9121 (N_9121,N_6543,N_5115);
nand U9122 (N_9122,N_7102,N_5093);
and U9123 (N_9123,N_5795,N_7437);
and U9124 (N_9124,N_5583,N_5063);
or U9125 (N_9125,N_6683,N_6693);
and U9126 (N_9126,N_5737,N_7326);
nor U9127 (N_9127,N_7144,N_5422);
and U9128 (N_9128,N_5831,N_7362);
nor U9129 (N_9129,N_6296,N_6297);
and U9130 (N_9130,N_5391,N_5331);
nand U9131 (N_9131,N_5581,N_5891);
or U9132 (N_9132,N_6346,N_5889);
nand U9133 (N_9133,N_5952,N_6241);
nand U9134 (N_9134,N_6773,N_5032);
nand U9135 (N_9135,N_6100,N_7188);
nand U9136 (N_9136,N_6286,N_6623);
nand U9137 (N_9137,N_6092,N_5189);
nor U9138 (N_9138,N_5904,N_7060);
and U9139 (N_9139,N_5723,N_5877);
nand U9140 (N_9140,N_5615,N_7299);
and U9141 (N_9141,N_7222,N_5506);
and U9142 (N_9142,N_5935,N_7023);
nor U9143 (N_9143,N_5515,N_7184);
nor U9144 (N_9144,N_6126,N_6781);
nand U9145 (N_9145,N_6734,N_6091);
nor U9146 (N_9146,N_6181,N_6433);
or U9147 (N_9147,N_5412,N_5751);
nor U9148 (N_9148,N_6847,N_7073);
nor U9149 (N_9149,N_6887,N_7285);
and U9150 (N_9150,N_6216,N_7232);
nor U9151 (N_9151,N_7220,N_5344);
or U9152 (N_9152,N_6395,N_5342);
or U9153 (N_9153,N_6045,N_5835);
nand U9154 (N_9154,N_5207,N_6566);
or U9155 (N_9155,N_5550,N_7027);
nor U9156 (N_9156,N_7368,N_7036);
and U9157 (N_9157,N_7481,N_6226);
and U9158 (N_9158,N_7419,N_6711);
nand U9159 (N_9159,N_5903,N_5112);
nand U9160 (N_9160,N_5502,N_5803);
or U9161 (N_9161,N_6976,N_5326);
xor U9162 (N_9162,N_5601,N_5892);
nand U9163 (N_9163,N_7232,N_5456);
nand U9164 (N_9164,N_6898,N_5447);
and U9165 (N_9165,N_6604,N_5867);
nor U9166 (N_9166,N_5890,N_6308);
and U9167 (N_9167,N_5563,N_5144);
and U9168 (N_9168,N_5190,N_7365);
nor U9169 (N_9169,N_5760,N_5736);
or U9170 (N_9170,N_6629,N_6146);
or U9171 (N_9171,N_6665,N_6834);
and U9172 (N_9172,N_6310,N_5944);
and U9173 (N_9173,N_5890,N_5976);
and U9174 (N_9174,N_6577,N_7401);
nor U9175 (N_9175,N_6036,N_6745);
nand U9176 (N_9176,N_7240,N_5411);
nor U9177 (N_9177,N_7180,N_6400);
and U9178 (N_9178,N_5338,N_6440);
nand U9179 (N_9179,N_7440,N_6520);
nor U9180 (N_9180,N_6607,N_5215);
nor U9181 (N_9181,N_6009,N_5689);
nand U9182 (N_9182,N_7097,N_5036);
and U9183 (N_9183,N_7120,N_5093);
and U9184 (N_9184,N_7401,N_6870);
or U9185 (N_9185,N_5091,N_7279);
and U9186 (N_9186,N_6405,N_7098);
or U9187 (N_9187,N_6169,N_5997);
and U9188 (N_9188,N_5560,N_6849);
and U9189 (N_9189,N_5705,N_5528);
nor U9190 (N_9190,N_5748,N_5894);
nor U9191 (N_9191,N_5868,N_6390);
nor U9192 (N_9192,N_5868,N_6479);
xnor U9193 (N_9193,N_5110,N_5605);
and U9194 (N_9194,N_6698,N_5623);
nor U9195 (N_9195,N_6740,N_7482);
or U9196 (N_9196,N_6994,N_6557);
nand U9197 (N_9197,N_6393,N_6698);
and U9198 (N_9198,N_5858,N_5157);
nand U9199 (N_9199,N_5458,N_5773);
nor U9200 (N_9200,N_5284,N_5507);
or U9201 (N_9201,N_6363,N_6750);
and U9202 (N_9202,N_6629,N_5309);
nand U9203 (N_9203,N_6545,N_5567);
and U9204 (N_9204,N_5618,N_6354);
or U9205 (N_9205,N_5975,N_6783);
and U9206 (N_9206,N_7280,N_6979);
nor U9207 (N_9207,N_6396,N_6276);
nor U9208 (N_9208,N_6691,N_5694);
nand U9209 (N_9209,N_6346,N_6380);
and U9210 (N_9210,N_6865,N_5250);
nand U9211 (N_9211,N_6646,N_6210);
and U9212 (N_9212,N_6422,N_7440);
nand U9213 (N_9213,N_6841,N_5946);
xnor U9214 (N_9214,N_6437,N_7124);
nand U9215 (N_9215,N_6507,N_7429);
and U9216 (N_9216,N_5754,N_6193);
nor U9217 (N_9217,N_7234,N_5199);
or U9218 (N_9218,N_6745,N_7149);
and U9219 (N_9219,N_5550,N_6121);
nand U9220 (N_9220,N_5082,N_6351);
nand U9221 (N_9221,N_5464,N_6402);
and U9222 (N_9222,N_6688,N_5358);
or U9223 (N_9223,N_5441,N_6857);
or U9224 (N_9224,N_6555,N_5562);
nor U9225 (N_9225,N_6756,N_6291);
and U9226 (N_9226,N_6943,N_5143);
nor U9227 (N_9227,N_5473,N_7074);
and U9228 (N_9228,N_5590,N_7183);
or U9229 (N_9229,N_5947,N_5326);
nand U9230 (N_9230,N_5603,N_6511);
or U9231 (N_9231,N_6311,N_5677);
nand U9232 (N_9232,N_6608,N_5840);
nand U9233 (N_9233,N_7450,N_6272);
or U9234 (N_9234,N_5944,N_6613);
nor U9235 (N_9235,N_5557,N_6673);
and U9236 (N_9236,N_5163,N_6127);
nor U9237 (N_9237,N_5915,N_6745);
nand U9238 (N_9238,N_6585,N_7475);
nor U9239 (N_9239,N_6033,N_6830);
nor U9240 (N_9240,N_5986,N_5434);
and U9241 (N_9241,N_6441,N_5944);
nor U9242 (N_9242,N_5346,N_5218);
or U9243 (N_9243,N_5982,N_5600);
and U9244 (N_9244,N_5589,N_7081);
and U9245 (N_9245,N_5051,N_6738);
or U9246 (N_9246,N_7008,N_6281);
and U9247 (N_9247,N_5452,N_5303);
nor U9248 (N_9248,N_6805,N_7234);
nand U9249 (N_9249,N_6641,N_6848);
or U9250 (N_9250,N_6927,N_5362);
xor U9251 (N_9251,N_6570,N_6322);
nor U9252 (N_9252,N_5255,N_5844);
nand U9253 (N_9253,N_6870,N_5232);
nor U9254 (N_9254,N_7244,N_5114);
or U9255 (N_9255,N_5615,N_6610);
nor U9256 (N_9256,N_6598,N_5955);
nand U9257 (N_9257,N_5366,N_5987);
or U9258 (N_9258,N_6368,N_6821);
xor U9259 (N_9259,N_6220,N_7382);
or U9260 (N_9260,N_6422,N_5053);
nor U9261 (N_9261,N_6422,N_7449);
nor U9262 (N_9262,N_7047,N_5365);
and U9263 (N_9263,N_7405,N_6006);
nand U9264 (N_9264,N_5569,N_6662);
and U9265 (N_9265,N_6541,N_6469);
or U9266 (N_9266,N_7035,N_6677);
and U9267 (N_9267,N_6981,N_6189);
or U9268 (N_9268,N_6475,N_6974);
or U9269 (N_9269,N_6309,N_6628);
nand U9270 (N_9270,N_7125,N_5122);
nor U9271 (N_9271,N_5026,N_7158);
nand U9272 (N_9272,N_5749,N_6402);
or U9273 (N_9273,N_6804,N_6091);
or U9274 (N_9274,N_6834,N_6080);
nand U9275 (N_9275,N_7464,N_6367);
or U9276 (N_9276,N_5613,N_6999);
nor U9277 (N_9277,N_5952,N_7367);
nor U9278 (N_9278,N_7236,N_6516);
or U9279 (N_9279,N_6825,N_7454);
or U9280 (N_9280,N_6589,N_7495);
or U9281 (N_9281,N_5138,N_6581);
nor U9282 (N_9282,N_5499,N_6941);
nand U9283 (N_9283,N_6557,N_5079);
or U9284 (N_9284,N_5554,N_6292);
and U9285 (N_9285,N_5060,N_5570);
and U9286 (N_9286,N_6731,N_5988);
or U9287 (N_9287,N_7205,N_5815);
nor U9288 (N_9288,N_6359,N_6226);
nand U9289 (N_9289,N_5631,N_6413);
nand U9290 (N_9290,N_6019,N_6579);
nor U9291 (N_9291,N_5036,N_5293);
and U9292 (N_9292,N_6066,N_6193);
and U9293 (N_9293,N_5993,N_6438);
nand U9294 (N_9294,N_5766,N_5246);
or U9295 (N_9295,N_6390,N_5375);
and U9296 (N_9296,N_5173,N_7088);
nand U9297 (N_9297,N_6550,N_6398);
and U9298 (N_9298,N_5124,N_6840);
or U9299 (N_9299,N_6521,N_5327);
or U9300 (N_9300,N_7487,N_6926);
nand U9301 (N_9301,N_7461,N_6092);
nand U9302 (N_9302,N_6884,N_6795);
and U9303 (N_9303,N_6715,N_6554);
nand U9304 (N_9304,N_7260,N_5629);
and U9305 (N_9305,N_5490,N_6972);
nor U9306 (N_9306,N_6278,N_7489);
nand U9307 (N_9307,N_6164,N_6338);
nor U9308 (N_9308,N_6111,N_7106);
nand U9309 (N_9309,N_6331,N_6199);
nand U9310 (N_9310,N_6669,N_6285);
or U9311 (N_9311,N_6303,N_6044);
or U9312 (N_9312,N_6697,N_7097);
or U9313 (N_9313,N_5438,N_5548);
or U9314 (N_9314,N_6389,N_6463);
nor U9315 (N_9315,N_5351,N_5560);
or U9316 (N_9316,N_5134,N_6916);
nor U9317 (N_9317,N_5634,N_6563);
nor U9318 (N_9318,N_5940,N_6687);
and U9319 (N_9319,N_6113,N_5347);
nor U9320 (N_9320,N_5653,N_6000);
nand U9321 (N_9321,N_5192,N_6423);
or U9322 (N_9322,N_5039,N_7369);
or U9323 (N_9323,N_7316,N_5724);
nand U9324 (N_9324,N_7415,N_7346);
nor U9325 (N_9325,N_5552,N_7298);
and U9326 (N_9326,N_5096,N_5905);
and U9327 (N_9327,N_6623,N_5565);
nor U9328 (N_9328,N_5793,N_7405);
nor U9329 (N_9329,N_7018,N_5723);
nand U9330 (N_9330,N_7436,N_5366);
and U9331 (N_9331,N_5025,N_5234);
and U9332 (N_9332,N_5589,N_5421);
or U9333 (N_9333,N_5026,N_7425);
or U9334 (N_9334,N_7027,N_5069);
or U9335 (N_9335,N_7363,N_7284);
and U9336 (N_9336,N_6100,N_7270);
and U9337 (N_9337,N_6518,N_6928);
or U9338 (N_9338,N_5264,N_7339);
and U9339 (N_9339,N_6470,N_5187);
nor U9340 (N_9340,N_7317,N_5815);
or U9341 (N_9341,N_7479,N_5604);
and U9342 (N_9342,N_6389,N_6327);
nor U9343 (N_9343,N_7144,N_6955);
nor U9344 (N_9344,N_7015,N_6037);
xor U9345 (N_9345,N_5754,N_7278);
and U9346 (N_9346,N_7435,N_7111);
nor U9347 (N_9347,N_6322,N_6533);
nand U9348 (N_9348,N_6594,N_6147);
nor U9349 (N_9349,N_7398,N_6226);
or U9350 (N_9350,N_6880,N_6899);
nand U9351 (N_9351,N_6406,N_6772);
or U9352 (N_9352,N_5628,N_6328);
and U9353 (N_9353,N_6664,N_6213);
nor U9354 (N_9354,N_6692,N_6017);
and U9355 (N_9355,N_6723,N_5988);
or U9356 (N_9356,N_6814,N_5725);
nor U9357 (N_9357,N_5441,N_6956);
and U9358 (N_9358,N_5639,N_5096);
and U9359 (N_9359,N_6273,N_5266);
nor U9360 (N_9360,N_6340,N_5605);
and U9361 (N_9361,N_5552,N_5950);
or U9362 (N_9362,N_5777,N_6124);
nor U9363 (N_9363,N_6227,N_5037);
and U9364 (N_9364,N_5844,N_6937);
nand U9365 (N_9365,N_6474,N_7425);
nand U9366 (N_9366,N_5492,N_5164);
nand U9367 (N_9367,N_7231,N_7156);
nor U9368 (N_9368,N_5585,N_5215);
or U9369 (N_9369,N_5914,N_5722);
or U9370 (N_9370,N_6024,N_6119);
or U9371 (N_9371,N_5143,N_7072);
and U9372 (N_9372,N_6792,N_7376);
nand U9373 (N_9373,N_7203,N_5698);
xnor U9374 (N_9374,N_7189,N_5028);
nor U9375 (N_9375,N_5306,N_5084);
or U9376 (N_9376,N_5064,N_6432);
nand U9377 (N_9377,N_6700,N_7198);
or U9378 (N_9378,N_7261,N_6226);
and U9379 (N_9379,N_6903,N_5193);
or U9380 (N_9380,N_5550,N_5220);
and U9381 (N_9381,N_5987,N_7406);
or U9382 (N_9382,N_6266,N_5904);
nand U9383 (N_9383,N_5432,N_7434);
or U9384 (N_9384,N_5113,N_5780);
nand U9385 (N_9385,N_6966,N_5803);
nor U9386 (N_9386,N_7074,N_5754);
or U9387 (N_9387,N_6333,N_6760);
nand U9388 (N_9388,N_6310,N_6998);
nor U9389 (N_9389,N_5614,N_5374);
nand U9390 (N_9390,N_5287,N_6989);
nand U9391 (N_9391,N_6004,N_5853);
xnor U9392 (N_9392,N_5177,N_6814);
and U9393 (N_9393,N_6447,N_6127);
and U9394 (N_9394,N_6411,N_6789);
nand U9395 (N_9395,N_6075,N_5766);
nand U9396 (N_9396,N_6099,N_6057);
nand U9397 (N_9397,N_5824,N_6513);
nand U9398 (N_9398,N_7202,N_5759);
or U9399 (N_9399,N_6780,N_6421);
nand U9400 (N_9400,N_6969,N_6506);
nor U9401 (N_9401,N_6400,N_6370);
or U9402 (N_9402,N_5705,N_5749);
and U9403 (N_9403,N_6937,N_6685);
or U9404 (N_9404,N_5608,N_5312);
nand U9405 (N_9405,N_5697,N_6545);
or U9406 (N_9406,N_5897,N_5154);
or U9407 (N_9407,N_6090,N_6737);
nor U9408 (N_9408,N_7381,N_5208);
nand U9409 (N_9409,N_5607,N_7118);
and U9410 (N_9410,N_5360,N_5710);
and U9411 (N_9411,N_6112,N_6340);
or U9412 (N_9412,N_5913,N_5934);
nand U9413 (N_9413,N_6431,N_5768);
and U9414 (N_9414,N_5740,N_5942);
or U9415 (N_9415,N_6582,N_5623);
nand U9416 (N_9416,N_6632,N_6806);
or U9417 (N_9417,N_6819,N_7242);
nor U9418 (N_9418,N_5297,N_6795);
or U9419 (N_9419,N_6839,N_7232);
nor U9420 (N_9420,N_5247,N_7390);
nand U9421 (N_9421,N_6241,N_7078);
nand U9422 (N_9422,N_5478,N_5099);
nor U9423 (N_9423,N_6139,N_7169);
nand U9424 (N_9424,N_5783,N_5207);
and U9425 (N_9425,N_5387,N_5121);
nand U9426 (N_9426,N_6558,N_6599);
nor U9427 (N_9427,N_5504,N_6769);
nand U9428 (N_9428,N_6951,N_6239);
and U9429 (N_9429,N_5917,N_5139);
or U9430 (N_9430,N_6462,N_5594);
nand U9431 (N_9431,N_6285,N_5648);
and U9432 (N_9432,N_6739,N_5735);
and U9433 (N_9433,N_5948,N_5739);
nand U9434 (N_9434,N_6743,N_6829);
and U9435 (N_9435,N_7067,N_7159);
nor U9436 (N_9436,N_5323,N_6775);
or U9437 (N_9437,N_5565,N_6235);
nor U9438 (N_9438,N_7374,N_5579);
or U9439 (N_9439,N_7082,N_7158);
nand U9440 (N_9440,N_5446,N_6335);
and U9441 (N_9441,N_6538,N_6750);
nor U9442 (N_9442,N_7109,N_5107);
or U9443 (N_9443,N_6886,N_7384);
nand U9444 (N_9444,N_6602,N_6184);
nor U9445 (N_9445,N_6794,N_5663);
or U9446 (N_9446,N_5707,N_5695);
nand U9447 (N_9447,N_5973,N_6227);
or U9448 (N_9448,N_6586,N_5388);
nand U9449 (N_9449,N_5910,N_7424);
or U9450 (N_9450,N_6866,N_6988);
xor U9451 (N_9451,N_5097,N_5316);
and U9452 (N_9452,N_6264,N_5730);
or U9453 (N_9453,N_6600,N_5959);
and U9454 (N_9454,N_6137,N_5997);
or U9455 (N_9455,N_6353,N_5205);
nand U9456 (N_9456,N_5156,N_6082);
nor U9457 (N_9457,N_5739,N_5562);
nor U9458 (N_9458,N_7004,N_7330);
or U9459 (N_9459,N_6883,N_6870);
xnor U9460 (N_9460,N_6485,N_5582);
nand U9461 (N_9461,N_5211,N_5719);
and U9462 (N_9462,N_5569,N_6865);
and U9463 (N_9463,N_7411,N_6909);
or U9464 (N_9464,N_6181,N_5963);
and U9465 (N_9465,N_5953,N_5310);
and U9466 (N_9466,N_5798,N_6224);
nand U9467 (N_9467,N_6779,N_5498);
nand U9468 (N_9468,N_7046,N_7064);
and U9469 (N_9469,N_5676,N_5242);
and U9470 (N_9470,N_5474,N_5736);
and U9471 (N_9471,N_7211,N_7338);
nor U9472 (N_9472,N_5542,N_5576);
and U9473 (N_9473,N_6662,N_5205);
and U9474 (N_9474,N_5171,N_6170);
nand U9475 (N_9475,N_6175,N_7286);
and U9476 (N_9476,N_6189,N_5761);
nand U9477 (N_9477,N_6435,N_5170);
and U9478 (N_9478,N_5147,N_6438);
nor U9479 (N_9479,N_5718,N_5102);
or U9480 (N_9480,N_6450,N_7019);
nor U9481 (N_9481,N_6432,N_6289);
or U9482 (N_9482,N_6426,N_7022);
or U9483 (N_9483,N_7114,N_7481);
and U9484 (N_9484,N_6156,N_5776);
nor U9485 (N_9485,N_6687,N_6961);
or U9486 (N_9486,N_6064,N_6421);
or U9487 (N_9487,N_5979,N_6150);
and U9488 (N_9488,N_6340,N_6680);
nor U9489 (N_9489,N_5459,N_5314);
and U9490 (N_9490,N_6998,N_6542);
nand U9491 (N_9491,N_6760,N_5561);
nand U9492 (N_9492,N_7102,N_5716);
and U9493 (N_9493,N_5303,N_6788);
or U9494 (N_9494,N_5845,N_5730);
nor U9495 (N_9495,N_5822,N_6649);
nand U9496 (N_9496,N_5462,N_5924);
and U9497 (N_9497,N_5990,N_6715);
nand U9498 (N_9498,N_5806,N_6617);
nand U9499 (N_9499,N_6208,N_5341);
or U9500 (N_9500,N_6429,N_5152);
nand U9501 (N_9501,N_5661,N_5818);
or U9502 (N_9502,N_6749,N_6795);
or U9503 (N_9503,N_7414,N_7426);
nand U9504 (N_9504,N_7317,N_7143);
or U9505 (N_9505,N_6396,N_5471);
nand U9506 (N_9506,N_7480,N_6877);
nand U9507 (N_9507,N_5958,N_5784);
or U9508 (N_9508,N_5635,N_5493);
or U9509 (N_9509,N_5092,N_5422);
nand U9510 (N_9510,N_5969,N_7034);
nor U9511 (N_9511,N_7427,N_7415);
or U9512 (N_9512,N_6255,N_5735);
and U9513 (N_9513,N_6753,N_6098);
nand U9514 (N_9514,N_5023,N_5444);
nor U9515 (N_9515,N_6524,N_7385);
nor U9516 (N_9516,N_5422,N_5163);
and U9517 (N_9517,N_6628,N_6005);
nand U9518 (N_9518,N_5419,N_5958);
and U9519 (N_9519,N_5450,N_5263);
nand U9520 (N_9520,N_5671,N_5084);
nand U9521 (N_9521,N_6105,N_7316);
nor U9522 (N_9522,N_7288,N_5746);
xnor U9523 (N_9523,N_6148,N_6606);
nand U9524 (N_9524,N_6814,N_5566);
nand U9525 (N_9525,N_7230,N_7132);
nor U9526 (N_9526,N_6865,N_7204);
and U9527 (N_9527,N_7385,N_7361);
nand U9528 (N_9528,N_6208,N_6098);
or U9529 (N_9529,N_7199,N_6368);
nand U9530 (N_9530,N_5680,N_5316);
and U9531 (N_9531,N_5705,N_5930);
and U9532 (N_9532,N_7040,N_6739);
nor U9533 (N_9533,N_6893,N_5988);
and U9534 (N_9534,N_5899,N_6232);
nor U9535 (N_9535,N_5688,N_5595);
nor U9536 (N_9536,N_6588,N_6739);
nand U9537 (N_9537,N_5578,N_5412);
or U9538 (N_9538,N_5896,N_5604);
and U9539 (N_9539,N_6683,N_5191);
or U9540 (N_9540,N_5529,N_6326);
and U9541 (N_9541,N_6137,N_6909);
and U9542 (N_9542,N_5415,N_6412);
or U9543 (N_9543,N_6026,N_6002);
nor U9544 (N_9544,N_5662,N_6366);
and U9545 (N_9545,N_5619,N_7017);
or U9546 (N_9546,N_5065,N_6747);
nor U9547 (N_9547,N_6437,N_5934);
and U9548 (N_9548,N_6512,N_7229);
and U9549 (N_9549,N_6735,N_6834);
and U9550 (N_9550,N_6796,N_5665);
nor U9551 (N_9551,N_5230,N_5088);
and U9552 (N_9552,N_5914,N_5216);
nor U9553 (N_9553,N_6970,N_6178);
and U9554 (N_9554,N_5163,N_5401);
nor U9555 (N_9555,N_7453,N_6657);
nor U9556 (N_9556,N_6293,N_6076);
nor U9557 (N_9557,N_5619,N_5741);
and U9558 (N_9558,N_6410,N_7076);
and U9559 (N_9559,N_7106,N_6339);
and U9560 (N_9560,N_5515,N_5890);
or U9561 (N_9561,N_6918,N_5327);
nor U9562 (N_9562,N_6547,N_7091);
or U9563 (N_9563,N_7360,N_5844);
nand U9564 (N_9564,N_7330,N_6299);
or U9565 (N_9565,N_5428,N_6107);
nand U9566 (N_9566,N_6601,N_7292);
nor U9567 (N_9567,N_7413,N_5660);
nor U9568 (N_9568,N_6199,N_6113);
nor U9569 (N_9569,N_6520,N_6098);
or U9570 (N_9570,N_6219,N_7443);
nor U9571 (N_9571,N_6306,N_7337);
nand U9572 (N_9572,N_6647,N_5292);
nor U9573 (N_9573,N_6247,N_6144);
nand U9574 (N_9574,N_5884,N_7176);
nand U9575 (N_9575,N_5366,N_5372);
and U9576 (N_9576,N_5098,N_5279);
or U9577 (N_9577,N_6750,N_6021);
or U9578 (N_9578,N_7070,N_6893);
and U9579 (N_9579,N_6430,N_7062);
and U9580 (N_9580,N_5327,N_5341);
or U9581 (N_9581,N_7246,N_6007);
and U9582 (N_9582,N_6048,N_5151);
or U9583 (N_9583,N_7238,N_6620);
or U9584 (N_9584,N_6104,N_5676);
nor U9585 (N_9585,N_6039,N_5936);
or U9586 (N_9586,N_5319,N_5852);
nor U9587 (N_9587,N_6782,N_6211);
and U9588 (N_9588,N_5588,N_5208);
or U9589 (N_9589,N_7181,N_5643);
or U9590 (N_9590,N_6069,N_7493);
and U9591 (N_9591,N_7375,N_7436);
nand U9592 (N_9592,N_6880,N_6929);
or U9593 (N_9593,N_5561,N_7105);
and U9594 (N_9594,N_6560,N_5170);
nand U9595 (N_9595,N_7385,N_5177);
nor U9596 (N_9596,N_5530,N_6057);
and U9597 (N_9597,N_6497,N_5594);
or U9598 (N_9598,N_5033,N_6640);
or U9599 (N_9599,N_7278,N_5805);
nand U9600 (N_9600,N_6721,N_6629);
nor U9601 (N_9601,N_7127,N_6900);
or U9602 (N_9602,N_5886,N_5702);
xor U9603 (N_9603,N_5078,N_7461);
nand U9604 (N_9604,N_6435,N_6193);
nor U9605 (N_9605,N_6284,N_6724);
and U9606 (N_9606,N_6421,N_6762);
xor U9607 (N_9607,N_6003,N_5641);
nand U9608 (N_9608,N_5866,N_7496);
nand U9609 (N_9609,N_5706,N_6282);
or U9610 (N_9610,N_5968,N_7349);
nand U9611 (N_9611,N_7474,N_7245);
or U9612 (N_9612,N_7247,N_6062);
and U9613 (N_9613,N_7404,N_6336);
nor U9614 (N_9614,N_5634,N_5286);
nand U9615 (N_9615,N_5651,N_5068);
and U9616 (N_9616,N_5641,N_5659);
nor U9617 (N_9617,N_7099,N_6520);
and U9618 (N_9618,N_5968,N_5958);
and U9619 (N_9619,N_7050,N_7145);
nor U9620 (N_9620,N_7208,N_5095);
and U9621 (N_9621,N_5403,N_6463);
or U9622 (N_9622,N_6674,N_6513);
or U9623 (N_9623,N_5929,N_5396);
nand U9624 (N_9624,N_7057,N_6805);
nor U9625 (N_9625,N_7016,N_6087);
nand U9626 (N_9626,N_5233,N_5169);
or U9627 (N_9627,N_6669,N_7015);
nor U9628 (N_9628,N_5176,N_5173);
or U9629 (N_9629,N_6770,N_5723);
or U9630 (N_9630,N_5815,N_6283);
and U9631 (N_9631,N_6989,N_6720);
and U9632 (N_9632,N_7381,N_7337);
and U9633 (N_9633,N_6738,N_5209);
and U9634 (N_9634,N_5611,N_5698);
nor U9635 (N_9635,N_5111,N_5827);
or U9636 (N_9636,N_6765,N_5467);
nand U9637 (N_9637,N_6872,N_6005);
nor U9638 (N_9638,N_5965,N_7428);
or U9639 (N_9639,N_5225,N_5989);
nor U9640 (N_9640,N_6205,N_7427);
nand U9641 (N_9641,N_6945,N_7227);
nor U9642 (N_9642,N_5396,N_5891);
nor U9643 (N_9643,N_5742,N_5052);
or U9644 (N_9644,N_6531,N_5950);
and U9645 (N_9645,N_7121,N_7265);
nand U9646 (N_9646,N_5539,N_5140);
and U9647 (N_9647,N_5538,N_5336);
or U9648 (N_9648,N_6803,N_6283);
and U9649 (N_9649,N_6113,N_6723);
or U9650 (N_9650,N_6442,N_5187);
or U9651 (N_9651,N_5245,N_7319);
nand U9652 (N_9652,N_7121,N_5805);
nor U9653 (N_9653,N_6210,N_5906);
nor U9654 (N_9654,N_6477,N_5512);
and U9655 (N_9655,N_6002,N_5011);
or U9656 (N_9656,N_5876,N_5074);
or U9657 (N_9657,N_5309,N_5587);
nor U9658 (N_9658,N_6130,N_7239);
and U9659 (N_9659,N_6912,N_7085);
nor U9660 (N_9660,N_6338,N_6367);
xor U9661 (N_9661,N_7184,N_5063);
nand U9662 (N_9662,N_5850,N_5552);
nand U9663 (N_9663,N_6739,N_6794);
or U9664 (N_9664,N_5340,N_5130);
nand U9665 (N_9665,N_6028,N_6911);
nand U9666 (N_9666,N_5625,N_5798);
nor U9667 (N_9667,N_5086,N_6860);
and U9668 (N_9668,N_5862,N_6608);
nand U9669 (N_9669,N_7008,N_5604);
nor U9670 (N_9670,N_7129,N_7253);
or U9671 (N_9671,N_6980,N_7390);
and U9672 (N_9672,N_7410,N_5114);
and U9673 (N_9673,N_6010,N_5609);
xor U9674 (N_9674,N_5625,N_6264);
nor U9675 (N_9675,N_6916,N_5775);
nand U9676 (N_9676,N_6282,N_6710);
and U9677 (N_9677,N_7081,N_6275);
nand U9678 (N_9678,N_7261,N_7208);
or U9679 (N_9679,N_6083,N_5366);
and U9680 (N_9680,N_5355,N_5670);
or U9681 (N_9681,N_6988,N_5921);
nor U9682 (N_9682,N_7266,N_5929);
nor U9683 (N_9683,N_7325,N_5747);
nand U9684 (N_9684,N_5946,N_6313);
nand U9685 (N_9685,N_6379,N_6095);
and U9686 (N_9686,N_6098,N_5665);
and U9687 (N_9687,N_5865,N_5517);
and U9688 (N_9688,N_6356,N_5224);
nand U9689 (N_9689,N_5108,N_6752);
nor U9690 (N_9690,N_6821,N_6594);
nor U9691 (N_9691,N_7470,N_5440);
nand U9692 (N_9692,N_5538,N_7354);
or U9693 (N_9693,N_5161,N_5582);
and U9694 (N_9694,N_5731,N_6355);
or U9695 (N_9695,N_5741,N_6732);
nand U9696 (N_9696,N_6630,N_7455);
and U9697 (N_9697,N_5745,N_6092);
nand U9698 (N_9698,N_5676,N_5996);
and U9699 (N_9699,N_5620,N_5927);
nand U9700 (N_9700,N_5401,N_5824);
nor U9701 (N_9701,N_6017,N_6636);
or U9702 (N_9702,N_7217,N_5928);
or U9703 (N_9703,N_6200,N_5125);
nand U9704 (N_9704,N_6540,N_7147);
and U9705 (N_9705,N_5387,N_5815);
or U9706 (N_9706,N_7360,N_6995);
nor U9707 (N_9707,N_5396,N_5990);
nand U9708 (N_9708,N_5392,N_5434);
nor U9709 (N_9709,N_5521,N_6431);
or U9710 (N_9710,N_5006,N_7486);
nand U9711 (N_9711,N_6633,N_5148);
and U9712 (N_9712,N_6500,N_5014);
and U9713 (N_9713,N_5741,N_5867);
and U9714 (N_9714,N_5717,N_6115);
nor U9715 (N_9715,N_5375,N_5500);
and U9716 (N_9716,N_6857,N_6401);
nor U9717 (N_9717,N_6154,N_5419);
nor U9718 (N_9718,N_5010,N_6128);
nor U9719 (N_9719,N_6958,N_7398);
nand U9720 (N_9720,N_5300,N_6152);
and U9721 (N_9721,N_6229,N_6518);
nand U9722 (N_9722,N_6424,N_7172);
nand U9723 (N_9723,N_6525,N_6483);
nor U9724 (N_9724,N_5448,N_5462);
nand U9725 (N_9725,N_5426,N_6134);
nand U9726 (N_9726,N_5568,N_5908);
nand U9727 (N_9727,N_5048,N_6112);
and U9728 (N_9728,N_5438,N_6485);
nor U9729 (N_9729,N_5401,N_5496);
nor U9730 (N_9730,N_6919,N_5048);
nor U9731 (N_9731,N_6890,N_6638);
nor U9732 (N_9732,N_5144,N_5536);
nor U9733 (N_9733,N_7121,N_7041);
and U9734 (N_9734,N_7253,N_7123);
and U9735 (N_9735,N_6968,N_7046);
nand U9736 (N_9736,N_7185,N_6657);
nor U9737 (N_9737,N_7172,N_5851);
and U9738 (N_9738,N_5365,N_6061);
nand U9739 (N_9739,N_5522,N_5560);
nand U9740 (N_9740,N_6774,N_6794);
and U9741 (N_9741,N_7497,N_6570);
nand U9742 (N_9742,N_6547,N_5250);
nand U9743 (N_9743,N_6413,N_6737);
or U9744 (N_9744,N_6713,N_6285);
nor U9745 (N_9745,N_5301,N_5750);
nor U9746 (N_9746,N_5899,N_5853);
nand U9747 (N_9747,N_6950,N_7345);
and U9748 (N_9748,N_5334,N_5721);
nand U9749 (N_9749,N_5157,N_5153);
and U9750 (N_9750,N_6811,N_6263);
nand U9751 (N_9751,N_5871,N_6918);
and U9752 (N_9752,N_5301,N_6667);
or U9753 (N_9753,N_6185,N_5101);
or U9754 (N_9754,N_7156,N_7422);
nor U9755 (N_9755,N_5623,N_6305);
or U9756 (N_9756,N_7094,N_5119);
nand U9757 (N_9757,N_6236,N_6639);
and U9758 (N_9758,N_7266,N_6720);
nand U9759 (N_9759,N_6573,N_7303);
or U9760 (N_9760,N_5932,N_6925);
or U9761 (N_9761,N_5176,N_7453);
nor U9762 (N_9762,N_5833,N_6508);
and U9763 (N_9763,N_6724,N_7275);
or U9764 (N_9764,N_6261,N_6088);
nand U9765 (N_9765,N_5671,N_5872);
nor U9766 (N_9766,N_6500,N_5204);
and U9767 (N_9767,N_6254,N_5859);
or U9768 (N_9768,N_5178,N_7226);
nor U9769 (N_9769,N_6214,N_6840);
and U9770 (N_9770,N_6102,N_7154);
and U9771 (N_9771,N_5953,N_5403);
or U9772 (N_9772,N_5813,N_7029);
nor U9773 (N_9773,N_6160,N_6158);
and U9774 (N_9774,N_6439,N_6411);
nand U9775 (N_9775,N_6968,N_7179);
nand U9776 (N_9776,N_7233,N_6889);
or U9777 (N_9777,N_5543,N_5388);
nand U9778 (N_9778,N_5424,N_5511);
and U9779 (N_9779,N_6499,N_6615);
nand U9780 (N_9780,N_6005,N_5315);
nand U9781 (N_9781,N_6277,N_5163);
or U9782 (N_9782,N_5894,N_6594);
and U9783 (N_9783,N_7462,N_6504);
and U9784 (N_9784,N_6826,N_7352);
and U9785 (N_9785,N_6872,N_6508);
or U9786 (N_9786,N_5021,N_5859);
nor U9787 (N_9787,N_5346,N_5546);
nor U9788 (N_9788,N_6844,N_6423);
and U9789 (N_9789,N_5987,N_6318);
or U9790 (N_9790,N_7273,N_6517);
nand U9791 (N_9791,N_6864,N_6315);
nand U9792 (N_9792,N_5253,N_6995);
nand U9793 (N_9793,N_6851,N_5932);
and U9794 (N_9794,N_5840,N_5638);
nor U9795 (N_9795,N_6136,N_6399);
or U9796 (N_9796,N_7323,N_5762);
nor U9797 (N_9797,N_7153,N_5865);
or U9798 (N_9798,N_5853,N_6275);
nor U9799 (N_9799,N_5652,N_6068);
nor U9800 (N_9800,N_5193,N_6238);
nand U9801 (N_9801,N_5062,N_7058);
nor U9802 (N_9802,N_5340,N_6551);
nor U9803 (N_9803,N_6366,N_5541);
or U9804 (N_9804,N_7433,N_6292);
and U9805 (N_9805,N_5938,N_6703);
or U9806 (N_9806,N_6226,N_7227);
xnor U9807 (N_9807,N_6569,N_5000);
or U9808 (N_9808,N_5165,N_7012);
nand U9809 (N_9809,N_5232,N_5138);
nor U9810 (N_9810,N_7222,N_6188);
nor U9811 (N_9811,N_5474,N_6619);
nor U9812 (N_9812,N_6532,N_5693);
or U9813 (N_9813,N_6518,N_5289);
nor U9814 (N_9814,N_5033,N_6251);
nand U9815 (N_9815,N_7107,N_6602);
nand U9816 (N_9816,N_7345,N_6076);
and U9817 (N_9817,N_7324,N_6658);
or U9818 (N_9818,N_6251,N_5457);
nor U9819 (N_9819,N_5722,N_5756);
and U9820 (N_9820,N_7440,N_5791);
nand U9821 (N_9821,N_6963,N_6844);
nor U9822 (N_9822,N_6205,N_5683);
nor U9823 (N_9823,N_6872,N_5292);
and U9824 (N_9824,N_6225,N_7107);
or U9825 (N_9825,N_6734,N_7439);
nor U9826 (N_9826,N_7177,N_5547);
nor U9827 (N_9827,N_7004,N_6635);
and U9828 (N_9828,N_5872,N_5514);
and U9829 (N_9829,N_6653,N_7019);
nor U9830 (N_9830,N_5089,N_7481);
or U9831 (N_9831,N_5550,N_6478);
nor U9832 (N_9832,N_5078,N_6325);
or U9833 (N_9833,N_6113,N_6233);
nor U9834 (N_9834,N_5190,N_5638);
or U9835 (N_9835,N_5498,N_7190);
and U9836 (N_9836,N_6787,N_6748);
or U9837 (N_9837,N_5194,N_6886);
nor U9838 (N_9838,N_5212,N_5724);
or U9839 (N_9839,N_7415,N_5605);
nor U9840 (N_9840,N_7142,N_7225);
nor U9841 (N_9841,N_6731,N_5215);
and U9842 (N_9842,N_6549,N_5810);
or U9843 (N_9843,N_7484,N_6001);
and U9844 (N_9844,N_7090,N_5086);
nor U9845 (N_9845,N_6219,N_6993);
or U9846 (N_9846,N_6069,N_5180);
and U9847 (N_9847,N_6888,N_7123);
nand U9848 (N_9848,N_6388,N_5694);
nor U9849 (N_9849,N_5760,N_7057);
xnor U9850 (N_9850,N_6192,N_6274);
or U9851 (N_9851,N_6491,N_5117);
or U9852 (N_9852,N_6950,N_5606);
nor U9853 (N_9853,N_6975,N_6373);
or U9854 (N_9854,N_7114,N_6973);
nor U9855 (N_9855,N_6406,N_7320);
and U9856 (N_9856,N_5233,N_6044);
nand U9857 (N_9857,N_6250,N_5526);
nand U9858 (N_9858,N_5558,N_6957);
nor U9859 (N_9859,N_5973,N_5061);
or U9860 (N_9860,N_5478,N_6021);
nand U9861 (N_9861,N_7401,N_5250);
and U9862 (N_9862,N_6938,N_6903);
nor U9863 (N_9863,N_5768,N_5797);
nor U9864 (N_9864,N_6989,N_5048);
nand U9865 (N_9865,N_6407,N_7265);
nand U9866 (N_9866,N_5709,N_5606);
nor U9867 (N_9867,N_5794,N_6065);
or U9868 (N_9868,N_5444,N_7423);
and U9869 (N_9869,N_6510,N_6919);
nand U9870 (N_9870,N_7224,N_5194);
nor U9871 (N_9871,N_5001,N_5654);
nor U9872 (N_9872,N_6010,N_6273);
or U9873 (N_9873,N_6316,N_6647);
and U9874 (N_9874,N_5022,N_5933);
nand U9875 (N_9875,N_5144,N_6088);
and U9876 (N_9876,N_6355,N_6787);
nor U9877 (N_9877,N_6531,N_7254);
nand U9878 (N_9878,N_6853,N_6833);
and U9879 (N_9879,N_5190,N_5161);
nor U9880 (N_9880,N_5460,N_6968);
and U9881 (N_9881,N_6718,N_6608);
and U9882 (N_9882,N_6787,N_6536);
nand U9883 (N_9883,N_5632,N_7038);
or U9884 (N_9884,N_5082,N_6761);
nor U9885 (N_9885,N_6798,N_7465);
or U9886 (N_9886,N_6808,N_5353);
or U9887 (N_9887,N_6727,N_7435);
nand U9888 (N_9888,N_5589,N_5707);
and U9889 (N_9889,N_6961,N_6564);
or U9890 (N_9890,N_5650,N_6106);
nor U9891 (N_9891,N_6150,N_6282);
and U9892 (N_9892,N_6897,N_5681);
and U9893 (N_9893,N_6478,N_5130);
or U9894 (N_9894,N_5365,N_7031);
nand U9895 (N_9895,N_6768,N_7159);
nand U9896 (N_9896,N_6312,N_5978);
nand U9897 (N_9897,N_5511,N_5643);
and U9898 (N_9898,N_5108,N_7466);
or U9899 (N_9899,N_6539,N_7356);
or U9900 (N_9900,N_5460,N_7387);
and U9901 (N_9901,N_7137,N_5498);
nand U9902 (N_9902,N_5232,N_5309);
nor U9903 (N_9903,N_6331,N_6332);
nand U9904 (N_9904,N_5970,N_6921);
or U9905 (N_9905,N_7360,N_7211);
or U9906 (N_9906,N_6267,N_6811);
and U9907 (N_9907,N_6292,N_7001);
and U9908 (N_9908,N_7024,N_5303);
nor U9909 (N_9909,N_6679,N_5160);
and U9910 (N_9910,N_6942,N_7139);
or U9911 (N_9911,N_5875,N_5559);
or U9912 (N_9912,N_5522,N_5633);
nor U9913 (N_9913,N_5238,N_6828);
and U9914 (N_9914,N_6508,N_5412);
or U9915 (N_9915,N_5553,N_7496);
nand U9916 (N_9916,N_7401,N_5569);
or U9917 (N_9917,N_5925,N_6834);
and U9918 (N_9918,N_5037,N_6538);
nor U9919 (N_9919,N_6567,N_6527);
nand U9920 (N_9920,N_5769,N_6177);
or U9921 (N_9921,N_6418,N_5443);
nor U9922 (N_9922,N_5238,N_5751);
and U9923 (N_9923,N_6521,N_7207);
nand U9924 (N_9924,N_5033,N_6257);
and U9925 (N_9925,N_5158,N_5932);
and U9926 (N_9926,N_6697,N_7151);
or U9927 (N_9927,N_5544,N_6447);
nand U9928 (N_9928,N_6471,N_6420);
or U9929 (N_9929,N_5522,N_5976);
nand U9930 (N_9930,N_6150,N_6405);
nor U9931 (N_9931,N_6424,N_6522);
nor U9932 (N_9932,N_7334,N_7015);
nor U9933 (N_9933,N_5679,N_5835);
or U9934 (N_9934,N_7057,N_6936);
or U9935 (N_9935,N_5559,N_6600);
nand U9936 (N_9936,N_6420,N_7372);
and U9937 (N_9937,N_7248,N_5911);
and U9938 (N_9938,N_5173,N_6303);
nand U9939 (N_9939,N_6956,N_5656);
or U9940 (N_9940,N_6124,N_7165);
or U9941 (N_9941,N_5012,N_7419);
or U9942 (N_9942,N_6076,N_5877);
nand U9943 (N_9943,N_7267,N_5696);
or U9944 (N_9944,N_6546,N_7050);
nand U9945 (N_9945,N_5019,N_6059);
nand U9946 (N_9946,N_5882,N_5873);
or U9947 (N_9947,N_7416,N_5474);
xor U9948 (N_9948,N_5783,N_5219);
nor U9949 (N_9949,N_7042,N_7262);
and U9950 (N_9950,N_5227,N_5766);
or U9951 (N_9951,N_6829,N_5983);
and U9952 (N_9952,N_5041,N_5147);
and U9953 (N_9953,N_7350,N_7059);
and U9954 (N_9954,N_5420,N_5777);
nand U9955 (N_9955,N_5493,N_6414);
nand U9956 (N_9956,N_5029,N_6568);
and U9957 (N_9957,N_7267,N_6773);
nand U9958 (N_9958,N_5942,N_7213);
nor U9959 (N_9959,N_5961,N_5200);
or U9960 (N_9960,N_6095,N_6559);
and U9961 (N_9961,N_7003,N_6376);
nor U9962 (N_9962,N_5924,N_6982);
nand U9963 (N_9963,N_6194,N_6256);
xnor U9964 (N_9964,N_7208,N_5013);
nor U9965 (N_9965,N_6557,N_7183);
nand U9966 (N_9966,N_5868,N_7437);
nand U9967 (N_9967,N_6525,N_7326);
nor U9968 (N_9968,N_5778,N_7026);
or U9969 (N_9969,N_5435,N_7468);
nor U9970 (N_9970,N_5707,N_6928);
nor U9971 (N_9971,N_6411,N_6840);
and U9972 (N_9972,N_6189,N_5801);
and U9973 (N_9973,N_5157,N_7028);
or U9974 (N_9974,N_7108,N_6257);
and U9975 (N_9975,N_6233,N_5432);
nand U9976 (N_9976,N_6258,N_6464);
and U9977 (N_9977,N_5306,N_5104);
nor U9978 (N_9978,N_5669,N_7361);
and U9979 (N_9979,N_6172,N_6622);
nand U9980 (N_9980,N_5304,N_6141);
nor U9981 (N_9981,N_7118,N_5061);
and U9982 (N_9982,N_6457,N_6838);
and U9983 (N_9983,N_5626,N_6348);
and U9984 (N_9984,N_7127,N_7161);
nand U9985 (N_9985,N_6268,N_5951);
nor U9986 (N_9986,N_5482,N_6787);
nand U9987 (N_9987,N_6217,N_5522);
nand U9988 (N_9988,N_7438,N_6503);
and U9989 (N_9989,N_7137,N_6097);
and U9990 (N_9990,N_5014,N_6763);
or U9991 (N_9991,N_5157,N_5415);
or U9992 (N_9992,N_6281,N_5035);
and U9993 (N_9993,N_6714,N_6928);
and U9994 (N_9994,N_5697,N_6862);
and U9995 (N_9995,N_7421,N_5946);
nand U9996 (N_9996,N_5077,N_6044);
and U9997 (N_9997,N_6918,N_7243);
nand U9998 (N_9998,N_6313,N_6379);
nor U9999 (N_9999,N_7318,N_6782);
and UO_0 (O_0,N_9571,N_7938);
or UO_1 (O_1,N_9581,N_8519);
nor UO_2 (O_2,N_7912,N_9659);
nand UO_3 (O_3,N_9208,N_9544);
or UO_4 (O_4,N_7902,N_9677);
nand UO_5 (O_5,N_8313,N_8425);
and UO_6 (O_6,N_9287,N_8947);
or UO_7 (O_7,N_8049,N_8727);
or UO_8 (O_8,N_8260,N_8142);
nor UO_9 (O_9,N_8786,N_8466);
and UO_10 (O_10,N_9793,N_8985);
nand UO_11 (O_11,N_9718,N_9462);
and UO_12 (O_12,N_7726,N_9080);
nor UO_13 (O_13,N_9833,N_8428);
and UO_14 (O_14,N_9383,N_8081);
nor UO_15 (O_15,N_8792,N_8318);
nand UO_16 (O_16,N_8654,N_7553);
nor UO_17 (O_17,N_7819,N_9706);
nand UO_18 (O_18,N_9487,N_8168);
nand UO_19 (O_19,N_7592,N_9745);
or UO_20 (O_20,N_8910,N_9855);
or UO_21 (O_21,N_8427,N_9825);
or UO_22 (O_22,N_8934,N_8093);
or UO_23 (O_23,N_8671,N_9503);
xor UO_24 (O_24,N_8320,N_7882);
nand UO_25 (O_25,N_8605,N_9961);
nor UO_26 (O_26,N_8137,N_8590);
or UO_27 (O_27,N_9130,N_8381);
nor UO_28 (O_28,N_8303,N_8082);
nor UO_29 (O_29,N_9001,N_9430);
and UO_30 (O_30,N_8909,N_9176);
or UO_31 (O_31,N_9940,N_7834);
nor UO_32 (O_32,N_8310,N_8461);
nand UO_33 (O_33,N_7674,N_8784);
or UO_34 (O_34,N_9134,N_9442);
or UO_35 (O_35,N_9580,N_9167);
nand UO_36 (O_36,N_9350,N_8973);
and UO_37 (O_37,N_9140,N_8588);
nor UO_38 (O_38,N_9570,N_9780);
nand UO_39 (O_39,N_8709,N_8202);
nand UO_40 (O_40,N_8366,N_8402);
nand UO_41 (O_41,N_8764,N_8562);
nor UO_42 (O_42,N_8743,N_7616);
or UO_43 (O_43,N_8702,N_8656);
nand UO_44 (O_44,N_9372,N_8420);
nor UO_45 (O_45,N_7949,N_7919);
or UO_46 (O_46,N_7530,N_9055);
nand UO_47 (O_47,N_7851,N_8338);
or UO_48 (O_48,N_8056,N_7754);
and UO_49 (O_49,N_7898,N_9108);
nor UO_50 (O_50,N_8210,N_9872);
and UO_51 (O_51,N_9906,N_8876);
nand UO_52 (O_52,N_7599,N_7782);
nor UO_53 (O_53,N_8437,N_8959);
and UO_54 (O_54,N_8760,N_9364);
and UO_55 (O_55,N_9199,N_9559);
nand UO_56 (O_56,N_7994,N_9636);
xnor UO_57 (O_57,N_8679,N_7733);
nor UO_58 (O_58,N_7612,N_7789);
or UO_59 (O_59,N_9841,N_8109);
and UO_60 (O_60,N_8031,N_8383);
or UO_61 (O_61,N_9010,N_9076);
nand UO_62 (O_62,N_8359,N_8261);
or UO_63 (O_63,N_9719,N_8548);
nor UO_64 (O_64,N_7904,N_9107);
nor UO_65 (O_65,N_9754,N_7868);
and UO_66 (O_66,N_9952,N_8148);
and UO_67 (O_67,N_8875,N_7929);
or UO_68 (O_68,N_9276,N_9895);
xnor UO_69 (O_69,N_8323,N_9510);
nand UO_70 (O_70,N_9813,N_8620);
nand UO_71 (O_71,N_8287,N_8066);
nor UO_72 (O_72,N_8482,N_8350);
nand UO_73 (O_73,N_8933,N_7812);
xnor UO_74 (O_74,N_9908,N_8996);
or UO_75 (O_75,N_8074,N_8255);
nor UO_76 (O_76,N_7531,N_9060);
or UO_77 (O_77,N_9909,N_8854);
nand UO_78 (O_78,N_7846,N_8232);
nor UO_79 (O_79,N_7661,N_9365);
and UO_80 (O_80,N_9241,N_8440);
and UO_81 (O_81,N_9903,N_8882);
nor UO_82 (O_82,N_7710,N_8751);
nor UO_83 (O_83,N_8516,N_8607);
nand UO_84 (O_84,N_9550,N_9099);
nor UO_85 (O_85,N_8669,N_8829);
or UO_86 (O_86,N_9876,N_8517);
or UO_87 (O_87,N_9911,N_9264);
nand UO_88 (O_88,N_8668,N_8922);
nor UO_89 (O_89,N_8853,N_8489);
and UO_90 (O_90,N_7738,N_8906);
or UO_91 (O_91,N_9464,N_7961);
nor UO_92 (O_92,N_9824,N_9786);
nor UO_93 (O_93,N_8227,N_7793);
and UO_94 (O_94,N_9970,N_9905);
nand UO_95 (O_95,N_9574,N_9697);
nor UO_96 (O_96,N_8724,N_9516);
nor UO_97 (O_97,N_9238,N_8980);
and UO_98 (O_98,N_7686,N_9349);
and UO_99 (O_99,N_8094,N_9561);
nand UO_100 (O_100,N_9837,N_8932);
nand UO_101 (O_101,N_8042,N_8463);
or UO_102 (O_102,N_8895,N_9842);
nand UO_103 (O_103,N_9293,N_8887);
or UO_104 (O_104,N_9897,N_9727);
or UO_105 (O_105,N_7838,N_9930);
or UO_106 (O_106,N_7984,N_7758);
nor UO_107 (O_107,N_7887,N_8872);
or UO_108 (O_108,N_7817,N_7593);
nand UO_109 (O_109,N_8067,N_7958);
nand UO_110 (O_110,N_8083,N_7610);
nor UO_111 (O_111,N_9759,N_7897);
nor UO_112 (O_112,N_9377,N_9007);
nor UO_113 (O_113,N_8475,N_8803);
nor UO_114 (O_114,N_7600,N_9644);
nand UO_115 (O_115,N_9476,N_9686);
nor UO_116 (O_116,N_8448,N_9030);
or UO_117 (O_117,N_8237,N_8016);
or UO_118 (O_118,N_9450,N_8936);
nand UO_119 (O_119,N_8289,N_9846);
or UO_120 (O_120,N_9454,N_8115);
nor UO_121 (O_121,N_7922,N_9640);
and UO_122 (O_122,N_8911,N_7878);
nand UO_123 (O_123,N_9734,N_7700);
and UO_124 (O_124,N_9986,N_9654);
xnor UO_125 (O_125,N_8271,N_9221);
or UO_126 (O_126,N_8358,N_8116);
and UO_127 (O_127,N_9589,N_9353);
nand UO_128 (O_128,N_9035,N_9771);
nand UO_129 (O_129,N_8086,N_9845);
or UO_130 (O_130,N_8849,N_9071);
nand UO_131 (O_131,N_9843,N_9434);
nor UO_132 (O_132,N_9411,N_7893);
xnor UO_133 (O_133,N_8581,N_8672);
or UO_134 (O_134,N_7840,N_9712);
and UO_135 (O_135,N_9963,N_8737);
xor UO_136 (O_136,N_8987,N_9165);
nor UO_137 (O_137,N_9693,N_9358);
and UO_138 (O_138,N_8617,N_8152);
and UO_139 (O_139,N_7697,N_7970);
or UO_140 (O_140,N_7895,N_9506);
or UO_141 (O_141,N_9344,N_9133);
nor UO_142 (O_142,N_7565,N_8307);
or UO_143 (O_143,N_9115,N_9122);
and UO_144 (O_144,N_9301,N_8953);
nand UO_145 (O_145,N_8663,N_9072);
or UO_146 (O_146,N_9057,N_9881);
nor UO_147 (O_147,N_7881,N_8376);
and UO_148 (O_148,N_9203,N_9960);
and UO_149 (O_149,N_9614,N_9146);
or UO_150 (O_150,N_9950,N_9689);
nor UO_151 (O_151,N_9191,N_9973);
nor UO_152 (O_152,N_7656,N_9106);
nand UO_153 (O_153,N_9048,N_8367);
nand UO_154 (O_154,N_8883,N_9894);
nand UO_155 (O_155,N_8711,N_7648);
nand UO_156 (O_156,N_8057,N_7857);
nor UO_157 (O_157,N_8648,N_8174);
and UO_158 (O_158,N_8575,N_8843);
nor UO_159 (O_159,N_8185,N_7535);
and UO_160 (O_160,N_7785,N_7936);
nor UO_161 (O_161,N_9817,N_8962);
or UO_162 (O_162,N_8154,N_8403);
nor UO_163 (O_163,N_8881,N_7832);
and UO_164 (O_164,N_9660,N_7559);
or UO_165 (O_165,N_8008,N_9242);
nand UO_166 (O_166,N_7644,N_9101);
and UO_167 (O_167,N_9765,N_8337);
nor UO_168 (O_168,N_9747,N_7571);
nor UO_169 (O_169,N_9066,N_9231);
nor UO_170 (O_170,N_9956,N_9585);
nand UO_171 (O_171,N_8378,N_9838);
nor UO_172 (O_172,N_8612,N_9619);
nor UO_173 (O_173,N_9814,N_9000);
or UO_174 (O_174,N_9187,N_8631);
xor UO_175 (O_175,N_7753,N_8326);
nor UO_176 (O_176,N_9091,N_8828);
or UO_177 (O_177,N_7876,N_8469);
nor UO_178 (O_178,N_8963,N_9114);
nor UO_179 (O_179,N_9310,N_8537);
and UO_180 (O_180,N_9529,N_9914);
and UO_181 (O_181,N_9576,N_9233);
and UO_182 (O_182,N_7512,N_8951);
nor UO_183 (O_183,N_7652,N_8385);
nand UO_184 (O_184,N_8815,N_7569);
and UO_185 (O_185,N_7960,N_8741);
nand UO_186 (O_186,N_9965,N_8190);
nand UO_187 (O_187,N_8496,N_9514);
or UO_188 (O_188,N_9641,N_8034);
nand UO_189 (O_189,N_7605,N_7532);
and UO_190 (O_190,N_9426,N_8479);
nor UO_191 (O_191,N_9998,N_9920);
or UO_192 (O_192,N_9482,N_9999);
nor UO_193 (O_193,N_7997,N_9286);
xor UO_194 (O_194,N_9338,N_8890);
nor UO_195 (O_195,N_8369,N_8543);
or UO_196 (O_196,N_9112,N_8293);
nand UO_197 (O_197,N_9145,N_9306);
and UO_198 (O_198,N_8561,N_9275);
or UO_199 (O_199,N_9764,N_7811);
or UO_200 (O_200,N_9971,N_9156);
xor UO_201 (O_201,N_7801,N_9179);
nand UO_202 (O_202,N_8652,N_9877);
and UO_203 (O_203,N_7705,N_9210);
and UO_204 (O_204,N_9994,N_8915);
and UO_205 (O_205,N_9505,N_9456);
nor UO_206 (O_206,N_9588,N_8673);
and UO_207 (O_207,N_7803,N_8602);
or UO_208 (O_208,N_7988,N_8226);
or UO_209 (O_209,N_8546,N_8111);
and UO_210 (O_210,N_9595,N_8344);
nor UO_211 (O_211,N_9412,N_9110);
nor UO_212 (O_212,N_8823,N_8865);
and UO_213 (O_213,N_7708,N_9535);
or UO_214 (O_214,N_8306,N_9945);
and UO_215 (O_215,N_8619,N_8270);
and UO_216 (O_216,N_9702,N_9768);
nand UO_217 (O_217,N_8001,N_9398);
or UO_218 (O_218,N_7871,N_7792);
nor UO_219 (O_219,N_9530,N_8248);
and UO_220 (O_220,N_9135,N_8222);
nand UO_221 (O_221,N_8451,N_9951);
and UO_222 (O_222,N_9681,N_8242);
and UO_223 (O_223,N_9847,N_8462);
nand UO_224 (O_224,N_9189,N_7673);
and UO_225 (O_225,N_8166,N_8062);
nor UO_226 (O_226,N_9009,N_8935);
nand UO_227 (O_227,N_9586,N_9651);
and UO_228 (O_228,N_7815,N_9031);
xnor UO_229 (O_229,N_9161,N_9262);
and UO_230 (O_230,N_9878,N_8609);
nand UO_231 (O_231,N_8308,N_9710);
nor UO_232 (O_232,N_9065,N_8643);
or UO_233 (O_233,N_8208,N_8052);
nand UO_234 (O_234,N_9796,N_9992);
nor UO_235 (O_235,N_9974,N_9739);
and UO_236 (O_236,N_8972,N_8811);
and UO_237 (O_237,N_9169,N_9003);
or UO_238 (O_238,N_9495,N_8090);
or UO_239 (O_239,N_8627,N_7609);
nor UO_240 (O_240,N_8777,N_8015);
nand UO_241 (O_241,N_9451,N_8742);
nor UO_242 (O_242,N_7845,N_8921);
or UO_243 (O_243,N_9781,N_9446);
nand UO_244 (O_244,N_8691,N_8674);
or UO_245 (O_245,N_7722,N_9818);
or UO_246 (O_246,N_8520,N_7784);
or UO_247 (O_247,N_7990,N_9705);
nor UO_248 (O_248,N_9407,N_9033);
nand UO_249 (O_249,N_7719,N_9160);
nand UO_250 (O_250,N_9700,N_9483);
nand UO_251 (O_251,N_8259,N_9272);
nand UO_252 (O_252,N_9429,N_8867);
and UO_253 (O_253,N_9853,N_9501);
nor UO_254 (O_254,N_7730,N_8613);
or UO_255 (O_255,N_8597,N_8201);
and UO_256 (O_256,N_8304,N_7947);
or UO_257 (O_257,N_7767,N_8079);
nor UO_258 (O_258,N_9722,N_9389);
and UO_259 (O_259,N_8916,N_9691);
nor UO_260 (O_260,N_8263,N_8256);
nor UO_261 (O_261,N_8397,N_8719);
nor UO_262 (O_262,N_9069,N_9590);
nand UO_263 (O_263,N_9937,N_7611);
and UO_264 (O_264,N_9246,N_8230);
nor UO_265 (O_265,N_9798,N_9333);
nor UO_266 (O_266,N_8856,N_8219);
or UO_267 (O_267,N_7714,N_8738);
nor UO_268 (O_268,N_9744,N_9117);
or UO_269 (O_269,N_8641,N_7880);
or UO_270 (O_270,N_8974,N_9014);
and UO_271 (O_271,N_7826,N_9621);
nand UO_272 (O_272,N_7540,N_9041);
or UO_273 (O_273,N_8472,N_7854);
or UO_274 (O_274,N_8228,N_9043);
and UO_275 (O_275,N_9315,N_8013);
nor UO_276 (O_276,N_8703,N_9247);
xnor UO_277 (O_277,N_7776,N_8923);
nor UO_278 (O_278,N_8851,N_9159);
nor UO_279 (O_279,N_7809,N_9475);
and UO_280 (O_280,N_7794,N_9849);
nor UO_281 (O_281,N_7561,N_9525);
nor UO_282 (O_282,N_9664,N_8113);
or UO_283 (O_283,N_8370,N_9005);
and UO_284 (O_284,N_7901,N_9982);
nand UO_285 (O_285,N_8276,N_8594);
nand UO_286 (O_286,N_8362,N_7933);
nor UO_287 (O_287,N_7944,N_8273);
and UO_288 (O_288,N_8110,N_9207);
or UO_289 (O_289,N_8838,N_7796);
or UO_290 (O_290,N_9511,N_7770);
and UO_291 (O_291,N_9356,N_8407);
nand UO_292 (O_292,N_9447,N_8464);
nor UO_293 (O_293,N_8950,N_9673);
nand UO_294 (O_294,N_9969,N_9892);
and UO_295 (O_295,N_7798,N_9193);
nand UO_296 (O_296,N_8690,N_8536);
nand UO_297 (O_297,N_8436,N_9980);
nor UO_298 (O_298,N_9694,N_8863);
and UO_299 (O_299,N_9282,N_9594);
and UO_300 (O_300,N_8162,N_7536);
or UO_301 (O_301,N_7576,N_8840);
nor UO_302 (O_302,N_9256,N_8000);
nand UO_303 (O_303,N_9981,N_9488);
nand UO_304 (O_304,N_8192,N_8329);
nor UO_305 (O_305,N_8623,N_9886);
and UO_306 (O_306,N_9624,N_8697);
or UO_307 (O_307,N_9564,N_8107);
nor UO_308 (O_308,N_9936,N_8503);
nand UO_309 (O_309,N_9360,N_9224);
xor UO_310 (O_310,N_8297,N_7704);
nor UO_311 (O_311,N_9183,N_8589);
nor UO_312 (O_312,N_8637,N_9313);
or UO_313 (O_313,N_9240,N_9320);
nor UO_314 (O_314,N_9804,N_9541);
or UO_315 (O_315,N_8091,N_8744);
nand UO_316 (O_316,N_9216,N_9491);
or UO_317 (O_317,N_9717,N_9889);
or UO_318 (O_318,N_8340,N_8802);
or UO_319 (O_319,N_9124,N_9870);
or UO_320 (O_320,N_8651,N_8797);
nor UO_321 (O_321,N_8640,N_8745);
and UO_322 (O_322,N_9284,N_9753);
nand UO_323 (O_323,N_8141,N_7830);
nor UO_324 (O_324,N_8127,N_8993);
nand UO_325 (O_325,N_8756,N_8145);
or UO_326 (O_326,N_9551,N_7667);
or UO_327 (O_327,N_8006,N_7608);
or UO_328 (O_328,N_7790,N_9004);
or UO_329 (O_329,N_9730,N_8434);
nand UO_330 (O_330,N_9283,N_8591);
and UO_331 (O_331,N_9863,N_9649);
and UO_332 (O_332,N_9883,N_9896);
or UO_333 (O_333,N_8371,N_7856);
nor UO_334 (O_334,N_9778,N_9204);
and UO_335 (O_335,N_9835,N_8610);
or UO_336 (O_336,N_8655,N_7509);
nand UO_337 (O_337,N_9391,N_8822);
nor UO_338 (O_338,N_8132,N_8398);
and UO_339 (O_339,N_9288,N_8284);
nand UO_340 (O_340,N_9336,N_8179);
nand UO_341 (O_341,N_8707,N_9016);
or UO_342 (O_342,N_8522,N_8636);
xor UO_343 (O_343,N_8501,N_7603);
or UO_344 (O_344,N_8164,N_8723);
nand UO_345 (O_345,N_7588,N_8047);
and UO_346 (O_346,N_8010,N_8146);
and UO_347 (O_347,N_8483,N_8021);
nand UO_348 (O_348,N_7558,N_9404);
and UO_349 (O_349,N_8125,N_9954);
and UO_350 (O_350,N_8975,N_7703);
nand UO_351 (O_351,N_8924,N_7516);
nor UO_352 (O_352,N_8382,N_8040);
nand UO_353 (O_353,N_8258,N_8732);
nor UO_354 (O_354,N_8862,N_9471);
and UO_355 (O_355,N_7642,N_7715);
nand UO_356 (O_356,N_8790,N_7615);
and UO_357 (O_357,N_8136,N_9683);
or UO_358 (O_358,N_7843,N_8106);
nor UO_359 (O_359,N_8955,N_9195);
and UO_360 (O_360,N_8846,N_8624);
and UO_361 (O_361,N_9844,N_8130);
nand UO_362 (O_362,N_9642,N_8353);
or UO_363 (O_363,N_8905,N_8269);
or UO_364 (O_364,N_8002,N_9815);
and UO_365 (O_365,N_9173,N_8423);
nand UO_366 (O_366,N_8585,N_7914);
nor UO_367 (O_367,N_9128,N_8526);
and UO_368 (O_368,N_7825,N_9334);
and UO_369 (O_369,N_9512,N_7954);
nand UO_370 (O_370,N_7556,N_8170);
or UO_371 (O_371,N_8728,N_7731);
nor UO_372 (O_372,N_9109,N_9271);
nand UO_373 (O_373,N_9968,N_9746);
or UO_374 (O_374,N_8505,N_9695);
nor UO_375 (O_375,N_9791,N_9228);
nand UO_376 (O_376,N_9898,N_7890);
nor UO_377 (O_377,N_7542,N_9939);
nand UO_378 (O_378,N_7723,N_9834);
nand UO_379 (O_379,N_8073,N_8465);
and UO_380 (O_380,N_7850,N_9490);
or UO_381 (O_381,N_7818,N_9987);
and UO_382 (O_382,N_9439,N_8611);
or UO_383 (O_383,N_8979,N_8285);
nor UO_384 (O_384,N_8704,N_8254);
or UO_385 (O_385,N_8864,N_8291);
and UO_386 (O_386,N_9543,N_8433);
and UO_387 (O_387,N_8386,N_8100);
or UO_388 (O_388,N_9045,N_8981);
nand UO_389 (O_389,N_9259,N_7788);
nor UO_390 (O_390,N_8312,N_7810);
nand UO_391 (O_391,N_8649,N_7965);
nor UO_392 (O_392,N_9655,N_7757);
and UO_393 (O_393,N_9023,N_9147);
or UO_394 (O_394,N_7595,N_8220);
nand UO_395 (O_395,N_9629,N_9604);
nand UO_396 (O_396,N_8681,N_9502);
nor UO_397 (O_397,N_9254,N_9704);
or UO_398 (O_398,N_9387,N_9139);
nand UO_399 (O_399,N_8061,N_7590);
nand UO_400 (O_400,N_9552,N_9931);
nor UO_401 (O_401,N_8044,N_7650);
nor UO_402 (O_402,N_7573,N_9489);
and UO_403 (O_403,N_7732,N_9767);
and UO_404 (O_404,N_9304,N_9050);
nand UO_405 (O_405,N_9486,N_9011);
or UO_406 (O_406,N_9612,N_9402);
nor UO_407 (O_407,N_7602,N_8188);
nor UO_408 (O_408,N_9465,N_8429);
nor UO_409 (O_409,N_8529,N_7614);
nand UO_410 (O_410,N_9184,N_9562);
or UO_411 (O_411,N_8249,N_9738);
or UO_412 (O_412,N_9361,N_7980);
and UO_413 (O_413,N_9626,N_8638);
or UO_414 (O_414,N_9947,N_9202);
nand UO_415 (O_415,N_8294,N_9557);
nand UO_416 (O_416,N_7597,N_8267);
nand UO_417 (O_417,N_9504,N_8839);
nand UO_418 (O_418,N_9458,N_7563);
nor UO_419 (O_419,N_7501,N_8492);
xnor UO_420 (O_420,N_8579,N_9639);
and UO_421 (O_421,N_9251,N_7539);
nand UO_422 (O_422,N_8776,N_9943);
or UO_423 (O_423,N_8346,N_8327);
nand UO_424 (O_424,N_8494,N_9285);
xor UO_425 (O_425,N_8076,N_9281);
and UO_426 (O_426,N_9335,N_9369);
or UO_427 (O_427,N_9913,N_7950);
nor UO_428 (O_428,N_9696,N_8969);
nor UO_429 (O_429,N_9800,N_7908);
nand UO_430 (O_430,N_8169,N_8808);
nand UO_431 (O_431,N_8506,N_9959);
nand UO_432 (O_432,N_8907,N_9723);
xnor UO_433 (O_433,N_9556,N_9790);
nor UO_434 (O_434,N_8244,N_8504);
and UO_435 (O_435,N_9729,N_9498);
nand UO_436 (O_436,N_9280,N_9953);
or UO_437 (O_437,N_8582,N_9784);
nor UO_438 (O_438,N_7505,N_9017);
and UO_439 (O_439,N_8595,N_9972);
nand UO_440 (O_440,N_7665,N_8938);
nor UO_441 (O_441,N_8357,N_8518);
and UO_442 (O_442,N_8858,N_8439);
and UO_443 (O_443,N_7601,N_9805);
nand UO_444 (O_444,N_9674,N_8873);
or UO_445 (O_445,N_9234,N_8454);
nand UO_446 (O_446,N_7967,N_9680);
nor UO_447 (O_447,N_8578,N_9020);
and UO_448 (O_448,N_9608,N_8372);
or UO_449 (O_449,N_7645,N_9865);
and UO_450 (O_450,N_9311,N_9307);
or UO_451 (O_451,N_8432,N_8171);
nand UO_452 (O_452,N_8471,N_7623);
and UO_453 (O_453,N_7655,N_7735);
nor UO_454 (O_454,N_8629,N_9265);
and UO_455 (O_455,N_7751,N_8901);
and UO_456 (O_456,N_8685,N_7783);
nand UO_457 (O_457,N_9047,N_8525);
and UO_458 (O_458,N_7606,N_8512);
and UO_459 (O_459,N_8213,N_7734);
and UO_460 (O_460,N_8749,N_8759);
or UO_461 (O_461,N_8527,N_9270);
or UO_462 (O_462,N_9770,N_8859);
and UO_463 (O_463,N_7907,N_9915);
and UO_464 (O_464,N_9685,N_8161);
nor UO_465 (O_465,N_9116,N_8941);
or UO_466 (O_466,N_8946,N_7632);
nor UO_467 (O_467,N_8758,N_9996);
nor UO_468 (O_468,N_8622,N_8055);
or UO_469 (O_469,N_8976,N_8241);
nor UO_470 (O_470,N_8957,N_7515);
nand UO_471 (O_471,N_7749,N_8621);
and UO_472 (O_472,N_9527,N_8818);
nand UO_473 (O_473,N_7800,N_7909);
or UO_474 (O_474,N_9657,N_9609);
and UO_475 (O_475,N_8361,N_9616);
or UO_476 (O_476,N_8186,N_7762);
and UO_477 (O_477,N_8559,N_7635);
nor UO_478 (O_478,N_7678,N_9941);
nand UO_479 (O_479,N_9597,N_8399);
and UO_480 (O_480,N_9049,N_8236);
nand UO_481 (O_481,N_8319,N_7831);
nor UO_482 (O_482,N_8592,N_9775);
nor UO_483 (O_483,N_9257,N_9403);
or UO_484 (O_484,N_9445,N_9875);
nor UO_485 (O_485,N_9728,N_8120);
and UO_486 (O_486,N_9096,N_9816);
nor UO_487 (O_487,N_8983,N_7677);
nor UO_488 (O_488,N_9643,N_7799);
nor UO_489 (O_489,N_9255,N_7568);
nor UO_490 (O_490,N_8274,N_9324);
nand UO_491 (O_491,N_9467,N_8835);
and UO_492 (O_492,N_8874,N_7872);
nand UO_493 (O_493,N_9823,N_9266);
and UO_494 (O_494,N_9230,N_8752);
nor UO_495 (O_495,N_9039,N_9013);
nand UO_496 (O_496,N_8701,N_9185);
nand UO_497 (O_497,N_7666,N_8007);
nand UO_498 (O_498,N_7720,N_9910);
nand UO_499 (O_499,N_8481,N_9463);
nor UO_500 (O_500,N_8059,N_9181);
or UO_501 (O_501,N_7824,N_9749);
and UO_502 (O_502,N_9171,N_8675);
or UO_503 (O_503,N_8354,N_7663);
nor UO_504 (O_504,N_9603,N_8027);
nor UO_505 (O_505,N_9563,N_8003);
or UO_506 (O_506,N_8278,N_7574);
or UO_507 (O_507,N_8836,N_8603);
and UO_508 (O_508,N_9785,N_9158);
nand UO_509 (O_509,N_8288,N_9901);
nand UO_510 (O_510,N_8217,N_8689);
and UO_511 (O_511,N_9792,N_8343);
nand UO_512 (O_512,N_9537,N_9237);
nor UO_513 (O_513,N_8814,N_9417);
and UO_514 (O_514,N_8415,N_8309);
or UO_515 (O_515,N_8450,N_8314);
nand UO_516 (O_516,N_8688,N_8404);
nor UO_517 (O_517,N_8060,N_8301);
or UO_518 (O_518,N_7688,N_9967);
or UO_519 (O_519,N_8355,N_8245);
xnor UO_520 (O_520,N_7528,N_8114);
and UO_521 (O_521,N_8426,N_9410);
nor UO_522 (O_522,N_8410,N_8138);
and UO_523 (O_523,N_9789,N_8457);
nor UO_524 (O_524,N_9774,N_9725);
nor UO_525 (O_525,N_8214,N_8195);
or UO_526 (O_526,N_8224,N_7739);
or UO_527 (O_527,N_9188,N_8364);
nand UO_528 (O_528,N_9277,N_8153);
or UO_529 (O_529,N_9085,N_8966);
and UO_530 (O_530,N_7816,N_7756);
or UO_531 (O_531,N_7518,N_8720);
or UO_532 (O_532,N_9370,N_9367);
and UO_533 (O_533,N_9025,N_8424);
or UO_534 (O_534,N_9569,N_8687);
nor UO_535 (O_535,N_8601,N_8869);
and UO_536 (O_536,N_9121,N_7684);
xor UO_537 (O_537,N_7930,N_9297);
and UO_538 (O_538,N_9888,N_8533);
or UO_539 (O_539,N_9545,N_7504);
nand UO_540 (O_540,N_7619,N_9715);
nand UO_541 (O_541,N_8124,N_8032);
nor UO_542 (O_542,N_8332,N_7903);
nand UO_543 (O_543,N_9752,N_9218);
and UO_544 (O_544,N_9979,N_8468);
nor UO_545 (O_545,N_9422,N_8948);
nor UO_546 (O_546,N_8341,N_9912);
nor UO_547 (O_547,N_9305,N_9480);
nand UO_548 (O_548,N_8077,N_9008);
nand UO_549 (O_549,N_7637,N_8769);
nor UO_550 (O_550,N_9743,N_9864);
nor UO_551 (O_551,N_9648,N_9997);
nand UO_552 (O_552,N_9322,N_7764);
or UO_553 (O_553,N_9572,N_7560);
nor UO_554 (O_554,N_9587,N_9568);
nor UO_555 (O_555,N_9382,N_9086);
nor UO_556 (O_556,N_8122,N_8712);
and UO_557 (O_557,N_8305,N_8104);
nand UO_558 (O_558,N_8216,N_9617);
and UO_559 (O_559,N_9596,N_7523);
and UO_560 (O_560,N_9783,N_9806);
and UO_561 (O_561,N_7668,N_8630);
or UO_562 (O_562,N_9175,N_9037);
or UO_563 (O_563,N_8204,N_9907);
nand UO_564 (O_564,N_7693,N_9194);
nor UO_565 (O_565,N_7971,N_8809);
nand UO_566 (O_566,N_7724,N_8286);
nand UO_567 (O_567,N_8264,N_9602);
and UO_568 (O_568,N_9352,N_8406);
and UO_569 (O_569,N_9736,N_8568);
or UO_570 (O_570,N_9152,N_9850);
nand UO_571 (O_571,N_7546,N_9524);
or UO_572 (O_572,N_8197,N_9082);
or UO_573 (O_573,N_7769,N_9902);
nand UO_574 (O_574,N_8279,N_9312);
or UO_575 (O_575,N_9212,N_9002);
and UO_576 (O_576,N_7946,N_8335);
nand UO_577 (O_577,N_7526,N_7543);
and UO_578 (O_578,N_9484,N_7579);
and UO_579 (O_579,N_8998,N_8566);
nor UO_580 (O_580,N_8896,N_9460);
nor UO_581 (O_581,N_9220,N_8747);
and UO_582 (O_582,N_9565,N_9857);
and UO_583 (O_583,N_7695,N_7959);
nand UO_584 (O_584,N_8816,N_8495);
nand UO_585 (O_585,N_9326,N_9645);
nand UO_586 (O_586,N_9073,N_7502);
nand UO_587 (O_587,N_8140,N_9500);
nand UO_588 (O_588,N_8499,N_8826);
nand UO_589 (O_589,N_9390,N_8647);
nand UO_590 (O_590,N_8817,N_8714);
nand UO_591 (O_591,N_8348,N_8356);
or UO_592 (O_592,N_8658,N_7837);
nand UO_593 (O_593,N_8984,N_9687);
and UO_594 (O_594,N_9308,N_8878);
nand UO_595 (O_595,N_9123,N_7510);
or UO_596 (O_596,N_9539,N_9938);
nor UO_597 (O_597,N_9141,N_8158);
and UO_598 (O_598,N_9425,N_7805);
or UO_599 (O_599,N_9087,N_9405);
nor UO_600 (O_600,N_9090,N_8788);
nor UO_601 (O_601,N_9531,N_8734);
nand UO_602 (O_602,N_8417,N_9517);
nor UO_603 (O_603,N_7952,N_8928);
xor UO_604 (O_604,N_7774,N_8128);
or UO_605 (O_605,N_8772,N_7987);
and UO_606 (O_606,N_8473,N_8740);
or UO_607 (O_607,N_7916,N_7634);
nand UO_608 (O_608,N_7982,N_9143);
nor UO_609 (O_609,N_9578,N_9225);
and UO_610 (O_610,N_9720,N_7989);
and UO_611 (O_611,N_8708,N_8035);
nand UO_612 (O_612,N_9862,N_9290);
and UO_613 (O_613,N_8650,N_9309);
or UO_614 (O_614,N_9478,N_8544);
or UO_615 (O_615,N_7617,N_8408);
or UO_616 (O_616,N_8748,N_8196);
nor UO_617 (O_617,N_9600,N_9890);
and UO_618 (O_618,N_9547,N_8474);
and UO_619 (O_619,N_9461,N_8670);
nand UO_620 (O_620,N_8857,N_7575);
and UO_621 (O_621,N_9245,N_9493);
nor UO_622 (O_622,N_7658,N_8990);
and UO_623 (O_623,N_8509,N_8292);
and UO_624 (O_624,N_9679,N_8135);
or UO_625 (O_625,N_8553,N_9497);
nand UO_626 (O_626,N_8695,N_9170);
nand UO_627 (O_627,N_9515,N_9385);
and UO_628 (O_628,N_9274,N_9396);
nand UO_629 (O_629,N_8283,N_8710);
or UO_630 (O_630,N_8488,N_7578);
nor UO_631 (O_631,N_8870,N_7676);
or UO_632 (O_632,N_8995,N_8085);
or UO_633 (O_633,N_8486,N_7647);
nor UO_634 (O_634,N_8025,N_9591);
nand UO_635 (O_635,N_9481,N_7891);
nor UO_636 (O_636,N_8225,N_8485);
nor UO_637 (O_637,N_8847,N_9345);
nor UO_638 (O_638,N_8129,N_8063);
or UO_639 (O_639,N_7955,N_8456);
nand UO_640 (O_640,N_9150,N_8721);
nand UO_641 (O_641,N_8296,N_7591);
or UO_642 (O_642,N_9026,N_9605);
nor UO_643 (O_643,N_7827,N_7896);
or UO_644 (O_644,N_8713,N_9455);
nand UO_645 (O_645,N_8510,N_9296);
nor UO_646 (O_646,N_7956,N_8952);
or UO_647 (O_647,N_7636,N_9757);
nor UO_648 (O_648,N_9468,N_8586);
and UO_649 (O_649,N_8763,N_9018);
nor UO_650 (O_650,N_9182,N_9132);
and UO_651 (O_651,N_8534,N_8556);
nand UO_652 (O_652,N_8441,N_8877);
and UO_653 (O_653,N_9138,N_9869);
or UO_654 (O_654,N_8334,N_7630);
nand UO_655 (O_655,N_7519,N_7580);
and UO_656 (O_656,N_8038,N_9991);
and UO_657 (O_657,N_9708,N_8089);
or UO_658 (O_658,N_9214,N_9661);
or UO_659 (O_659,N_8540,N_8753);
nand UO_660 (O_660,N_8683,N_9083);
nor UO_661 (O_661,N_8960,N_8005);
nand UO_662 (O_662,N_7981,N_9519);
nand UO_663 (O_663,N_7849,N_8994);
and UO_664 (O_664,N_8087,N_9222);
nand UO_665 (O_665,N_9542,N_9144);
and UO_666 (O_666,N_9802,N_7624);
and UO_667 (O_667,N_8807,N_8902);
and UO_668 (O_668,N_9810,N_8435);
or UO_669 (O_669,N_7942,N_8253);
or UO_670 (O_670,N_7775,N_9359);
and UO_671 (O_671,N_8223,N_8438);
and UO_672 (O_672,N_9413,N_9113);
and UO_673 (O_673,N_7701,N_8065);
nor UO_674 (O_674,N_7983,N_9226);
nand UO_675 (O_675,N_9215,N_8266);
nand UO_676 (O_676,N_9703,N_9229);
nand UO_677 (O_677,N_9735,N_7620);
nand UO_678 (O_678,N_9638,N_7917);
nand UO_679 (O_679,N_9059,N_8231);
or UO_680 (O_680,N_9388,N_9093);
and UO_681 (O_681,N_8762,N_9630);
and UO_682 (O_682,N_8604,N_9533);
nand UO_683 (O_683,N_8507,N_8899);
nand UO_684 (O_684,N_9637,N_9851);
nor UO_685 (O_685,N_8555,N_7741);
nor UO_686 (O_686,N_9357,N_8247);
and UO_687 (O_687,N_7685,N_8467);
nand UO_688 (O_688,N_7687,N_8088);
nor UO_689 (O_689,N_9104,N_8502);
or UO_690 (O_690,N_8238,N_8978);
nor UO_691 (O_691,N_8351,N_7589);
nor UO_692 (O_692,N_8058,N_9958);
nand UO_693 (O_693,N_8912,N_7842);
and UO_694 (O_694,N_9466,N_8653);
or UO_695 (O_695,N_9692,N_8277);
or UO_696 (O_696,N_9758,N_9263);
or UO_697 (O_697,N_8487,N_8131);
and UO_698 (O_698,N_8191,N_8167);
or UO_699 (O_699,N_8024,N_9707);
nand UO_700 (O_700,N_8780,N_9440);
and UO_701 (O_701,N_7836,N_8860);
nor UO_702 (O_702,N_9151,N_8694);
or UO_703 (O_703,N_9618,N_8182);
nand UO_704 (O_704,N_8178,N_9957);
nor UO_705 (O_705,N_8806,N_9522);
nand UO_706 (O_706,N_8419,N_7807);
nor UO_707 (O_707,N_9432,N_8295);
or UO_708 (O_708,N_7533,N_8773);
and UO_709 (O_709,N_9111,N_7839);
or UO_710 (O_710,N_9916,N_9190);
or UO_711 (O_711,N_9435,N_7996);
nand UO_712 (O_712,N_8218,N_8360);
and UO_713 (O_713,N_9698,N_8477);
nand UO_714 (O_714,N_9149,N_9354);
nor UO_715 (O_715,N_7986,N_8642);
and UO_716 (O_716,N_9078,N_9347);
nand UO_717 (O_717,N_7583,N_8147);
or UO_718 (O_718,N_8345,N_9021);
nand UO_719 (O_719,N_9097,N_9428);
and UO_720 (O_720,N_9470,N_8325);
or UO_721 (O_721,N_7594,N_7545);
nand UO_722 (O_722,N_8036,N_7985);
nand UO_723 (O_723,N_9300,N_8498);
nand UO_724 (O_724,N_8392,N_9538);
nor UO_725 (O_725,N_8019,N_7978);
nand UO_726 (O_726,N_9092,N_7649);
and UO_727 (O_727,N_8850,N_8616);
nor UO_728 (O_728,N_9858,N_7527);
and UO_729 (O_729,N_9829,N_9613);
nand UO_730 (O_730,N_8989,N_7672);
nand UO_731 (O_731,N_8149,N_7835);
and UO_732 (O_732,N_7889,N_9408);
nor UO_733 (O_733,N_9507,N_8317);
and UO_734 (O_734,N_8470,N_9343);
and UO_735 (O_735,N_9560,N_8886);
nand UO_736 (O_736,N_9006,N_8401);
or UO_737 (O_737,N_8508,N_8930);
and UO_738 (O_738,N_9201,N_9666);
nand UO_739 (O_739,N_8235,N_9485);
and UO_740 (O_740,N_8892,N_7729);
or UO_741 (O_741,N_9332,N_9874);
nand UO_742 (O_742,N_7866,N_8885);
and UO_743 (O_743,N_9536,N_9248);
nand UO_744 (O_744,N_8693,N_7823);
nor UO_745 (O_745,N_8660,N_8330);
nor UO_746 (O_746,N_9615,N_7828);
nand UO_747 (O_747,N_8324,N_8009);
or UO_748 (O_748,N_8400,N_9075);
or UO_749 (O_749,N_9762,N_9601);
or UO_750 (O_750,N_8888,N_9070);
and UO_751 (O_751,N_7927,N_9948);
nand UO_752 (O_752,N_9607,N_7659);
or UO_753 (O_753,N_9633,N_8961);
nand UO_754 (O_754,N_8699,N_9386);
nand UO_755 (O_755,N_8280,N_8409);
or UO_756 (O_756,N_8163,N_7847);
or UO_757 (O_757,N_9826,N_8731);
and UO_758 (O_758,N_8725,N_8956);
nand UO_759 (O_759,N_8583,N_8414);
and UO_760 (O_760,N_8598,N_8387);
nand UO_761 (O_761,N_7848,N_8810);
nor UO_762 (O_762,N_9646,N_9839);
or UO_763 (O_763,N_8453,N_9955);
and UO_764 (O_764,N_8041,N_9269);
nor UO_765 (O_765,N_9394,N_8080);
or UO_766 (O_766,N_8390,N_8262);
and UO_767 (O_767,N_9374,N_7943);
nand UO_768 (O_768,N_9095,N_9341);
and UO_769 (O_769,N_9213,N_8889);
or UO_770 (O_770,N_9866,N_7888);
nand UO_771 (O_771,N_7541,N_9022);
and UO_772 (O_772,N_7681,N_8377);
nand UO_773 (O_773,N_9922,N_9244);
or UO_774 (O_774,N_8193,N_8944);
nor UO_775 (O_775,N_8841,N_8026);
and UO_776 (O_776,N_8405,N_9261);
nor UO_777 (O_777,N_7627,N_9196);
or UO_778 (O_778,N_9378,N_9062);
and UO_779 (O_779,N_9098,N_9379);
and UO_780 (O_780,N_8391,N_9418);
and UO_781 (O_781,N_9119,N_7750);
and UO_782 (O_782,N_7683,N_8099);
and UO_783 (O_783,N_9038,N_8717);
or UO_784 (O_784,N_7945,N_8240);
or UO_785 (O_785,N_8374,N_9976);
nand UO_786 (O_786,N_8584,N_9227);
nand UO_787 (O_787,N_8144,N_8715);
or UO_788 (O_788,N_8422,N_7679);
or UO_789 (O_789,N_9925,N_7717);
or UO_790 (O_790,N_8634,N_8119);
nor UO_791 (O_791,N_8117,N_7671);
and UO_792 (O_792,N_9917,N_7884);
nand UO_793 (O_793,N_7507,N_9131);
nand UO_794 (O_794,N_9061,N_7711);
nor UO_795 (O_795,N_8608,N_8336);
nand UO_796 (O_796,N_9019,N_9079);
and UO_797 (O_797,N_8368,N_8339);
nor UO_798 (O_798,N_8991,N_9828);
and UO_799 (O_799,N_8967,N_9840);
and UO_800 (O_800,N_8446,N_8160);
or UO_801 (O_801,N_8528,N_7915);
and UO_802 (O_802,N_8903,N_8785);
nand UO_803 (O_803,N_7694,N_9136);
and UO_804 (O_804,N_8234,N_9628);
nor UO_805 (O_805,N_9040,N_8833);
nor UO_806 (O_806,N_7538,N_7968);
and UO_807 (O_807,N_8789,N_9209);
nand UO_808 (O_808,N_8667,N_9724);
nor UO_809 (O_809,N_7804,N_8842);
nand UO_810 (O_810,N_7795,N_8416);
nor UO_811 (O_811,N_8573,N_8644);
nand UO_812 (O_812,N_8600,N_9223);
or UO_813 (O_813,N_9794,N_8239);
nand UO_814 (O_814,N_8898,N_9325);
nand UO_815 (O_815,N_9620,N_9174);
and UO_816 (O_816,N_8039,N_7791);
or UO_817 (O_817,N_9831,N_8275);
or UO_818 (O_818,N_8150,N_9154);
or UO_819 (O_819,N_9582,N_8557);
and UO_820 (O_820,N_9027,N_8207);
or UO_821 (O_821,N_8761,N_9807);
and UO_822 (O_822,N_9526,N_9808);
or UO_823 (O_823,N_7906,N_7707);
and UO_824 (O_824,N_9355,N_7669);
and UO_825 (O_825,N_8175,N_7822);
or UO_826 (O_826,N_9164,N_8821);
and UO_827 (O_827,N_8824,N_8831);
nand UO_828 (O_828,N_8484,N_7964);
nand UO_829 (O_829,N_7973,N_9200);
and UO_830 (O_830,N_8813,N_8615);
nor UO_831 (O_831,N_9583,N_8480);
or UO_832 (O_832,N_9232,N_8331);
nor UO_833 (O_833,N_7638,N_8799);
nand UO_834 (O_834,N_9811,N_9219);
and UO_835 (O_835,N_9670,N_8676);
nor UO_836 (O_836,N_9625,N_9457);
nand UO_837 (O_837,N_7821,N_9584);
nand UO_838 (O_838,N_7555,N_8105);
and UO_839 (O_839,N_9635,N_8316);
or UO_840 (O_840,N_9477,N_8965);
nand UO_841 (O_841,N_8754,N_8200);
and UO_842 (O_842,N_8913,N_8606);
nand UO_843 (O_843,N_8793,N_9820);
or UO_844 (O_844,N_9094,N_8535);
or UO_845 (O_845,N_8118,N_8730);
and UO_846 (O_846,N_7550,N_9822);
nand UO_847 (O_847,N_9662,N_8029);
nand UO_848 (O_848,N_9258,N_9289);
or UO_849 (O_849,N_8596,N_9197);
and UO_850 (O_850,N_9942,N_7780);
nor UO_851 (O_851,N_7761,N_9267);
nor UO_852 (O_852,N_8302,N_9761);
and UO_853 (O_853,N_8682,N_8491);
nand UO_854 (O_854,N_9964,N_9701);
nand UO_855 (O_855,N_7993,N_9647);
or UO_856 (O_856,N_9988,N_8139);
and UO_857 (O_857,N_7709,N_8490);
and UO_858 (O_858,N_8252,N_9756);
and UO_859 (O_859,N_7859,N_9294);
nor UO_860 (O_860,N_9074,N_9342);
and UO_861 (O_861,N_7948,N_9924);
nor UO_862 (O_862,N_8686,N_7974);
or UO_863 (O_863,N_7745,N_9406);
nor UO_864 (O_864,N_8143,N_8078);
or UO_865 (O_865,N_8265,N_8739);
and UO_866 (O_866,N_9423,N_9153);
and UO_867 (O_867,N_7660,N_8268);
nand UO_868 (O_868,N_9279,N_9830);
nand UO_869 (O_869,N_9779,N_9373);
nand UO_870 (O_870,N_8781,N_7923);
and UO_871 (O_871,N_9946,N_9496);
nand UO_872 (O_872,N_7855,N_8908);
and UO_873 (O_873,N_7585,N_8871);
and UO_874 (O_874,N_9126,N_9180);
and UO_875 (O_875,N_9933,N_7874);
xnor UO_876 (O_876,N_9236,N_9298);
nor UO_877 (O_877,N_7625,N_9848);
or UO_878 (O_878,N_8290,N_9599);
and UO_879 (O_879,N_8560,N_8476);
nand UO_880 (O_880,N_9675,N_8447);
or UO_881 (O_881,N_8997,N_9051);
or UO_882 (O_882,N_7924,N_7514);
nand UO_883 (O_883,N_9977,N_7779);
or UO_884 (O_884,N_8970,N_7873);
nor UO_885 (O_885,N_8037,N_8282);
nor UO_886 (O_886,N_7657,N_7905);
nor UO_887 (O_887,N_9868,N_8045);
nand UO_888 (O_888,N_9887,N_9371);
nand UO_889 (O_889,N_8971,N_8389);
nand UO_890 (O_890,N_9318,N_9366);
nand UO_891 (O_891,N_7875,N_9801);
and UO_892 (O_892,N_8092,N_7736);
and UO_893 (O_893,N_8199,N_9521);
nor UO_894 (O_894,N_8733,N_9314);
nor UO_895 (O_895,N_8134,N_9157);
nand UO_896 (O_896,N_8639,N_7867);
nor UO_897 (O_897,N_8891,N_7529);
nor UO_898 (O_898,N_9376,N_7587);
and UO_899 (O_899,N_7651,N_8521);
and UO_900 (O_900,N_8299,N_9443);
nand UO_901 (O_901,N_9927,N_7921);
and UO_902 (O_902,N_9827,N_7742);
nor UO_903 (O_903,N_8513,N_9782);
or UO_904 (O_904,N_7633,N_8861);
nor UO_905 (O_905,N_9323,N_8778);
nor UO_906 (O_906,N_9363,N_8523);
or UO_907 (O_907,N_8943,N_9867);
or UO_908 (O_908,N_9711,N_8445);
nor UO_909 (O_909,N_8070,N_8497);
or UO_910 (O_910,N_9102,N_8982);
nand UO_911 (O_911,N_7534,N_8698);
or UO_912 (O_912,N_7883,N_9741);
or UO_913 (O_913,N_8661,N_8333);
nand UO_914 (O_914,N_9769,N_9766);
nor UO_915 (O_915,N_9611,N_8795);
nand UO_916 (O_916,N_7939,N_9012);
nand UO_917 (O_917,N_9579,N_9015);
or UO_918 (O_918,N_7765,N_9509);
nor UO_919 (O_919,N_9330,N_8157);
nand UO_920 (O_920,N_9384,N_8766);
nor UO_921 (O_921,N_7771,N_9206);
or UO_922 (O_922,N_9966,N_7766);
or UO_923 (O_923,N_7662,N_8645);
or UO_924 (O_924,N_7877,N_7596);
or UO_925 (O_925,N_9172,N_8571);
nor UO_926 (O_926,N_8394,N_9508);
nor UO_927 (O_927,N_8363,N_8380);
and UO_928 (O_928,N_8541,N_7737);
nand UO_929 (O_929,N_9885,N_9499);
nand UO_930 (O_930,N_9575,N_8159);
nor UO_931 (O_931,N_9469,N_9260);
or UO_932 (O_932,N_8493,N_8926);
nand UO_933 (O_933,N_7513,N_7743);
and UO_934 (O_934,N_9652,N_7992);
nand UO_935 (O_935,N_7979,N_7931);
and UO_936 (O_936,N_8812,N_8352);
nand UO_937 (O_937,N_7721,N_7682);
or UO_938 (O_938,N_8012,N_7511);
nor UO_939 (O_939,N_8431,N_9978);
and UO_940 (O_940,N_7748,N_9733);
nor UO_941 (O_941,N_8126,N_8251);
nor UO_942 (O_942,N_7969,N_9125);
nand UO_943 (O_943,N_7957,N_9235);
nor UO_944 (O_944,N_7862,N_7863);
xnor UO_945 (O_945,N_9773,N_8937);
nor UO_946 (O_946,N_9668,N_7937);
and UO_947 (O_947,N_9742,N_8662);
and UO_948 (O_948,N_8384,N_8375);
nand UO_949 (O_949,N_7698,N_9437);
and UO_950 (O_950,N_8570,N_8388);
nand UO_951 (O_951,N_9631,N_7598);
and UO_952 (O_952,N_8108,N_7829);
or UO_953 (O_953,N_9919,N_7692);
nor UO_954 (O_954,N_9120,N_8189);
or UO_955 (O_955,N_9032,N_8900);
nor UO_956 (O_956,N_8444,N_9162);
or UO_957 (O_957,N_9249,N_8298);
nor UO_958 (O_958,N_7935,N_9492);
nor UO_959 (O_959,N_9737,N_8180);
and UO_960 (O_960,N_8311,N_9751);
or UO_961 (O_961,N_7562,N_9893);
or UO_962 (O_962,N_9854,N_9441);
and UO_963 (O_963,N_8187,N_7577);
nor UO_964 (O_964,N_9750,N_8834);
nand UO_965 (O_965,N_7547,N_7564);
and UO_966 (O_966,N_7772,N_7503);
or UO_967 (O_967,N_9714,N_8177);
and UO_968 (O_968,N_8830,N_8054);
and UO_969 (O_969,N_9415,N_9105);
or UO_970 (O_970,N_8565,N_9540);
nand UO_971 (O_971,N_9409,N_9063);
nand UO_972 (O_972,N_7557,N_9346);
or UO_973 (O_973,N_7934,N_7706);
nor UO_974 (O_974,N_8075,N_9036);
nand UO_975 (O_975,N_8750,N_9678);
nor UO_976 (O_976,N_9879,N_8819);
nand UO_977 (O_977,N_7781,N_9268);
nor UO_978 (O_978,N_9178,N_9532);
and UO_979 (O_979,N_9054,N_7654);
or UO_980 (O_980,N_9339,N_9278);
nand UO_981 (O_981,N_8272,N_8837);
nor UO_982 (O_982,N_7628,N_7725);
nor UO_983 (O_983,N_9419,N_7689);
nor UO_984 (O_984,N_7699,N_8300);
and UO_985 (O_985,N_8677,N_9990);
nand UO_986 (O_986,N_9676,N_9089);
nand UO_987 (O_987,N_9029,N_7680);
or UO_988 (O_988,N_8205,N_9474);
nand UO_989 (O_989,N_9534,N_7524);
and UO_990 (O_990,N_9053,N_8452);
nand UO_991 (O_991,N_8614,N_9684);
nand UO_992 (O_992,N_8102,N_9064);
nor UO_993 (O_993,N_9669,N_9395);
or UO_994 (O_994,N_9348,N_8033);
nor UO_995 (O_995,N_8539,N_9880);
and UO_996 (O_996,N_8735,N_7759);
and UO_997 (O_997,N_9573,N_8051);
nor UO_998 (O_998,N_7932,N_8992);
or UO_999 (O_999,N_9518,N_9553);
nand UO_1000 (O_1000,N_7778,N_7852);
or UO_1001 (O_1001,N_7584,N_8718);
nor UO_1002 (O_1002,N_9929,N_8365);
nor UO_1003 (O_1003,N_7976,N_7629);
and UO_1004 (O_1004,N_8246,N_8023);
or UO_1005 (O_1005,N_7641,N_7910);
and UO_1006 (O_1006,N_8787,N_8798);
or UO_1007 (O_1007,N_8347,N_9421);
nor UO_1008 (O_1008,N_7626,N_9928);
or UO_1009 (O_1009,N_8215,N_9494);
nor UO_1010 (O_1010,N_9024,N_7718);
nand UO_1011 (O_1011,N_9129,N_7913);
and UO_1012 (O_1012,N_9243,N_9882);
nor UO_1013 (O_1013,N_8209,N_9393);
nand UO_1014 (O_1014,N_9431,N_9856);
and UO_1015 (O_1015,N_8716,N_8925);
and UO_1016 (O_1016,N_7844,N_9672);
and UO_1017 (O_1017,N_8097,N_7773);
nor UO_1018 (O_1018,N_8046,N_8659);
nor UO_1019 (O_1019,N_7940,N_8852);
and UO_1020 (O_1020,N_9622,N_8626);
and UO_1021 (O_1021,N_9392,N_7777);
nor UO_1022 (O_1022,N_9088,N_7506);
nand UO_1023 (O_1023,N_8212,N_7586);
nand UO_1024 (O_1024,N_8914,N_8593);
nor UO_1025 (O_1025,N_8206,N_8919);
and UO_1026 (O_1026,N_8563,N_8050);
and UO_1027 (O_1027,N_9250,N_8940);
and UO_1028 (O_1028,N_8599,N_8478);
and UO_1029 (O_1029,N_9566,N_8511);
and UO_1030 (O_1030,N_9397,N_8665);
nor UO_1031 (O_1031,N_9716,N_8574);
nand UO_1032 (O_1032,N_9148,N_9084);
and UO_1033 (O_1033,N_7814,N_8373);
and UO_1034 (O_1034,N_9832,N_9932);
or UO_1035 (O_1035,N_7728,N_9787);
nand UO_1036 (O_1036,N_8770,N_9812);
nor UO_1037 (O_1037,N_8999,N_8552);
nand UO_1038 (O_1038,N_9137,N_9993);
and UO_1039 (O_1039,N_7899,N_7918);
and UO_1040 (O_1040,N_8729,N_8538);
nor UO_1041 (O_1041,N_9799,N_8576);
nand UO_1042 (O_1042,N_9058,N_8030);
nand UO_1043 (O_1043,N_8664,N_7670);
nor UO_1044 (O_1044,N_9650,N_8460);
nor UO_1045 (O_1045,N_9427,N_8514);
nor UO_1046 (O_1046,N_8567,N_8443);
xnor UO_1047 (O_1047,N_8072,N_8411);
and UO_1048 (O_1048,N_7858,N_9192);
or UO_1049 (O_1049,N_8929,N_8918);
nand UO_1050 (O_1050,N_8155,N_7640);
nand UO_1051 (O_1051,N_9081,N_9690);
nand UO_1052 (O_1052,N_8071,N_9688);
and UO_1053 (O_1053,N_9861,N_8328);
nor UO_1054 (O_1054,N_9667,N_8736);
nand UO_1055 (O_1055,N_7975,N_8515);
nand UO_1056 (O_1056,N_8791,N_7554);
or UO_1057 (O_1057,N_9459,N_8779);
and UO_1058 (O_1058,N_9975,N_9523);
and UO_1059 (O_1059,N_9949,N_7607);
nand UO_1060 (O_1060,N_7552,N_7953);
nand UO_1061 (O_1061,N_9610,N_9567);
or UO_1062 (O_1062,N_8988,N_7746);
nor UO_1063 (O_1063,N_9142,N_8804);
xor UO_1064 (O_1064,N_8172,N_7716);
nor UO_1065 (O_1065,N_9118,N_9211);
nand UO_1066 (O_1066,N_7522,N_9362);
nor UO_1067 (O_1067,N_9163,N_9453);
nor UO_1068 (O_1068,N_7653,N_9473);
or UO_1069 (O_1069,N_9328,N_8281);
nor UO_1070 (O_1070,N_8825,N_8349);
or UO_1071 (O_1071,N_9327,N_7727);
nand UO_1072 (O_1072,N_9292,N_7500);
and UO_1073 (O_1073,N_9375,N_9186);
nor UO_1074 (O_1074,N_8500,N_8635);
or UO_1075 (O_1075,N_9984,N_8430);
and UO_1076 (O_1076,N_7820,N_9295);
and UO_1077 (O_1077,N_9623,N_9340);
nor UO_1078 (O_1078,N_9709,N_9420);
and UO_1079 (O_1079,N_8322,N_8181);
nand UO_1080 (O_1080,N_7853,N_9891);
or UO_1081 (O_1081,N_9755,N_9052);
and UO_1082 (O_1082,N_8767,N_8945);
and UO_1083 (O_1083,N_7548,N_9884);
and UO_1084 (O_1084,N_7570,N_8580);
nand UO_1085 (O_1085,N_8395,N_8101);
or UO_1086 (O_1086,N_8977,N_8068);
or UO_1087 (O_1087,N_7768,N_8832);
or UO_1088 (O_1088,N_8156,N_8550);
nand UO_1089 (O_1089,N_9198,N_8547);
nor UO_1090 (O_1090,N_9546,N_9989);
or UO_1091 (O_1091,N_9424,N_9433);
nor UO_1092 (O_1092,N_9329,N_9918);
nand UO_1093 (O_1093,N_8879,N_9944);
nand UO_1094 (O_1094,N_9665,N_9177);
and UO_1095 (O_1095,N_9803,N_8939);
xnor UO_1096 (O_1096,N_7928,N_8257);
and UO_1097 (O_1097,N_8564,N_9836);
and UO_1098 (O_1098,N_9337,N_8705);
or UO_1099 (O_1099,N_9479,N_8893);
or UO_1100 (O_1100,N_7998,N_7664);
and UO_1101 (O_1101,N_7951,N_9797);
nand UO_1102 (O_1102,N_8551,N_8805);
or UO_1103 (O_1103,N_9548,N_9217);
or UO_1104 (O_1104,N_8771,N_8628);
nor UO_1105 (O_1105,N_9520,N_8198);
nor UO_1106 (O_1106,N_7551,N_9316);
nand UO_1107 (O_1107,N_9449,N_7567);
and UO_1108 (O_1108,N_8421,N_9593);
nand UO_1109 (O_1109,N_8011,N_7841);
and UO_1110 (O_1110,N_8184,N_7537);
nand UO_1111 (O_1111,N_9042,N_8229);
or UO_1112 (O_1112,N_8183,N_8722);
and UO_1113 (O_1113,N_7864,N_8103);
and UO_1114 (O_1114,N_9028,N_9381);
nor UO_1115 (O_1115,N_7926,N_8211);
nor UO_1116 (O_1116,N_8123,N_9627);
or UO_1117 (O_1117,N_8726,N_9732);
nor UO_1118 (O_1118,N_8755,N_9962);
or UO_1119 (O_1119,N_8646,N_8459);
or UO_1120 (O_1120,N_9899,N_7604);
nand UO_1121 (O_1121,N_9663,N_8868);
and UO_1122 (O_1122,N_9317,N_7763);
and UO_1123 (O_1123,N_9472,N_9873);
nand UO_1124 (O_1124,N_9166,N_8554);
nand UO_1125 (O_1125,N_7712,N_8680);
or UO_1126 (O_1126,N_9795,N_9438);
nand UO_1127 (O_1127,N_8043,N_7869);
or UO_1128 (O_1128,N_7966,N_9321);
or UO_1129 (O_1129,N_7691,N_8455);
and UO_1130 (O_1130,N_9303,N_8549);
nor UO_1131 (O_1131,N_9252,N_8625);
and UO_1132 (O_1132,N_8545,N_9554);
and UO_1133 (O_1133,N_8986,N_8558);
nor UO_1134 (O_1134,N_9558,N_9444);
and UO_1135 (O_1135,N_7886,N_8569);
and UO_1136 (O_1136,N_8004,N_7696);
or UO_1137 (O_1137,N_9934,N_7860);
or UO_1138 (O_1138,N_9721,N_8796);
nor UO_1139 (O_1139,N_7702,N_9592);
nand UO_1140 (O_1140,N_8315,N_7755);
or UO_1141 (O_1141,N_7622,N_9598);
nand UO_1142 (O_1142,N_8618,N_7963);
or UO_1143 (O_1143,N_8678,N_8931);
nor UO_1144 (O_1144,N_7675,N_8018);
nand UO_1145 (O_1145,N_9904,N_8855);
nor UO_1146 (O_1146,N_8657,N_7991);
and UO_1147 (O_1147,N_8165,N_9068);
or UO_1148 (O_1148,N_9900,N_7760);
nor UO_1149 (O_1149,N_9351,N_7618);
and UO_1150 (O_1150,N_9302,N_7544);
nand UO_1151 (O_1151,N_8194,N_7892);
or UO_1152 (O_1152,N_7813,N_8112);
and UO_1153 (O_1153,N_8866,N_9448);
xor UO_1154 (O_1154,N_9995,N_8768);
nor UO_1155 (O_1155,N_9860,N_7525);
nor UO_1156 (O_1156,N_9331,N_8632);
nor UO_1157 (O_1157,N_8844,N_8053);
nand UO_1158 (O_1158,N_8765,N_8098);
nor UO_1159 (O_1159,N_9168,N_7566);
and UO_1160 (O_1160,N_7582,N_8173);
or UO_1161 (O_1161,N_9871,N_8442);
nor UO_1162 (O_1162,N_7870,N_9606);
nor UO_1163 (O_1163,N_9046,N_9416);
nand UO_1164 (O_1164,N_8017,N_8949);
nor UO_1165 (O_1165,N_9653,N_7879);
nand UO_1166 (O_1166,N_9852,N_8572);
and UO_1167 (O_1167,N_8530,N_8532);
nand UO_1168 (O_1168,N_9777,N_7920);
nor UO_1169 (O_1169,N_9760,N_9549);
nor UO_1170 (O_1170,N_7802,N_8884);
or UO_1171 (O_1171,N_7646,N_7613);
nor UO_1172 (O_1172,N_8542,N_7713);
and UO_1173 (O_1173,N_8783,N_9513);
and UO_1174 (O_1174,N_8958,N_8794);
nor UO_1175 (O_1175,N_8746,N_8014);
nand UO_1176 (O_1176,N_8022,N_8233);
or UO_1177 (O_1177,N_9414,N_8121);
or UO_1178 (O_1178,N_7941,N_8801);
and UO_1179 (O_1179,N_8782,N_8964);
or UO_1180 (O_1180,N_8706,N_9985);
and UO_1181 (O_1181,N_9935,N_9713);
and UO_1182 (O_1182,N_8942,N_7962);
or UO_1183 (O_1183,N_9399,N_7900);
and UO_1184 (O_1184,N_9699,N_8920);
nand UO_1185 (O_1185,N_8413,N_9034);
or UO_1186 (O_1186,N_7747,N_9632);
and UO_1187 (O_1187,N_8666,N_7885);
nand UO_1188 (O_1188,N_7865,N_9401);
and UO_1189 (O_1189,N_9253,N_9983);
nand UO_1190 (O_1190,N_9819,N_8342);
and UO_1191 (O_1191,N_8418,N_9127);
nor UO_1192 (O_1192,N_9056,N_7690);
nor UO_1193 (O_1193,N_8633,N_7621);
nand UO_1194 (O_1194,N_9926,N_7861);
xor UO_1195 (O_1195,N_7508,N_8396);
nand UO_1196 (O_1196,N_8250,N_8692);
or UO_1197 (O_1197,N_7911,N_9656);
nor UO_1198 (O_1198,N_8133,N_8524);
and UO_1199 (O_1199,N_9859,N_9155);
and UO_1200 (O_1200,N_9368,N_9921);
nand UO_1201 (O_1201,N_7643,N_8048);
nor UO_1202 (O_1202,N_9380,N_7631);
or UO_1203 (O_1203,N_9436,N_9239);
nor UO_1204 (O_1204,N_8904,N_9291);
and UO_1205 (O_1205,N_9748,N_9731);
and UO_1206 (O_1206,N_7549,N_8845);
or UO_1207 (O_1207,N_8020,N_8880);
nor UO_1208 (O_1208,N_8827,N_9067);
or UO_1209 (O_1209,N_8696,N_8449);
nand UO_1210 (O_1210,N_8243,N_7740);
and UO_1211 (O_1211,N_8084,N_9682);
and UO_1212 (O_1212,N_9671,N_8321);
and UO_1213 (O_1213,N_7581,N_9788);
and UO_1214 (O_1214,N_9205,N_9273);
nor UO_1215 (O_1215,N_9776,N_8096);
or UO_1216 (O_1216,N_9658,N_7572);
nor UO_1217 (O_1217,N_8684,N_9740);
nand UO_1218 (O_1218,N_9763,N_9103);
and UO_1219 (O_1219,N_9809,N_9923);
nand UO_1220 (O_1220,N_8379,N_7972);
nand UO_1221 (O_1221,N_8095,N_9044);
nor UO_1222 (O_1222,N_7977,N_8775);
nand UO_1223 (O_1223,N_7521,N_8968);
nand UO_1224 (O_1224,N_7517,N_8203);
nand UO_1225 (O_1225,N_7995,N_7787);
nor UO_1226 (O_1226,N_8820,N_8151);
nand UO_1227 (O_1227,N_9577,N_8587);
nand UO_1228 (O_1228,N_8412,N_7925);
or UO_1229 (O_1229,N_8954,N_7639);
nor UO_1230 (O_1230,N_9528,N_8774);
nor UO_1231 (O_1231,N_7833,N_8176);
or UO_1232 (O_1232,N_8757,N_8700);
or UO_1233 (O_1233,N_8221,N_7808);
and UO_1234 (O_1234,N_7752,N_8577);
or UO_1235 (O_1235,N_9452,N_9772);
nand UO_1236 (O_1236,N_9400,N_8393);
nor UO_1237 (O_1237,N_8897,N_8917);
nand UO_1238 (O_1238,N_8800,N_8069);
nand UO_1239 (O_1239,N_8064,N_7744);
or UO_1240 (O_1240,N_7999,N_9821);
nand UO_1241 (O_1241,N_9319,N_7806);
nor UO_1242 (O_1242,N_8531,N_8894);
or UO_1243 (O_1243,N_9077,N_7894);
nand UO_1244 (O_1244,N_7797,N_9100);
nand UO_1245 (O_1245,N_8848,N_7786);
nand UO_1246 (O_1246,N_9726,N_8028);
or UO_1247 (O_1247,N_7520,N_8927);
nand UO_1248 (O_1248,N_8458,N_9555);
nor UO_1249 (O_1249,N_9299,N_9634);
nand UO_1250 (O_1250,N_8616,N_8511);
nand UO_1251 (O_1251,N_8516,N_7520);
and UO_1252 (O_1252,N_8769,N_7931);
nor UO_1253 (O_1253,N_9373,N_8292);
and UO_1254 (O_1254,N_7501,N_9351);
and UO_1255 (O_1255,N_9169,N_9173);
or UO_1256 (O_1256,N_8732,N_7827);
or UO_1257 (O_1257,N_9235,N_7743);
and UO_1258 (O_1258,N_9944,N_9379);
nor UO_1259 (O_1259,N_8095,N_8308);
nand UO_1260 (O_1260,N_8594,N_7587);
and UO_1261 (O_1261,N_7610,N_7669);
nor UO_1262 (O_1262,N_8422,N_8902);
nor UO_1263 (O_1263,N_9865,N_7657);
nor UO_1264 (O_1264,N_8085,N_9981);
nor UO_1265 (O_1265,N_8318,N_9015);
nor UO_1266 (O_1266,N_7523,N_8410);
and UO_1267 (O_1267,N_9646,N_9658);
nand UO_1268 (O_1268,N_9566,N_8485);
and UO_1269 (O_1269,N_8174,N_9640);
or UO_1270 (O_1270,N_8188,N_9600);
nand UO_1271 (O_1271,N_9529,N_9959);
nand UO_1272 (O_1272,N_9699,N_8973);
nand UO_1273 (O_1273,N_8522,N_9987);
and UO_1274 (O_1274,N_8115,N_8015);
and UO_1275 (O_1275,N_9226,N_9633);
nor UO_1276 (O_1276,N_7774,N_8476);
and UO_1277 (O_1277,N_8643,N_9340);
nand UO_1278 (O_1278,N_8077,N_9831);
nor UO_1279 (O_1279,N_8214,N_9915);
and UO_1280 (O_1280,N_7896,N_8546);
and UO_1281 (O_1281,N_9714,N_8443);
or UO_1282 (O_1282,N_7618,N_8639);
and UO_1283 (O_1283,N_8977,N_8745);
nand UO_1284 (O_1284,N_8556,N_9887);
and UO_1285 (O_1285,N_9514,N_9072);
nand UO_1286 (O_1286,N_9117,N_8319);
nand UO_1287 (O_1287,N_8705,N_9103);
nand UO_1288 (O_1288,N_8243,N_8716);
or UO_1289 (O_1289,N_9494,N_9240);
nand UO_1290 (O_1290,N_7681,N_7662);
or UO_1291 (O_1291,N_7818,N_9190);
or UO_1292 (O_1292,N_8544,N_7618);
nor UO_1293 (O_1293,N_8630,N_9335);
and UO_1294 (O_1294,N_9266,N_7629);
and UO_1295 (O_1295,N_7662,N_7763);
and UO_1296 (O_1296,N_9125,N_8962);
nor UO_1297 (O_1297,N_9605,N_9879);
and UO_1298 (O_1298,N_8892,N_7790);
nor UO_1299 (O_1299,N_9423,N_9226);
or UO_1300 (O_1300,N_9758,N_9095);
and UO_1301 (O_1301,N_8847,N_8864);
nor UO_1302 (O_1302,N_8896,N_8091);
and UO_1303 (O_1303,N_8166,N_9994);
nand UO_1304 (O_1304,N_8320,N_9987);
nand UO_1305 (O_1305,N_8541,N_8906);
or UO_1306 (O_1306,N_9932,N_8878);
nor UO_1307 (O_1307,N_9946,N_8189);
nand UO_1308 (O_1308,N_9317,N_8410);
and UO_1309 (O_1309,N_8423,N_7807);
or UO_1310 (O_1310,N_8255,N_8527);
nand UO_1311 (O_1311,N_9437,N_7524);
or UO_1312 (O_1312,N_9172,N_8092);
nor UO_1313 (O_1313,N_7749,N_8203);
nor UO_1314 (O_1314,N_7862,N_9139);
nand UO_1315 (O_1315,N_8234,N_8807);
xnor UO_1316 (O_1316,N_7782,N_9014);
and UO_1317 (O_1317,N_9751,N_8212);
and UO_1318 (O_1318,N_9030,N_7950);
or UO_1319 (O_1319,N_9562,N_7727);
or UO_1320 (O_1320,N_9595,N_8446);
and UO_1321 (O_1321,N_8715,N_7517);
and UO_1322 (O_1322,N_7579,N_8561);
or UO_1323 (O_1323,N_9344,N_8349);
nor UO_1324 (O_1324,N_8037,N_7623);
nand UO_1325 (O_1325,N_7751,N_9302);
and UO_1326 (O_1326,N_8533,N_9357);
nand UO_1327 (O_1327,N_7934,N_8700);
nand UO_1328 (O_1328,N_9902,N_8987);
and UO_1329 (O_1329,N_8565,N_9371);
nand UO_1330 (O_1330,N_8235,N_8471);
nand UO_1331 (O_1331,N_9602,N_7810);
and UO_1332 (O_1332,N_9362,N_9230);
and UO_1333 (O_1333,N_7796,N_8749);
nor UO_1334 (O_1334,N_8566,N_9741);
nand UO_1335 (O_1335,N_7674,N_7607);
nand UO_1336 (O_1336,N_9085,N_8213);
nand UO_1337 (O_1337,N_8306,N_8480);
and UO_1338 (O_1338,N_7692,N_8172);
nand UO_1339 (O_1339,N_9295,N_7590);
and UO_1340 (O_1340,N_9810,N_7765);
nor UO_1341 (O_1341,N_7840,N_7606);
or UO_1342 (O_1342,N_8955,N_7895);
nor UO_1343 (O_1343,N_9248,N_9477);
and UO_1344 (O_1344,N_9186,N_8332);
or UO_1345 (O_1345,N_8010,N_9083);
nand UO_1346 (O_1346,N_7581,N_9449);
and UO_1347 (O_1347,N_9797,N_9706);
and UO_1348 (O_1348,N_9808,N_7960);
nor UO_1349 (O_1349,N_8930,N_8717);
and UO_1350 (O_1350,N_8704,N_9875);
or UO_1351 (O_1351,N_8996,N_8457);
and UO_1352 (O_1352,N_9590,N_8617);
or UO_1353 (O_1353,N_8138,N_8580);
nor UO_1354 (O_1354,N_9862,N_8294);
nor UO_1355 (O_1355,N_7582,N_8250);
or UO_1356 (O_1356,N_8567,N_8491);
and UO_1357 (O_1357,N_9424,N_9110);
xor UO_1358 (O_1358,N_9316,N_8023);
nand UO_1359 (O_1359,N_9902,N_8562);
nor UO_1360 (O_1360,N_8692,N_9837);
nor UO_1361 (O_1361,N_8641,N_8176);
and UO_1362 (O_1362,N_8800,N_8162);
xnor UO_1363 (O_1363,N_9930,N_8521);
nor UO_1364 (O_1364,N_8588,N_8294);
or UO_1365 (O_1365,N_7750,N_9426);
nand UO_1366 (O_1366,N_8345,N_9815);
nand UO_1367 (O_1367,N_7922,N_7537);
or UO_1368 (O_1368,N_8107,N_7794);
nand UO_1369 (O_1369,N_9267,N_7618);
or UO_1370 (O_1370,N_8664,N_9869);
nand UO_1371 (O_1371,N_9654,N_8502);
and UO_1372 (O_1372,N_9999,N_8174);
nor UO_1373 (O_1373,N_8659,N_8543);
and UO_1374 (O_1374,N_9099,N_9879);
xnor UO_1375 (O_1375,N_9878,N_8714);
nand UO_1376 (O_1376,N_7988,N_7861);
nor UO_1377 (O_1377,N_9573,N_9751);
or UO_1378 (O_1378,N_9729,N_9725);
and UO_1379 (O_1379,N_7612,N_7815);
or UO_1380 (O_1380,N_9546,N_7821);
and UO_1381 (O_1381,N_7635,N_7819);
or UO_1382 (O_1382,N_8274,N_9316);
nor UO_1383 (O_1383,N_8726,N_8222);
and UO_1384 (O_1384,N_7577,N_9116);
nor UO_1385 (O_1385,N_9834,N_8006);
nand UO_1386 (O_1386,N_8662,N_9306);
or UO_1387 (O_1387,N_8653,N_9563);
nand UO_1388 (O_1388,N_8851,N_9214);
or UO_1389 (O_1389,N_9298,N_7512);
nand UO_1390 (O_1390,N_9305,N_7783);
nand UO_1391 (O_1391,N_9228,N_7968);
nor UO_1392 (O_1392,N_9152,N_8790);
nor UO_1393 (O_1393,N_7723,N_8160);
or UO_1394 (O_1394,N_8962,N_8172);
nand UO_1395 (O_1395,N_8935,N_8905);
nand UO_1396 (O_1396,N_7675,N_7762);
and UO_1397 (O_1397,N_9957,N_7835);
nor UO_1398 (O_1398,N_9474,N_8162);
and UO_1399 (O_1399,N_8790,N_8142);
or UO_1400 (O_1400,N_8007,N_9226);
nor UO_1401 (O_1401,N_8120,N_7947);
nand UO_1402 (O_1402,N_8651,N_8036);
or UO_1403 (O_1403,N_9249,N_9468);
nand UO_1404 (O_1404,N_9277,N_7936);
nor UO_1405 (O_1405,N_7530,N_7883);
nand UO_1406 (O_1406,N_9616,N_9387);
nor UO_1407 (O_1407,N_8121,N_9807);
and UO_1408 (O_1408,N_7658,N_9917);
and UO_1409 (O_1409,N_7987,N_7657);
nor UO_1410 (O_1410,N_8977,N_9724);
and UO_1411 (O_1411,N_9831,N_7550);
nand UO_1412 (O_1412,N_9336,N_8070);
and UO_1413 (O_1413,N_9290,N_7738);
and UO_1414 (O_1414,N_9765,N_9747);
or UO_1415 (O_1415,N_7776,N_9450);
nor UO_1416 (O_1416,N_9543,N_8915);
nand UO_1417 (O_1417,N_8871,N_9077);
nand UO_1418 (O_1418,N_9731,N_9767);
nor UO_1419 (O_1419,N_8382,N_7829);
and UO_1420 (O_1420,N_8618,N_8035);
nor UO_1421 (O_1421,N_9790,N_9900);
or UO_1422 (O_1422,N_8321,N_9334);
or UO_1423 (O_1423,N_9755,N_8529);
and UO_1424 (O_1424,N_8713,N_8773);
and UO_1425 (O_1425,N_8897,N_8336);
nor UO_1426 (O_1426,N_9681,N_9253);
and UO_1427 (O_1427,N_7820,N_9823);
or UO_1428 (O_1428,N_9922,N_8130);
or UO_1429 (O_1429,N_9508,N_7600);
nand UO_1430 (O_1430,N_9861,N_7776);
nor UO_1431 (O_1431,N_9561,N_9531);
or UO_1432 (O_1432,N_8970,N_9077);
or UO_1433 (O_1433,N_9728,N_9047);
and UO_1434 (O_1434,N_8804,N_8387);
or UO_1435 (O_1435,N_9246,N_9755);
and UO_1436 (O_1436,N_9291,N_9180);
nand UO_1437 (O_1437,N_9335,N_7597);
or UO_1438 (O_1438,N_8983,N_9701);
nor UO_1439 (O_1439,N_9449,N_8719);
nor UO_1440 (O_1440,N_8409,N_7580);
or UO_1441 (O_1441,N_8051,N_8385);
or UO_1442 (O_1442,N_8199,N_8628);
nor UO_1443 (O_1443,N_9804,N_9003);
xnor UO_1444 (O_1444,N_9385,N_8891);
and UO_1445 (O_1445,N_8233,N_7691);
nand UO_1446 (O_1446,N_8270,N_7884);
nand UO_1447 (O_1447,N_8093,N_9564);
or UO_1448 (O_1448,N_9392,N_8690);
nor UO_1449 (O_1449,N_7803,N_9979);
or UO_1450 (O_1450,N_9061,N_8152);
or UO_1451 (O_1451,N_8757,N_7835);
and UO_1452 (O_1452,N_9768,N_7531);
and UO_1453 (O_1453,N_8655,N_7590);
and UO_1454 (O_1454,N_8199,N_9652);
nand UO_1455 (O_1455,N_7829,N_9568);
nand UO_1456 (O_1456,N_9374,N_8150);
nor UO_1457 (O_1457,N_8149,N_9039);
or UO_1458 (O_1458,N_8949,N_9425);
and UO_1459 (O_1459,N_9810,N_8459);
nor UO_1460 (O_1460,N_8116,N_8200);
or UO_1461 (O_1461,N_9273,N_7711);
and UO_1462 (O_1462,N_9055,N_8532);
nor UO_1463 (O_1463,N_7672,N_8429);
nor UO_1464 (O_1464,N_7665,N_9381);
and UO_1465 (O_1465,N_9307,N_9090);
and UO_1466 (O_1466,N_7990,N_9270);
nor UO_1467 (O_1467,N_7975,N_8503);
nor UO_1468 (O_1468,N_8170,N_8297);
nor UO_1469 (O_1469,N_8440,N_7718);
nor UO_1470 (O_1470,N_8682,N_7510);
or UO_1471 (O_1471,N_9851,N_9481);
and UO_1472 (O_1472,N_8470,N_7675);
and UO_1473 (O_1473,N_9502,N_9349);
nand UO_1474 (O_1474,N_8167,N_9013);
or UO_1475 (O_1475,N_8692,N_8155);
nand UO_1476 (O_1476,N_7598,N_9731);
nand UO_1477 (O_1477,N_8121,N_7878);
nand UO_1478 (O_1478,N_8298,N_8529);
nand UO_1479 (O_1479,N_9668,N_8217);
nand UO_1480 (O_1480,N_8540,N_9754);
nor UO_1481 (O_1481,N_8597,N_8447);
and UO_1482 (O_1482,N_8427,N_7683);
and UO_1483 (O_1483,N_8363,N_9430);
or UO_1484 (O_1484,N_9802,N_9831);
nor UO_1485 (O_1485,N_8452,N_9825);
and UO_1486 (O_1486,N_9962,N_7847);
nand UO_1487 (O_1487,N_9546,N_8763);
and UO_1488 (O_1488,N_8243,N_7631);
nand UO_1489 (O_1489,N_8454,N_9522);
nor UO_1490 (O_1490,N_9532,N_8215);
or UO_1491 (O_1491,N_8741,N_9556);
and UO_1492 (O_1492,N_8645,N_8761);
nor UO_1493 (O_1493,N_8843,N_8036);
nand UO_1494 (O_1494,N_9304,N_9511);
and UO_1495 (O_1495,N_8337,N_8599);
nand UO_1496 (O_1496,N_8220,N_9783);
nand UO_1497 (O_1497,N_8634,N_9198);
nor UO_1498 (O_1498,N_8372,N_8942);
nor UO_1499 (O_1499,N_7624,N_9054);
endmodule