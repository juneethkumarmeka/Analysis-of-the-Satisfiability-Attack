module basic_750_5000_1000_5_levels_5xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
and U0 (N_0,In_419,In_654);
or U1 (N_1,In_80,In_64);
and U2 (N_2,In_568,In_635);
nor U3 (N_3,In_457,In_28);
nand U4 (N_4,In_733,In_567);
nor U5 (N_5,In_103,In_431);
nand U6 (N_6,In_174,In_686);
and U7 (N_7,In_200,In_328);
nand U8 (N_8,In_475,In_362);
and U9 (N_9,In_44,In_310);
nand U10 (N_10,In_344,In_641);
and U11 (N_11,In_651,In_433);
or U12 (N_12,In_721,In_94);
nor U13 (N_13,In_681,In_560);
nand U14 (N_14,In_519,In_474);
and U15 (N_15,In_77,In_435);
or U16 (N_16,In_525,In_143);
and U17 (N_17,In_26,In_218);
nor U18 (N_18,In_645,In_239);
or U19 (N_19,In_327,In_11);
nor U20 (N_20,In_380,In_219);
or U21 (N_21,In_452,In_570);
xor U22 (N_22,In_450,In_281);
nor U23 (N_23,In_550,In_365);
and U24 (N_24,In_125,In_267);
or U25 (N_25,In_273,In_2);
nor U26 (N_26,In_132,In_366);
nor U27 (N_27,In_27,In_79);
or U28 (N_28,In_677,In_115);
or U29 (N_29,In_159,In_575);
nor U30 (N_30,In_65,In_551);
and U31 (N_31,In_264,In_287);
and U32 (N_32,In_694,In_32);
or U33 (N_33,In_726,In_153);
or U34 (N_34,In_165,In_356);
nand U35 (N_35,In_173,In_675);
nor U36 (N_36,In_34,In_97);
or U37 (N_37,In_361,In_92);
nor U38 (N_38,In_417,In_680);
and U39 (N_39,In_43,In_89);
nand U40 (N_40,In_60,In_322);
or U41 (N_41,In_496,In_478);
nand U42 (N_42,In_701,In_368);
xor U43 (N_43,In_113,In_195);
nand U44 (N_44,In_707,In_81);
xor U45 (N_45,In_737,In_313);
nor U46 (N_46,In_364,In_597);
or U47 (N_47,In_710,In_454);
nand U48 (N_48,In_491,In_42);
and U49 (N_49,In_446,In_449);
nor U50 (N_50,In_352,In_277);
nand U51 (N_51,In_52,In_226);
and U52 (N_52,In_91,In_745);
and U53 (N_53,In_590,In_552);
and U54 (N_54,In_99,In_208);
or U55 (N_55,In_544,In_418);
or U56 (N_56,In_326,In_594);
and U57 (N_57,In_293,In_579);
or U58 (N_58,In_439,In_220);
and U59 (N_59,In_512,In_378);
nor U60 (N_60,In_407,In_718);
nor U61 (N_61,In_600,In_516);
nand U62 (N_62,In_485,In_342);
or U63 (N_63,In_655,In_390);
xor U64 (N_64,In_448,In_319);
nor U65 (N_65,In_347,In_324);
or U66 (N_66,In_129,In_574);
or U67 (N_67,In_16,In_460);
nand U68 (N_68,In_316,In_526);
or U69 (N_69,In_257,In_229);
and U70 (N_70,In_614,In_687);
and U71 (N_71,In_467,In_540);
nor U72 (N_72,In_527,In_705);
or U73 (N_73,In_430,In_628);
xnor U74 (N_74,In_702,In_468);
xor U75 (N_75,In_302,In_217);
nand U76 (N_76,In_397,In_672);
and U77 (N_77,In_695,In_509);
nand U78 (N_78,In_41,In_228);
nor U79 (N_79,In_351,In_375);
nand U80 (N_80,In_154,In_345);
and U81 (N_81,In_533,In_379);
nor U82 (N_82,In_39,In_558);
and U83 (N_83,In_615,In_40);
or U84 (N_84,In_255,In_329);
nand U85 (N_85,In_48,In_522);
nand U86 (N_86,In_679,In_472);
nor U87 (N_87,In_238,In_246);
nand U88 (N_88,In_96,In_507);
nand U89 (N_89,In_160,In_295);
or U90 (N_90,In_384,In_86);
and U91 (N_91,In_740,In_411);
nor U92 (N_92,In_306,In_673);
nand U93 (N_93,In_8,In_725);
and U94 (N_94,In_652,In_688);
or U95 (N_95,In_214,In_684);
nand U96 (N_96,In_206,In_225);
xnor U97 (N_97,In_555,In_339);
or U98 (N_98,In_301,In_172);
or U99 (N_99,In_31,In_330);
or U100 (N_100,In_249,In_331);
nor U101 (N_101,In_501,In_74);
nand U102 (N_102,In_88,In_205);
nand U103 (N_103,In_396,In_294);
and U104 (N_104,In_458,In_481);
or U105 (N_105,In_398,In_196);
and U106 (N_106,In_466,In_489);
nor U107 (N_107,In_631,In_105);
nand U108 (N_108,In_323,In_367);
or U109 (N_109,In_744,In_395);
or U110 (N_110,In_563,In_640);
xnor U111 (N_111,In_711,In_176);
nand U112 (N_112,In_576,In_134);
and U113 (N_113,In_336,In_290);
nor U114 (N_114,In_280,In_199);
xnor U115 (N_115,In_618,In_676);
nor U116 (N_116,In_500,In_167);
nor U117 (N_117,In_646,In_235);
xor U118 (N_118,In_377,In_95);
nor U119 (N_119,In_639,In_469);
or U120 (N_120,In_657,In_498);
or U121 (N_121,In_572,In_423);
and U122 (N_122,In_437,In_538);
or U123 (N_123,In_182,In_545);
xor U124 (N_124,In_170,In_181);
and U125 (N_125,In_162,In_197);
xor U126 (N_126,In_604,In_739);
nand U127 (N_127,In_6,In_237);
or U128 (N_128,In_547,In_282);
or U129 (N_129,In_186,In_633);
or U130 (N_130,In_389,In_497);
nor U131 (N_131,In_494,In_157);
nor U132 (N_132,In_625,In_559);
nor U133 (N_133,In_341,In_297);
nor U134 (N_134,In_506,In_272);
nor U135 (N_135,In_643,In_689);
nor U136 (N_136,In_122,In_296);
or U137 (N_137,In_488,In_135);
and U138 (N_138,In_114,In_401);
nand U139 (N_139,In_57,In_175);
nor U140 (N_140,In_338,In_391);
nand U141 (N_141,In_268,In_127);
or U142 (N_142,In_653,In_265);
and U143 (N_143,In_158,In_748);
nand U144 (N_144,In_82,In_201);
nor U145 (N_145,In_671,In_429);
or U146 (N_146,In_72,In_164);
xnor U147 (N_147,In_514,In_402);
or U148 (N_148,In_300,In_150);
or U149 (N_149,In_566,In_37);
nor U150 (N_150,In_9,In_393);
nand U151 (N_151,In_562,In_17);
xnor U152 (N_152,In_578,In_256);
nor U153 (N_153,In_424,In_586);
and U154 (N_154,In_23,In_678);
and U155 (N_155,In_528,In_589);
nor U156 (N_156,In_470,In_722);
and U157 (N_157,In_253,In_535);
nand U158 (N_158,In_703,In_110);
nor U159 (N_159,In_337,In_656);
or U160 (N_160,In_529,In_732);
nand U161 (N_161,In_148,In_36);
and U162 (N_162,In_691,In_699);
nand U163 (N_163,In_731,In_193);
nor U164 (N_164,In_612,In_325);
nand U165 (N_165,In_479,In_142);
and U166 (N_166,In_664,In_622);
nor U167 (N_167,In_697,In_649);
xor U168 (N_168,In_333,In_119);
and U169 (N_169,In_595,In_388);
and U170 (N_170,In_659,In_582);
nand U171 (N_171,In_569,In_447);
or U172 (N_172,In_444,In_29);
and U173 (N_173,In_236,In_359);
nand U174 (N_174,In_521,In_55);
xor U175 (N_175,In_462,In_598);
or U176 (N_176,In_620,In_719);
or U177 (N_177,In_505,In_62);
or U178 (N_178,In_605,In_240);
nor U179 (N_179,In_156,In_185);
and U180 (N_180,In_416,In_203);
nand U181 (N_181,In_147,In_53);
and U182 (N_182,In_495,In_692);
and U183 (N_183,In_215,In_247);
and U184 (N_184,In_536,In_30);
and U185 (N_185,In_248,In_123);
and U186 (N_186,In_665,In_585);
nand U187 (N_187,In_473,In_285);
nand U188 (N_188,In_627,In_7);
nor U189 (N_189,In_670,In_354);
nand U190 (N_190,In_727,In_106);
or U191 (N_191,In_611,In_145);
nor U192 (N_192,In_262,In_376);
xor U193 (N_193,In_592,In_116);
nand U194 (N_194,In_713,In_374);
or U195 (N_195,In_276,In_685);
nor U196 (N_196,In_21,In_292);
nand U197 (N_197,In_480,In_161);
and U198 (N_198,In_108,In_15);
or U199 (N_199,In_318,In_621);
nor U200 (N_200,In_465,In_71);
nand U201 (N_201,In_392,In_606);
nor U202 (N_202,In_674,In_412);
nor U203 (N_203,In_371,In_171);
nand U204 (N_204,In_549,In_486);
and U205 (N_205,In_245,In_212);
xor U206 (N_206,In_534,In_548);
nand U207 (N_207,In_714,In_67);
and U208 (N_208,In_224,In_211);
or U209 (N_209,In_373,In_487);
or U210 (N_210,In_386,In_73);
xor U211 (N_211,In_149,In_139);
nor U212 (N_212,In_350,In_482);
or U213 (N_213,In_503,In_204);
nand U214 (N_214,In_405,In_138);
and U215 (N_215,In_629,In_434);
or U216 (N_216,In_194,In_510);
nand U217 (N_217,In_613,In_177);
and U218 (N_218,In_729,In_537);
or U219 (N_219,In_413,In_54);
and U220 (N_220,In_422,In_704);
or U221 (N_221,In_133,In_603);
nor U222 (N_222,In_141,In_724);
and U223 (N_223,In_252,In_230);
nor U224 (N_224,In_553,In_298);
xor U225 (N_225,In_308,In_189);
and U226 (N_226,In_24,In_227);
and U227 (N_227,In_144,In_523);
nor U228 (N_228,In_188,In_554);
and U229 (N_229,In_314,In_288);
or U230 (N_230,In_696,In_124);
and U231 (N_231,In_455,In_436);
nor U232 (N_232,In_630,In_573);
nand U233 (N_233,In_637,In_291);
nor U234 (N_234,In_241,In_546);
and U235 (N_235,In_484,In_109);
nand U236 (N_236,In_101,In_5);
nand U237 (N_237,In_168,In_140);
and U238 (N_238,In_394,In_191);
xor U239 (N_239,In_266,In_524);
or U240 (N_240,In_111,In_438);
or U241 (N_241,In_464,In_63);
nor U242 (N_242,In_321,In_187);
xor U243 (N_243,In_209,In_584);
nor U244 (N_244,In_118,In_432);
nor U245 (N_245,In_440,In_299);
or U246 (N_246,In_610,In_504);
xor U247 (N_247,In_409,In_320);
or U248 (N_248,In_84,In_286);
nor U249 (N_249,In_624,In_508);
or U250 (N_250,In_369,In_38);
and U251 (N_251,In_445,In_90);
or U252 (N_252,In_233,In_743);
nand U253 (N_253,In_104,In_210);
or U254 (N_254,In_483,In_642);
and U255 (N_255,In_408,In_511);
nor U256 (N_256,In_68,In_355);
nand U257 (N_257,In_107,In_442);
xnor U258 (N_258,In_131,In_258);
or U259 (N_259,In_541,In_18);
nand U260 (N_260,In_658,In_234);
nand U261 (N_261,In_121,In_735);
nand U262 (N_262,In_530,In_137);
nand U263 (N_263,In_1,In_93);
nand U264 (N_264,In_357,In_564);
nand U265 (N_265,In_499,In_730);
nand U266 (N_266,In_22,In_85);
nand U267 (N_267,In_358,In_202);
or U268 (N_268,In_166,In_542);
nand U269 (N_269,In_83,In_14);
and U270 (N_270,In_593,In_728);
and U271 (N_271,In_619,In_451);
or U272 (N_272,In_117,In_736);
nor U273 (N_273,In_35,In_274);
nand U274 (N_274,In_556,In_179);
or U275 (N_275,In_660,In_647);
nor U276 (N_276,In_66,In_349);
and U277 (N_277,In_78,In_477);
and U278 (N_278,In_155,In_404);
xor U279 (N_279,In_403,In_425);
nand U280 (N_280,In_25,In_539);
nor U281 (N_281,In_311,In_45);
and U282 (N_282,In_588,In_581);
nor U283 (N_283,In_269,In_231);
nand U284 (N_284,In_56,In_463);
nand U285 (N_285,In_120,In_644);
xnor U286 (N_286,In_250,In_98);
nand U287 (N_287,In_662,In_348);
xor U288 (N_288,In_4,In_599);
nor U289 (N_289,In_381,In_259);
xor U290 (N_290,In_683,In_720);
nand U291 (N_291,In_626,In_47);
and U292 (N_292,In_58,In_747);
or U293 (N_293,In_661,In_441);
and U294 (N_294,In_242,In_415);
xnor U295 (N_295,In_609,In_515);
xnor U296 (N_296,In_360,In_741);
or U297 (N_297,In_410,In_532);
nand U298 (N_298,In_580,In_387);
nand U299 (N_299,In_583,In_146);
or U300 (N_300,In_275,In_715);
or U301 (N_301,In_10,In_693);
nand U302 (N_302,In_616,In_283);
nand U303 (N_303,In_243,In_634);
xnor U304 (N_304,In_50,In_623);
nor U305 (N_305,In_700,In_420);
nor U306 (N_306,In_461,In_383);
nor U307 (N_307,In_400,In_19);
or U308 (N_308,In_663,In_363);
nand U309 (N_309,In_638,In_307);
nor U310 (N_310,In_370,In_304);
xor U311 (N_311,In_192,In_577);
nand U312 (N_312,In_561,In_270);
nand U313 (N_313,In_668,In_207);
nand U314 (N_314,In_399,In_87);
nor U315 (N_315,In_492,In_709);
nor U316 (N_316,In_669,In_261);
nand U317 (N_317,In_184,In_602);
nand U318 (N_318,In_608,In_232);
or U319 (N_319,In_49,In_263);
or U320 (N_320,In_667,In_251);
nand U321 (N_321,In_706,In_46);
or U322 (N_322,In_75,In_309);
or U323 (N_323,In_213,In_698);
nor U324 (N_324,In_632,In_601);
nor U325 (N_325,In_617,In_346);
and U326 (N_326,In_650,In_557);
and U327 (N_327,In_278,In_636);
and U328 (N_328,In_428,In_221);
xor U329 (N_329,In_12,In_471);
or U330 (N_330,In_385,In_690);
or U331 (N_331,In_216,In_749);
or U332 (N_332,In_151,In_565);
nor U333 (N_333,In_303,In_260);
or U334 (N_334,In_128,In_738);
nor U335 (N_335,In_335,In_382);
and U336 (N_336,In_682,In_69);
xnor U337 (N_337,In_490,In_305);
and U338 (N_338,In_59,In_152);
nand U339 (N_339,In_0,In_223);
or U340 (N_340,In_244,In_112);
and U341 (N_341,In_543,In_493);
or U342 (N_342,In_648,In_502);
xnor U343 (N_343,In_254,In_61);
nor U344 (N_344,In_317,In_271);
and U345 (N_345,In_100,In_426);
or U346 (N_346,In_20,In_178);
nand U347 (N_347,In_531,In_315);
and U348 (N_348,In_289,In_518);
and U349 (N_349,In_180,In_591);
or U350 (N_350,In_51,In_421);
or U351 (N_351,In_717,In_742);
nand U352 (N_352,In_3,In_708);
and U353 (N_353,In_453,In_169);
nor U354 (N_354,In_406,In_587);
nand U355 (N_355,In_353,In_414);
nor U356 (N_356,In_13,In_513);
nand U357 (N_357,In_126,In_427);
nor U358 (N_358,In_343,In_372);
nor U359 (N_359,In_666,In_596);
and U360 (N_360,In_136,In_716);
or U361 (N_361,In_334,In_190);
xnor U362 (N_362,In_76,In_459);
or U363 (N_363,In_476,In_712);
nand U364 (N_364,In_198,In_312);
and U365 (N_365,In_607,In_70);
or U366 (N_366,In_130,In_340);
and U367 (N_367,In_734,In_102);
and U368 (N_368,In_284,In_332);
nand U369 (N_369,In_520,In_222);
nand U370 (N_370,In_456,In_517);
nand U371 (N_371,In_746,In_723);
or U372 (N_372,In_443,In_279);
and U373 (N_373,In_163,In_183);
nor U374 (N_374,In_33,In_571);
nand U375 (N_375,In_712,In_394);
nand U376 (N_376,In_350,In_5);
nand U377 (N_377,In_461,In_566);
nand U378 (N_378,In_660,In_305);
nor U379 (N_379,In_396,In_547);
and U380 (N_380,In_688,In_119);
nand U381 (N_381,In_347,In_676);
nand U382 (N_382,In_86,In_601);
nor U383 (N_383,In_421,In_66);
nand U384 (N_384,In_291,In_242);
or U385 (N_385,In_73,In_388);
nor U386 (N_386,In_657,In_291);
nor U387 (N_387,In_80,In_624);
xor U388 (N_388,In_376,In_157);
nand U389 (N_389,In_69,In_527);
xnor U390 (N_390,In_412,In_460);
xor U391 (N_391,In_413,In_390);
nand U392 (N_392,In_30,In_502);
and U393 (N_393,In_265,In_626);
nor U394 (N_394,In_152,In_567);
nand U395 (N_395,In_155,In_163);
and U396 (N_396,In_292,In_621);
nor U397 (N_397,In_489,In_529);
or U398 (N_398,In_627,In_57);
and U399 (N_399,In_263,In_134);
nor U400 (N_400,In_488,In_341);
nand U401 (N_401,In_649,In_430);
or U402 (N_402,In_663,In_417);
nand U403 (N_403,In_53,In_487);
and U404 (N_404,In_736,In_242);
nand U405 (N_405,In_267,In_332);
nand U406 (N_406,In_529,In_405);
xor U407 (N_407,In_46,In_11);
or U408 (N_408,In_95,In_240);
nor U409 (N_409,In_156,In_371);
nand U410 (N_410,In_332,In_386);
nand U411 (N_411,In_472,In_717);
and U412 (N_412,In_256,In_528);
and U413 (N_413,In_689,In_453);
or U414 (N_414,In_92,In_303);
or U415 (N_415,In_597,In_264);
nand U416 (N_416,In_657,In_573);
or U417 (N_417,In_42,In_220);
nand U418 (N_418,In_159,In_121);
nand U419 (N_419,In_240,In_513);
nand U420 (N_420,In_100,In_330);
xor U421 (N_421,In_461,In_5);
and U422 (N_422,In_371,In_18);
and U423 (N_423,In_522,In_137);
nor U424 (N_424,In_512,In_257);
xor U425 (N_425,In_612,In_132);
nand U426 (N_426,In_386,In_726);
or U427 (N_427,In_246,In_346);
xnor U428 (N_428,In_346,In_309);
or U429 (N_429,In_130,In_579);
or U430 (N_430,In_493,In_738);
and U431 (N_431,In_43,In_735);
xor U432 (N_432,In_107,In_41);
or U433 (N_433,In_454,In_705);
nor U434 (N_434,In_242,In_564);
or U435 (N_435,In_106,In_476);
nor U436 (N_436,In_476,In_457);
xnor U437 (N_437,In_186,In_595);
xnor U438 (N_438,In_443,In_219);
and U439 (N_439,In_87,In_69);
nand U440 (N_440,In_601,In_508);
and U441 (N_441,In_41,In_486);
nor U442 (N_442,In_622,In_36);
nor U443 (N_443,In_633,In_80);
or U444 (N_444,In_465,In_75);
and U445 (N_445,In_342,In_491);
nor U446 (N_446,In_92,In_337);
and U447 (N_447,In_415,In_19);
nor U448 (N_448,In_565,In_372);
nand U449 (N_449,In_514,In_308);
nor U450 (N_450,In_277,In_635);
nand U451 (N_451,In_619,In_201);
and U452 (N_452,In_233,In_272);
nor U453 (N_453,In_574,In_689);
xnor U454 (N_454,In_555,In_661);
nand U455 (N_455,In_145,In_29);
or U456 (N_456,In_204,In_183);
nand U457 (N_457,In_8,In_298);
nor U458 (N_458,In_100,In_673);
or U459 (N_459,In_700,In_670);
or U460 (N_460,In_165,In_208);
nand U461 (N_461,In_628,In_651);
nand U462 (N_462,In_5,In_573);
nand U463 (N_463,In_94,In_513);
or U464 (N_464,In_173,In_429);
nand U465 (N_465,In_226,In_63);
xor U466 (N_466,In_260,In_387);
and U467 (N_467,In_376,In_103);
or U468 (N_468,In_530,In_45);
xor U469 (N_469,In_671,In_481);
and U470 (N_470,In_722,In_684);
and U471 (N_471,In_297,In_230);
and U472 (N_472,In_274,In_276);
nand U473 (N_473,In_747,In_196);
nand U474 (N_474,In_518,In_557);
and U475 (N_475,In_133,In_570);
and U476 (N_476,In_521,In_626);
and U477 (N_477,In_211,In_99);
or U478 (N_478,In_294,In_28);
and U479 (N_479,In_32,In_728);
and U480 (N_480,In_645,In_582);
and U481 (N_481,In_244,In_485);
nand U482 (N_482,In_578,In_461);
and U483 (N_483,In_725,In_446);
and U484 (N_484,In_85,In_395);
nand U485 (N_485,In_426,In_367);
or U486 (N_486,In_470,In_169);
nor U487 (N_487,In_601,In_133);
xor U488 (N_488,In_519,In_276);
nor U489 (N_489,In_579,In_729);
xor U490 (N_490,In_744,In_564);
or U491 (N_491,In_204,In_304);
xor U492 (N_492,In_240,In_625);
and U493 (N_493,In_211,In_398);
nor U494 (N_494,In_485,In_501);
or U495 (N_495,In_556,In_662);
or U496 (N_496,In_205,In_427);
and U497 (N_497,In_337,In_695);
nand U498 (N_498,In_539,In_197);
and U499 (N_499,In_277,In_330);
nor U500 (N_500,In_737,In_460);
or U501 (N_501,In_634,In_413);
and U502 (N_502,In_470,In_315);
nand U503 (N_503,In_134,In_455);
or U504 (N_504,In_409,In_739);
xnor U505 (N_505,In_307,In_48);
or U506 (N_506,In_55,In_102);
and U507 (N_507,In_213,In_386);
and U508 (N_508,In_346,In_404);
or U509 (N_509,In_521,In_719);
and U510 (N_510,In_534,In_697);
or U511 (N_511,In_534,In_683);
or U512 (N_512,In_514,In_377);
nand U513 (N_513,In_24,In_9);
nor U514 (N_514,In_537,In_211);
nand U515 (N_515,In_23,In_708);
or U516 (N_516,In_309,In_352);
or U517 (N_517,In_582,In_496);
and U518 (N_518,In_384,In_351);
and U519 (N_519,In_714,In_50);
and U520 (N_520,In_612,In_218);
or U521 (N_521,In_267,In_87);
nand U522 (N_522,In_29,In_665);
nand U523 (N_523,In_481,In_379);
nand U524 (N_524,In_560,In_65);
nor U525 (N_525,In_312,In_573);
or U526 (N_526,In_535,In_482);
nor U527 (N_527,In_635,In_431);
and U528 (N_528,In_348,In_571);
nor U529 (N_529,In_476,In_361);
nand U530 (N_530,In_620,In_737);
nor U531 (N_531,In_408,In_88);
nor U532 (N_532,In_577,In_477);
nand U533 (N_533,In_326,In_648);
or U534 (N_534,In_588,In_257);
nor U535 (N_535,In_502,In_403);
xor U536 (N_536,In_312,In_739);
and U537 (N_537,In_118,In_106);
xor U538 (N_538,In_124,In_153);
or U539 (N_539,In_374,In_87);
nand U540 (N_540,In_0,In_396);
xnor U541 (N_541,In_220,In_445);
or U542 (N_542,In_393,In_519);
nor U543 (N_543,In_352,In_624);
xor U544 (N_544,In_454,In_149);
nand U545 (N_545,In_164,In_138);
nor U546 (N_546,In_625,In_641);
xor U547 (N_547,In_123,In_676);
xnor U548 (N_548,In_344,In_302);
and U549 (N_549,In_336,In_638);
nor U550 (N_550,In_440,In_48);
or U551 (N_551,In_732,In_307);
nor U552 (N_552,In_417,In_215);
or U553 (N_553,In_748,In_39);
or U554 (N_554,In_743,In_293);
nand U555 (N_555,In_288,In_191);
nand U556 (N_556,In_418,In_353);
and U557 (N_557,In_87,In_585);
or U558 (N_558,In_224,In_366);
nand U559 (N_559,In_695,In_37);
and U560 (N_560,In_106,In_126);
nand U561 (N_561,In_680,In_632);
and U562 (N_562,In_660,In_632);
or U563 (N_563,In_558,In_262);
nand U564 (N_564,In_563,In_296);
nand U565 (N_565,In_393,In_513);
nand U566 (N_566,In_219,In_480);
and U567 (N_567,In_212,In_60);
and U568 (N_568,In_558,In_187);
nand U569 (N_569,In_273,In_313);
xor U570 (N_570,In_51,In_492);
nand U571 (N_571,In_114,In_593);
nor U572 (N_572,In_212,In_387);
nor U573 (N_573,In_418,In_532);
nand U574 (N_574,In_452,In_153);
nor U575 (N_575,In_433,In_523);
nand U576 (N_576,In_112,In_743);
nand U577 (N_577,In_108,In_722);
and U578 (N_578,In_461,In_119);
and U579 (N_579,In_132,In_263);
nor U580 (N_580,In_167,In_293);
nor U581 (N_581,In_187,In_278);
nand U582 (N_582,In_104,In_691);
or U583 (N_583,In_580,In_633);
nand U584 (N_584,In_127,In_79);
or U585 (N_585,In_89,In_85);
nand U586 (N_586,In_429,In_523);
or U587 (N_587,In_195,In_329);
nand U588 (N_588,In_1,In_707);
or U589 (N_589,In_320,In_651);
nand U590 (N_590,In_240,In_111);
or U591 (N_591,In_682,In_349);
or U592 (N_592,In_676,In_302);
xor U593 (N_593,In_189,In_311);
nand U594 (N_594,In_14,In_0);
and U595 (N_595,In_704,In_121);
nand U596 (N_596,In_615,In_579);
xor U597 (N_597,In_532,In_578);
nand U598 (N_598,In_432,In_275);
nand U599 (N_599,In_366,In_3);
nor U600 (N_600,In_619,In_272);
nand U601 (N_601,In_301,In_620);
nand U602 (N_602,In_143,In_364);
and U603 (N_603,In_742,In_282);
nand U604 (N_604,In_731,In_353);
or U605 (N_605,In_311,In_564);
nand U606 (N_606,In_400,In_107);
and U607 (N_607,In_128,In_323);
nor U608 (N_608,In_688,In_302);
nor U609 (N_609,In_702,In_446);
xor U610 (N_610,In_209,In_419);
and U611 (N_611,In_255,In_725);
xnor U612 (N_612,In_442,In_214);
xnor U613 (N_613,In_623,In_275);
xnor U614 (N_614,In_7,In_198);
nor U615 (N_615,In_321,In_562);
nand U616 (N_616,In_145,In_211);
xnor U617 (N_617,In_468,In_426);
nand U618 (N_618,In_382,In_411);
nand U619 (N_619,In_179,In_508);
and U620 (N_620,In_711,In_147);
nor U621 (N_621,In_399,In_551);
nand U622 (N_622,In_197,In_93);
or U623 (N_623,In_726,In_691);
nor U624 (N_624,In_369,In_14);
nor U625 (N_625,In_57,In_182);
and U626 (N_626,In_732,In_248);
or U627 (N_627,In_226,In_488);
nand U628 (N_628,In_714,In_716);
xor U629 (N_629,In_347,In_514);
nor U630 (N_630,In_440,In_271);
nand U631 (N_631,In_3,In_582);
and U632 (N_632,In_304,In_508);
nor U633 (N_633,In_30,In_293);
nand U634 (N_634,In_35,In_376);
or U635 (N_635,In_452,In_679);
nor U636 (N_636,In_524,In_102);
or U637 (N_637,In_34,In_594);
or U638 (N_638,In_520,In_152);
or U639 (N_639,In_715,In_314);
nor U640 (N_640,In_749,In_188);
nand U641 (N_641,In_172,In_601);
nor U642 (N_642,In_474,In_432);
nor U643 (N_643,In_421,In_2);
or U644 (N_644,In_278,In_443);
nor U645 (N_645,In_502,In_674);
or U646 (N_646,In_52,In_706);
nand U647 (N_647,In_530,In_108);
nor U648 (N_648,In_32,In_36);
nor U649 (N_649,In_414,In_421);
nand U650 (N_650,In_447,In_77);
or U651 (N_651,In_735,In_45);
xor U652 (N_652,In_50,In_456);
nor U653 (N_653,In_459,In_219);
and U654 (N_654,In_444,In_361);
or U655 (N_655,In_65,In_138);
nor U656 (N_656,In_19,In_298);
and U657 (N_657,In_609,In_391);
xnor U658 (N_658,In_316,In_455);
nor U659 (N_659,In_585,In_410);
nor U660 (N_660,In_510,In_232);
nor U661 (N_661,In_709,In_178);
and U662 (N_662,In_106,In_373);
nor U663 (N_663,In_126,In_322);
nor U664 (N_664,In_232,In_453);
and U665 (N_665,In_72,In_120);
or U666 (N_666,In_342,In_334);
and U667 (N_667,In_233,In_711);
or U668 (N_668,In_258,In_617);
nand U669 (N_669,In_87,In_679);
and U670 (N_670,In_397,In_438);
or U671 (N_671,In_481,In_512);
or U672 (N_672,In_454,In_37);
nor U673 (N_673,In_536,In_260);
and U674 (N_674,In_408,In_46);
nand U675 (N_675,In_407,In_675);
nor U676 (N_676,In_553,In_341);
or U677 (N_677,In_481,In_362);
or U678 (N_678,In_679,In_689);
or U679 (N_679,In_568,In_394);
and U680 (N_680,In_526,In_22);
nand U681 (N_681,In_107,In_678);
nand U682 (N_682,In_2,In_118);
nand U683 (N_683,In_496,In_378);
or U684 (N_684,In_410,In_2);
nand U685 (N_685,In_28,In_552);
and U686 (N_686,In_504,In_508);
nand U687 (N_687,In_594,In_448);
nand U688 (N_688,In_669,In_248);
and U689 (N_689,In_328,In_705);
or U690 (N_690,In_58,In_693);
nor U691 (N_691,In_625,In_551);
nor U692 (N_692,In_154,In_587);
nand U693 (N_693,In_264,In_748);
nor U694 (N_694,In_101,In_698);
nor U695 (N_695,In_682,In_514);
nand U696 (N_696,In_410,In_289);
nand U697 (N_697,In_595,In_428);
nand U698 (N_698,In_518,In_359);
or U699 (N_699,In_195,In_352);
or U700 (N_700,In_670,In_427);
and U701 (N_701,In_281,In_272);
nor U702 (N_702,In_623,In_539);
nor U703 (N_703,In_36,In_584);
or U704 (N_704,In_161,In_414);
nor U705 (N_705,In_123,In_200);
nand U706 (N_706,In_678,In_464);
or U707 (N_707,In_402,In_73);
nor U708 (N_708,In_491,In_415);
xor U709 (N_709,In_52,In_584);
xor U710 (N_710,In_718,In_595);
nand U711 (N_711,In_538,In_576);
nand U712 (N_712,In_10,In_589);
and U713 (N_713,In_595,In_248);
and U714 (N_714,In_75,In_163);
nor U715 (N_715,In_571,In_110);
nand U716 (N_716,In_395,In_376);
and U717 (N_717,In_472,In_477);
or U718 (N_718,In_490,In_134);
and U719 (N_719,In_572,In_313);
or U720 (N_720,In_309,In_553);
or U721 (N_721,In_43,In_338);
nor U722 (N_722,In_296,In_704);
and U723 (N_723,In_371,In_1);
xnor U724 (N_724,In_332,In_395);
nand U725 (N_725,In_468,In_84);
nor U726 (N_726,In_352,In_247);
nor U727 (N_727,In_226,In_503);
nand U728 (N_728,In_418,In_566);
and U729 (N_729,In_568,In_82);
and U730 (N_730,In_212,In_76);
and U731 (N_731,In_142,In_728);
nor U732 (N_732,In_606,In_457);
or U733 (N_733,In_506,In_322);
and U734 (N_734,In_48,In_587);
or U735 (N_735,In_278,In_378);
and U736 (N_736,In_267,In_659);
or U737 (N_737,In_139,In_658);
or U738 (N_738,In_138,In_327);
nor U739 (N_739,In_83,In_394);
nor U740 (N_740,In_674,In_279);
nor U741 (N_741,In_344,In_461);
nand U742 (N_742,In_61,In_221);
and U743 (N_743,In_398,In_395);
and U744 (N_744,In_639,In_537);
xor U745 (N_745,In_557,In_214);
and U746 (N_746,In_472,In_667);
xnor U747 (N_747,In_396,In_546);
xor U748 (N_748,In_224,In_110);
or U749 (N_749,In_279,In_644);
nor U750 (N_750,In_93,In_343);
xor U751 (N_751,In_501,In_30);
nand U752 (N_752,In_126,In_749);
and U753 (N_753,In_283,In_259);
xnor U754 (N_754,In_672,In_48);
nor U755 (N_755,In_363,In_212);
nor U756 (N_756,In_271,In_120);
and U757 (N_757,In_255,In_309);
xor U758 (N_758,In_726,In_245);
or U759 (N_759,In_726,In_303);
nand U760 (N_760,In_244,In_459);
nand U761 (N_761,In_153,In_588);
and U762 (N_762,In_408,In_563);
nand U763 (N_763,In_154,In_544);
and U764 (N_764,In_135,In_253);
or U765 (N_765,In_490,In_181);
nor U766 (N_766,In_214,In_10);
nor U767 (N_767,In_174,In_732);
or U768 (N_768,In_694,In_212);
or U769 (N_769,In_694,In_629);
nor U770 (N_770,In_267,In_724);
or U771 (N_771,In_8,In_93);
nand U772 (N_772,In_557,In_34);
xor U773 (N_773,In_325,In_428);
or U774 (N_774,In_419,In_27);
or U775 (N_775,In_714,In_271);
xnor U776 (N_776,In_733,In_540);
nor U777 (N_777,In_400,In_67);
nand U778 (N_778,In_289,In_735);
or U779 (N_779,In_203,In_631);
nand U780 (N_780,In_78,In_289);
and U781 (N_781,In_27,In_617);
or U782 (N_782,In_590,In_478);
and U783 (N_783,In_280,In_516);
nand U784 (N_784,In_153,In_590);
and U785 (N_785,In_711,In_291);
nand U786 (N_786,In_501,In_297);
nand U787 (N_787,In_412,In_687);
or U788 (N_788,In_696,In_225);
nor U789 (N_789,In_79,In_131);
xnor U790 (N_790,In_30,In_32);
xnor U791 (N_791,In_279,In_718);
nand U792 (N_792,In_75,In_460);
or U793 (N_793,In_365,In_437);
nor U794 (N_794,In_144,In_491);
and U795 (N_795,In_562,In_373);
xnor U796 (N_796,In_0,In_191);
nor U797 (N_797,In_389,In_721);
or U798 (N_798,In_316,In_31);
or U799 (N_799,In_311,In_627);
nor U800 (N_800,In_63,In_722);
or U801 (N_801,In_204,In_715);
nor U802 (N_802,In_279,In_286);
or U803 (N_803,In_203,In_73);
xor U804 (N_804,In_419,In_379);
nor U805 (N_805,In_17,In_34);
nor U806 (N_806,In_262,In_321);
nand U807 (N_807,In_152,In_703);
or U808 (N_808,In_288,In_400);
and U809 (N_809,In_616,In_606);
nor U810 (N_810,In_624,In_366);
nor U811 (N_811,In_661,In_330);
or U812 (N_812,In_350,In_485);
nor U813 (N_813,In_337,In_1);
and U814 (N_814,In_518,In_385);
xor U815 (N_815,In_24,In_571);
and U816 (N_816,In_314,In_662);
xnor U817 (N_817,In_474,In_489);
xor U818 (N_818,In_688,In_216);
and U819 (N_819,In_735,In_58);
and U820 (N_820,In_204,In_297);
nand U821 (N_821,In_487,In_149);
nor U822 (N_822,In_93,In_67);
xnor U823 (N_823,In_525,In_14);
nand U824 (N_824,In_263,In_335);
nor U825 (N_825,In_613,In_371);
or U826 (N_826,In_191,In_61);
nand U827 (N_827,In_20,In_592);
or U828 (N_828,In_524,In_423);
and U829 (N_829,In_686,In_269);
nand U830 (N_830,In_552,In_746);
or U831 (N_831,In_151,In_622);
and U832 (N_832,In_480,In_703);
or U833 (N_833,In_229,In_299);
or U834 (N_834,In_206,In_257);
nor U835 (N_835,In_560,In_725);
nand U836 (N_836,In_39,In_556);
and U837 (N_837,In_53,In_445);
nor U838 (N_838,In_686,In_455);
nand U839 (N_839,In_686,In_457);
nor U840 (N_840,In_583,In_239);
and U841 (N_841,In_711,In_714);
xor U842 (N_842,In_249,In_419);
or U843 (N_843,In_78,In_170);
or U844 (N_844,In_351,In_647);
nand U845 (N_845,In_470,In_741);
nand U846 (N_846,In_257,In_98);
nand U847 (N_847,In_53,In_73);
nand U848 (N_848,In_668,In_335);
and U849 (N_849,In_568,In_267);
nand U850 (N_850,In_308,In_674);
or U851 (N_851,In_146,In_587);
xor U852 (N_852,In_134,In_728);
or U853 (N_853,In_571,In_182);
or U854 (N_854,In_3,In_394);
nand U855 (N_855,In_73,In_275);
nand U856 (N_856,In_371,In_152);
and U857 (N_857,In_213,In_611);
or U858 (N_858,In_177,In_242);
nand U859 (N_859,In_391,In_425);
nand U860 (N_860,In_1,In_723);
nand U861 (N_861,In_113,In_48);
and U862 (N_862,In_663,In_681);
and U863 (N_863,In_28,In_515);
nand U864 (N_864,In_224,In_162);
and U865 (N_865,In_328,In_134);
and U866 (N_866,In_743,In_18);
nor U867 (N_867,In_12,In_636);
or U868 (N_868,In_584,In_445);
and U869 (N_869,In_521,In_34);
xnor U870 (N_870,In_204,In_360);
nand U871 (N_871,In_250,In_298);
nor U872 (N_872,In_131,In_373);
xnor U873 (N_873,In_4,In_624);
or U874 (N_874,In_198,In_508);
or U875 (N_875,In_746,In_32);
and U876 (N_876,In_472,In_497);
and U877 (N_877,In_328,In_601);
nand U878 (N_878,In_626,In_544);
or U879 (N_879,In_259,In_732);
or U880 (N_880,In_331,In_284);
or U881 (N_881,In_335,In_272);
xnor U882 (N_882,In_611,In_587);
or U883 (N_883,In_16,In_181);
nand U884 (N_884,In_235,In_352);
or U885 (N_885,In_663,In_357);
xor U886 (N_886,In_134,In_152);
nor U887 (N_887,In_579,In_72);
or U888 (N_888,In_112,In_255);
nor U889 (N_889,In_369,In_418);
nand U890 (N_890,In_112,In_178);
or U891 (N_891,In_79,In_443);
nor U892 (N_892,In_353,In_226);
nand U893 (N_893,In_114,In_664);
nand U894 (N_894,In_98,In_715);
and U895 (N_895,In_549,In_660);
or U896 (N_896,In_30,In_484);
nand U897 (N_897,In_251,In_625);
or U898 (N_898,In_741,In_552);
or U899 (N_899,In_523,In_496);
nand U900 (N_900,In_643,In_268);
or U901 (N_901,In_59,In_297);
and U902 (N_902,In_314,In_417);
nand U903 (N_903,In_723,In_186);
nand U904 (N_904,In_171,In_388);
nor U905 (N_905,In_165,In_220);
nor U906 (N_906,In_291,In_397);
and U907 (N_907,In_509,In_291);
or U908 (N_908,In_292,In_586);
and U909 (N_909,In_4,In_144);
and U910 (N_910,In_10,In_478);
xor U911 (N_911,In_363,In_536);
nor U912 (N_912,In_500,In_612);
nand U913 (N_913,In_140,In_306);
or U914 (N_914,In_623,In_213);
and U915 (N_915,In_724,In_346);
or U916 (N_916,In_434,In_204);
xor U917 (N_917,In_448,In_115);
nand U918 (N_918,In_697,In_745);
or U919 (N_919,In_539,In_628);
nand U920 (N_920,In_106,In_686);
and U921 (N_921,In_138,In_570);
and U922 (N_922,In_569,In_141);
or U923 (N_923,In_666,In_640);
nor U924 (N_924,In_442,In_264);
nor U925 (N_925,In_594,In_405);
xor U926 (N_926,In_170,In_258);
or U927 (N_927,In_33,In_211);
xor U928 (N_928,In_655,In_242);
nor U929 (N_929,In_691,In_649);
nor U930 (N_930,In_445,In_401);
and U931 (N_931,In_700,In_16);
xnor U932 (N_932,In_658,In_232);
or U933 (N_933,In_277,In_7);
or U934 (N_934,In_634,In_346);
or U935 (N_935,In_320,In_366);
nor U936 (N_936,In_554,In_267);
and U937 (N_937,In_612,In_433);
or U938 (N_938,In_333,In_701);
and U939 (N_939,In_190,In_653);
nor U940 (N_940,In_631,In_494);
nand U941 (N_941,In_564,In_359);
or U942 (N_942,In_638,In_4);
nand U943 (N_943,In_33,In_126);
xnor U944 (N_944,In_584,In_587);
and U945 (N_945,In_394,In_409);
nand U946 (N_946,In_472,In_532);
nor U947 (N_947,In_457,In_627);
nand U948 (N_948,In_366,In_490);
nand U949 (N_949,In_114,In_635);
nand U950 (N_950,In_727,In_6);
and U951 (N_951,In_183,In_648);
nand U952 (N_952,In_27,In_552);
nand U953 (N_953,In_617,In_545);
or U954 (N_954,In_64,In_370);
nand U955 (N_955,In_111,In_625);
and U956 (N_956,In_704,In_394);
and U957 (N_957,In_367,In_519);
nor U958 (N_958,In_610,In_114);
and U959 (N_959,In_612,In_276);
xnor U960 (N_960,In_407,In_154);
nand U961 (N_961,In_552,In_247);
and U962 (N_962,In_617,In_228);
nand U963 (N_963,In_577,In_490);
or U964 (N_964,In_569,In_113);
nand U965 (N_965,In_468,In_444);
nor U966 (N_966,In_321,In_235);
and U967 (N_967,In_503,In_627);
nand U968 (N_968,In_415,In_456);
xor U969 (N_969,In_470,In_591);
or U970 (N_970,In_131,In_468);
or U971 (N_971,In_152,In_698);
or U972 (N_972,In_58,In_437);
nor U973 (N_973,In_68,In_261);
or U974 (N_974,In_434,In_601);
nand U975 (N_975,In_246,In_269);
and U976 (N_976,In_535,In_467);
nor U977 (N_977,In_11,In_432);
nor U978 (N_978,In_32,In_154);
xor U979 (N_979,In_663,In_273);
or U980 (N_980,In_103,In_400);
nor U981 (N_981,In_411,In_91);
or U982 (N_982,In_395,In_631);
or U983 (N_983,In_606,In_198);
nand U984 (N_984,In_520,In_518);
nand U985 (N_985,In_34,In_398);
nand U986 (N_986,In_413,In_378);
and U987 (N_987,In_367,In_44);
and U988 (N_988,In_137,In_409);
nor U989 (N_989,In_276,In_207);
nand U990 (N_990,In_669,In_222);
or U991 (N_991,In_287,In_689);
and U992 (N_992,In_372,In_611);
or U993 (N_993,In_427,In_715);
nand U994 (N_994,In_342,In_674);
nand U995 (N_995,In_700,In_678);
or U996 (N_996,In_693,In_25);
nand U997 (N_997,In_287,In_529);
nor U998 (N_998,In_412,In_211);
or U999 (N_999,In_722,In_278);
xnor U1000 (N_1000,N_427,N_682);
and U1001 (N_1001,N_71,N_0);
xnor U1002 (N_1002,N_65,N_401);
or U1003 (N_1003,N_149,N_463);
xor U1004 (N_1004,N_569,N_482);
and U1005 (N_1005,N_827,N_756);
nor U1006 (N_1006,N_155,N_951);
nor U1007 (N_1007,N_672,N_646);
or U1008 (N_1008,N_189,N_285);
nand U1009 (N_1009,N_616,N_791);
or U1010 (N_1010,N_859,N_941);
nand U1011 (N_1011,N_627,N_478);
nor U1012 (N_1012,N_954,N_28);
xnor U1013 (N_1013,N_665,N_464);
or U1014 (N_1014,N_391,N_146);
nand U1015 (N_1015,N_380,N_303);
nor U1016 (N_1016,N_7,N_499);
nor U1017 (N_1017,N_578,N_563);
or U1018 (N_1018,N_789,N_233);
or U1019 (N_1019,N_943,N_89);
nor U1020 (N_1020,N_144,N_322);
nor U1021 (N_1021,N_942,N_436);
or U1022 (N_1022,N_325,N_449);
or U1023 (N_1023,N_535,N_444);
nor U1024 (N_1024,N_680,N_57);
and U1025 (N_1025,N_767,N_892);
nor U1026 (N_1026,N_784,N_424);
and U1027 (N_1027,N_173,N_925);
and U1028 (N_1028,N_373,N_824);
xor U1029 (N_1029,N_504,N_485);
nand U1030 (N_1030,N_126,N_640);
nor U1031 (N_1031,N_545,N_678);
or U1032 (N_1032,N_390,N_918);
nor U1033 (N_1033,N_115,N_377);
nor U1034 (N_1034,N_240,N_817);
and U1035 (N_1035,N_628,N_602);
and U1036 (N_1036,N_119,N_281);
nand U1037 (N_1037,N_739,N_447);
nand U1038 (N_1038,N_179,N_656);
or U1039 (N_1039,N_592,N_333);
or U1040 (N_1040,N_428,N_572);
or U1041 (N_1041,N_435,N_429);
and U1042 (N_1042,N_216,N_777);
xnor U1043 (N_1043,N_68,N_22);
nor U1044 (N_1044,N_721,N_979);
nand U1045 (N_1045,N_417,N_465);
or U1046 (N_1046,N_225,N_278);
nand U1047 (N_1047,N_926,N_663);
nor U1048 (N_1048,N_669,N_700);
xor U1049 (N_1049,N_127,N_116);
and U1050 (N_1050,N_922,N_612);
or U1051 (N_1051,N_154,N_328);
nor U1052 (N_1052,N_272,N_714);
nor U1053 (N_1053,N_555,N_691);
nor U1054 (N_1054,N_99,N_981);
or U1055 (N_1055,N_805,N_245);
xor U1056 (N_1056,N_101,N_198);
or U1057 (N_1057,N_75,N_5);
and U1058 (N_1058,N_176,N_354);
or U1059 (N_1059,N_566,N_231);
nor U1060 (N_1060,N_654,N_120);
xor U1061 (N_1061,N_746,N_630);
or U1062 (N_1062,N_603,N_413);
and U1063 (N_1063,N_871,N_736);
and U1064 (N_1064,N_802,N_58);
xnor U1065 (N_1065,N_431,N_929);
nand U1066 (N_1066,N_617,N_803);
or U1067 (N_1067,N_192,N_526);
or U1068 (N_1068,N_542,N_765);
xor U1069 (N_1069,N_170,N_534);
or U1070 (N_1070,N_622,N_423);
and U1071 (N_1071,N_912,N_932);
nor U1072 (N_1072,N_34,N_952);
and U1073 (N_1073,N_600,N_341);
nor U1074 (N_1074,N_843,N_324);
nor U1075 (N_1075,N_226,N_2);
nand U1076 (N_1076,N_854,N_122);
nand U1077 (N_1077,N_171,N_206);
and U1078 (N_1078,N_598,N_456);
or U1079 (N_1079,N_904,N_106);
xnor U1080 (N_1080,N_883,N_561);
nor U1081 (N_1081,N_634,N_906);
or U1082 (N_1082,N_840,N_232);
xor U1083 (N_1083,N_987,N_933);
nand U1084 (N_1084,N_402,N_426);
nor U1085 (N_1085,N_406,N_935);
or U1086 (N_1086,N_317,N_410);
nor U1087 (N_1087,N_610,N_381);
nand U1088 (N_1088,N_78,N_698);
nor U1089 (N_1089,N_386,N_481);
nand U1090 (N_1090,N_894,N_946);
nand U1091 (N_1091,N_641,N_543);
nor U1092 (N_1092,N_919,N_55);
nor U1093 (N_1093,N_183,N_974);
nor U1094 (N_1094,N_1,N_438);
or U1095 (N_1095,N_15,N_4);
nor U1096 (N_1096,N_108,N_350);
xor U1097 (N_1097,N_313,N_755);
nand U1098 (N_1098,N_923,N_342);
nor U1099 (N_1099,N_897,N_114);
and U1100 (N_1100,N_418,N_597);
or U1101 (N_1101,N_732,N_666);
or U1102 (N_1102,N_46,N_551);
nor U1103 (N_1103,N_934,N_728);
nor U1104 (N_1104,N_707,N_227);
nand U1105 (N_1105,N_422,N_986);
and U1106 (N_1106,N_331,N_409);
nor U1107 (N_1107,N_506,N_957);
nor U1108 (N_1108,N_706,N_584);
and U1109 (N_1109,N_743,N_870);
nand U1110 (N_1110,N_441,N_488);
nand U1111 (N_1111,N_270,N_782);
nand U1112 (N_1112,N_754,N_967);
xor U1113 (N_1113,N_913,N_443);
or U1114 (N_1114,N_87,N_515);
or U1115 (N_1115,N_604,N_924);
nand U1116 (N_1116,N_236,N_958);
nand U1117 (N_1117,N_693,N_93);
and U1118 (N_1118,N_964,N_780);
xnor U1119 (N_1119,N_623,N_838);
and U1120 (N_1120,N_970,N_667);
or U1121 (N_1121,N_549,N_833);
or U1122 (N_1122,N_73,N_588);
and U1123 (N_1123,N_483,N_959);
nor U1124 (N_1124,N_512,N_842);
and U1125 (N_1125,N_692,N_294);
and U1126 (N_1126,N_52,N_117);
and U1127 (N_1127,N_845,N_676);
nand U1128 (N_1128,N_375,N_983);
nor U1129 (N_1129,N_397,N_237);
nor U1130 (N_1130,N_14,N_865);
and U1131 (N_1131,N_786,N_323);
or U1132 (N_1132,N_168,N_374);
and U1133 (N_1133,N_813,N_914);
nor U1134 (N_1134,N_516,N_971);
or U1135 (N_1135,N_948,N_265);
nand U1136 (N_1136,N_775,N_234);
xnor U1137 (N_1137,N_367,N_460);
and U1138 (N_1138,N_212,N_20);
nand U1139 (N_1139,N_383,N_498);
or U1140 (N_1140,N_857,N_348);
nand U1141 (N_1141,N_306,N_927);
nor U1142 (N_1142,N_880,N_528);
or U1143 (N_1143,N_276,N_205);
nand U1144 (N_1144,N_66,N_82);
nand U1145 (N_1145,N_886,N_993);
nor U1146 (N_1146,N_379,N_243);
nand U1147 (N_1147,N_875,N_560);
and U1148 (N_1148,N_486,N_586);
or U1149 (N_1149,N_162,N_972);
nor U1150 (N_1150,N_961,N_411);
or U1151 (N_1151,N_188,N_518);
nand U1152 (N_1152,N_257,N_21);
nor U1153 (N_1153,N_662,N_302);
nand U1154 (N_1154,N_466,N_445);
nand U1155 (N_1155,N_163,N_79);
nor U1156 (N_1156,N_420,N_30);
nor U1157 (N_1157,N_145,N_214);
nand U1158 (N_1158,N_585,N_25);
xor U1159 (N_1159,N_249,N_361);
and U1160 (N_1160,N_928,N_42);
nor U1161 (N_1161,N_131,N_36);
nor U1162 (N_1162,N_384,N_157);
nand U1163 (N_1163,N_292,N_98);
nor U1164 (N_1164,N_267,N_547);
nor U1165 (N_1165,N_264,N_32);
or U1166 (N_1166,N_757,N_242);
and U1167 (N_1167,N_91,N_901);
nand U1168 (N_1168,N_621,N_844);
nand U1169 (N_1169,N_273,N_658);
nand U1170 (N_1170,N_694,N_29);
nor U1171 (N_1171,N_989,N_363);
nand U1172 (N_1172,N_811,N_439);
nand U1173 (N_1173,N_23,N_151);
nor U1174 (N_1174,N_864,N_856);
or U1175 (N_1175,N_858,N_320);
nand U1176 (N_1176,N_920,N_262);
nand U1177 (N_1177,N_741,N_175);
nand U1178 (N_1178,N_810,N_56);
nor U1179 (N_1179,N_102,N_31);
and U1180 (N_1180,N_725,N_636);
nand U1181 (N_1181,N_152,N_298);
and U1182 (N_1182,N_148,N_679);
nand U1183 (N_1183,N_724,N_462);
nand U1184 (N_1184,N_812,N_13);
nor U1185 (N_1185,N_197,N_289);
nand U1186 (N_1186,N_546,N_795);
nor U1187 (N_1187,N_771,N_105);
nor U1188 (N_1188,N_657,N_966);
or U1189 (N_1189,N_11,N_531);
nor U1190 (N_1190,N_329,N_12);
nor U1191 (N_1191,N_508,N_147);
or U1192 (N_1192,N_254,N_10);
and U1193 (N_1193,N_873,N_635);
and U1194 (N_1194,N_632,N_358);
nor U1195 (N_1195,N_737,N_203);
nand U1196 (N_1196,N_454,N_394);
nor U1197 (N_1197,N_915,N_469);
or U1198 (N_1198,N_984,N_625);
nor U1199 (N_1199,N_839,N_251);
or U1200 (N_1200,N_210,N_853);
xnor U1201 (N_1201,N_991,N_684);
xor U1202 (N_1202,N_207,N_309);
nand U1203 (N_1203,N_570,N_717);
or U1204 (N_1204,N_818,N_338);
nand U1205 (N_1205,N_310,N_299);
or U1206 (N_1206,N_850,N_893);
and U1207 (N_1207,N_752,N_167);
and U1208 (N_1208,N_86,N_712);
or U1209 (N_1209,N_710,N_467);
or U1210 (N_1210,N_740,N_288);
nand U1211 (N_1211,N_969,N_365);
or U1212 (N_1212,N_644,N_977);
nand U1213 (N_1213,N_209,N_138);
or U1214 (N_1214,N_540,N_100);
nand U1215 (N_1215,N_174,N_200);
and U1216 (N_1216,N_129,N_793);
nor U1217 (N_1217,N_474,N_589);
nor U1218 (N_1218,N_671,N_594);
or U1219 (N_1219,N_573,N_318);
or U1220 (N_1220,N_419,N_533);
nor U1221 (N_1221,N_351,N_316);
nor U1222 (N_1222,N_530,N_497);
or U1223 (N_1223,N_815,N_84);
xor U1224 (N_1224,N_779,N_936);
and U1225 (N_1225,N_955,N_219);
nand U1226 (N_1226,N_246,N_142);
nand U1227 (N_1227,N_90,N_260);
or U1228 (N_1228,N_172,N_911);
nor U1229 (N_1229,N_295,N_185);
xor U1230 (N_1230,N_62,N_500);
xnor U1231 (N_1231,N_403,N_290);
xnor U1232 (N_1232,N_557,N_639);
or U1233 (N_1233,N_502,N_238);
nor U1234 (N_1234,N_790,N_125);
nor U1235 (N_1235,N_523,N_937);
and U1236 (N_1236,N_655,N_799);
or U1237 (N_1237,N_885,N_809);
nor U1238 (N_1238,N_768,N_221);
xnor U1239 (N_1239,N_769,N_266);
nor U1240 (N_1240,N_976,N_283);
and U1241 (N_1241,N_800,N_269);
nand U1242 (N_1242,N_683,N_816);
nand U1243 (N_1243,N_607,N_501);
nand U1244 (N_1244,N_473,N_711);
nor U1245 (N_1245,N_822,N_327);
nor U1246 (N_1246,N_554,N_74);
nand U1247 (N_1247,N_253,N_284);
and U1248 (N_1248,N_583,N_280);
and U1249 (N_1249,N_581,N_356);
or U1250 (N_1250,N_773,N_388);
nand U1251 (N_1251,N_279,N_564);
xor U1252 (N_1252,N_965,N_567);
or U1253 (N_1253,N_490,N_297);
nor U1254 (N_1254,N_806,N_369);
nor U1255 (N_1255,N_118,N_143);
nand U1256 (N_1256,N_440,N_994);
nand U1257 (N_1257,N_182,N_8);
nand U1258 (N_1258,N_268,N_81);
or U1259 (N_1259,N_368,N_876);
nand U1260 (N_1260,N_695,N_686);
nor U1261 (N_1261,N_228,N_177);
nor U1262 (N_1262,N_51,N_293);
and U1263 (N_1263,N_613,N_405);
xor U1264 (N_1264,N_437,N_455);
nand U1265 (N_1265,N_718,N_988);
xnor U1266 (N_1266,N_421,N_733);
nand U1267 (N_1267,N_701,N_618);
nand U1268 (N_1268,N_869,N_608);
nand U1269 (N_1269,N_235,N_121);
and U1270 (N_1270,N_399,N_763);
xor U1271 (N_1271,N_186,N_713);
or U1272 (N_1272,N_631,N_334);
or U1273 (N_1273,N_215,N_997);
or U1274 (N_1274,N_213,N_985);
nor U1275 (N_1275,N_18,N_72);
nand U1276 (N_1276,N_643,N_624);
and U1277 (N_1277,N_263,N_591);
nor U1278 (N_1278,N_801,N_256);
and U1279 (N_1279,N_944,N_826);
nand U1280 (N_1280,N_975,N_376);
and U1281 (N_1281,N_472,N_664);
nor U1282 (N_1282,N_514,N_690);
or U1283 (N_1283,N_872,N_165);
or U1284 (N_1284,N_459,N_787);
xor U1285 (N_1285,N_953,N_61);
xor U1286 (N_1286,N_576,N_448);
nor U1287 (N_1287,N_250,N_606);
or U1288 (N_1288,N_352,N_193);
xnor U1289 (N_1289,N_404,N_863);
or U1290 (N_1290,N_615,N_804);
nand U1291 (N_1291,N_962,N_807);
nand U1292 (N_1292,N_9,N_336);
nand U1293 (N_1293,N_161,N_371);
nor U1294 (N_1294,N_689,N_239);
nand U1295 (N_1295,N_848,N_687);
nor U1296 (N_1296,N_909,N_275);
and U1297 (N_1297,N_494,N_300);
and U1298 (N_1298,N_389,N_311);
nor U1299 (N_1299,N_370,N_868);
and U1300 (N_1300,N_626,N_681);
or U1301 (N_1301,N_524,N_675);
or U1302 (N_1302,N_208,N_837);
nor U1303 (N_1303,N_24,N_575);
and U1304 (N_1304,N_830,N_255);
nand U1305 (N_1305,N_723,N_532);
and U1306 (N_1306,N_751,N_261);
nor U1307 (N_1307,N_582,N_308);
xnor U1308 (N_1308,N_783,N_150);
or U1309 (N_1309,N_230,N_851);
xor U1310 (N_1310,N_393,N_510);
and U1311 (N_1311,N_762,N_109);
or U1312 (N_1312,N_708,N_907);
nor U1313 (N_1313,N_64,N_940);
and U1314 (N_1314,N_513,N_366);
nand U1315 (N_1315,N_6,N_614);
nor U1316 (N_1316,N_593,N_947);
nor U1317 (N_1317,N_541,N_330);
nand U1318 (N_1318,N_748,N_425);
or U1319 (N_1319,N_550,N_896);
xnor U1320 (N_1320,N_178,N_450);
nor U1321 (N_1321,N_905,N_978);
nand U1322 (N_1322,N_702,N_889);
and U1323 (N_1323,N_949,N_647);
xor U1324 (N_1324,N_866,N_651);
nand U1325 (N_1325,N_900,N_396);
nand U1326 (N_1326,N_895,N_76);
nand U1327 (N_1327,N_312,N_94);
nor U1328 (N_1328,N_128,N_135);
or U1329 (N_1329,N_38,N_734);
and U1330 (N_1330,N_385,N_705);
nor U1331 (N_1331,N_517,N_855);
and U1332 (N_1332,N_59,N_525);
and U1333 (N_1333,N_139,N_956);
nand U1334 (N_1334,N_796,N_17);
or U1335 (N_1335,N_998,N_629);
nor U1336 (N_1336,N_758,N_355);
nand U1337 (N_1337,N_744,N_111);
nor U1338 (N_1338,N_877,N_874);
nor U1339 (N_1339,N_878,N_191);
or U1340 (N_1340,N_80,N_574);
nor U1341 (N_1341,N_479,N_794);
or U1342 (N_1342,N_699,N_785);
or U1343 (N_1343,N_457,N_107);
nor U1344 (N_1344,N_496,N_339);
nor U1345 (N_1345,N_67,N_766);
nor U1346 (N_1346,N_609,N_759);
nand U1347 (N_1347,N_852,N_963);
and U1348 (N_1348,N_387,N_476);
xor U1349 (N_1349,N_596,N_287);
and U1350 (N_1350,N_982,N_85);
and U1351 (N_1351,N_434,N_742);
and U1352 (N_1352,N_770,N_750);
nor U1353 (N_1353,N_343,N_670);
or U1354 (N_1354,N_653,N_619);
nand U1355 (N_1355,N_247,N_315);
nor U1356 (N_1356,N_611,N_652);
xor U1357 (N_1357,N_565,N_44);
or U1358 (N_1358,N_346,N_112);
nor U1359 (N_1359,N_735,N_160);
xnor U1360 (N_1360,N_841,N_360);
nor U1361 (N_1361,N_537,N_319);
nor U1362 (N_1362,N_696,N_709);
and U1363 (N_1363,N_938,N_507);
nor U1364 (N_1364,N_595,N_529);
nand U1365 (N_1365,N_903,N_492);
nor U1366 (N_1366,N_642,N_158);
or U1367 (N_1367,N_980,N_808);
or U1368 (N_1368,N_35,N_180);
or U1369 (N_1369,N_867,N_69);
or U1370 (N_1370,N_83,N_552);
nor U1371 (N_1371,N_820,N_54);
nor U1372 (N_1372,N_190,N_849);
or U1373 (N_1373,N_832,N_400);
and U1374 (N_1374,N_660,N_415);
and U1375 (N_1375,N_747,N_321);
or U1376 (N_1376,N_659,N_562);
xor U1377 (N_1377,N_685,N_489);
and U1378 (N_1378,N_184,N_568);
nand U1379 (N_1379,N_730,N_950);
or U1380 (N_1380,N_879,N_156);
xnor U1381 (N_1381,N_814,N_673);
xor U1382 (N_1382,N_697,N_677);
xor U1383 (N_1383,N_722,N_835);
and U1384 (N_1384,N_556,N_195);
nor U1385 (N_1385,N_202,N_77);
and U1386 (N_1386,N_891,N_797);
nand U1387 (N_1387,N_764,N_314);
and U1388 (N_1388,N_648,N_211);
nor U1389 (N_1389,N_505,N_223);
or U1390 (N_1390,N_282,N_60);
nand U1391 (N_1391,N_973,N_164);
nor U1392 (N_1392,N_908,N_92);
or U1393 (N_1393,N_475,N_493);
and U1394 (N_1394,N_633,N_860);
nand U1395 (N_1395,N_511,N_939);
nand U1396 (N_1396,N_345,N_347);
nor U1397 (N_1397,N_430,N_218);
or U1398 (N_1398,N_137,N_113);
and U1399 (N_1399,N_491,N_123);
nand U1400 (N_1400,N_521,N_749);
nor U1401 (N_1401,N_720,N_577);
nand U1402 (N_1402,N_945,N_398);
nor U1403 (N_1403,N_761,N_831);
nor U1404 (N_1404,N_372,N_638);
and U1405 (N_1405,N_519,N_362);
and U1406 (N_1406,N_204,N_364);
and U1407 (N_1407,N_432,N_259);
nand U1408 (N_1408,N_548,N_798);
or U1409 (N_1409,N_487,N_846);
or U1410 (N_1410,N_27,N_353);
nor U1411 (N_1411,N_296,N_63);
nand U1412 (N_1412,N_587,N_271);
and U1413 (N_1413,N_477,N_326);
and U1414 (N_1414,N_930,N_453);
and U1415 (N_1415,N_544,N_650);
or U1416 (N_1416,N_899,N_199);
or U1417 (N_1417,N_990,N_719);
nand U1418 (N_1418,N_41,N_407);
nor U1419 (N_1419,N_992,N_495);
nand U1420 (N_1420,N_130,N_590);
and U1421 (N_1421,N_229,N_446);
and U1422 (N_1422,N_834,N_286);
and U1423 (N_1423,N_760,N_43);
and U1424 (N_1424,N_252,N_668);
nor U1425 (N_1425,N_503,N_140);
nor U1426 (N_1426,N_882,N_166);
xor U1427 (N_1427,N_509,N_776);
nor U1428 (N_1428,N_96,N_37);
nand U1429 (N_1429,N_715,N_649);
or U1430 (N_1430,N_461,N_220);
or U1431 (N_1431,N_716,N_887);
or U1432 (N_1432,N_571,N_458);
nor U1433 (N_1433,N_50,N_70);
xor U1434 (N_1434,N_821,N_416);
nor U1435 (N_1435,N_274,N_960);
nand U1436 (N_1436,N_729,N_580);
and U1437 (N_1437,N_412,N_103);
xnor U1438 (N_1438,N_217,N_442);
nor U1439 (N_1439,N_703,N_201);
nor U1440 (N_1440,N_359,N_605);
or U1441 (N_1441,N_132,N_470);
and U1442 (N_1442,N_995,N_241);
or U1443 (N_1443,N_395,N_110);
nand U1444 (N_1444,N_745,N_738);
or U1445 (N_1445,N_414,N_731);
nand U1446 (N_1446,N_33,N_527);
nand U1447 (N_1447,N_104,N_39);
and U1448 (N_1448,N_357,N_291);
nor U1449 (N_1449,N_53,N_553);
nand U1450 (N_1450,N_599,N_898);
or U1451 (N_1451,N_522,N_836);
or U1452 (N_1452,N_774,N_408);
or U1453 (N_1453,N_88,N_97);
and U1454 (N_1454,N_968,N_26);
nand U1455 (N_1455,N_277,N_484);
xnor U1456 (N_1456,N_159,N_392);
nand U1457 (N_1457,N_704,N_620);
nor U1458 (N_1458,N_95,N_196);
or U1459 (N_1459,N_305,N_559);
xor U1460 (N_1460,N_884,N_888);
xnor U1461 (N_1461,N_881,N_753);
or U1462 (N_1462,N_141,N_3);
and U1463 (N_1463,N_823,N_910);
or U1464 (N_1464,N_244,N_579);
xor U1465 (N_1465,N_601,N_169);
nand U1466 (N_1466,N_222,N_45);
or U1467 (N_1467,N_153,N_301);
and U1468 (N_1468,N_433,N_996);
or U1469 (N_1469,N_781,N_47);
nand U1470 (N_1470,N_916,N_194);
xnor U1471 (N_1471,N_902,N_480);
nor U1472 (N_1472,N_661,N_136);
or U1473 (N_1473,N_772,N_468);
or U1474 (N_1474,N_471,N_788);
and U1475 (N_1475,N_536,N_726);
nor U1476 (N_1476,N_452,N_332);
nand U1477 (N_1477,N_778,N_862);
nand U1478 (N_1478,N_999,N_181);
nor U1479 (N_1479,N_40,N_337);
nor U1480 (N_1480,N_340,N_890);
xnor U1481 (N_1481,N_16,N_825);
xor U1482 (N_1482,N_819,N_49);
or U1483 (N_1483,N_307,N_829);
nand U1484 (N_1484,N_187,N_637);
nand U1485 (N_1485,N_792,N_727);
nor U1486 (N_1486,N_917,N_921);
nor U1487 (N_1487,N_931,N_349);
xor U1488 (N_1488,N_645,N_19);
and U1489 (N_1489,N_558,N_124);
nand U1490 (N_1490,N_134,N_847);
and U1491 (N_1491,N_538,N_451);
nand U1492 (N_1492,N_520,N_539);
and U1493 (N_1493,N_248,N_861);
nand U1494 (N_1494,N_258,N_674);
or U1495 (N_1495,N_382,N_335);
and U1496 (N_1496,N_224,N_344);
and U1497 (N_1497,N_48,N_688);
or U1498 (N_1498,N_133,N_378);
nand U1499 (N_1499,N_828,N_304);
or U1500 (N_1500,N_168,N_584);
and U1501 (N_1501,N_407,N_960);
nor U1502 (N_1502,N_178,N_680);
or U1503 (N_1503,N_212,N_68);
nor U1504 (N_1504,N_764,N_861);
nor U1505 (N_1505,N_752,N_400);
and U1506 (N_1506,N_938,N_68);
or U1507 (N_1507,N_609,N_815);
nor U1508 (N_1508,N_954,N_20);
nor U1509 (N_1509,N_652,N_834);
and U1510 (N_1510,N_239,N_163);
xor U1511 (N_1511,N_616,N_461);
and U1512 (N_1512,N_10,N_217);
xnor U1513 (N_1513,N_997,N_188);
nand U1514 (N_1514,N_493,N_128);
xor U1515 (N_1515,N_268,N_198);
nand U1516 (N_1516,N_312,N_528);
nor U1517 (N_1517,N_750,N_728);
and U1518 (N_1518,N_199,N_416);
nand U1519 (N_1519,N_195,N_417);
nand U1520 (N_1520,N_989,N_434);
and U1521 (N_1521,N_596,N_944);
and U1522 (N_1522,N_609,N_1);
or U1523 (N_1523,N_491,N_517);
or U1524 (N_1524,N_278,N_215);
nand U1525 (N_1525,N_110,N_939);
or U1526 (N_1526,N_940,N_378);
nand U1527 (N_1527,N_581,N_114);
xnor U1528 (N_1528,N_568,N_942);
nor U1529 (N_1529,N_366,N_655);
and U1530 (N_1530,N_95,N_92);
or U1531 (N_1531,N_207,N_475);
xor U1532 (N_1532,N_181,N_631);
and U1533 (N_1533,N_30,N_11);
and U1534 (N_1534,N_980,N_968);
xor U1535 (N_1535,N_780,N_31);
nor U1536 (N_1536,N_601,N_333);
nand U1537 (N_1537,N_515,N_977);
nand U1538 (N_1538,N_876,N_885);
or U1539 (N_1539,N_101,N_802);
and U1540 (N_1540,N_577,N_44);
nor U1541 (N_1541,N_566,N_923);
and U1542 (N_1542,N_70,N_429);
xor U1543 (N_1543,N_530,N_619);
nand U1544 (N_1544,N_764,N_311);
or U1545 (N_1545,N_265,N_845);
or U1546 (N_1546,N_798,N_746);
and U1547 (N_1547,N_108,N_681);
nand U1548 (N_1548,N_935,N_622);
nand U1549 (N_1549,N_958,N_159);
nand U1550 (N_1550,N_74,N_446);
nand U1551 (N_1551,N_833,N_157);
or U1552 (N_1552,N_711,N_747);
nor U1553 (N_1553,N_558,N_117);
and U1554 (N_1554,N_263,N_130);
nor U1555 (N_1555,N_216,N_525);
or U1556 (N_1556,N_469,N_756);
xnor U1557 (N_1557,N_37,N_65);
nor U1558 (N_1558,N_367,N_45);
or U1559 (N_1559,N_213,N_266);
xnor U1560 (N_1560,N_546,N_340);
nand U1561 (N_1561,N_69,N_795);
nor U1562 (N_1562,N_91,N_944);
and U1563 (N_1563,N_348,N_338);
or U1564 (N_1564,N_992,N_36);
or U1565 (N_1565,N_176,N_754);
xor U1566 (N_1566,N_634,N_268);
nor U1567 (N_1567,N_974,N_531);
and U1568 (N_1568,N_421,N_996);
nor U1569 (N_1569,N_496,N_699);
nor U1570 (N_1570,N_325,N_961);
nor U1571 (N_1571,N_616,N_463);
and U1572 (N_1572,N_841,N_749);
and U1573 (N_1573,N_242,N_291);
nand U1574 (N_1574,N_896,N_202);
nor U1575 (N_1575,N_416,N_478);
nand U1576 (N_1576,N_735,N_156);
nor U1577 (N_1577,N_943,N_519);
nor U1578 (N_1578,N_938,N_928);
nor U1579 (N_1579,N_634,N_810);
xor U1580 (N_1580,N_675,N_877);
and U1581 (N_1581,N_588,N_895);
or U1582 (N_1582,N_761,N_251);
nor U1583 (N_1583,N_988,N_302);
nor U1584 (N_1584,N_992,N_83);
nor U1585 (N_1585,N_271,N_499);
nand U1586 (N_1586,N_175,N_928);
nand U1587 (N_1587,N_402,N_526);
or U1588 (N_1588,N_250,N_85);
or U1589 (N_1589,N_674,N_52);
or U1590 (N_1590,N_808,N_466);
and U1591 (N_1591,N_38,N_258);
nand U1592 (N_1592,N_851,N_644);
and U1593 (N_1593,N_420,N_951);
or U1594 (N_1594,N_408,N_891);
and U1595 (N_1595,N_902,N_386);
nand U1596 (N_1596,N_706,N_57);
nor U1597 (N_1597,N_429,N_845);
nor U1598 (N_1598,N_556,N_105);
or U1599 (N_1599,N_416,N_75);
nand U1600 (N_1600,N_7,N_494);
or U1601 (N_1601,N_80,N_684);
xor U1602 (N_1602,N_117,N_646);
nand U1603 (N_1603,N_79,N_9);
and U1604 (N_1604,N_905,N_854);
and U1605 (N_1605,N_82,N_474);
nand U1606 (N_1606,N_791,N_417);
or U1607 (N_1607,N_305,N_933);
or U1608 (N_1608,N_700,N_993);
xnor U1609 (N_1609,N_94,N_52);
nor U1610 (N_1610,N_65,N_600);
nand U1611 (N_1611,N_272,N_178);
nor U1612 (N_1612,N_203,N_927);
or U1613 (N_1613,N_399,N_382);
xnor U1614 (N_1614,N_439,N_351);
nand U1615 (N_1615,N_89,N_31);
or U1616 (N_1616,N_483,N_839);
or U1617 (N_1617,N_794,N_795);
or U1618 (N_1618,N_222,N_199);
or U1619 (N_1619,N_929,N_481);
nor U1620 (N_1620,N_52,N_18);
or U1621 (N_1621,N_159,N_938);
and U1622 (N_1622,N_281,N_375);
nor U1623 (N_1623,N_280,N_149);
xnor U1624 (N_1624,N_404,N_247);
nor U1625 (N_1625,N_659,N_773);
or U1626 (N_1626,N_946,N_268);
or U1627 (N_1627,N_373,N_428);
nand U1628 (N_1628,N_953,N_874);
nor U1629 (N_1629,N_791,N_132);
and U1630 (N_1630,N_187,N_35);
nand U1631 (N_1631,N_496,N_656);
nor U1632 (N_1632,N_649,N_84);
nor U1633 (N_1633,N_117,N_632);
or U1634 (N_1634,N_769,N_142);
nor U1635 (N_1635,N_851,N_983);
nand U1636 (N_1636,N_45,N_190);
or U1637 (N_1637,N_146,N_100);
xor U1638 (N_1638,N_633,N_497);
xnor U1639 (N_1639,N_657,N_951);
nor U1640 (N_1640,N_558,N_92);
nor U1641 (N_1641,N_230,N_911);
or U1642 (N_1642,N_355,N_551);
or U1643 (N_1643,N_374,N_491);
nand U1644 (N_1644,N_966,N_211);
nor U1645 (N_1645,N_928,N_687);
nor U1646 (N_1646,N_478,N_856);
and U1647 (N_1647,N_470,N_661);
and U1648 (N_1648,N_515,N_942);
and U1649 (N_1649,N_621,N_525);
and U1650 (N_1650,N_473,N_893);
nand U1651 (N_1651,N_233,N_71);
nor U1652 (N_1652,N_859,N_622);
and U1653 (N_1653,N_892,N_474);
xnor U1654 (N_1654,N_754,N_924);
or U1655 (N_1655,N_241,N_6);
xnor U1656 (N_1656,N_254,N_588);
nand U1657 (N_1657,N_797,N_982);
nand U1658 (N_1658,N_728,N_273);
or U1659 (N_1659,N_539,N_671);
and U1660 (N_1660,N_980,N_653);
nor U1661 (N_1661,N_504,N_870);
nor U1662 (N_1662,N_516,N_476);
nor U1663 (N_1663,N_89,N_429);
or U1664 (N_1664,N_100,N_520);
nand U1665 (N_1665,N_709,N_760);
xor U1666 (N_1666,N_572,N_607);
nor U1667 (N_1667,N_752,N_563);
or U1668 (N_1668,N_264,N_443);
or U1669 (N_1669,N_674,N_201);
nand U1670 (N_1670,N_546,N_873);
or U1671 (N_1671,N_78,N_834);
or U1672 (N_1672,N_725,N_587);
nand U1673 (N_1673,N_592,N_440);
nor U1674 (N_1674,N_975,N_377);
nand U1675 (N_1675,N_210,N_713);
nor U1676 (N_1676,N_582,N_449);
nor U1677 (N_1677,N_849,N_561);
or U1678 (N_1678,N_809,N_163);
and U1679 (N_1679,N_386,N_249);
and U1680 (N_1680,N_348,N_17);
and U1681 (N_1681,N_295,N_262);
nand U1682 (N_1682,N_530,N_924);
xor U1683 (N_1683,N_302,N_272);
nor U1684 (N_1684,N_290,N_234);
nand U1685 (N_1685,N_819,N_439);
and U1686 (N_1686,N_563,N_618);
or U1687 (N_1687,N_276,N_714);
nor U1688 (N_1688,N_14,N_135);
and U1689 (N_1689,N_616,N_97);
nor U1690 (N_1690,N_131,N_282);
nor U1691 (N_1691,N_531,N_249);
nor U1692 (N_1692,N_630,N_196);
xnor U1693 (N_1693,N_128,N_775);
and U1694 (N_1694,N_772,N_370);
or U1695 (N_1695,N_253,N_166);
or U1696 (N_1696,N_989,N_277);
and U1697 (N_1697,N_696,N_784);
and U1698 (N_1698,N_552,N_902);
nor U1699 (N_1699,N_301,N_539);
or U1700 (N_1700,N_420,N_418);
and U1701 (N_1701,N_749,N_183);
nor U1702 (N_1702,N_489,N_790);
nor U1703 (N_1703,N_51,N_234);
xnor U1704 (N_1704,N_16,N_508);
or U1705 (N_1705,N_992,N_553);
nor U1706 (N_1706,N_204,N_303);
nand U1707 (N_1707,N_928,N_720);
or U1708 (N_1708,N_388,N_710);
nand U1709 (N_1709,N_194,N_166);
xor U1710 (N_1710,N_304,N_189);
and U1711 (N_1711,N_717,N_563);
nor U1712 (N_1712,N_133,N_814);
and U1713 (N_1713,N_151,N_777);
xor U1714 (N_1714,N_740,N_494);
and U1715 (N_1715,N_950,N_439);
nand U1716 (N_1716,N_688,N_917);
or U1717 (N_1717,N_624,N_564);
nand U1718 (N_1718,N_840,N_314);
or U1719 (N_1719,N_257,N_145);
nor U1720 (N_1720,N_329,N_689);
nor U1721 (N_1721,N_930,N_722);
nand U1722 (N_1722,N_690,N_151);
nor U1723 (N_1723,N_71,N_273);
or U1724 (N_1724,N_701,N_291);
nor U1725 (N_1725,N_46,N_791);
or U1726 (N_1726,N_449,N_279);
or U1727 (N_1727,N_755,N_576);
xnor U1728 (N_1728,N_425,N_667);
nor U1729 (N_1729,N_197,N_277);
and U1730 (N_1730,N_755,N_84);
nand U1731 (N_1731,N_905,N_48);
and U1732 (N_1732,N_818,N_611);
nand U1733 (N_1733,N_285,N_174);
and U1734 (N_1734,N_303,N_763);
or U1735 (N_1735,N_567,N_735);
and U1736 (N_1736,N_91,N_807);
nor U1737 (N_1737,N_881,N_599);
xor U1738 (N_1738,N_364,N_776);
nand U1739 (N_1739,N_946,N_363);
nor U1740 (N_1740,N_717,N_549);
or U1741 (N_1741,N_568,N_961);
or U1742 (N_1742,N_998,N_909);
nand U1743 (N_1743,N_601,N_451);
and U1744 (N_1744,N_939,N_990);
xor U1745 (N_1745,N_467,N_699);
or U1746 (N_1746,N_8,N_966);
nand U1747 (N_1747,N_547,N_651);
nor U1748 (N_1748,N_970,N_424);
nand U1749 (N_1749,N_368,N_652);
xor U1750 (N_1750,N_966,N_946);
nor U1751 (N_1751,N_726,N_809);
and U1752 (N_1752,N_803,N_787);
xnor U1753 (N_1753,N_181,N_435);
nand U1754 (N_1754,N_46,N_106);
or U1755 (N_1755,N_600,N_681);
nor U1756 (N_1756,N_85,N_496);
and U1757 (N_1757,N_302,N_428);
nand U1758 (N_1758,N_154,N_714);
and U1759 (N_1759,N_228,N_492);
and U1760 (N_1760,N_900,N_313);
or U1761 (N_1761,N_661,N_998);
nand U1762 (N_1762,N_257,N_900);
or U1763 (N_1763,N_941,N_47);
xor U1764 (N_1764,N_953,N_48);
xor U1765 (N_1765,N_404,N_107);
and U1766 (N_1766,N_185,N_778);
nand U1767 (N_1767,N_93,N_607);
nand U1768 (N_1768,N_282,N_329);
nor U1769 (N_1769,N_186,N_855);
nand U1770 (N_1770,N_403,N_707);
nand U1771 (N_1771,N_376,N_311);
nand U1772 (N_1772,N_665,N_765);
or U1773 (N_1773,N_38,N_709);
nand U1774 (N_1774,N_671,N_232);
nand U1775 (N_1775,N_301,N_38);
xor U1776 (N_1776,N_958,N_818);
nor U1777 (N_1777,N_475,N_771);
or U1778 (N_1778,N_232,N_94);
nand U1779 (N_1779,N_159,N_77);
and U1780 (N_1780,N_671,N_66);
xnor U1781 (N_1781,N_210,N_470);
and U1782 (N_1782,N_498,N_189);
nand U1783 (N_1783,N_932,N_841);
and U1784 (N_1784,N_902,N_591);
nor U1785 (N_1785,N_774,N_354);
or U1786 (N_1786,N_401,N_83);
nor U1787 (N_1787,N_617,N_569);
nand U1788 (N_1788,N_301,N_265);
nor U1789 (N_1789,N_342,N_241);
or U1790 (N_1790,N_967,N_164);
nand U1791 (N_1791,N_400,N_557);
xnor U1792 (N_1792,N_424,N_728);
nor U1793 (N_1793,N_719,N_478);
and U1794 (N_1794,N_812,N_35);
nand U1795 (N_1795,N_996,N_422);
xor U1796 (N_1796,N_49,N_617);
or U1797 (N_1797,N_164,N_920);
and U1798 (N_1798,N_895,N_981);
nor U1799 (N_1799,N_238,N_870);
nand U1800 (N_1800,N_157,N_491);
and U1801 (N_1801,N_758,N_859);
nand U1802 (N_1802,N_119,N_200);
or U1803 (N_1803,N_829,N_459);
or U1804 (N_1804,N_708,N_798);
nor U1805 (N_1805,N_141,N_652);
and U1806 (N_1806,N_228,N_77);
nand U1807 (N_1807,N_232,N_630);
and U1808 (N_1808,N_614,N_572);
nand U1809 (N_1809,N_168,N_886);
or U1810 (N_1810,N_254,N_120);
nand U1811 (N_1811,N_631,N_962);
nand U1812 (N_1812,N_842,N_68);
xor U1813 (N_1813,N_103,N_600);
nor U1814 (N_1814,N_626,N_988);
or U1815 (N_1815,N_730,N_269);
nor U1816 (N_1816,N_746,N_705);
and U1817 (N_1817,N_925,N_379);
nand U1818 (N_1818,N_44,N_664);
and U1819 (N_1819,N_957,N_548);
nor U1820 (N_1820,N_595,N_881);
nor U1821 (N_1821,N_448,N_939);
xnor U1822 (N_1822,N_486,N_622);
and U1823 (N_1823,N_713,N_526);
nand U1824 (N_1824,N_185,N_896);
nor U1825 (N_1825,N_580,N_172);
or U1826 (N_1826,N_962,N_997);
nor U1827 (N_1827,N_85,N_535);
or U1828 (N_1828,N_36,N_398);
nand U1829 (N_1829,N_836,N_362);
or U1830 (N_1830,N_219,N_65);
xnor U1831 (N_1831,N_865,N_146);
nor U1832 (N_1832,N_453,N_132);
xnor U1833 (N_1833,N_751,N_181);
or U1834 (N_1834,N_182,N_799);
nand U1835 (N_1835,N_525,N_673);
or U1836 (N_1836,N_952,N_211);
nand U1837 (N_1837,N_516,N_705);
xor U1838 (N_1838,N_3,N_51);
nor U1839 (N_1839,N_128,N_350);
nand U1840 (N_1840,N_118,N_932);
nor U1841 (N_1841,N_557,N_889);
nand U1842 (N_1842,N_612,N_541);
and U1843 (N_1843,N_251,N_495);
nand U1844 (N_1844,N_105,N_805);
nand U1845 (N_1845,N_40,N_836);
nor U1846 (N_1846,N_129,N_700);
and U1847 (N_1847,N_71,N_208);
nor U1848 (N_1848,N_277,N_154);
nand U1849 (N_1849,N_905,N_756);
xor U1850 (N_1850,N_615,N_824);
and U1851 (N_1851,N_529,N_143);
nand U1852 (N_1852,N_335,N_256);
nor U1853 (N_1853,N_452,N_621);
and U1854 (N_1854,N_6,N_761);
nor U1855 (N_1855,N_552,N_422);
or U1856 (N_1856,N_947,N_9);
xor U1857 (N_1857,N_364,N_8);
nand U1858 (N_1858,N_151,N_935);
xor U1859 (N_1859,N_464,N_586);
nor U1860 (N_1860,N_555,N_944);
nand U1861 (N_1861,N_882,N_662);
and U1862 (N_1862,N_131,N_170);
nand U1863 (N_1863,N_173,N_111);
xor U1864 (N_1864,N_80,N_223);
or U1865 (N_1865,N_665,N_674);
nor U1866 (N_1866,N_848,N_557);
and U1867 (N_1867,N_721,N_669);
or U1868 (N_1868,N_436,N_516);
xnor U1869 (N_1869,N_454,N_668);
nor U1870 (N_1870,N_903,N_36);
nor U1871 (N_1871,N_489,N_896);
nand U1872 (N_1872,N_447,N_721);
nor U1873 (N_1873,N_964,N_133);
nand U1874 (N_1874,N_153,N_936);
nand U1875 (N_1875,N_210,N_564);
xor U1876 (N_1876,N_168,N_705);
and U1877 (N_1877,N_66,N_859);
and U1878 (N_1878,N_86,N_967);
or U1879 (N_1879,N_174,N_602);
nor U1880 (N_1880,N_255,N_883);
nor U1881 (N_1881,N_4,N_721);
nor U1882 (N_1882,N_758,N_777);
or U1883 (N_1883,N_582,N_51);
and U1884 (N_1884,N_808,N_553);
or U1885 (N_1885,N_357,N_472);
nor U1886 (N_1886,N_900,N_827);
nand U1887 (N_1887,N_866,N_595);
xnor U1888 (N_1888,N_871,N_766);
xnor U1889 (N_1889,N_653,N_311);
nor U1890 (N_1890,N_550,N_439);
xor U1891 (N_1891,N_621,N_796);
and U1892 (N_1892,N_264,N_464);
or U1893 (N_1893,N_912,N_867);
nand U1894 (N_1894,N_426,N_388);
or U1895 (N_1895,N_645,N_370);
nand U1896 (N_1896,N_784,N_31);
nor U1897 (N_1897,N_894,N_812);
nor U1898 (N_1898,N_848,N_404);
nand U1899 (N_1899,N_572,N_168);
nor U1900 (N_1900,N_369,N_326);
nand U1901 (N_1901,N_721,N_277);
and U1902 (N_1902,N_741,N_774);
or U1903 (N_1903,N_574,N_454);
and U1904 (N_1904,N_296,N_622);
or U1905 (N_1905,N_376,N_260);
and U1906 (N_1906,N_753,N_671);
xnor U1907 (N_1907,N_10,N_164);
or U1908 (N_1908,N_652,N_412);
and U1909 (N_1909,N_352,N_685);
xor U1910 (N_1910,N_686,N_449);
and U1911 (N_1911,N_333,N_835);
xor U1912 (N_1912,N_69,N_812);
and U1913 (N_1913,N_597,N_807);
or U1914 (N_1914,N_397,N_2);
nor U1915 (N_1915,N_602,N_34);
nor U1916 (N_1916,N_646,N_916);
and U1917 (N_1917,N_333,N_742);
and U1918 (N_1918,N_533,N_107);
and U1919 (N_1919,N_8,N_979);
or U1920 (N_1920,N_626,N_396);
nor U1921 (N_1921,N_405,N_521);
or U1922 (N_1922,N_787,N_24);
nor U1923 (N_1923,N_762,N_95);
nand U1924 (N_1924,N_862,N_782);
nand U1925 (N_1925,N_333,N_687);
nor U1926 (N_1926,N_918,N_721);
and U1927 (N_1927,N_587,N_866);
nor U1928 (N_1928,N_1,N_416);
nor U1929 (N_1929,N_769,N_196);
nor U1930 (N_1930,N_660,N_759);
nor U1931 (N_1931,N_698,N_256);
and U1932 (N_1932,N_24,N_889);
and U1933 (N_1933,N_2,N_465);
and U1934 (N_1934,N_948,N_852);
nor U1935 (N_1935,N_34,N_228);
nor U1936 (N_1936,N_91,N_317);
or U1937 (N_1937,N_257,N_922);
or U1938 (N_1938,N_806,N_778);
and U1939 (N_1939,N_747,N_272);
xor U1940 (N_1940,N_530,N_317);
nor U1941 (N_1941,N_774,N_650);
nor U1942 (N_1942,N_671,N_700);
or U1943 (N_1943,N_952,N_706);
nor U1944 (N_1944,N_544,N_40);
nand U1945 (N_1945,N_33,N_255);
xnor U1946 (N_1946,N_179,N_614);
or U1947 (N_1947,N_309,N_938);
and U1948 (N_1948,N_926,N_409);
nand U1949 (N_1949,N_483,N_442);
or U1950 (N_1950,N_839,N_322);
or U1951 (N_1951,N_712,N_450);
nand U1952 (N_1952,N_833,N_151);
and U1953 (N_1953,N_994,N_755);
xnor U1954 (N_1954,N_521,N_825);
and U1955 (N_1955,N_754,N_3);
or U1956 (N_1956,N_253,N_66);
and U1957 (N_1957,N_228,N_290);
nand U1958 (N_1958,N_612,N_518);
and U1959 (N_1959,N_58,N_230);
or U1960 (N_1960,N_518,N_105);
nor U1961 (N_1961,N_30,N_983);
nor U1962 (N_1962,N_529,N_954);
nand U1963 (N_1963,N_654,N_239);
nor U1964 (N_1964,N_675,N_621);
nand U1965 (N_1965,N_257,N_766);
and U1966 (N_1966,N_702,N_404);
nor U1967 (N_1967,N_602,N_954);
nor U1968 (N_1968,N_856,N_69);
nand U1969 (N_1969,N_192,N_404);
nor U1970 (N_1970,N_386,N_732);
nor U1971 (N_1971,N_990,N_546);
nand U1972 (N_1972,N_265,N_680);
nor U1973 (N_1973,N_745,N_948);
nand U1974 (N_1974,N_285,N_372);
and U1975 (N_1975,N_866,N_50);
or U1976 (N_1976,N_724,N_708);
nor U1977 (N_1977,N_2,N_930);
or U1978 (N_1978,N_148,N_454);
xnor U1979 (N_1979,N_467,N_256);
nand U1980 (N_1980,N_184,N_914);
nand U1981 (N_1981,N_634,N_937);
or U1982 (N_1982,N_315,N_150);
or U1983 (N_1983,N_514,N_560);
and U1984 (N_1984,N_205,N_740);
nor U1985 (N_1985,N_302,N_98);
and U1986 (N_1986,N_355,N_258);
nand U1987 (N_1987,N_165,N_484);
and U1988 (N_1988,N_418,N_415);
nand U1989 (N_1989,N_846,N_935);
nand U1990 (N_1990,N_153,N_232);
and U1991 (N_1991,N_546,N_850);
nor U1992 (N_1992,N_506,N_539);
and U1993 (N_1993,N_34,N_286);
xnor U1994 (N_1994,N_688,N_344);
nor U1995 (N_1995,N_491,N_386);
and U1996 (N_1996,N_105,N_372);
and U1997 (N_1997,N_120,N_145);
nand U1998 (N_1998,N_106,N_14);
or U1999 (N_1999,N_471,N_230);
xnor U2000 (N_2000,N_1776,N_1475);
or U2001 (N_2001,N_1889,N_1841);
nand U2002 (N_2002,N_1975,N_1223);
nor U2003 (N_2003,N_1898,N_1431);
or U2004 (N_2004,N_1266,N_1699);
and U2005 (N_2005,N_1255,N_1429);
nand U2006 (N_2006,N_1456,N_1376);
nand U2007 (N_2007,N_1234,N_1936);
and U2008 (N_2008,N_1476,N_1779);
nor U2009 (N_2009,N_1031,N_1311);
and U2010 (N_2010,N_1291,N_1228);
nand U2011 (N_2011,N_1704,N_1408);
and U2012 (N_2012,N_1585,N_1319);
or U2013 (N_2013,N_1063,N_1661);
nand U2014 (N_2014,N_1143,N_1347);
nor U2015 (N_2015,N_1672,N_1034);
or U2016 (N_2016,N_1486,N_1589);
and U2017 (N_2017,N_1999,N_1618);
or U2018 (N_2018,N_1494,N_1281);
nor U2019 (N_2019,N_1225,N_1395);
and U2020 (N_2020,N_1771,N_1335);
and U2021 (N_2021,N_1501,N_1949);
and U2022 (N_2022,N_1533,N_1306);
nand U2023 (N_2023,N_1108,N_1194);
and U2024 (N_2024,N_1753,N_1890);
and U2025 (N_2025,N_1263,N_1768);
and U2026 (N_2026,N_1605,N_1010);
or U2027 (N_2027,N_1328,N_1440);
nand U2028 (N_2028,N_1430,N_1750);
nand U2029 (N_2029,N_1612,N_1561);
or U2030 (N_2030,N_1356,N_1535);
and U2031 (N_2031,N_1229,N_1198);
and U2032 (N_2032,N_1235,N_1277);
nand U2033 (N_2033,N_1979,N_1098);
and U2034 (N_2034,N_1379,N_1652);
nor U2035 (N_2035,N_1287,N_1482);
nand U2036 (N_2036,N_1237,N_1847);
and U2037 (N_2037,N_1368,N_1427);
nor U2038 (N_2038,N_1338,N_1327);
and U2039 (N_2039,N_1591,N_1109);
and U2040 (N_2040,N_1659,N_1913);
or U2041 (N_2041,N_1906,N_1880);
nor U2042 (N_2042,N_1901,N_1732);
and U2043 (N_2043,N_1537,N_1226);
nor U2044 (N_2044,N_1514,N_1353);
and U2045 (N_2045,N_1869,N_1744);
nor U2046 (N_2046,N_1997,N_1496);
or U2047 (N_2047,N_1657,N_1918);
nand U2048 (N_2048,N_1624,N_1608);
and U2049 (N_2049,N_1726,N_1660);
nand U2050 (N_2050,N_1003,N_1286);
xor U2051 (N_2051,N_1354,N_1176);
nand U2052 (N_2052,N_1013,N_1484);
or U2053 (N_2053,N_1682,N_1819);
nand U2054 (N_2054,N_1487,N_1520);
nor U2055 (N_2055,N_1619,N_1643);
and U2056 (N_2056,N_1043,N_1828);
nor U2057 (N_2057,N_1763,N_1530);
and U2058 (N_2058,N_1444,N_1056);
nand U2059 (N_2059,N_1911,N_1305);
nor U2060 (N_2060,N_1665,N_1500);
nor U2061 (N_2061,N_1859,N_1713);
and U2062 (N_2062,N_1360,N_1565);
xor U2063 (N_2063,N_1217,N_1320);
nor U2064 (N_2064,N_1441,N_1212);
nand U2065 (N_2065,N_1468,N_1173);
or U2066 (N_2066,N_1460,N_1697);
or U2067 (N_2067,N_1649,N_1593);
nand U2068 (N_2068,N_1271,N_1739);
nor U2069 (N_2069,N_1413,N_1493);
and U2070 (N_2070,N_1445,N_1887);
xnor U2071 (N_2071,N_1821,N_1769);
nor U2072 (N_2072,N_1128,N_1965);
and U2073 (N_2073,N_1510,N_1443);
xor U2074 (N_2074,N_1791,N_1982);
nor U2075 (N_2075,N_1762,N_1012);
nor U2076 (N_2076,N_1703,N_1380);
and U2077 (N_2077,N_1384,N_1323);
and U2078 (N_2078,N_1386,N_1688);
or U2079 (N_2079,N_1896,N_1946);
nor U2080 (N_2080,N_1206,N_1939);
nand U2081 (N_2081,N_1680,N_1049);
and U2082 (N_2082,N_1187,N_1943);
nand U2083 (N_2083,N_1477,N_1086);
xnor U2084 (N_2084,N_1976,N_1213);
and U2085 (N_2085,N_1352,N_1015);
or U2086 (N_2086,N_1282,N_1199);
or U2087 (N_2087,N_1696,N_1724);
or U2088 (N_2088,N_1546,N_1935);
nor U2089 (N_2089,N_1813,N_1960);
nor U2090 (N_2090,N_1170,N_1362);
or U2091 (N_2091,N_1833,N_1942);
or U2092 (N_2092,N_1417,N_1528);
nand U2093 (N_2093,N_1645,N_1937);
xnor U2094 (N_2094,N_1861,N_1256);
or U2095 (N_2095,N_1160,N_1967);
nor U2096 (N_2096,N_1106,N_1866);
nand U2097 (N_2097,N_1785,N_1519);
nor U2098 (N_2098,N_1595,N_1656);
nor U2099 (N_2099,N_1601,N_1978);
nor U2100 (N_2100,N_1089,N_1558);
or U2101 (N_2101,N_1590,N_1433);
and U2102 (N_2102,N_1518,N_1425);
or U2103 (N_2103,N_1919,N_1893);
nor U2104 (N_2104,N_1471,N_1100);
xnor U2105 (N_2105,N_1342,N_1285);
and U2106 (N_2106,N_1868,N_1243);
or U2107 (N_2107,N_1647,N_1358);
nor U2108 (N_2108,N_1584,N_1127);
and U2109 (N_2109,N_1250,N_1723);
and U2110 (N_2110,N_1721,N_1559);
xor U2111 (N_2111,N_1862,N_1473);
nand U2112 (N_2112,N_1130,N_1382);
or U2113 (N_2113,N_1451,N_1857);
xor U2114 (N_2114,N_1592,N_1599);
xor U2115 (N_2115,N_1567,N_1046);
or U2116 (N_2116,N_1693,N_1808);
or U2117 (N_2117,N_1834,N_1236);
nand U2118 (N_2118,N_1815,N_1525);
nand U2119 (N_2119,N_1941,N_1845);
nand U2120 (N_2120,N_1884,N_1416);
or U2121 (N_2121,N_1509,N_1930);
nor U2122 (N_2122,N_1956,N_1921);
nand U2123 (N_2123,N_1094,N_1747);
or U2124 (N_2124,N_1614,N_1016);
or U2125 (N_2125,N_1773,N_1414);
nor U2126 (N_2126,N_1905,N_1071);
or U2127 (N_2127,N_1527,N_1515);
nand U2128 (N_2128,N_1298,N_1505);
or U2129 (N_2129,N_1393,N_1695);
nor U2130 (N_2130,N_1961,N_1453);
or U2131 (N_2131,N_1208,N_1994);
nand U2132 (N_2132,N_1800,N_1827);
or U2133 (N_2133,N_1992,N_1093);
or U2134 (N_2134,N_1728,N_1372);
and U2135 (N_2135,N_1251,N_1267);
or U2136 (N_2136,N_1481,N_1265);
nand U2137 (N_2137,N_1120,N_1953);
nor U2138 (N_2138,N_1774,N_1420);
nand U2139 (N_2139,N_1014,N_1539);
or U2140 (N_2140,N_1066,N_1080);
or U2141 (N_2141,N_1302,N_1111);
nor U2142 (N_2142,N_1415,N_1041);
nor U2143 (N_2143,N_1172,N_1099);
or U2144 (N_2144,N_1268,N_1474);
xnor U2145 (N_2145,N_1787,N_1945);
nor U2146 (N_2146,N_1081,N_1597);
nor U2147 (N_2147,N_1050,N_1995);
or U2148 (N_2148,N_1465,N_1262);
and U2149 (N_2149,N_1606,N_1466);
nand U2150 (N_2150,N_1694,N_1947);
xnor U2151 (N_2151,N_1784,N_1439);
nand U2152 (N_2152,N_1708,N_1264);
xor U2153 (N_2153,N_1838,N_1725);
xor U2154 (N_2154,N_1547,N_1908);
xor U2155 (N_2155,N_1087,N_1853);
nand U2156 (N_2156,N_1782,N_1394);
xor U2157 (N_2157,N_1240,N_1326);
nor U2158 (N_2158,N_1200,N_1712);
nand U2159 (N_2159,N_1163,N_1238);
nor U2160 (N_2160,N_1793,N_1432);
and U2161 (N_2161,N_1736,N_1634);
nand U2162 (N_2162,N_1818,N_1761);
nor U2163 (N_2163,N_1863,N_1367);
nand U2164 (N_2164,N_1702,N_1400);
nor U2165 (N_2165,N_1646,N_1715);
xor U2166 (N_2166,N_1042,N_1166);
xor U2167 (N_2167,N_1344,N_1783);
nand U2168 (N_2168,N_1454,N_1058);
nor U2169 (N_2169,N_1290,N_1575);
and U2170 (N_2170,N_1572,N_1650);
nor U2171 (N_2171,N_1403,N_1141);
nor U2172 (N_2172,N_1824,N_1716);
nand U2173 (N_2173,N_1180,N_1745);
nor U2174 (N_2174,N_1900,N_1125);
and U2175 (N_2175,N_1743,N_1934);
nor U2176 (N_2176,N_1741,N_1681);
or U2177 (N_2177,N_1436,N_1830);
and U2178 (N_2178,N_1147,N_1698);
and U2179 (N_2179,N_1090,N_1801);
nand U2180 (N_2180,N_1405,N_1553);
or U2181 (N_2181,N_1877,N_1249);
and U2182 (N_2182,N_1545,N_1511);
and U2183 (N_2183,N_1580,N_1447);
xnor U2184 (N_2184,N_1331,N_1182);
or U2185 (N_2185,N_1790,N_1806);
nand U2186 (N_2186,N_1038,N_1574);
or U2187 (N_2187,N_1304,N_1966);
nand U2188 (N_2188,N_1734,N_1951);
nand U2189 (N_2189,N_1024,N_1222);
or U2190 (N_2190,N_1563,N_1067);
and U2191 (N_2191,N_1419,N_1987);
nand U2192 (N_2192,N_1759,N_1873);
nand U2193 (N_2193,N_1437,N_1462);
or U2194 (N_2194,N_1507,N_1219);
nand U2195 (N_2195,N_1107,N_1516);
xnor U2196 (N_2196,N_1810,N_1274);
nor U2197 (N_2197,N_1028,N_1065);
nand U2198 (N_2198,N_1571,N_1259);
nor U2199 (N_2199,N_1749,N_1714);
nor U2200 (N_2200,N_1668,N_1635);
xor U2201 (N_2201,N_1371,N_1438);
nand U2202 (N_2202,N_1917,N_1835);
and U2203 (N_2203,N_1142,N_1005);
or U2204 (N_2204,N_1927,N_1188);
or U2205 (N_2205,N_1727,N_1875);
xor U2206 (N_2206,N_1020,N_1114);
and U2207 (N_2207,N_1879,N_1766);
nand U2208 (N_2208,N_1381,N_1296);
nand U2209 (N_2209,N_1689,N_1678);
and U2210 (N_2210,N_1581,N_1280);
nor U2211 (N_2211,N_1955,N_1018);
nor U2212 (N_2212,N_1637,N_1512);
and U2213 (N_2213,N_1310,N_1370);
and U2214 (N_2214,N_1276,N_1241);
nor U2215 (N_2215,N_1137,N_1675);
or U2216 (N_2216,N_1498,N_1991);
or U2217 (N_2217,N_1390,N_1532);
or U2218 (N_2218,N_1330,N_1174);
nor U2219 (N_2219,N_1555,N_1490);
nor U2220 (N_2220,N_1780,N_1004);
and U2221 (N_2221,N_1588,N_1369);
nand U2222 (N_2222,N_1168,N_1710);
and U2223 (N_2223,N_1644,N_1165);
and U2224 (N_2224,N_1191,N_1933);
nand U2225 (N_2225,N_1129,N_1722);
nand U2226 (N_2226,N_1136,N_1464);
nand U2227 (N_2227,N_1816,N_1077);
nor U2228 (N_2228,N_1506,N_1061);
nor U2229 (N_2229,N_1551,N_1526);
nand U2230 (N_2230,N_1151,N_1928);
and U2231 (N_2231,N_1653,N_1074);
nand U2232 (N_2232,N_1556,N_1626);
nor U2233 (N_2233,N_1088,N_1118);
nand U2234 (N_2234,N_1974,N_1085);
and U2235 (N_2235,N_1765,N_1795);
or U2236 (N_2236,N_1993,N_1489);
or U2237 (N_2237,N_1201,N_1169);
and U2238 (N_2238,N_1383,N_1117);
nand U2239 (N_2239,N_1092,N_1711);
nand U2240 (N_2240,N_1984,N_1822);
and U2241 (N_2241,N_1959,N_1124);
and U2242 (N_2242,N_1632,N_1638);
nor U2243 (N_2243,N_1073,N_1220);
nand U2244 (N_2244,N_1452,N_1521);
and U2245 (N_2245,N_1598,N_1258);
or U2246 (N_2246,N_1625,N_1864);
and U2247 (N_2247,N_1811,N_1078);
and U2248 (N_2248,N_1449,N_1876);
nand U2249 (N_2249,N_1871,N_1664);
and U2250 (N_2250,N_1197,N_1190);
or U2251 (N_2251,N_1303,N_1971);
xnor U2252 (N_2252,N_1562,N_1154);
and U2253 (N_2253,N_1651,N_1836);
and U2254 (N_2254,N_1629,N_1275);
or U2255 (N_2255,N_1435,N_1973);
and U2256 (N_2256,N_1273,N_1426);
or U2257 (N_2257,N_1642,N_1210);
nor U2258 (N_2258,N_1115,N_1002);
or U2259 (N_2259,N_1792,N_1297);
nor U2260 (N_2260,N_1740,N_1628);
or U2261 (N_2261,N_1990,N_1504);
nand U2262 (N_2262,N_1348,N_1705);
and U2263 (N_2263,N_1463,N_1448);
nand U2264 (N_2264,N_1903,N_1627);
nand U2265 (N_2265,N_1522,N_1922);
xor U2266 (N_2266,N_1045,N_1144);
xor U2267 (N_2267,N_1852,N_1329);
nand U2268 (N_2268,N_1940,N_1209);
and U2269 (N_2269,N_1026,N_1897);
xor U2270 (N_2270,N_1972,N_1019);
nor U2271 (N_2271,N_1798,N_1428);
nor U2272 (N_2272,N_1301,N_1121);
nor U2273 (N_2273,N_1033,N_1531);
or U2274 (N_2274,N_1288,N_1399);
or U2275 (N_2275,N_1397,N_1832);
and U2276 (N_2276,N_1669,N_1543);
nand U2277 (N_2277,N_1044,N_1039);
or U2278 (N_2278,N_1602,N_1434);
nand U2279 (N_2279,N_1060,N_1692);
or U2280 (N_2280,N_1874,N_1760);
xnor U2281 (N_2281,N_1185,N_1239);
and U2282 (N_2282,N_1181,N_1719);
nand U2283 (N_2283,N_1340,N_1929);
and U2284 (N_2284,N_1270,N_1673);
and U2285 (N_2285,N_1097,N_1735);
or U2286 (N_2286,N_1257,N_1186);
nand U2287 (N_2287,N_1321,N_1772);
nor U2288 (N_2288,N_1729,N_1684);
and U2289 (N_2289,N_1211,N_1232);
and U2290 (N_2290,N_1594,N_1882);
nand U2291 (N_2291,N_1398,N_1583);
nand U2292 (N_2292,N_1122,N_1796);
xnor U2293 (N_2293,N_1817,N_1805);
nand U2294 (N_2294,N_1915,N_1640);
or U2295 (N_2295,N_1756,N_1148);
or U2296 (N_2296,N_1872,N_1391);
nand U2297 (N_2297,N_1192,N_1570);
nand U2298 (N_2298,N_1022,N_1324);
nor U2299 (N_2299,N_1885,N_1245);
and U2300 (N_2300,N_1478,N_1387);
or U2301 (N_2301,N_1881,N_1569);
nand U2302 (N_2302,N_1529,N_1051);
or U2303 (N_2303,N_1079,N_1396);
or U2304 (N_2304,N_1377,N_1224);
or U2305 (N_2305,N_1135,N_1068);
nor U2306 (N_2306,N_1737,N_1706);
xor U2307 (N_2307,N_1964,N_1389);
nand U2308 (N_2308,N_1731,N_1549);
xnor U2309 (N_2309,N_1138,N_1278);
nor U2310 (N_2310,N_1985,N_1683);
nor U2311 (N_2311,N_1839,N_1767);
nor U2312 (N_2312,N_1809,N_1284);
nor U2313 (N_2313,N_1891,N_1076);
nand U2314 (N_2314,N_1295,N_1218);
and U2315 (N_2315,N_1854,N_1542);
and U2316 (N_2316,N_1582,N_1253);
and U2317 (N_2317,N_1064,N_1047);
or U2318 (N_2318,N_1084,N_1030);
nand U2319 (N_2319,N_1962,N_1021);
or U2320 (N_2320,N_1814,N_1754);
and U2321 (N_2321,N_1164,N_1343);
and U2322 (N_2322,N_1586,N_1242);
nand U2323 (N_2323,N_1177,N_1254);
and U2324 (N_2324,N_1070,N_1804);
nand U2325 (N_2325,N_1269,N_1667);
nand U2326 (N_2326,N_1910,N_1925);
xnor U2327 (N_2327,N_1621,N_1252);
nor U2328 (N_2328,N_1133,N_1540);
nor U2329 (N_2329,N_1202,N_1317);
and U2330 (N_2330,N_1523,N_1161);
xor U2331 (N_2331,N_1479,N_1293);
or U2332 (N_2332,N_1325,N_1848);
nand U2333 (N_2333,N_1346,N_1989);
nand U2334 (N_2334,N_1069,N_1011);
or U2335 (N_2335,N_1145,N_1422);
nand U2336 (N_2336,N_1576,N_1001);
nand U2337 (N_2337,N_1958,N_1374);
or U2338 (N_2338,N_1844,N_1424);
nor U2339 (N_2339,N_1053,N_1062);
nor U2340 (N_2340,N_1162,N_1227);
and U2341 (N_2341,N_1502,N_1912);
nand U2342 (N_2342,N_1691,N_1679);
nand U2343 (N_2343,N_1467,N_1566);
and U2344 (N_2344,N_1931,N_1183);
nor U2345 (N_2345,N_1718,N_1544);
or U2346 (N_2346,N_1455,N_1052);
nand U2347 (N_2347,N_1924,N_1865);
xor U2348 (N_2348,N_1957,N_1920);
nand U2349 (N_2349,N_1411,N_1778);
or U2350 (N_2350,N_1837,N_1671);
xnor U2351 (N_2351,N_1587,N_1986);
nand U2352 (N_2352,N_1373,N_1799);
xnor U2353 (N_2353,N_1914,N_1025);
nand U2354 (N_2354,N_1091,N_1923);
and U2355 (N_2355,N_1184,N_1336);
or U2356 (N_2356,N_1167,N_1639);
and U2357 (N_2357,N_1777,N_1623);
or U2358 (N_2358,N_1006,N_1205);
nand U2359 (N_2359,N_1846,N_1812);
and U2360 (N_2360,N_1007,N_1700);
xor U2361 (N_2361,N_1054,N_1513);
nand U2362 (N_2362,N_1663,N_1662);
nand U2363 (N_2363,N_1797,N_1472);
xor U2364 (N_2364,N_1495,N_1641);
or U2365 (N_2365,N_1707,N_1620);
nand U2366 (N_2366,N_1607,N_1573);
nand U2367 (N_2367,N_1888,N_1996);
or U2368 (N_2368,N_1630,N_1450);
nor U2369 (N_2369,N_1503,N_1195);
nand U2370 (N_2370,N_1322,N_1159);
or U2371 (N_2371,N_1981,N_1552);
nor U2372 (N_2372,N_1345,N_1083);
nand U2373 (N_2373,N_1483,N_1146);
nor U2374 (N_2374,N_1407,N_1216);
or U2375 (N_2375,N_1977,N_1341);
and U2376 (N_2376,N_1375,N_1916);
and U2377 (N_2377,N_1365,N_1894);
or U2378 (N_2378,N_1579,N_1843);
nand U2379 (N_2379,N_1826,N_1855);
or U2380 (N_2380,N_1717,N_1690);
xor U2381 (N_2381,N_1899,N_1339);
or U2382 (N_2382,N_1457,N_1541);
nand U2383 (N_2383,N_1082,N_1119);
xnor U2384 (N_2384,N_1536,N_1446);
or U2385 (N_2385,N_1421,N_1459);
nor U2386 (N_2386,N_1907,N_1152);
xnor U2387 (N_2387,N_1480,N_1131);
or U2388 (N_2388,N_1858,N_1823);
or U2389 (N_2389,N_1102,N_1175);
or U2390 (N_2390,N_1560,N_1775);
nand U2391 (N_2391,N_1105,N_1568);
nand U2392 (N_2392,N_1458,N_1850);
nor U2393 (N_2393,N_1781,N_1538);
nor U2394 (N_2394,N_1048,N_1676);
nand U2395 (N_2395,N_1364,N_1289);
nand U2396 (N_2396,N_1687,N_1307);
or U2397 (N_2397,N_1072,N_1548);
nor U2398 (N_2398,N_1658,N_1361);
or U2399 (N_2399,N_1596,N_1831);
and U2400 (N_2400,N_1631,N_1231);
nor U2401 (N_2401,N_1221,N_1802);
and U2402 (N_2402,N_1000,N_1755);
xnor U2403 (N_2403,N_1230,N_1112);
nand U2404 (N_2404,N_1485,N_1385);
and U2405 (N_2405,N_1292,N_1534);
or U2406 (N_2406,N_1488,N_1751);
or U2407 (N_2407,N_1789,N_1337);
and U2408 (N_2408,N_1315,N_1564);
nand U2409 (N_2409,N_1418,N_1392);
or U2410 (N_2410,N_1742,N_1359);
or U2411 (N_2411,N_1609,N_1248);
or U2412 (N_2412,N_1104,N_1313);
nor U2413 (N_2413,N_1110,N_1770);
and U2414 (N_2414,N_1892,N_1171);
nand U2415 (N_2415,N_1156,N_1948);
and U2416 (N_2416,N_1807,N_1709);
nor U2417 (N_2417,N_1648,N_1764);
nor U2418 (N_2418,N_1611,N_1333);
nor U2419 (N_2419,N_1261,N_1746);
or U2420 (N_2420,N_1207,N_1851);
or U2421 (N_2421,N_1178,N_1883);
or U2422 (N_2422,N_1193,N_1686);
or U2423 (N_2423,N_1442,N_1674);
xnor U2424 (N_2424,N_1926,N_1134);
nor U2425 (N_2425,N_1730,N_1179);
nor U2426 (N_2426,N_1870,N_1189);
or U2427 (N_2427,N_1349,N_1334);
and U2428 (N_2428,N_1357,N_1008);
nor U2429 (N_2429,N_1968,N_1401);
or U2430 (N_2430,N_1139,N_1260);
and U2431 (N_2431,N_1654,N_1247);
nor U2432 (N_2432,N_1932,N_1423);
nor U2433 (N_2433,N_1895,N_1738);
nor U2434 (N_2434,N_1757,N_1318);
nor U2435 (N_2435,N_1944,N_1616);
or U2436 (N_2436,N_1300,N_1153);
or U2437 (N_2437,N_1517,N_1366);
nand U2438 (N_2438,N_1860,N_1113);
and U2439 (N_2439,N_1491,N_1350);
or U2440 (N_2440,N_1840,N_1617);
nor U2441 (N_2441,N_1040,N_1469);
xnor U2442 (N_2442,N_1312,N_1557);
nand U2443 (N_2443,N_1023,N_1272);
nand U2444 (N_2444,N_1035,N_1279);
nand U2445 (N_2445,N_1158,N_1406);
nor U2446 (N_2446,N_1470,N_1554);
and U2447 (N_2447,N_1410,N_1748);
or U2448 (N_2448,N_1196,N_1029);
nor U2449 (N_2449,N_1215,N_1059);
nor U2450 (N_2450,N_1103,N_1009);
and U2451 (N_2451,N_1622,N_1954);
nand U2452 (N_2452,N_1037,N_1983);
nand U2453 (N_2453,N_1788,N_1132);
or U2454 (N_2454,N_1314,N_1636);
or U2455 (N_2455,N_1701,N_1096);
nand U2456 (N_2456,N_1363,N_1613);
and U2457 (N_2457,N_1508,N_1283);
and U2458 (N_2458,N_1204,N_1842);
or U2459 (N_2459,N_1980,N_1149);
or U2460 (N_2460,N_1332,N_1758);
or U2461 (N_2461,N_1032,N_1524);
nor U2462 (N_2462,N_1825,N_1878);
or U2463 (N_2463,N_1670,N_1499);
nor U2464 (N_2464,N_1578,N_1388);
and U2465 (N_2465,N_1412,N_1938);
or U2466 (N_2466,N_1351,N_1909);
nand U2467 (N_2467,N_1157,N_1402);
nand U2468 (N_2468,N_1655,N_1856);
or U2469 (N_2469,N_1203,N_1902);
or U2470 (N_2470,N_1233,N_1720);
nand U2471 (N_2471,N_1904,N_1294);
and U2472 (N_2472,N_1820,N_1308);
and U2473 (N_2473,N_1123,N_1461);
nand U2474 (N_2474,N_1867,N_1036);
nand U2475 (N_2475,N_1095,N_1970);
nor U2476 (N_2476,N_1017,N_1155);
nand U2477 (N_2477,N_1988,N_1600);
nor U2478 (N_2478,N_1677,N_1299);
and U2479 (N_2479,N_1150,N_1355);
nand U2480 (N_2480,N_1316,N_1409);
and U2481 (N_2481,N_1849,N_1214);
nand U2482 (N_2482,N_1057,N_1246);
or U2483 (N_2483,N_1492,N_1998);
and U2484 (N_2484,N_1055,N_1886);
xor U2485 (N_2485,N_1577,N_1604);
nor U2486 (N_2486,N_1950,N_1952);
or U2487 (N_2487,N_1497,N_1244);
or U2488 (N_2488,N_1126,N_1101);
nor U2489 (N_2489,N_1685,N_1116);
nand U2490 (N_2490,N_1803,N_1027);
xor U2491 (N_2491,N_1610,N_1603);
nand U2492 (N_2492,N_1733,N_1140);
or U2493 (N_2493,N_1829,N_1752);
and U2494 (N_2494,N_1550,N_1786);
and U2495 (N_2495,N_1309,N_1633);
and U2496 (N_2496,N_1378,N_1075);
nand U2497 (N_2497,N_1404,N_1963);
nand U2498 (N_2498,N_1615,N_1666);
nand U2499 (N_2499,N_1969,N_1794);
and U2500 (N_2500,N_1051,N_1130);
nand U2501 (N_2501,N_1278,N_1812);
nand U2502 (N_2502,N_1072,N_1583);
xnor U2503 (N_2503,N_1480,N_1359);
nand U2504 (N_2504,N_1287,N_1571);
and U2505 (N_2505,N_1001,N_1227);
or U2506 (N_2506,N_1702,N_1138);
nand U2507 (N_2507,N_1012,N_1952);
nor U2508 (N_2508,N_1855,N_1223);
and U2509 (N_2509,N_1779,N_1458);
and U2510 (N_2510,N_1898,N_1593);
or U2511 (N_2511,N_1218,N_1853);
nand U2512 (N_2512,N_1153,N_1290);
or U2513 (N_2513,N_1835,N_1402);
and U2514 (N_2514,N_1253,N_1346);
nand U2515 (N_2515,N_1041,N_1317);
or U2516 (N_2516,N_1967,N_1325);
or U2517 (N_2517,N_1798,N_1397);
and U2518 (N_2518,N_1816,N_1385);
or U2519 (N_2519,N_1162,N_1026);
and U2520 (N_2520,N_1577,N_1107);
nor U2521 (N_2521,N_1355,N_1621);
or U2522 (N_2522,N_1270,N_1776);
and U2523 (N_2523,N_1726,N_1033);
or U2524 (N_2524,N_1588,N_1174);
xor U2525 (N_2525,N_1661,N_1935);
nand U2526 (N_2526,N_1644,N_1939);
nand U2527 (N_2527,N_1564,N_1174);
nand U2528 (N_2528,N_1348,N_1699);
and U2529 (N_2529,N_1016,N_1889);
nor U2530 (N_2530,N_1779,N_1672);
and U2531 (N_2531,N_1605,N_1494);
nand U2532 (N_2532,N_1095,N_1389);
nor U2533 (N_2533,N_1473,N_1208);
nor U2534 (N_2534,N_1529,N_1603);
nor U2535 (N_2535,N_1764,N_1067);
nor U2536 (N_2536,N_1642,N_1819);
nand U2537 (N_2537,N_1761,N_1296);
nor U2538 (N_2538,N_1243,N_1933);
nor U2539 (N_2539,N_1728,N_1641);
or U2540 (N_2540,N_1752,N_1149);
nand U2541 (N_2541,N_1471,N_1795);
nor U2542 (N_2542,N_1650,N_1608);
nor U2543 (N_2543,N_1240,N_1959);
or U2544 (N_2544,N_1559,N_1373);
or U2545 (N_2545,N_1104,N_1380);
nand U2546 (N_2546,N_1558,N_1929);
or U2547 (N_2547,N_1400,N_1295);
nand U2548 (N_2548,N_1567,N_1245);
nand U2549 (N_2549,N_1584,N_1793);
nand U2550 (N_2550,N_1056,N_1988);
and U2551 (N_2551,N_1707,N_1742);
nor U2552 (N_2552,N_1292,N_1399);
xnor U2553 (N_2553,N_1976,N_1245);
nor U2554 (N_2554,N_1817,N_1344);
and U2555 (N_2555,N_1789,N_1853);
nor U2556 (N_2556,N_1645,N_1881);
and U2557 (N_2557,N_1845,N_1438);
nor U2558 (N_2558,N_1107,N_1691);
nor U2559 (N_2559,N_1328,N_1689);
nor U2560 (N_2560,N_1080,N_1258);
nand U2561 (N_2561,N_1496,N_1258);
or U2562 (N_2562,N_1541,N_1683);
and U2563 (N_2563,N_1827,N_1024);
nand U2564 (N_2564,N_1185,N_1147);
or U2565 (N_2565,N_1801,N_1376);
nor U2566 (N_2566,N_1546,N_1385);
nor U2567 (N_2567,N_1930,N_1346);
nor U2568 (N_2568,N_1013,N_1036);
nand U2569 (N_2569,N_1052,N_1349);
nand U2570 (N_2570,N_1605,N_1194);
and U2571 (N_2571,N_1438,N_1961);
or U2572 (N_2572,N_1550,N_1943);
or U2573 (N_2573,N_1335,N_1696);
nand U2574 (N_2574,N_1868,N_1557);
or U2575 (N_2575,N_1022,N_1712);
or U2576 (N_2576,N_1623,N_1189);
nand U2577 (N_2577,N_1100,N_1392);
and U2578 (N_2578,N_1952,N_1710);
and U2579 (N_2579,N_1792,N_1148);
or U2580 (N_2580,N_1493,N_1694);
nand U2581 (N_2581,N_1690,N_1326);
and U2582 (N_2582,N_1542,N_1028);
nand U2583 (N_2583,N_1804,N_1370);
nor U2584 (N_2584,N_1283,N_1292);
xnor U2585 (N_2585,N_1590,N_1711);
nor U2586 (N_2586,N_1451,N_1555);
or U2587 (N_2587,N_1219,N_1463);
and U2588 (N_2588,N_1860,N_1129);
and U2589 (N_2589,N_1370,N_1634);
nor U2590 (N_2590,N_1813,N_1630);
and U2591 (N_2591,N_1723,N_1408);
or U2592 (N_2592,N_1757,N_1258);
and U2593 (N_2593,N_1406,N_1504);
nor U2594 (N_2594,N_1066,N_1780);
and U2595 (N_2595,N_1246,N_1891);
nand U2596 (N_2596,N_1040,N_1829);
nor U2597 (N_2597,N_1466,N_1331);
nor U2598 (N_2598,N_1632,N_1639);
nand U2599 (N_2599,N_1862,N_1676);
and U2600 (N_2600,N_1006,N_1203);
or U2601 (N_2601,N_1266,N_1859);
nor U2602 (N_2602,N_1643,N_1305);
xor U2603 (N_2603,N_1292,N_1774);
nand U2604 (N_2604,N_1571,N_1549);
nor U2605 (N_2605,N_1278,N_1374);
and U2606 (N_2606,N_1608,N_1097);
or U2607 (N_2607,N_1182,N_1726);
and U2608 (N_2608,N_1412,N_1288);
nand U2609 (N_2609,N_1727,N_1527);
or U2610 (N_2610,N_1776,N_1811);
nor U2611 (N_2611,N_1710,N_1635);
and U2612 (N_2612,N_1597,N_1073);
nor U2613 (N_2613,N_1191,N_1888);
or U2614 (N_2614,N_1196,N_1277);
and U2615 (N_2615,N_1027,N_1502);
nor U2616 (N_2616,N_1992,N_1960);
and U2617 (N_2617,N_1083,N_1002);
nand U2618 (N_2618,N_1616,N_1090);
and U2619 (N_2619,N_1826,N_1280);
or U2620 (N_2620,N_1085,N_1866);
nor U2621 (N_2621,N_1680,N_1322);
nor U2622 (N_2622,N_1094,N_1406);
and U2623 (N_2623,N_1172,N_1383);
nor U2624 (N_2624,N_1835,N_1227);
and U2625 (N_2625,N_1495,N_1245);
and U2626 (N_2626,N_1193,N_1195);
nor U2627 (N_2627,N_1990,N_1533);
nand U2628 (N_2628,N_1845,N_1554);
or U2629 (N_2629,N_1726,N_1794);
nor U2630 (N_2630,N_1987,N_1615);
and U2631 (N_2631,N_1561,N_1015);
nor U2632 (N_2632,N_1029,N_1851);
nand U2633 (N_2633,N_1106,N_1572);
xor U2634 (N_2634,N_1793,N_1425);
or U2635 (N_2635,N_1340,N_1665);
xor U2636 (N_2636,N_1516,N_1964);
and U2637 (N_2637,N_1208,N_1733);
and U2638 (N_2638,N_1526,N_1586);
or U2639 (N_2639,N_1971,N_1585);
and U2640 (N_2640,N_1364,N_1183);
nand U2641 (N_2641,N_1115,N_1141);
and U2642 (N_2642,N_1769,N_1723);
nand U2643 (N_2643,N_1046,N_1969);
nor U2644 (N_2644,N_1909,N_1433);
nand U2645 (N_2645,N_1648,N_1115);
nor U2646 (N_2646,N_1790,N_1915);
or U2647 (N_2647,N_1233,N_1482);
and U2648 (N_2648,N_1440,N_1137);
nor U2649 (N_2649,N_1456,N_1708);
nand U2650 (N_2650,N_1767,N_1099);
nor U2651 (N_2651,N_1613,N_1896);
nand U2652 (N_2652,N_1606,N_1660);
or U2653 (N_2653,N_1701,N_1694);
nand U2654 (N_2654,N_1877,N_1044);
nand U2655 (N_2655,N_1793,N_1192);
xor U2656 (N_2656,N_1317,N_1583);
or U2657 (N_2657,N_1811,N_1030);
and U2658 (N_2658,N_1122,N_1621);
nand U2659 (N_2659,N_1988,N_1377);
and U2660 (N_2660,N_1276,N_1310);
nand U2661 (N_2661,N_1039,N_1122);
xor U2662 (N_2662,N_1218,N_1359);
or U2663 (N_2663,N_1898,N_1319);
nand U2664 (N_2664,N_1379,N_1660);
nor U2665 (N_2665,N_1876,N_1490);
nor U2666 (N_2666,N_1175,N_1849);
xnor U2667 (N_2667,N_1086,N_1757);
nand U2668 (N_2668,N_1616,N_1070);
or U2669 (N_2669,N_1592,N_1286);
or U2670 (N_2670,N_1926,N_1528);
or U2671 (N_2671,N_1122,N_1194);
or U2672 (N_2672,N_1151,N_1599);
or U2673 (N_2673,N_1139,N_1501);
and U2674 (N_2674,N_1450,N_1767);
and U2675 (N_2675,N_1834,N_1342);
nand U2676 (N_2676,N_1628,N_1961);
and U2677 (N_2677,N_1923,N_1265);
nor U2678 (N_2678,N_1011,N_1312);
nor U2679 (N_2679,N_1165,N_1319);
and U2680 (N_2680,N_1508,N_1673);
and U2681 (N_2681,N_1666,N_1252);
nor U2682 (N_2682,N_1100,N_1399);
and U2683 (N_2683,N_1132,N_1093);
nand U2684 (N_2684,N_1832,N_1378);
and U2685 (N_2685,N_1447,N_1279);
nor U2686 (N_2686,N_1579,N_1889);
or U2687 (N_2687,N_1842,N_1310);
or U2688 (N_2688,N_1861,N_1638);
xor U2689 (N_2689,N_1434,N_1530);
nand U2690 (N_2690,N_1965,N_1253);
and U2691 (N_2691,N_1392,N_1824);
or U2692 (N_2692,N_1710,N_1785);
and U2693 (N_2693,N_1855,N_1953);
nor U2694 (N_2694,N_1212,N_1985);
nor U2695 (N_2695,N_1247,N_1104);
nand U2696 (N_2696,N_1823,N_1182);
nor U2697 (N_2697,N_1280,N_1419);
nand U2698 (N_2698,N_1204,N_1582);
or U2699 (N_2699,N_1966,N_1886);
and U2700 (N_2700,N_1256,N_1695);
nand U2701 (N_2701,N_1578,N_1576);
nand U2702 (N_2702,N_1967,N_1269);
or U2703 (N_2703,N_1573,N_1405);
or U2704 (N_2704,N_1371,N_1272);
or U2705 (N_2705,N_1259,N_1401);
nor U2706 (N_2706,N_1421,N_1507);
nor U2707 (N_2707,N_1855,N_1583);
nor U2708 (N_2708,N_1450,N_1394);
and U2709 (N_2709,N_1678,N_1202);
or U2710 (N_2710,N_1898,N_1639);
xor U2711 (N_2711,N_1993,N_1423);
and U2712 (N_2712,N_1619,N_1679);
nand U2713 (N_2713,N_1821,N_1115);
or U2714 (N_2714,N_1552,N_1025);
nand U2715 (N_2715,N_1180,N_1890);
and U2716 (N_2716,N_1223,N_1190);
nand U2717 (N_2717,N_1489,N_1880);
or U2718 (N_2718,N_1097,N_1909);
xnor U2719 (N_2719,N_1574,N_1629);
and U2720 (N_2720,N_1075,N_1249);
and U2721 (N_2721,N_1035,N_1364);
nand U2722 (N_2722,N_1141,N_1841);
nand U2723 (N_2723,N_1646,N_1167);
nor U2724 (N_2724,N_1891,N_1548);
or U2725 (N_2725,N_1828,N_1291);
nand U2726 (N_2726,N_1100,N_1340);
nand U2727 (N_2727,N_1850,N_1459);
nor U2728 (N_2728,N_1280,N_1575);
nand U2729 (N_2729,N_1561,N_1626);
and U2730 (N_2730,N_1727,N_1445);
nor U2731 (N_2731,N_1649,N_1296);
nand U2732 (N_2732,N_1674,N_1837);
xnor U2733 (N_2733,N_1781,N_1075);
nand U2734 (N_2734,N_1875,N_1626);
or U2735 (N_2735,N_1189,N_1075);
and U2736 (N_2736,N_1901,N_1299);
and U2737 (N_2737,N_1324,N_1838);
nand U2738 (N_2738,N_1245,N_1415);
nor U2739 (N_2739,N_1286,N_1897);
and U2740 (N_2740,N_1888,N_1914);
and U2741 (N_2741,N_1750,N_1182);
nor U2742 (N_2742,N_1888,N_1912);
and U2743 (N_2743,N_1664,N_1548);
xor U2744 (N_2744,N_1083,N_1719);
nor U2745 (N_2745,N_1942,N_1696);
and U2746 (N_2746,N_1442,N_1891);
xor U2747 (N_2747,N_1908,N_1213);
nor U2748 (N_2748,N_1169,N_1454);
and U2749 (N_2749,N_1650,N_1892);
and U2750 (N_2750,N_1761,N_1490);
xor U2751 (N_2751,N_1916,N_1293);
nand U2752 (N_2752,N_1213,N_1132);
nand U2753 (N_2753,N_1895,N_1691);
or U2754 (N_2754,N_1330,N_1085);
xor U2755 (N_2755,N_1165,N_1563);
and U2756 (N_2756,N_1426,N_1921);
or U2757 (N_2757,N_1656,N_1230);
nor U2758 (N_2758,N_1531,N_1918);
xor U2759 (N_2759,N_1574,N_1072);
or U2760 (N_2760,N_1066,N_1205);
or U2761 (N_2761,N_1920,N_1196);
and U2762 (N_2762,N_1771,N_1528);
nand U2763 (N_2763,N_1998,N_1169);
or U2764 (N_2764,N_1229,N_1235);
xnor U2765 (N_2765,N_1515,N_1478);
and U2766 (N_2766,N_1006,N_1365);
and U2767 (N_2767,N_1714,N_1446);
nor U2768 (N_2768,N_1584,N_1673);
xor U2769 (N_2769,N_1265,N_1567);
nor U2770 (N_2770,N_1174,N_1186);
nand U2771 (N_2771,N_1803,N_1959);
nand U2772 (N_2772,N_1245,N_1393);
and U2773 (N_2773,N_1637,N_1593);
or U2774 (N_2774,N_1329,N_1133);
nand U2775 (N_2775,N_1294,N_1631);
xor U2776 (N_2776,N_1334,N_1545);
nand U2777 (N_2777,N_1113,N_1421);
and U2778 (N_2778,N_1690,N_1643);
nor U2779 (N_2779,N_1085,N_1839);
or U2780 (N_2780,N_1903,N_1371);
and U2781 (N_2781,N_1742,N_1721);
nand U2782 (N_2782,N_1939,N_1092);
nor U2783 (N_2783,N_1486,N_1508);
or U2784 (N_2784,N_1062,N_1228);
nor U2785 (N_2785,N_1673,N_1902);
nor U2786 (N_2786,N_1322,N_1242);
nand U2787 (N_2787,N_1942,N_1558);
nand U2788 (N_2788,N_1528,N_1767);
or U2789 (N_2789,N_1070,N_1648);
nor U2790 (N_2790,N_1605,N_1158);
nor U2791 (N_2791,N_1702,N_1083);
and U2792 (N_2792,N_1105,N_1856);
nand U2793 (N_2793,N_1144,N_1572);
nand U2794 (N_2794,N_1613,N_1736);
and U2795 (N_2795,N_1978,N_1009);
nor U2796 (N_2796,N_1835,N_1094);
nand U2797 (N_2797,N_1019,N_1237);
nand U2798 (N_2798,N_1421,N_1873);
and U2799 (N_2799,N_1970,N_1574);
xnor U2800 (N_2800,N_1724,N_1367);
nand U2801 (N_2801,N_1059,N_1509);
xnor U2802 (N_2802,N_1590,N_1827);
nand U2803 (N_2803,N_1691,N_1384);
xnor U2804 (N_2804,N_1035,N_1567);
nand U2805 (N_2805,N_1371,N_1345);
and U2806 (N_2806,N_1990,N_1223);
and U2807 (N_2807,N_1643,N_1228);
nor U2808 (N_2808,N_1064,N_1927);
and U2809 (N_2809,N_1880,N_1989);
nand U2810 (N_2810,N_1224,N_1465);
or U2811 (N_2811,N_1285,N_1507);
or U2812 (N_2812,N_1148,N_1824);
nor U2813 (N_2813,N_1975,N_1443);
or U2814 (N_2814,N_1169,N_1815);
or U2815 (N_2815,N_1470,N_1567);
nand U2816 (N_2816,N_1031,N_1123);
nand U2817 (N_2817,N_1381,N_1733);
nor U2818 (N_2818,N_1649,N_1689);
or U2819 (N_2819,N_1299,N_1840);
xnor U2820 (N_2820,N_1048,N_1470);
or U2821 (N_2821,N_1326,N_1835);
nor U2822 (N_2822,N_1769,N_1212);
nand U2823 (N_2823,N_1327,N_1011);
nand U2824 (N_2824,N_1023,N_1666);
and U2825 (N_2825,N_1554,N_1214);
and U2826 (N_2826,N_1971,N_1340);
or U2827 (N_2827,N_1235,N_1026);
or U2828 (N_2828,N_1800,N_1145);
xor U2829 (N_2829,N_1146,N_1653);
nor U2830 (N_2830,N_1347,N_1378);
nor U2831 (N_2831,N_1873,N_1683);
or U2832 (N_2832,N_1170,N_1711);
nor U2833 (N_2833,N_1047,N_1181);
nor U2834 (N_2834,N_1300,N_1633);
and U2835 (N_2835,N_1104,N_1145);
nand U2836 (N_2836,N_1223,N_1504);
nor U2837 (N_2837,N_1557,N_1845);
nor U2838 (N_2838,N_1378,N_1911);
nor U2839 (N_2839,N_1939,N_1480);
and U2840 (N_2840,N_1000,N_1096);
nor U2841 (N_2841,N_1035,N_1227);
or U2842 (N_2842,N_1585,N_1259);
or U2843 (N_2843,N_1483,N_1882);
xnor U2844 (N_2844,N_1493,N_1466);
nor U2845 (N_2845,N_1147,N_1956);
nor U2846 (N_2846,N_1453,N_1813);
xor U2847 (N_2847,N_1251,N_1852);
xor U2848 (N_2848,N_1433,N_1633);
xnor U2849 (N_2849,N_1008,N_1120);
nand U2850 (N_2850,N_1109,N_1696);
nand U2851 (N_2851,N_1699,N_1083);
nor U2852 (N_2852,N_1099,N_1038);
nand U2853 (N_2853,N_1864,N_1996);
or U2854 (N_2854,N_1715,N_1122);
nand U2855 (N_2855,N_1992,N_1512);
nand U2856 (N_2856,N_1703,N_1137);
nor U2857 (N_2857,N_1206,N_1199);
or U2858 (N_2858,N_1034,N_1180);
and U2859 (N_2859,N_1277,N_1272);
xor U2860 (N_2860,N_1862,N_1479);
nor U2861 (N_2861,N_1129,N_1239);
or U2862 (N_2862,N_1175,N_1066);
nor U2863 (N_2863,N_1178,N_1731);
or U2864 (N_2864,N_1485,N_1627);
or U2865 (N_2865,N_1033,N_1097);
nor U2866 (N_2866,N_1648,N_1687);
nor U2867 (N_2867,N_1471,N_1578);
xor U2868 (N_2868,N_1602,N_1923);
or U2869 (N_2869,N_1389,N_1515);
nand U2870 (N_2870,N_1261,N_1487);
nor U2871 (N_2871,N_1862,N_1675);
nand U2872 (N_2872,N_1665,N_1458);
nor U2873 (N_2873,N_1562,N_1641);
nand U2874 (N_2874,N_1715,N_1184);
and U2875 (N_2875,N_1500,N_1913);
nor U2876 (N_2876,N_1396,N_1065);
nor U2877 (N_2877,N_1394,N_1971);
nand U2878 (N_2878,N_1651,N_1375);
and U2879 (N_2879,N_1710,N_1486);
nand U2880 (N_2880,N_1539,N_1983);
and U2881 (N_2881,N_1270,N_1554);
nor U2882 (N_2882,N_1548,N_1462);
nand U2883 (N_2883,N_1929,N_1366);
nand U2884 (N_2884,N_1255,N_1542);
and U2885 (N_2885,N_1848,N_1851);
nand U2886 (N_2886,N_1968,N_1322);
and U2887 (N_2887,N_1804,N_1658);
nand U2888 (N_2888,N_1946,N_1762);
or U2889 (N_2889,N_1413,N_1365);
nor U2890 (N_2890,N_1622,N_1759);
nor U2891 (N_2891,N_1402,N_1283);
nand U2892 (N_2892,N_1759,N_1387);
nor U2893 (N_2893,N_1369,N_1218);
nor U2894 (N_2894,N_1895,N_1533);
nand U2895 (N_2895,N_1405,N_1729);
xnor U2896 (N_2896,N_1482,N_1532);
and U2897 (N_2897,N_1761,N_1865);
nand U2898 (N_2898,N_1161,N_1458);
nand U2899 (N_2899,N_1980,N_1302);
nand U2900 (N_2900,N_1903,N_1819);
nand U2901 (N_2901,N_1313,N_1550);
xnor U2902 (N_2902,N_1532,N_1621);
or U2903 (N_2903,N_1844,N_1762);
nor U2904 (N_2904,N_1141,N_1397);
and U2905 (N_2905,N_1928,N_1351);
or U2906 (N_2906,N_1991,N_1169);
xor U2907 (N_2907,N_1955,N_1573);
xnor U2908 (N_2908,N_1044,N_1971);
or U2909 (N_2909,N_1488,N_1933);
nor U2910 (N_2910,N_1155,N_1051);
and U2911 (N_2911,N_1373,N_1030);
nand U2912 (N_2912,N_1048,N_1835);
nor U2913 (N_2913,N_1637,N_1516);
and U2914 (N_2914,N_1821,N_1800);
and U2915 (N_2915,N_1801,N_1636);
and U2916 (N_2916,N_1604,N_1513);
xnor U2917 (N_2917,N_1742,N_1094);
nor U2918 (N_2918,N_1620,N_1735);
nand U2919 (N_2919,N_1687,N_1511);
and U2920 (N_2920,N_1417,N_1741);
or U2921 (N_2921,N_1404,N_1886);
or U2922 (N_2922,N_1306,N_1721);
nand U2923 (N_2923,N_1736,N_1394);
or U2924 (N_2924,N_1594,N_1903);
or U2925 (N_2925,N_1863,N_1100);
nor U2926 (N_2926,N_1833,N_1706);
nor U2927 (N_2927,N_1207,N_1255);
nand U2928 (N_2928,N_1481,N_1143);
nand U2929 (N_2929,N_1251,N_1618);
nand U2930 (N_2930,N_1015,N_1741);
or U2931 (N_2931,N_1917,N_1380);
and U2932 (N_2932,N_1929,N_1808);
or U2933 (N_2933,N_1478,N_1293);
nand U2934 (N_2934,N_1548,N_1073);
nand U2935 (N_2935,N_1136,N_1538);
or U2936 (N_2936,N_1936,N_1359);
nor U2937 (N_2937,N_1464,N_1551);
and U2938 (N_2938,N_1547,N_1187);
nor U2939 (N_2939,N_1444,N_1339);
nand U2940 (N_2940,N_1273,N_1488);
and U2941 (N_2941,N_1207,N_1238);
nor U2942 (N_2942,N_1246,N_1744);
and U2943 (N_2943,N_1243,N_1009);
nor U2944 (N_2944,N_1814,N_1376);
or U2945 (N_2945,N_1076,N_1041);
or U2946 (N_2946,N_1760,N_1767);
or U2947 (N_2947,N_1567,N_1119);
xor U2948 (N_2948,N_1350,N_1632);
and U2949 (N_2949,N_1105,N_1217);
and U2950 (N_2950,N_1206,N_1554);
nor U2951 (N_2951,N_1076,N_1362);
xor U2952 (N_2952,N_1256,N_1175);
and U2953 (N_2953,N_1933,N_1054);
or U2954 (N_2954,N_1576,N_1175);
or U2955 (N_2955,N_1634,N_1428);
nand U2956 (N_2956,N_1024,N_1751);
nor U2957 (N_2957,N_1679,N_1178);
and U2958 (N_2958,N_1224,N_1125);
xor U2959 (N_2959,N_1940,N_1396);
or U2960 (N_2960,N_1006,N_1430);
and U2961 (N_2961,N_1091,N_1352);
or U2962 (N_2962,N_1507,N_1649);
xor U2963 (N_2963,N_1506,N_1064);
nor U2964 (N_2964,N_1498,N_1688);
and U2965 (N_2965,N_1229,N_1496);
nor U2966 (N_2966,N_1321,N_1260);
nor U2967 (N_2967,N_1921,N_1938);
or U2968 (N_2968,N_1166,N_1554);
nand U2969 (N_2969,N_1681,N_1309);
or U2970 (N_2970,N_1726,N_1738);
and U2971 (N_2971,N_1006,N_1177);
xor U2972 (N_2972,N_1537,N_1763);
and U2973 (N_2973,N_1192,N_1436);
nor U2974 (N_2974,N_1942,N_1647);
nand U2975 (N_2975,N_1863,N_1225);
nand U2976 (N_2976,N_1209,N_1217);
nor U2977 (N_2977,N_1924,N_1206);
or U2978 (N_2978,N_1547,N_1608);
nor U2979 (N_2979,N_1155,N_1809);
and U2980 (N_2980,N_1381,N_1880);
nand U2981 (N_2981,N_1351,N_1061);
nor U2982 (N_2982,N_1869,N_1183);
xnor U2983 (N_2983,N_1114,N_1982);
or U2984 (N_2984,N_1092,N_1661);
nand U2985 (N_2985,N_1407,N_1187);
or U2986 (N_2986,N_1648,N_1943);
nand U2987 (N_2987,N_1967,N_1050);
and U2988 (N_2988,N_1292,N_1643);
or U2989 (N_2989,N_1931,N_1099);
and U2990 (N_2990,N_1871,N_1601);
or U2991 (N_2991,N_1999,N_1338);
nor U2992 (N_2992,N_1921,N_1127);
nor U2993 (N_2993,N_1383,N_1303);
and U2994 (N_2994,N_1944,N_1361);
or U2995 (N_2995,N_1832,N_1972);
nand U2996 (N_2996,N_1248,N_1610);
or U2997 (N_2997,N_1517,N_1866);
or U2998 (N_2998,N_1064,N_1291);
or U2999 (N_2999,N_1525,N_1916);
xor U3000 (N_3000,N_2199,N_2815);
nand U3001 (N_3001,N_2753,N_2589);
and U3002 (N_3002,N_2288,N_2069);
nand U3003 (N_3003,N_2134,N_2270);
or U3004 (N_3004,N_2120,N_2600);
nand U3005 (N_3005,N_2625,N_2327);
nand U3006 (N_3006,N_2263,N_2894);
nand U3007 (N_3007,N_2216,N_2629);
xor U3008 (N_3008,N_2287,N_2395);
and U3009 (N_3009,N_2247,N_2444);
or U3010 (N_3010,N_2739,N_2141);
nand U3011 (N_3011,N_2361,N_2713);
and U3012 (N_3012,N_2569,N_2382);
nand U3013 (N_3013,N_2766,N_2927);
or U3014 (N_3014,N_2283,N_2236);
nand U3015 (N_3015,N_2539,N_2292);
nand U3016 (N_3016,N_2295,N_2635);
xor U3017 (N_3017,N_2044,N_2404);
or U3018 (N_3018,N_2850,N_2594);
nor U3019 (N_3019,N_2093,N_2091);
nor U3020 (N_3020,N_2061,N_2279);
and U3021 (N_3021,N_2155,N_2585);
nand U3022 (N_3022,N_2343,N_2325);
nor U3023 (N_3023,N_2450,N_2750);
nand U3024 (N_3024,N_2062,N_2023);
nand U3025 (N_3025,N_2043,N_2519);
nand U3026 (N_3026,N_2415,N_2597);
nand U3027 (N_3027,N_2246,N_2743);
nor U3028 (N_3028,N_2363,N_2650);
xor U3029 (N_3029,N_2700,N_2873);
nand U3030 (N_3030,N_2866,N_2803);
or U3031 (N_3031,N_2830,N_2009);
or U3032 (N_3032,N_2747,N_2478);
nor U3033 (N_3033,N_2016,N_2063);
xnor U3034 (N_3034,N_2353,N_2997);
nor U3035 (N_3035,N_2692,N_2150);
or U3036 (N_3036,N_2552,N_2869);
xnor U3037 (N_3037,N_2416,N_2936);
nor U3038 (N_3038,N_2621,N_2748);
nand U3039 (N_3039,N_2351,N_2790);
nand U3040 (N_3040,N_2469,N_2052);
nor U3041 (N_3041,N_2948,N_2724);
and U3042 (N_3042,N_2110,N_2514);
xnor U3043 (N_3043,N_2309,N_2034);
or U3044 (N_3044,N_2065,N_2423);
xor U3045 (N_3045,N_2067,N_2767);
xor U3046 (N_3046,N_2173,N_2699);
and U3047 (N_3047,N_2687,N_2522);
and U3048 (N_3048,N_2860,N_2880);
and U3049 (N_3049,N_2223,N_2544);
or U3050 (N_3050,N_2542,N_2959);
and U3051 (N_3051,N_2234,N_2268);
or U3052 (N_3052,N_2842,N_2992);
nor U3053 (N_3053,N_2780,N_2314);
or U3054 (N_3054,N_2546,N_2810);
nor U3055 (N_3055,N_2411,N_2933);
nand U3056 (N_3056,N_2525,N_2112);
and U3057 (N_3057,N_2328,N_2647);
and U3058 (N_3058,N_2427,N_2963);
or U3059 (N_3059,N_2549,N_2235);
nand U3060 (N_3060,N_2432,N_2829);
and U3061 (N_3061,N_2904,N_2111);
or U3062 (N_3062,N_2551,N_2332);
xnor U3063 (N_3063,N_2886,N_2964);
nand U3064 (N_3064,N_2291,N_2367);
nand U3065 (N_3065,N_2072,N_2045);
and U3066 (N_3066,N_2082,N_2147);
or U3067 (N_3067,N_2706,N_2186);
or U3068 (N_3068,N_2162,N_2012);
nor U3069 (N_3069,N_2505,N_2655);
or U3070 (N_3070,N_2922,N_2376);
nand U3071 (N_3071,N_2387,N_2489);
xnor U3072 (N_3072,N_2897,N_2153);
nor U3073 (N_3073,N_2165,N_2050);
nor U3074 (N_3074,N_2042,N_2709);
nor U3075 (N_3075,N_2078,N_2077);
nand U3076 (N_3076,N_2584,N_2819);
nand U3077 (N_3077,N_2560,N_2211);
and U3078 (N_3078,N_2939,N_2108);
nand U3079 (N_3079,N_2466,N_2280);
and U3080 (N_3080,N_2499,N_2547);
and U3081 (N_3081,N_2051,N_2123);
and U3082 (N_3082,N_2137,N_2430);
nor U3083 (N_3083,N_2758,N_2720);
nand U3084 (N_3084,N_2675,N_2100);
nor U3085 (N_3085,N_2929,N_2437);
nor U3086 (N_3086,N_2285,N_2229);
or U3087 (N_3087,N_2431,N_2126);
and U3088 (N_3088,N_2422,N_2393);
or U3089 (N_3089,N_2386,N_2824);
nor U3090 (N_3090,N_2220,N_2953);
and U3091 (N_3091,N_2985,N_2660);
and U3092 (N_3092,N_2540,N_2474);
nand U3093 (N_3093,N_2070,N_2443);
nand U3094 (N_3094,N_2098,N_2035);
and U3095 (N_3095,N_2172,N_2438);
nand U3096 (N_3096,N_2302,N_2374);
nor U3097 (N_3097,N_2508,N_2218);
nand U3098 (N_3098,N_2973,N_2618);
nand U3099 (N_3099,N_2663,N_2426);
nor U3100 (N_3100,N_2058,N_2079);
nor U3101 (N_3101,N_2678,N_2403);
or U3102 (N_3102,N_2795,N_2490);
nor U3103 (N_3103,N_2520,N_2662);
or U3104 (N_3104,N_2734,N_2686);
and U3105 (N_3105,N_2916,N_2406);
nor U3106 (N_3106,N_2901,N_2360);
and U3107 (N_3107,N_2669,N_2745);
or U3108 (N_3108,N_2467,N_2512);
and U3109 (N_3109,N_2782,N_2844);
and U3110 (N_3110,N_2366,N_2733);
nor U3111 (N_3111,N_2510,N_2825);
and U3112 (N_3112,N_2994,N_2611);
nand U3113 (N_3113,N_2884,N_2591);
xnor U3114 (N_3114,N_2746,N_2846);
nand U3115 (N_3115,N_2129,N_2148);
nand U3116 (N_3116,N_2693,N_2588);
nand U3117 (N_3117,N_2381,N_2476);
and U3118 (N_3118,N_2785,N_2250);
or U3119 (N_3119,N_2481,N_2945);
or U3120 (N_3120,N_2011,N_2947);
or U3121 (N_3121,N_2348,N_2852);
or U3122 (N_3122,N_2380,N_2461);
and U3123 (N_3123,N_2176,N_2170);
and U3124 (N_3124,N_2728,N_2167);
nor U3125 (N_3125,N_2337,N_2056);
or U3126 (N_3126,N_2949,N_2410);
and U3127 (N_3127,N_2541,N_2164);
and U3128 (N_3128,N_2741,N_2762);
nand U3129 (N_3129,N_2453,N_2861);
or U3130 (N_3130,N_2980,N_2344);
nor U3131 (N_3131,N_2193,N_2641);
nor U3132 (N_3132,N_2987,N_2837);
nand U3133 (N_3133,N_2119,N_2131);
and U3134 (N_3134,N_2049,N_2041);
or U3135 (N_3135,N_2666,N_2602);
nor U3136 (N_3136,N_2856,N_2583);
or U3137 (N_3137,N_2265,N_2527);
nand U3138 (N_3138,N_2418,N_2817);
nand U3139 (N_3139,N_2708,N_2071);
or U3140 (N_3140,N_2735,N_2269);
or U3141 (N_3141,N_2075,N_2972);
and U3142 (N_3142,N_2048,N_2849);
nand U3143 (N_3143,N_2854,N_2968);
nor U3144 (N_3144,N_2457,N_2826);
and U3145 (N_3145,N_2214,N_2197);
nand U3146 (N_3146,N_2255,N_2446);
nor U3147 (N_3147,N_2232,N_2695);
nand U3148 (N_3148,N_2240,N_2046);
and U3149 (N_3149,N_2967,N_2339);
or U3150 (N_3150,N_2731,N_2357);
xnor U3151 (N_3151,N_2175,N_2310);
xor U3152 (N_3152,N_2491,N_2862);
nor U3153 (N_3153,N_2350,N_2094);
xor U3154 (N_3154,N_2354,N_2590);
nor U3155 (N_3155,N_2838,N_2937);
nand U3156 (N_3156,N_2931,N_2952);
nand U3157 (N_3157,N_2145,N_2483);
or U3158 (N_3158,N_2482,N_2352);
or U3159 (N_3159,N_2978,N_2631);
or U3160 (N_3160,N_2245,N_2191);
and U3161 (N_3161,N_2614,N_2778);
and U3162 (N_3162,N_2832,N_2847);
nor U3163 (N_3163,N_2801,N_2694);
nor U3164 (N_3164,N_2993,N_2412);
xor U3165 (N_3165,N_2524,N_2441);
and U3166 (N_3166,N_2681,N_2607);
nor U3167 (N_3167,N_2005,N_2304);
nor U3168 (N_3168,N_2535,N_2646);
nand U3169 (N_3169,N_2400,N_2598);
or U3170 (N_3170,N_2113,N_2651);
nor U3171 (N_3171,N_2417,N_2447);
or U3172 (N_3172,N_2941,N_2433);
nor U3173 (N_3173,N_2096,N_2492);
xnor U3174 (N_3174,N_2823,N_2106);
nor U3175 (N_3175,N_2143,N_2809);
or U3176 (N_3176,N_2715,N_2299);
nand U3177 (N_3177,N_2317,N_2135);
or U3178 (N_3178,N_2306,N_2974);
and U3179 (N_3179,N_2887,N_2771);
nor U3180 (N_3180,N_2996,N_2434);
nand U3181 (N_3181,N_2454,N_2813);
nand U3182 (N_3182,N_2338,N_2924);
and U3183 (N_3183,N_2772,N_2375);
nor U3184 (N_3184,N_2870,N_2217);
or U3185 (N_3185,N_2800,N_2981);
or U3186 (N_3186,N_2789,N_2875);
nand U3187 (N_3187,N_2811,N_2168);
nor U3188 (N_3188,N_2909,N_2455);
nand U3189 (N_3189,N_2362,N_2388);
xor U3190 (N_3190,N_2623,N_2190);
and U3191 (N_3191,N_2840,N_2272);
or U3192 (N_3192,N_2534,N_2448);
or U3193 (N_3193,N_2572,N_2054);
nand U3194 (N_3194,N_2301,N_2315);
or U3195 (N_3195,N_2064,N_2845);
xor U3196 (N_3196,N_2567,N_2683);
and U3197 (N_3197,N_2892,N_2877);
nand U3198 (N_3198,N_2596,N_2526);
and U3199 (N_3199,N_2127,N_2725);
or U3200 (N_3200,N_2806,N_2359);
nor U3201 (N_3201,N_2898,N_2961);
or U3202 (N_3202,N_2452,N_2274);
xor U3203 (N_3203,N_2495,N_2321);
nand U3204 (N_3204,N_2765,N_2798);
nand U3205 (N_3205,N_2865,N_2885);
and U3206 (N_3206,N_2133,N_2580);
nor U3207 (N_3207,N_2773,N_2679);
and U3208 (N_3208,N_2032,N_2958);
nor U3209 (N_3209,N_2221,N_2730);
or U3210 (N_3210,N_2358,N_2521);
or U3211 (N_3211,N_2289,N_2084);
nor U3212 (N_3212,N_2297,N_2156);
or U3213 (N_3213,N_2872,N_2039);
or U3214 (N_3214,N_2515,N_2528);
nand U3215 (N_3215,N_2341,N_2755);
nand U3216 (N_3216,N_2074,N_2073);
nand U3217 (N_3217,N_2013,N_2424);
nor U3218 (N_3218,N_2595,N_2570);
nand U3219 (N_3219,N_2969,N_2468);
or U3220 (N_3220,N_2083,N_2021);
nand U3221 (N_3221,N_2557,N_2639);
or U3222 (N_3222,N_2578,N_2575);
nand U3223 (N_3223,N_2857,N_2905);
nand U3224 (N_3224,N_2209,N_2970);
nand U3225 (N_3225,N_2346,N_2494);
or U3226 (N_3226,N_2037,N_2930);
or U3227 (N_3227,N_2060,N_2312);
and U3228 (N_3228,N_2896,N_2889);
and U3229 (N_3229,N_2435,N_2159);
or U3230 (N_3230,N_2533,N_2919);
or U3231 (N_3231,N_2227,N_2258);
or U3232 (N_3232,N_2334,N_2727);
xor U3233 (N_3233,N_2429,N_2576);
nor U3234 (N_3234,N_2900,N_2685);
nor U3235 (N_3235,N_2022,N_2207);
nand U3236 (N_3236,N_2883,N_2226);
nor U3237 (N_3237,N_2702,N_2445);
or U3238 (N_3238,N_2210,N_2006);
nand U3239 (N_3239,N_2744,N_2821);
nand U3240 (N_3240,N_2200,N_2068);
or U3241 (N_3241,N_2355,N_2053);
or U3242 (N_3242,N_2726,N_2248);
nand U3243 (N_3243,N_2564,N_2657);
nand U3244 (N_3244,N_2036,N_2237);
xor U3245 (N_3245,N_2116,N_2178);
or U3246 (N_3246,N_2506,N_2238);
nand U3247 (N_3247,N_2910,N_2105);
nor U3248 (N_3248,N_2373,N_2488);
and U3249 (N_3249,N_2389,N_2398);
nor U3250 (N_3250,N_2954,N_2473);
or U3251 (N_3251,N_2899,N_2665);
or U3252 (N_3252,N_2462,N_2254);
xor U3253 (N_3253,N_2493,N_2076);
nor U3254 (N_3254,N_2703,N_2977);
nand U3255 (N_3255,N_2776,N_2950);
and U3256 (N_3256,N_2960,N_2277);
nand U3257 (N_3257,N_2554,N_2764);
and U3258 (N_3258,N_2464,N_2169);
xor U3259 (N_3259,N_2836,N_2463);
and U3260 (N_3260,N_2719,N_2257);
xnor U3261 (N_3261,N_2117,N_2787);
nor U3262 (N_3262,N_2878,N_2957);
and U3263 (N_3263,N_2252,N_2982);
or U3264 (N_3264,N_2436,N_2517);
nand U3265 (N_3265,N_2305,N_2293);
nand U3266 (N_3266,N_2523,N_2017);
and U3267 (N_3267,N_2440,N_2859);
and U3268 (N_3268,N_2729,N_2636);
or U3269 (N_3269,N_2260,N_2956);
nor U3270 (N_3270,N_2322,N_2059);
nand U3271 (N_3271,N_2251,N_2089);
nor U3272 (N_3272,N_2749,N_2951);
and U3273 (N_3273,N_2907,N_2763);
and U3274 (N_3274,N_2477,N_2802);
nor U3275 (N_3275,N_2278,N_2989);
nor U3276 (N_3276,N_2784,N_2654);
nand U3277 (N_3277,N_2616,N_2777);
nand U3278 (N_3278,N_2653,N_2608);
and U3279 (N_3279,N_2485,N_2736);
xor U3280 (N_3280,N_2814,N_2808);
or U3281 (N_3281,N_2313,N_2303);
nor U3282 (N_3282,N_2101,N_2273);
nor U3283 (N_3283,N_2047,N_2498);
and U3284 (N_3284,N_2384,N_2475);
and U3285 (N_3285,N_2668,N_2827);
or U3286 (N_3286,N_2031,N_2871);
nor U3287 (N_3287,N_2599,N_2874);
nor U3288 (N_3288,N_2171,N_2356);
and U3289 (N_3289,N_2722,N_2645);
and U3290 (N_3290,N_2912,N_2697);
nor U3291 (N_3291,N_2691,N_2090);
nor U3292 (N_3292,N_2807,N_2563);
nor U3293 (N_3293,N_2192,N_2030);
or U3294 (N_3294,N_2613,N_2586);
nand U3295 (N_3295,N_2561,N_2876);
nor U3296 (N_3296,N_2080,N_2984);
nor U3297 (N_3297,N_2449,N_2818);
xnor U3298 (N_3298,N_2264,N_2504);
nor U3299 (N_3299,N_2760,N_2562);
nand U3300 (N_3300,N_2181,N_2673);
or U3301 (N_3301,N_2307,N_2935);
and U3302 (N_3302,N_2319,N_2109);
and U3303 (N_3303,N_2055,N_2003);
and U3304 (N_3304,N_2125,N_2228);
nand U3305 (N_3305,N_2414,N_2834);
nand U3306 (N_3306,N_2369,N_2442);
nand U3307 (N_3307,N_2532,N_2027);
and U3308 (N_3308,N_2333,N_2835);
xor U3309 (N_3309,N_2975,N_2925);
nor U3310 (N_3310,N_2470,N_2550);
or U3311 (N_3311,N_2225,N_2007);
xnor U3312 (N_3312,N_2378,N_2831);
nand U3313 (N_3313,N_2995,N_2224);
and U3314 (N_3314,N_2243,N_2188);
nor U3315 (N_3315,N_2509,N_2717);
or U3316 (N_3316,N_2266,N_2511);
and U3317 (N_3317,N_2256,N_2710);
or U3318 (N_3318,N_2843,N_2775);
nor U3319 (N_3319,N_2066,N_2316);
xnor U3320 (N_3320,N_2940,N_2617);
xnor U3321 (N_3321,N_2918,N_2841);
or U3322 (N_3322,N_2020,N_2913);
xnor U3323 (N_3323,N_2401,N_2204);
and U3324 (N_3324,N_2132,N_2010);
or U3325 (N_3325,N_2128,N_2342);
nor U3326 (N_3326,N_2456,N_2026);
nor U3327 (N_3327,N_2480,N_2965);
nor U3328 (N_3328,N_2425,N_2943);
nand U3329 (N_3329,N_2737,N_2115);
or U3330 (N_3330,N_2095,N_2839);
nand U3331 (N_3331,N_2379,N_2926);
nand U3332 (N_3332,N_2057,N_2548);
nor U3333 (N_3333,N_2507,N_2121);
and U3334 (N_3334,N_2704,N_2259);
xor U3335 (N_3335,N_2915,N_2976);
and U3336 (N_3336,N_2140,N_2428);
or U3337 (N_3337,N_2868,N_2986);
nor U3338 (N_3338,N_2282,N_2160);
xor U3339 (N_3339,N_2705,N_2215);
nand U3340 (N_3340,N_2212,N_2472);
or U3341 (N_3341,N_2122,N_2104);
and U3342 (N_3342,N_2604,N_2555);
and U3343 (N_3343,N_2684,N_2497);
or U3344 (N_3344,N_2769,N_2331);
nor U3345 (N_3345,N_2920,N_2628);
and U3346 (N_3346,N_2962,N_2372);
nand U3347 (N_3347,N_2024,N_2275);
nor U3348 (N_3348,N_2500,N_2391);
xor U3349 (N_3349,N_2002,N_2902);
nand U3350 (N_3350,N_2187,N_2637);
or U3351 (N_3351,N_2543,N_2139);
or U3352 (N_3352,N_2324,N_2674);
nor U3353 (N_3353,N_2603,N_2081);
and U3354 (N_3354,N_2882,N_2182);
and U3355 (N_3355,N_2318,N_2040);
nor U3356 (N_3356,N_2102,N_2579);
nand U3357 (N_3357,N_2848,N_2999);
nor U3358 (N_3358,N_2788,N_2015);
or U3359 (N_3359,N_2502,N_2183);
nor U3360 (N_3360,N_2242,N_2938);
and U3361 (N_3361,N_2833,N_2759);
nand U3362 (N_3362,N_2670,N_2088);
and U3363 (N_3363,N_2479,N_2465);
xor U3364 (N_3364,N_2157,N_2619);
and U3365 (N_3365,N_2680,N_2000);
and U3366 (N_3366,N_2677,N_2336);
or U3367 (N_3367,N_2537,N_2891);
nand U3368 (N_3368,N_2791,N_2556);
and U3369 (N_3369,N_2484,N_2701);
nand U3370 (N_3370,N_2349,N_2718);
and U3371 (N_3371,N_2364,N_2368);
nand U3372 (N_3372,N_2103,N_2971);
or U3373 (N_3373,N_2652,N_2858);
xor U3374 (N_3374,N_2149,N_2408);
nor U3375 (N_3375,N_2231,N_2195);
xor U3376 (N_3376,N_2656,N_2142);
and U3377 (N_3377,N_2851,N_2659);
and U3378 (N_3378,N_2714,N_2955);
xnor U3379 (N_3379,N_2086,N_2796);
nand U3380 (N_3380,N_2300,N_2107);
and U3381 (N_3381,N_2213,N_2184);
and U3382 (N_3382,N_2138,N_2676);
xnor U3383 (N_3383,N_2723,N_2262);
nand U3384 (N_3384,N_2460,N_2756);
or U3385 (N_3385,N_2752,N_2179);
xor U3386 (N_3386,N_2205,N_2863);
or U3387 (N_3387,N_2879,N_2166);
nor U3388 (N_3388,N_2638,N_2163);
or U3389 (N_3389,N_2601,N_2185);
or U3390 (N_3390,N_2624,N_2249);
or U3391 (N_3391,N_2308,N_2370);
or U3392 (N_3392,N_2593,N_2592);
nand U3393 (N_3393,N_2014,N_2087);
nor U3394 (N_3394,N_2696,N_2893);
and U3395 (N_3395,N_2487,N_2581);
nand U3396 (N_3396,N_2419,N_2864);
or U3397 (N_3397,N_2392,N_2921);
nand U3398 (N_3398,N_2241,N_2545);
nor U3399 (N_3399,N_2501,N_2587);
nor U3400 (N_3400,N_2151,N_2559);
xnor U3401 (N_3401,N_2627,N_2740);
or U3402 (N_3402,N_2394,N_2712);
xor U3403 (N_3403,N_2124,N_2664);
nor U3404 (N_3404,N_2486,N_2805);
or U3405 (N_3405,N_2711,N_2405);
and U3406 (N_3406,N_2296,N_2198);
and U3407 (N_3407,N_2038,N_2085);
nor U3408 (N_3408,N_2661,N_2794);
or U3409 (N_3409,N_2643,N_2732);
nand U3410 (N_3410,N_2018,N_2397);
nor U3411 (N_3411,N_2001,N_2738);
xor U3412 (N_3412,N_2667,N_2320);
nand U3413 (N_3413,N_2371,N_2816);
and U3414 (N_3414,N_2201,N_2329);
nand U3415 (N_3415,N_2294,N_2610);
or U3416 (N_3416,N_2914,N_2154);
or U3417 (N_3417,N_2853,N_2158);
and U3418 (N_3418,N_2144,N_2496);
and U3419 (N_3419,N_2906,N_2253);
nand U3420 (N_3420,N_2136,N_2612);
nand U3421 (N_3421,N_2458,N_2029);
or U3422 (N_3422,N_2281,N_2658);
xnor U3423 (N_3423,N_2233,N_2689);
xor U3424 (N_3424,N_2622,N_2377);
xor U3425 (N_3425,N_2267,N_2707);
nand U3426 (N_3426,N_2630,N_2615);
nor U3427 (N_3427,N_2439,N_2908);
or U3428 (N_3428,N_2340,N_2385);
nand U3429 (N_3429,N_2751,N_2152);
or U3430 (N_3430,N_2530,N_2399);
or U3431 (N_3431,N_2761,N_2516);
or U3432 (N_3432,N_2895,N_2503);
nand U3433 (N_3433,N_2632,N_2928);
nor U3434 (N_3434,N_2208,N_2742);
nor U3435 (N_3435,N_2271,N_2130);
nor U3436 (N_3436,N_2323,N_2311);
or U3437 (N_3437,N_2983,N_2290);
nand U3438 (N_3438,N_2531,N_2793);
or U3439 (N_3439,N_2558,N_2609);
nand U3440 (N_3440,N_2536,N_2513);
and U3441 (N_3441,N_2903,N_2390);
nor U3442 (N_3442,N_2917,N_2177);
xnor U3443 (N_3443,N_2407,N_2239);
or U3444 (N_3444,N_2345,N_2222);
nand U3445 (N_3445,N_2008,N_2161);
and U3446 (N_3446,N_2451,N_2383);
or U3447 (N_3447,N_2990,N_2518);
or U3448 (N_3448,N_2754,N_2786);
nand U3449 (N_3449,N_2261,N_2529);
nor U3450 (N_3450,N_2409,N_2716);
xor U3451 (N_3451,N_2988,N_2206);
xnor U3452 (N_3452,N_2792,N_2998);
xor U3453 (N_3453,N_2326,N_2768);
nor U3454 (N_3454,N_2019,N_2890);
and U3455 (N_3455,N_2025,N_2538);
nand U3456 (N_3456,N_2923,N_2779);
xor U3457 (N_3457,N_2888,N_2196);
or U3458 (N_3458,N_2781,N_2979);
or U3459 (N_3459,N_2099,N_2620);
and U3460 (N_3460,N_2114,N_2721);
or U3461 (N_3461,N_2932,N_2180);
or U3462 (N_3462,N_2966,N_2413);
xnor U3463 (N_3463,N_2626,N_2276);
xor U3464 (N_3464,N_2881,N_2671);
nand U3465 (N_3465,N_2991,N_2553);
nor U3466 (N_3466,N_2634,N_2867);
or U3467 (N_3467,N_2330,N_2946);
and U3468 (N_3468,N_2644,N_2420);
nand U3469 (N_3469,N_2298,N_2934);
xor U3470 (N_3470,N_2230,N_2347);
nor U3471 (N_3471,N_2574,N_2335);
xor U3472 (N_3472,N_2244,N_2202);
nand U3473 (N_3473,N_2757,N_2284);
nor U3474 (N_3474,N_2797,N_2566);
nand U3475 (N_3475,N_2640,N_2004);
nor U3476 (N_3476,N_2146,N_2855);
or U3477 (N_3477,N_2421,N_2820);
and U3478 (N_3478,N_2774,N_2944);
and U3479 (N_3479,N_2565,N_2118);
and U3480 (N_3480,N_2286,N_2648);
nor U3481 (N_3481,N_2573,N_2582);
nand U3482 (N_3482,N_2189,N_2783);
or U3483 (N_3483,N_2672,N_2822);
or U3484 (N_3484,N_2804,N_2682);
nand U3485 (N_3485,N_2688,N_2033);
nand U3486 (N_3486,N_2365,N_2577);
or U3487 (N_3487,N_2812,N_2606);
and U3488 (N_3488,N_2770,N_2174);
or U3489 (N_3489,N_2698,N_2194);
and U3490 (N_3490,N_2396,N_2642);
nor U3491 (N_3491,N_2568,N_2942);
or U3492 (N_3492,N_2459,N_2690);
nand U3493 (N_3493,N_2571,N_2911);
and U3494 (N_3494,N_2028,N_2828);
xnor U3495 (N_3495,N_2402,N_2649);
nor U3496 (N_3496,N_2097,N_2799);
nor U3497 (N_3497,N_2219,N_2605);
nand U3498 (N_3498,N_2471,N_2203);
or U3499 (N_3499,N_2092,N_2633);
nand U3500 (N_3500,N_2921,N_2565);
nor U3501 (N_3501,N_2127,N_2430);
or U3502 (N_3502,N_2721,N_2013);
nand U3503 (N_3503,N_2433,N_2018);
nor U3504 (N_3504,N_2988,N_2364);
and U3505 (N_3505,N_2570,N_2738);
and U3506 (N_3506,N_2712,N_2930);
and U3507 (N_3507,N_2523,N_2374);
or U3508 (N_3508,N_2396,N_2892);
nor U3509 (N_3509,N_2676,N_2362);
and U3510 (N_3510,N_2060,N_2197);
and U3511 (N_3511,N_2840,N_2935);
xnor U3512 (N_3512,N_2253,N_2041);
nand U3513 (N_3513,N_2651,N_2078);
nor U3514 (N_3514,N_2853,N_2658);
and U3515 (N_3515,N_2608,N_2862);
or U3516 (N_3516,N_2391,N_2421);
nand U3517 (N_3517,N_2042,N_2735);
nor U3518 (N_3518,N_2388,N_2899);
xnor U3519 (N_3519,N_2795,N_2285);
and U3520 (N_3520,N_2706,N_2024);
and U3521 (N_3521,N_2448,N_2987);
or U3522 (N_3522,N_2310,N_2928);
and U3523 (N_3523,N_2824,N_2034);
nand U3524 (N_3524,N_2834,N_2090);
xnor U3525 (N_3525,N_2710,N_2632);
xor U3526 (N_3526,N_2109,N_2554);
or U3527 (N_3527,N_2155,N_2481);
nand U3528 (N_3528,N_2282,N_2957);
and U3529 (N_3529,N_2758,N_2247);
xor U3530 (N_3530,N_2357,N_2932);
nor U3531 (N_3531,N_2516,N_2813);
xnor U3532 (N_3532,N_2232,N_2169);
nand U3533 (N_3533,N_2545,N_2645);
nand U3534 (N_3534,N_2307,N_2591);
or U3535 (N_3535,N_2884,N_2326);
or U3536 (N_3536,N_2316,N_2824);
nor U3537 (N_3537,N_2481,N_2747);
or U3538 (N_3538,N_2664,N_2195);
nand U3539 (N_3539,N_2411,N_2649);
or U3540 (N_3540,N_2391,N_2640);
and U3541 (N_3541,N_2321,N_2670);
nand U3542 (N_3542,N_2186,N_2972);
nand U3543 (N_3543,N_2280,N_2050);
nor U3544 (N_3544,N_2638,N_2079);
or U3545 (N_3545,N_2102,N_2568);
or U3546 (N_3546,N_2435,N_2782);
nor U3547 (N_3547,N_2328,N_2662);
or U3548 (N_3548,N_2909,N_2317);
or U3549 (N_3549,N_2835,N_2121);
and U3550 (N_3550,N_2869,N_2482);
nand U3551 (N_3551,N_2286,N_2141);
or U3552 (N_3552,N_2927,N_2476);
or U3553 (N_3553,N_2217,N_2261);
or U3554 (N_3554,N_2469,N_2839);
nand U3555 (N_3555,N_2854,N_2199);
or U3556 (N_3556,N_2702,N_2844);
nor U3557 (N_3557,N_2439,N_2927);
or U3558 (N_3558,N_2288,N_2523);
or U3559 (N_3559,N_2937,N_2804);
nor U3560 (N_3560,N_2258,N_2573);
nand U3561 (N_3561,N_2665,N_2424);
and U3562 (N_3562,N_2037,N_2574);
and U3563 (N_3563,N_2182,N_2510);
and U3564 (N_3564,N_2025,N_2632);
nand U3565 (N_3565,N_2259,N_2267);
and U3566 (N_3566,N_2991,N_2311);
or U3567 (N_3567,N_2827,N_2947);
and U3568 (N_3568,N_2947,N_2514);
or U3569 (N_3569,N_2792,N_2683);
nand U3570 (N_3570,N_2040,N_2620);
nand U3571 (N_3571,N_2178,N_2609);
and U3572 (N_3572,N_2915,N_2094);
nor U3573 (N_3573,N_2316,N_2341);
xor U3574 (N_3574,N_2437,N_2219);
nor U3575 (N_3575,N_2203,N_2161);
nand U3576 (N_3576,N_2419,N_2264);
or U3577 (N_3577,N_2840,N_2758);
xnor U3578 (N_3578,N_2281,N_2522);
and U3579 (N_3579,N_2863,N_2442);
or U3580 (N_3580,N_2686,N_2428);
nand U3581 (N_3581,N_2052,N_2742);
or U3582 (N_3582,N_2096,N_2869);
nor U3583 (N_3583,N_2111,N_2728);
or U3584 (N_3584,N_2262,N_2009);
nand U3585 (N_3585,N_2402,N_2861);
nand U3586 (N_3586,N_2430,N_2760);
and U3587 (N_3587,N_2851,N_2111);
or U3588 (N_3588,N_2119,N_2576);
nor U3589 (N_3589,N_2453,N_2535);
and U3590 (N_3590,N_2980,N_2823);
or U3591 (N_3591,N_2257,N_2460);
nor U3592 (N_3592,N_2741,N_2904);
nand U3593 (N_3593,N_2002,N_2123);
or U3594 (N_3594,N_2751,N_2720);
and U3595 (N_3595,N_2329,N_2227);
nand U3596 (N_3596,N_2495,N_2651);
xnor U3597 (N_3597,N_2233,N_2319);
and U3598 (N_3598,N_2091,N_2764);
and U3599 (N_3599,N_2065,N_2929);
nor U3600 (N_3600,N_2125,N_2641);
or U3601 (N_3601,N_2951,N_2923);
xor U3602 (N_3602,N_2327,N_2390);
or U3603 (N_3603,N_2558,N_2586);
nor U3604 (N_3604,N_2633,N_2810);
nor U3605 (N_3605,N_2538,N_2921);
and U3606 (N_3606,N_2856,N_2956);
and U3607 (N_3607,N_2833,N_2544);
and U3608 (N_3608,N_2699,N_2244);
nor U3609 (N_3609,N_2452,N_2874);
nor U3610 (N_3610,N_2402,N_2363);
and U3611 (N_3611,N_2941,N_2296);
nor U3612 (N_3612,N_2494,N_2140);
and U3613 (N_3613,N_2026,N_2358);
or U3614 (N_3614,N_2530,N_2242);
nand U3615 (N_3615,N_2854,N_2907);
nor U3616 (N_3616,N_2680,N_2278);
or U3617 (N_3617,N_2019,N_2530);
and U3618 (N_3618,N_2736,N_2952);
and U3619 (N_3619,N_2850,N_2824);
or U3620 (N_3620,N_2982,N_2292);
nand U3621 (N_3621,N_2605,N_2710);
and U3622 (N_3622,N_2762,N_2730);
xnor U3623 (N_3623,N_2601,N_2790);
and U3624 (N_3624,N_2165,N_2448);
xor U3625 (N_3625,N_2321,N_2691);
nor U3626 (N_3626,N_2443,N_2938);
nor U3627 (N_3627,N_2001,N_2039);
nor U3628 (N_3628,N_2270,N_2953);
and U3629 (N_3629,N_2725,N_2243);
xor U3630 (N_3630,N_2116,N_2224);
nor U3631 (N_3631,N_2223,N_2525);
nand U3632 (N_3632,N_2931,N_2140);
nand U3633 (N_3633,N_2292,N_2819);
or U3634 (N_3634,N_2970,N_2106);
nand U3635 (N_3635,N_2725,N_2594);
or U3636 (N_3636,N_2137,N_2278);
nor U3637 (N_3637,N_2033,N_2765);
nand U3638 (N_3638,N_2536,N_2443);
nor U3639 (N_3639,N_2721,N_2300);
nand U3640 (N_3640,N_2397,N_2278);
nor U3641 (N_3641,N_2431,N_2598);
nand U3642 (N_3642,N_2504,N_2049);
or U3643 (N_3643,N_2086,N_2575);
or U3644 (N_3644,N_2739,N_2091);
and U3645 (N_3645,N_2214,N_2589);
xor U3646 (N_3646,N_2576,N_2802);
and U3647 (N_3647,N_2611,N_2110);
nand U3648 (N_3648,N_2389,N_2209);
or U3649 (N_3649,N_2902,N_2156);
or U3650 (N_3650,N_2096,N_2859);
nor U3651 (N_3651,N_2524,N_2652);
nand U3652 (N_3652,N_2496,N_2369);
nor U3653 (N_3653,N_2959,N_2357);
or U3654 (N_3654,N_2760,N_2879);
or U3655 (N_3655,N_2994,N_2667);
or U3656 (N_3656,N_2958,N_2787);
nand U3657 (N_3657,N_2025,N_2688);
xnor U3658 (N_3658,N_2264,N_2625);
or U3659 (N_3659,N_2851,N_2131);
or U3660 (N_3660,N_2722,N_2332);
or U3661 (N_3661,N_2733,N_2693);
xnor U3662 (N_3662,N_2613,N_2081);
nor U3663 (N_3663,N_2769,N_2557);
nand U3664 (N_3664,N_2293,N_2635);
or U3665 (N_3665,N_2278,N_2418);
and U3666 (N_3666,N_2304,N_2133);
or U3667 (N_3667,N_2824,N_2741);
and U3668 (N_3668,N_2977,N_2671);
and U3669 (N_3669,N_2710,N_2798);
nand U3670 (N_3670,N_2491,N_2643);
xnor U3671 (N_3671,N_2908,N_2675);
nand U3672 (N_3672,N_2857,N_2833);
nor U3673 (N_3673,N_2005,N_2878);
xor U3674 (N_3674,N_2414,N_2423);
or U3675 (N_3675,N_2980,N_2260);
xnor U3676 (N_3676,N_2021,N_2848);
and U3677 (N_3677,N_2082,N_2526);
nor U3678 (N_3678,N_2553,N_2279);
or U3679 (N_3679,N_2088,N_2229);
xnor U3680 (N_3680,N_2666,N_2205);
nand U3681 (N_3681,N_2091,N_2455);
nor U3682 (N_3682,N_2695,N_2218);
xor U3683 (N_3683,N_2119,N_2760);
or U3684 (N_3684,N_2911,N_2420);
nand U3685 (N_3685,N_2633,N_2234);
and U3686 (N_3686,N_2419,N_2138);
xor U3687 (N_3687,N_2027,N_2825);
or U3688 (N_3688,N_2783,N_2763);
xnor U3689 (N_3689,N_2973,N_2231);
and U3690 (N_3690,N_2730,N_2984);
and U3691 (N_3691,N_2140,N_2340);
nor U3692 (N_3692,N_2114,N_2122);
nand U3693 (N_3693,N_2415,N_2537);
nand U3694 (N_3694,N_2972,N_2425);
and U3695 (N_3695,N_2501,N_2709);
xnor U3696 (N_3696,N_2400,N_2659);
and U3697 (N_3697,N_2565,N_2619);
xnor U3698 (N_3698,N_2042,N_2933);
or U3699 (N_3699,N_2625,N_2914);
or U3700 (N_3700,N_2810,N_2338);
xor U3701 (N_3701,N_2009,N_2003);
nand U3702 (N_3702,N_2134,N_2606);
nand U3703 (N_3703,N_2343,N_2262);
and U3704 (N_3704,N_2400,N_2176);
nor U3705 (N_3705,N_2315,N_2502);
nor U3706 (N_3706,N_2588,N_2792);
and U3707 (N_3707,N_2856,N_2539);
xnor U3708 (N_3708,N_2420,N_2060);
nand U3709 (N_3709,N_2283,N_2912);
nand U3710 (N_3710,N_2814,N_2567);
nand U3711 (N_3711,N_2538,N_2719);
nand U3712 (N_3712,N_2984,N_2361);
and U3713 (N_3713,N_2522,N_2896);
and U3714 (N_3714,N_2907,N_2290);
nor U3715 (N_3715,N_2594,N_2592);
nand U3716 (N_3716,N_2788,N_2836);
nor U3717 (N_3717,N_2364,N_2393);
xor U3718 (N_3718,N_2313,N_2922);
nor U3719 (N_3719,N_2705,N_2915);
xnor U3720 (N_3720,N_2073,N_2802);
or U3721 (N_3721,N_2507,N_2351);
nor U3722 (N_3722,N_2439,N_2125);
nor U3723 (N_3723,N_2679,N_2102);
and U3724 (N_3724,N_2101,N_2226);
and U3725 (N_3725,N_2121,N_2257);
and U3726 (N_3726,N_2877,N_2105);
xnor U3727 (N_3727,N_2871,N_2574);
and U3728 (N_3728,N_2625,N_2329);
nor U3729 (N_3729,N_2234,N_2249);
and U3730 (N_3730,N_2248,N_2879);
nand U3731 (N_3731,N_2640,N_2543);
nor U3732 (N_3732,N_2755,N_2501);
and U3733 (N_3733,N_2243,N_2873);
or U3734 (N_3734,N_2992,N_2580);
nor U3735 (N_3735,N_2509,N_2132);
or U3736 (N_3736,N_2237,N_2966);
nand U3737 (N_3737,N_2647,N_2511);
nand U3738 (N_3738,N_2471,N_2167);
nand U3739 (N_3739,N_2979,N_2506);
and U3740 (N_3740,N_2124,N_2114);
or U3741 (N_3741,N_2679,N_2100);
and U3742 (N_3742,N_2063,N_2791);
nand U3743 (N_3743,N_2782,N_2697);
and U3744 (N_3744,N_2526,N_2577);
nand U3745 (N_3745,N_2175,N_2115);
nand U3746 (N_3746,N_2951,N_2736);
xnor U3747 (N_3747,N_2501,N_2252);
nand U3748 (N_3748,N_2276,N_2881);
nor U3749 (N_3749,N_2975,N_2880);
xnor U3750 (N_3750,N_2149,N_2530);
nand U3751 (N_3751,N_2946,N_2508);
nor U3752 (N_3752,N_2670,N_2611);
nand U3753 (N_3753,N_2172,N_2766);
nor U3754 (N_3754,N_2732,N_2229);
or U3755 (N_3755,N_2706,N_2717);
nand U3756 (N_3756,N_2211,N_2389);
and U3757 (N_3757,N_2586,N_2299);
and U3758 (N_3758,N_2607,N_2229);
nand U3759 (N_3759,N_2716,N_2082);
and U3760 (N_3760,N_2979,N_2560);
nor U3761 (N_3761,N_2227,N_2488);
and U3762 (N_3762,N_2838,N_2403);
or U3763 (N_3763,N_2889,N_2055);
nand U3764 (N_3764,N_2479,N_2321);
or U3765 (N_3765,N_2283,N_2202);
nand U3766 (N_3766,N_2360,N_2006);
or U3767 (N_3767,N_2888,N_2780);
nand U3768 (N_3768,N_2368,N_2883);
nand U3769 (N_3769,N_2964,N_2392);
nor U3770 (N_3770,N_2957,N_2519);
nand U3771 (N_3771,N_2937,N_2833);
nand U3772 (N_3772,N_2003,N_2784);
and U3773 (N_3773,N_2591,N_2764);
nor U3774 (N_3774,N_2787,N_2587);
nand U3775 (N_3775,N_2719,N_2200);
or U3776 (N_3776,N_2035,N_2100);
nor U3777 (N_3777,N_2789,N_2222);
nand U3778 (N_3778,N_2089,N_2246);
nor U3779 (N_3779,N_2511,N_2121);
nand U3780 (N_3780,N_2108,N_2031);
or U3781 (N_3781,N_2727,N_2239);
and U3782 (N_3782,N_2353,N_2626);
nand U3783 (N_3783,N_2159,N_2933);
nor U3784 (N_3784,N_2316,N_2318);
or U3785 (N_3785,N_2702,N_2412);
or U3786 (N_3786,N_2245,N_2766);
nand U3787 (N_3787,N_2546,N_2449);
and U3788 (N_3788,N_2324,N_2676);
or U3789 (N_3789,N_2600,N_2638);
xor U3790 (N_3790,N_2604,N_2181);
or U3791 (N_3791,N_2312,N_2980);
or U3792 (N_3792,N_2322,N_2449);
or U3793 (N_3793,N_2944,N_2869);
xnor U3794 (N_3794,N_2171,N_2784);
and U3795 (N_3795,N_2186,N_2310);
nand U3796 (N_3796,N_2444,N_2847);
xor U3797 (N_3797,N_2007,N_2386);
nor U3798 (N_3798,N_2789,N_2357);
nand U3799 (N_3799,N_2586,N_2363);
nor U3800 (N_3800,N_2814,N_2096);
nor U3801 (N_3801,N_2000,N_2403);
nand U3802 (N_3802,N_2080,N_2208);
or U3803 (N_3803,N_2958,N_2763);
or U3804 (N_3804,N_2726,N_2453);
or U3805 (N_3805,N_2773,N_2320);
and U3806 (N_3806,N_2465,N_2689);
nand U3807 (N_3807,N_2128,N_2438);
xor U3808 (N_3808,N_2843,N_2682);
nor U3809 (N_3809,N_2847,N_2165);
xnor U3810 (N_3810,N_2341,N_2067);
nor U3811 (N_3811,N_2521,N_2732);
nor U3812 (N_3812,N_2639,N_2910);
nor U3813 (N_3813,N_2692,N_2126);
or U3814 (N_3814,N_2508,N_2273);
nand U3815 (N_3815,N_2109,N_2621);
or U3816 (N_3816,N_2507,N_2609);
nor U3817 (N_3817,N_2746,N_2710);
and U3818 (N_3818,N_2772,N_2505);
and U3819 (N_3819,N_2199,N_2471);
xor U3820 (N_3820,N_2855,N_2844);
nor U3821 (N_3821,N_2341,N_2245);
and U3822 (N_3822,N_2265,N_2066);
xnor U3823 (N_3823,N_2378,N_2669);
nor U3824 (N_3824,N_2602,N_2390);
nor U3825 (N_3825,N_2526,N_2485);
xor U3826 (N_3826,N_2162,N_2066);
and U3827 (N_3827,N_2527,N_2917);
or U3828 (N_3828,N_2190,N_2213);
and U3829 (N_3829,N_2253,N_2726);
and U3830 (N_3830,N_2430,N_2643);
and U3831 (N_3831,N_2255,N_2830);
nand U3832 (N_3832,N_2690,N_2042);
nand U3833 (N_3833,N_2211,N_2819);
nor U3834 (N_3834,N_2669,N_2483);
nand U3835 (N_3835,N_2416,N_2926);
nand U3836 (N_3836,N_2820,N_2059);
or U3837 (N_3837,N_2779,N_2740);
nand U3838 (N_3838,N_2533,N_2392);
xor U3839 (N_3839,N_2566,N_2790);
nand U3840 (N_3840,N_2293,N_2324);
and U3841 (N_3841,N_2193,N_2507);
nand U3842 (N_3842,N_2000,N_2802);
xnor U3843 (N_3843,N_2504,N_2437);
xor U3844 (N_3844,N_2219,N_2892);
nor U3845 (N_3845,N_2142,N_2218);
and U3846 (N_3846,N_2320,N_2821);
nor U3847 (N_3847,N_2402,N_2150);
nor U3848 (N_3848,N_2904,N_2300);
nand U3849 (N_3849,N_2656,N_2559);
or U3850 (N_3850,N_2758,N_2161);
nand U3851 (N_3851,N_2624,N_2189);
and U3852 (N_3852,N_2565,N_2173);
and U3853 (N_3853,N_2693,N_2139);
and U3854 (N_3854,N_2335,N_2782);
xnor U3855 (N_3855,N_2886,N_2811);
nor U3856 (N_3856,N_2173,N_2992);
and U3857 (N_3857,N_2011,N_2197);
nor U3858 (N_3858,N_2686,N_2194);
and U3859 (N_3859,N_2930,N_2025);
or U3860 (N_3860,N_2448,N_2814);
nor U3861 (N_3861,N_2998,N_2033);
xor U3862 (N_3862,N_2710,N_2028);
nand U3863 (N_3863,N_2519,N_2740);
and U3864 (N_3864,N_2852,N_2542);
or U3865 (N_3865,N_2250,N_2181);
and U3866 (N_3866,N_2669,N_2257);
nor U3867 (N_3867,N_2188,N_2087);
nor U3868 (N_3868,N_2259,N_2276);
nor U3869 (N_3869,N_2356,N_2039);
or U3870 (N_3870,N_2258,N_2798);
nand U3871 (N_3871,N_2458,N_2676);
and U3872 (N_3872,N_2099,N_2787);
or U3873 (N_3873,N_2325,N_2391);
and U3874 (N_3874,N_2612,N_2171);
and U3875 (N_3875,N_2691,N_2269);
or U3876 (N_3876,N_2478,N_2222);
nand U3877 (N_3877,N_2852,N_2428);
or U3878 (N_3878,N_2291,N_2864);
nor U3879 (N_3879,N_2731,N_2657);
and U3880 (N_3880,N_2918,N_2460);
nor U3881 (N_3881,N_2866,N_2581);
nor U3882 (N_3882,N_2033,N_2676);
xor U3883 (N_3883,N_2425,N_2144);
xor U3884 (N_3884,N_2606,N_2057);
or U3885 (N_3885,N_2485,N_2520);
xor U3886 (N_3886,N_2983,N_2131);
nand U3887 (N_3887,N_2617,N_2421);
nand U3888 (N_3888,N_2297,N_2194);
xor U3889 (N_3889,N_2793,N_2995);
nand U3890 (N_3890,N_2250,N_2399);
nand U3891 (N_3891,N_2521,N_2150);
or U3892 (N_3892,N_2124,N_2960);
xnor U3893 (N_3893,N_2614,N_2681);
nand U3894 (N_3894,N_2281,N_2732);
or U3895 (N_3895,N_2867,N_2468);
nor U3896 (N_3896,N_2786,N_2852);
or U3897 (N_3897,N_2178,N_2109);
nor U3898 (N_3898,N_2538,N_2879);
and U3899 (N_3899,N_2841,N_2815);
and U3900 (N_3900,N_2320,N_2113);
and U3901 (N_3901,N_2719,N_2482);
or U3902 (N_3902,N_2067,N_2991);
nand U3903 (N_3903,N_2364,N_2690);
nor U3904 (N_3904,N_2130,N_2154);
and U3905 (N_3905,N_2519,N_2070);
nand U3906 (N_3906,N_2305,N_2564);
xnor U3907 (N_3907,N_2367,N_2539);
nor U3908 (N_3908,N_2840,N_2522);
and U3909 (N_3909,N_2770,N_2073);
and U3910 (N_3910,N_2359,N_2757);
or U3911 (N_3911,N_2047,N_2768);
or U3912 (N_3912,N_2337,N_2442);
xor U3913 (N_3913,N_2005,N_2797);
and U3914 (N_3914,N_2078,N_2591);
or U3915 (N_3915,N_2216,N_2553);
nand U3916 (N_3916,N_2984,N_2151);
nand U3917 (N_3917,N_2453,N_2442);
nor U3918 (N_3918,N_2675,N_2597);
nand U3919 (N_3919,N_2748,N_2039);
xnor U3920 (N_3920,N_2857,N_2028);
or U3921 (N_3921,N_2042,N_2927);
xor U3922 (N_3922,N_2231,N_2256);
or U3923 (N_3923,N_2896,N_2318);
or U3924 (N_3924,N_2667,N_2908);
nand U3925 (N_3925,N_2231,N_2398);
nor U3926 (N_3926,N_2150,N_2954);
and U3927 (N_3927,N_2800,N_2680);
or U3928 (N_3928,N_2616,N_2292);
or U3929 (N_3929,N_2808,N_2067);
nand U3930 (N_3930,N_2931,N_2580);
and U3931 (N_3931,N_2186,N_2527);
xnor U3932 (N_3932,N_2590,N_2093);
and U3933 (N_3933,N_2486,N_2389);
or U3934 (N_3934,N_2881,N_2973);
nand U3935 (N_3935,N_2409,N_2142);
or U3936 (N_3936,N_2051,N_2852);
or U3937 (N_3937,N_2221,N_2325);
and U3938 (N_3938,N_2207,N_2683);
nor U3939 (N_3939,N_2840,N_2844);
nor U3940 (N_3940,N_2740,N_2165);
nand U3941 (N_3941,N_2235,N_2057);
or U3942 (N_3942,N_2785,N_2030);
or U3943 (N_3943,N_2089,N_2159);
nand U3944 (N_3944,N_2242,N_2762);
or U3945 (N_3945,N_2293,N_2419);
xnor U3946 (N_3946,N_2239,N_2832);
and U3947 (N_3947,N_2001,N_2045);
or U3948 (N_3948,N_2100,N_2680);
nor U3949 (N_3949,N_2565,N_2275);
nand U3950 (N_3950,N_2142,N_2499);
and U3951 (N_3951,N_2100,N_2286);
and U3952 (N_3952,N_2713,N_2499);
or U3953 (N_3953,N_2528,N_2356);
or U3954 (N_3954,N_2805,N_2122);
and U3955 (N_3955,N_2374,N_2447);
or U3956 (N_3956,N_2590,N_2859);
or U3957 (N_3957,N_2957,N_2140);
nand U3958 (N_3958,N_2706,N_2864);
and U3959 (N_3959,N_2983,N_2679);
nor U3960 (N_3960,N_2946,N_2858);
or U3961 (N_3961,N_2539,N_2576);
and U3962 (N_3962,N_2882,N_2979);
and U3963 (N_3963,N_2092,N_2159);
or U3964 (N_3964,N_2450,N_2749);
nand U3965 (N_3965,N_2796,N_2776);
or U3966 (N_3966,N_2176,N_2677);
xor U3967 (N_3967,N_2073,N_2378);
nor U3968 (N_3968,N_2974,N_2709);
or U3969 (N_3969,N_2675,N_2520);
nor U3970 (N_3970,N_2066,N_2680);
and U3971 (N_3971,N_2554,N_2792);
or U3972 (N_3972,N_2718,N_2042);
and U3973 (N_3973,N_2399,N_2484);
nand U3974 (N_3974,N_2454,N_2441);
nand U3975 (N_3975,N_2282,N_2661);
nand U3976 (N_3976,N_2461,N_2693);
and U3977 (N_3977,N_2363,N_2016);
nor U3978 (N_3978,N_2310,N_2798);
and U3979 (N_3979,N_2109,N_2292);
xor U3980 (N_3980,N_2932,N_2946);
or U3981 (N_3981,N_2517,N_2354);
and U3982 (N_3982,N_2239,N_2836);
and U3983 (N_3983,N_2639,N_2320);
nor U3984 (N_3984,N_2938,N_2206);
nor U3985 (N_3985,N_2476,N_2572);
nand U3986 (N_3986,N_2124,N_2362);
nor U3987 (N_3987,N_2363,N_2180);
xor U3988 (N_3988,N_2684,N_2979);
and U3989 (N_3989,N_2742,N_2945);
xor U3990 (N_3990,N_2919,N_2511);
nand U3991 (N_3991,N_2092,N_2824);
or U3992 (N_3992,N_2800,N_2694);
nand U3993 (N_3993,N_2684,N_2282);
nand U3994 (N_3994,N_2540,N_2501);
nor U3995 (N_3995,N_2265,N_2562);
nand U3996 (N_3996,N_2806,N_2003);
or U3997 (N_3997,N_2220,N_2536);
and U3998 (N_3998,N_2726,N_2594);
or U3999 (N_3999,N_2268,N_2403);
and U4000 (N_4000,N_3588,N_3669);
nor U4001 (N_4001,N_3036,N_3843);
nand U4002 (N_4002,N_3603,N_3979);
and U4003 (N_4003,N_3319,N_3642);
and U4004 (N_4004,N_3412,N_3228);
nor U4005 (N_4005,N_3810,N_3494);
nor U4006 (N_4006,N_3812,N_3419);
nand U4007 (N_4007,N_3311,N_3636);
and U4008 (N_4008,N_3251,N_3238);
nand U4009 (N_4009,N_3960,N_3671);
or U4010 (N_4010,N_3602,N_3911);
nand U4011 (N_4011,N_3512,N_3284);
nand U4012 (N_4012,N_3692,N_3770);
xnor U4013 (N_4013,N_3594,N_3431);
nand U4014 (N_4014,N_3143,N_3490);
or U4015 (N_4015,N_3520,N_3651);
or U4016 (N_4016,N_3532,N_3461);
or U4017 (N_4017,N_3971,N_3105);
nand U4018 (N_4018,N_3151,N_3368);
nor U4019 (N_4019,N_3179,N_3241);
xor U4020 (N_4020,N_3556,N_3427);
xor U4021 (N_4021,N_3759,N_3043);
nor U4022 (N_4022,N_3069,N_3680);
or U4023 (N_4023,N_3965,N_3548);
or U4024 (N_4024,N_3549,N_3360);
nor U4025 (N_4025,N_3455,N_3046);
or U4026 (N_4026,N_3044,N_3698);
xor U4027 (N_4027,N_3270,N_3689);
nor U4028 (N_4028,N_3744,N_3183);
or U4029 (N_4029,N_3621,N_3060);
nand U4030 (N_4030,N_3531,N_3972);
xnor U4031 (N_4031,N_3868,N_3558);
nor U4032 (N_4032,N_3630,N_3954);
nand U4033 (N_4033,N_3609,N_3479);
nor U4034 (N_4034,N_3087,N_3802);
or U4035 (N_4035,N_3236,N_3795);
and U4036 (N_4036,N_3392,N_3202);
and U4037 (N_4037,N_3216,N_3010);
or U4038 (N_4038,N_3581,N_3233);
nand U4039 (N_4039,N_3535,N_3656);
and U4040 (N_4040,N_3554,N_3413);
nor U4041 (N_4041,N_3130,N_3464);
and U4042 (N_4042,N_3242,N_3645);
and U4043 (N_4043,N_3700,N_3204);
nand U4044 (N_4044,N_3871,N_3415);
and U4045 (N_4045,N_3779,N_3847);
or U4046 (N_4046,N_3154,N_3780);
nor U4047 (N_4047,N_3774,N_3855);
nor U4048 (N_4048,N_3953,N_3369);
nand U4049 (N_4049,N_3090,N_3816);
nor U4050 (N_4050,N_3222,N_3612);
and U4051 (N_4051,N_3343,N_3212);
or U4052 (N_4052,N_3467,N_3113);
nor U4053 (N_4053,N_3463,N_3002);
nor U4054 (N_4054,N_3095,N_3758);
nand U4055 (N_4055,N_3137,N_3207);
nor U4056 (N_4056,N_3437,N_3654);
nand U4057 (N_4057,N_3731,N_3018);
nand U4058 (N_4058,N_3539,N_3796);
nand U4059 (N_4059,N_3966,N_3666);
nand U4060 (N_4060,N_3144,N_3823);
and U4061 (N_4061,N_3356,N_3511);
or U4062 (N_4062,N_3746,N_3434);
xor U4063 (N_4063,N_3540,N_3742);
nor U4064 (N_4064,N_3587,N_3836);
or U4065 (N_4065,N_3443,N_3310);
nor U4066 (N_4066,N_3142,N_3957);
xor U4067 (N_4067,N_3566,N_3178);
or U4068 (N_4068,N_3628,N_3834);
nor U4069 (N_4069,N_3385,N_3777);
and U4070 (N_4070,N_3844,N_3301);
nand U4071 (N_4071,N_3955,N_3472);
nor U4072 (N_4072,N_3266,N_3153);
nand U4073 (N_4073,N_3734,N_3793);
xnor U4074 (N_4074,N_3590,N_3527);
nor U4075 (N_4075,N_3277,N_3752);
nand U4076 (N_4076,N_3889,N_3396);
or U4077 (N_4077,N_3295,N_3918);
nor U4078 (N_4078,N_3003,N_3948);
nand U4079 (N_4079,N_3832,N_3996);
or U4080 (N_4080,N_3004,N_3093);
or U4081 (N_4081,N_3712,N_3167);
or U4082 (N_4082,N_3842,N_3880);
or U4083 (N_4083,N_3023,N_3318);
nand U4084 (N_4084,N_3862,N_3045);
or U4085 (N_4085,N_3940,N_3380);
or U4086 (N_4086,N_3593,N_3345);
and U4087 (N_4087,N_3033,N_3229);
or U4088 (N_4088,N_3405,N_3273);
nor U4089 (N_4089,N_3323,N_3173);
nand U4090 (N_4090,N_3870,N_3987);
nor U4091 (N_4091,N_3975,N_3803);
and U4092 (N_4092,N_3882,N_3097);
nor U4093 (N_4093,N_3613,N_3348);
or U4094 (N_4094,N_3324,N_3243);
or U4095 (N_4095,N_3287,N_3361);
or U4096 (N_4096,N_3353,N_3357);
or U4097 (N_4097,N_3608,N_3509);
nand U4098 (N_4098,N_3622,N_3508);
or U4099 (N_4099,N_3976,N_3504);
or U4100 (N_4100,N_3077,N_3468);
and U4101 (N_4101,N_3120,N_3696);
nor U4102 (N_4102,N_3568,N_3985);
nor U4103 (N_4103,N_3322,N_3344);
xnor U4104 (N_4104,N_3124,N_3007);
nor U4105 (N_4105,N_3248,N_3756);
nand U4106 (N_4106,N_3278,N_3737);
and U4107 (N_4107,N_3833,N_3435);
and U4108 (N_4108,N_3579,N_3571);
nor U4109 (N_4109,N_3271,N_3114);
and U4110 (N_4110,N_3677,N_3340);
and U4111 (N_4111,N_3122,N_3325);
and U4112 (N_4112,N_3668,N_3474);
nand U4113 (N_4113,N_3339,N_3992);
nand U4114 (N_4114,N_3984,N_3279);
or U4115 (N_4115,N_3377,N_3422);
and U4116 (N_4116,N_3252,N_3768);
and U4117 (N_4117,N_3150,N_3533);
and U4118 (N_4118,N_3049,N_3705);
nand U4119 (N_4119,N_3393,N_3063);
and U4120 (N_4120,N_3126,N_3115);
nor U4121 (N_4121,N_3961,N_3051);
nand U4122 (N_4122,N_3619,N_3281);
and U4123 (N_4123,N_3896,N_3838);
or U4124 (N_4124,N_3291,N_3713);
nor U4125 (N_4125,N_3331,N_3061);
or U4126 (N_4126,N_3224,N_3928);
nand U4127 (N_4127,N_3272,N_3168);
nand U4128 (N_4128,N_3264,N_3121);
nor U4129 (N_4129,N_3119,N_3958);
and U4130 (N_4130,N_3190,N_3657);
nor U4131 (N_4131,N_3280,N_3764);
nor U4132 (N_4132,N_3403,N_3687);
nor U4133 (N_4133,N_3521,N_3573);
xnor U4134 (N_4134,N_3038,N_3986);
or U4135 (N_4135,N_3219,N_3553);
nor U4136 (N_4136,N_3232,N_3686);
or U4137 (N_4137,N_3177,N_3606);
xnor U4138 (N_4138,N_3326,N_3840);
nand U4139 (N_4139,N_3788,N_3000);
or U4140 (N_4140,N_3863,N_3516);
nor U4141 (N_4141,N_3306,N_3785);
and U4142 (N_4142,N_3883,N_3854);
and U4143 (N_4143,N_3198,N_3555);
and U4144 (N_4144,N_3626,N_3104);
or U4145 (N_4145,N_3035,N_3635);
nand U4146 (N_4146,N_3931,N_3817);
and U4147 (N_4147,N_3445,N_3933);
or U4148 (N_4148,N_3011,N_3034);
nor U4149 (N_4149,N_3830,N_3110);
or U4150 (N_4150,N_3416,N_3309);
or U4151 (N_4151,N_3522,N_3265);
and U4152 (N_4152,N_3754,N_3818);
nor U4153 (N_4153,N_3483,N_3433);
or U4154 (N_4154,N_3876,N_3864);
or U4155 (N_4155,N_3374,N_3262);
nor U4156 (N_4156,N_3194,N_3086);
nor U4157 (N_4157,N_3544,N_3491);
or U4158 (N_4158,N_3902,N_3952);
and U4159 (N_4159,N_3980,N_3592);
nor U4160 (N_4160,N_3366,N_3096);
nand U4161 (N_4161,N_3787,N_3417);
and U4162 (N_4162,N_3565,N_3223);
nor U4163 (N_4163,N_3254,N_3282);
nor U4164 (N_4164,N_3389,N_3586);
nor U4165 (N_4165,N_3644,N_3302);
xnor U4166 (N_4166,N_3719,N_3714);
nand U4167 (N_4167,N_3359,N_3773);
or U4168 (N_4168,N_3943,N_3446);
or U4169 (N_4169,N_3249,N_3991);
nand U4170 (N_4170,N_3170,N_3199);
nor U4171 (N_4171,N_3017,N_3885);
nor U4172 (N_4172,N_3599,N_3525);
nand U4173 (N_4173,N_3267,N_3798);
or U4174 (N_4174,N_3926,N_3056);
and U4175 (N_4175,N_3459,N_3921);
nand U4176 (N_4176,N_3016,N_3342);
and U4177 (N_4177,N_3808,N_3012);
nand U4178 (N_4178,N_3886,N_3672);
or U4179 (N_4179,N_3849,N_3906);
and U4180 (N_4180,N_3716,N_3998);
nand U4181 (N_4181,N_3074,N_3576);
nand U4182 (N_4182,N_3428,N_3268);
nand U4183 (N_4183,N_3729,N_3505);
or U4184 (N_4184,N_3538,N_3552);
nand U4185 (N_4185,N_3245,N_3103);
and U4186 (N_4186,N_3988,N_3217);
nor U4187 (N_4187,N_3767,N_3032);
or U4188 (N_4188,N_3561,N_3047);
nor U4189 (N_4189,N_3073,N_3037);
or U4190 (N_4190,N_3589,N_3523);
or U4191 (N_4191,N_3425,N_3959);
nand U4192 (N_4192,N_3372,N_3909);
nor U4193 (N_4193,N_3296,N_3230);
xor U4194 (N_4194,N_3418,N_3208);
and U4195 (N_4195,N_3649,N_3676);
and U4196 (N_4196,N_3934,N_3820);
nand U4197 (N_4197,N_3009,N_3977);
and U4198 (N_4198,N_3912,N_3187);
or U4199 (N_4199,N_3949,N_3064);
nand U4200 (N_4200,N_3999,N_3724);
and U4201 (N_4201,N_3888,N_3465);
nand U4202 (N_4202,N_3171,N_3660);
nor U4203 (N_4203,N_3510,N_3691);
nor U4204 (N_4204,N_3730,N_3530);
nand U4205 (N_4205,N_3327,N_3076);
xnor U4206 (N_4206,N_3702,N_3725);
nand U4207 (N_4207,N_3312,N_3085);
nor U4208 (N_4208,N_3182,N_3081);
or U4209 (N_4209,N_3776,N_3653);
and U4210 (N_4210,N_3709,N_3028);
nor U4211 (N_4211,N_3210,N_3543);
or U4212 (N_4212,N_3790,N_3276);
nor U4213 (N_4213,N_3717,N_3867);
nand U4214 (N_4214,N_3292,N_3237);
and U4215 (N_4215,N_3062,N_3457);
nor U4216 (N_4216,N_3815,N_3701);
nor U4217 (N_4217,N_3813,N_3070);
nor U4218 (N_4218,N_3316,N_3710);
xor U4219 (N_4219,N_3444,N_3946);
xor U4220 (N_4220,N_3022,N_3188);
and U4221 (N_4221,N_3584,N_3100);
and U4222 (N_4222,N_3983,N_3735);
or U4223 (N_4223,N_3524,N_3895);
nand U4224 (N_4224,N_3835,N_3797);
or U4225 (N_4225,N_3778,N_3874);
nand U4226 (N_4226,N_3160,N_3694);
or U4227 (N_4227,N_3399,N_3024);
nand U4228 (N_4228,N_3638,N_3400);
nand U4229 (N_4229,N_3355,N_3395);
nand U4230 (N_4230,N_3493,N_3050);
or U4231 (N_4231,N_3424,N_3501);
or U4232 (N_4232,N_3226,N_3439);
or U4233 (N_4233,N_3006,N_3440);
and U4234 (N_4234,N_3580,N_3567);
nor U4235 (N_4235,N_3806,N_3873);
xor U4236 (N_4236,N_3629,N_3495);
nand U4237 (N_4237,N_3745,N_3891);
nor U4238 (N_4238,N_3235,N_3460);
xor U4239 (N_4239,N_3378,N_3469);
nand U4240 (N_4240,N_3286,N_3411);
or U4241 (N_4241,N_3381,N_3487);
and U4242 (N_4242,N_3333,N_3578);
and U4243 (N_4243,N_3106,N_3517);
nand U4244 (N_4244,N_3846,N_3174);
or U4245 (N_4245,N_3658,N_3995);
or U4246 (N_4246,N_3477,N_3244);
nand U4247 (N_4247,N_3211,N_3111);
or U4248 (N_4248,N_3175,N_3614);
or U4249 (N_4249,N_3577,N_3390);
or U4250 (N_4250,N_3901,N_3591);
nand U4251 (N_4251,N_3195,N_3898);
and U4252 (N_4252,N_3781,N_3920);
nor U4253 (N_4253,N_3853,N_3877);
nor U4254 (N_4254,N_3757,N_3157);
nand U4255 (N_4255,N_3547,N_3488);
or U4256 (N_4256,N_3132,N_3409);
xnor U4257 (N_4257,N_3789,N_3486);
nand U4258 (N_4258,N_3337,N_3913);
xor U4259 (N_4259,N_3450,N_3828);
nor U4260 (N_4260,N_3072,N_3969);
or U4261 (N_4261,N_3726,N_3894);
xor U4262 (N_4262,N_3866,N_3117);
or U4263 (N_4263,N_3382,N_3367);
or U4264 (N_4264,N_3401,N_3620);
xor U4265 (N_4265,N_3583,N_3947);
or U4266 (N_4266,N_3447,N_3564);
and U4267 (N_4267,N_3935,N_3181);
nor U4268 (N_4268,N_3763,N_3304);
nor U4269 (N_4269,N_3507,N_3218);
and U4270 (N_4270,N_3082,N_3821);
nor U4271 (N_4271,N_3951,N_3290);
nand U4272 (N_4272,N_3829,N_3938);
nand U4273 (N_4273,N_3346,N_3956);
nor U4274 (N_4274,N_3197,N_3336);
and U4275 (N_4275,N_3970,N_3482);
and U4276 (N_4276,N_3030,N_3088);
and U4277 (N_4277,N_3053,N_3740);
nor U4278 (N_4278,N_3839,N_3640);
nand U4279 (N_4279,N_3155,N_3029);
and U4280 (N_4280,N_3852,N_3632);
nand U4281 (N_4281,N_3080,N_3663);
nor U4282 (N_4282,N_3127,N_3159);
xor U4283 (N_4283,N_3362,N_3827);
or U4284 (N_4284,N_3321,N_3145);
nor U4285 (N_4285,N_3350,N_3600);
or U4286 (N_4286,N_3135,N_3805);
and U4287 (N_4287,N_3376,N_3528);
or U4288 (N_4288,N_3604,N_3068);
nor U4289 (N_4289,N_3247,N_3307);
nor U4290 (N_4290,N_3025,N_3274);
nor U4291 (N_4291,N_3013,N_3426);
nor U4292 (N_4292,N_3430,N_3670);
and U4293 (N_4293,N_3625,N_3231);
or U4294 (N_4294,N_3667,N_3406);
and U4295 (N_4295,N_3518,N_3192);
nand U4296 (N_4296,N_3989,N_3066);
or U4297 (N_4297,N_3536,N_3596);
xnor U4298 (N_4298,N_3263,N_3941);
or U4299 (N_4299,N_3582,N_3749);
or U4300 (N_4300,N_3526,N_3314);
nand U4301 (N_4301,N_3682,N_3020);
nor U4302 (N_4302,N_3647,N_3001);
nand U4303 (N_4303,N_3618,N_3156);
or U4304 (N_4304,N_3545,N_3769);
nand U4305 (N_4305,N_3598,N_3129);
nor U4306 (N_4306,N_3225,N_3476);
and U4307 (N_4307,N_3165,N_3837);
nor U4308 (N_4308,N_3633,N_3929);
or U4309 (N_4309,N_3048,N_3052);
nor U4310 (N_4310,N_3775,N_3610);
or U4311 (N_4311,N_3466,N_3529);
nand U4312 (N_4312,N_3704,N_3220);
or U4313 (N_4313,N_3299,N_3332);
nor U4314 (N_4314,N_3643,N_3101);
nand U4315 (N_4315,N_3615,N_3451);
xor U4316 (N_4316,N_3293,N_3605);
or U4317 (N_4317,N_3240,N_3239);
nor U4318 (N_4318,N_3964,N_3041);
nor U4319 (N_4319,N_3040,N_3695);
nor U4320 (N_4320,N_3027,N_3804);
nand U4321 (N_4321,N_3456,N_3675);
and U4322 (N_4322,N_3711,N_3917);
or U4323 (N_4323,N_3498,N_3075);
nor U4324 (N_4324,N_3897,N_3308);
xnor U4325 (N_4325,N_3485,N_3572);
or U4326 (N_4326,N_3707,N_3910);
nor U4327 (N_4327,N_3283,N_3039);
nand U4328 (N_4328,N_3189,N_3706);
nor U4329 (N_4329,N_3149,N_3685);
and U4330 (N_4330,N_3108,N_3634);
nor U4331 (N_4331,N_3506,N_3213);
nor U4332 (N_4332,N_3963,N_3169);
nand U4333 (N_4333,N_3720,N_3631);
nor U4334 (N_4334,N_3721,N_3936);
or U4335 (N_4335,N_3246,N_3285);
nor U4336 (N_4336,N_3750,N_3761);
and U4337 (N_4337,N_3462,N_3099);
xnor U4338 (N_4338,N_3652,N_3484);
nand U4339 (N_4339,N_3394,N_3923);
and U4340 (N_4340,N_3215,N_3499);
nand U4341 (N_4341,N_3722,N_3848);
nand U4342 (N_4342,N_3858,N_3794);
nand U4343 (N_4343,N_3908,N_3470);
nor U4344 (N_4344,N_3765,N_3193);
nor U4345 (N_4345,N_3743,N_3384);
nor U4346 (N_4346,N_3180,N_3261);
and U4347 (N_4347,N_3221,N_3055);
xnor U4348 (N_4348,N_3162,N_3981);
nand U4349 (N_4349,N_3503,N_3098);
or U4350 (N_4350,N_3831,N_3026);
or U4351 (N_4351,N_3471,N_3397);
or U4352 (N_4352,N_3563,N_3728);
or U4353 (N_4353,N_3015,N_3708);
and U4354 (N_4354,N_3607,N_3442);
nor U4355 (N_4355,N_3365,N_3201);
nor U4356 (N_4356,N_3845,N_3519);
or U4357 (N_4357,N_3341,N_3005);
or U4358 (N_4358,N_3617,N_3347);
nor U4359 (N_4359,N_3650,N_3313);
and U4360 (N_4360,N_3370,N_3305);
nand U4361 (N_4361,N_3407,N_3616);
nor U4362 (N_4362,N_3489,N_3739);
xor U4363 (N_4363,N_3138,N_3927);
or U4364 (N_4364,N_3083,N_3865);
or U4365 (N_4365,N_3388,N_3408);
nor U4366 (N_4366,N_3627,N_3136);
nor U4367 (N_4367,N_3674,N_3480);
nand U4368 (N_4368,N_3298,N_3771);
or U4369 (N_4369,N_3661,N_3693);
nor U4370 (N_4370,N_3534,N_3079);
nor U4371 (N_4371,N_3715,N_3930);
xor U4372 (N_4372,N_3205,N_3328);
nand U4373 (N_4373,N_3665,N_3514);
and U4374 (N_4374,N_3990,N_3684);
nand U4375 (N_4375,N_3574,N_3537);
and U4376 (N_4376,N_3881,N_3560);
and U4377 (N_4377,N_3557,N_3690);
nand U4378 (N_4378,N_3078,N_3067);
nand U4379 (N_4379,N_3732,N_3784);
nor U4380 (N_4380,N_3875,N_3379);
nor U4381 (N_4381,N_3611,N_3914);
or U4382 (N_4382,N_3059,N_3646);
or U4383 (N_4383,N_3297,N_3887);
and U4384 (N_4384,N_3791,N_3163);
nand U4385 (N_4385,N_3227,N_3112);
nor U4386 (N_4386,N_3819,N_3391);
or U4387 (N_4387,N_3751,N_3260);
nand U4388 (N_4388,N_3250,N_3801);
or U4389 (N_4389,N_3166,N_3900);
and U4390 (N_4390,N_3454,N_3057);
and U4391 (N_4391,N_3133,N_3107);
nand U4392 (N_4392,N_3116,N_3747);
or U4393 (N_4393,N_3639,N_3317);
and U4394 (N_4394,N_3659,N_3008);
nand U4395 (N_4395,N_3860,N_3915);
nand U4396 (N_4396,N_3905,N_3448);
or U4397 (N_4397,N_3982,N_3071);
or U4398 (N_4398,N_3497,N_3903);
nor U4399 (N_4399,N_3354,N_3699);
or U4400 (N_4400,N_3973,N_3623);
xnor U4401 (N_4401,N_3209,N_3257);
nor U4402 (N_4402,N_3932,N_3799);
nand U4403 (N_4403,N_3733,N_3423);
nand U4404 (N_4404,N_3783,N_3595);
or U4405 (N_4405,N_3824,N_3939);
xor U4406 (N_4406,N_3678,N_3358);
nand U4407 (N_4407,N_3892,N_3962);
or U4408 (N_4408,N_3158,N_3879);
nor U4409 (N_4409,N_3703,N_3338);
nor U4410 (N_4410,N_3161,N_3924);
or U4411 (N_4411,N_3569,N_3515);
and U4412 (N_4412,N_3475,N_3502);
nor U4413 (N_4413,N_3432,N_3125);
and U4414 (N_4414,N_3420,N_3562);
nor U4415 (N_4415,N_3942,N_3184);
or U4416 (N_4416,N_3131,N_3019);
or U4417 (N_4417,N_3429,N_3139);
nor U4418 (N_4418,N_3058,N_3258);
nand U4419 (N_4419,N_3859,N_3772);
or U4420 (N_4420,N_3031,N_3937);
and U4421 (N_4421,N_3861,N_3089);
nand U4422 (N_4422,N_3500,N_3320);
nor U4423 (N_4423,N_3513,N_3148);
nand U4424 (N_4424,N_3092,N_3481);
or U4425 (N_4425,N_3597,N_3869);
nor U4426 (N_4426,N_3727,N_3123);
xnor U4427 (N_4427,N_3206,N_3748);
nor U4428 (N_4428,N_3185,N_3807);
nand U4429 (N_4429,N_3496,N_3054);
or U4430 (N_4430,N_3414,N_3792);
and U4431 (N_4431,N_3575,N_3662);
nor U4432 (N_4432,N_3814,N_3335);
nor U4433 (N_4433,N_3559,N_3851);
or U4434 (N_4434,N_3825,N_3681);
nand U4435 (N_4435,N_3164,N_3351);
nand U4436 (N_4436,N_3919,N_3809);
nor U4437 (N_4437,N_3315,N_3303);
or U4438 (N_4438,N_3762,N_3492);
or U4439 (N_4439,N_3893,N_3449);
nand U4440 (N_4440,N_3176,N_3857);
and U4441 (N_4441,N_3200,N_3550);
and U4442 (N_4442,N_3822,N_3925);
nand U4443 (N_4443,N_3383,N_3782);
nand U4444 (N_4444,N_3850,N_3736);
and U4445 (N_4445,N_3436,N_3766);
nor U4446 (N_4446,N_3551,N_3330);
nand U4447 (N_4447,N_3118,N_3196);
nand U4448 (N_4448,N_3259,N_3253);
and U4449 (N_4449,N_3841,N_3453);
or U4450 (N_4450,N_3473,N_3140);
or U4451 (N_4451,N_3452,N_3234);
or U4452 (N_4452,N_3546,N_3723);
nand U4453 (N_4453,N_3997,N_3373);
nor U4454 (N_4454,N_3300,N_3826);
nor U4455 (N_4455,N_3585,N_3288);
nand U4456 (N_4456,N_3760,N_3146);
nor U4457 (N_4457,N_3974,N_3994);
nand U4458 (N_4458,N_3065,N_3856);
and U4459 (N_4459,N_3375,N_3128);
or U4460 (N_4460,N_3094,N_3289);
nand U4461 (N_4461,N_3683,N_3441);
nor U4462 (N_4462,N_3329,N_3648);
and U4463 (N_4463,N_3697,N_3978);
nor U4464 (N_4464,N_3152,N_3042);
nor U4465 (N_4465,N_3458,N_3398);
nor U4466 (N_4466,N_3404,N_3014);
nand U4467 (N_4467,N_3641,N_3084);
xor U4468 (N_4468,N_3738,N_3624);
or U4469 (N_4469,N_3109,N_3944);
nand U4470 (N_4470,N_3371,N_3945);
nor U4471 (N_4471,N_3410,N_3386);
and U4472 (N_4472,N_3601,N_3172);
nand U4473 (N_4473,N_3664,N_3275);
nor U4474 (N_4474,N_3688,N_3203);
or U4475 (N_4475,N_3968,N_3679);
nor U4476 (N_4476,N_3890,N_3542);
or U4477 (N_4477,N_3147,N_3387);
and U4478 (N_4478,N_3021,N_3967);
or U4479 (N_4479,N_3334,N_3541);
nor U4480 (N_4480,N_3294,N_3907);
or U4481 (N_4481,N_3904,N_3363);
nor U4482 (N_4482,N_3878,N_3673);
and U4483 (N_4483,N_3256,N_3352);
nand U4484 (N_4484,N_3800,N_3872);
or U4485 (N_4485,N_3478,N_3186);
nor U4486 (N_4486,N_3884,N_3091);
and U4487 (N_4487,N_3811,N_3655);
nand U4488 (N_4488,N_3141,N_3364);
or U4489 (N_4489,N_3349,N_3922);
and U4490 (N_4490,N_3637,N_3993);
or U4491 (N_4491,N_3741,N_3755);
and U4492 (N_4492,N_3191,N_3421);
nand U4493 (N_4493,N_3916,N_3570);
nand U4494 (N_4494,N_3786,N_3134);
nor U4495 (N_4495,N_3102,N_3899);
nand U4496 (N_4496,N_3950,N_3402);
xnor U4497 (N_4497,N_3718,N_3438);
or U4498 (N_4498,N_3214,N_3269);
and U4499 (N_4499,N_3255,N_3753);
and U4500 (N_4500,N_3324,N_3907);
xnor U4501 (N_4501,N_3612,N_3225);
or U4502 (N_4502,N_3573,N_3158);
xor U4503 (N_4503,N_3431,N_3104);
xor U4504 (N_4504,N_3821,N_3627);
nand U4505 (N_4505,N_3982,N_3155);
and U4506 (N_4506,N_3490,N_3697);
or U4507 (N_4507,N_3792,N_3612);
and U4508 (N_4508,N_3959,N_3253);
nor U4509 (N_4509,N_3312,N_3341);
or U4510 (N_4510,N_3052,N_3879);
nor U4511 (N_4511,N_3686,N_3272);
nand U4512 (N_4512,N_3778,N_3418);
and U4513 (N_4513,N_3301,N_3365);
nand U4514 (N_4514,N_3438,N_3563);
xor U4515 (N_4515,N_3545,N_3637);
or U4516 (N_4516,N_3531,N_3994);
nand U4517 (N_4517,N_3899,N_3046);
and U4518 (N_4518,N_3768,N_3948);
xnor U4519 (N_4519,N_3135,N_3767);
nand U4520 (N_4520,N_3590,N_3320);
nor U4521 (N_4521,N_3640,N_3371);
and U4522 (N_4522,N_3269,N_3677);
or U4523 (N_4523,N_3115,N_3223);
nor U4524 (N_4524,N_3041,N_3596);
nand U4525 (N_4525,N_3873,N_3012);
and U4526 (N_4526,N_3090,N_3606);
xnor U4527 (N_4527,N_3754,N_3077);
xor U4528 (N_4528,N_3616,N_3689);
nand U4529 (N_4529,N_3629,N_3772);
and U4530 (N_4530,N_3721,N_3885);
or U4531 (N_4531,N_3070,N_3005);
nand U4532 (N_4532,N_3784,N_3052);
nor U4533 (N_4533,N_3659,N_3748);
or U4534 (N_4534,N_3774,N_3537);
and U4535 (N_4535,N_3776,N_3961);
or U4536 (N_4536,N_3532,N_3696);
nand U4537 (N_4537,N_3617,N_3233);
and U4538 (N_4538,N_3676,N_3399);
or U4539 (N_4539,N_3155,N_3110);
nand U4540 (N_4540,N_3548,N_3545);
and U4541 (N_4541,N_3405,N_3999);
xnor U4542 (N_4542,N_3830,N_3422);
nor U4543 (N_4543,N_3358,N_3472);
nor U4544 (N_4544,N_3347,N_3351);
nor U4545 (N_4545,N_3776,N_3266);
nand U4546 (N_4546,N_3735,N_3627);
xor U4547 (N_4547,N_3486,N_3646);
nand U4548 (N_4548,N_3796,N_3330);
nand U4549 (N_4549,N_3320,N_3520);
and U4550 (N_4550,N_3224,N_3986);
nand U4551 (N_4551,N_3381,N_3646);
nand U4552 (N_4552,N_3503,N_3388);
nand U4553 (N_4553,N_3113,N_3808);
or U4554 (N_4554,N_3787,N_3912);
and U4555 (N_4555,N_3310,N_3901);
and U4556 (N_4556,N_3514,N_3040);
and U4557 (N_4557,N_3077,N_3495);
nor U4558 (N_4558,N_3624,N_3173);
nor U4559 (N_4559,N_3905,N_3478);
nand U4560 (N_4560,N_3521,N_3170);
nor U4561 (N_4561,N_3140,N_3626);
or U4562 (N_4562,N_3573,N_3814);
and U4563 (N_4563,N_3422,N_3192);
nor U4564 (N_4564,N_3314,N_3430);
nor U4565 (N_4565,N_3777,N_3296);
and U4566 (N_4566,N_3635,N_3899);
or U4567 (N_4567,N_3144,N_3814);
or U4568 (N_4568,N_3099,N_3924);
nand U4569 (N_4569,N_3818,N_3520);
nor U4570 (N_4570,N_3558,N_3368);
xnor U4571 (N_4571,N_3781,N_3646);
or U4572 (N_4572,N_3905,N_3067);
or U4573 (N_4573,N_3851,N_3273);
and U4574 (N_4574,N_3436,N_3910);
nand U4575 (N_4575,N_3594,N_3005);
and U4576 (N_4576,N_3058,N_3733);
or U4577 (N_4577,N_3745,N_3541);
xor U4578 (N_4578,N_3879,N_3232);
or U4579 (N_4579,N_3295,N_3581);
nand U4580 (N_4580,N_3162,N_3747);
nor U4581 (N_4581,N_3521,N_3235);
and U4582 (N_4582,N_3468,N_3786);
xor U4583 (N_4583,N_3410,N_3441);
nand U4584 (N_4584,N_3718,N_3196);
and U4585 (N_4585,N_3851,N_3276);
or U4586 (N_4586,N_3709,N_3703);
nand U4587 (N_4587,N_3311,N_3241);
nand U4588 (N_4588,N_3586,N_3147);
xnor U4589 (N_4589,N_3564,N_3190);
and U4590 (N_4590,N_3615,N_3809);
nor U4591 (N_4591,N_3122,N_3979);
and U4592 (N_4592,N_3884,N_3218);
or U4593 (N_4593,N_3618,N_3846);
nand U4594 (N_4594,N_3169,N_3806);
and U4595 (N_4595,N_3504,N_3297);
or U4596 (N_4596,N_3026,N_3467);
and U4597 (N_4597,N_3516,N_3864);
or U4598 (N_4598,N_3082,N_3692);
or U4599 (N_4599,N_3463,N_3924);
and U4600 (N_4600,N_3784,N_3780);
nand U4601 (N_4601,N_3396,N_3649);
and U4602 (N_4602,N_3731,N_3051);
or U4603 (N_4603,N_3951,N_3890);
nor U4604 (N_4604,N_3815,N_3304);
and U4605 (N_4605,N_3609,N_3736);
and U4606 (N_4606,N_3143,N_3001);
nand U4607 (N_4607,N_3387,N_3130);
nand U4608 (N_4608,N_3944,N_3032);
or U4609 (N_4609,N_3219,N_3109);
or U4610 (N_4610,N_3831,N_3705);
and U4611 (N_4611,N_3149,N_3984);
or U4612 (N_4612,N_3976,N_3909);
or U4613 (N_4613,N_3991,N_3597);
nand U4614 (N_4614,N_3676,N_3661);
nand U4615 (N_4615,N_3409,N_3695);
xnor U4616 (N_4616,N_3947,N_3670);
and U4617 (N_4617,N_3904,N_3611);
nor U4618 (N_4618,N_3513,N_3010);
nor U4619 (N_4619,N_3311,N_3839);
nand U4620 (N_4620,N_3709,N_3981);
xnor U4621 (N_4621,N_3460,N_3053);
and U4622 (N_4622,N_3461,N_3466);
nand U4623 (N_4623,N_3793,N_3614);
and U4624 (N_4624,N_3411,N_3551);
nand U4625 (N_4625,N_3973,N_3519);
and U4626 (N_4626,N_3043,N_3990);
and U4627 (N_4627,N_3949,N_3731);
and U4628 (N_4628,N_3053,N_3726);
xor U4629 (N_4629,N_3600,N_3992);
or U4630 (N_4630,N_3570,N_3690);
xnor U4631 (N_4631,N_3539,N_3422);
nand U4632 (N_4632,N_3347,N_3120);
and U4633 (N_4633,N_3678,N_3315);
nand U4634 (N_4634,N_3244,N_3203);
or U4635 (N_4635,N_3370,N_3286);
or U4636 (N_4636,N_3560,N_3462);
nand U4637 (N_4637,N_3545,N_3715);
or U4638 (N_4638,N_3587,N_3222);
nand U4639 (N_4639,N_3915,N_3506);
nor U4640 (N_4640,N_3368,N_3260);
nand U4641 (N_4641,N_3497,N_3631);
nor U4642 (N_4642,N_3730,N_3648);
and U4643 (N_4643,N_3292,N_3221);
xor U4644 (N_4644,N_3619,N_3577);
and U4645 (N_4645,N_3944,N_3970);
nand U4646 (N_4646,N_3378,N_3634);
nor U4647 (N_4647,N_3078,N_3418);
or U4648 (N_4648,N_3255,N_3259);
nand U4649 (N_4649,N_3301,N_3434);
nor U4650 (N_4650,N_3396,N_3357);
nor U4651 (N_4651,N_3916,N_3323);
and U4652 (N_4652,N_3557,N_3649);
and U4653 (N_4653,N_3171,N_3194);
nand U4654 (N_4654,N_3569,N_3945);
and U4655 (N_4655,N_3910,N_3338);
nor U4656 (N_4656,N_3795,N_3345);
nand U4657 (N_4657,N_3462,N_3696);
nand U4658 (N_4658,N_3100,N_3614);
nor U4659 (N_4659,N_3573,N_3535);
nor U4660 (N_4660,N_3816,N_3127);
nor U4661 (N_4661,N_3364,N_3824);
nand U4662 (N_4662,N_3530,N_3398);
and U4663 (N_4663,N_3421,N_3895);
and U4664 (N_4664,N_3901,N_3959);
nor U4665 (N_4665,N_3691,N_3106);
nor U4666 (N_4666,N_3436,N_3150);
nor U4667 (N_4667,N_3616,N_3860);
and U4668 (N_4668,N_3837,N_3240);
and U4669 (N_4669,N_3396,N_3501);
nand U4670 (N_4670,N_3066,N_3929);
nand U4671 (N_4671,N_3614,N_3032);
nand U4672 (N_4672,N_3361,N_3346);
nand U4673 (N_4673,N_3600,N_3825);
nand U4674 (N_4674,N_3899,N_3646);
nand U4675 (N_4675,N_3327,N_3770);
nor U4676 (N_4676,N_3783,N_3876);
nand U4677 (N_4677,N_3984,N_3136);
or U4678 (N_4678,N_3745,N_3801);
nor U4679 (N_4679,N_3703,N_3219);
and U4680 (N_4680,N_3137,N_3215);
nand U4681 (N_4681,N_3969,N_3004);
nand U4682 (N_4682,N_3234,N_3706);
or U4683 (N_4683,N_3369,N_3102);
nand U4684 (N_4684,N_3665,N_3470);
nor U4685 (N_4685,N_3404,N_3207);
nand U4686 (N_4686,N_3584,N_3213);
nand U4687 (N_4687,N_3216,N_3135);
nand U4688 (N_4688,N_3423,N_3622);
and U4689 (N_4689,N_3160,N_3528);
or U4690 (N_4690,N_3304,N_3630);
nor U4691 (N_4691,N_3293,N_3755);
or U4692 (N_4692,N_3096,N_3551);
nor U4693 (N_4693,N_3062,N_3823);
nand U4694 (N_4694,N_3905,N_3599);
and U4695 (N_4695,N_3770,N_3804);
or U4696 (N_4696,N_3904,N_3873);
or U4697 (N_4697,N_3538,N_3177);
or U4698 (N_4698,N_3711,N_3455);
or U4699 (N_4699,N_3808,N_3893);
nor U4700 (N_4700,N_3558,N_3017);
and U4701 (N_4701,N_3999,N_3918);
nand U4702 (N_4702,N_3666,N_3960);
nand U4703 (N_4703,N_3544,N_3786);
nand U4704 (N_4704,N_3516,N_3256);
xor U4705 (N_4705,N_3021,N_3496);
nand U4706 (N_4706,N_3244,N_3638);
or U4707 (N_4707,N_3663,N_3757);
nand U4708 (N_4708,N_3081,N_3801);
nor U4709 (N_4709,N_3791,N_3956);
and U4710 (N_4710,N_3388,N_3809);
or U4711 (N_4711,N_3833,N_3881);
and U4712 (N_4712,N_3335,N_3862);
nor U4713 (N_4713,N_3355,N_3400);
nand U4714 (N_4714,N_3085,N_3170);
nor U4715 (N_4715,N_3562,N_3460);
xor U4716 (N_4716,N_3986,N_3467);
nor U4717 (N_4717,N_3373,N_3060);
nand U4718 (N_4718,N_3535,N_3930);
and U4719 (N_4719,N_3348,N_3989);
nand U4720 (N_4720,N_3727,N_3412);
nand U4721 (N_4721,N_3238,N_3183);
and U4722 (N_4722,N_3612,N_3042);
nor U4723 (N_4723,N_3591,N_3576);
and U4724 (N_4724,N_3805,N_3827);
and U4725 (N_4725,N_3002,N_3389);
nand U4726 (N_4726,N_3985,N_3261);
nand U4727 (N_4727,N_3722,N_3430);
and U4728 (N_4728,N_3481,N_3606);
or U4729 (N_4729,N_3567,N_3041);
and U4730 (N_4730,N_3032,N_3736);
nand U4731 (N_4731,N_3743,N_3257);
xor U4732 (N_4732,N_3592,N_3485);
nand U4733 (N_4733,N_3156,N_3889);
or U4734 (N_4734,N_3479,N_3117);
and U4735 (N_4735,N_3553,N_3878);
nand U4736 (N_4736,N_3764,N_3034);
and U4737 (N_4737,N_3495,N_3364);
nor U4738 (N_4738,N_3571,N_3543);
nor U4739 (N_4739,N_3961,N_3001);
and U4740 (N_4740,N_3345,N_3724);
nor U4741 (N_4741,N_3857,N_3770);
and U4742 (N_4742,N_3437,N_3045);
and U4743 (N_4743,N_3171,N_3775);
and U4744 (N_4744,N_3598,N_3853);
nor U4745 (N_4745,N_3116,N_3355);
and U4746 (N_4746,N_3209,N_3100);
nand U4747 (N_4747,N_3832,N_3675);
and U4748 (N_4748,N_3436,N_3315);
or U4749 (N_4749,N_3466,N_3673);
or U4750 (N_4750,N_3484,N_3656);
and U4751 (N_4751,N_3221,N_3069);
nor U4752 (N_4752,N_3123,N_3591);
or U4753 (N_4753,N_3122,N_3599);
or U4754 (N_4754,N_3588,N_3760);
and U4755 (N_4755,N_3436,N_3172);
or U4756 (N_4756,N_3466,N_3312);
and U4757 (N_4757,N_3115,N_3686);
nand U4758 (N_4758,N_3800,N_3063);
and U4759 (N_4759,N_3119,N_3558);
or U4760 (N_4760,N_3387,N_3481);
xnor U4761 (N_4761,N_3524,N_3801);
and U4762 (N_4762,N_3482,N_3198);
nand U4763 (N_4763,N_3676,N_3196);
nor U4764 (N_4764,N_3032,N_3788);
nand U4765 (N_4765,N_3165,N_3426);
nand U4766 (N_4766,N_3285,N_3578);
and U4767 (N_4767,N_3149,N_3130);
nand U4768 (N_4768,N_3099,N_3911);
and U4769 (N_4769,N_3316,N_3019);
xor U4770 (N_4770,N_3263,N_3827);
or U4771 (N_4771,N_3566,N_3002);
or U4772 (N_4772,N_3784,N_3910);
and U4773 (N_4773,N_3541,N_3402);
and U4774 (N_4774,N_3250,N_3070);
or U4775 (N_4775,N_3601,N_3242);
nor U4776 (N_4776,N_3209,N_3134);
and U4777 (N_4777,N_3928,N_3894);
nand U4778 (N_4778,N_3115,N_3764);
nor U4779 (N_4779,N_3141,N_3157);
nor U4780 (N_4780,N_3466,N_3069);
nor U4781 (N_4781,N_3921,N_3436);
xnor U4782 (N_4782,N_3768,N_3026);
or U4783 (N_4783,N_3755,N_3971);
nor U4784 (N_4784,N_3607,N_3367);
or U4785 (N_4785,N_3382,N_3571);
or U4786 (N_4786,N_3447,N_3838);
and U4787 (N_4787,N_3958,N_3248);
xor U4788 (N_4788,N_3825,N_3570);
and U4789 (N_4789,N_3666,N_3152);
and U4790 (N_4790,N_3941,N_3697);
and U4791 (N_4791,N_3638,N_3769);
or U4792 (N_4792,N_3084,N_3402);
nand U4793 (N_4793,N_3313,N_3592);
and U4794 (N_4794,N_3837,N_3241);
nor U4795 (N_4795,N_3613,N_3325);
and U4796 (N_4796,N_3193,N_3654);
and U4797 (N_4797,N_3988,N_3950);
nand U4798 (N_4798,N_3256,N_3851);
and U4799 (N_4799,N_3622,N_3233);
or U4800 (N_4800,N_3485,N_3934);
xnor U4801 (N_4801,N_3441,N_3080);
nand U4802 (N_4802,N_3953,N_3405);
xor U4803 (N_4803,N_3209,N_3541);
nor U4804 (N_4804,N_3740,N_3425);
nand U4805 (N_4805,N_3596,N_3778);
nand U4806 (N_4806,N_3851,N_3448);
and U4807 (N_4807,N_3246,N_3750);
and U4808 (N_4808,N_3022,N_3317);
and U4809 (N_4809,N_3849,N_3791);
and U4810 (N_4810,N_3342,N_3550);
nand U4811 (N_4811,N_3120,N_3384);
nor U4812 (N_4812,N_3787,N_3719);
nand U4813 (N_4813,N_3598,N_3034);
nand U4814 (N_4814,N_3294,N_3417);
and U4815 (N_4815,N_3101,N_3472);
or U4816 (N_4816,N_3801,N_3064);
or U4817 (N_4817,N_3425,N_3784);
xor U4818 (N_4818,N_3939,N_3013);
nand U4819 (N_4819,N_3502,N_3058);
or U4820 (N_4820,N_3268,N_3278);
or U4821 (N_4821,N_3811,N_3649);
and U4822 (N_4822,N_3020,N_3831);
xor U4823 (N_4823,N_3278,N_3071);
and U4824 (N_4824,N_3501,N_3194);
and U4825 (N_4825,N_3028,N_3568);
xor U4826 (N_4826,N_3744,N_3466);
and U4827 (N_4827,N_3137,N_3079);
nor U4828 (N_4828,N_3381,N_3967);
or U4829 (N_4829,N_3202,N_3366);
and U4830 (N_4830,N_3719,N_3254);
and U4831 (N_4831,N_3533,N_3884);
xor U4832 (N_4832,N_3678,N_3450);
nor U4833 (N_4833,N_3607,N_3311);
nor U4834 (N_4834,N_3441,N_3323);
or U4835 (N_4835,N_3693,N_3912);
nand U4836 (N_4836,N_3251,N_3865);
or U4837 (N_4837,N_3123,N_3089);
and U4838 (N_4838,N_3729,N_3914);
nor U4839 (N_4839,N_3390,N_3334);
and U4840 (N_4840,N_3966,N_3570);
nand U4841 (N_4841,N_3036,N_3253);
and U4842 (N_4842,N_3546,N_3797);
nor U4843 (N_4843,N_3865,N_3319);
and U4844 (N_4844,N_3713,N_3351);
and U4845 (N_4845,N_3621,N_3809);
or U4846 (N_4846,N_3057,N_3073);
or U4847 (N_4847,N_3088,N_3054);
nand U4848 (N_4848,N_3231,N_3332);
nor U4849 (N_4849,N_3057,N_3430);
nand U4850 (N_4850,N_3939,N_3372);
and U4851 (N_4851,N_3827,N_3217);
and U4852 (N_4852,N_3774,N_3016);
nand U4853 (N_4853,N_3894,N_3197);
nor U4854 (N_4854,N_3112,N_3048);
nand U4855 (N_4855,N_3543,N_3421);
nor U4856 (N_4856,N_3222,N_3416);
xnor U4857 (N_4857,N_3961,N_3930);
nand U4858 (N_4858,N_3760,N_3179);
or U4859 (N_4859,N_3494,N_3885);
nor U4860 (N_4860,N_3942,N_3789);
and U4861 (N_4861,N_3932,N_3949);
nand U4862 (N_4862,N_3135,N_3570);
nor U4863 (N_4863,N_3026,N_3182);
nand U4864 (N_4864,N_3805,N_3947);
xnor U4865 (N_4865,N_3073,N_3183);
nor U4866 (N_4866,N_3504,N_3165);
and U4867 (N_4867,N_3725,N_3309);
nor U4868 (N_4868,N_3647,N_3701);
nor U4869 (N_4869,N_3344,N_3801);
nand U4870 (N_4870,N_3747,N_3278);
nand U4871 (N_4871,N_3086,N_3847);
xor U4872 (N_4872,N_3166,N_3639);
nor U4873 (N_4873,N_3295,N_3341);
or U4874 (N_4874,N_3232,N_3630);
nand U4875 (N_4875,N_3405,N_3609);
or U4876 (N_4876,N_3103,N_3596);
or U4877 (N_4877,N_3300,N_3498);
and U4878 (N_4878,N_3888,N_3740);
nor U4879 (N_4879,N_3667,N_3263);
and U4880 (N_4880,N_3165,N_3268);
or U4881 (N_4881,N_3402,N_3210);
nor U4882 (N_4882,N_3694,N_3686);
nand U4883 (N_4883,N_3896,N_3210);
nand U4884 (N_4884,N_3311,N_3456);
and U4885 (N_4885,N_3119,N_3608);
xor U4886 (N_4886,N_3195,N_3988);
nor U4887 (N_4887,N_3842,N_3597);
and U4888 (N_4888,N_3863,N_3976);
nor U4889 (N_4889,N_3212,N_3025);
nor U4890 (N_4890,N_3634,N_3127);
or U4891 (N_4891,N_3119,N_3702);
or U4892 (N_4892,N_3810,N_3567);
or U4893 (N_4893,N_3780,N_3441);
and U4894 (N_4894,N_3608,N_3034);
or U4895 (N_4895,N_3377,N_3941);
or U4896 (N_4896,N_3827,N_3651);
nor U4897 (N_4897,N_3992,N_3010);
and U4898 (N_4898,N_3853,N_3711);
or U4899 (N_4899,N_3023,N_3903);
nor U4900 (N_4900,N_3509,N_3775);
or U4901 (N_4901,N_3783,N_3281);
nand U4902 (N_4902,N_3024,N_3837);
and U4903 (N_4903,N_3480,N_3591);
nor U4904 (N_4904,N_3715,N_3195);
or U4905 (N_4905,N_3143,N_3761);
nor U4906 (N_4906,N_3720,N_3288);
and U4907 (N_4907,N_3902,N_3544);
nand U4908 (N_4908,N_3788,N_3897);
nor U4909 (N_4909,N_3245,N_3822);
nand U4910 (N_4910,N_3919,N_3231);
nor U4911 (N_4911,N_3990,N_3222);
and U4912 (N_4912,N_3676,N_3698);
nor U4913 (N_4913,N_3149,N_3586);
nor U4914 (N_4914,N_3364,N_3660);
nor U4915 (N_4915,N_3353,N_3675);
nand U4916 (N_4916,N_3207,N_3114);
nor U4917 (N_4917,N_3615,N_3704);
or U4918 (N_4918,N_3253,N_3362);
and U4919 (N_4919,N_3698,N_3532);
nand U4920 (N_4920,N_3654,N_3243);
nor U4921 (N_4921,N_3787,N_3304);
nor U4922 (N_4922,N_3400,N_3569);
nor U4923 (N_4923,N_3199,N_3573);
nor U4924 (N_4924,N_3675,N_3395);
xor U4925 (N_4925,N_3896,N_3371);
nand U4926 (N_4926,N_3763,N_3699);
nand U4927 (N_4927,N_3555,N_3508);
or U4928 (N_4928,N_3416,N_3231);
and U4929 (N_4929,N_3613,N_3957);
and U4930 (N_4930,N_3684,N_3433);
and U4931 (N_4931,N_3143,N_3434);
nor U4932 (N_4932,N_3490,N_3664);
xor U4933 (N_4933,N_3726,N_3286);
xor U4934 (N_4934,N_3998,N_3808);
nand U4935 (N_4935,N_3029,N_3483);
or U4936 (N_4936,N_3406,N_3318);
xnor U4937 (N_4937,N_3330,N_3790);
nand U4938 (N_4938,N_3657,N_3129);
or U4939 (N_4939,N_3339,N_3932);
nor U4940 (N_4940,N_3410,N_3835);
nand U4941 (N_4941,N_3286,N_3852);
nor U4942 (N_4942,N_3423,N_3454);
nor U4943 (N_4943,N_3679,N_3919);
or U4944 (N_4944,N_3591,N_3778);
nand U4945 (N_4945,N_3684,N_3082);
or U4946 (N_4946,N_3982,N_3274);
or U4947 (N_4947,N_3249,N_3020);
nand U4948 (N_4948,N_3350,N_3822);
xor U4949 (N_4949,N_3864,N_3958);
and U4950 (N_4950,N_3119,N_3388);
nand U4951 (N_4951,N_3189,N_3646);
and U4952 (N_4952,N_3993,N_3227);
and U4953 (N_4953,N_3308,N_3110);
or U4954 (N_4954,N_3385,N_3693);
nor U4955 (N_4955,N_3011,N_3237);
nand U4956 (N_4956,N_3751,N_3109);
xor U4957 (N_4957,N_3576,N_3192);
and U4958 (N_4958,N_3498,N_3171);
nor U4959 (N_4959,N_3309,N_3127);
and U4960 (N_4960,N_3616,N_3569);
or U4961 (N_4961,N_3704,N_3301);
and U4962 (N_4962,N_3598,N_3462);
and U4963 (N_4963,N_3834,N_3105);
nor U4964 (N_4964,N_3369,N_3636);
nand U4965 (N_4965,N_3650,N_3725);
and U4966 (N_4966,N_3082,N_3567);
and U4967 (N_4967,N_3394,N_3906);
or U4968 (N_4968,N_3845,N_3875);
and U4969 (N_4969,N_3478,N_3356);
nor U4970 (N_4970,N_3768,N_3757);
nor U4971 (N_4971,N_3618,N_3310);
nand U4972 (N_4972,N_3327,N_3120);
nor U4973 (N_4973,N_3452,N_3859);
nand U4974 (N_4974,N_3647,N_3673);
nor U4975 (N_4975,N_3941,N_3089);
or U4976 (N_4976,N_3908,N_3389);
or U4977 (N_4977,N_3922,N_3632);
xor U4978 (N_4978,N_3396,N_3201);
or U4979 (N_4979,N_3408,N_3416);
xor U4980 (N_4980,N_3907,N_3928);
and U4981 (N_4981,N_3490,N_3480);
or U4982 (N_4982,N_3301,N_3284);
nand U4983 (N_4983,N_3561,N_3036);
xor U4984 (N_4984,N_3226,N_3904);
and U4985 (N_4985,N_3554,N_3456);
or U4986 (N_4986,N_3790,N_3211);
nand U4987 (N_4987,N_3452,N_3706);
nor U4988 (N_4988,N_3011,N_3570);
xnor U4989 (N_4989,N_3526,N_3527);
nand U4990 (N_4990,N_3044,N_3246);
nand U4991 (N_4991,N_3733,N_3623);
or U4992 (N_4992,N_3689,N_3979);
or U4993 (N_4993,N_3541,N_3937);
nor U4994 (N_4994,N_3121,N_3899);
nor U4995 (N_4995,N_3297,N_3576);
nand U4996 (N_4996,N_3973,N_3075);
and U4997 (N_4997,N_3217,N_3186);
nor U4998 (N_4998,N_3293,N_3353);
and U4999 (N_4999,N_3256,N_3279);
and UO_0 (O_0,N_4431,N_4775);
nand UO_1 (O_1,N_4769,N_4170);
xor UO_2 (O_2,N_4210,N_4260);
and UO_3 (O_3,N_4747,N_4103);
or UO_4 (O_4,N_4726,N_4911);
and UO_5 (O_5,N_4615,N_4494);
nor UO_6 (O_6,N_4645,N_4846);
and UO_7 (O_7,N_4398,N_4995);
xor UO_8 (O_8,N_4045,N_4575);
xnor UO_9 (O_9,N_4887,N_4857);
xor UO_10 (O_10,N_4930,N_4740);
nor UO_11 (O_11,N_4607,N_4734);
or UO_12 (O_12,N_4416,N_4519);
and UO_13 (O_13,N_4858,N_4498);
nor UO_14 (O_14,N_4327,N_4359);
nand UO_15 (O_15,N_4903,N_4097);
nand UO_16 (O_16,N_4397,N_4859);
nor UO_17 (O_17,N_4298,N_4776);
or UO_18 (O_18,N_4446,N_4670);
xor UO_19 (O_19,N_4383,N_4493);
or UO_20 (O_20,N_4000,N_4815);
and UO_21 (O_21,N_4269,N_4014);
or UO_22 (O_22,N_4121,N_4888);
or UO_23 (O_23,N_4410,N_4104);
or UO_24 (O_24,N_4276,N_4419);
nand UO_25 (O_25,N_4457,N_4074);
or UO_26 (O_26,N_4291,N_4990);
nand UO_27 (O_27,N_4186,N_4301);
or UO_28 (O_28,N_4316,N_4277);
or UO_29 (O_29,N_4056,N_4566);
xor UO_30 (O_30,N_4009,N_4418);
nand UO_31 (O_31,N_4439,N_4490);
and UO_32 (O_32,N_4019,N_4790);
xor UO_33 (O_33,N_4484,N_4534);
nand UO_34 (O_34,N_4515,N_4626);
and UO_35 (O_35,N_4060,N_4263);
and UO_36 (O_36,N_4375,N_4025);
nor UO_37 (O_37,N_4448,N_4785);
nand UO_38 (O_38,N_4989,N_4317);
xor UO_39 (O_39,N_4255,N_4117);
and UO_40 (O_40,N_4611,N_4133);
or UO_41 (O_41,N_4308,N_4055);
or UO_42 (O_42,N_4706,N_4681);
and UO_43 (O_43,N_4346,N_4666);
nor UO_44 (O_44,N_4052,N_4884);
and UO_45 (O_45,N_4355,N_4279);
or UO_46 (O_46,N_4703,N_4651);
or UO_47 (O_47,N_4042,N_4915);
or UO_48 (O_48,N_4364,N_4078);
nor UO_49 (O_49,N_4798,N_4280);
nor UO_50 (O_50,N_4219,N_4763);
or UO_51 (O_51,N_4605,N_4780);
xnor UO_52 (O_52,N_4131,N_4230);
and UO_53 (O_53,N_4576,N_4046);
and UO_54 (O_54,N_4122,N_4142);
nor UO_55 (O_55,N_4556,N_4179);
and UO_56 (O_56,N_4270,N_4345);
or UO_57 (O_57,N_4167,N_4601);
and UO_58 (O_58,N_4169,N_4433);
or UO_59 (O_59,N_4467,N_4095);
or UO_60 (O_60,N_4223,N_4328);
nor UO_61 (O_61,N_4907,N_4744);
and UO_62 (O_62,N_4402,N_4340);
or UO_63 (O_63,N_4459,N_4671);
nand UO_64 (O_64,N_4486,N_4211);
nand UO_65 (O_65,N_4401,N_4783);
nand UO_66 (O_66,N_4246,N_4509);
or UO_67 (O_67,N_4971,N_4200);
or UO_68 (O_68,N_4144,N_4682);
or UO_69 (O_69,N_4933,N_4109);
or UO_70 (O_70,N_4756,N_4668);
or UO_71 (O_71,N_4113,N_4480);
or UO_72 (O_72,N_4158,N_4898);
nand UO_73 (O_73,N_4384,N_4295);
or UO_74 (O_74,N_4112,N_4156);
nand UO_75 (O_75,N_4172,N_4175);
nor UO_76 (O_76,N_4313,N_4017);
and UO_77 (O_77,N_4202,N_4426);
and UO_78 (O_78,N_4141,N_4176);
and UO_79 (O_79,N_4686,N_4201);
or UO_80 (O_80,N_4228,N_4361);
or UO_81 (O_81,N_4207,N_4595);
xnor UO_82 (O_82,N_4238,N_4466);
nor UO_83 (O_83,N_4960,N_4369);
and UO_84 (O_84,N_4565,N_4733);
or UO_85 (O_85,N_4570,N_4393);
nor UO_86 (O_86,N_4043,N_4928);
or UO_87 (O_87,N_4648,N_4227);
nand UO_88 (O_88,N_4127,N_4979);
nor UO_89 (O_89,N_4525,N_4792);
nand UO_90 (O_90,N_4106,N_4016);
and UO_91 (O_91,N_4994,N_4244);
or UO_92 (O_92,N_4463,N_4126);
and UO_93 (O_93,N_4654,N_4901);
xor UO_94 (O_94,N_4116,N_4386);
and UO_95 (O_95,N_4413,N_4076);
nand UO_96 (O_96,N_4011,N_4587);
nand UO_97 (O_97,N_4717,N_4869);
and UO_98 (O_98,N_4289,N_4378);
nor UO_99 (O_99,N_4661,N_4475);
or UO_100 (O_100,N_4069,N_4006);
xnor UO_101 (O_101,N_4786,N_4900);
or UO_102 (O_102,N_4522,N_4745);
or UO_103 (O_103,N_4603,N_4973);
or UO_104 (O_104,N_4083,N_4759);
nand UO_105 (O_105,N_4927,N_4892);
and UO_106 (O_106,N_4329,N_4412);
nor UO_107 (O_107,N_4941,N_4312);
or UO_108 (O_108,N_4264,N_4497);
or UO_109 (O_109,N_4456,N_4347);
or UO_110 (O_110,N_4921,N_4487);
nand UO_111 (O_111,N_4482,N_4067);
nor UO_112 (O_112,N_4198,N_4975);
nand UO_113 (O_113,N_4986,N_4472);
and UO_114 (O_114,N_4018,N_4988);
nor UO_115 (O_115,N_4580,N_4377);
xor UO_116 (O_116,N_4325,N_4254);
nor UO_117 (O_117,N_4914,N_4504);
nor UO_118 (O_118,N_4394,N_4005);
or UO_119 (O_119,N_4797,N_4796);
and UO_120 (O_120,N_4704,N_4940);
nor UO_121 (O_121,N_4387,N_4677);
or UO_122 (O_122,N_4385,N_4180);
and UO_123 (O_123,N_4166,N_4943);
nand UO_124 (O_124,N_4469,N_4065);
nor UO_125 (O_125,N_4962,N_4080);
nand UO_126 (O_126,N_4920,N_4349);
and UO_127 (O_127,N_4062,N_4068);
nor UO_128 (O_128,N_4008,N_4174);
nor UO_129 (O_129,N_4523,N_4559);
nand UO_130 (O_130,N_4217,N_4602);
and UO_131 (O_131,N_4689,N_4100);
nor UO_132 (O_132,N_4321,N_4022);
nand UO_133 (O_133,N_4157,N_4249);
and UO_134 (O_134,N_4588,N_4058);
xor UO_135 (O_135,N_4360,N_4500);
and UO_136 (O_136,N_4800,N_4718);
and UO_137 (O_137,N_4814,N_4038);
or UO_138 (O_138,N_4878,N_4372);
nor UO_139 (O_139,N_4715,N_4114);
xor UO_140 (O_140,N_4934,N_4627);
or UO_141 (O_141,N_4508,N_4947);
and UO_142 (O_142,N_4512,N_4503);
and UO_143 (O_143,N_4631,N_4030);
nor UO_144 (O_144,N_4477,N_4552);
nand UO_145 (O_145,N_4765,N_4248);
and UO_146 (O_146,N_4963,N_4404);
nor UO_147 (O_147,N_4510,N_4949);
nand UO_148 (O_148,N_4581,N_4791);
or UO_149 (O_149,N_4388,N_4367);
nor UO_150 (O_150,N_4417,N_4481);
nand UO_151 (O_151,N_4855,N_4513);
and UO_152 (O_152,N_4282,N_4558);
xnor UO_153 (O_153,N_4315,N_4243);
nand UO_154 (O_154,N_4337,N_4954);
nor UO_155 (O_155,N_4902,N_4272);
or UO_156 (O_156,N_4091,N_4267);
or UO_157 (O_157,N_4352,N_4048);
or UO_158 (O_158,N_4777,N_4411);
nand UO_159 (O_159,N_4739,N_4425);
or UO_160 (O_160,N_4057,N_4820);
xnor UO_161 (O_161,N_4090,N_4643);
or UO_162 (O_162,N_4698,N_4445);
nand UO_163 (O_163,N_4787,N_4817);
nand UO_164 (O_164,N_4598,N_4320);
and UO_165 (O_165,N_4707,N_4948);
nand UO_166 (O_166,N_4119,N_4281);
xor UO_167 (O_167,N_4444,N_4592);
or UO_168 (O_168,N_4610,N_4098);
xnor UO_169 (O_169,N_4543,N_4978);
nand UO_170 (O_170,N_4001,N_4102);
nor UO_171 (O_171,N_4662,N_4904);
or UO_172 (O_172,N_4604,N_4845);
xor UO_173 (O_173,N_4035,N_4146);
and UO_174 (O_174,N_4816,N_4118);
nand UO_175 (O_175,N_4306,N_4932);
nand UO_176 (O_176,N_4760,N_4899);
xnor UO_177 (O_177,N_4574,N_4140);
and UO_178 (O_178,N_4350,N_4124);
or UO_179 (O_179,N_4597,N_4163);
xnor UO_180 (O_180,N_4297,N_4652);
and UO_181 (O_181,N_4343,N_4222);
xnor UO_182 (O_182,N_4958,N_4415);
and UO_183 (O_183,N_4010,N_4205);
xnor UO_184 (O_184,N_4951,N_4036);
nor UO_185 (O_185,N_4268,N_4518);
or UO_186 (O_186,N_4134,N_4129);
nand UO_187 (O_187,N_4538,N_4633);
nor UO_188 (O_188,N_4086,N_4256);
and UO_189 (O_189,N_4488,N_4299);
nand UO_190 (O_190,N_4409,N_4624);
nor UO_191 (O_191,N_4373,N_4583);
nor UO_192 (O_192,N_4047,N_4586);
nand UO_193 (O_193,N_4547,N_4632);
nor UO_194 (O_194,N_4465,N_4204);
or UO_195 (O_195,N_4096,N_4591);
xnor UO_196 (O_196,N_4980,N_4891);
or UO_197 (O_197,N_4053,N_4403);
nor UO_198 (O_198,N_4961,N_4473);
or UO_199 (O_199,N_4357,N_4309);
nand UO_200 (O_200,N_4985,N_4033);
or UO_201 (O_201,N_4572,N_4724);
or UO_202 (O_202,N_4685,N_4723);
nand UO_203 (O_203,N_4007,N_4694);
and UO_204 (O_204,N_4063,N_4533);
or UO_205 (O_205,N_4619,N_4655);
or UO_206 (O_206,N_4240,N_4614);
nor UO_207 (O_207,N_4746,N_4839);
nand UO_208 (O_208,N_4709,N_4391);
nand UO_209 (O_209,N_4208,N_4041);
nor UO_210 (O_210,N_4753,N_4981);
nor UO_211 (O_211,N_4913,N_4271);
nand UO_212 (O_212,N_4185,N_4319);
xnor UO_213 (O_213,N_4049,N_4969);
nor UO_214 (O_214,N_4752,N_4420);
or UO_215 (O_215,N_4965,N_4236);
xor UO_216 (O_216,N_4061,N_4909);
and UO_217 (O_217,N_4082,N_4189);
nor UO_218 (O_218,N_4827,N_4774);
or UO_219 (O_219,N_4802,N_4916);
nand UO_220 (O_220,N_4294,N_4843);
nand UO_221 (O_221,N_4507,N_4606);
and UO_222 (O_222,N_4532,N_4365);
xor UO_223 (O_223,N_4004,N_4089);
xnor UO_224 (O_224,N_4395,N_4261);
or UO_225 (O_225,N_4535,N_4600);
nand UO_226 (O_226,N_4873,N_4748);
and UO_227 (O_227,N_4665,N_4031);
or UO_228 (O_228,N_4077,N_4883);
nor UO_229 (O_229,N_4324,N_4370);
or UO_230 (O_230,N_4870,N_4612);
and UO_231 (O_231,N_4819,N_4242);
and UO_232 (O_232,N_4101,N_4154);
nor UO_233 (O_233,N_4435,N_4190);
or UO_234 (O_234,N_4865,N_4310);
and UO_235 (O_235,N_4381,N_4303);
and UO_236 (O_236,N_4302,N_4919);
nor UO_237 (O_237,N_4669,N_4620);
and UO_238 (O_238,N_4946,N_4245);
or UO_239 (O_239,N_4613,N_4721);
or UO_240 (O_240,N_4257,N_4695);
xor UO_241 (O_241,N_4164,N_4560);
xor UO_242 (O_242,N_4075,N_4987);
nand UO_243 (O_243,N_4770,N_4646);
nor UO_244 (O_244,N_4524,N_4437);
and UO_245 (O_245,N_4288,N_4897);
and UO_246 (O_246,N_4203,N_4856);
nor UO_247 (O_247,N_4637,N_4339);
nand UO_248 (O_248,N_4521,N_4300);
and UO_249 (O_249,N_4194,N_4374);
or UO_250 (O_250,N_4054,N_4561);
or UO_251 (O_251,N_4218,N_4772);
nand UO_252 (O_252,N_4983,N_4768);
nand UO_253 (O_253,N_4697,N_4161);
nor UO_254 (O_254,N_4735,N_4696);
and UO_255 (O_255,N_4640,N_4461);
nor UO_256 (O_256,N_4278,N_4429);
xor UO_257 (O_257,N_4224,N_4801);
or UO_258 (O_258,N_4977,N_4546);
nand UO_259 (O_259,N_4729,N_4550);
nand UO_260 (O_260,N_4766,N_4910);
nor UO_261 (O_261,N_4476,N_4738);
xor UO_262 (O_262,N_4722,N_4483);
or UO_263 (O_263,N_4929,N_4924);
nand UO_264 (O_264,N_4366,N_4471);
xor UO_265 (O_265,N_4656,N_4183);
xor UO_266 (O_266,N_4639,N_4608);
nand UO_267 (O_267,N_4235,N_4823);
nand UO_268 (O_268,N_4599,N_4020);
nor UO_269 (O_269,N_4758,N_4710);
xnor UO_270 (O_270,N_4285,N_4779);
nand UO_271 (O_271,N_4931,N_4489);
or UO_272 (O_272,N_4622,N_4392);
or UO_273 (O_273,N_4192,N_4024);
and UO_274 (O_274,N_4453,N_4092);
nor UO_275 (O_275,N_4545,N_4649);
nand UO_276 (O_276,N_4537,N_4806);
nor UO_277 (O_277,N_4332,N_4214);
nand UO_278 (O_278,N_4807,N_4216);
xnor UO_279 (O_279,N_4209,N_4750);
nor UO_280 (O_280,N_4539,N_4585);
and UO_281 (O_281,N_4432,N_4937);
nor UO_282 (O_282,N_4834,N_4436);
and UO_283 (O_283,N_4451,N_4353);
and UO_284 (O_284,N_4982,N_4809);
or UO_285 (O_285,N_4700,N_4623);
nor UO_286 (O_286,N_4132,N_4452);
nand UO_287 (O_287,N_4757,N_4195);
nor UO_288 (O_288,N_4474,N_4795);
xor UO_289 (O_289,N_4713,N_4749);
and UO_290 (O_290,N_4028,N_4831);
or UO_291 (O_291,N_4778,N_4253);
nand UO_292 (O_292,N_4330,N_4866);
and UO_293 (O_293,N_4885,N_4462);
nand UO_294 (O_294,N_4553,N_4782);
nand UO_295 (O_295,N_4442,N_4344);
xor UO_296 (O_296,N_4356,N_4773);
nor UO_297 (O_297,N_4993,N_4862);
xor UO_298 (O_298,N_4021,N_4896);
or UO_299 (O_299,N_4283,N_4754);
or UO_300 (O_300,N_4673,N_4099);
and UO_301 (O_301,N_4305,N_4318);
nand UO_302 (O_302,N_4781,N_4247);
nand UO_303 (O_303,N_4621,N_4485);
or UO_304 (O_304,N_4151,N_4348);
or UO_305 (O_305,N_4657,N_4527);
or UO_306 (O_306,N_4842,N_4070);
or UO_307 (O_307,N_4771,N_4590);
nand UO_308 (O_308,N_4578,N_4551);
or UO_309 (O_309,N_4712,N_4860);
nand UO_310 (O_310,N_4259,N_4196);
nand UO_311 (O_311,N_4968,N_4678);
and UO_312 (O_312,N_4742,N_4826);
xor UO_313 (O_313,N_4147,N_4991);
or UO_314 (O_314,N_4567,N_4972);
nor UO_315 (O_315,N_4691,N_4821);
and UO_316 (O_316,N_4221,N_4935);
xor UO_317 (O_317,N_4066,N_4225);
nor UO_318 (O_318,N_4322,N_4793);
or UO_319 (O_319,N_4877,N_4634);
nand UO_320 (O_320,N_4362,N_4193);
nand UO_321 (O_321,N_4026,N_4853);
and UO_322 (O_322,N_4531,N_4926);
nand UO_323 (O_323,N_4160,N_4212);
or UO_324 (O_324,N_4514,N_4848);
nand UO_325 (O_325,N_4501,N_4880);
or UO_326 (O_326,N_4864,N_4912);
xnor UO_327 (O_327,N_4159,N_4882);
xor UO_328 (O_328,N_4274,N_4275);
and UO_329 (O_329,N_4861,N_4447);
and UO_330 (O_330,N_4794,N_4844);
and UO_331 (O_331,N_4908,N_4400);
and UO_332 (O_332,N_4148,N_4799);
nand UO_333 (O_333,N_4568,N_4191);
nand UO_334 (O_334,N_4833,N_4818);
nand UO_335 (O_335,N_4761,N_4804);
nor UO_336 (O_336,N_4495,N_4690);
nor UO_337 (O_337,N_4434,N_4414);
and UO_338 (O_338,N_4389,N_4215);
nor UO_339 (O_339,N_4996,N_4479);
nand UO_340 (O_340,N_4582,N_4307);
nand UO_341 (O_341,N_4334,N_4110);
or UO_342 (O_342,N_4732,N_4725);
xor UO_343 (O_343,N_4079,N_4629);
nand UO_344 (O_344,N_4502,N_4239);
or UO_345 (O_345,N_4520,N_4636);
nor UO_346 (O_346,N_4549,N_4813);
or UO_347 (O_347,N_4379,N_4338);
and UO_348 (O_348,N_4563,N_4674);
nor UO_349 (O_349,N_4918,N_4663);
or UO_350 (O_350,N_4784,N_4087);
xor UO_351 (O_351,N_4071,N_4094);
nand UO_352 (O_352,N_4408,N_4331);
and UO_353 (O_353,N_4832,N_4679);
or UO_354 (O_354,N_4177,N_4618);
or UO_355 (O_355,N_4829,N_4311);
and UO_356 (O_356,N_4135,N_4755);
nor UO_357 (O_357,N_4213,N_4491);
or UO_358 (O_358,N_4967,N_4584);
or UO_359 (O_359,N_4326,N_4013);
nand UO_360 (O_360,N_4917,N_4676);
nand UO_361 (O_361,N_4423,N_4764);
nor UO_362 (O_362,N_4455,N_4130);
nand UO_363 (O_363,N_4064,N_4659);
nor UO_364 (O_364,N_4849,N_4950);
and UO_365 (O_365,N_4894,N_4998);
and UO_366 (O_366,N_4788,N_4032);
nand UO_367 (O_367,N_4557,N_4072);
nand UO_368 (O_368,N_4577,N_4617);
nand UO_369 (O_369,N_4959,N_4838);
or UO_370 (O_370,N_4984,N_4737);
nand UO_371 (O_371,N_4241,N_4380);
or UO_372 (O_372,N_4730,N_4736);
and UO_373 (O_373,N_4505,N_4751);
nand UO_374 (O_374,N_4206,N_4296);
xnor UO_375 (O_375,N_4850,N_4037);
nor UO_376 (O_376,N_4139,N_4964);
nor UO_377 (O_377,N_4162,N_4232);
and UO_378 (O_378,N_4081,N_4262);
nand UO_379 (O_379,N_4667,N_4905);
nand UO_380 (O_380,N_4441,N_4182);
nand UO_381 (O_381,N_4231,N_4825);
nand UO_382 (O_382,N_4427,N_4390);
or UO_383 (O_383,N_4234,N_4406);
and UO_384 (O_384,N_4371,N_4233);
and UO_385 (O_385,N_4644,N_4727);
nand UO_386 (O_386,N_4470,N_4555);
xor UO_387 (O_387,N_4810,N_4573);
nor UO_388 (O_388,N_4108,N_4970);
nand UO_389 (O_389,N_4593,N_4692);
or UO_390 (O_390,N_4530,N_4464);
and UO_391 (O_391,N_4939,N_4852);
or UO_392 (O_392,N_4496,N_4675);
nand UO_393 (O_393,N_4625,N_4683);
nand UO_394 (O_394,N_4699,N_4428);
or UO_395 (O_395,N_4863,N_4171);
or UO_396 (O_396,N_4867,N_4803);
xnor UO_397 (O_397,N_4153,N_4088);
or UO_398 (O_398,N_4528,N_4847);
or UO_399 (O_399,N_4711,N_4138);
or UO_400 (O_400,N_4841,N_4424);
and UO_401 (O_401,N_4705,N_4714);
nor UO_402 (O_402,N_4945,N_4105);
nor UO_403 (O_403,N_4579,N_4178);
or UO_404 (O_404,N_4450,N_4630);
nand UO_405 (O_405,N_4516,N_4039);
nand UO_406 (O_406,N_4893,N_4719);
or UO_407 (O_407,N_4716,N_4029);
or UO_408 (O_408,N_4728,N_4889);
or UO_409 (O_409,N_4701,N_4084);
nand UO_410 (O_410,N_4137,N_4944);
or UO_411 (O_411,N_4229,N_4955);
nor UO_412 (O_412,N_4237,N_4376);
nand UO_413 (O_413,N_4672,N_4828);
or UO_414 (O_414,N_4430,N_4854);
nor UO_415 (O_415,N_4073,N_4762);
or UO_416 (O_416,N_4906,N_4890);
and UO_417 (O_417,N_4421,N_4548);
nor UO_418 (O_418,N_4879,N_4368);
nand UO_419 (O_419,N_4155,N_4407);
nor UO_420 (O_420,N_4293,N_4868);
and UO_421 (O_421,N_4454,N_4250);
and UO_422 (O_422,N_4438,N_4059);
and UO_423 (O_423,N_4422,N_4638);
nor UO_424 (O_424,N_4351,N_4128);
nand UO_425 (O_425,N_4149,N_4252);
and UO_426 (O_426,N_4616,N_4107);
and UO_427 (O_427,N_4399,N_4184);
xor UO_428 (O_428,N_4658,N_4187);
and UO_429 (O_429,N_4999,N_4342);
nor UO_430 (O_430,N_4286,N_4554);
nor UO_431 (O_431,N_4875,N_4323);
xnor UO_432 (O_432,N_4596,N_4822);
xnor UO_433 (O_433,N_4688,N_4966);
and UO_434 (O_434,N_4468,N_4922);
or UO_435 (O_435,N_4886,N_4382);
xor UO_436 (O_436,N_4542,N_4478);
xnor UO_437 (O_437,N_4571,N_4440);
nand UO_438 (O_438,N_4143,N_4635);
and UO_439 (O_439,N_4499,N_4023);
and UO_440 (O_440,N_4836,N_4012);
and UO_441 (O_441,N_4647,N_4292);
nand UO_442 (O_442,N_4199,N_4871);
nor UO_443 (O_443,N_4336,N_4152);
and UO_444 (O_444,N_4258,N_4284);
nand UO_445 (O_445,N_4743,N_4526);
and UO_446 (O_446,N_4653,N_4641);
xnor UO_447 (O_447,N_4314,N_4517);
nand UO_448 (O_448,N_4953,N_4974);
nor UO_449 (O_449,N_4173,N_4506);
nand UO_450 (O_450,N_4812,N_4811);
or UO_451 (O_451,N_4789,N_4664);
nor UO_452 (O_452,N_4564,N_4544);
nand UO_453 (O_453,N_4363,N_4492);
nand UO_454 (O_454,N_4895,N_4805);
or UO_455 (O_455,N_4562,N_4015);
or UO_456 (O_456,N_4354,N_4093);
or UO_457 (O_457,N_4541,N_4835);
xor UO_458 (O_458,N_4830,N_4824);
nand UO_459 (O_459,N_4660,N_4226);
nor UO_460 (O_460,N_4511,N_4003);
and UO_461 (O_461,N_4458,N_4304);
nand UO_462 (O_462,N_4872,N_4702);
nand UO_463 (O_463,N_4123,N_4808);
nor UO_464 (O_464,N_4720,N_4290);
or UO_465 (O_465,N_4405,N_4992);
nor UO_466 (O_466,N_4956,N_4027);
and UO_467 (O_467,N_4536,N_4876);
xor UO_468 (O_468,N_4044,N_4684);
or UO_469 (O_469,N_4002,N_4837);
nand UO_470 (O_470,N_4609,N_4168);
and UO_471 (O_471,N_4881,N_4687);
nand UO_472 (O_472,N_4936,N_4396);
or UO_473 (O_473,N_4273,N_4851);
nor UO_474 (O_474,N_4287,N_4111);
and UO_475 (O_475,N_4741,N_4085);
and UO_476 (O_476,N_4220,N_4050);
or UO_477 (O_477,N_4942,N_4874);
or UO_478 (O_478,N_4443,N_4051);
nor UO_479 (O_479,N_4333,N_4976);
or UO_480 (O_480,N_4594,N_4650);
nand UO_481 (O_481,N_4957,N_4449);
and UO_482 (O_482,N_4938,N_4265);
nor UO_483 (O_483,N_4952,N_4569);
nand UO_484 (O_484,N_4136,N_4540);
or UO_485 (O_485,N_4188,N_4145);
nand UO_486 (O_486,N_4589,N_4642);
and UO_487 (O_487,N_4460,N_4150);
nor UO_488 (O_488,N_4731,N_4708);
or UO_489 (O_489,N_4341,N_4628);
xnor UO_490 (O_490,N_4358,N_4529);
or UO_491 (O_491,N_4251,N_4181);
or UO_492 (O_492,N_4997,N_4335);
nand UO_493 (O_493,N_4120,N_4840);
nand UO_494 (O_494,N_4925,N_4266);
or UO_495 (O_495,N_4197,N_4680);
and UO_496 (O_496,N_4115,N_4125);
nor UO_497 (O_497,N_4693,N_4923);
or UO_498 (O_498,N_4034,N_4040);
nand UO_499 (O_499,N_4767,N_4165);
or UO_500 (O_500,N_4220,N_4667);
and UO_501 (O_501,N_4686,N_4345);
xor UO_502 (O_502,N_4009,N_4201);
nor UO_503 (O_503,N_4214,N_4864);
and UO_504 (O_504,N_4894,N_4759);
and UO_505 (O_505,N_4651,N_4975);
nor UO_506 (O_506,N_4698,N_4449);
nor UO_507 (O_507,N_4428,N_4595);
or UO_508 (O_508,N_4364,N_4725);
nor UO_509 (O_509,N_4351,N_4435);
nor UO_510 (O_510,N_4998,N_4797);
and UO_511 (O_511,N_4328,N_4283);
and UO_512 (O_512,N_4329,N_4983);
nand UO_513 (O_513,N_4007,N_4943);
and UO_514 (O_514,N_4411,N_4955);
or UO_515 (O_515,N_4579,N_4369);
nand UO_516 (O_516,N_4952,N_4038);
and UO_517 (O_517,N_4100,N_4822);
and UO_518 (O_518,N_4892,N_4884);
nor UO_519 (O_519,N_4896,N_4461);
or UO_520 (O_520,N_4051,N_4347);
xnor UO_521 (O_521,N_4261,N_4166);
and UO_522 (O_522,N_4877,N_4908);
nand UO_523 (O_523,N_4959,N_4234);
nand UO_524 (O_524,N_4411,N_4653);
nor UO_525 (O_525,N_4506,N_4216);
and UO_526 (O_526,N_4972,N_4201);
nor UO_527 (O_527,N_4762,N_4370);
or UO_528 (O_528,N_4000,N_4778);
or UO_529 (O_529,N_4621,N_4572);
nor UO_530 (O_530,N_4308,N_4205);
nand UO_531 (O_531,N_4739,N_4485);
nand UO_532 (O_532,N_4978,N_4322);
and UO_533 (O_533,N_4867,N_4841);
and UO_534 (O_534,N_4979,N_4552);
nand UO_535 (O_535,N_4267,N_4853);
or UO_536 (O_536,N_4126,N_4211);
nor UO_537 (O_537,N_4950,N_4376);
nor UO_538 (O_538,N_4381,N_4388);
or UO_539 (O_539,N_4430,N_4097);
xor UO_540 (O_540,N_4939,N_4070);
and UO_541 (O_541,N_4207,N_4487);
and UO_542 (O_542,N_4455,N_4242);
or UO_543 (O_543,N_4412,N_4201);
xor UO_544 (O_544,N_4321,N_4230);
nand UO_545 (O_545,N_4256,N_4582);
nor UO_546 (O_546,N_4244,N_4034);
and UO_547 (O_547,N_4631,N_4836);
and UO_548 (O_548,N_4187,N_4925);
nand UO_549 (O_549,N_4953,N_4076);
xnor UO_550 (O_550,N_4681,N_4229);
and UO_551 (O_551,N_4656,N_4936);
nor UO_552 (O_552,N_4575,N_4749);
nor UO_553 (O_553,N_4799,N_4329);
nor UO_554 (O_554,N_4005,N_4086);
nand UO_555 (O_555,N_4681,N_4471);
nor UO_556 (O_556,N_4770,N_4411);
and UO_557 (O_557,N_4448,N_4545);
nor UO_558 (O_558,N_4894,N_4017);
or UO_559 (O_559,N_4758,N_4121);
or UO_560 (O_560,N_4320,N_4063);
or UO_561 (O_561,N_4559,N_4036);
nand UO_562 (O_562,N_4039,N_4703);
and UO_563 (O_563,N_4894,N_4057);
or UO_564 (O_564,N_4134,N_4629);
nand UO_565 (O_565,N_4350,N_4084);
nor UO_566 (O_566,N_4138,N_4099);
or UO_567 (O_567,N_4061,N_4138);
xor UO_568 (O_568,N_4248,N_4621);
nor UO_569 (O_569,N_4694,N_4794);
xnor UO_570 (O_570,N_4557,N_4213);
nor UO_571 (O_571,N_4496,N_4665);
nor UO_572 (O_572,N_4472,N_4988);
and UO_573 (O_573,N_4309,N_4756);
nor UO_574 (O_574,N_4297,N_4648);
or UO_575 (O_575,N_4265,N_4430);
nand UO_576 (O_576,N_4265,N_4905);
or UO_577 (O_577,N_4194,N_4697);
xnor UO_578 (O_578,N_4746,N_4967);
or UO_579 (O_579,N_4284,N_4580);
nor UO_580 (O_580,N_4966,N_4416);
xnor UO_581 (O_581,N_4143,N_4427);
nand UO_582 (O_582,N_4942,N_4221);
or UO_583 (O_583,N_4044,N_4170);
and UO_584 (O_584,N_4222,N_4034);
xor UO_585 (O_585,N_4006,N_4987);
nand UO_586 (O_586,N_4384,N_4668);
and UO_587 (O_587,N_4010,N_4882);
and UO_588 (O_588,N_4657,N_4304);
nand UO_589 (O_589,N_4843,N_4855);
nor UO_590 (O_590,N_4163,N_4871);
nor UO_591 (O_591,N_4473,N_4566);
xor UO_592 (O_592,N_4777,N_4234);
and UO_593 (O_593,N_4457,N_4221);
and UO_594 (O_594,N_4418,N_4592);
nand UO_595 (O_595,N_4086,N_4362);
or UO_596 (O_596,N_4118,N_4970);
nor UO_597 (O_597,N_4880,N_4162);
nor UO_598 (O_598,N_4873,N_4035);
nand UO_599 (O_599,N_4863,N_4085);
nor UO_600 (O_600,N_4673,N_4561);
nand UO_601 (O_601,N_4659,N_4920);
xnor UO_602 (O_602,N_4938,N_4007);
nand UO_603 (O_603,N_4595,N_4509);
or UO_604 (O_604,N_4751,N_4546);
and UO_605 (O_605,N_4417,N_4441);
nor UO_606 (O_606,N_4250,N_4314);
or UO_607 (O_607,N_4894,N_4060);
nand UO_608 (O_608,N_4720,N_4956);
and UO_609 (O_609,N_4412,N_4146);
xor UO_610 (O_610,N_4013,N_4474);
or UO_611 (O_611,N_4771,N_4319);
and UO_612 (O_612,N_4238,N_4318);
nor UO_613 (O_613,N_4158,N_4928);
nor UO_614 (O_614,N_4649,N_4911);
or UO_615 (O_615,N_4226,N_4032);
nand UO_616 (O_616,N_4597,N_4292);
or UO_617 (O_617,N_4700,N_4572);
or UO_618 (O_618,N_4521,N_4133);
nor UO_619 (O_619,N_4261,N_4604);
nand UO_620 (O_620,N_4688,N_4000);
nor UO_621 (O_621,N_4721,N_4383);
and UO_622 (O_622,N_4548,N_4392);
or UO_623 (O_623,N_4300,N_4888);
or UO_624 (O_624,N_4626,N_4096);
nand UO_625 (O_625,N_4120,N_4261);
nor UO_626 (O_626,N_4310,N_4414);
or UO_627 (O_627,N_4560,N_4569);
or UO_628 (O_628,N_4296,N_4699);
and UO_629 (O_629,N_4970,N_4862);
or UO_630 (O_630,N_4489,N_4418);
and UO_631 (O_631,N_4970,N_4947);
or UO_632 (O_632,N_4769,N_4339);
nor UO_633 (O_633,N_4532,N_4815);
nor UO_634 (O_634,N_4260,N_4742);
or UO_635 (O_635,N_4595,N_4240);
nand UO_636 (O_636,N_4655,N_4498);
nand UO_637 (O_637,N_4559,N_4850);
or UO_638 (O_638,N_4766,N_4649);
or UO_639 (O_639,N_4591,N_4268);
xor UO_640 (O_640,N_4957,N_4351);
xor UO_641 (O_641,N_4525,N_4736);
nor UO_642 (O_642,N_4350,N_4695);
nand UO_643 (O_643,N_4608,N_4836);
or UO_644 (O_644,N_4226,N_4780);
and UO_645 (O_645,N_4775,N_4200);
nand UO_646 (O_646,N_4188,N_4154);
nor UO_647 (O_647,N_4640,N_4504);
nand UO_648 (O_648,N_4126,N_4607);
and UO_649 (O_649,N_4361,N_4655);
nor UO_650 (O_650,N_4616,N_4022);
or UO_651 (O_651,N_4231,N_4108);
nand UO_652 (O_652,N_4187,N_4992);
nand UO_653 (O_653,N_4769,N_4496);
and UO_654 (O_654,N_4213,N_4810);
xnor UO_655 (O_655,N_4585,N_4306);
nor UO_656 (O_656,N_4703,N_4809);
nor UO_657 (O_657,N_4288,N_4534);
nand UO_658 (O_658,N_4276,N_4440);
and UO_659 (O_659,N_4425,N_4872);
and UO_660 (O_660,N_4760,N_4560);
nand UO_661 (O_661,N_4875,N_4569);
nor UO_662 (O_662,N_4512,N_4945);
or UO_663 (O_663,N_4771,N_4435);
and UO_664 (O_664,N_4176,N_4666);
nand UO_665 (O_665,N_4002,N_4575);
xor UO_666 (O_666,N_4794,N_4532);
or UO_667 (O_667,N_4488,N_4672);
xor UO_668 (O_668,N_4553,N_4250);
nor UO_669 (O_669,N_4397,N_4230);
and UO_670 (O_670,N_4304,N_4618);
nor UO_671 (O_671,N_4754,N_4167);
and UO_672 (O_672,N_4284,N_4184);
xor UO_673 (O_673,N_4254,N_4386);
xor UO_674 (O_674,N_4508,N_4911);
nor UO_675 (O_675,N_4612,N_4406);
xor UO_676 (O_676,N_4790,N_4128);
nand UO_677 (O_677,N_4272,N_4233);
nand UO_678 (O_678,N_4344,N_4958);
nand UO_679 (O_679,N_4803,N_4118);
nand UO_680 (O_680,N_4582,N_4320);
xnor UO_681 (O_681,N_4953,N_4086);
or UO_682 (O_682,N_4834,N_4007);
nor UO_683 (O_683,N_4241,N_4137);
nor UO_684 (O_684,N_4988,N_4986);
and UO_685 (O_685,N_4888,N_4506);
and UO_686 (O_686,N_4323,N_4099);
or UO_687 (O_687,N_4114,N_4439);
nand UO_688 (O_688,N_4094,N_4973);
xnor UO_689 (O_689,N_4915,N_4781);
nand UO_690 (O_690,N_4929,N_4200);
nor UO_691 (O_691,N_4845,N_4953);
nor UO_692 (O_692,N_4515,N_4587);
xor UO_693 (O_693,N_4820,N_4447);
and UO_694 (O_694,N_4698,N_4029);
and UO_695 (O_695,N_4834,N_4313);
and UO_696 (O_696,N_4623,N_4183);
and UO_697 (O_697,N_4157,N_4931);
and UO_698 (O_698,N_4314,N_4915);
and UO_699 (O_699,N_4632,N_4758);
and UO_700 (O_700,N_4322,N_4874);
or UO_701 (O_701,N_4106,N_4983);
nand UO_702 (O_702,N_4484,N_4943);
nand UO_703 (O_703,N_4247,N_4251);
xor UO_704 (O_704,N_4705,N_4053);
nor UO_705 (O_705,N_4740,N_4379);
and UO_706 (O_706,N_4833,N_4078);
nor UO_707 (O_707,N_4949,N_4391);
nor UO_708 (O_708,N_4687,N_4712);
xnor UO_709 (O_709,N_4780,N_4625);
or UO_710 (O_710,N_4178,N_4378);
and UO_711 (O_711,N_4278,N_4106);
nor UO_712 (O_712,N_4886,N_4602);
nand UO_713 (O_713,N_4195,N_4076);
or UO_714 (O_714,N_4316,N_4186);
or UO_715 (O_715,N_4250,N_4686);
and UO_716 (O_716,N_4705,N_4497);
nand UO_717 (O_717,N_4653,N_4960);
and UO_718 (O_718,N_4065,N_4295);
nand UO_719 (O_719,N_4438,N_4178);
nand UO_720 (O_720,N_4799,N_4447);
nand UO_721 (O_721,N_4187,N_4995);
and UO_722 (O_722,N_4493,N_4521);
nand UO_723 (O_723,N_4261,N_4288);
nor UO_724 (O_724,N_4731,N_4991);
nand UO_725 (O_725,N_4832,N_4235);
and UO_726 (O_726,N_4527,N_4302);
nand UO_727 (O_727,N_4134,N_4893);
and UO_728 (O_728,N_4340,N_4305);
nor UO_729 (O_729,N_4355,N_4394);
nor UO_730 (O_730,N_4942,N_4451);
and UO_731 (O_731,N_4057,N_4555);
nor UO_732 (O_732,N_4789,N_4867);
xnor UO_733 (O_733,N_4130,N_4442);
nand UO_734 (O_734,N_4420,N_4913);
nand UO_735 (O_735,N_4533,N_4038);
nand UO_736 (O_736,N_4656,N_4810);
or UO_737 (O_737,N_4138,N_4687);
nor UO_738 (O_738,N_4729,N_4580);
xnor UO_739 (O_739,N_4875,N_4832);
and UO_740 (O_740,N_4706,N_4447);
or UO_741 (O_741,N_4112,N_4471);
or UO_742 (O_742,N_4714,N_4236);
nor UO_743 (O_743,N_4266,N_4345);
or UO_744 (O_744,N_4174,N_4237);
nor UO_745 (O_745,N_4338,N_4941);
nor UO_746 (O_746,N_4192,N_4038);
nor UO_747 (O_747,N_4748,N_4964);
nand UO_748 (O_748,N_4824,N_4577);
nor UO_749 (O_749,N_4587,N_4053);
and UO_750 (O_750,N_4897,N_4602);
nand UO_751 (O_751,N_4841,N_4241);
xor UO_752 (O_752,N_4217,N_4708);
and UO_753 (O_753,N_4687,N_4368);
and UO_754 (O_754,N_4820,N_4393);
nand UO_755 (O_755,N_4420,N_4095);
nor UO_756 (O_756,N_4873,N_4624);
and UO_757 (O_757,N_4480,N_4812);
xnor UO_758 (O_758,N_4864,N_4641);
nand UO_759 (O_759,N_4492,N_4004);
and UO_760 (O_760,N_4066,N_4437);
nor UO_761 (O_761,N_4926,N_4200);
and UO_762 (O_762,N_4076,N_4048);
nand UO_763 (O_763,N_4957,N_4404);
nor UO_764 (O_764,N_4386,N_4572);
nor UO_765 (O_765,N_4766,N_4360);
nand UO_766 (O_766,N_4300,N_4513);
and UO_767 (O_767,N_4547,N_4235);
and UO_768 (O_768,N_4370,N_4045);
or UO_769 (O_769,N_4559,N_4793);
or UO_770 (O_770,N_4448,N_4541);
xor UO_771 (O_771,N_4190,N_4095);
nor UO_772 (O_772,N_4711,N_4499);
or UO_773 (O_773,N_4010,N_4284);
nor UO_774 (O_774,N_4386,N_4186);
or UO_775 (O_775,N_4080,N_4779);
nand UO_776 (O_776,N_4670,N_4145);
nor UO_777 (O_777,N_4930,N_4325);
xnor UO_778 (O_778,N_4165,N_4689);
and UO_779 (O_779,N_4465,N_4192);
nor UO_780 (O_780,N_4768,N_4518);
nand UO_781 (O_781,N_4594,N_4620);
nand UO_782 (O_782,N_4052,N_4599);
or UO_783 (O_783,N_4896,N_4759);
or UO_784 (O_784,N_4589,N_4983);
nand UO_785 (O_785,N_4552,N_4943);
nand UO_786 (O_786,N_4388,N_4503);
and UO_787 (O_787,N_4080,N_4970);
or UO_788 (O_788,N_4426,N_4561);
xnor UO_789 (O_789,N_4366,N_4931);
nor UO_790 (O_790,N_4478,N_4267);
nand UO_791 (O_791,N_4303,N_4131);
or UO_792 (O_792,N_4053,N_4161);
nand UO_793 (O_793,N_4818,N_4956);
nand UO_794 (O_794,N_4922,N_4298);
nor UO_795 (O_795,N_4238,N_4211);
nor UO_796 (O_796,N_4298,N_4628);
and UO_797 (O_797,N_4463,N_4010);
or UO_798 (O_798,N_4071,N_4767);
or UO_799 (O_799,N_4213,N_4457);
nor UO_800 (O_800,N_4826,N_4013);
and UO_801 (O_801,N_4637,N_4744);
nor UO_802 (O_802,N_4271,N_4564);
nand UO_803 (O_803,N_4577,N_4595);
nor UO_804 (O_804,N_4946,N_4218);
xor UO_805 (O_805,N_4811,N_4174);
nand UO_806 (O_806,N_4761,N_4726);
and UO_807 (O_807,N_4887,N_4179);
nor UO_808 (O_808,N_4872,N_4573);
nor UO_809 (O_809,N_4261,N_4269);
or UO_810 (O_810,N_4305,N_4594);
nor UO_811 (O_811,N_4975,N_4990);
or UO_812 (O_812,N_4122,N_4233);
nor UO_813 (O_813,N_4986,N_4312);
or UO_814 (O_814,N_4884,N_4163);
nand UO_815 (O_815,N_4805,N_4544);
nand UO_816 (O_816,N_4718,N_4381);
nor UO_817 (O_817,N_4792,N_4097);
nor UO_818 (O_818,N_4036,N_4353);
and UO_819 (O_819,N_4097,N_4919);
nor UO_820 (O_820,N_4876,N_4257);
or UO_821 (O_821,N_4616,N_4066);
nor UO_822 (O_822,N_4935,N_4077);
nand UO_823 (O_823,N_4171,N_4662);
xor UO_824 (O_824,N_4025,N_4651);
nor UO_825 (O_825,N_4646,N_4759);
or UO_826 (O_826,N_4306,N_4644);
and UO_827 (O_827,N_4809,N_4370);
nor UO_828 (O_828,N_4937,N_4029);
or UO_829 (O_829,N_4617,N_4705);
and UO_830 (O_830,N_4488,N_4164);
or UO_831 (O_831,N_4678,N_4845);
nor UO_832 (O_832,N_4439,N_4992);
xor UO_833 (O_833,N_4647,N_4025);
or UO_834 (O_834,N_4193,N_4985);
nand UO_835 (O_835,N_4599,N_4338);
or UO_836 (O_836,N_4287,N_4261);
or UO_837 (O_837,N_4109,N_4841);
xor UO_838 (O_838,N_4034,N_4384);
or UO_839 (O_839,N_4766,N_4784);
xnor UO_840 (O_840,N_4201,N_4315);
nand UO_841 (O_841,N_4392,N_4444);
nand UO_842 (O_842,N_4325,N_4802);
nand UO_843 (O_843,N_4254,N_4599);
nor UO_844 (O_844,N_4765,N_4540);
or UO_845 (O_845,N_4409,N_4571);
nand UO_846 (O_846,N_4509,N_4398);
xnor UO_847 (O_847,N_4510,N_4707);
and UO_848 (O_848,N_4374,N_4957);
xor UO_849 (O_849,N_4032,N_4564);
and UO_850 (O_850,N_4592,N_4333);
nand UO_851 (O_851,N_4560,N_4435);
nand UO_852 (O_852,N_4233,N_4872);
nor UO_853 (O_853,N_4067,N_4164);
nand UO_854 (O_854,N_4047,N_4577);
nand UO_855 (O_855,N_4700,N_4093);
or UO_856 (O_856,N_4718,N_4831);
nor UO_857 (O_857,N_4743,N_4969);
and UO_858 (O_858,N_4193,N_4885);
nor UO_859 (O_859,N_4514,N_4207);
and UO_860 (O_860,N_4694,N_4035);
or UO_861 (O_861,N_4672,N_4778);
nor UO_862 (O_862,N_4511,N_4189);
or UO_863 (O_863,N_4065,N_4733);
nor UO_864 (O_864,N_4027,N_4833);
and UO_865 (O_865,N_4193,N_4240);
or UO_866 (O_866,N_4184,N_4296);
and UO_867 (O_867,N_4196,N_4590);
nand UO_868 (O_868,N_4464,N_4750);
and UO_869 (O_869,N_4043,N_4941);
nor UO_870 (O_870,N_4070,N_4331);
and UO_871 (O_871,N_4529,N_4756);
xor UO_872 (O_872,N_4571,N_4087);
nor UO_873 (O_873,N_4892,N_4962);
and UO_874 (O_874,N_4215,N_4315);
nand UO_875 (O_875,N_4008,N_4710);
nand UO_876 (O_876,N_4455,N_4162);
nor UO_877 (O_877,N_4009,N_4874);
xor UO_878 (O_878,N_4400,N_4504);
nand UO_879 (O_879,N_4277,N_4557);
and UO_880 (O_880,N_4349,N_4111);
xnor UO_881 (O_881,N_4650,N_4373);
or UO_882 (O_882,N_4633,N_4051);
nor UO_883 (O_883,N_4284,N_4589);
nor UO_884 (O_884,N_4456,N_4908);
or UO_885 (O_885,N_4094,N_4226);
or UO_886 (O_886,N_4490,N_4566);
nor UO_887 (O_887,N_4684,N_4800);
xor UO_888 (O_888,N_4244,N_4916);
nor UO_889 (O_889,N_4306,N_4394);
or UO_890 (O_890,N_4296,N_4957);
nand UO_891 (O_891,N_4491,N_4310);
and UO_892 (O_892,N_4704,N_4925);
or UO_893 (O_893,N_4459,N_4465);
nor UO_894 (O_894,N_4636,N_4470);
xnor UO_895 (O_895,N_4151,N_4832);
or UO_896 (O_896,N_4190,N_4228);
nor UO_897 (O_897,N_4896,N_4530);
nor UO_898 (O_898,N_4435,N_4092);
or UO_899 (O_899,N_4284,N_4621);
or UO_900 (O_900,N_4928,N_4156);
or UO_901 (O_901,N_4307,N_4531);
and UO_902 (O_902,N_4376,N_4906);
xor UO_903 (O_903,N_4781,N_4720);
and UO_904 (O_904,N_4870,N_4597);
and UO_905 (O_905,N_4344,N_4959);
and UO_906 (O_906,N_4251,N_4325);
and UO_907 (O_907,N_4257,N_4392);
nor UO_908 (O_908,N_4183,N_4229);
nor UO_909 (O_909,N_4768,N_4352);
nor UO_910 (O_910,N_4608,N_4996);
nand UO_911 (O_911,N_4674,N_4030);
or UO_912 (O_912,N_4078,N_4279);
and UO_913 (O_913,N_4088,N_4782);
nand UO_914 (O_914,N_4733,N_4834);
nor UO_915 (O_915,N_4580,N_4481);
or UO_916 (O_916,N_4563,N_4700);
or UO_917 (O_917,N_4232,N_4190);
xor UO_918 (O_918,N_4779,N_4477);
or UO_919 (O_919,N_4201,N_4589);
and UO_920 (O_920,N_4060,N_4428);
nor UO_921 (O_921,N_4608,N_4266);
or UO_922 (O_922,N_4340,N_4846);
or UO_923 (O_923,N_4299,N_4730);
or UO_924 (O_924,N_4067,N_4674);
or UO_925 (O_925,N_4768,N_4892);
nor UO_926 (O_926,N_4955,N_4431);
or UO_927 (O_927,N_4643,N_4943);
and UO_928 (O_928,N_4833,N_4467);
or UO_929 (O_929,N_4016,N_4189);
and UO_930 (O_930,N_4323,N_4908);
nand UO_931 (O_931,N_4888,N_4917);
and UO_932 (O_932,N_4214,N_4603);
and UO_933 (O_933,N_4840,N_4860);
nand UO_934 (O_934,N_4643,N_4487);
nand UO_935 (O_935,N_4722,N_4275);
or UO_936 (O_936,N_4982,N_4337);
nand UO_937 (O_937,N_4380,N_4869);
or UO_938 (O_938,N_4080,N_4921);
nand UO_939 (O_939,N_4284,N_4273);
nand UO_940 (O_940,N_4763,N_4026);
or UO_941 (O_941,N_4840,N_4054);
nor UO_942 (O_942,N_4241,N_4186);
nor UO_943 (O_943,N_4142,N_4444);
xor UO_944 (O_944,N_4152,N_4543);
and UO_945 (O_945,N_4653,N_4529);
or UO_946 (O_946,N_4089,N_4330);
and UO_947 (O_947,N_4034,N_4928);
nand UO_948 (O_948,N_4624,N_4966);
nor UO_949 (O_949,N_4836,N_4430);
nand UO_950 (O_950,N_4003,N_4988);
or UO_951 (O_951,N_4502,N_4266);
nor UO_952 (O_952,N_4598,N_4440);
or UO_953 (O_953,N_4898,N_4778);
nor UO_954 (O_954,N_4232,N_4078);
nor UO_955 (O_955,N_4568,N_4798);
and UO_956 (O_956,N_4743,N_4194);
and UO_957 (O_957,N_4653,N_4433);
xor UO_958 (O_958,N_4242,N_4346);
nor UO_959 (O_959,N_4263,N_4145);
nor UO_960 (O_960,N_4185,N_4879);
and UO_961 (O_961,N_4628,N_4330);
xnor UO_962 (O_962,N_4522,N_4322);
or UO_963 (O_963,N_4144,N_4487);
or UO_964 (O_964,N_4740,N_4030);
or UO_965 (O_965,N_4484,N_4035);
nand UO_966 (O_966,N_4747,N_4297);
nand UO_967 (O_967,N_4812,N_4520);
nand UO_968 (O_968,N_4931,N_4783);
xnor UO_969 (O_969,N_4692,N_4281);
and UO_970 (O_970,N_4649,N_4109);
and UO_971 (O_971,N_4840,N_4199);
and UO_972 (O_972,N_4716,N_4177);
nand UO_973 (O_973,N_4838,N_4942);
and UO_974 (O_974,N_4987,N_4391);
nand UO_975 (O_975,N_4143,N_4965);
nor UO_976 (O_976,N_4052,N_4233);
nor UO_977 (O_977,N_4120,N_4076);
or UO_978 (O_978,N_4057,N_4873);
or UO_979 (O_979,N_4154,N_4214);
nand UO_980 (O_980,N_4513,N_4861);
nand UO_981 (O_981,N_4516,N_4279);
nor UO_982 (O_982,N_4888,N_4421);
nand UO_983 (O_983,N_4872,N_4765);
or UO_984 (O_984,N_4380,N_4532);
xnor UO_985 (O_985,N_4849,N_4165);
or UO_986 (O_986,N_4132,N_4995);
nand UO_987 (O_987,N_4469,N_4454);
and UO_988 (O_988,N_4957,N_4717);
and UO_989 (O_989,N_4693,N_4855);
nor UO_990 (O_990,N_4299,N_4406);
nand UO_991 (O_991,N_4869,N_4949);
nand UO_992 (O_992,N_4105,N_4502);
nor UO_993 (O_993,N_4830,N_4506);
and UO_994 (O_994,N_4822,N_4382);
or UO_995 (O_995,N_4391,N_4374);
xor UO_996 (O_996,N_4906,N_4454);
nand UO_997 (O_997,N_4472,N_4071);
nand UO_998 (O_998,N_4017,N_4685);
nand UO_999 (O_999,N_4218,N_4051);
endmodule