module basic_3000_30000_3500_5_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
nand U0 (N_0,In_1360,In_1916);
nand U1 (N_1,In_2086,In_2809);
or U2 (N_2,In_1572,In_738);
or U3 (N_3,In_1198,In_156);
xnor U4 (N_4,In_1442,In_2664);
nor U5 (N_5,In_1702,In_2440);
nor U6 (N_6,In_1141,In_1739);
nand U7 (N_7,In_921,In_354);
xor U8 (N_8,In_2810,In_1196);
nor U9 (N_9,In_190,In_425);
nor U10 (N_10,In_2030,In_988);
nand U11 (N_11,In_923,In_480);
xor U12 (N_12,In_2831,In_2042);
nand U13 (N_13,In_2988,In_1811);
xnor U14 (N_14,In_2800,In_407);
xor U15 (N_15,In_1236,In_2136);
nor U16 (N_16,In_1097,In_552);
xnor U17 (N_17,In_1305,In_659);
xnor U18 (N_18,In_691,In_2911);
and U19 (N_19,In_584,In_896);
nor U20 (N_20,In_224,In_1491);
xnor U21 (N_21,In_638,In_2494);
xor U22 (N_22,In_9,In_2002);
xor U23 (N_23,In_2053,In_222);
nand U24 (N_24,In_2408,In_1448);
xor U25 (N_25,In_1072,In_2355);
nand U26 (N_26,In_2660,In_1477);
nand U27 (N_27,In_620,In_574);
and U28 (N_28,In_1210,In_2108);
xnor U29 (N_29,In_1584,In_2533);
nand U30 (N_30,In_1436,In_237);
nor U31 (N_31,In_1770,In_1663);
xor U32 (N_32,In_677,In_2931);
xnor U33 (N_33,In_684,In_999);
xor U34 (N_34,In_2986,In_23);
nor U35 (N_35,In_2389,In_2492);
or U36 (N_36,In_720,In_472);
xor U37 (N_37,In_2903,In_86);
and U38 (N_38,In_1242,In_2701);
xor U39 (N_39,In_1175,In_513);
nor U40 (N_40,In_2825,In_2849);
and U41 (N_41,In_2006,In_1293);
nand U42 (N_42,In_2959,In_2569);
and U43 (N_43,In_475,In_2134);
nand U44 (N_44,In_2535,In_359);
nand U45 (N_45,In_2137,In_2348);
nand U46 (N_46,In_2364,In_551);
or U47 (N_47,In_997,In_1324);
or U48 (N_48,In_1506,In_2901);
and U49 (N_49,In_1283,In_2278);
and U50 (N_50,In_482,In_1250);
xnor U51 (N_51,In_2785,In_990);
nand U52 (N_52,In_1984,In_2674);
or U53 (N_53,In_651,In_395);
and U54 (N_54,In_1886,In_1567);
xnor U55 (N_55,In_2550,In_1214);
and U56 (N_56,In_670,In_2294);
and U57 (N_57,In_2586,In_1775);
xnor U58 (N_58,In_2105,In_2705);
xor U59 (N_59,In_1762,In_2944);
and U60 (N_60,In_424,In_1077);
nand U61 (N_61,In_2438,In_1553);
nand U62 (N_62,In_2595,In_256);
and U63 (N_63,In_641,In_2433);
nor U64 (N_64,In_1009,In_1372);
nand U65 (N_65,In_1426,In_2430);
nor U66 (N_66,In_2017,In_1847);
xor U67 (N_67,In_2806,In_1776);
nand U68 (N_68,In_2425,In_1706);
nor U69 (N_69,In_594,In_1517);
and U70 (N_70,In_1086,In_216);
nor U71 (N_71,In_1381,In_949);
or U72 (N_72,In_823,In_2119);
nand U73 (N_73,In_1824,In_1605);
or U74 (N_74,In_645,In_2422);
nor U75 (N_75,In_51,In_1885);
and U76 (N_76,In_2401,In_2754);
nand U77 (N_77,In_891,In_2194);
xor U78 (N_78,In_1649,In_2565);
xnor U79 (N_79,In_2366,In_2193);
xor U80 (N_80,In_2387,In_2678);
nor U81 (N_81,In_352,In_1037);
or U82 (N_82,In_2204,In_488);
xnor U83 (N_83,In_2324,In_567);
and U84 (N_84,In_2669,In_1264);
or U85 (N_85,In_711,In_2253);
nor U86 (N_86,In_2094,In_2585);
nor U87 (N_87,In_2034,In_2215);
or U88 (N_88,In_540,In_1846);
xnor U89 (N_89,In_2682,In_1493);
nor U90 (N_90,In_1716,In_1058);
or U91 (N_91,In_402,In_2515);
or U92 (N_92,In_2750,In_2673);
nand U93 (N_93,In_1364,In_84);
nand U94 (N_94,In_575,In_47);
nand U95 (N_95,In_1505,In_1760);
or U96 (N_96,In_1528,In_2591);
nor U97 (N_97,In_2715,In_379);
nand U98 (N_98,In_2117,In_1371);
or U99 (N_99,In_193,In_283);
xor U100 (N_100,In_1667,In_2556);
nor U101 (N_101,In_515,In_2311);
and U102 (N_102,In_604,In_1551);
and U103 (N_103,In_1286,In_2263);
nor U104 (N_104,In_933,In_1400);
xnor U105 (N_105,In_511,In_1073);
and U106 (N_106,In_2416,In_1335);
nor U107 (N_107,In_110,In_1231);
nor U108 (N_108,In_2829,In_564);
nand U109 (N_109,In_2512,In_1511);
or U110 (N_110,In_1799,In_2172);
nand U111 (N_111,In_2460,In_2141);
nand U112 (N_112,In_1578,In_2784);
xor U113 (N_113,In_1986,In_2449);
or U114 (N_114,In_2342,In_1905);
nand U115 (N_115,In_2917,In_1970);
nand U116 (N_116,In_209,In_907);
or U117 (N_117,In_2381,In_63);
nor U118 (N_118,In_1162,In_185);
and U119 (N_119,In_523,In_1880);
nor U120 (N_120,In_189,In_559);
nor U121 (N_121,In_446,In_957);
nand U122 (N_122,In_8,In_757);
nand U123 (N_123,In_2457,In_1414);
nand U124 (N_124,In_1951,In_2485);
xnor U125 (N_125,In_1127,In_974);
nor U126 (N_126,In_2361,In_581);
and U127 (N_127,In_788,In_1587);
or U128 (N_128,In_2611,In_592);
and U129 (N_129,In_734,In_806);
and U130 (N_130,In_1096,In_661);
xnor U131 (N_131,In_825,In_2890);
nor U132 (N_132,In_49,In_1806);
nand U133 (N_133,In_2327,In_1140);
nand U134 (N_134,In_1566,In_2865);
nor U135 (N_135,In_2851,In_1615);
and U136 (N_136,In_1326,In_1378);
and U137 (N_137,In_2662,In_672);
xor U138 (N_138,In_674,In_611);
and U139 (N_139,In_439,In_998);
and U140 (N_140,In_1819,In_2158);
nor U141 (N_141,In_862,In_1248);
nor U142 (N_142,In_1105,In_2582);
nor U143 (N_143,In_1919,In_1212);
and U144 (N_144,In_1173,In_1499);
xnor U145 (N_145,In_1366,In_42);
nor U146 (N_146,In_1321,In_1415);
nand U147 (N_147,In_1100,In_375);
or U148 (N_148,In_218,In_2157);
and U149 (N_149,In_2292,In_2385);
xnor U150 (N_150,In_2641,In_1425);
nand U151 (N_151,In_2719,In_2804);
xnor U152 (N_152,In_1380,In_2623);
xnor U153 (N_153,In_2922,In_2548);
and U154 (N_154,In_1390,In_50);
nor U155 (N_155,In_2801,In_633);
nand U156 (N_156,In_2943,In_1546);
and U157 (N_157,In_2722,In_2538);
or U158 (N_158,In_2333,In_1056);
xor U159 (N_159,In_243,In_1808);
or U160 (N_160,In_499,In_750);
nand U161 (N_161,In_1818,In_2124);
xnor U162 (N_162,In_52,In_2060);
nor U163 (N_163,In_184,In_87);
and U164 (N_164,In_920,In_872);
or U165 (N_165,In_2863,In_2270);
or U166 (N_166,In_1855,In_2646);
and U167 (N_167,In_2966,In_1518);
nand U168 (N_168,In_1660,In_1256);
or U169 (N_169,In_285,In_1385);
nor U170 (N_170,In_1482,In_24);
and U171 (N_171,In_883,In_1969);
xnor U172 (N_172,In_1948,In_1298);
and U173 (N_173,In_2041,In_1202);
and U174 (N_174,In_2773,In_214);
xor U175 (N_175,In_2087,In_1642);
or U176 (N_176,In_104,In_1132);
and U177 (N_177,In_541,In_1512);
nor U178 (N_178,In_1875,In_269);
xnor U179 (N_179,In_2073,In_839);
or U180 (N_180,In_247,In_2968);
nand U181 (N_181,In_2313,In_2111);
nand U182 (N_182,In_1756,In_2298);
nor U183 (N_183,In_1745,In_2468);
xnor U184 (N_184,In_2828,In_1558);
xnor U185 (N_185,In_212,In_1085);
and U186 (N_186,In_2789,In_2970);
and U187 (N_187,In_2523,In_2072);
xnor U188 (N_188,In_2207,In_2603);
and U189 (N_189,In_1606,In_1979);
nand U190 (N_190,In_204,In_2596);
nand U191 (N_191,In_1750,In_2875);
and U192 (N_192,In_2409,In_1873);
and U193 (N_193,In_637,In_1592);
nor U194 (N_194,In_2350,In_98);
xnor U195 (N_195,In_1237,In_2707);
or U196 (N_196,In_2549,In_2403);
xor U197 (N_197,In_724,In_1774);
and U198 (N_198,In_2162,In_849);
xnor U199 (N_199,In_2628,In_1475);
xor U200 (N_200,In_2918,In_2915);
nor U201 (N_201,In_969,In_1996);
or U202 (N_202,In_890,In_1942);
nor U203 (N_203,In_2935,In_827);
nand U204 (N_204,In_875,In_2467);
xnor U205 (N_205,In_2496,In_2534);
or U206 (N_206,In_1150,In_1177);
and U207 (N_207,In_1710,In_1523);
xnor U208 (N_208,In_2827,In_1608);
and U209 (N_209,In_1458,In_2772);
nand U210 (N_210,In_1229,In_502);
xor U211 (N_211,In_634,In_1165);
nor U212 (N_212,In_1461,In_444);
nand U213 (N_213,In_1035,In_2228);
and U214 (N_214,In_1797,In_1301);
nand U215 (N_215,In_1252,In_295);
xor U216 (N_216,In_984,In_2394);
and U217 (N_217,In_2266,In_2452);
nand U218 (N_218,In_139,In_2268);
or U219 (N_219,In_1532,In_2599);
and U220 (N_220,In_445,In_693);
or U221 (N_221,In_1272,In_1620);
nand U222 (N_222,In_477,In_1912);
and U223 (N_223,In_400,In_1557);
nand U224 (N_224,In_1598,In_1866);
or U225 (N_225,In_1720,In_1836);
and U226 (N_226,In_2873,In_2652);
nor U227 (N_227,In_174,In_1950);
nand U228 (N_228,In_869,In_336);
and U229 (N_229,In_639,In_625);
xor U230 (N_230,In_1920,In_2584);
xnor U231 (N_231,In_688,In_62);
nand U232 (N_232,In_2615,In_1330);
xor U233 (N_233,In_1722,In_162);
xor U234 (N_234,In_2372,In_2127);
xnor U235 (N_235,In_1675,In_1467);
nand U236 (N_236,In_2131,In_1845);
nand U237 (N_237,In_1831,In_1555);
nor U238 (N_238,In_588,In_2315);
nand U239 (N_239,In_1148,In_1023);
or U240 (N_240,In_2781,In_1123);
nor U241 (N_241,In_1306,In_1643);
nand U242 (N_242,In_1652,In_629);
nand U243 (N_243,In_2335,In_173);
and U244 (N_244,In_506,In_2690);
and U245 (N_245,In_2798,In_483);
nand U246 (N_246,In_2428,In_2469);
xnor U247 (N_247,In_731,In_2888);
or U248 (N_248,In_1524,In_353);
or U249 (N_249,In_1794,In_1695);
and U250 (N_250,In_2256,In_1471);
and U251 (N_251,In_1373,In_341);
or U252 (N_252,In_2067,In_368);
and U253 (N_253,In_662,In_2767);
nand U254 (N_254,In_1787,In_361);
nand U255 (N_255,In_982,In_2606);
nand U256 (N_256,In_2720,In_2638);
nand U257 (N_257,In_178,In_942);
nor U258 (N_258,In_1707,In_573);
or U259 (N_259,In_2564,In_260);
nor U260 (N_260,In_1176,In_2122);
nand U261 (N_261,In_1342,In_2741);
and U262 (N_262,In_1358,In_1392);
xor U263 (N_263,In_1561,In_1136);
or U264 (N_264,In_713,In_1693);
or U265 (N_265,In_1868,In_300);
nor U266 (N_266,In_1815,In_366);
and U267 (N_267,In_207,In_2483);
and U268 (N_268,In_970,In_2693);
xnor U269 (N_269,In_1405,In_2214);
xor U270 (N_270,In_1893,In_314);
nor U271 (N_271,In_1998,In_697);
and U272 (N_272,In_2459,In_2503);
xor U273 (N_273,In_1375,In_1904);
nor U274 (N_274,In_2349,In_580);
nand U275 (N_275,In_369,In_195);
and U276 (N_276,In_373,In_851);
and U277 (N_277,In_1357,In_649);
and U278 (N_278,In_2580,In_2198);
or U279 (N_279,In_986,In_2790);
nand U280 (N_280,In_2530,In_2223);
nand U281 (N_281,In_2985,In_2151);
nand U282 (N_282,In_1768,In_1648);
xnor U283 (N_283,In_1267,In_2390);
nor U284 (N_284,In_2993,In_1903);
nand U285 (N_285,In_981,In_1317);
or U286 (N_286,In_440,In_2012);
nor U287 (N_287,In_1792,In_155);
and U288 (N_288,In_137,In_1851);
nor U289 (N_289,In_1657,In_1311);
nand U290 (N_290,In_2893,In_2761);
nor U291 (N_291,In_2926,In_2532);
and U292 (N_292,In_1325,In_1758);
nor U293 (N_293,In_1068,In_2008);
or U294 (N_294,In_2044,In_27);
xnor U295 (N_295,In_384,In_78);
or U296 (N_296,In_1895,In_121);
and U297 (N_297,In_1925,In_874);
nand U298 (N_298,In_1694,In_2511);
and U299 (N_299,In_610,In_2419);
nand U300 (N_300,In_2818,In_1402);
and U301 (N_301,In_2451,In_1600);
nand U302 (N_302,In_2484,In_2631);
nand U303 (N_303,In_1391,In_2112);
xor U304 (N_304,In_1839,In_2153);
or U305 (N_305,In_1991,In_1501);
or U306 (N_306,In_505,In_1931);
nand U307 (N_307,In_2259,In_142);
or U308 (N_308,In_1914,In_2411);
and U309 (N_309,In_2553,In_943);
nor U310 (N_310,In_2144,In_2125);
nor U311 (N_311,In_433,In_2659);
xor U312 (N_312,In_698,In_2161);
xnor U313 (N_313,In_1790,In_2844);
or U314 (N_314,In_1673,In_2116);
xor U315 (N_315,In_884,In_778);
and U316 (N_316,In_1939,In_962);
or U317 (N_317,In_1533,In_2003);
xnor U318 (N_318,In_1536,In_1370);
xor U319 (N_319,In_2129,In_1275);
nand U320 (N_320,In_1732,In_805);
xnor U321 (N_321,In_297,In_2681);
xor U322 (N_322,In_168,In_529);
nor U323 (N_323,In_699,In_2597);
xor U324 (N_324,In_2517,In_550);
nor U325 (N_325,In_164,In_1021);
nand U326 (N_326,In_221,In_2814);
nor U327 (N_327,In_763,In_2883);
xnor U328 (N_328,In_2021,In_1701);
nand U329 (N_329,In_263,In_1352);
or U330 (N_330,In_2453,In_593);
nand U331 (N_331,In_725,In_2149);
nor U332 (N_332,In_2946,In_1435);
or U333 (N_333,In_1046,In_329);
and U334 (N_334,In_2380,In_1539);
nor U335 (N_335,In_1336,In_945);
xnor U336 (N_336,In_1308,In_2588);
xor U337 (N_337,In_394,In_2028);
xnor U338 (N_338,In_1987,In_423);
nor U339 (N_339,In_1676,In_1923);
nor U340 (N_340,In_2442,In_2032);
nor U341 (N_341,In_1222,In_1227);
and U342 (N_342,In_2739,In_801);
nor U343 (N_343,In_2326,In_449);
xor U344 (N_344,In_723,In_249);
xor U345 (N_345,In_1947,In_1469);
xor U346 (N_346,In_1091,In_356);
or U347 (N_347,In_55,In_2482);
nand U348 (N_348,In_1929,In_1069);
nor U349 (N_349,In_1502,In_1946);
nand U350 (N_350,In_2885,In_2774);
nand U351 (N_351,In_2651,In_646);
or U352 (N_352,In_210,In_2896);
xnor U353 (N_353,In_2080,In_2027);
nand U354 (N_354,In_422,In_2264);
or U355 (N_355,In_898,In_1120);
or U356 (N_356,In_2793,In_2300);
and U357 (N_357,In_1788,In_1757);
and U358 (N_358,In_2843,In_1698);
and U359 (N_359,In_2920,In_2872);
and U360 (N_360,In_11,In_696);
nor U361 (N_361,In_1130,In_1971);
xnor U362 (N_362,In_987,In_663);
xor U363 (N_363,In_1821,In_961);
and U364 (N_364,In_977,In_1934);
and U365 (N_365,In_1447,In_2964);
xor U366 (N_366,In_312,In_844);
and U367 (N_367,In_1007,In_1463);
or U368 (N_368,In_251,In_2991);
or U369 (N_369,In_279,In_950);
and U370 (N_370,In_1044,In_2730);
xor U371 (N_371,In_231,In_1483);
nand U372 (N_372,In_2527,In_2634);
and U373 (N_373,In_2639,In_1852);
nand U374 (N_374,In_673,In_1179);
nand U375 (N_375,In_1459,In_1737);
nor U376 (N_376,In_1801,In_2692);
nor U377 (N_377,In_2206,In_2057);
nand U378 (N_378,In_1688,In_2960);
or U379 (N_379,In_2466,In_1954);
or U380 (N_380,In_1060,In_2925);
nor U381 (N_381,In_2933,In_2953);
xnor U382 (N_382,In_1257,In_364);
nand U383 (N_383,In_2617,In_1901);
xor U384 (N_384,In_1974,In_1274);
nor U385 (N_385,In_814,In_2842);
or U386 (N_386,In_1441,In_2543);
or U387 (N_387,In_188,In_702);
nor U388 (N_388,In_2076,In_274);
or U389 (N_389,In_2813,In_1258);
xnor U390 (N_390,In_1633,In_2402);
nand U391 (N_391,In_2643,In_5);
or U392 (N_392,In_1235,In_1853);
nand U393 (N_393,In_1396,In_331);
nand U394 (N_394,In_2272,In_1115);
or U395 (N_395,In_1327,In_1464);
nand U396 (N_396,In_1485,In_2627);
or U397 (N_397,In_1356,In_798);
nor U398 (N_398,In_1940,In_2344);
or U399 (N_399,In_2899,In_2473);
or U400 (N_400,In_595,In_809);
nor U401 (N_401,In_766,In_2587);
nand U402 (N_402,In_2365,In_1936);
xnor U403 (N_403,In_853,In_810);
xnor U404 (N_404,In_1446,In_1423);
nor U405 (N_405,In_2299,In_1090);
and U406 (N_406,In_924,In_76);
nand U407 (N_407,In_1225,In_1771);
and U408 (N_408,In_1027,In_1409);
and U409 (N_409,In_2984,In_208);
nand U410 (N_410,In_351,In_701);
nor U411 (N_411,In_1753,In_320);
or U412 (N_412,In_1238,In_270);
or U413 (N_413,In_315,In_1602);
or U414 (N_414,In_1245,In_2213);
and U415 (N_415,In_632,In_1190);
and U416 (N_416,In_1348,In_873);
nor U417 (N_417,In_2269,In_668);
and U418 (N_418,In_334,In_1583);
or U419 (N_419,In_335,In_2765);
or U420 (N_420,In_159,In_271);
nand U421 (N_421,In_1455,In_128);
xor U422 (N_422,In_979,In_1050);
nand U423 (N_423,In_2540,In_2520);
xor U424 (N_424,In_1055,In_25);
or U425 (N_425,In_2497,In_1922);
and U426 (N_426,In_861,In_1353);
nand U427 (N_427,In_2637,In_765);
and U428 (N_428,In_1544,In_1629);
nor U429 (N_429,In_776,In_2656);
nor U430 (N_430,In_2011,In_1167);
nor U431 (N_431,In_153,In_870);
nand U432 (N_432,In_2519,In_2329);
or U433 (N_433,In_733,In_937);
nor U434 (N_434,In_228,In_215);
nand U435 (N_435,In_570,In_124);
nor U436 (N_436,In_141,In_10);
or U437 (N_437,In_736,In_1443);
nor U438 (N_438,In_1266,In_254);
nand U439 (N_439,In_2839,In_793);
xnor U440 (N_440,In_2531,In_507);
and U441 (N_441,In_1662,In_266);
nor U442 (N_442,In_2794,In_1133);
and U443 (N_443,In_2514,In_2636);
nor U444 (N_444,In_1376,In_2205);
and U445 (N_445,In_1783,In_2091);
nor U446 (N_446,In_1647,In_1419);
nand U447 (N_447,In_1717,In_1010);
and U448 (N_448,In_6,In_172);
xnor U449 (N_449,In_1387,In_1755);
or U450 (N_450,In_2229,In_2501);
nand U451 (N_451,In_1661,In_888);
nor U452 (N_452,In_1014,In_2224);
nand U453 (N_453,In_556,In_1589);
or U454 (N_454,In_457,In_1444);
nor U455 (N_455,In_2826,In_2846);
nand U456 (N_456,In_1128,In_2330);
or U457 (N_457,In_992,In_817);
xnor U458 (N_458,In_2123,In_238);
and U459 (N_459,In_1457,In_2441);
and U460 (N_460,In_1273,In_2051);
xnor U461 (N_461,In_2358,In_2293);
and U462 (N_462,In_548,In_1842);
and U463 (N_463,In_1084,In_689);
nand U464 (N_464,In_1692,In_690);
nor U465 (N_465,In_2328,In_1725);
nor U466 (N_466,In_605,In_347);
nor U467 (N_467,In_1197,In_2574);
or U468 (N_468,In_1782,In_2928);
and U469 (N_469,In_1408,In_119);
nand U470 (N_470,In_2322,In_1896);
nor U471 (N_471,In_2747,In_1961);
nor U472 (N_472,In_66,In_2762);
xnor U473 (N_473,In_2850,In_1285);
and U474 (N_474,In_508,In_2019);
and U475 (N_475,In_728,In_2861);
and U476 (N_476,In_1881,In_2462);
nor U477 (N_477,In_273,In_281);
xnor U478 (N_478,In_2504,In_2963);
xnor U479 (N_479,In_2434,In_2886);
and U480 (N_480,In_236,In_2823);
nor U481 (N_481,In_2895,In_2780);
and U482 (N_482,In_2235,In_2035);
xor U483 (N_483,In_54,In_913);
or U484 (N_484,In_2495,In_2536);
or U485 (N_485,In_2887,In_1254);
nand U486 (N_486,In_1193,In_2188);
nand U487 (N_487,In_932,In_1080);
or U488 (N_488,In_1837,In_452);
nand U489 (N_489,In_2095,In_1063);
and U490 (N_490,In_2238,In_2797);
nor U491 (N_491,In_2261,In_2649);
and U492 (N_492,In_2957,In_758);
or U493 (N_493,In_1144,In_2479);
nor U494 (N_494,In_1681,In_404);
nand U495 (N_495,In_2697,In_307);
and U496 (N_496,In_1045,In_455);
nand U497 (N_497,In_67,In_177);
and U498 (N_498,In_1569,In_1843);
and U499 (N_499,In_2220,In_2316);
xnor U500 (N_500,In_2562,In_1389);
and U501 (N_501,In_2276,In_374);
and U502 (N_502,In_2868,In_928);
nor U503 (N_503,In_808,In_2472);
nor U504 (N_504,In_2277,In_1460);
or U505 (N_505,In_1111,In_2165);
and U506 (N_506,In_2100,In_528);
xnor U507 (N_507,In_1051,In_2647);
nand U508 (N_508,In_2209,In_2219);
nand U509 (N_509,In_2783,In_1205);
or U510 (N_510,In_2120,In_2320);
or U511 (N_511,In_1966,In_2982);
or U512 (N_512,In_2642,In_2216);
or U513 (N_513,In_2581,In_700);
nand U514 (N_514,In_2176,In_1181);
and U515 (N_515,In_1430,In_1398);
and U516 (N_516,In_678,In_3);
and U517 (N_517,In_1560,In_1169);
xnor U518 (N_518,In_2132,In_2847);
nand U519 (N_519,In_301,In_1634);
and U520 (N_520,In_2305,In_1344);
xor U521 (N_521,In_2724,In_1048);
xnor U522 (N_522,In_2729,In_2371);
nor U523 (N_523,In_2306,In_618);
nand U524 (N_524,In_1840,In_1967);
and U525 (N_525,In_783,In_1395);
nor U526 (N_526,In_414,In_2249);
nand U527 (N_527,In_2170,In_275);
nor U528 (N_528,In_1221,In_485);
nand U529 (N_529,In_2561,In_495);
or U530 (N_530,In_1208,In_892);
xnor U531 (N_531,In_1654,In_2152);
xor U532 (N_532,In_357,In_756);
and U533 (N_533,In_1319,In_145);
and U534 (N_534,In_1593,In_2558);
xor U535 (N_535,In_1804,In_2420);
xor U536 (N_536,In_2845,In_2241);
xor U537 (N_537,In_2480,In_1714);
nor U538 (N_538,In_199,In_2481);
or U539 (N_539,In_2323,In_82);
xnor U540 (N_540,In_233,In_2869);
or U541 (N_541,In_561,In_365);
xnor U542 (N_542,In_2735,In_1738);
nand U543 (N_543,In_1333,In_642);
and U544 (N_544,In_836,In_837);
and U545 (N_545,In_2745,In_393);
xnor U546 (N_546,In_2791,In_1070);
and U547 (N_547,In_735,In_2362);
and U548 (N_548,In_1708,In_333);
nor U549 (N_549,In_833,In_1307);
or U550 (N_550,In_1427,In_1339);
nand U551 (N_551,In_2083,In_818);
nor U552 (N_552,In_2068,In_1883);
xor U553 (N_553,In_1713,In_909);
xor U554 (N_554,In_1057,In_348);
and U555 (N_555,In_2318,In_2871);
nand U556 (N_556,In_1182,In_784);
nor U557 (N_557,In_1472,In_2560);
or U558 (N_558,In_2099,In_2169);
xnor U559 (N_559,In_1607,In_288);
nand U560 (N_560,In_143,In_621);
nand U561 (N_561,In_2396,In_1204);
xnor U562 (N_562,In_2317,In_1424);
nand U563 (N_563,In_1052,In_383);
nor U564 (N_564,In_903,In_1071);
xor U565 (N_565,In_2274,In_2128);
xnor U566 (N_566,In_103,In_127);
nand U567 (N_567,In_501,In_1594);
nand U568 (N_568,In_264,In_2471);
nor U569 (N_569,In_1029,In_653);
nand U570 (N_570,In_2413,In_2231);
or U571 (N_571,In_1418,In_61);
xnor U572 (N_572,In_1478,In_1036);
nand U573 (N_573,In_122,In_120);
nand U574 (N_574,In_1440,In_519);
nand U575 (N_575,In_899,In_148);
nor U576 (N_576,In_2179,In_2539);
nand U577 (N_577,In_2456,In_2513);
xor U578 (N_578,In_2275,In_1278);
nor U579 (N_579,In_2291,In_239);
xor U580 (N_580,In_1937,In_526);
and U581 (N_581,In_2677,In_1684);
nor U582 (N_582,In_2653,In_747);
or U583 (N_583,In_2732,In_2341);
and U584 (N_584,In_1296,In_2196);
xnor U585 (N_585,In_2889,In_4);
xor U586 (N_586,In_654,In_846);
or U587 (N_587,In_2879,In_2601);
nand U588 (N_588,In_958,In_2633);
or U589 (N_589,In_43,In_412);
or U590 (N_590,In_2995,In_708);
nor U591 (N_591,In_2516,In_2190);
xnor U592 (N_592,In_2180,In_2786);
and U593 (N_593,In_2431,In_876);
nand U594 (N_594,In_1577,In_740);
xor U595 (N_595,In_1779,In_1059);
nor U596 (N_596,In_2178,In_1312);
nor U597 (N_597,In_31,In_612);
or U598 (N_598,In_2109,In_2302);
nand U599 (N_599,In_1399,In_2375);
and U600 (N_600,In_2163,In_785);
and U601 (N_601,In_1240,In_1433);
and U602 (N_602,In_1599,In_1889);
nor U603 (N_603,In_2436,In_255);
nor U604 (N_604,In_767,In_1382);
nand U605 (N_605,In_1924,In_1064);
and U606 (N_606,In_1363,In_2183);
nand U607 (N_607,In_205,In_569);
nand U608 (N_608,In_56,In_2343);
xnor U609 (N_609,In_1752,In_169);
nor U610 (N_610,In_1913,In_2225);
xor U611 (N_611,In_40,In_2838);
nor U612 (N_612,In_664,In_349);
nor U613 (N_613,In_2771,In_1580);
and U614 (N_614,In_2836,In_2740);
nand U615 (N_615,In_2001,In_1597);
nand U616 (N_616,In_2775,In_695);
xnor U617 (N_617,In_1001,In_2731);
xor U618 (N_618,In_290,In_1907);
and U619 (N_619,In_1726,In_1146);
nor U620 (N_620,In_1462,In_754);
xnor U621 (N_621,In_1476,In_1246);
and U622 (N_622,In_497,In_2212);
or U623 (N_623,In_2426,In_2589);
nor U624 (N_624,In_2061,In_859);
or U625 (N_625,In_1420,In_1172);
or U626 (N_626,In_1089,In_2749);
nand U627 (N_627,In_901,In_1576);
and U628 (N_628,In_2702,In_1259);
xor U629 (N_629,In_1030,In_2725);
nor U630 (N_630,In_650,In_560);
xor U631 (N_631,In_161,In_2542);
nor U632 (N_632,In_991,In_1975);
nand U633 (N_633,In_2414,In_1552);
and U634 (N_634,In_2082,In_2974);
or U635 (N_635,In_665,In_1671);
nand U636 (N_636,In_2703,In_1864);
nand U637 (N_637,In_2555,In_1754);
or U638 (N_638,In_2738,In_1340);
or U639 (N_639,In_2308,In_252);
or U640 (N_640,In_1042,In_1610);
xor U641 (N_641,In_261,In_2242);
nor U642 (N_642,In_2075,In_980);
nor U643 (N_643,In_2078,In_1451);
nand U644 (N_644,In_1749,In_1094);
or U645 (N_645,In_2185,In_1345);
and U646 (N_646,In_1740,In_2951);
or U647 (N_647,In_835,In_812);
nand U648 (N_648,In_435,In_181);
and U649 (N_649,In_2427,In_1092);
or U650 (N_650,In_1117,In_340);
nand U651 (N_651,In_1727,In_1316);
nand U652 (N_652,In_1011,In_2279);
nand U653 (N_653,In_183,In_131);
and U654 (N_654,In_1134,In_259);
nor U655 (N_655,In_432,In_1571);
xor U656 (N_656,In_590,In_1489);
nor U657 (N_657,In_1962,In_781);
nor U658 (N_658,In_1786,In_1268);
xnor U659 (N_659,In_1184,In_2992);
nand U660 (N_660,In_732,In_1005);
xnor U661 (N_661,In_154,In_685);
nand U662 (N_662,In_490,In_1802);
xnor U663 (N_663,In_500,In_562);
xor U664 (N_664,In_72,In_0);
xnor U665 (N_665,In_1062,In_1521);
nand U666 (N_666,In_123,In_2488);
xor U667 (N_667,In_2004,In_2572);
nor U668 (N_668,In_2937,In_2622);
nor U669 (N_669,In_1535,In_985);
or U670 (N_670,In_420,In_676);
xnor U671 (N_671,In_2866,In_346);
nand U672 (N_672,In_902,In_1854);
and U673 (N_673,In_1361,In_2619);
nand U674 (N_674,In_470,In_675);
and U675 (N_675,In_607,In_126);
and U676 (N_676,In_563,In_1049);
xnor U677 (N_677,In_2945,In_2280);
nor U678 (N_678,In_2417,In_512);
and U679 (N_679,In_2718,In_832);
and U680 (N_680,In_669,In_2544);
and U681 (N_681,In_2189,In_1174);
xnor U682 (N_682,In_886,In_2952);
and U683 (N_683,In_804,In_2064);
xor U684 (N_684,In_391,In_622);
nor U685 (N_685,In_158,In_2281);
nor U686 (N_686,In_2687,In_2029);
xnor U687 (N_687,In_1980,In_321);
or U688 (N_688,In_1495,In_729);
nand U689 (N_689,In_815,In_292);
nor U690 (N_690,In_1158,In_2612);
and U691 (N_691,In_1988,In_2246);
or U692 (N_692,In_647,In_1581);
and U693 (N_693,In_2036,In_1926);
or U694 (N_694,In_327,In_2133);
and U695 (N_695,In_2575,In_1575);
xnor U696 (N_696,In_2607,In_1183);
and U697 (N_697,In_1322,In_813);
xor U698 (N_698,In_1249,In_880);
nor U699 (N_699,In_1261,In_2038);
or U700 (N_700,In_234,In_410);
nand U701 (N_701,In_2526,In_2140);
nor U702 (N_702,In_2421,In_1565);
nand U703 (N_703,In_2388,In_2546);
nor U704 (N_704,In_2821,In_577);
and U705 (N_705,In_187,In_739);
nor U706 (N_706,In_2458,In_135);
nor U707 (N_707,In_2805,In_1941);
and U708 (N_708,In_461,In_644);
nor U709 (N_709,In_2378,In_1809);
or U710 (N_710,In_2626,In_834);
or U711 (N_711,In_182,In_782);
xnor U712 (N_712,In_2769,In_2833);
or U713 (N_713,In_1705,In_1848);
nor U714 (N_714,In_323,In_1679);
nor U715 (N_715,In_521,In_1498);
and U716 (N_716,In_191,In_1000);
and U717 (N_717,In_1943,In_1156);
or U718 (N_718,In_1026,In_1087);
nand U719 (N_719,In_1365,In_978);
and U720 (N_720,In_1891,In_2445);
and U721 (N_721,In_1411,In_565);
nand U722 (N_722,In_1299,In_709);
nand U723 (N_723,In_771,In_2616);
xnor U724 (N_724,In_1730,In_679);
nand U725 (N_725,In_1910,In_2766);
nand U726 (N_726,In_2962,In_2854);
nor U727 (N_727,In_1742,In_419);
nand U728 (N_728,In_1972,In_585);
nor U729 (N_729,In_2948,In_2712);
or U730 (N_730,In_1473,In_2424);
nor U731 (N_731,In_838,In_1061);
xor U732 (N_732,In_2251,In_545);
and U733 (N_733,In_1484,In_557);
and U734 (N_734,In_2150,In_2912);
or U735 (N_735,In_176,In_1949);
nor U736 (N_736,In_1816,In_2071);
and U737 (N_737,In_1468,In_1012);
xnor U738 (N_738,In_860,In_1829);
or U739 (N_739,In_1351,In_630);
nor U740 (N_740,In_2613,In_2713);
xnor U741 (N_741,In_2245,In_1686);
or U742 (N_742,In_140,In_2967);
or U743 (N_743,In_1530,In_2084);
nand U744 (N_744,In_1689,In_2448);
or U745 (N_745,In_2486,In_372);
xnor U746 (N_746,In_1263,In_759);
nor U747 (N_747,In_931,In_318);
or U748 (N_748,In_617,In_777);
and U749 (N_749,In_232,In_2559);
and U750 (N_750,In_309,In_1614);
and U751 (N_751,In_2181,In_442);
xnor U752 (N_752,In_1277,In_1088);
or U753 (N_753,In_1865,In_1765);
nor U754 (N_754,In_1718,In_2676);
and U755 (N_755,In_1860,In_2217);
and U756 (N_756,In_426,In_1480);
xnor U757 (N_757,In_887,In_2524);
or U758 (N_758,In_1294,In_968);
nand U759 (N_759,In_2050,In_2691);
or U760 (N_760,In_773,In_1219);
xnor U761 (N_761,In_2894,In_1228);
nor U762 (N_762,In_1932,In_789);
and U763 (N_763,In_1683,In_1313);
nor U764 (N_764,In_1206,In_1066);
nand U765 (N_765,In_2373,In_1412);
or U766 (N_766,In_1659,In_2675);
or U767 (N_767,In_623,In_1751);
nor U768 (N_768,In_2807,In_2347);
xnor U769 (N_769,In_2498,In_2429);
or U770 (N_770,In_476,In_919);
and U771 (N_771,In_1990,In_1122);
and U772 (N_772,In_257,In_2777);
and U773 (N_773,In_2054,In_1908);
nor U774 (N_774,In_2906,In_70);
and U775 (N_775,In_7,In_2285);
xor U776 (N_776,In_1022,In_2590);
or U777 (N_777,In_1189,In_1563);
nor U778 (N_778,In_1582,In_109);
nor U779 (N_779,In_451,In_2882);
and U780 (N_780,In_2927,In_456);
or U781 (N_781,In_1421,In_2858);
or U782 (N_782,In_376,In_385);
nand U783 (N_783,In_579,In_345);
nand U784 (N_784,In_1744,In_1810);
or U785 (N_785,In_828,In_388);
nand U786 (N_786,In_2924,In_889);
nor U787 (N_787,In_94,In_1107);
nand U788 (N_788,In_1841,In_466);
nor U789 (N_789,In_2618,In_2635);
nand U790 (N_790,In_2470,In_1915);
or U791 (N_791,In_1288,In_2583);
and U792 (N_792,In_447,In_2999);
nand U793 (N_793,In_305,In_227);
or U794 (N_794,In_2,In_2552);
nand U795 (N_795,In_2423,In_2391);
xnor U796 (N_796,In_299,In_583);
nand U797 (N_797,In_1869,In_401);
and U798 (N_798,In_1276,In_2499);
or U799 (N_799,In_2525,In_606);
xnor U800 (N_800,In_956,In_2648);
and U801 (N_801,In_1508,In_1766);
xor U802 (N_802,In_481,In_29);
nor U803 (N_803,In_681,In_1729);
nor U804 (N_804,In_289,In_2052);
nor U805 (N_805,In_925,In_166);
or U806 (N_806,In_1978,In_2138);
or U807 (N_807,In_1157,In_1888);
or U808 (N_808,In_1636,In_1777);
nor U809 (N_809,In_1284,In_596);
and U810 (N_810,In_2579,In_217);
and U811 (N_811,In_77,In_2369);
or U812 (N_812,In_478,In_2755);
and U813 (N_813,In_996,In_1858);
or U814 (N_814,In_250,In_1232);
xnor U815 (N_815,In_302,In_905);
nand U816 (N_816,In_2287,In_74);
and U817 (N_817,In_1013,In_1812);
or U818 (N_818,In_2024,In_17);
nor U819 (N_819,In_12,In_1076);
xor U820 (N_820,In_2763,In_2862);
xor U821 (N_821,In_1796,In_1354);
and U822 (N_822,In_2186,In_2812);
nand U823 (N_823,In_1639,In_726);
and U824 (N_824,In_975,In_2288);
nor U825 (N_825,In_2367,In_100);
nand U826 (N_826,In_794,In_1002);
xor U827 (N_827,In_1825,In_1791);
nor U828 (N_828,In_2013,In_1006);
and U829 (N_829,In_1884,In_1622);
and U830 (N_830,In_944,In_2840);
nand U831 (N_831,In_742,In_658);
or U832 (N_832,In_1004,In_1867);
or U833 (N_833,In_2878,In_2130);
xor U834 (N_834,In_1406,In_2733);
nand U835 (N_835,In_399,In_1403);
and U836 (N_836,In_566,In_2630);
or U837 (N_837,In_1793,In_1763);
nand U838 (N_838,In_2950,In_2644);
and U839 (N_839,In_213,In_965);
or U840 (N_840,In_2592,In_83);
xnor U841 (N_841,In_845,In_1159);
and U842 (N_842,In_125,In_1509);
nand U843 (N_843,In_2655,In_2891);
and U844 (N_844,In_2598,In_2696);
nand U845 (N_845,In_2529,In_857);
nor U846 (N_846,In_1909,In_910);
nand U847 (N_847,In_65,In_2939);
nand U848 (N_848,In_1666,In_2090);
or U849 (N_849,In_1187,In_948);
or U850 (N_850,In_769,In_2248);
xnor U851 (N_851,In_392,In_2788);
nor U852 (N_852,In_850,In_1828);
xor U853 (N_853,In_2444,In_1338);
or U854 (N_854,In_1613,In_167);
nand U855 (N_855,In_2716,In_1217);
xnor U856 (N_856,In_922,In_1985);
xor U857 (N_857,In_1239,In_1194);
nand U858 (N_858,In_36,In_703);
and U859 (N_859,In_2014,In_2803);
and U860 (N_860,In_2247,In_245);
or U861 (N_861,In_53,In_2476);
xor U862 (N_862,In_363,In_2443);
nor U863 (N_863,In_325,In_2455);
or U864 (N_864,In_2704,In_462);
and U865 (N_865,In_362,In_1712);
and U866 (N_866,In_2257,In_994);
nor U867 (N_867,In_1665,In_1520);
or U868 (N_868,In_1761,In_816);
and U869 (N_869,In_1935,In_966);
xor U870 (N_870,In_108,In_2508);
or U871 (N_871,In_2727,In_2567);
or U872 (N_872,In_856,In_2621);
nor U873 (N_873,In_536,In_1618);
xor U874 (N_874,In_2779,In_745);
nand U875 (N_875,In_1554,In_1160);
and U876 (N_876,In_1672,In_2941);
nand U877 (N_877,In_2521,In_2092);
or U878 (N_878,In_1164,In_112);
xor U879 (N_879,In_2142,In_894);
and U880 (N_880,In_1585,In_332);
and U881 (N_881,In_1525,In_2221);
xor U882 (N_882,In_780,In_2670);
nor U883 (N_883,In_2066,In_350);
nand U884 (N_884,In_165,In_2368);
nand U885 (N_885,In_1835,In_2898);
nand U886 (N_886,In_1780,In_1767);
nor U887 (N_887,In_304,In_2191);
nor U888 (N_888,In_1721,In_820);
or U889 (N_889,In_555,In_2088);
or U890 (N_890,In_527,In_2684);
nor U891 (N_891,In_330,In_601);
nand U892 (N_892,In_102,In_1215);
nand U893 (N_893,In_1466,In_35);
nand U894 (N_894,In_2192,In_504);
and U895 (N_895,In_319,In_30);
and U896 (N_896,In_1538,In_286);
xnor U897 (N_897,In_2356,In_1432);
nor U898 (N_898,In_542,In_2657);
nor U899 (N_899,In_316,In_48);
nor U900 (N_900,In_1347,In_13);
or U901 (N_901,In_1997,In_2016);
nor U902 (N_902,In_1188,In_2304);
xnor U903 (N_903,In_33,In_377);
nand U904 (N_904,In_2309,In_2352);
xor U905 (N_905,In_683,In_2679);
or U906 (N_906,In_960,In_530);
or U907 (N_907,In_1668,In_1075);
nor U908 (N_908,In_1747,In_1481);
xor U909 (N_909,In_2841,In_2243);
nand U910 (N_910,In_2173,In_284);
or U911 (N_911,In_484,In_1724);
nand U912 (N_912,In_2464,In_2295);
nor U913 (N_913,In_2489,In_608);
and U914 (N_914,In_1832,In_2742);
nor U915 (N_915,In_2166,In_1397);
xor U916 (N_916,In_2258,In_1233);
or U917 (N_917,In_1927,In_2977);
nand U918 (N_918,In_1149,In_1989);
nor U919 (N_919,In_1251,In_1616);
nand U920 (N_920,In_2359,In_115);
nor U921 (N_921,In_69,In_460);
nand U922 (N_922,In_431,In_2255);
nor U923 (N_923,In_753,In_522);
nor U924 (N_924,In_847,In_58);
and U925 (N_925,In_2680,In_2020);
xor U926 (N_926,In_885,In_831);
nor U927 (N_927,In_1515,In_2155);
or U928 (N_928,In_413,In_1850);
and U929 (N_929,In_2998,In_2936);
nand U930 (N_930,In_2958,In_1870);
nor U931 (N_931,In_2154,In_2577);
nand U932 (N_932,In_276,In_1394);
nor U933 (N_933,In_277,In_2852);
and U934 (N_934,In_941,In_1703);
and U935 (N_935,In_1126,In_947);
xnor U936 (N_936,In_865,In_1145);
nor U937 (N_937,In_1295,In_1496);
or U938 (N_938,In_2250,In_2683);
or U939 (N_939,In_2446,In_772);
or U940 (N_940,In_1677,In_1124);
nand U941 (N_941,In_2537,In_871);
nand U942 (N_942,In_223,In_1281);
and U943 (N_943,In_133,In_971);
and U944 (N_944,In_2354,In_614);
or U945 (N_945,In_2500,In_427);
and U946 (N_946,In_2033,In_1329);
xor U947 (N_947,In_2233,In_150);
or U948 (N_948,In_1103,In_2557);
nor U949 (N_949,In_1320,In_2065);
nor U950 (N_950,In_180,In_2824);
nand U951 (N_951,In_458,In_1226);
nand U952 (N_952,In_2541,In_589);
or U953 (N_953,In_1079,In_737);
nand U954 (N_954,In_1155,In_2792);
and U955 (N_955,In_525,In_1025);
or U956 (N_956,In_2023,In_1032);
or U957 (N_957,In_976,In_803);
nand U958 (N_958,In_1260,In_707);
and U959 (N_959,In_1170,In_278);
or U960 (N_960,In_287,In_454);
and U961 (N_961,In_2107,In_908);
xnor U962 (N_962,In_326,In_866);
and U963 (N_963,In_1289,In_2310);
nor U964 (N_964,In_1516,In_533);
nor U965 (N_965,In_1262,In_1270);
nor U966 (N_966,In_282,In_1166);
nor U967 (N_967,In_2714,In_1218);
and U968 (N_968,In_602,In_936);
and U969 (N_969,In_2770,In_179);
or U970 (N_970,In_459,In_95);
nor U971 (N_971,In_1911,In_531);
or U972 (N_972,In_203,In_656);
xnor U973 (N_973,In_687,In_1534);
nor U974 (N_974,In_2325,In_1015);
xnor U975 (N_975,In_2671,In_1545);
or U976 (N_976,In_1031,In_543);
nor U977 (N_977,In_2254,In_1759);
or U978 (N_978,In_1304,In_2593);
nor U979 (N_979,In_749,In_1687);
nor U980 (N_980,In_2666,In_2077);
nand U981 (N_981,In_2098,In_2751);
and U982 (N_982,In_1368,In_2640);
nor U983 (N_983,In_293,In_2734);
nor U984 (N_984,In_1098,In_1043);
xor U985 (N_985,In_954,In_926);
or U986 (N_986,In_2286,In_240);
nor U987 (N_987,In_2976,In_2756);
nor U988 (N_988,In_2916,In_811);
or U989 (N_989,In_258,In_692);
and U990 (N_990,In_1255,In_1386);
nor U991 (N_991,In_2980,In_160);
and U992 (N_992,In_1109,In_1699);
and U993 (N_993,In_517,In_2923);
nand U994 (N_994,In_344,In_1139);
nand U995 (N_995,In_2624,In_1332);
or U996 (N_996,In_2097,In_1456);
xor U997 (N_997,In_197,In_1789);
and U998 (N_998,In_586,In_244);
nor U999 (N_999,In_2187,In_2282);
nor U1000 (N_1000,In_2620,In_1452);
or U1001 (N_1001,In_911,In_2197);
nor U1002 (N_1002,In_39,In_2782);
nand U1003 (N_1003,In_469,In_626);
xor U1004 (N_1004,In_2370,In_464);
nor U1005 (N_1005,In_2200,In_2376);
and U1006 (N_1006,In_1209,In_1644);
xor U1007 (N_1007,In_1416,In_2474);
xnor U1008 (N_1008,In_387,In_303);
or U1009 (N_1009,In_2811,In_1417);
nand U1010 (N_1010,In_895,In_940);
nand U1011 (N_1011,In_509,In_640);
or U1012 (N_1012,In_1112,In_2222);
nor U1013 (N_1013,In_1637,In_2600);
nor U1014 (N_1014,In_741,In_744);
nand U1015 (N_1015,In_2711,In_2218);
nand U1016 (N_1016,In_2147,In_1861);
xor U1017 (N_1017,In_1626,In_535);
xor U1018 (N_1018,In_2156,In_1454);
nand U1019 (N_1019,In_2398,In_1334);
nand U1020 (N_1020,In_253,In_32);
and U1021 (N_1021,In_416,In_75);
nand U1022 (N_1022,In_1604,In_1008);
nor U1023 (N_1023,In_1367,In_229);
xnor U1024 (N_1024,In_138,In_342);
xnor U1025 (N_1025,In_403,In_2848);
nand U1026 (N_1026,In_429,In_1955);
nor U1027 (N_1027,In_2979,In_1624);
or U1028 (N_1028,In_1549,In_1827);
nand U1029 (N_1029,In_1680,In_1595);
nor U1030 (N_1030,In_1438,In_2079);
and U1031 (N_1031,In_2093,In_2748);
nor U1032 (N_1032,In_434,In_587);
and U1033 (N_1033,In_2284,In_2965);
nor U1034 (N_1034,In_443,In_1522);
nor U1035 (N_1035,In_746,In_1343);
nor U1036 (N_1036,In_1890,In_2175);
or U1037 (N_1037,In_655,In_2658);
or U1038 (N_1038,In_717,In_2244);
xor U1039 (N_1039,In_2708,In_1669);
xnor U1040 (N_1040,In_1723,In_1253);
or U1041 (N_1041,In_211,In_2709);
or U1042 (N_1042,In_1121,In_2892);
nor U1043 (N_1043,In_2418,In_498);
or U1044 (N_1044,In_1769,In_934);
or U1045 (N_1045,In_196,In_682);
or U1046 (N_1046,In_2795,In_863);
nand U1047 (N_1047,In_852,In_1814);
or U1048 (N_1048,In_1161,In_175);
or U1049 (N_1049,In_496,In_748);
nor U1050 (N_1050,In_2184,In_1003);
xor U1051 (N_1051,In_200,In_219);
nand U1052 (N_1052,In_296,In_600);
nand U1053 (N_1053,In_2314,In_2000);
nor U1054 (N_1054,In_144,In_2081);
or U1055 (N_1055,In_2723,In_2400);
xor U1056 (N_1056,In_1882,In_492);
and U1057 (N_1057,In_972,In_779);
nand U1058 (N_1058,In_2874,In_616);
nand U1059 (N_1059,In_1429,In_1640);
nand U1060 (N_1060,In_864,In_1099);
xnor U1061 (N_1061,In_2260,In_553);
and U1062 (N_1062,In_1269,In_1933);
nand U1063 (N_1063,In_1733,In_2039);
nand U1064 (N_1064,In_2139,In_1995);
or U1065 (N_1065,In_1817,In_959);
or U1066 (N_1066,In_983,In_1562);
nor U1067 (N_1067,In_2942,In_1930);
nand U1068 (N_1068,In_2816,In_1826);
nor U1069 (N_1069,In_2135,In_2661);
xor U1070 (N_1070,In_2290,In_2493);
nor U1071 (N_1071,In_2764,In_202);
and U1072 (N_1072,In_311,In_313);
nand U1073 (N_1073,In_1635,In_101);
nor U1074 (N_1074,In_2382,In_1129);
or U1075 (N_1075,In_544,In_2397);
nand U1076 (N_1076,In_946,In_2940);
or U1077 (N_1077,In_2410,In_1047);
nor U1078 (N_1078,In_308,In_92);
and U1079 (N_1079,In_1038,In_97);
or U1080 (N_1080,In_1152,In_1638);
nand U1081 (N_1081,In_2961,In_2415);
nand U1082 (N_1082,In_20,In_486);
nor U1083 (N_1083,In_790,In_2386);
nor U1084 (N_1084,In_230,In_1570);
and U1085 (N_1085,In_1093,In_1486);
nor U1086 (N_1086,In_2148,In_716);
nand U1087 (N_1087,In_2645,In_2908);
nor U1088 (N_1088,In_280,In_2346);
nand U1089 (N_1089,In_246,In_1807);
nor U1090 (N_1090,In_705,In_1147);
and U1091 (N_1091,In_1303,In_912);
or U1092 (N_1092,In_712,In_2126);
or U1093 (N_1093,In_2614,In_1033);
and U1094 (N_1094,In_1656,In_918);
xnor U1095 (N_1095,In_743,In_2168);
or U1096 (N_1096,In_627,In_474);
and U1097 (N_1097,In_355,In_792);
xnor U1098 (N_1098,In_599,In_706);
nand U1099 (N_1099,In_2753,In_2240);
xnor U1100 (N_1100,In_2118,In_2267);
nand U1101 (N_1101,In_68,In_993);
or U1102 (N_1102,In_91,In_2969);
xnor U1103 (N_1103,In_2576,In_111);
nand U1104 (N_1104,In_1748,In_2568);
or U1105 (N_1105,In_2336,In_106);
nand U1106 (N_1106,In_1291,In_1894);
nand U1107 (N_1107,In_1772,In_900);
or U1108 (N_1108,In_194,In_317);
and U1109 (N_1109,In_2685,In_2043);
or U1110 (N_1110,In_2106,In_1383);
nand U1111 (N_1111,In_1265,In_2164);
nor U1112 (N_1112,In_1192,In_2856);
and U1113 (N_1113,In_1548,In_2056);
and U1114 (N_1114,In_81,In_1191);
xor U1115 (N_1115,In_1564,In_1856);
nand U1116 (N_1116,In_206,In_415);
xor U1117 (N_1117,In_1862,In_1938);
nor U1118 (N_1118,In_2973,In_667);
nand U1119 (N_1119,In_1279,In_322);
nor U1120 (N_1120,In_186,In_1838);
and U1121 (N_1121,In_572,In_1118);
xor U1122 (N_1122,In_534,In_518);
xor U1123 (N_1123,In_1627,In_493);
or U1124 (N_1124,In_90,In_881);
nand U1125 (N_1125,In_1540,In_151);
and U1126 (N_1126,In_409,In_418);
or U1127 (N_1127,In_1510,In_1497);
nor U1128 (N_1128,In_1664,In_715);
nand U1129 (N_1129,In_2759,In_636);
nand U1130 (N_1130,In_916,In_2334);
nand U1131 (N_1131,In_1994,In_1670);
xnor U1132 (N_1132,In_1431,In_2239);
nor U1133 (N_1133,In_408,In_1);
and U1134 (N_1134,In_1892,In_2297);
and U1135 (N_1135,In_1953,In_2919);
xnor U1136 (N_1136,In_2340,In_686);
xor U1137 (N_1137,In_1805,In_225);
or U1138 (N_1138,In_1785,In_2379);
xor U1139 (N_1139,In_2629,In_1309);
and U1140 (N_1140,In_2227,In_2332);
and U1141 (N_1141,In_1163,In_2799);
nor U1142 (N_1142,In_830,In_1203);
or U1143 (N_1143,In_2145,In_1151);
xor U1144 (N_1144,In_582,In_1168);
xnor U1145 (N_1145,In_2689,In_1959);
nor U1146 (N_1146,In_1323,In_2232);
nand U1147 (N_1147,In_797,In_938);
xnor U1148 (N_1148,In_1211,In_1900);
and U1149 (N_1149,In_1823,In_2721);
and U1150 (N_1150,In_791,In_1612);
or U1151 (N_1151,In_1131,In_514);
or U1152 (N_1152,In_1709,In_1542);
nor U1153 (N_1153,In_1104,In_96);
xor U1154 (N_1154,In_628,In_1992);
nand U1155 (N_1155,In_57,In_1822);
nor U1156 (N_1156,In_1906,In_468);
and U1157 (N_1157,In_1247,In_235);
nor U1158 (N_1158,In_1547,In_398);
nor U1159 (N_1159,In_2160,In_370);
nand U1160 (N_1160,In_248,In_371);
nor U1161 (N_1161,In_1579,In_635);
nor U1162 (N_1162,In_1658,In_265);
or U1163 (N_1163,In_1878,In_2048);
or U1164 (N_1164,In_2758,In_1746);
or U1165 (N_1165,In_1590,In_730);
xor U1166 (N_1166,In_2760,In_1287);
and U1167 (N_1167,In_822,In_840);
or U1168 (N_1168,In_2914,In_1428);
xnor U1169 (N_1169,In_15,In_2997);
or U1170 (N_1170,In_1574,In_2015);
nand U1171 (N_1171,In_955,In_1678);
xnor U1172 (N_1172,In_2554,In_2930);
xnor U1173 (N_1173,In_2796,In_473);
and U1174 (N_1174,In_939,In_760);
nand U1175 (N_1175,In_1207,In_2632);
and U1176 (N_1176,In_774,In_2728);
xnor U1177 (N_1177,In_2665,In_2236);
nand U1178 (N_1178,In_2405,In_904);
or U1179 (N_1179,In_1734,In_2594);
nor U1180 (N_1180,In_2321,In_2502);
nor U1181 (N_1181,In_1280,In_1899);
and U1182 (N_1182,In_2089,In_2237);
and U1183 (N_1183,In_59,In_38);
nor U1184 (N_1184,In_786,In_1331);
xnor U1185 (N_1185,In_538,In_1437);
or U1186 (N_1186,In_819,In_1230);
nand U1187 (N_1187,In_571,In_2897);
xnor U1188 (N_1188,In_1711,In_1982);
nand U1189 (N_1189,In_1016,In_2778);
xor U1190 (N_1190,In_113,In_694);
nor U1191 (N_1191,In_2465,In_2074);
xnor U1192 (N_1192,In_2208,In_2201);
or U1193 (N_1193,In_1651,In_1349);
or U1194 (N_1194,In_1500,In_1201);
nand U1195 (N_1195,In_2837,In_2507);
xor U1196 (N_1196,In_2938,In_2047);
and U1197 (N_1197,In_2757,In_2510);
nor U1198 (N_1198,In_1697,In_1125);
nand U1199 (N_1199,In_1019,In_1488);
and U1200 (N_1200,In_1617,In_524);
and U1201 (N_1201,In_1921,In_2121);
nor U1202 (N_1202,In_1282,In_367);
or U1203 (N_1203,In_2978,In_2262);
xnor U1204 (N_1204,In_107,In_963);
and U1205 (N_1205,In_714,In_1359);
or U1206 (N_1206,In_64,In_2743);
and U1207 (N_1207,In_1704,In_893);
nor U1208 (N_1208,In_1465,In_2700);
xnor U1209 (N_1209,In_1957,In_1778);
xor U1210 (N_1210,In_800,In_2663);
or U1211 (N_1211,In_1065,In_752);
and U1212 (N_1212,In_1106,In_2578);
xnor U1213 (N_1213,In_2699,In_1968);
xor U1214 (N_1214,In_1874,In_430);
and U1215 (N_1215,In_643,In_2905);
and U1216 (N_1216,In_34,In_1434);
and U1217 (N_1217,In_2994,In_930);
nor U1218 (N_1218,In_1243,In_1186);
nor U1219 (N_1219,In_136,In_134);
or U1220 (N_1220,In_824,In_1876);
nor U1221 (N_1221,In_1741,In_1388);
xnor U1222 (N_1222,In_467,In_2406);
nor U1223 (N_1223,In_1135,In_2694);
or U1224 (N_1224,In_117,In_1216);
xor U1225 (N_1225,In_1337,In_268);
nor U1226 (N_1226,In_1445,In_294);
xnor U1227 (N_1227,In_2907,In_1795);
and U1228 (N_1228,In_510,In_1346);
nor U1229 (N_1229,In_1143,In_1632);
and U1230 (N_1230,In_718,In_2746);
nand U1231 (N_1231,In_2686,In_1887);
and U1232 (N_1232,In_1067,In_2005);
nor U1233 (N_1233,In_489,In_2289);
nor U1234 (N_1234,In_1736,In_1450);
or U1235 (N_1235,In_450,In_2167);
xor U1236 (N_1236,In_2787,In_2491);
xnor U1237 (N_1237,In_2900,In_619);
nor U1238 (N_1238,In_2545,In_2230);
nand U1239 (N_1239,In_1619,In_841);
and U1240 (N_1240,In_88,In_1830);
xnor U1241 (N_1241,In_2296,In_132);
and U1242 (N_1242,In_2104,In_2904);
nor U1243 (N_1243,In_914,In_1138);
and U1244 (N_1244,In_2363,In_1039);
nand U1245 (N_1245,In_2475,In_272);
nor U1246 (N_1246,In_1820,In_85);
nor U1247 (N_1247,In_787,In_660);
or U1248 (N_1248,In_1180,In_80);
and U1249 (N_1249,In_2983,In_719);
nand U1250 (N_1250,In_1834,In_2226);
and U1251 (N_1251,In_1803,In_14);
nor U1252 (N_1252,In_2855,In_491);
nand U1253 (N_1253,In_1224,In_1507);
nand U1254 (N_1254,In_157,In_796);
or U1255 (N_1255,In_1609,In_1573);
xnor U1256 (N_1256,In_381,In_897);
nor U1257 (N_1257,In_615,In_1690);
nor U1258 (N_1258,In_929,In_22);
nor U1259 (N_1259,In_1952,In_848);
xor U1260 (N_1260,In_2909,In_1220);
nor U1261 (N_1261,In_241,In_1877);
and U1262 (N_1262,In_927,In_2407);
xor U1263 (N_1263,In_163,In_826);
xor U1264 (N_1264,In_487,In_1965);
and U1265 (N_1265,In_2884,In_2744);
and U1266 (N_1266,In_624,In_520);
xnor U1267 (N_1267,In_2412,In_171);
or U1268 (N_1268,In_2018,In_2506);
and U1269 (N_1269,In_380,In_1449);
nand U1270 (N_1270,In_2776,In_2360);
xnor U1271 (N_1271,In_2547,In_2834);
and U1272 (N_1272,In_2062,In_2522);
xnor U1273 (N_1273,In_437,In_1116);
xnor U1274 (N_1274,In_1813,In_855);
nor U1275 (N_1275,In_2602,In_328);
xnor U1276 (N_1276,In_2202,In_2303);
xor U1277 (N_1277,In_1646,In_2505);
and U1278 (N_1278,In_360,In_479);
nand U1279 (N_1279,In_1603,In_1863);
nand U1280 (N_1280,In_598,In_1543);
nand U1281 (N_1281,In_2461,In_105);
xor U1282 (N_1282,In_2668,In_1041);
and U1283 (N_1283,In_428,In_2450);
or U1284 (N_1284,In_1355,In_1735);
nor U1285 (N_1285,In_1630,In_2025);
nand U1286 (N_1286,In_1199,In_953);
xnor U1287 (N_1287,In_2987,In_2608);
nor U1288 (N_1288,In_73,In_116);
nor U1289 (N_1289,In_2518,In_2736);
nand U1290 (N_1290,In_71,In_146);
or U1291 (N_1291,In_436,In_503);
or U1292 (N_1292,In_727,In_1490);
and U1293 (N_1293,In_2040,In_2210);
and U1294 (N_1294,In_1999,In_405);
nor U1295 (N_1295,In_1492,In_1611);
and U1296 (N_1296,In_2477,In_1743);
nand U1297 (N_1297,In_1302,In_2265);
or U1298 (N_1298,In_915,In_2393);
nand U1299 (N_1299,In_242,In_591);
or U1300 (N_1300,In_2174,In_1731);
xor U1301 (N_1301,In_89,In_421);
or U1302 (N_1302,In_1514,In_761);
nor U1303 (N_1303,In_1413,In_1271);
nand U1304 (N_1304,In_386,In_2182);
xnor U1305 (N_1305,In_1137,In_2528);
nand U1306 (N_1306,In_1341,In_1529);
or U1307 (N_1307,In_631,In_2252);
and U1308 (N_1308,In_448,In_609);
and U1309 (N_1309,In_1550,In_1784);
nor U1310 (N_1310,In_1527,In_1470);
nor U1311 (N_1311,In_2949,In_60);
xnor U1312 (N_1312,In_1653,In_1541);
or U1313 (N_1313,In_770,In_2860);
xnor U1314 (N_1314,In_129,In_597);
xor U1315 (N_1315,In_226,In_1110);
xor U1316 (N_1316,In_1833,In_1685);
xnor U1317 (N_1317,In_1108,In_2752);
nand U1318 (N_1318,In_1631,In_842);
and U1319 (N_1319,In_1113,In_453);
nand U1320 (N_1320,In_1976,In_1963);
xor U1321 (N_1321,In_378,In_1018);
or U1322 (N_1322,In_952,In_16);
nand U1323 (N_1323,In_2910,In_1153);
or U1324 (N_1324,In_1844,In_41);
and U1325 (N_1325,In_795,In_2880);
or U1326 (N_1326,In_2710,In_2802);
nand U1327 (N_1327,In_2864,In_1973);
xnor U1328 (N_1328,In_1362,In_1310);
nor U1329 (N_1329,In_2307,In_1315);
nand U1330 (N_1330,In_2490,In_989);
and U1331 (N_1331,In_964,In_1034);
nor U1332 (N_1332,In_1519,In_799);
xor U1333 (N_1333,In_2384,In_2604);
xnor U1334 (N_1334,In_1241,In_843);
nand U1335 (N_1335,In_147,In_1300);
or U1336 (N_1336,In_1223,In_1095);
and U1337 (N_1337,In_1928,In_1020);
nand U1338 (N_1338,In_2830,In_406);
or U1339 (N_1339,In_1142,In_1078);
nor U1340 (N_1340,In_751,In_2876);
or U1341 (N_1341,In_554,In_1531);
nor U1342 (N_1342,In_1185,In_995);
nand U1343 (N_1343,In_2463,In_2103);
nand U1344 (N_1344,In_1623,In_2447);
nor U1345 (N_1345,In_2399,In_2672);
and U1346 (N_1346,In_44,In_2319);
nand U1347 (N_1347,In_2007,In_762);
xnor U1348 (N_1348,In_1588,In_396);
nand U1349 (N_1349,In_1114,In_382);
or U1350 (N_1350,In_1074,In_1537);
and U1351 (N_1351,In_1504,In_2478);
nor U1352 (N_1352,In_652,In_1764);
xnor U1353 (N_1353,In_2870,In_768);
xnor U1354 (N_1354,In_37,In_2859);
or U1355 (N_1355,In_1556,In_1290);
nor U1356 (N_1356,In_1494,In_1081);
nand U1357 (N_1357,In_1101,In_549);
nand U1358 (N_1358,In_1964,In_2377);
or U1359 (N_1359,In_2058,In_1586);
or U1360 (N_1360,In_2171,In_2688);
and U1361 (N_1361,In_2726,In_2357);
nand U1362 (N_1362,In_807,In_858);
xor U1363 (N_1363,In_2096,In_19);
and U1364 (N_1364,In_2981,In_438);
nor U1365 (N_1365,In_465,In_722);
nor U1366 (N_1366,In_558,In_2022);
or U1367 (N_1367,In_2768,In_2026);
nor U1368 (N_1368,In_2009,In_1601);
and U1369 (N_1369,In_1503,In_1800);
nor U1370 (N_1370,In_358,In_1328);
nand U1371 (N_1371,In_879,In_1700);
and U1372 (N_1372,In_324,In_338);
nand U1373 (N_1373,In_291,In_343);
or U1374 (N_1374,In_2737,In_906);
and U1375 (N_1375,In_463,In_397);
xnor U1376 (N_1376,In_2990,In_79);
and U1377 (N_1377,In_2509,In_546);
or U1378 (N_1378,In_1859,In_2820);
nor U1379 (N_1379,In_2395,In_1568);
nand U1380 (N_1380,In_2177,In_2353);
nor U1381 (N_1381,In_1422,In_2956);
or U1382 (N_1382,In_2113,In_1526);
and U1383 (N_1383,In_1944,In_306);
or U1384 (N_1384,In_1234,In_1993);
xor U1385 (N_1385,In_2566,In_46);
or U1386 (N_1386,In_1983,In_2283);
nor U1387 (N_1387,In_2695,In_1682);
or U1388 (N_1388,In_967,In_2972);
nand U1389 (N_1389,In_1781,In_2437);
nand U1390 (N_1390,In_1674,In_867);
nand U1391 (N_1391,In_2877,In_2301);
or U1392 (N_1392,In_2069,In_2063);
and U1393 (N_1393,In_262,In_2374);
nor U1394 (N_1394,In_2435,In_2115);
and U1395 (N_1395,In_192,In_1591);
nand U1396 (N_1396,In_1655,In_2570);
and U1397 (N_1397,In_2832,In_878);
or U1398 (N_1398,In_2143,In_1054);
nor U1399 (N_1399,In_2331,In_2454);
nand U1400 (N_1400,In_1596,In_1897);
and U1401 (N_1401,In_2101,In_2932);
and U1402 (N_1402,In_1178,In_2717);
or U1403 (N_1403,In_2605,In_2271);
and U1404 (N_1404,In_1119,In_2857);
or U1405 (N_1405,In_578,In_704);
xor U1406 (N_1406,In_935,In_93);
nand U1407 (N_1407,In_441,In_2698);
or U1408 (N_1408,In_2159,In_710);
nand U1409 (N_1409,In_2345,In_2819);
or U1410 (N_1410,In_1715,In_1083);
or U1411 (N_1411,In_310,In_1053);
and U1412 (N_1412,In_1917,In_516);
or U1413 (N_1413,In_2835,In_2059);
or U1414 (N_1414,In_2934,In_1857);
or U1415 (N_1415,In_2881,In_2211);
nor U1416 (N_1416,In_1872,In_2971);
or U1417 (N_1417,In_1393,In_390);
xor U1418 (N_1418,In_951,In_2085);
xnor U1419 (N_1419,In_1407,In_2010);
nor U1420 (N_1420,In_1017,In_2339);
xnor U1421 (N_1421,In_1691,In_2055);
nand U1422 (N_1422,In_2808,In_267);
or U1423 (N_1423,In_2954,In_2195);
and U1424 (N_1424,In_1453,In_2110);
or U1425 (N_1425,In_2203,In_471);
xor U1426 (N_1426,In_2867,In_829);
and U1427 (N_1427,In_821,In_1628);
or U1428 (N_1428,In_1958,In_2432);
nor U1429 (N_1429,In_337,In_298);
nand U1430 (N_1430,In_1645,In_973);
or U1431 (N_1431,In_1171,In_882);
nor U1432 (N_1432,In_802,In_417);
and U1433 (N_1433,In_1849,In_2650);
xor U1434 (N_1434,In_1384,In_1213);
nor U1435 (N_1435,In_389,In_1379);
nand U1436 (N_1436,In_2913,In_648);
or U1437 (N_1437,In_99,In_1028);
or U1438 (N_1438,In_1918,In_1696);
nand U1439 (N_1439,In_2337,In_26);
or U1440 (N_1440,In_1945,In_2199);
and U1441 (N_1441,In_2404,In_1350);
and U1442 (N_1442,In_2392,In_2609);
or U1443 (N_1443,In_1439,In_2822);
and U1444 (N_1444,In_18,In_532);
or U1445 (N_1445,In_1297,In_130);
xnor U1446 (N_1446,In_21,In_2921);
xnor U1447 (N_1447,In_2551,In_1871);
or U1448 (N_1448,In_2487,In_2114);
nand U1449 (N_1449,In_2045,In_539);
nand U1450 (N_1450,In_1314,In_2625);
xnor U1451 (N_1451,In_657,In_2706);
or U1452 (N_1452,In_1981,In_568);
or U1453 (N_1453,In_868,In_764);
xnor U1454 (N_1454,In_494,In_1024);
or U1455 (N_1455,In_1404,In_152);
and U1456 (N_1456,In_1200,In_1879);
nand U1457 (N_1457,In_1474,In_201);
nand U1458 (N_1458,In_755,In_2049);
xnor U1459 (N_1459,In_2947,In_721);
or U1460 (N_1460,In_1377,In_114);
xor U1461 (N_1461,In_537,In_2902);
nor U1462 (N_1462,In_28,In_1040);
xnor U1463 (N_1463,In_2338,In_2996);
nand U1464 (N_1464,In_1956,In_1728);
nand U1465 (N_1465,In_1641,In_1082);
nand U1466 (N_1466,In_2654,In_1773);
nand U1467 (N_1467,In_547,In_1401);
and U1468 (N_1468,In_170,In_45);
or U1469 (N_1469,In_1798,In_2312);
or U1470 (N_1470,In_1410,In_2102);
or U1471 (N_1471,In_2070,In_2853);
xnor U1472 (N_1472,In_680,In_1977);
or U1473 (N_1473,In_2046,In_671);
xor U1474 (N_1474,In_149,In_613);
or U1475 (N_1475,In_198,In_2146);
nor U1476 (N_1476,In_2667,In_2610);
nand U1477 (N_1477,In_2929,In_339);
xnor U1478 (N_1478,In_917,In_1487);
or U1479 (N_1479,In_2573,In_2815);
nor U1480 (N_1480,In_1902,In_2031);
xor U1481 (N_1481,In_2571,In_1559);
nor U1482 (N_1482,In_411,In_2955);
and U1483 (N_1483,In_1154,In_2383);
nand U1484 (N_1484,In_877,In_854);
nor U1485 (N_1485,In_2817,In_1513);
and U1486 (N_1486,In_2351,In_118);
and U1487 (N_1487,In_2563,In_666);
nor U1488 (N_1488,In_1318,In_2439);
xor U1489 (N_1489,In_1195,In_1292);
and U1490 (N_1490,In_1102,In_1374);
or U1491 (N_1491,In_1898,In_576);
nor U1492 (N_1492,In_1650,In_1960);
nor U1493 (N_1493,In_2989,In_1719);
and U1494 (N_1494,In_1621,In_603);
xor U1495 (N_1495,In_1625,In_2975);
nand U1496 (N_1496,In_1369,In_1244);
or U1497 (N_1497,In_2234,In_2273);
xnor U1498 (N_1498,In_2037,In_775);
nand U1499 (N_1499,In_220,In_1479);
and U1500 (N_1500,In_946,In_1100);
nor U1501 (N_1501,In_1322,In_649);
xnor U1502 (N_1502,In_2861,In_2758);
nand U1503 (N_1503,In_2882,In_2493);
and U1504 (N_1504,In_2053,In_877);
or U1505 (N_1505,In_622,In_761);
xor U1506 (N_1506,In_1998,In_598);
nor U1507 (N_1507,In_2098,In_1373);
and U1508 (N_1508,In_1437,In_1852);
xnor U1509 (N_1509,In_2108,In_1839);
xnor U1510 (N_1510,In_996,In_566);
nor U1511 (N_1511,In_400,In_1713);
or U1512 (N_1512,In_2835,In_1007);
xnor U1513 (N_1513,In_1335,In_2483);
or U1514 (N_1514,In_398,In_2469);
nand U1515 (N_1515,In_2746,In_941);
nand U1516 (N_1516,In_343,In_802);
or U1517 (N_1517,In_295,In_1102);
and U1518 (N_1518,In_2826,In_1135);
nand U1519 (N_1519,In_2025,In_581);
nor U1520 (N_1520,In_970,In_2490);
nand U1521 (N_1521,In_286,In_2648);
and U1522 (N_1522,In_2865,In_910);
xnor U1523 (N_1523,In_1299,In_1789);
nor U1524 (N_1524,In_1267,In_2481);
nand U1525 (N_1525,In_852,In_891);
or U1526 (N_1526,In_406,In_2347);
xnor U1527 (N_1527,In_2341,In_2764);
and U1528 (N_1528,In_287,In_889);
and U1529 (N_1529,In_1655,In_1459);
nand U1530 (N_1530,In_2149,In_315);
and U1531 (N_1531,In_1031,In_261);
or U1532 (N_1532,In_2599,In_235);
or U1533 (N_1533,In_2717,In_2392);
nor U1534 (N_1534,In_1144,In_952);
xnor U1535 (N_1535,In_1540,In_1170);
and U1536 (N_1536,In_2500,In_2209);
nor U1537 (N_1537,In_1051,In_439);
and U1538 (N_1538,In_545,In_1267);
and U1539 (N_1539,In_303,In_1529);
and U1540 (N_1540,In_1451,In_2412);
xnor U1541 (N_1541,In_2983,In_1285);
and U1542 (N_1542,In_2352,In_479);
or U1543 (N_1543,In_587,In_928);
nor U1544 (N_1544,In_1079,In_2969);
nand U1545 (N_1545,In_1862,In_824);
nand U1546 (N_1546,In_1664,In_983);
nor U1547 (N_1547,In_1642,In_187);
and U1548 (N_1548,In_226,In_2576);
nand U1549 (N_1549,In_472,In_1861);
and U1550 (N_1550,In_2384,In_2991);
nor U1551 (N_1551,In_2258,In_615);
or U1552 (N_1552,In_1285,In_1120);
or U1553 (N_1553,In_92,In_477);
nand U1554 (N_1554,In_1679,In_231);
xor U1555 (N_1555,In_1551,In_1414);
nand U1556 (N_1556,In_2537,In_2469);
nand U1557 (N_1557,In_1644,In_1254);
xnor U1558 (N_1558,In_2839,In_634);
nor U1559 (N_1559,In_617,In_672);
and U1560 (N_1560,In_1832,In_1062);
and U1561 (N_1561,In_2366,In_1381);
and U1562 (N_1562,In_1495,In_1374);
xor U1563 (N_1563,In_184,In_2278);
nand U1564 (N_1564,In_2988,In_767);
nand U1565 (N_1565,In_1307,In_1047);
and U1566 (N_1566,In_1429,In_276);
nor U1567 (N_1567,In_1537,In_2011);
nand U1568 (N_1568,In_407,In_762);
xnor U1569 (N_1569,In_1760,In_2145);
nor U1570 (N_1570,In_1499,In_1928);
nor U1571 (N_1571,In_1418,In_2582);
nor U1572 (N_1572,In_335,In_1294);
or U1573 (N_1573,In_2467,In_1732);
nor U1574 (N_1574,In_1423,In_2228);
xor U1575 (N_1575,In_2513,In_1941);
nand U1576 (N_1576,In_841,In_1651);
nor U1577 (N_1577,In_437,In_1579);
nor U1578 (N_1578,In_1188,In_2832);
xnor U1579 (N_1579,In_111,In_1144);
or U1580 (N_1580,In_582,In_69);
or U1581 (N_1581,In_1292,In_2806);
or U1582 (N_1582,In_1220,In_1103);
or U1583 (N_1583,In_2832,In_432);
and U1584 (N_1584,In_1072,In_1750);
nand U1585 (N_1585,In_175,In_1420);
or U1586 (N_1586,In_821,In_2457);
or U1587 (N_1587,In_1092,In_2974);
nand U1588 (N_1588,In_1092,In_800);
nand U1589 (N_1589,In_2228,In_2071);
xnor U1590 (N_1590,In_857,In_1029);
and U1591 (N_1591,In_2519,In_296);
xnor U1592 (N_1592,In_1927,In_356);
xor U1593 (N_1593,In_1868,In_1867);
or U1594 (N_1594,In_385,In_13);
and U1595 (N_1595,In_1886,In_2237);
and U1596 (N_1596,In_1915,In_1445);
or U1597 (N_1597,In_1414,In_1062);
or U1598 (N_1598,In_2138,In_2803);
nand U1599 (N_1599,In_1131,In_2209);
nand U1600 (N_1600,In_2116,In_115);
nand U1601 (N_1601,In_2147,In_624);
and U1602 (N_1602,In_963,In_603);
nor U1603 (N_1603,In_2840,In_1649);
and U1604 (N_1604,In_950,In_2353);
nor U1605 (N_1605,In_883,In_1115);
and U1606 (N_1606,In_2183,In_1527);
and U1607 (N_1607,In_2600,In_1717);
nor U1608 (N_1608,In_446,In_2721);
nor U1609 (N_1609,In_1735,In_1790);
and U1610 (N_1610,In_1087,In_2565);
nand U1611 (N_1611,In_2882,In_558);
nor U1612 (N_1612,In_2106,In_1774);
xor U1613 (N_1613,In_1427,In_162);
nor U1614 (N_1614,In_1691,In_2840);
nor U1615 (N_1615,In_2439,In_587);
nor U1616 (N_1616,In_2540,In_643);
nor U1617 (N_1617,In_2814,In_195);
and U1618 (N_1618,In_2294,In_2819);
and U1619 (N_1619,In_2316,In_783);
nor U1620 (N_1620,In_2320,In_2554);
or U1621 (N_1621,In_2129,In_1973);
nand U1622 (N_1622,In_1326,In_1950);
or U1623 (N_1623,In_1031,In_504);
or U1624 (N_1624,In_2113,In_2908);
xnor U1625 (N_1625,In_1531,In_2047);
or U1626 (N_1626,In_1009,In_1213);
or U1627 (N_1627,In_2330,In_2688);
xnor U1628 (N_1628,In_192,In_2258);
nor U1629 (N_1629,In_2897,In_2551);
and U1630 (N_1630,In_138,In_1004);
and U1631 (N_1631,In_834,In_807);
nand U1632 (N_1632,In_1535,In_1189);
nand U1633 (N_1633,In_1432,In_1035);
or U1634 (N_1634,In_1583,In_1030);
xnor U1635 (N_1635,In_2075,In_205);
xnor U1636 (N_1636,In_469,In_2781);
and U1637 (N_1637,In_1282,In_164);
or U1638 (N_1638,In_469,In_1680);
and U1639 (N_1639,In_1591,In_1211);
nor U1640 (N_1640,In_2609,In_404);
and U1641 (N_1641,In_1305,In_342);
nand U1642 (N_1642,In_1669,In_2655);
xor U1643 (N_1643,In_996,In_2093);
nor U1644 (N_1644,In_252,In_332);
and U1645 (N_1645,In_1862,In_2651);
and U1646 (N_1646,In_790,In_2731);
nand U1647 (N_1647,In_2019,In_2642);
and U1648 (N_1648,In_1986,In_2119);
xor U1649 (N_1649,In_2314,In_2202);
or U1650 (N_1650,In_2245,In_1145);
or U1651 (N_1651,In_2668,In_929);
nand U1652 (N_1652,In_1378,In_1233);
and U1653 (N_1653,In_2866,In_2791);
nand U1654 (N_1654,In_1138,In_1817);
nor U1655 (N_1655,In_1994,In_2037);
nor U1656 (N_1656,In_2273,In_1306);
nand U1657 (N_1657,In_1450,In_2899);
nand U1658 (N_1658,In_2227,In_1640);
nor U1659 (N_1659,In_2693,In_1221);
nand U1660 (N_1660,In_2809,In_2844);
xnor U1661 (N_1661,In_641,In_252);
and U1662 (N_1662,In_1981,In_2387);
nor U1663 (N_1663,In_2532,In_1972);
and U1664 (N_1664,In_2689,In_1252);
or U1665 (N_1665,In_389,In_2374);
nor U1666 (N_1666,In_2413,In_1631);
xnor U1667 (N_1667,In_1988,In_2397);
and U1668 (N_1668,In_1182,In_960);
and U1669 (N_1669,In_640,In_1951);
and U1670 (N_1670,In_2771,In_1211);
xnor U1671 (N_1671,In_829,In_922);
and U1672 (N_1672,In_1858,In_2438);
nor U1673 (N_1673,In_725,In_1715);
or U1674 (N_1674,In_341,In_716);
xor U1675 (N_1675,In_964,In_868);
xnor U1676 (N_1676,In_2679,In_1892);
or U1677 (N_1677,In_2562,In_1701);
nand U1678 (N_1678,In_1406,In_2709);
nand U1679 (N_1679,In_212,In_466);
and U1680 (N_1680,In_2431,In_1136);
nor U1681 (N_1681,In_2744,In_551);
xor U1682 (N_1682,In_2995,In_2412);
nand U1683 (N_1683,In_831,In_664);
xor U1684 (N_1684,In_646,In_108);
nor U1685 (N_1685,In_1771,In_281);
and U1686 (N_1686,In_2739,In_2980);
or U1687 (N_1687,In_2359,In_2130);
or U1688 (N_1688,In_2090,In_2193);
and U1689 (N_1689,In_1316,In_1954);
or U1690 (N_1690,In_1845,In_1218);
or U1691 (N_1691,In_854,In_482);
or U1692 (N_1692,In_2310,In_860);
xnor U1693 (N_1693,In_388,In_938);
nor U1694 (N_1694,In_1735,In_2805);
and U1695 (N_1695,In_868,In_921);
nor U1696 (N_1696,In_2050,In_2778);
xor U1697 (N_1697,In_2472,In_788);
or U1698 (N_1698,In_484,In_1628);
xnor U1699 (N_1699,In_297,In_152);
nor U1700 (N_1700,In_701,In_1296);
xnor U1701 (N_1701,In_927,In_336);
nor U1702 (N_1702,In_340,In_2374);
xor U1703 (N_1703,In_452,In_1080);
or U1704 (N_1704,In_2168,In_2012);
xor U1705 (N_1705,In_1375,In_1310);
and U1706 (N_1706,In_2336,In_1589);
xor U1707 (N_1707,In_1309,In_279);
nor U1708 (N_1708,In_1138,In_1347);
xnor U1709 (N_1709,In_1846,In_2302);
or U1710 (N_1710,In_2673,In_680);
or U1711 (N_1711,In_2723,In_1480);
nand U1712 (N_1712,In_1018,In_633);
nand U1713 (N_1713,In_2162,In_1089);
xor U1714 (N_1714,In_2317,In_1681);
xor U1715 (N_1715,In_13,In_2436);
nor U1716 (N_1716,In_2240,In_934);
nand U1717 (N_1717,In_976,In_1945);
xnor U1718 (N_1718,In_690,In_33);
xor U1719 (N_1719,In_414,In_2068);
or U1720 (N_1720,In_347,In_1678);
xor U1721 (N_1721,In_2913,In_1038);
or U1722 (N_1722,In_2372,In_1550);
nor U1723 (N_1723,In_1749,In_2700);
or U1724 (N_1724,In_248,In_2890);
nor U1725 (N_1725,In_1094,In_585);
nor U1726 (N_1726,In_2202,In_2814);
and U1727 (N_1727,In_2950,In_2123);
and U1728 (N_1728,In_44,In_2899);
nand U1729 (N_1729,In_2959,In_1669);
nand U1730 (N_1730,In_1747,In_2360);
or U1731 (N_1731,In_1893,In_2340);
nand U1732 (N_1732,In_304,In_849);
and U1733 (N_1733,In_2021,In_1117);
xnor U1734 (N_1734,In_490,In_1421);
and U1735 (N_1735,In_2569,In_950);
nor U1736 (N_1736,In_1992,In_1047);
and U1737 (N_1737,In_2224,In_454);
or U1738 (N_1738,In_2804,In_613);
nand U1739 (N_1739,In_304,In_883);
and U1740 (N_1740,In_575,In_2311);
or U1741 (N_1741,In_1313,In_1094);
xor U1742 (N_1742,In_309,In_1331);
nand U1743 (N_1743,In_1690,In_1110);
and U1744 (N_1744,In_509,In_1233);
or U1745 (N_1745,In_2501,In_1006);
nor U1746 (N_1746,In_2385,In_933);
nand U1747 (N_1747,In_284,In_215);
and U1748 (N_1748,In_700,In_138);
nand U1749 (N_1749,In_187,In_1940);
and U1750 (N_1750,In_2695,In_838);
nor U1751 (N_1751,In_819,In_2168);
xor U1752 (N_1752,In_1582,In_1535);
or U1753 (N_1753,In_2059,In_728);
or U1754 (N_1754,In_666,In_2179);
nand U1755 (N_1755,In_1581,In_1084);
xor U1756 (N_1756,In_2844,In_2466);
nor U1757 (N_1757,In_2396,In_1930);
or U1758 (N_1758,In_1502,In_2946);
or U1759 (N_1759,In_1689,In_1077);
nor U1760 (N_1760,In_781,In_933);
and U1761 (N_1761,In_2114,In_371);
or U1762 (N_1762,In_456,In_2981);
nor U1763 (N_1763,In_1425,In_2527);
and U1764 (N_1764,In_655,In_1929);
nor U1765 (N_1765,In_2073,In_1089);
nand U1766 (N_1766,In_1143,In_2625);
or U1767 (N_1767,In_1532,In_1768);
nor U1768 (N_1768,In_2599,In_13);
nand U1769 (N_1769,In_2535,In_2969);
nand U1770 (N_1770,In_1134,In_2721);
and U1771 (N_1771,In_1094,In_2461);
nor U1772 (N_1772,In_879,In_562);
xnor U1773 (N_1773,In_402,In_2188);
and U1774 (N_1774,In_2976,In_1506);
or U1775 (N_1775,In_1728,In_911);
or U1776 (N_1776,In_2662,In_1724);
nand U1777 (N_1777,In_2892,In_1586);
nand U1778 (N_1778,In_1475,In_1743);
nor U1779 (N_1779,In_2588,In_1915);
xor U1780 (N_1780,In_2691,In_658);
and U1781 (N_1781,In_2242,In_2198);
and U1782 (N_1782,In_199,In_757);
nor U1783 (N_1783,In_1009,In_2046);
xnor U1784 (N_1784,In_2351,In_1417);
or U1785 (N_1785,In_2165,In_1146);
xnor U1786 (N_1786,In_2278,In_1829);
nor U1787 (N_1787,In_2989,In_937);
nor U1788 (N_1788,In_606,In_406);
or U1789 (N_1789,In_1175,In_225);
nand U1790 (N_1790,In_2833,In_1150);
or U1791 (N_1791,In_287,In_892);
nand U1792 (N_1792,In_1746,In_1891);
xnor U1793 (N_1793,In_2871,In_2783);
xor U1794 (N_1794,In_1018,In_1112);
and U1795 (N_1795,In_816,In_50);
and U1796 (N_1796,In_1303,In_1343);
and U1797 (N_1797,In_2091,In_481);
or U1798 (N_1798,In_460,In_2843);
and U1799 (N_1799,In_1642,In_283);
or U1800 (N_1800,In_389,In_2576);
or U1801 (N_1801,In_276,In_620);
nor U1802 (N_1802,In_2121,In_897);
and U1803 (N_1803,In_1495,In_2070);
nand U1804 (N_1804,In_2373,In_1208);
or U1805 (N_1805,In_1402,In_2466);
and U1806 (N_1806,In_234,In_856);
xnor U1807 (N_1807,In_658,In_749);
nand U1808 (N_1808,In_2114,In_275);
nand U1809 (N_1809,In_1419,In_2526);
xnor U1810 (N_1810,In_996,In_843);
or U1811 (N_1811,In_2083,In_598);
and U1812 (N_1812,In_2170,In_2267);
nand U1813 (N_1813,In_830,In_1311);
nor U1814 (N_1814,In_1380,In_425);
xnor U1815 (N_1815,In_2233,In_1253);
xor U1816 (N_1816,In_538,In_438);
nor U1817 (N_1817,In_2427,In_986);
nor U1818 (N_1818,In_966,In_2930);
and U1819 (N_1819,In_2232,In_2288);
or U1820 (N_1820,In_2032,In_1813);
nor U1821 (N_1821,In_1177,In_2304);
or U1822 (N_1822,In_2369,In_2532);
and U1823 (N_1823,In_815,In_28);
or U1824 (N_1824,In_198,In_498);
nand U1825 (N_1825,In_175,In_2560);
and U1826 (N_1826,In_1797,In_1407);
or U1827 (N_1827,In_2755,In_249);
and U1828 (N_1828,In_920,In_2422);
nor U1829 (N_1829,In_421,In_1380);
nor U1830 (N_1830,In_1833,In_823);
nor U1831 (N_1831,In_2081,In_2832);
xnor U1832 (N_1832,In_1679,In_2799);
and U1833 (N_1833,In_104,In_2685);
nand U1834 (N_1834,In_2639,In_2508);
and U1835 (N_1835,In_1163,In_829);
and U1836 (N_1836,In_1180,In_2740);
xnor U1837 (N_1837,In_2232,In_428);
nor U1838 (N_1838,In_1655,In_2101);
or U1839 (N_1839,In_223,In_1523);
xnor U1840 (N_1840,In_663,In_2394);
or U1841 (N_1841,In_1518,In_1933);
nand U1842 (N_1842,In_123,In_1605);
xnor U1843 (N_1843,In_870,In_695);
xor U1844 (N_1844,In_626,In_2283);
nor U1845 (N_1845,In_1623,In_2);
and U1846 (N_1846,In_1675,In_1415);
xnor U1847 (N_1847,In_422,In_1895);
nand U1848 (N_1848,In_2516,In_133);
xor U1849 (N_1849,In_82,In_1870);
nand U1850 (N_1850,In_1016,In_1740);
xor U1851 (N_1851,In_1871,In_1756);
nor U1852 (N_1852,In_1748,In_1115);
xor U1853 (N_1853,In_2990,In_1981);
or U1854 (N_1854,In_336,In_454);
nand U1855 (N_1855,In_2275,In_88);
nand U1856 (N_1856,In_276,In_1984);
xor U1857 (N_1857,In_675,In_114);
nor U1858 (N_1858,In_485,In_666);
or U1859 (N_1859,In_2347,In_735);
nor U1860 (N_1860,In_2589,In_2163);
and U1861 (N_1861,In_1412,In_2348);
or U1862 (N_1862,In_786,In_288);
nor U1863 (N_1863,In_1520,In_960);
and U1864 (N_1864,In_200,In_1763);
xor U1865 (N_1865,In_2035,In_2037);
nor U1866 (N_1866,In_1157,In_242);
nand U1867 (N_1867,In_325,In_522);
nor U1868 (N_1868,In_2419,In_1595);
or U1869 (N_1869,In_2523,In_2248);
and U1870 (N_1870,In_2304,In_539);
xnor U1871 (N_1871,In_1391,In_1028);
xnor U1872 (N_1872,In_2616,In_1060);
or U1873 (N_1873,In_2167,In_2514);
nand U1874 (N_1874,In_289,In_2423);
and U1875 (N_1875,In_1758,In_597);
xnor U1876 (N_1876,In_2497,In_2912);
or U1877 (N_1877,In_1397,In_82);
xnor U1878 (N_1878,In_801,In_2685);
and U1879 (N_1879,In_1185,In_1547);
and U1880 (N_1880,In_1241,In_2208);
nor U1881 (N_1881,In_33,In_1751);
nor U1882 (N_1882,In_717,In_1619);
or U1883 (N_1883,In_1944,In_2876);
nor U1884 (N_1884,In_1107,In_2147);
or U1885 (N_1885,In_2956,In_1334);
nor U1886 (N_1886,In_914,In_2980);
xnor U1887 (N_1887,In_1808,In_1606);
or U1888 (N_1888,In_307,In_2055);
and U1889 (N_1889,In_2081,In_1755);
nand U1890 (N_1890,In_1841,In_1972);
xnor U1891 (N_1891,In_1724,In_1802);
xor U1892 (N_1892,In_106,In_55);
xnor U1893 (N_1893,In_100,In_938);
xnor U1894 (N_1894,In_2156,In_2204);
nand U1895 (N_1895,In_830,In_2675);
xnor U1896 (N_1896,In_1759,In_2477);
xor U1897 (N_1897,In_2071,In_191);
nand U1898 (N_1898,In_2996,In_943);
or U1899 (N_1899,In_2116,In_1072);
and U1900 (N_1900,In_275,In_2400);
nor U1901 (N_1901,In_2704,In_389);
nor U1902 (N_1902,In_956,In_1087);
or U1903 (N_1903,In_2069,In_2826);
xor U1904 (N_1904,In_40,In_1434);
or U1905 (N_1905,In_698,In_1584);
nor U1906 (N_1906,In_2687,In_1600);
nand U1907 (N_1907,In_1937,In_2931);
xnor U1908 (N_1908,In_1043,In_353);
xnor U1909 (N_1909,In_1530,In_791);
nor U1910 (N_1910,In_1549,In_2612);
nand U1911 (N_1911,In_1145,In_262);
and U1912 (N_1912,In_202,In_2174);
nand U1913 (N_1913,In_90,In_2800);
and U1914 (N_1914,In_1348,In_943);
and U1915 (N_1915,In_787,In_1117);
nand U1916 (N_1916,In_2993,In_233);
or U1917 (N_1917,In_1485,In_1049);
nor U1918 (N_1918,In_2327,In_30);
nor U1919 (N_1919,In_1703,In_1463);
xor U1920 (N_1920,In_361,In_2081);
nor U1921 (N_1921,In_2092,In_2790);
or U1922 (N_1922,In_1400,In_683);
or U1923 (N_1923,In_2458,In_1611);
or U1924 (N_1924,In_53,In_1805);
xnor U1925 (N_1925,In_1925,In_392);
nor U1926 (N_1926,In_1518,In_2464);
nor U1927 (N_1927,In_2196,In_1601);
nor U1928 (N_1928,In_1294,In_1797);
nand U1929 (N_1929,In_1553,In_1258);
and U1930 (N_1930,In_2285,In_2700);
xnor U1931 (N_1931,In_1750,In_1873);
and U1932 (N_1932,In_2543,In_38);
and U1933 (N_1933,In_152,In_1835);
nand U1934 (N_1934,In_1781,In_60);
nand U1935 (N_1935,In_1680,In_331);
or U1936 (N_1936,In_2423,In_23);
nand U1937 (N_1937,In_1924,In_1368);
or U1938 (N_1938,In_2379,In_207);
nand U1939 (N_1939,In_868,In_1279);
nor U1940 (N_1940,In_1785,In_1560);
nor U1941 (N_1941,In_2892,In_26);
nand U1942 (N_1942,In_574,In_2539);
and U1943 (N_1943,In_2871,In_790);
and U1944 (N_1944,In_1996,In_2491);
and U1945 (N_1945,In_2956,In_2296);
nand U1946 (N_1946,In_788,In_777);
xor U1947 (N_1947,In_1872,In_860);
and U1948 (N_1948,In_1977,In_1105);
nand U1949 (N_1949,In_1907,In_854);
and U1950 (N_1950,In_2218,In_2584);
or U1951 (N_1951,In_846,In_1516);
and U1952 (N_1952,In_2099,In_2266);
or U1953 (N_1953,In_2804,In_2758);
xor U1954 (N_1954,In_2694,In_1035);
nor U1955 (N_1955,In_2659,In_182);
nand U1956 (N_1956,In_229,In_2208);
nand U1957 (N_1957,In_732,In_1691);
nand U1958 (N_1958,In_1162,In_584);
and U1959 (N_1959,In_1710,In_2608);
or U1960 (N_1960,In_684,In_698);
nor U1961 (N_1961,In_1471,In_219);
or U1962 (N_1962,In_1147,In_2454);
xnor U1963 (N_1963,In_930,In_2981);
nand U1964 (N_1964,In_345,In_1324);
or U1965 (N_1965,In_2324,In_1837);
xnor U1966 (N_1966,In_796,In_1407);
nor U1967 (N_1967,In_2873,In_2759);
or U1968 (N_1968,In_719,In_685);
and U1969 (N_1969,In_1530,In_311);
xnor U1970 (N_1970,In_128,In_1884);
and U1971 (N_1971,In_1048,In_1981);
and U1972 (N_1972,In_1666,In_2171);
and U1973 (N_1973,In_1913,In_2057);
or U1974 (N_1974,In_2215,In_1252);
and U1975 (N_1975,In_1091,In_2168);
and U1976 (N_1976,In_1521,In_1201);
nand U1977 (N_1977,In_480,In_1675);
nor U1978 (N_1978,In_1907,In_1817);
and U1979 (N_1979,In_2226,In_86);
and U1980 (N_1980,In_2156,In_2891);
xor U1981 (N_1981,In_2090,In_1650);
xor U1982 (N_1982,In_993,In_410);
nor U1983 (N_1983,In_2733,In_700);
nor U1984 (N_1984,In_2793,In_1576);
nand U1985 (N_1985,In_1063,In_1053);
and U1986 (N_1986,In_1498,In_1228);
or U1987 (N_1987,In_2415,In_1585);
xnor U1988 (N_1988,In_69,In_1061);
nand U1989 (N_1989,In_526,In_1459);
and U1990 (N_1990,In_718,In_974);
nor U1991 (N_1991,In_2767,In_566);
nor U1992 (N_1992,In_1157,In_1298);
and U1993 (N_1993,In_726,In_1051);
nand U1994 (N_1994,In_1285,In_1759);
and U1995 (N_1995,In_2078,In_535);
xnor U1996 (N_1996,In_1388,In_1630);
or U1997 (N_1997,In_872,In_1465);
and U1998 (N_1998,In_1372,In_1071);
xor U1999 (N_1999,In_1139,In_2065);
xnor U2000 (N_2000,In_1917,In_2464);
nor U2001 (N_2001,In_1211,In_312);
and U2002 (N_2002,In_2688,In_2613);
xor U2003 (N_2003,In_202,In_2038);
xor U2004 (N_2004,In_2325,In_19);
and U2005 (N_2005,In_391,In_2937);
and U2006 (N_2006,In_2667,In_2119);
and U2007 (N_2007,In_1381,In_1623);
and U2008 (N_2008,In_1242,In_2981);
nand U2009 (N_2009,In_2651,In_2232);
xnor U2010 (N_2010,In_2954,In_254);
xor U2011 (N_2011,In_2225,In_2586);
nor U2012 (N_2012,In_836,In_1616);
nand U2013 (N_2013,In_76,In_2090);
xnor U2014 (N_2014,In_2024,In_1822);
or U2015 (N_2015,In_1488,In_2109);
or U2016 (N_2016,In_370,In_283);
or U2017 (N_2017,In_2588,In_1572);
and U2018 (N_2018,In_2676,In_2629);
or U2019 (N_2019,In_2039,In_2559);
and U2020 (N_2020,In_2877,In_1030);
or U2021 (N_2021,In_2574,In_1994);
and U2022 (N_2022,In_1031,In_1997);
nor U2023 (N_2023,In_2850,In_1733);
nand U2024 (N_2024,In_503,In_2442);
or U2025 (N_2025,In_221,In_320);
or U2026 (N_2026,In_1520,In_1130);
or U2027 (N_2027,In_1,In_440);
xnor U2028 (N_2028,In_1302,In_2571);
nand U2029 (N_2029,In_1947,In_1743);
xor U2030 (N_2030,In_2220,In_2523);
or U2031 (N_2031,In_1737,In_529);
nand U2032 (N_2032,In_1558,In_2783);
and U2033 (N_2033,In_1190,In_190);
and U2034 (N_2034,In_2241,In_2878);
xor U2035 (N_2035,In_436,In_2329);
xnor U2036 (N_2036,In_2903,In_277);
nor U2037 (N_2037,In_1470,In_1990);
or U2038 (N_2038,In_1809,In_888);
xor U2039 (N_2039,In_1809,In_1316);
xnor U2040 (N_2040,In_2664,In_2420);
nand U2041 (N_2041,In_2810,In_2790);
nor U2042 (N_2042,In_608,In_1460);
or U2043 (N_2043,In_2017,In_1825);
xor U2044 (N_2044,In_1875,In_2142);
nand U2045 (N_2045,In_2482,In_403);
and U2046 (N_2046,In_823,In_861);
and U2047 (N_2047,In_431,In_1956);
or U2048 (N_2048,In_1635,In_2130);
or U2049 (N_2049,In_1589,In_214);
xnor U2050 (N_2050,In_914,In_1147);
nand U2051 (N_2051,In_481,In_527);
nor U2052 (N_2052,In_1847,In_1762);
and U2053 (N_2053,In_1289,In_2306);
nor U2054 (N_2054,In_611,In_2344);
or U2055 (N_2055,In_2494,In_534);
xor U2056 (N_2056,In_836,In_1716);
or U2057 (N_2057,In_782,In_413);
nand U2058 (N_2058,In_2985,In_371);
xor U2059 (N_2059,In_1207,In_2623);
or U2060 (N_2060,In_1074,In_2324);
xor U2061 (N_2061,In_579,In_930);
and U2062 (N_2062,In_2914,In_2499);
or U2063 (N_2063,In_1432,In_1597);
nor U2064 (N_2064,In_2721,In_1748);
nor U2065 (N_2065,In_1104,In_1269);
or U2066 (N_2066,In_513,In_778);
xnor U2067 (N_2067,In_1396,In_2292);
nor U2068 (N_2068,In_2105,In_2947);
nor U2069 (N_2069,In_132,In_142);
nand U2070 (N_2070,In_181,In_395);
or U2071 (N_2071,In_662,In_855);
nand U2072 (N_2072,In_2851,In_2157);
and U2073 (N_2073,In_423,In_2005);
and U2074 (N_2074,In_1645,In_2386);
nand U2075 (N_2075,In_510,In_1206);
xnor U2076 (N_2076,In_48,In_2636);
nor U2077 (N_2077,In_1009,In_1528);
nor U2078 (N_2078,In_2096,In_1208);
xor U2079 (N_2079,In_383,In_6);
or U2080 (N_2080,In_1136,In_577);
nand U2081 (N_2081,In_269,In_1619);
or U2082 (N_2082,In_342,In_2385);
and U2083 (N_2083,In_606,In_578);
nand U2084 (N_2084,In_1971,In_2006);
xnor U2085 (N_2085,In_1530,In_535);
and U2086 (N_2086,In_285,In_1143);
nand U2087 (N_2087,In_1182,In_789);
and U2088 (N_2088,In_356,In_2083);
or U2089 (N_2089,In_808,In_1336);
or U2090 (N_2090,In_1806,In_2397);
or U2091 (N_2091,In_660,In_1898);
xnor U2092 (N_2092,In_2921,In_315);
nand U2093 (N_2093,In_2622,In_2739);
nand U2094 (N_2094,In_677,In_2208);
xnor U2095 (N_2095,In_287,In_1811);
and U2096 (N_2096,In_881,In_71);
or U2097 (N_2097,In_2077,In_1157);
nor U2098 (N_2098,In_736,In_2838);
xnor U2099 (N_2099,In_2294,In_1116);
or U2100 (N_2100,In_421,In_2962);
or U2101 (N_2101,In_678,In_2910);
nand U2102 (N_2102,In_71,In_310);
nor U2103 (N_2103,In_168,In_2197);
nor U2104 (N_2104,In_1944,In_2613);
or U2105 (N_2105,In_1996,In_1055);
or U2106 (N_2106,In_2415,In_362);
and U2107 (N_2107,In_1996,In_167);
xnor U2108 (N_2108,In_1328,In_162);
or U2109 (N_2109,In_627,In_2025);
nand U2110 (N_2110,In_2176,In_834);
or U2111 (N_2111,In_1512,In_2243);
nor U2112 (N_2112,In_2035,In_2104);
and U2113 (N_2113,In_2078,In_871);
nand U2114 (N_2114,In_856,In_223);
nand U2115 (N_2115,In_325,In_311);
nor U2116 (N_2116,In_2842,In_610);
and U2117 (N_2117,In_1108,In_468);
and U2118 (N_2118,In_1578,In_1453);
nand U2119 (N_2119,In_511,In_99);
or U2120 (N_2120,In_269,In_2177);
nor U2121 (N_2121,In_2715,In_71);
nor U2122 (N_2122,In_2761,In_110);
xnor U2123 (N_2123,In_2497,In_1879);
nor U2124 (N_2124,In_2852,In_2631);
and U2125 (N_2125,In_2395,In_1165);
nand U2126 (N_2126,In_2115,In_2595);
nand U2127 (N_2127,In_2047,In_892);
and U2128 (N_2128,In_1421,In_1500);
or U2129 (N_2129,In_2104,In_158);
or U2130 (N_2130,In_197,In_1482);
nand U2131 (N_2131,In_1989,In_1771);
or U2132 (N_2132,In_1600,In_1141);
xor U2133 (N_2133,In_779,In_2424);
and U2134 (N_2134,In_696,In_933);
xnor U2135 (N_2135,In_2988,In_2921);
nand U2136 (N_2136,In_1341,In_437);
and U2137 (N_2137,In_533,In_1429);
xnor U2138 (N_2138,In_1731,In_813);
nor U2139 (N_2139,In_466,In_2952);
nor U2140 (N_2140,In_635,In_128);
and U2141 (N_2141,In_499,In_2804);
nand U2142 (N_2142,In_2638,In_2994);
nand U2143 (N_2143,In_2885,In_367);
nand U2144 (N_2144,In_233,In_1798);
nand U2145 (N_2145,In_2304,In_745);
nor U2146 (N_2146,In_2199,In_840);
xnor U2147 (N_2147,In_1344,In_1237);
nand U2148 (N_2148,In_715,In_2390);
nand U2149 (N_2149,In_1201,In_1818);
nor U2150 (N_2150,In_2290,In_870);
or U2151 (N_2151,In_2958,In_2851);
and U2152 (N_2152,In_1154,In_2398);
nand U2153 (N_2153,In_539,In_1713);
nor U2154 (N_2154,In_991,In_2170);
xnor U2155 (N_2155,In_1440,In_2371);
nor U2156 (N_2156,In_798,In_2637);
or U2157 (N_2157,In_1260,In_855);
and U2158 (N_2158,In_2817,In_2908);
nand U2159 (N_2159,In_400,In_2044);
or U2160 (N_2160,In_973,In_1591);
xor U2161 (N_2161,In_1868,In_2147);
or U2162 (N_2162,In_1717,In_1163);
xor U2163 (N_2163,In_1937,In_12);
and U2164 (N_2164,In_2023,In_73);
and U2165 (N_2165,In_666,In_2008);
nor U2166 (N_2166,In_2920,In_1213);
and U2167 (N_2167,In_1026,In_2148);
or U2168 (N_2168,In_2122,In_263);
or U2169 (N_2169,In_1085,In_223);
nand U2170 (N_2170,In_2271,In_584);
or U2171 (N_2171,In_2840,In_2746);
xor U2172 (N_2172,In_565,In_702);
and U2173 (N_2173,In_136,In_1884);
nand U2174 (N_2174,In_2765,In_956);
xor U2175 (N_2175,In_268,In_2824);
or U2176 (N_2176,In_2586,In_149);
or U2177 (N_2177,In_2391,In_832);
xnor U2178 (N_2178,In_2432,In_2378);
or U2179 (N_2179,In_1464,In_2270);
xnor U2180 (N_2180,In_2476,In_1232);
nand U2181 (N_2181,In_2082,In_1296);
and U2182 (N_2182,In_681,In_1689);
or U2183 (N_2183,In_2636,In_2029);
and U2184 (N_2184,In_1807,In_2116);
nor U2185 (N_2185,In_2456,In_1244);
and U2186 (N_2186,In_1676,In_1549);
nor U2187 (N_2187,In_2017,In_441);
nor U2188 (N_2188,In_924,In_418);
nor U2189 (N_2189,In_1159,In_1372);
nor U2190 (N_2190,In_2426,In_111);
nor U2191 (N_2191,In_1483,In_274);
or U2192 (N_2192,In_1422,In_2400);
nor U2193 (N_2193,In_2834,In_2102);
nor U2194 (N_2194,In_454,In_739);
or U2195 (N_2195,In_559,In_2767);
nand U2196 (N_2196,In_366,In_12);
xnor U2197 (N_2197,In_361,In_1803);
or U2198 (N_2198,In_823,In_1774);
nor U2199 (N_2199,In_1894,In_2219);
nand U2200 (N_2200,In_811,In_2716);
and U2201 (N_2201,In_767,In_1043);
xnor U2202 (N_2202,In_947,In_2);
nor U2203 (N_2203,In_950,In_888);
and U2204 (N_2204,In_2440,In_2834);
nor U2205 (N_2205,In_1157,In_706);
or U2206 (N_2206,In_1912,In_1936);
nand U2207 (N_2207,In_726,In_2847);
nor U2208 (N_2208,In_2102,In_949);
and U2209 (N_2209,In_754,In_1199);
nor U2210 (N_2210,In_1422,In_635);
nor U2211 (N_2211,In_1654,In_128);
nor U2212 (N_2212,In_2812,In_934);
xor U2213 (N_2213,In_1817,In_332);
or U2214 (N_2214,In_2436,In_1297);
nand U2215 (N_2215,In_1930,In_1977);
and U2216 (N_2216,In_2197,In_1270);
and U2217 (N_2217,In_143,In_2951);
and U2218 (N_2218,In_2210,In_2808);
or U2219 (N_2219,In_2221,In_481);
xnor U2220 (N_2220,In_1435,In_2301);
nand U2221 (N_2221,In_2033,In_1429);
and U2222 (N_2222,In_2065,In_2490);
nand U2223 (N_2223,In_1054,In_1131);
nor U2224 (N_2224,In_437,In_1965);
nor U2225 (N_2225,In_2862,In_1424);
xnor U2226 (N_2226,In_760,In_714);
nor U2227 (N_2227,In_2641,In_1396);
nor U2228 (N_2228,In_2076,In_2610);
and U2229 (N_2229,In_819,In_1425);
xnor U2230 (N_2230,In_675,In_189);
and U2231 (N_2231,In_1852,In_1742);
and U2232 (N_2232,In_1731,In_1600);
nor U2233 (N_2233,In_473,In_2201);
and U2234 (N_2234,In_1515,In_2448);
or U2235 (N_2235,In_576,In_2177);
or U2236 (N_2236,In_195,In_1738);
or U2237 (N_2237,In_1847,In_16);
and U2238 (N_2238,In_2818,In_1822);
nand U2239 (N_2239,In_2610,In_2333);
and U2240 (N_2240,In_2218,In_2159);
and U2241 (N_2241,In_638,In_2910);
and U2242 (N_2242,In_0,In_1534);
xor U2243 (N_2243,In_340,In_168);
nand U2244 (N_2244,In_2237,In_487);
or U2245 (N_2245,In_654,In_1279);
xor U2246 (N_2246,In_2462,In_1485);
xor U2247 (N_2247,In_2806,In_1586);
nor U2248 (N_2248,In_1961,In_2941);
nand U2249 (N_2249,In_558,In_1430);
nor U2250 (N_2250,In_992,In_1535);
and U2251 (N_2251,In_2604,In_2731);
xnor U2252 (N_2252,In_919,In_67);
nand U2253 (N_2253,In_1007,In_378);
nor U2254 (N_2254,In_2880,In_1429);
nand U2255 (N_2255,In_1659,In_2924);
xor U2256 (N_2256,In_2646,In_1973);
or U2257 (N_2257,In_2106,In_596);
or U2258 (N_2258,In_1201,In_1949);
and U2259 (N_2259,In_2316,In_2671);
nand U2260 (N_2260,In_2738,In_2217);
nor U2261 (N_2261,In_2277,In_1631);
xor U2262 (N_2262,In_2110,In_722);
and U2263 (N_2263,In_1432,In_864);
nor U2264 (N_2264,In_2469,In_1817);
nor U2265 (N_2265,In_2730,In_2603);
xnor U2266 (N_2266,In_527,In_2502);
nand U2267 (N_2267,In_1538,In_2123);
nor U2268 (N_2268,In_611,In_2604);
nor U2269 (N_2269,In_484,In_657);
or U2270 (N_2270,In_401,In_2839);
and U2271 (N_2271,In_2231,In_1222);
xnor U2272 (N_2272,In_1457,In_2650);
xor U2273 (N_2273,In_2298,In_2231);
xor U2274 (N_2274,In_2615,In_1585);
nor U2275 (N_2275,In_2275,In_199);
or U2276 (N_2276,In_601,In_184);
and U2277 (N_2277,In_225,In_1645);
and U2278 (N_2278,In_2867,In_2816);
and U2279 (N_2279,In_1761,In_2426);
or U2280 (N_2280,In_2953,In_1677);
nor U2281 (N_2281,In_2355,In_2119);
nor U2282 (N_2282,In_857,In_2834);
nand U2283 (N_2283,In_1167,In_1517);
xor U2284 (N_2284,In_1950,In_2355);
or U2285 (N_2285,In_820,In_2566);
nand U2286 (N_2286,In_163,In_1037);
nor U2287 (N_2287,In_223,In_2214);
xor U2288 (N_2288,In_773,In_2733);
nor U2289 (N_2289,In_314,In_2601);
and U2290 (N_2290,In_2372,In_1822);
nor U2291 (N_2291,In_2205,In_2174);
nor U2292 (N_2292,In_1489,In_1895);
and U2293 (N_2293,In_759,In_1330);
nor U2294 (N_2294,In_1887,In_1842);
nor U2295 (N_2295,In_2808,In_1289);
or U2296 (N_2296,In_1528,In_2402);
nand U2297 (N_2297,In_1039,In_1394);
nand U2298 (N_2298,In_2838,In_2995);
or U2299 (N_2299,In_768,In_1793);
and U2300 (N_2300,In_2258,In_1483);
or U2301 (N_2301,In_2758,In_688);
nor U2302 (N_2302,In_2884,In_1622);
and U2303 (N_2303,In_809,In_2123);
and U2304 (N_2304,In_1440,In_909);
nand U2305 (N_2305,In_2978,In_462);
xor U2306 (N_2306,In_334,In_2980);
and U2307 (N_2307,In_147,In_2632);
and U2308 (N_2308,In_699,In_1517);
or U2309 (N_2309,In_1065,In_2989);
xnor U2310 (N_2310,In_2014,In_401);
or U2311 (N_2311,In_478,In_305);
nor U2312 (N_2312,In_1825,In_816);
xnor U2313 (N_2313,In_501,In_2777);
nand U2314 (N_2314,In_2942,In_2668);
or U2315 (N_2315,In_1246,In_2761);
or U2316 (N_2316,In_437,In_2586);
xnor U2317 (N_2317,In_818,In_1002);
nand U2318 (N_2318,In_1291,In_2989);
or U2319 (N_2319,In_2218,In_2713);
nor U2320 (N_2320,In_2746,In_2139);
and U2321 (N_2321,In_2669,In_2338);
nor U2322 (N_2322,In_2144,In_2062);
or U2323 (N_2323,In_2916,In_680);
or U2324 (N_2324,In_1826,In_987);
xnor U2325 (N_2325,In_367,In_831);
nor U2326 (N_2326,In_1983,In_590);
nand U2327 (N_2327,In_1352,In_2016);
nand U2328 (N_2328,In_1782,In_533);
nand U2329 (N_2329,In_20,In_444);
and U2330 (N_2330,In_85,In_539);
and U2331 (N_2331,In_1158,In_122);
nand U2332 (N_2332,In_1717,In_2556);
xnor U2333 (N_2333,In_1109,In_2204);
or U2334 (N_2334,In_2394,In_1822);
and U2335 (N_2335,In_1728,In_223);
nor U2336 (N_2336,In_218,In_1737);
nor U2337 (N_2337,In_1592,In_201);
nor U2338 (N_2338,In_518,In_1003);
xnor U2339 (N_2339,In_2804,In_1913);
and U2340 (N_2340,In_2480,In_540);
and U2341 (N_2341,In_820,In_122);
nand U2342 (N_2342,In_778,In_2189);
nand U2343 (N_2343,In_1469,In_2641);
nand U2344 (N_2344,In_1799,In_2776);
nor U2345 (N_2345,In_2052,In_640);
xor U2346 (N_2346,In_723,In_2806);
xor U2347 (N_2347,In_987,In_2463);
xnor U2348 (N_2348,In_950,In_2552);
xnor U2349 (N_2349,In_296,In_2956);
or U2350 (N_2350,In_1733,In_661);
nor U2351 (N_2351,In_400,In_2194);
xnor U2352 (N_2352,In_102,In_1728);
nor U2353 (N_2353,In_2434,In_892);
xor U2354 (N_2354,In_801,In_391);
nor U2355 (N_2355,In_2701,In_520);
nand U2356 (N_2356,In_307,In_1764);
nor U2357 (N_2357,In_2445,In_1153);
nor U2358 (N_2358,In_2140,In_2060);
nand U2359 (N_2359,In_344,In_883);
xor U2360 (N_2360,In_1039,In_2943);
nand U2361 (N_2361,In_2158,In_429);
nand U2362 (N_2362,In_1725,In_550);
nand U2363 (N_2363,In_1128,In_962);
xor U2364 (N_2364,In_734,In_2339);
xor U2365 (N_2365,In_2068,In_4);
xor U2366 (N_2366,In_1553,In_790);
nor U2367 (N_2367,In_1760,In_494);
and U2368 (N_2368,In_1635,In_2896);
xor U2369 (N_2369,In_2125,In_338);
and U2370 (N_2370,In_1243,In_1540);
xor U2371 (N_2371,In_1266,In_829);
nand U2372 (N_2372,In_2276,In_2516);
nor U2373 (N_2373,In_1588,In_2162);
nor U2374 (N_2374,In_1357,In_2993);
nor U2375 (N_2375,In_1669,In_188);
and U2376 (N_2376,In_2491,In_1475);
or U2377 (N_2377,In_1180,In_387);
nor U2378 (N_2378,In_931,In_2135);
and U2379 (N_2379,In_2850,In_661);
and U2380 (N_2380,In_2370,In_1173);
and U2381 (N_2381,In_2677,In_1331);
nand U2382 (N_2382,In_2425,In_1540);
nand U2383 (N_2383,In_556,In_925);
nand U2384 (N_2384,In_1101,In_2934);
xor U2385 (N_2385,In_1920,In_994);
and U2386 (N_2386,In_91,In_2314);
or U2387 (N_2387,In_1400,In_1178);
and U2388 (N_2388,In_305,In_1077);
nor U2389 (N_2389,In_2503,In_798);
and U2390 (N_2390,In_1832,In_2182);
nand U2391 (N_2391,In_658,In_962);
nor U2392 (N_2392,In_1432,In_1476);
nor U2393 (N_2393,In_2914,In_2447);
nor U2394 (N_2394,In_2028,In_502);
nor U2395 (N_2395,In_81,In_1729);
xor U2396 (N_2396,In_175,In_954);
and U2397 (N_2397,In_1664,In_633);
and U2398 (N_2398,In_2750,In_1875);
nand U2399 (N_2399,In_1360,In_388);
nor U2400 (N_2400,In_792,In_2781);
xor U2401 (N_2401,In_1063,In_2147);
or U2402 (N_2402,In_130,In_933);
nor U2403 (N_2403,In_283,In_679);
nand U2404 (N_2404,In_756,In_228);
xnor U2405 (N_2405,In_2441,In_2279);
or U2406 (N_2406,In_2220,In_929);
or U2407 (N_2407,In_2063,In_434);
and U2408 (N_2408,In_1145,In_427);
and U2409 (N_2409,In_2291,In_169);
nor U2410 (N_2410,In_1018,In_1919);
xor U2411 (N_2411,In_1302,In_166);
xnor U2412 (N_2412,In_1826,In_41);
or U2413 (N_2413,In_437,In_748);
nor U2414 (N_2414,In_894,In_1346);
nand U2415 (N_2415,In_2183,In_1795);
and U2416 (N_2416,In_685,In_607);
or U2417 (N_2417,In_1908,In_704);
nor U2418 (N_2418,In_2289,In_705);
or U2419 (N_2419,In_1987,In_1957);
or U2420 (N_2420,In_1798,In_797);
nor U2421 (N_2421,In_1343,In_2938);
xor U2422 (N_2422,In_1559,In_173);
xor U2423 (N_2423,In_1596,In_1999);
xor U2424 (N_2424,In_2986,In_2336);
or U2425 (N_2425,In_880,In_2027);
nor U2426 (N_2426,In_2211,In_2197);
and U2427 (N_2427,In_904,In_2040);
nor U2428 (N_2428,In_1778,In_2018);
and U2429 (N_2429,In_2440,In_529);
nand U2430 (N_2430,In_108,In_2600);
or U2431 (N_2431,In_800,In_2234);
and U2432 (N_2432,In_1292,In_1507);
nor U2433 (N_2433,In_2708,In_471);
and U2434 (N_2434,In_2859,In_639);
nor U2435 (N_2435,In_161,In_1658);
nor U2436 (N_2436,In_239,In_2100);
or U2437 (N_2437,In_1855,In_123);
xnor U2438 (N_2438,In_2056,In_175);
and U2439 (N_2439,In_2123,In_1062);
xor U2440 (N_2440,In_2355,In_1034);
nand U2441 (N_2441,In_1083,In_1851);
and U2442 (N_2442,In_772,In_1205);
nor U2443 (N_2443,In_2487,In_211);
xor U2444 (N_2444,In_2485,In_283);
or U2445 (N_2445,In_1662,In_991);
xor U2446 (N_2446,In_734,In_204);
or U2447 (N_2447,In_585,In_1878);
nor U2448 (N_2448,In_1777,In_1732);
nand U2449 (N_2449,In_2749,In_2545);
nand U2450 (N_2450,In_2452,In_949);
and U2451 (N_2451,In_828,In_1782);
nor U2452 (N_2452,In_1760,In_2944);
or U2453 (N_2453,In_2510,In_1639);
nand U2454 (N_2454,In_1288,In_1449);
nor U2455 (N_2455,In_2871,In_1950);
or U2456 (N_2456,In_2506,In_1326);
and U2457 (N_2457,In_1336,In_1590);
nor U2458 (N_2458,In_1596,In_1516);
and U2459 (N_2459,In_515,In_2290);
nand U2460 (N_2460,In_796,In_2470);
nor U2461 (N_2461,In_2141,In_1351);
or U2462 (N_2462,In_430,In_2633);
or U2463 (N_2463,In_686,In_1456);
and U2464 (N_2464,In_927,In_534);
xor U2465 (N_2465,In_826,In_205);
and U2466 (N_2466,In_1931,In_1732);
and U2467 (N_2467,In_2726,In_573);
or U2468 (N_2468,In_1698,In_831);
xor U2469 (N_2469,In_45,In_1543);
and U2470 (N_2470,In_746,In_1168);
nand U2471 (N_2471,In_1455,In_2437);
nand U2472 (N_2472,In_1585,In_201);
xor U2473 (N_2473,In_161,In_2534);
xor U2474 (N_2474,In_2397,In_1280);
and U2475 (N_2475,In_1326,In_1124);
nor U2476 (N_2476,In_1198,In_731);
nand U2477 (N_2477,In_2129,In_2890);
xor U2478 (N_2478,In_2662,In_1954);
nor U2479 (N_2479,In_913,In_551);
nand U2480 (N_2480,In_343,In_1531);
nor U2481 (N_2481,In_2716,In_517);
nand U2482 (N_2482,In_2157,In_1872);
or U2483 (N_2483,In_1562,In_957);
or U2484 (N_2484,In_2771,In_2897);
or U2485 (N_2485,In_2085,In_2296);
nor U2486 (N_2486,In_839,In_2137);
xor U2487 (N_2487,In_2488,In_2601);
nand U2488 (N_2488,In_1634,In_1246);
nor U2489 (N_2489,In_2869,In_595);
or U2490 (N_2490,In_2482,In_2992);
or U2491 (N_2491,In_1365,In_1351);
and U2492 (N_2492,In_2430,In_2995);
and U2493 (N_2493,In_1699,In_934);
nor U2494 (N_2494,In_39,In_2239);
nor U2495 (N_2495,In_2761,In_2544);
and U2496 (N_2496,In_900,In_1072);
nand U2497 (N_2497,In_1060,In_1160);
or U2498 (N_2498,In_949,In_494);
xnor U2499 (N_2499,In_967,In_2763);
nor U2500 (N_2500,In_2070,In_2455);
nand U2501 (N_2501,In_2527,In_2056);
and U2502 (N_2502,In_1125,In_682);
nor U2503 (N_2503,In_2421,In_778);
and U2504 (N_2504,In_482,In_2475);
nand U2505 (N_2505,In_988,In_2035);
nand U2506 (N_2506,In_1118,In_745);
xor U2507 (N_2507,In_2818,In_1459);
nor U2508 (N_2508,In_1390,In_897);
xor U2509 (N_2509,In_519,In_34);
and U2510 (N_2510,In_1821,In_1789);
nor U2511 (N_2511,In_902,In_1383);
and U2512 (N_2512,In_280,In_926);
and U2513 (N_2513,In_163,In_1451);
nor U2514 (N_2514,In_652,In_2830);
or U2515 (N_2515,In_2264,In_1217);
xnor U2516 (N_2516,In_1652,In_2136);
or U2517 (N_2517,In_1913,In_1437);
nor U2518 (N_2518,In_2085,In_873);
nand U2519 (N_2519,In_2151,In_860);
nand U2520 (N_2520,In_917,In_895);
or U2521 (N_2521,In_2011,In_2606);
nor U2522 (N_2522,In_2582,In_2319);
xnor U2523 (N_2523,In_114,In_1945);
nand U2524 (N_2524,In_144,In_236);
or U2525 (N_2525,In_2139,In_2797);
nor U2526 (N_2526,In_1758,In_2668);
nor U2527 (N_2527,In_820,In_744);
or U2528 (N_2528,In_774,In_1951);
xor U2529 (N_2529,In_1014,In_1809);
nand U2530 (N_2530,In_1350,In_1042);
or U2531 (N_2531,In_876,In_830);
nor U2532 (N_2532,In_1473,In_1827);
and U2533 (N_2533,In_2844,In_1575);
nor U2534 (N_2534,In_1597,In_1923);
and U2535 (N_2535,In_2747,In_718);
and U2536 (N_2536,In_1442,In_1138);
or U2537 (N_2537,In_926,In_1698);
or U2538 (N_2538,In_1687,In_2474);
xor U2539 (N_2539,In_2982,In_497);
or U2540 (N_2540,In_71,In_105);
xnor U2541 (N_2541,In_492,In_1370);
nand U2542 (N_2542,In_1815,In_903);
nand U2543 (N_2543,In_1783,In_688);
and U2544 (N_2544,In_2525,In_1379);
and U2545 (N_2545,In_366,In_152);
nor U2546 (N_2546,In_1572,In_2925);
xnor U2547 (N_2547,In_2361,In_2620);
xnor U2548 (N_2548,In_2306,In_2088);
and U2549 (N_2549,In_755,In_2400);
or U2550 (N_2550,In_712,In_327);
nand U2551 (N_2551,In_597,In_1808);
xor U2552 (N_2552,In_1577,In_344);
and U2553 (N_2553,In_1395,In_302);
nand U2554 (N_2554,In_1171,In_861);
nor U2555 (N_2555,In_776,In_889);
nand U2556 (N_2556,In_233,In_2693);
nand U2557 (N_2557,In_579,In_296);
nand U2558 (N_2558,In_2472,In_606);
and U2559 (N_2559,In_409,In_1592);
and U2560 (N_2560,In_244,In_1343);
nor U2561 (N_2561,In_2393,In_1930);
xnor U2562 (N_2562,In_9,In_2225);
or U2563 (N_2563,In_1453,In_494);
nand U2564 (N_2564,In_2577,In_2077);
and U2565 (N_2565,In_472,In_2517);
nand U2566 (N_2566,In_1246,In_2605);
and U2567 (N_2567,In_2194,In_2552);
nand U2568 (N_2568,In_119,In_1012);
nor U2569 (N_2569,In_1476,In_529);
nand U2570 (N_2570,In_2589,In_1893);
and U2571 (N_2571,In_1437,In_832);
or U2572 (N_2572,In_1007,In_2916);
nor U2573 (N_2573,In_771,In_1680);
nor U2574 (N_2574,In_1839,In_702);
xnor U2575 (N_2575,In_488,In_2966);
xnor U2576 (N_2576,In_1041,In_2798);
nand U2577 (N_2577,In_1541,In_1648);
nor U2578 (N_2578,In_2827,In_799);
and U2579 (N_2579,In_1449,In_2551);
nor U2580 (N_2580,In_2277,In_514);
nand U2581 (N_2581,In_2061,In_2512);
xor U2582 (N_2582,In_2170,In_1372);
nand U2583 (N_2583,In_758,In_1700);
nand U2584 (N_2584,In_2697,In_1030);
and U2585 (N_2585,In_619,In_1312);
nor U2586 (N_2586,In_600,In_557);
nand U2587 (N_2587,In_222,In_652);
or U2588 (N_2588,In_408,In_530);
and U2589 (N_2589,In_1132,In_668);
or U2590 (N_2590,In_2395,In_1321);
and U2591 (N_2591,In_2827,In_2384);
nor U2592 (N_2592,In_330,In_1339);
nand U2593 (N_2593,In_1899,In_1474);
nand U2594 (N_2594,In_768,In_1549);
nor U2595 (N_2595,In_1637,In_896);
or U2596 (N_2596,In_2132,In_263);
nor U2597 (N_2597,In_2735,In_2265);
xor U2598 (N_2598,In_1715,In_898);
nor U2599 (N_2599,In_159,In_743);
xor U2600 (N_2600,In_576,In_2828);
nand U2601 (N_2601,In_1219,In_716);
and U2602 (N_2602,In_2777,In_30);
nor U2603 (N_2603,In_1094,In_471);
or U2604 (N_2604,In_406,In_2589);
xor U2605 (N_2605,In_2461,In_2559);
xor U2606 (N_2606,In_2868,In_1837);
nand U2607 (N_2607,In_2921,In_2856);
nand U2608 (N_2608,In_2222,In_2182);
and U2609 (N_2609,In_851,In_446);
nor U2610 (N_2610,In_1568,In_255);
or U2611 (N_2611,In_2944,In_2683);
nor U2612 (N_2612,In_810,In_878);
or U2613 (N_2613,In_519,In_206);
or U2614 (N_2614,In_804,In_2897);
and U2615 (N_2615,In_918,In_1379);
or U2616 (N_2616,In_2104,In_93);
nor U2617 (N_2617,In_1014,In_715);
nor U2618 (N_2618,In_2867,In_786);
nor U2619 (N_2619,In_960,In_896);
and U2620 (N_2620,In_1930,In_156);
xor U2621 (N_2621,In_2432,In_404);
xnor U2622 (N_2622,In_249,In_2081);
nor U2623 (N_2623,In_707,In_421);
nor U2624 (N_2624,In_1705,In_31);
nand U2625 (N_2625,In_2748,In_2863);
nand U2626 (N_2626,In_635,In_1547);
or U2627 (N_2627,In_559,In_684);
or U2628 (N_2628,In_135,In_1963);
and U2629 (N_2629,In_2384,In_348);
or U2630 (N_2630,In_2664,In_1919);
nand U2631 (N_2631,In_180,In_602);
xor U2632 (N_2632,In_75,In_1432);
nand U2633 (N_2633,In_2595,In_1796);
and U2634 (N_2634,In_2065,In_2550);
and U2635 (N_2635,In_2879,In_495);
or U2636 (N_2636,In_1411,In_830);
nand U2637 (N_2637,In_570,In_2172);
nand U2638 (N_2638,In_2004,In_950);
nand U2639 (N_2639,In_2897,In_1796);
or U2640 (N_2640,In_1594,In_357);
or U2641 (N_2641,In_1408,In_1486);
and U2642 (N_2642,In_817,In_977);
nor U2643 (N_2643,In_2080,In_2273);
xnor U2644 (N_2644,In_1293,In_1317);
and U2645 (N_2645,In_1158,In_1321);
nor U2646 (N_2646,In_1098,In_1581);
or U2647 (N_2647,In_259,In_2086);
xor U2648 (N_2648,In_204,In_2926);
and U2649 (N_2649,In_718,In_62);
xor U2650 (N_2650,In_1681,In_1459);
nand U2651 (N_2651,In_2909,In_2187);
nand U2652 (N_2652,In_101,In_2544);
nand U2653 (N_2653,In_2907,In_1938);
nor U2654 (N_2654,In_2955,In_1150);
nor U2655 (N_2655,In_1838,In_37);
nor U2656 (N_2656,In_2427,In_1417);
xnor U2657 (N_2657,In_886,In_2499);
xnor U2658 (N_2658,In_2208,In_1918);
xor U2659 (N_2659,In_2470,In_2511);
or U2660 (N_2660,In_2364,In_1165);
and U2661 (N_2661,In_808,In_1663);
xor U2662 (N_2662,In_715,In_1388);
xnor U2663 (N_2663,In_1349,In_1267);
nand U2664 (N_2664,In_887,In_2340);
xor U2665 (N_2665,In_1075,In_511);
nand U2666 (N_2666,In_2749,In_1750);
xor U2667 (N_2667,In_2078,In_330);
nor U2668 (N_2668,In_1745,In_804);
nor U2669 (N_2669,In_940,In_952);
xnor U2670 (N_2670,In_1399,In_1232);
or U2671 (N_2671,In_2145,In_180);
or U2672 (N_2672,In_2155,In_800);
xor U2673 (N_2673,In_2975,In_1111);
nor U2674 (N_2674,In_1064,In_248);
nand U2675 (N_2675,In_688,In_2713);
nand U2676 (N_2676,In_2043,In_1584);
and U2677 (N_2677,In_2371,In_802);
or U2678 (N_2678,In_2544,In_312);
nand U2679 (N_2679,In_2492,In_2707);
and U2680 (N_2680,In_766,In_1911);
and U2681 (N_2681,In_1915,In_1159);
or U2682 (N_2682,In_653,In_561);
xnor U2683 (N_2683,In_2106,In_698);
nor U2684 (N_2684,In_1348,In_54);
or U2685 (N_2685,In_2666,In_1693);
nand U2686 (N_2686,In_2700,In_273);
nor U2687 (N_2687,In_2515,In_2867);
nor U2688 (N_2688,In_214,In_1895);
xor U2689 (N_2689,In_1240,In_2787);
xor U2690 (N_2690,In_2465,In_311);
or U2691 (N_2691,In_1390,In_1062);
xnor U2692 (N_2692,In_1547,In_661);
nand U2693 (N_2693,In_2882,In_2894);
nor U2694 (N_2694,In_398,In_1293);
or U2695 (N_2695,In_157,In_44);
or U2696 (N_2696,In_77,In_2656);
nand U2697 (N_2697,In_2984,In_752);
nand U2698 (N_2698,In_1404,In_78);
xor U2699 (N_2699,In_697,In_1953);
nor U2700 (N_2700,In_26,In_727);
nor U2701 (N_2701,In_2982,In_177);
xnor U2702 (N_2702,In_2628,In_806);
nor U2703 (N_2703,In_777,In_2659);
and U2704 (N_2704,In_1288,In_155);
nor U2705 (N_2705,In_1607,In_1831);
and U2706 (N_2706,In_1448,In_643);
xor U2707 (N_2707,In_2728,In_1415);
and U2708 (N_2708,In_2351,In_184);
xor U2709 (N_2709,In_1999,In_2568);
nor U2710 (N_2710,In_1198,In_1042);
nand U2711 (N_2711,In_926,In_956);
nor U2712 (N_2712,In_1361,In_638);
or U2713 (N_2713,In_2679,In_2247);
xor U2714 (N_2714,In_303,In_680);
xor U2715 (N_2715,In_2713,In_805);
or U2716 (N_2716,In_183,In_2964);
or U2717 (N_2717,In_2750,In_2973);
nand U2718 (N_2718,In_2307,In_516);
and U2719 (N_2719,In_1449,In_716);
or U2720 (N_2720,In_1973,In_2096);
xor U2721 (N_2721,In_955,In_1402);
nor U2722 (N_2722,In_2026,In_246);
xnor U2723 (N_2723,In_102,In_298);
or U2724 (N_2724,In_2870,In_1952);
nor U2725 (N_2725,In_1743,In_1244);
nor U2726 (N_2726,In_2477,In_860);
nor U2727 (N_2727,In_2343,In_1731);
nand U2728 (N_2728,In_1995,In_1545);
xnor U2729 (N_2729,In_660,In_203);
nor U2730 (N_2730,In_1505,In_788);
nand U2731 (N_2731,In_2971,In_2936);
nand U2732 (N_2732,In_264,In_90);
xor U2733 (N_2733,In_2938,In_2622);
nor U2734 (N_2734,In_2980,In_2462);
nand U2735 (N_2735,In_487,In_195);
xor U2736 (N_2736,In_1200,In_1193);
nor U2737 (N_2737,In_2941,In_2751);
and U2738 (N_2738,In_1579,In_2455);
or U2739 (N_2739,In_33,In_2270);
nand U2740 (N_2740,In_605,In_1013);
nor U2741 (N_2741,In_1845,In_985);
xor U2742 (N_2742,In_1318,In_768);
and U2743 (N_2743,In_1295,In_2773);
and U2744 (N_2744,In_1534,In_1954);
or U2745 (N_2745,In_363,In_2190);
nor U2746 (N_2746,In_2042,In_1103);
nand U2747 (N_2747,In_1719,In_2755);
nor U2748 (N_2748,In_2288,In_756);
xnor U2749 (N_2749,In_1055,In_1662);
xor U2750 (N_2750,In_42,In_1868);
nor U2751 (N_2751,In_843,In_252);
xnor U2752 (N_2752,In_2544,In_1501);
and U2753 (N_2753,In_1170,In_391);
nor U2754 (N_2754,In_2890,In_785);
nand U2755 (N_2755,In_2398,In_2970);
and U2756 (N_2756,In_1355,In_1119);
nor U2757 (N_2757,In_694,In_870);
nand U2758 (N_2758,In_2722,In_1166);
and U2759 (N_2759,In_2055,In_649);
and U2760 (N_2760,In_761,In_1890);
or U2761 (N_2761,In_230,In_2295);
nand U2762 (N_2762,In_1529,In_509);
nand U2763 (N_2763,In_683,In_2548);
xnor U2764 (N_2764,In_1727,In_994);
or U2765 (N_2765,In_496,In_119);
nor U2766 (N_2766,In_1673,In_380);
xor U2767 (N_2767,In_1684,In_760);
or U2768 (N_2768,In_959,In_1827);
nor U2769 (N_2769,In_1351,In_2844);
or U2770 (N_2770,In_2432,In_122);
xor U2771 (N_2771,In_1833,In_2474);
nand U2772 (N_2772,In_1550,In_813);
and U2773 (N_2773,In_393,In_288);
nand U2774 (N_2774,In_1305,In_215);
xnor U2775 (N_2775,In_2422,In_2661);
nand U2776 (N_2776,In_2550,In_2194);
or U2777 (N_2777,In_2747,In_2984);
nand U2778 (N_2778,In_828,In_2368);
xnor U2779 (N_2779,In_2525,In_372);
nand U2780 (N_2780,In_2377,In_2240);
xnor U2781 (N_2781,In_538,In_302);
nor U2782 (N_2782,In_654,In_409);
nand U2783 (N_2783,In_1483,In_562);
and U2784 (N_2784,In_2648,In_2262);
nand U2785 (N_2785,In_225,In_1041);
xnor U2786 (N_2786,In_1082,In_497);
nor U2787 (N_2787,In_225,In_2358);
xnor U2788 (N_2788,In_2100,In_1166);
and U2789 (N_2789,In_585,In_936);
xor U2790 (N_2790,In_2196,In_2013);
nand U2791 (N_2791,In_791,In_2340);
nand U2792 (N_2792,In_909,In_2418);
and U2793 (N_2793,In_1567,In_1071);
nand U2794 (N_2794,In_2618,In_1153);
or U2795 (N_2795,In_492,In_573);
xor U2796 (N_2796,In_1790,In_2109);
or U2797 (N_2797,In_2163,In_870);
nand U2798 (N_2798,In_2140,In_1757);
nand U2799 (N_2799,In_338,In_2748);
xor U2800 (N_2800,In_1315,In_1687);
nand U2801 (N_2801,In_461,In_1618);
xor U2802 (N_2802,In_2892,In_1547);
or U2803 (N_2803,In_116,In_1058);
nand U2804 (N_2804,In_2866,In_303);
nor U2805 (N_2805,In_1191,In_2349);
nor U2806 (N_2806,In_848,In_2940);
nor U2807 (N_2807,In_491,In_819);
nor U2808 (N_2808,In_2927,In_301);
nor U2809 (N_2809,In_1174,In_2452);
nor U2810 (N_2810,In_1839,In_511);
or U2811 (N_2811,In_465,In_1909);
xnor U2812 (N_2812,In_1121,In_2102);
nand U2813 (N_2813,In_1759,In_943);
nor U2814 (N_2814,In_132,In_1014);
xor U2815 (N_2815,In_2465,In_2137);
nor U2816 (N_2816,In_1508,In_2110);
and U2817 (N_2817,In_2977,In_2680);
or U2818 (N_2818,In_2889,In_2208);
and U2819 (N_2819,In_1684,In_2916);
nand U2820 (N_2820,In_1642,In_1254);
xnor U2821 (N_2821,In_2222,In_2091);
and U2822 (N_2822,In_44,In_1835);
nor U2823 (N_2823,In_1839,In_919);
and U2824 (N_2824,In_12,In_1393);
xor U2825 (N_2825,In_2138,In_2411);
and U2826 (N_2826,In_1833,In_2362);
xnor U2827 (N_2827,In_1297,In_1909);
or U2828 (N_2828,In_1322,In_126);
or U2829 (N_2829,In_2455,In_1415);
nor U2830 (N_2830,In_1997,In_1816);
nor U2831 (N_2831,In_722,In_512);
and U2832 (N_2832,In_2772,In_86);
nor U2833 (N_2833,In_2749,In_390);
and U2834 (N_2834,In_196,In_2217);
and U2835 (N_2835,In_2096,In_2919);
nand U2836 (N_2836,In_2289,In_466);
and U2837 (N_2837,In_830,In_2215);
xor U2838 (N_2838,In_1261,In_414);
nand U2839 (N_2839,In_2676,In_204);
nor U2840 (N_2840,In_1972,In_2575);
nor U2841 (N_2841,In_644,In_2638);
xor U2842 (N_2842,In_2553,In_2634);
nor U2843 (N_2843,In_2370,In_2032);
nand U2844 (N_2844,In_662,In_784);
nor U2845 (N_2845,In_1331,In_2414);
xor U2846 (N_2846,In_1407,In_2631);
nor U2847 (N_2847,In_1098,In_775);
and U2848 (N_2848,In_1216,In_1665);
nor U2849 (N_2849,In_1224,In_1821);
nor U2850 (N_2850,In_2945,In_1422);
nor U2851 (N_2851,In_1519,In_1928);
nor U2852 (N_2852,In_2651,In_2734);
nor U2853 (N_2853,In_1437,In_1303);
nor U2854 (N_2854,In_2159,In_1746);
or U2855 (N_2855,In_2522,In_469);
nor U2856 (N_2856,In_1866,In_1939);
xnor U2857 (N_2857,In_608,In_2667);
or U2858 (N_2858,In_2415,In_130);
nand U2859 (N_2859,In_466,In_420);
and U2860 (N_2860,In_1002,In_1581);
nand U2861 (N_2861,In_1849,In_1741);
xnor U2862 (N_2862,In_701,In_937);
xnor U2863 (N_2863,In_1192,In_2534);
and U2864 (N_2864,In_187,In_2238);
or U2865 (N_2865,In_1371,In_1155);
nand U2866 (N_2866,In_1758,In_418);
and U2867 (N_2867,In_1702,In_2407);
nand U2868 (N_2868,In_1863,In_2816);
nor U2869 (N_2869,In_964,In_2466);
or U2870 (N_2870,In_2040,In_2374);
nand U2871 (N_2871,In_553,In_1196);
xnor U2872 (N_2872,In_207,In_1667);
or U2873 (N_2873,In_2088,In_1952);
nand U2874 (N_2874,In_88,In_1255);
nand U2875 (N_2875,In_2819,In_2434);
nor U2876 (N_2876,In_2082,In_1563);
or U2877 (N_2877,In_1914,In_1731);
and U2878 (N_2878,In_1169,In_1080);
and U2879 (N_2879,In_947,In_2458);
or U2880 (N_2880,In_2966,In_1363);
or U2881 (N_2881,In_1601,In_2400);
or U2882 (N_2882,In_48,In_1720);
nor U2883 (N_2883,In_1219,In_2972);
and U2884 (N_2884,In_357,In_903);
nor U2885 (N_2885,In_1031,In_2388);
xnor U2886 (N_2886,In_1502,In_1814);
or U2887 (N_2887,In_370,In_1543);
and U2888 (N_2888,In_411,In_70);
or U2889 (N_2889,In_2094,In_551);
and U2890 (N_2890,In_1966,In_1025);
xor U2891 (N_2891,In_561,In_1387);
xnor U2892 (N_2892,In_171,In_780);
xor U2893 (N_2893,In_1011,In_725);
or U2894 (N_2894,In_2757,In_1007);
and U2895 (N_2895,In_1742,In_2815);
xor U2896 (N_2896,In_2808,In_17);
nor U2897 (N_2897,In_834,In_1940);
nor U2898 (N_2898,In_1479,In_26);
and U2899 (N_2899,In_1138,In_346);
xnor U2900 (N_2900,In_1810,In_2141);
and U2901 (N_2901,In_1,In_2967);
nor U2902 (N_2902,In_468,In_235);
nand U2903 (N_2903,In_2390,In_276);
nand U2904 (N_2904,In_2484,In_1785);
nor U2905 (N_2905,In_2635,In_2443);
xor U2906 (N_2906,In_1645,In_292);
and U2907 (N_2907,In_783,In_2558);
and U2908 (N_2908,In_2905,In_1416);
and U2909 (N_2909,In_2130,In_2945);
nand U2910 (N_2910,In_766,In_2927);
and U2911 (N_2911,In_2771,In_907);
and U2912 (N_2912,In_1390,In_593);
or U2913 (N_2913,In_2483,In_650);
and U2914 (N_2914,In_2778,In_2337);
nand U2915 (N_2915,In_2191,In_298);
nand U2916 (N_2916,In_2598,In_604);
and U2917 (N_2917,In_542,In_2589);
xnor U2918 (N_2918,In_85,In_2901);
nor U2919 (N_2919,In_1481,In_1967);
nor U2920 (N_2920,In_1786,In_2892);
nand U2921 (N_2921,In_1870,In_971);
and U2922 (N_2922,In_104,In_2570);
nor U2923 (N_2923,In_1081,In_919);
xnor U2924 (N_2924,In_1203,In_1806);
or U2925 (N_2925,In_1778,In_1517);
nand U2926 (N_2926,In_2090,In_1228);
or U2927 (N_2927,In_764,In_1723);
or U2928 (N_2928,In_217,In_339);
and U2929 (N_2929,In_2951,In_1226);
and U2930 (N_2930,In_655,In_1509);
xnor U2931 (N_2931,In_581,In_2249);
nor U2932 (N_2932,In_118,In_352);
nor U2933 (N_2933,In_1251,In_2308);
or U2934 (N_2934,In_454,In_1851);
and U2935 (N_2935,In_2175,In_548);
nor U2936 (N_2936,In_1796,In_1684);
and U2937 (N_2937,In_372,In_2165);
nand U2938 (N_2938,In_1206,In_382);
xnor U2939 (N_2939,In_1256,In_2530);
or U2940 (N_2940,In_2882,In_650);
nand U2941 (N_2941,In_1421,In_1942);
xnor U2942 (N_2942,In_2368,In_703);
xnor U2943 (N_2943,In_1528,In_832);
or U2944 (N_2944,In_892,In_2322);
nor U2945 (N_2945,In_2151,In_2033);
or U2946 (N_2946,In_2102,In_607);
and U2947 (N_2947,In_2939,In_1927);
nor U2948 (N_2948,In_676,In_1485);
nor U2949 (N_2949,In_55,In_1211);
xnor U2950 (N_2950,In_1678,In_2222);
nor U2951 (N_2951,In_412,In_1251);
xor U2952 (N_2952,In_2559,In_2436);
nor U2953 (N_2953,In_2789,In_1576);
or U2954 (N_2954,In_2125,In_2079);
nand U2955 (N_2955,In_720,In_230);
nor U2956 (N_2956,In_2138,In_1987);
nor U2957 (N_2957,In_506,In_1081);
and U2958 (N_2958,In_1254,In_1850);
xnor U2959 (N_2959,In_748,In_1135);
and U2960 (N_2960,In_2279,In_838);
and U2961 (N_2961,In_1414,In_207);
xnor U2962 (N_2962,In_2837,In_1397);
xnor U2963 (N_2963,In_2310,In_2992);
or U2964 (N_2964,In_2472,In_1639);
or U2965 (N_2965,In_2700,In_266);
or U2966 (N_2966,In_972,In_2459);
and U2967 (N_2967,In_802,In_2525);
xnor U2968 (N_2968,In_1742,In_998);
nor U2969 (N_2969,In_2067,In_1045);
or U2970 (N_2970,In_1543,In_2278);
nor U2971 (N_2971,In_1767,In_1162);
or U2972 (N_2972,In_1256,In_2559);
nand U2973 (N_2973,In_928,In_380);
xor U2974 (N_2974,In_2426,In_2241);
xnor U2975 (N_2975,In_877,In_2845);
xor U2976 (N_2976,In_925,In_1435);
and U2977 (N_2977,In_817,In_1506);
or U2978 (N_2978,In_1150,In_2207);
nor U2979 (N_2979,In_643,In_1224);
nor U2980 (N_2980,In_2193,In_228);
xnor U2981 (N_2981,In_167,In_931);
nand U2982 (N_2982,In_549,In_2502);
nand U2983 (N_2983,In_271,In_2002);
nor U2984 (N_2984,In_1548,In_452);
or U2985 (N_2985,In_1902,In_2829);
nand U2986 (N_2986,In_2271,In_2284);
nand U2987 (N_2987,In_2891,In_2099);
nor U2988 (N_2988,In_2829,In_1577);
and U2989 (N_2989,In_2229,In_2810);
xor U2990 (N_2990,In_154,In_2553);
or U2991 (N_2991,In_1343,In_1043);
nor U2992 (N_2992,In_1358,In_1111);
or U2993 (N_2993,In_1852,In_44);
nor U2994 (N_2994,In_11,In_1588);
xor U2995 (N_2995,In_1058,In_518);
xnor U2996 (N_2996,In_1888,In_2741);
nand U2997 (N_2997,In_10,In_1109);
and U2998 (N_2998,In_1166,In_1098);
or U2999 (N_2999,In_1825,In_613);
and U3000 (N_3000,In_1664,In_1626);
xnor U3001 (N_3001,In_1256,In_1453);
and U3002 (N_3002,In_494,In_254);
and U3003 (N_3003,In_462,In_2448);
xnor U3004 (N_3004,In_1443,In_1395);
or U3005 (N_3005,In_2215,In_2513);
xor U3006 (N_3006,In_1755,In_2472);
xor U3007 (N_3007,In_17,In_1196);
and U3008 (N_3008,In_1841,In_969);
xor U3009 (N_3009,In_625,In_605);
xnor U3010 (N_3010,In_521,In_2189);
nand U3011 (N_3011,In_1180,In_2629);
or U3012 (N_3012,In_211,In_1128);
nor U3013 (N_3013,In_2100,In_2532);
xnor U3014 (N_3014,In_17,In_2369);
xnor U3015 (N_3015,In_1927,In_2771);
nor U3016 (N_3016,In_1733,In_2612);
nand U3017 (N_3017,In_1045,In_2176);
xnor U3018 (N_3018,In_1898,In_2496);
xnor U3019 (N_3019,In_1248,In_2956);
nand U3020 (N_3020,In_770,In_660);
xor U3021 (N_3021,In_772,In_494);
nor U3022 (N_3022,In_1153,In_909);
and U3023 (N_3023,In_2831,In_84);
or U3024 (N_3024,In_870,In_1497);
and U3025 (N_3025,In_718,In_612);
xor U3026 (N_3026,In_2552,In_469);
or U3027 (N_3027,In_2133,In_1834);
or U3028 (N_3028,In_1818,In_394);
or U3029 (N_3029,In_1063,In_2887);
and U3030 (N_3030,In_90,In_1982);
nand U3031 (N_3031,In_2341,In_1331);
nand U3032 (N_3032,In_1094,In_200);
or U3033 (N_3033,In_2411,In_764);
xnor U3034 (N_3034,In_62,In_395);
nand U3035 (N_3035,In_2059,In_2026);
or U3036 (N_3036,In_1267,In_774);
nor U3037 (N_3037,In_2482,In_957);
nand U3038 (N_3038,In_1751,In_2499);
nand U3039 (N_3039,In_1256,In_551);
xnor U3040 (N_3040,In_2243,In_6);
xor U3041 (N_3041,In_768,In_892);
xor U3042 (N_3042,In_1469,In_1414);
and U3043 (N_3043,In_2190,In_2116);
nand U3044 (N_3044,In_349,In_2947);
and U3045 (N_3045,In_1697,In_562);
nor U3046 (N_3046,In_448,In_2933);
nand U3047 (N_3047,In_846,In_2645);
nand U3048 (N_3048,In_2613,In_2533);
or U3049 (N_3049,In_2930,In_478);
xor U3050 (N_3050,In_2405,In_2711);
nand U3051 (N_3051,In_2104,In_2087);
nor U3052 (N_3052,In_754,In_2803);
or U3053 (N_3053,In_1809,In_464);
nor U3054 (N_3054,In_1800,In_2183);
and U3055 (N_3055,In_182,In_564);
nand U3056 (N_3056,In_2669,In_2528);
nand U3057 (N_3057,In_387,In_1086);
nor U3058 (N_3058,In_567,In_1673);
and U3059 (N_3059,In_1461,In_1914);
xnor U3060 (N_3060,In_192,In_1545);
nor U3061 (N_3061,In_2990,In_2612);
nand U3062 (N_3062,In_531,In_987);
or U3063 (N_3063,In_1336,In_2691);
nor U3064 (N_3064,In_2704,In_791);
xnor U3065 (N_3065,In_2466,In_2135);
and U3066 (N_3066,In_2909,In_1541);
and U3067 (N_3067,In_1532,In_143);
nor U3068 (N_3068,In_932,In_682);
nor U3069 (N_3069,In_1287,In_841);
xor U3070 (N_3070,In_2088,In_2336);
xnor U3071 (N_3071,In_2498,In_2349);
nor U3072 (N_3072,In_1141,In_2293);
nand U3073 (N_3073,In_469,In_2582);
or U3074 (N_3074,In_2423,In_2038);
nor U3075 (N_3075,In_1167,In_1260);
or U3076 (N_3076,In_719,In_2252);
or U3077 (N_3077,In_770,In_605);
nor U3078 (N_3078,In_438,In_2437);
xnor U3079 (N_3079,In_1706,In_470);
nand U3080 (N_3080,In_944,In_2086);
nor U3081 (N_3081,In_1911,In_2832);
xor U3082 (N_3082,In_1195,In_2473);
xnor U3083 (N_3083,In_2559,In_65);
nor U3084 (N_3084,In_2074,In_890);
nand U3085 (N_3085,In_424,In_2224);
nand U3086 (N_3086,In_2764,In_2712);
or U3087 (N_3087,In_189,In_1550);
or U3088 (N_3088,In_1859,In_823);
xor U3089 (N_3089,In_2642,In_393);
nand U3090 (N_3090,In_2959,In_2392);
or U3091 (N_3091,In_1906,In_207);
nor U3092 (N_3092,In_564,In_734);
or U3093 (N_3093,In_385,In_81);
and U3094 (N_3094,In_573,In_1842);
and U3095 (N_3095,In_21,In_2446);
xor U3096 (N_3096,In_1956,In_1470);
and U3097 (N_3097,In_2693,In_271);
and U3098 (N_3098,In_645,In_2297);
nand U3099 (N_3099,In_616,In_2654);
nor U3100 (N_3100,In_2996,In_1979);
and U3101 (N_3101,In_13,In_2242);
and U3102 (N_3102,In_1757,In_1475);
xor U3103 (N_3103,In_933,In_44);
or U3104 (N_3104,In_1706,In_1554);
xor U3105 (N_3105,In_1581,In_2136);
nor U3106 (N_3106,In_1785,In_2544);
or U3107 (N_3107,In_312,In_1466);
nand U3108 (N_3108,In_502,In_2091);
nand U3109 (N_3109,In_1778,In_412);
or U3110 (N_3110,In_2233,In_1224);
xor U3111 (N_3111,In_1150,In_1305);
xnor U3112 (N_3112,In_1400,In_220);
xor U3113 (N_3113,In_1159,In_566);
nand U3114 (N_3114,In_168,In_81);
nor U3115 (N_3115,In_1775,In_2566);
nand U3116 (N_3116,In_513,In_1618);
nand U3117 (N_3117,In_629,In_2093);
xor U3118 (N_3118,In_1181,In_1563);
nand U3119 (N_3119,In_1621,In_407);
and U3120 (N_3120,In_27,In_2895);
xnor U3121 (N_3121,In_1957,In_775);
or U3122 (N_3122,In_2210,In_2194);
or U3123 (N_3123,In_2970,In_1868);
or U3124 (N_3124,In_1297,In_1604);
or U3125 (N_3125,In_2605,In_2975);
or U3126 (N_3126,In_2071,In_2410);
nor U3127 (N_3127,In_2979,In_722);
nand U3128 (N_3128,In_1620,In_2369);
xor U3129 (N_3129,In_936,In_2022);
or U3130 (N_3130,In_1486,In_2257);
xnor U3131 (N_3131,In_2617,In_903);
nor U3132 (N_3132,In_1863,In_2644);
nor U3133 (N_3133,In_2283,In_2824);
nand U3134 (N_3134,In_110,In_2571);
nand U3135 (N_3135,In_2260,In_2636);
or U3136 (N_3136,In_1796,In_1134);
and U3137 (N_3137,In_767,In_2849);
nand U3138 (N_3138,In_1008,In_508);
nor U3139 (N_3139,In_70,In_2382);
xor U3140 (N_3140,In_2701,In_2364);
nor U3141 (N_3141,In_2185,In_2283);
nand U3142 (N_3142,In_2184,In_2870);
nand U3143 (N_3143,In_2064,In_2813);
nor U3144 (N_3144,In_205,In_561);
xnor U3145 (N_3145,In_2913,In_60);
and U3146 (N_3146,In_2140,In_2079);
xor U3147 (N_3147,In_335,In_158);
xnor U3148 (N_3148,In_2586,In_2980);
and U3149 (N_3149,In_1022,In_1817);
or U3150 (N_3150,In_1310,In_1855);
nor U3151 (N_3151,In_1683,In_2842);
xnor U3152 (N_3152,In_792,In_1068);
nor U3153 (N_3153,In_2541,In_884);
nor U3154 (N_3154,In_1855,In_2580);
or U3155 (N_3155,In_2101,In_2754);
xor U3156 (N_3156,In_2515,In_372);
or U3157 (N_3157,In_1453,In_1765);
or U3158 (N_3158,In_1630,In_1571);
nor U3159 (N_3159,In_1762,In_11);
and U3160 (N_3160,In_879,In_2835);
xor U3161 (N_3161,In_173,In_1188);
nand U3162 (N_3162,In_1027,In_1456);
and U3163 (N_3163,In_1451,In_2832);
and U3164 (N_3164,In_119,In_1914);
nand U3165 (N_3165,In_2082,In_327);
xnor U3166 (N_3166,In_2995,In_1940);
nand U3167 (N_3167,In_2358,In_254);
and U3168 (N_3168,In_2251,In_1823);
or U3169 (N_3169,In_2322,In_2698);
nor U3170 (N_3170,In_1714,In_778);
xnor U3171 (N_3171,In_2481,In_1555);
nor U3172 (N_3172,In_2966,In_1525);
xor U3173 (N_3173,In_1569,In_2840);
or U3174 (N_3174,In_417,In_668);
and U3175 (N_3175,In_1310,In_296);
nand U3176 (N_3176,In_1692,In_363);
and U3177 (N_3177,In_1161,In_2796);
or U3178 (N_3178,In_1629,In_2524);
nand U3179 (N_3179,In_204,In_2475);
nand U3180 (N_3180,In_790,In_15);
nor U3181 (N_3181,In_481,In_59);
nor U3182 (N_3182,In_446,In_2771);
nand U3183 (N_3183,In_1918,In_1263);
or U3184 (N_3184,In_2237,In_1988);
and U3185 (N_3185,In_1567,In_882);
or U3186 (N_3186,In_1409,In_2156);
or U3187 (N_3187,In_772,In_2106);
or U3188 (N_3188,In_2910,In_2551);
and U3189 (N_3189,In_281,In_1550);
xor U3190 (N_3190,In_514,In_2070);
xnor U3191 (N_3191,In_2828,In_1398);
xnor U3192 (N_3192,In_613,In_1972);
or U3193 (N_3193,In_1091,In_1139);
nand U3194 (N_3194,In_676,In_15);
or U3195 (N_3195,In_2003,In_2463);
and U3196 (N_3196,In_1398,In_1867);
nor U3197 (N_3197,In_2505,In_2223);
or U3198 (N_3198,In_845,In_2393);
nor U3199 (N_3199,In_2302,In_1935);
and U3200 (N_3200,In_1973,In_2385);
nand U3201 (N_3201,In_1774,In_2227);
nand U3202 (N_3202,In_1391,In_2831);
nand U3203 (N_3203,In_2972,In_706);
or U3204 (N_3204,In_2810,In_1949);
and U3205 (N_3205,In_502,In_824);
and U3206 (N_3206,In_976,In_1946);
nor U3207 (N_3207,In_459,In_2521);
or U3208 (N_3208,In_2514,In_642);
nand U3209 (N_3209,In_602,In_2935);
nand U3210 (N_3210,In_1445,In_1901);
xnor U3211 (N_3211,In_2791,In_2663);
nand U3212 (N_3212,In_2772,In_1298);
and U3213 (N_3213,In_2704,In_128);
nor U3214 (N_3214,In_1533,In_2047);
nand U3215 (N_3215,In_95,In_926);
nand U3216 (N_3216,In_2308,In_896);
xnor U3217 (N_3217,In_1733,In_1541);
or U3218 (N_3218,In_1737,In_2385);
xor U3219 (N_3219,In_1481,In_532);
xor U3220 (N_3220,In_1929,In_2721);
nor U3221 (N_3221,In_755,In_1891);
nor U3222 (N_3222,In_888,In_925);
and U3223 (N_3223,In_1831,In_1883);
nor U3224 (N_3224,In_2336,In_2670);
nand U3225 (N_3225,In_148,In_880);
or U3226 (N_3226,In_1415,In_1665);
nand U3227 (N_3227,In_1836,In_1934);
nand U3228 (N_3228,In_1497,In_696);
xor U3229 (N_3229,In_1162,In_1964);
nand U3230 (N_3230,In_3,In_460);
nor U3231 (N_3231,In_743,In_81);
xnor U3232 (N_3232,In_1262,In_480);
nand U3233 (N_3233,In_928,In_1966);
nor U3234 (N_3234,In_1705,In_862);
xor U3235 (N_3235,In_2099,In_2330);
xor U3236 (N_3236,In_909,In_421);
nor U3237 (N_3237,In_1336,In_33);
and U3238 (N_3238,In_2676,In_2759);
xnor U3239 (N_3239,In_2229,In_2236);
xnor U3240 (N_3240,In_2439,In_1708);
and U3241 (N_3241,In_66,In_1389);
or U3242 (N_3242,In_1690,In_2998);
or U3243 (N_3243,In_131,In_1913);
and U3244 (N_3244,In_1583,In_1499);
or U3245 (N_3245,In_2495,In_2483);
nand U3246 (N_3246,In_1157,In_2189);
nand U3247 (N_3247,In_1332,In_367);
or U3248 (N_3248,In_1470,In_647);
xor U3249 (N_3249,In_2577,In_217);
nand U3250 (N_3250,In_462,In_1911);
and U3251 (N_3251,In_1411,In_1180);
xnor U3252 (N_3252,In_625,In_1936);
nor U3253 (N_3253,In_486,In_1428);
or U3254 (N_3254,In_1855,In_148);
or U3255 (N_3255,In_210,In_1539);
xor U3256 (N_3256,In_1565,In_1623);
and U3257 (N_3257,In_2544,In_653);
and U3258 (N_3258,In_348,In_1653);
nand U3259 (N_3259,In_2623,In_2141);
or U3260 (N_3260,In_1953,In_777);
and U3261 (N_3261,In_2924,In_525);
xnor U3262 (N_3262,In_1984,In_1323);
xnor U3263 (N_3263,In_1218,In_1849);
nor U3264 (N_3264,In_1461,In_2174);
or U3265 (N_3265,In_1033,In_64);
nand U3266 (N_3266,In_2916,In_2915);
xor U3267 (N_3267,In_2051,In_562);
or U3268 (N_3268,In_1053,In_2468);
xor U3269 (N_3269,In_215,In_2414);
nor U3270 (N_3270,In_909,In_2288);
nand U3271 (N_3271,In_926,In_920);
nand U3272 (N_3272,In_344,In_2294);
xor U3273 (N_3273,In_748,In_1129);
xnor U3274 (N_3274,In_2495,In_588);
and U3275 (N_3275,In_1951,In_2400);
nand U3276 (N_3276,In_568,In_2681);
and U3277 (N_3277,In_905,In_1126);
nand U3278 (N_3278,In_593,In_761);
nor U3279 (N_3279,In_2982,In_1087);
and U3280 (N_3280,In_1649,In_1625);
xor U3281 (N_3281,In_985,In_511);
nand U3282 (N_3282,In_881,In_924);
xor U3283 (N_3283,In_2762,In_2420);
xor U3284 (N_3284,In_2056,In_971);
or U3285 (N_3285,In_1557,In_2217);
and U3286 (N_3286,In_1385,In_283);
xnor U3287 (N_3287,In_1023,In_2608);
xnor U3288 (N_3288,In_2359,In_2353);
nor U3289 (N_3289,In_848,In_2992);
nor U3290 (N_3290,In_2316,In_2400);
nand U3291 (N_3291,In_750,In_1802);
or U3292 (N_3292,In_2597,In_1617);
or U3293 (N_3293,In_559,In_422);
nor U3294 (N_3294,In_785,In_2961);
and U3295 (N_3295,In_138,In_2396);
or U3296 (N_3296,In_2871,In_2277);
and U3297 (N_3297,In_2271,In_2200);
and U3298 (N_3298,In_1541,In_1650);
or U3299 (N_3299,In_603,In_1386);
nor U3300 (N_3300,In_2850,In_556);
nor U3301 (N_3301,In_135,In_2868);
nand U3302 (N_3302,In_2208,In_2183);
or U3303 (N_3303,In_2172,In_2323);
nor U3304 (N_3304,In_623,In_1164);
and U3305 (N_3305,In_926,In_2002);
nand U3306 (N_3306,In_191,In_474);
nand U3307 (N_3307,In_724,In_172);
nor U3308 (N_3308,In_1710,In_1383);
nor U3309 (N_3309,In_343,In_2243);
and U3310 (N_3310,In_580,In_2414);
and U3311 (N_3311,In_2572,In_880);
or U3312 (N_3312,In_396,In_1442);
nor U3313 (N_3313,In_748,In_2855);
nand U3314 (N_3314,In_312,In_2548);
or U3315 (N_3315,In_1062,In_1331);
xor U3316 (N_3316,In_2122,In_1271);
nor U3317 (N_3317,In_1206,In_2323);
and U3318 (N_3318,In_994,In_1172);
nor U3319 (N_3319,In_47,In_2178);
nor U3320 (N_3320,In_360,In_1386);
or U3321 (N_3321,In_2357,In_613);
or U3322 (N_3322,In_1075,In_2636);
and U3323 (N_3323,In_1095,In_1904);
or U3324 (N_3324,In_130,In_1549);
and U3325 (N_3325,In_2730,In_2983);
or U3326 (N_3326,In_862,In_2638);
nand U3327 (N_3327,In_2805,In_1223);
and U3328 (N_3328,In_2965,In_835);
and U3329 (N_3329,In_2603,In_692);
nor U3330 (N_3330,In_402,In_2626);
or U3331 (N_3331,In_2440,In_1848);
nor U3332 (N_3332,In_2819,In_57);
and U3333 (N_3333,In_1208,In_1128);
or U3334 (N_3334,In_372,In_1654);
or U3335 (N_3335,In_1685,In_1213);
and U3336 (N_3336,In_1447,In_1314);
nand U3337 (N_3337,In_306,In_2993);
xor U3338 (N_3338,In_705,In_2299);
nand U3339 (N_3339,In_1893,In_20);
nor U3340 (N_3340,In_371,In_249);
or U3341 (N_3341,In_662,In_2042);
and U3342 (N_3342,In_224,In_2421);
xor U3343 (N_3343,In_2347,In_2365);
nand U3344 (N_3344,In_179,In_1260);
or U3345 (N_3345,In_2917,In_1379);
or U3346 (N_3346,In_1893,In_2838);
nand U3347 (N_3347,In_1128,In_2743);
xor U3348 (N_3348,In_2334,In_249);
nor U3349 (N_3349,In_2424,In_184);
nor U3350 (N_3350,In_2030,In_2231);
xnor U3351 (N_3351,In_1686,In_1129);
nor U3352 (N_3352,In_887,In_2286);
or U3353 (N_3353,In_1142,In_828);
or U3354 (N_3354,In_588,In_2951);
or U3355 (N_3355,In_1262,In_679);
nand U3356 (N_3356,In_2117,In_1784);
and U3357 (N_3357,In_2312,In_447);
nand U3358 (N_3358,In_1270,In_407);
or U3359 (N_3359,In_2166,In_853);
nand U3360 (N_3360,In_2157,In_48);
or U3361 (N_3361,In_485,In_1036);
or U3362 (N_3362,In_1273,In_471);
and U3363 (N_3363,In_2616,In_2685);
nand U3364 (N_3364,In_1837,In_1631);
nand U3365 (N_3365,In_97,In_2118);
or U3366 (N_3366,In_1736,In_2851);
nor U3367 (N_3367,In_1377,In_2906);
and U3368 (N_3368,In_1797,In_1423);
nand U3369 (N_3369,In_2805,In_2380);
nor U3370 (N_3370,In_2289,In_1808);
nor U3371 (N_3371,In_833,In_929);
or U3372 (N_3372,In_1276,In_1481);
nor U3373 (N_3373,In_281,In_2085);
nor U3374 (N_3374,In_214,In_2110);
nand U3375 (N_3375,In_15,In_646);
nand U3376 (N_3376,In_1508,In_464);
or U3377 (N_3377,In_39,In_1416);
nor U3378 (N_3378,In_121,In_522);
nand U3379 (N_3379,In_469,In_2158);
nand U3380 (N_3380,In_1474,In_2701);
xor U3381 (N_3381,In_2721,In_602);
or U3382 (N_3382,In_2,In_636);
and U3383 (N_3383,In_755,In_2858);
and U3384 (N_3384,In_918,In_832);
nand U3385 (N_3385,In_2194,In_2186);
and U3386 (N_3386,In_1897,In_694);
nor U3387 (N_3387,In_2781,In_1472);
xor U3388 (N_3388,In_1751,In_2168);
or U3389 (N_3389,In_1103,In_2737);
or U3390 (N_3390,In_2219,In_2628);
nor U3391 (N_3391,In_92,In_2980);
and U3392 (N_3392,In_1060,In_694);
and U3393 (N_3393,In_2658,In_2695);
and U3394 (N_3394,In_484,In_2249);
nand U3395 (N_3395,In_2689,In_2914);
nor U3396 (N_3396,In_2550,In_1277);
or U3397 (N_3397,In_1104,In_1822);
nor U3398 (N_3398,In_583,In_1022);
and U3399 (N_3399,In_2959,In_2268);
or U3400 (N_3400,In_1639,In_1595);
nand U3401 (N_3401,In_837,In_2332);
or U3402 (N_3402,In_1051,In_553);
or U3403 (N_3403,In_1795,In_1173);
nand U3404 (N_3404,In_280,In_1726);
xor U3405 (N_3405,In_406,In_752);
and U3406 (N_3406,In_1781,In_1398);
nor U3407 (N_3407,In_494,In_1748);
xor U3408 (N_3408,In_1751,In_1482);
xor U3409 (N_3409,In_2189,In_1090);
xnor U3410 (N_3410,In_2388,In_2341);
xnor U3411 (N_3411,In_1006,In_2350);
xor U3412 (N_3412,In_1324,In_2667);
or U3413 (N_3413,In_1270,In_2408);
nor U3414 (N_3414,In_800,In_397);
nand U3415 (N_3415,In_2941,In_1234);
nand U3416 (N_3416,In_249,In_1839);
or U3417 (N_3417,In_2620,In_290);
nor U3418 (N_3418,In_2912,In_412);
nor U3419 (N_3419,In_2067,In_515);
nand U3420 (N_3420,In_2815,In_2987);
nor U3421 (N_3421,In_2335,In_2253);
and U3422 (N_3422,In_1265,In_2514);
and U3423 (N_3423,In_1901,In_1053);
nand U3424 (N_3424,In_899,In_1382);
and U3425 (N_3425,In_913,In_793);
xor U3426 (N_3426,In_2746,In_297);
and U3427 (N_3427,In_2261,In_915);
and U3428 (N_3428,In_354,In_1115);
xnor U3429 (N_3429,In_1702,In_661);
nor U3430 (N_3430,In_1675,In_2021);
nand U3431 (N_3431,In_2383,In_2856);
xor U3432 (N_3432,In_2536,In_1418);
or U3433 (N_3433,In_1918,In_576);
and U3434 (N_3434,In_2455,In_1759);
xor U3435 (N_3435,In_1218,In_1679);
nand U3436 (N_3436,In_689,In_617);
or U3437 (N_3437,In_1880,In_355);
nor U3438 (N_3438,In_2431,In_1288);
xnor U3439 (N_3439,In_1463,In_795);
nand U3440 (N_3440,In_2947,In_2519);
nand U3441 (N_3441,In_1845,In_340);
xnor U3442 (N_3442,In_1744,In_2400);
nor U3443 (N_3443,In_90,In_1909);
or U3444 (N_3444,In_313,In_2538);
xnor U3445 (N_3445,In_2584,In_2080);
nand U3446 (N_3446,In_1305,In_2710);
xor U3447 (N_3447,In_850,In_598);
or U3448 (N_3448,In_2780,In_2896);
xnor U3449 (N_3449,In_1545,In_2057);
xnor U3450 (N_3450,In_2364,In_605);
nand U3451 (N_3451,In_63,In_1104);
nand U3452 (N_3452,In_1351,In_1223);
nor U3453 (N_3453,In_1998,In_1018);
nor U3454 (N_3454,In_2526,In_65);
xnor U3455 (N_3455,In_2948,In_813);
or U3456 (N_3456,In_2044,In_122);
nand U3457 (N_3457,In_924,In_886);
or U3458 (N_3458,In_1161,In_372);
xor U3459 (N_3459,In_2779,In_2852);
or U3460 (N_3460,In_758,In_1753);
and U3461 (N_3461,In_2401,In_1024);
nor U3462 (N_3462,In_411,In_1137);
and U3463 (N_3463,In_439,In_1622);
and U3464 (N_3464,In_1845,In_2556);
or U3465 (N_3465,In_1684,In_634);
nor U3466 (N_3466,In_1520,In_2106);
and U3467 (N_3467,In_81,In_1197);
nor U3468 (N_3468,In_803,In_1669);
xor U3469 (N_3469,In_397,In_1128);
nand U3470 (N_3470,In_2665,In_576);
nor U3471 (N_3471,In_1129,In_1003);
xor U3472 (N_3472,In_1412,In_1300);
or U3473 (N_3473,In_2575,In_338);
xnor U3474 (N_3474,In_1174,In_294);
xor U3475 (N_3475,In_2584,In_42);
or U3476 (N_3476,In_1854,In_2846);
and U3477 (N_3477,In_2940,In_1464);
xor U3478 (N_3478,In_1924,In_2941);
and U3479 (N_3479,In_533,In_2132);
xor U3480 (N_3480,In_1080,In_1823);
or U3481 (N_3481,In_1049,In_991);
xnor U3482 (N_3482,In_2846,In_1600);
nand U3483 (N_3483,In_343,In_1819);
or U3484 (N_3484,In_1454,In_337);
nor U3485 (N_3485,In_1051,In_2029);
and U3486 (N_3486,In_2718,In_2615);
nand U3487 (N_3487,In_316,In_1602);
xor U3488 (N_3488,In_2242,In_699);
or U3489 (N_3489,In_2636,In_1794);
or U3490 (N_3490,In_662,In_1001);
or U3491 (N_3491,In_2780,In_2298);
and U3492 (N_3492,In_1904,In_21);
or U3493 (N_3493,In_136,In_716);
xnor U3494 (N_3494,In_1006,In_1286);
and U3495 (N_3495,In_888,In_2763);
and U3496 (N_3496,In_643,In_2499);
nand U3497 (N_3497,In_972,In_1423);
nor U3498 (N_3498,In_1826,In_834);
or U3499 (N_3499,In_1602,In_2219);
xor U3500 (N_3500,In_1126,In_2237);
or U3501 (N_3501,In_1464,In_1721);
or U3502 (N_3502,In_2249,In_131);
and U3503 (N_3503,In_1279,In_1106);
or U3504 (N_3504,In_1290,In_2971);
or U3505 (N_3505,In_2874,In_116);
and U3506 (N_3506,In_168,In_390);
and U3507 (N_3507,In_2697,In_2985);
nor U3508 (N_3508,In_670,In_1988);
xnor U3509 (N_3509,In_1771,In_1642);
nand U3510 (N_3510,In_1569,In_2297);
nand U3511 (N_3511,In_73,In_564);
or U3512 (N_3512,In_1669,In_1716);
or U3513 (N_3513,In_2532,In_2318);
xor U3514 (N_3514,In_1383,In_666);
and U3515 (N_3515,In_2899,In_2339);
or U3516 (N_3516,In_2177,In_2646);
nor U3517 (N_3517,In_291,In_751);
or U3518 (N_3518,In_2419,In_920);
nand U3519 (N_3519,In_110,In_2782);
nand U3520 (N_3520,In_2077,In_2822);
nor U3521 (N_3521,In_2002,In_348);
or U3522 (N_3522,In_552,In_875);
nor U3523 (N_3523,In_2285,In_424);
xor U3524 (N_3524,In_874,In_1122);
and U3525 (N_3525,In_920,In_730);
nor U3526 (N_3526,In_709,In_2444);
nand U3527 (N_3527,In_1530,In_468);
or U3528 (N_3528,In_524,In_821);
nand U3529 (N_3529,In_243,In_1);
or U3530 (N_3530,In_1445,In_608);
xnor U3531 (N_3531,In_2220,In_743);
and U3532 (N_3532,In_2350,In_748);
xor U3533 (N_3533,In_178,In_847);
nand U3534 (N_3534,In_2134,In_2252);
or U3535 (N_3535,In_2975,In_679);
nor U3536 (N_3536,In_2273,In_2031);
nand U3537 (N_3537,In_2099,In_2833);
or U3538 (N_3538,In_970,In_2275);
or U3539 (N_3539,In_2941,In_168);
nand U3540 (N_3540,In_2779,In_303);
or U3541 (N_3541,In_141,In_513);
xnor U3542 (N_3542,In_456,In_1803);
nand U3543 (N_3543,In_2989,In_2314);
or U3544 (N_3544,In_926,In_741);
and U3545 (N_3545,In_213,In_1359);
or U3546 (N_3546,In_1013,In_118);
nor U3547 (N_3547,In_2544,In_1828);
xor U3548 (N_3548,In_2756,In_2582);
nand U3549 (N_3549,In_555,In_1762);
and U3550 (N_3550,In_2940,In_2416);
nor U3551 (N_3551,In_1351,In_915);
or U3552 (N_3552,In_812,In_1925);
nor U3553 (N_3553,In_70,In_2250);
xor U3554 (N_3554,In_584,In_661);
nand U3555 (N_3555,In_1759,In_1634);
nand U3556 (N_3556,In_2375,In_2854);
xnor U3557 (N_3557,In_2625,In_2251);
xnor U3558 (N_3558,In_1140,In_2301);
nand U3559 (N_3559,In_1993,In_198);
xnor U3560 (N_3560,In_2519,In_2518);
nand U3561 (N_3561,In_1751,In_1159);
xor U3562 (N_3562,In_2220,In_2299);
xor U3563 (N_3563,In_1990,In_2140);
and U3564 (N_3564,In_957,In_923);
or U3565 (N_3565,In_1471,In_442);
xnor U3566 (N_3566,In_2476,In_2986);
or U3567 (N_3567,In_1606,In_338);
or U3568 (N_3568,In_230,In_1403);
and U3569 (N_3569,In_794,In_1849);
xnor U3570 (N_3570,In_844,In_1837);
nor U3571 (N_3571,In_303,In_2666);
nor U3572 (N_3572,In_1466,In_762);
or U3573 (N_3573,In_428,In_745);
xnor U3574 (N_3574,In_53,In_2935);
xor U3575 (N_3575,In_922,In_1793);
nand U3576 (N_3576,In_590,In_1727);
xnor U3577 (N_3577,In_746,In_1514);
and U3578 (N_3578,In_2467,In_527);
xnor U3579 (N_3579,In_1127,In_1248);
nor U3580 (N_3580,In_2714,In_1833);
or U3581 (N_3581,In_332,In_423);
nand U3582 (N_3582,In_1395,In_2535);
or U3583 (N_3583,In_1760,In_176);
or U3584 (N_3584,In_2892,In_1864);
nand U3585 (N_3585,In_1685,In_1517);
nor U3586 (N_3586,In_2340,In_1063);
nor U3587 (N_3587,In_1595,In_544);
and U3588 (N_3588,In_59,In_57);
or U3589 (N_3589,In_897,In_2161);
nor U3590 (N_3590,In_1294,In_2415);
nor U3591 (N_3591,In_2638,In_1946);
xor U3592 (N_3592,In_1649,In_632);
xnor U3593 (N_3593,In_106,In_35);
or U3594 (N_3594,In_2677,In_1301);
nand U3595 (N_3595,In_235,In_1327);
xor U3596 (N_3596,In_964,In_2995);
and U3597 (N_3597,In_421,In_1429);
nor U3598 (N_3598,In_203,In_2540);
nand U3599 (N_3599,In_2059,In_1859);
or U3600 (N_3600,In_2570,In_2841);
nand U3601 (N_3601,In_1314,In_201);
xnor U3602 (N_3602,In_2393,In_150);
or U3603 (N_3603,In_1772,In_2029);
or U3604 (N_3604,In_2821,In_2648);
and U3605 (N_3605,In_573,In_584);
and U3606 (N_3606,In_2422,In_706);
nor U3607 (N_3607,In_624,In_2743);
xor U3608 (N_3608,In_1196,In_1376);
and U3609 (N_3609,In_1162,In_1170);
nand U3610 (N_3610,In_378,In_2216);
nor U3611 (N_3611,In_2107,In_1933);
or U3612 (N_3612,In_686,In_1639);
xor U3613 (N_3613,In_2421,In_2591);
and U3614 (N_3614,In_900,In_1025);
nand U3615 (N_3615,In_2524,In_30);
or U3616 (N_3616,In_1128,In_2866);
or U3617 (N_3617,In_1372,In_2200);
nor U3618 (N_3618,In_2722,In_2186);
nand U3619 (N_3619,In_1897,In_1730);
nand U3620 (N_3620,In_2208,In_574);
nand U3621 (N_3621,In_285,In_2445);
and U3622 (N_3622,In_2770,In_2672);
or U3623 (N_3623,In_2633,In_2922);
nand U3624 (N_3624,In_983,In_1291);
nor U3625 (N_3625,In_69,In_1124);
xor U3626 (N_3626,In_1223,In_2557);
xnor U3627 (N_3627,In_1490,In_1517);
and U3628 (N_3628,In_2954,In_1373);
nor U3629 (N_3629,In_2467,In_1403);
and U3630 (N_3630,In_2803,In_2799);
nand U3631 (N_3631,In_1162,In_217);
nand U3632 (N_3632,In_2726,In_2828);
and U3633 (N_3633,In_2522,In_2763);
xnor U3634 (N_3634,In_1007,In_361);
or U3635 (N_3635,In_1184,In_2635);
nor U3636 (N_3636,In_972,In_1113);
nor U3637 (N_3637,In_2478,In_2218);
xnor U3638 (N_3638,In_1446,In_1275);
and U3639 (N_3639,In_1131,In_1491);
xnor U3640 (N_3640,In_1484,In_2639);
nor U3641 (N_3641,In_194,In_1881);
xnor U3642 (N_3642,In_2990,In_1109);
or U3643 (N_3643,In_910,In_1806);
nand U3644 (N_3644,In_1704,In_2996);
or U3645 (N_3645,In_896,In_1176);
and U3646 (N_3646,In_2895,In_1234);
and U3647 (N_3647,In_2718,In_452);
or U3648 (N_3648,In_2339,In_1656);
xnor U3649 (N_3649,In_249,In_2412);
xor U3650 (N_3650,In_2380,In_369);
or U3651 (N_3651,In_0,In_2583);
or U3652 (N_3652,In_1952,In_1921);
and U3653 (N_3653,In_1237,In_827);
or U3654 (N_3654,In_362,In_1627);
or U3655 (N_3655,In_2371,In_409);
nor U3656 (N_3656,In_1123,In_1191);
and U3657 (N_3657,In_952,In_49);
or U3658 (N_3658,In_2341,In_1014);
and U3659 (N_3659,In_2063,In_1311);
xnor U3660 (N_3660,In_990,In_1185);
nor U3661 (N_3661,In_2178,In_1245);
nand U3662 (N_3662,In_1723,In_1576);
nor U3663 (N_3663,In_1982,In_2828);
nor U3664 (N_3664,In_2914,In_474);
and U3665 (N_3665,In_1441,In_1634);
nor U3666 (N_3666,In_212,In_2576);
nand U3667 (N_3667,In_68,In_2773);
and U3668 (N_3668,In_1141,In_955);
or U3669 (N_3669,In_1922,In_2750);
and U3670 (N_3670,In_1221,In_1745);
nor U3671 (N_3671,In_725,In_979);
nor U3672 (N_3672,In_849,In_251);
nand U3673 (N_3673,In_834,In_1312);
or U3674 (N_3674,In_2545,In_1816);
nor U3675 (N_3675,In_1966,In_1668);
or U3676 (N_3676,In_639,In_772);
or U3677 (N_3677,In_621,In_1599);
nand U3678 (N_3678,In_414,In_132);
or U3679 (N_3679,In_2501,In_2892);
or U3680 (N_3680,In_478,In_214);
or U3681 (N_3681,In_2992,In_2777);
nor U3682 (N_3682,In_1142,In_965);
nand U3683 (N_3683,In_1472,In_2421);
and U3684 (N_3684,In_933,In_1478);
nor U3685 (N_3685,In_786,In_1730);
nand U3686 (N_3686,In_2408,In_1763);
nand U3687 (N_3687,In_1566,In_2756);
nor U3688 (N_3688,In_2243,In_481);
nand U3689 (N_3689,In_1492,In_701);
xnor U3690 (N_3690,In_1866,In_2059);
nand U3691 (N_3691,In_305,In_2970);
xnor U3692 (N_3692,In_943,In_1235);
nand U3693 (N_3693,In_2060,In_1846);
xnor U3694 (N_3694,In_2657,In_1651);
nor U3695 (N_3695,In_2143,In_2647);
nor U3696 (N_3696,In_1287,In_731);
and U3697 (N_3697,In_374,In_30);
or U3698 (N_3698,In_1574,In_719);
nand U3699 (N_3699,In_1991,In_906);
nand U3700 (N_3700,In_2264,In_2274);
nand U3701 (N_3701,In_2296,In_474);
nor U3702 (N_3702,In_871,In_2549);
and U3703 (N_3703,In_2146,In_1386);
xnor U3704 (N_3704,In_609,In_2011);
and U3705 (N_3705,In_727,In_2510);
and U3706 (N_3706,In_1832,In_1511);
xor U3707 (N_3707,In_689,In_2978);
nand U3708 (N_3708,In_1161,In_1546);
xor U3709 (N_3709,In_1556,In_1259);
xor U3710 (N_3710,In_834,In_2082);
or U3711 (N_3711,In_2847,In_1366);
nand U3712 (N_3712,In_813,In_850);
nand U3713 (N_3713,In_1481,In_2686);
and U3714 (N_3714,In_1181,In_2100);
nand U3715 (N_3715,In_2357,In_813);
nor U3716 (N_3716,In_330,In_2854);
or U3717 (N_3717,In_826,In_1587);
or U3718 (N_3718,In_2769,In_2011);
and U3719 (N_3719,In_473,In_727);
or U3720 (N_3720,In_1354,In_2457);
nand U3721 (N_3721,In_916,In_2594);
and U3722 (N_3722,In_1050,In_217);
nor U3723 (N_3723,In_2213,In_2468);
nor U3724 (N_3724,In_126,In_2013);
xnor U3725 (N_3725,In_1225,In_1793);
nand U3726 (N_3726,In_562,In_1161);
nand U3727 (N_3727,In_2826,In_880);
xnor U3728 (N_3728,In_2783,In_197);
nor U3729 (N_3729,In_1540,In_2053);
and U3730 (N_3730,In_2187,In_1273);
nor U3731 (N_3731,In_131,In_2113);
and U3732 (N_3732,In_1516,In_1941);
nor U3733 (N_3733,In_534,In_1706);
and U3734 (N_3734,In_2225,In_114);
or U3735 (N_3735,In_2798,In_1784);
nand U3736 (N_3736,In_1921,In_2441);
or U3737 (N_3737,In_1359,In_2110);
nand U3738 (N_3738,In_2637,In_2114);
nor U3739 (N_3739,In_2342,In_2934);
or U3740 (N_3740,In_926,In_722);
xnor U3741 (N_3741,In_847,In_1281);
nand U3742 (N_3742,In_160,In_2199);
or U3743 (N_3743,In_2567,In_1351);
or U3744 (N_3744,In_2993,In_2816);
nand U3745 (N_3745,In_2218,In_1552);
nand U3746 (N_3746,In_2588,In_2623);
nor U3747 (N_3747,In_851,In_234);
nor U3748 (N_3748,In_423,In_782);
nor U3749 (N_3749,In_111,In_1019);
or U3750 (N_3750,In_382,In_840);
xnor U3751 (N_3751,In_2716,In_2885);
nand U3752 (N_3752,In_223,In_1674);
xor U3753 (N_3753,In_1129,In_2413);
or U3754 (N_3754,In_1501,In_1611);
and U3755 (N_3755,In_2752,In_1961);
nand U3756 (N_3756,In_2939,In_477);
xnor U3757 (N_3757,In_687,In_985);
xnor U3758 (N_3758,In_2950,In_1152);
nand U3759 (N_3759,In_2832,In_252);
and U3760 (N_3760,In_2941,In_2375);
and U3761 (N_3761,In_363,In_1614);
or U3762 (N_3762,In_369,In_594);
nand U3763 (N_3763,In_55,In_1425);
xnor U3764 (N_3764,In_1095,In_1183);
nand U3765 (N_3765,In_2946,In_2120);
nand U3766 (N_3766,In_249,In_483);
or U3767 (N_3767,In_2123,In_1358);
xor U3768 (N_3768,In_1049,In_2159);
and U3769 (N_3769,In_2283,In_761);
and U3770 (N_3770,In_2001,In_757);
and U3771 (N_3771,In_1800,In_1753);
nor U3772 (N_3772,In_2443,In_1503);
and U3773 (N_3773,In_189,In_13);
and U3774 (N_3774,In_1010,In_350);
or U3775 (N_3775,In_1747,In_532);
and U3776 (N_3776,In_158,In_2930);
nand U3777 (N_3777,In_1992,In_2950);
xor U3778 (N_3778,In_2481,In_1612);
and U3779 (N_3779,In_2479,In_210);
xnor U3780 (N_3780,In_329,In_1480);
xnor U3781 (N_3781,In_2854,In_2069);
nor U3782 (N_3782,In_2789,In_292);
and U3783 (N_3783,In_1892,In_1684);
or U3784 (N_3784,In_618,In_2048);
nand U3785 (N_3785,In_510,In_788);
nor U3786 (N_3786,In_2099,In_2045);
and U3787 (N_3787,In_1712,In_323);
or U3788 (N_3788,In_1976,In_1701);
nand U3789 (N_3789,In_316,In_620);
xnor U3790 (N_3790,In_1907,In_622);
and U3791 (N_3791,In_574,In_525);
nand U3792 (N_3792,In_2779,In_1400);
and U3793 (N_3793,In_363,In_2346);
nand U3794 (N_3794,In_2425,In_914);
and U3795 (N_3795,In_1418,In_384);
nor U3796 (N_3796,In_2198,In_2359);
xor U3797 (N_3797,In_331,In_1311);
nor U3798 (N_3798,In_2106,In_61);
and U3799 (N_3799,In_322,In_663);
or U3800 (N_3800,In_2906,In_249);
or U3801 (N_3801,In_1454,In_62);
nor U3802 (N_3802,In_324,In_1177);
and U3803 (N_3803,In_1248,In_318);
nor U3804 (N_3804,In_1128,In_268);
or U3805 (N_3805,In_967,In_927);
and U3806 (N_3806,In_1374,In_2887);
nand U3807 (N_3807,In_885,In_2629);
and U3808 (N_3808,In_2700,In_84);
and U3809 (N_3809,In_1250,In_2070);
and U3810 (N_3810,In_1846,In_2912);
or U3811 (N_3811,In_2025,In_1328);
nand U3812 (N_3812,In_2845,In_2631);
nand U3813 (N_3813,In_1729,In_860);
nand U3814 (N_3814,In_999,In_2045);
or U3815 (N_3815,In_987,In_375);
or U3816 (N_3816,In_1772,In_1891);
or U3817 (N_3817,In_2170,In_985);
and U3818 (N_3818,In_871,In_984);
or U3819 (N_3819,In_2352,In_2852);
nor U3820 (N_3820,In_568,In_89);
nand U3821 (N_3821,In_1177,In_785);
or U3822 (N_3822,In_400,In_2713);
xor U3823 (N_3823,In_2683,In_453);
xor U3824 (N_3824,In_2564,In_742);
xor U3825 (N_3825,In_2760,In_795);
nand U3826 (N_3826,In_679,In_1957);
nand U3827 (N_3827,In_487,In_490);
or U3828 (N_3828,In_411,In_557);
nand U3829 (N_3829,In_645,In_396);
xnor U3830 (N_3830,In_791,In_1318);
and U3831 (N_3831,In_2026,In_2835);
and U3832 (N_3832,In_1526,In_63);
nor U3833 (N_3833,In_567,In_2927);
and U3834 (N_3834,In_1210,In_2550);
or U3835 (N_3835,In_1856,In_8);
xor U3836 (N_3836,In_1887,In_1617);
and U3837 (N_3837,In_1111,In_948);
or U3838 (N_3838,In_597,In_97);
or U3839 (N_3839,In_1469,In_1505);
nand U3840 (N_3840,In_1209,In_1231);
or U3841 (N_3841,In_1161,In_1629);
xnor U3842 (N_3842,In_1204,In_1818);
xor U3843 (N_3843,In_1191,In_616);
and U3844 (N_3844,In_2119,In_732);
xor U3845 (N_3845,In_1574,In_1769);
xor U3846 (N_3846,In_1134,In_2511);
nor U3847 (N_3847,In_850,In_1978);
xor U3848 (N_3848,In_1188,In_1422);
nand U3849 (N_3849,In_1587,In_1777);
xnor U3850 (N_3850,In_1067,In_1280);
and U3851 (N_3851,In_2894,In_60);
xnor U3852 (N_3852,In_113,In_1013);
nor U3853 (N_3853,In_1206,In_2215);
and U3854 (N_3854,In_794,In_2948);
xor U3855 (N_3855,In_360,In_1219);
nor U3856 (N_3856,In_1693,In_2282);
or U3857 (N_3857,In_492,In_2729);
and U3858 (N_3858,In_959,In_1416);
xor U3859 (N_3859,In_455,In_526);
nor U3860 (N_3860,In_2804,In_1324);
nand U3861 (N_3861,In_1327,In_973);
xor U3862 (N_3862,In_2050,In_1262);
nand U3863 (N_3863,In_2845,In_1241);
and U3864 (N_3864,In_433,In_232);
and U3865 (N_3865,In_2794,In_1478);
or U3866 (N_3866,In_2526,In_2401);
nand U3867 (N_3867,In_221,In_1782);
nor U3868 (N_3868,In_2428,In_2430);
and U3869 (N_3869,In_1916,In_2142);
xnor U3870 (N_3870,In_1680,In_117);
xnor U3871 (N_3871,In_1322,In_1765);
nor U3872 (N_3872,In_1109,In_1263);
nor U3873 (N_3873,In_1364,In_237);
and U3874 (N_3874,In_2112,In_1567);
nand U3875 (N_3875,In_280,In_2993);
nand U3876 (N_3876,In_2294,In_2512);
or U3877 (N_3877,In_2211,In_480);
nand U3878 (N_3878,In_1855,In_1497);
xor U3879 (N_3879,In_4,In_1678);
nand U3880 (N_3880,In_567,In_1110);
or U3881 (N_3881,In_1532,In_2193);
nor U3882 (N_3882,In_2211,In_2607);
nor U3883 (N_3883,In_1979,In_2956);
and U3884 (N_3884,In_1925,In_1297);
nand U3885 (N_3885,In_2564,In_155);
or U3886 (N_3886,In_2444,In_797);
nor U3887 (N_3887,In_1641,In_345);
and U3888 (N_3888,In_2596,In_1413);
or U3889 (N_3889,In_933,In_514);
and U3890 (N_3890,In_1608,In_2001);
nand U3891 (N_3891,In_77,In_385);
or U3892 (N_3892,In_2036,In_669);
or U3893 (N_3893,In_1953,In_2412);
xor U3894 (N_3894,In_1726,In_865);
and U3895 (N_3895,In_1287,In_2508);
and U3896 (N_3896,In_406,In_955);
nand U3897 (N_3897,In_1751,In_920);
and U3898 (N_3898,In_529,In_2888);
and U3899 (N_3899,In_203,In_991);
xnor U3900 (N_3900,In_2977,In_2375);
nand U3901 (N_3901,In_310,In_776);
nor U3902 (N_3902,In_2302,In_1505);
or U3903 (N_3903,In_341,In_1492);
nor U3904 (N_3904,In_1340,In_2920);
nor U3905 (N_3905,In_1562,In_2807);
nor U3906 (N_3906,In_2671,In_2340);
nand U3907 (N_3907,In_783,In_2309);
or U3908 (N_3908,In_2142,In_80);
or U3909 (N_3909,In_1579,In_1114);
xnor U3910 (N_3910,In_960,In_794);
nand U3911 (N_3911,In_512,In_995);
nand U3912 (N_3912,In_2889,In_145);
nor U3913 (N_3913,In_2110,In_1490);
and U3914 (N_3914,In_2478,In_1887);
nor U3915 (N_3915,In_1398,In_2976);
nand U3916 (N_3916,In_545,In_2696);
xnor U3917 (N_3917,In_2143,In_217);
nand U3918 (N_3918,In_1693,In_2034);
nand U3919 (N_3919,In_775,In_2376);
nor U3920 (N_3920,In_2934,In_2525);
and U3921 (N_3921,In_2448,In_81);
xnor U3922 (N_3922,In_1434,In_2508);
nand U3923 (N_3923,In_1747,In_1163);
nand U3924 (N_3924,In_1998,In_1786);
or U3925 (N_3925,In_415,In_319);
or U3926 (N_3926,In_162,In_1051);
xor U3927 (N_3927,In_776,In_709);
nor U3928 (N_3928,In_2276,In_707);
nor U3929 (N_3929,In_148,In_2171);
nand U3930 (N_3930,In_1691,In_2859);
nand U3931 (N_3931,In_2604,In_1419);
nor U3932 (N_3932,In_122,In_623);
and U3933 (N_3933,In_590,In_1353);
or U3934 (N_3934,In_1617,In_70);
or U3935 (N_3935,In_1115,In_1849);
nand U3936 (N_3936,In_170,In_588);
nor U3937 (N_3937,In_2755,In_2391);
and U3938 (N_3938,In_2457,In_2658);
nand U3939 (N_3939,In_1906,In_1518);
and U3940 (N_3940,In_2255,In_2899);
nand U3941 (N_3941,In_39,In_536);
and U3942 (N_3942,In_929,In_55);
nand U3943 (N_3943,In_1922,In_411);
or U3944 (N_3944,In_2069,In_1228);
or U3945 (N_3945,In_2423,In_670);
nand U3946 (N_3946,In_2649,In_2893);
or U3947 (N_3947,In_679,In_2541);
nand U3948 (N_3948,In_2060,In_1748);
nor U3949 (N_3949,In_134,In_1816);
and U3950 (N_3950,In_2187,In_562);
and U3951 (N_3951,In_1365,In_784);
and U3952 (N_3952,In_1057,In_2190);
nor U3953 (N_3953,In_2897,In_1175);
or U3954 (N_3954,In_2729,In_2776);
nor U3955 (N_3955,In_786,In_1538);
xor U3956 (N_3956,In_1621,In_135);
nand U3957 (N_3957,In_2390,In_811);
and U3958 (N_3958,In_2805,In_108);
nor U3959 (N_3959,In_684,In_1874);
nor U3960 (N_3960,In_627,In_1856);
nor U3961 (N_3961,In_2524,In_1249);
nand U3962 (N_3962,In_1785,In_2291);
xor U3963 (N_3963,In_2385,In_2063);
or U3964 (N_3964,In_2794,In_542);
or U3965 (N_3965,In_1175,In_2653);
nand U3966 (N_3966,In_646,In_712);
or U3967 (N_3967,In_1500,In_1027);
or U3968 (N_3968,In_2696,In_76);
or U3969 (N_3969,In_2735,In_1105);
xnor U3970 (N_3970,In_2821,In_2078);
nand U3971 (N_3971,In_343,In_2769);
nor U3972 (N_3972,In_1497,In_1382);
xor U3973 (N_3973,In_461,In_706);
and U3974 (N_3974,In_1215,In_889);
or U3975 (N_3975,In_2393,In_811);
or U3976 (N_3976,In_228,In_578);
and U3977 (N_3977,In_1360,In_1562);
xor U3978 (N_3978,In_2152,In_2607);
nor U3979 (N_3979,In_1847,In_900);
nand U3980 (N_3980,In_528,In_219);
and U3981 (N_3981,In_1705,In_717);
xor U3982 (N_3982,In_1870,In_1077);
nand U3983 (N_3983,In_2277,In_2572);
xnor U3984 (N_3984,In_765,In_2985);
nand U3985 (N_3985,In_1450,In_1731);
or U3986 (N_3986,In_949,In_2734);
nor U3987 (N_3987,In_493,In_970);
nor U3988 (N_3988,In_1134,In_1512);
nand U3989 (N_3989,In_1848,In_1626);
nand U3990 (N_3990,In_54,In_1717);
nand U3991 (N_3991,In_2686,In_1813);
or U3992 (N_3992,In_1071,In_1213);
nand U3993 (N_3993,In_144,In_2228);
xnor U3994 (N_3994,In_1453,In_2673);
and U3995 (N_3995,In_130,In_1240);
and U3996 (N_3996,In_2822,In_1037);
xor U3997 (N_3997,In_1323,In_1613);
or U3998 (N_3998,In_1297,In_578);
or U3999 (N_3999,In_519,In_2782);
xnor U4000 (N_4000,In_2125,In_2717);
nand U4001 (N_4001,In_1708,In_1674);
or U4002 (N_4002,In_2833,In_2243);
xor U4003 (N_4003,In_871,In_465);
nand U4004 (N_4004,In_1855,In_545);
xor U4005 (N_4005,In_1191,In_1684);
xor U4006 (N_4006,In_323,In_2640);
nand U4007 (N_4007,In_2919,In_1604);
or U4008 (N_4008,In_1044,In_2413);
nor U4009 (N_4009,In_1001,In_1239);
nor U4010 (N_4010,In_619,In_2298);
and U4011 (N_4011,In_662,In_1561);
nor U4012 (N_4012,In_593,In_2573);
nand U4013 (N_4013,In_347,In_2894);
and U4014 (N_4014,In_1182,In_1202);
or U4015 (N_4015,In_211,In_1270);
xor U4016 (N_4016,In_2102,In_1193);
nor U4017 (N_4017,In_661,In_2212);
and U4018 (N_4018,In_1580,In_1506);
and U4019 (N_4019,In_1826,In_1205);
or U4020 (N_4020,In_1010,In_1085);
xor U4021 (N_4021,In_1674,In_279);
nand U4022 (N_4022,In_2871,In_2498);
nor U4023 (N_4023,In_2790,In_911);
xor U4024 (N_4024,In_138,In_2375);
nand U4025 (N_4025,In_1573,In_525);
and U4026 (N_4026,In_1718,In_524);
xor U4027 (N_4027,In_2659,In_437);
xnor U4028 (N_4028,In_2418,In_816);
nor U4029 (N_4029,In_384,In_208);
nand U4030 (N_4030,In_1446,In_22);
xnor U4031 (N_4031,In_1705,In_2707);
nor U4032 (N_4032,In_2914,In_874);
xnor U4033 (N_4033,In_1648,In_1546);
and U4034 (N_4034,In_2466,In_2596);
or U4035 (N_4035,In_948,In_2389);
xor U4036 (N_4036,In_2743,In_500);
nand U4037 (N_4037,In_198,In_1516);
and U4038 (N_4038,In_1599,In_2812);
nor U4039 (N_4039,In_1197,In_594);
or U4040 (N_4040,In_1091,In_2512);
or U4041 (N_4041,In_660,In_332);
nand U4042 (N_4042,In_434,In_1505);
or U4043 (N_4043,In_157,In_382);
or U4044 (N_4044,In_1685,In_1263);
xnor U4045 (N_4045,In_300,In_743);
and U4046 (N_4046,In_2870,In_274);
and U4047 (N_4047,In_843,In_2426);
nand U4048 (N_4048,In_2544,In_2752);
nor U4049 (N_4049,In_822,In_329);
nor U4050 (N_4050,In_1292,In_926);
nand U4051 (N_4051,In_986,In_1164);
nor U4052 (N_4052,In_1890,In_2964);
or U4053 (N_4053,In_1509,In_312);
xor U4054 (N_4054,In_1393,In_1233);
or U4055 (N_4055,In_215,In_524);
nand U4056 (N_4056,In_2322,In_1590);
and U4057 (N_4057,In_2293,In_1421);
nand U4058 (N_4058,In_1359,In_1670);
nand U4059 (N_4059,In_1018,In_2679);
nand U4060 (N_4060,In_435,In_83);
nand U4061 (N_4061,In_83,In_1691);
nand U4062 (N_4062,In_1123,In_2563);
nor U4063 (N_4063,In_1450,In_2479);
or U4064 (N_4064,In_1727,In_2451);
nand U4065 (N_4065,In_89,In_2327);
or U4066 (N_4066,In_401,In_1068);
nand U4067 (N_4067,In_2303,In_2601);
or U4068 (N_4068,In_427,In_2160);
and U4069 (N_4069,In_678,In_379);
nor U4070 (N_4070,In_1681,In_2320);
or U4071 (N_4071,In_627,In_2161);
nor U4072 (N_4072,In_1781,In_142);
or U4073 (N_4073,In_2621,In_646);
nor U4074 (N_4074,In_334,In_798);
nand U4075 (N_4075,In_2799,In_1267);
nand U4076 (N_4076,In_2441,In_2596);
or U4077 (N_4077,In_1964,In_2540);
nand U4078 (N_4078,In_1510,In_1065);
nor U4079 (N_4079,In_1230,In_882);
xor U4080 (N_4080,In_336,In_999);
nand U4081 (N_4081,In_582,In_2443);
nor U4082 (N_4082,In_860,In_999);
xor U4083 (N_4083,In_2833,In_282);
and U4084 (N_4084,In_1394,In_1435);
xnor U4085 (N_4085,In_1913,In_556);
xor U4086 (N_4086,In_2234,In_2473);
or U4087 (N_4087,In_1944,In_2171);
and U4088 (N_4088,In_1476,In_30);
or U4089 (N_4089,In_2744,In_2831);
xnor U4090 (N_4090,In_2851,In_1423);
or U4091 (N_4091,In_2351,In_473);
or U4092 (N_4092,In_418,In_276);
and U4093 (N_4093,In_1434,In_2465);
or U4094 (N_4094,In_2523,In_2706);
nand U4095 (N_4095,In_1643,In_1121);
nor U4096 (N_4096,In_214,In_2769);
nand U4097 (N_4097,In_98,In_681);
nand U4098 (N_4098,In_2413,In_1453);
or U4099 (N_4099,In_2184,In_961);
or U4100 (N_4100,In_1414,In_1812);
and U4101 (N_4101,In_1192,In_697);
or U4102 (N_4102,In_1431,In_2550);
nor U4103 (N_4103,In_1912,In_2601);
and U4104 (N_4104,In_799,In_2674);
nand U4105 (N_4105,In_178,In_2316);
or U4106 (N_4106,In_2215,In_1097);
xnor U4107 (N_4107,In_503,In_102);
nand U4108 (N_4108,In_2962,In_1169);
nand U4109 (N_4109,In_1267,In_2036);
or U4110 (N_4110,In_1329,In_1694);
nand U4111 (N_4111,In_2611,In_2975);
or U4112 (N_4112,In_2550,In_870);
and U4113 (N_4113,In_1317,In_2192);
xnor U4114 (N_4114,In_512,In_786);
or U4115 (N_4115,In_2735,In_2793);
xor U4116 (N_4116,In_178,In_2019);
and U4117 (N_4117,In_431,In_1375);
nand U4118 (N_4118,In_1871,In_1252);
and U4119 (N_4119,In_870,In_1636);
and U4120 (N_4120,In_1435,In_370);
or U4121 (N_4121,In_1168,In_917);
xnor U4122 (N_4122,In_1561,In_1948);
nand U4123 (N_4123,In_2725,In_860);
xnor U4124 (N_4124,In_2941,In_357);
nand U4125 (N_4125,In_984,In_1576);
or U4126 (N_4126,In_1241,In_306);
and U4127 (N_4127,In_1930,In_1525);
nand U4128 (N_4128,In_95,In_1738);
and U4129 (N_4129,In_2579,In_137);
and U4130 (N_4130,In_1124,In_2400);
xnor U4131 (N_4131,In_19,In_1644);
or U4132 (N_4132,In_503,In_2970);
nor U4133 (N_4133,In_284,In_2878);
nand U4134 (N_4134,In_2258,In_1752);
or U4135 (N_4135,In_1962,In_943);
and U4136 (N_4136,In_848,In_944);
nor U4137 (N_4137,In_2801,In_1311);
and U4138 (N_4138,In_564,In_498);
or U4139 (N_4139,In_230,In_1670);
xor U4140 (N_4140,In_713,In_939);
nand U4141 (N_4141,In_193,In_2703);
xnor U4142 (N_4142,In_783,In_1237);
and U4143 (N_4143,In_1597,In_2743);
and U4144 (N_4144,In_1582,In_2911);
nor U4145 (N_4145,In_912,In_2751);
or U4146 (N_4146,In_1816,In_2032);
nor U4147 (N_4147,In_1630,In_2859);
nand U4148 (N_4148,In_435,In_1548);
and U4149 (N_4149,In_2746,In_145);
or U4150 (N_4150,In_1308,In_1070);
and U4151 (N_4151,In_2843,In_1045);
xnor U4152 (N_4152,In_790,In_2710);
and U4153 (N_4153,In_1710,In_2251);
xnor U4154 (N_4154,In_2841,In_356);
or U4155 (N_4155,In_1643,In_2167);
nor U4156 (N_4156,In_2455,In_973);
and U4157 (N_4157,In_1382,In_1674);
nor U4158 (N_4158,In_840,In_1029);
or U4159 (N_4159,In_1457,In_937);
xor U4160 (N_4160,In_1308,In_1372);
nor U4161 (N_4161,In_608,In_2665);
or U4162 (N_4162,In_1609,In_2139);
xor U4163 (N_4163,In_1326,In_1945);
nand U4164 (N_4164,In_949,In_1901);
nor U4165 (N_4165,In_2375,In_1103);
xnor U4166 (N_4166,In_2378,In_2248);
nor U4167 (N_4167,In_1062,In_2266);
xor U4168 (N_4168,In_2004,In_2017);
and U4169 (N_4169,In_566,In_2091);
nor U4170 (N_4170,In_1272,In_1924);
nor U4171 (N_4171,In_2320,In_478);
xor U4172 (N_4172,In_1427,In_2500);
or U4173 (N_4173,In_2687,In_616);
nand U4174 (N_4174,In_1829,In_1223);
xor U4175 (N_4175,In_265,In_2421);
nand U4176 (N_4176,In_1942,In_2984);
nor U4177 (N_4177,In_2571,In_2691);
or U4178 (N_4178,In_1588,In_331);
or U4179 (N_4179,In_1016,In_1057);
or U4180 (N_4180,In_610,In_155);
nand U4181 (N_4181,In_813,In_2972);
or U4182 (N_4182,In_2311,In_2167);
or U4183 (N_4183,In_1086,In_1557);
or U4184 (N_4184,In_2806,In_1834);
xor U4185 (N_4185,In_2781,In_1084);
nor U4186 (N_4186,In_1239,In_656);
nand U4187 (N_4187,In_489,In_2037);
nor U4188 (N_4188,In_1206,In_447);
xnor U4189 (N_4189,In_176,In_2262);
xnor U4190 (N_4190,In_671,In_79);
xnor U4191 (N_4191,In_1542,In_1908);
nand U4192 (N_4192,In_1485,In_149);
nand U4193 (N_4193,In_2906,In_1684);
xnor U4194 (N_4194,In_2524,In_1996);
nand U4195 (N_4195,In_1805,In_2591);
xnor U4196 (N_4196,In_1569,In_590);
nand U4197 (N_4197,In_2780,In_1310);
and U4198 (N_4198,In_2238,In_1507);
or U4199 (N_4199,In_951,In_2078);
xor U4200 (N_4200,In_1979,In_1413);
or U4201 (N_4201,In_2373,In_2243);
or U4202 (N_4202,In_2182,In_823);
xnor U4203 (N_4203,In_2309,In_795);
nor U4204 (N_4204,In_8,In_2518);
and U4205 (N_4205,In_2666,In_2099);
nor U4206 (N_4206,In_33,In_100);
xnor U4207 (N_4207,In_449,In_1928);
nor U4208 (N_4208,In_505,In_1666);
xor U4209 (N_4209,In_895,In_925);
or U4210 (N_4210,In_1386,In_644);
nor U4211 (N_4211,In_969,In_2262);
xnor U4212 (N_4212,In_421,In_541);
xor U4213 (N_4213,In_2054,In_1125);
nand U4214 (N_4214,In_2014,In_1528);
and U4215 (N_4215,In_405,In_269);
xor U4216 (N_4216,In_1920,In_1874);
and U4217 (N_4217,In_66,In_2542);
nand U4218 (N_4218,In_2034,In_1919);
and U4219 (N_4219,In_1140,In_1132);
nor U4220 (N_4220,In_1037,In_643);
or U4221 (N_4221,In_1611,In_2459);
xnor U4222 (N_4222,In_145,In_1266);
xor U4223 (N_4223,In_2353,In_360);
xor U4224 (N_4224,In_281,In_1853);
nand U4225 (N_4225,In_2600,In_1529);
xor U4226 (N_4226,In_899,In_931);
nor U4227 (N_4227,In_2768,In_1013);
nand U4228 (N_4228,In_2020,In_2175);
nand U4229 (N_4229,In_31,In_333);
nor U4230 (N_4230,In_2186,In_1481);
xor U4231 (N_4231,In_1679,In_2859);
nor U4232 (N_4232,In_146,In_251);
and U4233 (N_4233,In_518,In_1199);
nor U4234 (N_4234,In_25,In_2911);
or U4235 (N_4235,In_2238,In_1368);
xor U4236 (N_4236,In_277,In_188);
xor U4237 (N_4237,In_1786,In_364);
or U4238 (N_4238,In_2664,In_834);
xor U4239 (N_4239,In_2721,In_2874);
xnor U4240 (N_4240,In_1173,In_2198);
or U4241 (N_4241,In_290,In_434);
or U4242 (N_4242,In_1116,In_234);
and U4243 (N_4243,In_1476,In_163);
or U4244 (N_4244,In_958,In_704);
nand U4245 (N_4245,In_2033,In_1925);
xor U4246 (N_4246,In_1518,In_729);
and U4247 (N_4247,In_615,In_2895);
xnor U4248 (N_4248,In_2644,In_2076);
xnor U4249 (N_4249,In_352,In_2153);
or U4250 (N_4250,In_138,In_1240);
nor U4251 (N_4251,In_2501,In_2409);
or U4252 (N_4252,In_2897,In_2982);
and U4253 (N_4253,In_695,In_847);
nor U4254 (N_4254,In_1558,In_1499);
nand U4255 (N_4255,In_1339,In_2560);
nand U4256 (N_4256,In_637,In_179);
or U4257 (N_4257,In_1,In_898);
and U4258 (N_4258,In_2907,In_2960);
and U4259 (N_4259,In_1228,In_2762);
nand U4260 (N_4260,In_1574,In_2126);
nor U4261 (N_4261,In_549,In_2099);
nor U4262 (N_4262,In_1287,In_862);
nand U4263 (N_4263,In_509,In_342);
or U4264 (N_4264,In_1256,In_245);
nor U4265 (N_4265,In_1968,In_1775);
xor U4266 (N_4266,In_2303,In_2123);
xor U4267 (N_4267,In_2519,In_1023);
nand U4268 (N_4268,In_712,In_1919);
and U4269 (N_4269,In_320,In_2683);
nor U4270 (N_4270,In_1997,In_2512);
or U4271 (N_4271,In_2141,In_1689);
or U4272 (N_4272,In_2953,In_2430);
nand U4273 (N_4273,In_2560,In_1474);
nor U4274 (N_4274,In_1507,In_1613);
nor U4275 (N_4275,In_1410,In_1187);
or U4276 (N_4276,In_2669,In_471);
or U4277 (N_4277,In_383,In_2804);
xnor U4278 (N_4278,In_2110,In_491);
or U4279 (N_4279,In_656,In_2186);
or U4280 (N_4280,In_561,In_2380);
or U4281 (N_4281,In_1472,In_249);
nand U4282 (N_4282,In_1496,In_773);
xnor U4283 (N_4283,In_1232,In_1647);
nand U4284 (N_4284,In_1891,In_38);
nand U4285 (N_4285,In_1499,In_1857);
or U4286 (N_4286,In_2418,In_663);
nand U4287 (N_4287,In_2015,In_1900);
or U4288 (N_4288,In_591,In_558);
nor U4289 (N_4289,In_686,In_719);
and U4290 (N_4290,In_66,In_1433);
nor U4291 (N_4291,In_528,In_1333);
xnor U4292 (N_4292,In_2816,In_1734);
nor U4293 (N_4293,In_572,In_1783);
and U4294 (N_4294,In_1366,In_1780);
nor U4295 (N_4295,In_2483,In_2265);
or U4296 (N_4296,In_2583,In_2909);
nor U4297 (N_4297,In_1305,In_909);
nor U4298 (N_4298,In_2378,In_1882);
nand U4299 (N_4299,In_981,In_1682);
xor U4300 (N_4300,In_1419,In_2196);
and U4301 (N_4301,In_770,In_1041);
or U4302 (N_4302,In_2326,In_1228);
nand U4303 (N_4303,In_2912,In_928);
xor U4304 (N_4304,In_2494,In_1865);
nor U4305 (N_4305,In_1256,In_1573);
nor U4306 (N_4306,In_693,In_1454);
nand U4307 (N_4307,In_714,In_2997);
nor U4308 (N_4308,In_454,In_2526);
xnor U4309 (N_4309,In_274,In_1663);
nor U4310 (N_4310,In_680,In_2435);
nand U4311 (N_4311,In_246,In_334);
nand U4312 (N_4312,In_1389,In_1395);
or U4313 (N_4313,In_431,In_2315);
and U4314 (N_4314,In_2107,In_1086);
or U4315 (N_4315,In_1481,In_1484);
nand U4316 (N_4316,In_2206,In_2596);
and U4317 (N_4317,In_1392,In_155);
or U4318 (N_4318,In_2026,In_1374);
nand U4319 (N_4319,In_1182,In_1724);
and U4320 (N_4320,In_1024,In_2836);
nand U4321 (N_4321,In_1300,In_987);
and U4322 (N_4322,In_574,In_658);
and U4323 (N_4323,In_1451,In_1458);
nand U4324 (N_4324,In_1144,In_1366);
and U4325 (N_4325,In_2635,In_1851);
nand U4326 (N_4326,In_1600,In_1279);
or U4327 (N_4327,In_1598,In_2060);
nand U4328 (N_4328,In_2912,In_1763);
and U4329 (N_4329,In_739,In_1610);
xor U4330 (N_4330,In_412,In_112);
nand U4331 (N_4331,In_530,In_2322);
nor U4332 (N_4332,In_237,In_241);
or U4333 (N_4333,In_1334,In_1041);
nor U4334 (N_4334,In_2127,In_1035);
nor U4335 (N_4335,In_2774,In_1582);
nor U4336 (N_4336,In_1617,In_1374);
nor U4337 (N_4337,In_203,In_1910);
nand U4338 (N_4338,In_2973,In_1408);
nand U4339 (N_4339,In_2247,In_821);
and U4340 (N_4340,In_1667,In_27);
nand U4341 (N_4341,In_2747,In_1583);
nor U4342 (N_4342,In_2803,In_255);
nor U4343 (N_4343,In_1049,In_2186);
xnor U4344 (N_4344,In_551,In_2469);
nor U4345 (N_4345,In_422,In_1509);
and U4346 (N_4346,In_305,In_1555);
xor U4347 (N_4347,In_1682,In_2404);
or U4348 (N_4348,In_2964,In_394);
nor U4349 (N_4349,In_837,In_2775);
and U4350 (N_4350,In_642,In_1319);
or U4351 (N_4351,In_1259,In_2193);
and U4352 (N_4352,In_2548,In_1414);
or U4353 (N_4353,In_1493,In_1690);
nand U4354 (N_4354,In_1862,In_2333);
nor U4355 (N_4355,In_2049,In_1107);
nand U4356 (N_4356,In_1306,In_2845);
nand U4357 (N_4357,In_114,In_1955);
or U4358 (N_4358,In_168,In_1417);
and U4359 (N_4359,In_1272,In_2569);
nand U4360 (N_4360,In_1591,In_703);
nand U4361 (N_4361,In_303,In_1559);
nor U4362 (N_4362,In_2013,In_2198);
nand U4363 (N_4363,In_551,In_1120);
and U4364 (N_4364,In_2890,In_1375);
xnor U4365 (N_4365,In_142,In_1696);
and U4366 (N_4366,In_1660,In_1720);
nand U4367 (N_4367,In_19,In_2261);
xnor U4368 (N_4368,In_2324,In_813);
xnor U4369 (N_4369,In_2104,In_2044);
and U4370 (N_4370,In_1998,In_2189);
or U4371 (N_4371,In_990,In_2764);
nand U4372 (N_4372,In_1638,In_1182);
or U4373 (N_4373,In_2164,In_1403);
or U4374 (N_4374,In_1854,In_765);
and U4375 (N_4375,In_2861,In_1961);
and U4376 (N_4376,In_2326,In_1140);
nand U4377 (N_4377,In_2144,In_2516);
and U4378 (N_4378,In_771,In_290);
and U4379 (N_4379,In_1529,In_1827);
nor U4380 (N_4380,In_967,In_2169);
nor U4381 (N_4381,In_2525,In_525);
nand U4382 (N_4382,In_2595,In_179);
xnor U4383 (N_4383,In_855,In_1594);
or U4384 (N_4384,In_1277,In_2528);
nor U4385 (N_4385,In_33,In_382);
and U4386 (N_4386,In_590,In_9);
or U4387 (N_4387,In_2274,In_1270);
nand U4388 (N_4388,In_2465,In_2408);
nand U4389 (N_4389,In_1515,In_1644);
and U4390 (N_4390,In_1710,In_521);
nand U4391 (N_4391,In_336,In_24);
and U4392 (N_4392,In_1108,In_2511);
nor U4393 (N_4393,In_2155,In_1284);
or U4394 (N_4394,In_760,In_1330);
nand U4395 (N_4395,In_2555,In_1019);
or U4396 (N_4396,In_2769,In_2055);
nand U4397 (N_4397,In_1732,In_2261);
or U4398 (N_4398,In_1211,In_264);
nand U4399 (N_4399,In_1889,In_1411);
nor U4400 (N_4400,In_304,In_267);
nand U4401 (N_4401,In_1081,In_2802);
xor U4402 (N_4402,In_1196,In_2607);
or U4403 (N_4403,In_2224,In_2106);
xnor U4404 (N_4404,In_1000,In_2209);
or U4405 (N_4405,In_1835,In_1035);
xor U4406 (N_4406,In_667,In_1405);
xor U4407 (N_4407,In_1356,In_636);
nand U4408 (N_4408,In_177,In_123);
or U4409 (N_4409,In_2277,In_1890);
xnor U4410 (N_4410,In_1108,In_1272);
or U4411 (N_4411,In_1781,In_1348);
or U4412 (N_4412,In_728,In_639);
nand U4413 (N_4413,In_2298,In_2199);
nand U4414 (N_4414,In_2214,In_1743);
nor U4415 (N_4415,In_838,In_2064);
nand U4416 (N_4416,In_2954,In_111);
xnor U4417 (N_4417,In_2142,In_2557);
nor U4418 (N_4418,In_1061,In_202);
or U4419 (N_4419,In_2872,In_1051);
and U4420 (N_4420,In_134,In_1864);
nor U4421 (N_4421,In_318,In_1564);
xor U4422 (N_4422,In_2184,In_1040);
nand U4423 (N_4423,In_900,In_1010);
or U4424 (N_4424,In_1701,In_261);
or U4425 (N_4425,In_822,In_362);
xor U4426 (N_4426,In_1242,In_2714);
xnor U4427 (N_4427,In_562,In_520);
and U4428 (N_4428,In_2095,In_36);
nor U4429 (N_4429,In_2374,In_263);
nand U4430 (N_4430,In_604,In_2353);
nor U4431 (N_4431,In_2138,In_419);
nand U4432 (N_4432,In_270,In_772);
and U4433 (N_4433,In_1083,In_1545);
nand U4434 (N_4434,In_1779,In_1091);
or U4435 (N_4435,In_410,In_1532);
nand U4436 (N_4436,In_988,In_1559);
or U4437 (N_4437,In_816,In_1537);
and U4438 (N_4438,In_2824,In_661);
xor U4439 (N_4439,In_1194,In_1546);
xnor U4440 (N_4440,In_2649,In_1119);
or U4441 (N_4441,In_498,In_700);
nor U4442 (N_4442,In_430,In_2093);
nor U4443 (N_4443,In_1203,In_2720);
nand U4444 (N_4444,In_2081,In_2885);
xnor U4445 (N_4445,In_2926,In_2740);
nor U4446 (N_4446,In_1123,In_2859);
xnor U4447 (N_4447,In_2270,In_277);
and U4448 (N_4448,In_939,In_1488);
or U4449 (N_4449,In_2915,In_864);
nand U4450 (N_4450,In_42,In_2155);
nand U4451 (N_4451,In_334,In_2544);
nor U4452 (N_4452,In_920,In_1851);
nand U4453 (N_4453,In_242,In_2849);
xor U4454 (N_4454,In_944,In_2196);
xnor U4455 (N_4455,In_2982,In_2299);
xnor U4456 (N_4456,In_652,In_2770);
or U4457 (N_4457,In_117,In_2467);
xor U4458 (N_4458,In_408,In_1575);
and U4459 (N_4459,In_343,In_2141);
xnor U4460 (N_4460,In_2501,In_2019);
or U4461 (N_4461,In_80,In_787);
nand U4462 (N_4462,In_334,In_2409);
xnor U4463 (N_4463,In_1005,In_1657);
nor U4464 (N_4464,In_367,In_1103);
nand U4465 (N_4465,In_1164,In_1409);
xnor U4466 (N_4466,In_2106,In_899);
and U4467 (N_4467,In_2903,In_2781);
or U4468 (N_4468,In_225,In_1795);
xnor U4469 (N_4469,In_1596,In_1500);
and U4470 (N_4470,In_1043,In_462);
or U4471 (N_4471,In_423,In_637);
and U4472 (N_4472,In_1166,In_2358);
xnor U4473 (N_4473,In_1890,In_197);
and U4474 (N_4474,In_2263,In_2455);
and U4475 (N_4475,In_193,In_637);
or U4476 (N_4476,In_1723,In_527);
nand U4477 (N_4477,In_2712,In_3);
nand U4478 (N_4478,In_1173,In_1158);
nor U4479 (N_4479,In_2859,In_2204);
xor U4480 (N_4480,In_227,In_2557);
or U4481 (N_4481,In_1325,In_1646);
and U4482 (N_4482,In_2943,In_2744);
or U4483 (N_4483,In_1238,In_1535);
or U4484 (N_4484,In_2035,In_2457);
and U4485 (N_4485,In_356,In_2814);
xnor U4486 (N_4486,In_621,In_1191);
and U4487 (N_4487,In_1558,In_2588);
nor U4488 (N_4488,In_296,In_1347);
nand U4489 (N_4489,In_1669,In_729);
xor U4490 (N_4490,In_2181,In_714);
nor U4491 (N_4491,In_320,In_2369);
nand U4492 (N_4492,In_1617,In_1795);
nand U4493 (N_4493,In_2959,In_145);
or U4494 (N_4494,In_319,In_2935);
nand U4495 (N_4495,In_2063,In_2879);
and U4496 (N_4496,In_1835,In_1691);
nand U4497 (N_4497,In_2158,In_2062);
or U4498 (N_4498,In_1091,In_1314);
xor U4499 (N_4499,In_2665,In_1729);
or U4500 (N_4500,In_87,In_961);
nand U4501 (N_4501,In_2210,In_546);
or U4502 (N_4502,In_257,In_93);
or U4503 (N_4503,In_857,In_2766);
xnor U4504 (N_4504,In_1481,In_1674);
or U4505 (N_4505,In_275,In_2653);
nor U4506 (N_4506,In_867,In_2835);
or U4507 (N_4507,In_1595,In_212);
and U4508 (N_4508,In_1683,In_1802);
xnor U4509 (N_4509,In_2911,In_296);
nor U4510 (N_4510,In_2677,In_1477);
nor U4511 (N_4511,In_2102,In_2240);
or U4512 (N_4512,In_508,In_2176);
or U4513 (N_4513,In_377,In_1323);
or U4514 (N_4514,In_2902,In_1418);
nand U4515 (N_4515,In_1704,In_1409);
or U4516 (N_4516,In_2994,In_220);
nand U4517 (N_4517,In_2711,In_580);
and U4518 (N_4518,In_2373,In_1306);
xor U4519 (N_4519,In_2134,In_1449);
nor U4520 (N_4520,In_2,In_1357);
and U4521 (N_4521,In_2223,In_1688);
xor U4522 (N_4522,In_1244,In_1550);
xor U4523 (N_4523,In_346,In_1418);
xnor U4524 (N_4524,In_2973,In_905);
and U4525 (N_4525,In_2871,In_289);
nor U4526 (N_4526,In_675,In_130);
xor U4527 (N_4527,In_2615,In_1969);
or U4528 (N_4528,In_2762,In_742);
and U4529 (N_4529,In_1088,In_1555);
nor U4530 (N_4530,In_2449,In_1735);
nand U4531 (N_4531,In_780,In_1368);
and U4532 (N_4532,In_1665,In_794);
xnor U4533 (N_4533,In_2832,In_2450);
xnor U4534 (N_4534,In_2431,In_2344);
nor U4535 (N_4535,In_225,In_2380);
nand U4536 (N_4536,In_1183,In_755);
nand U4537 (N_4537,In_1824,In_1947);
or U4538 (N_4538,In_1074,In_2872);
nand U4539 (N_4539,In_1109,In_139);
or U4540 (N_4540,In_2950,In_850);
or U4541 (N_4541,In_1657,In_1958);
or U4542 (N_4542,In_2761,In_283);
nand U4543 (N_4543,In_2886,In_984);
or U4544 (N_4544,In_2949,In_518);
or U4545 (N_4545,In_589,In_1854);
nor U4546 (N_4546,In_852,In_2716);
nor U4547 (N_4547,In_1236,In_674);
nand U4548 (N_4548,In_2330,In_2393);
or U4549 (N_4549,In_2361,In_1258);
nand U4550 (N_4550,In_121,In_2482);
nand U4551 (N_4551,In_1641,In_272);
nor U4552 (N_4552,In_294,In_1861);
nand U4553 (N_4553,In_959,In_2475);
nor U4554 (N_4554,In_2885,In_2641);
nand U4555 (N_4555,In_811,In_2724);
nor U4556 (N_4556,In_829,In_1391);
nor U4557 (N_4557,In_611,In_1246);
nand U4558 (N_4558,In_753,In_1258);
or U4559 (N_4559,In_54,In_1430);
nor U4560 (N_4560,In_1117,In_127);
and U4561 (N_4561,In_2243,In_2220);
nand U4562 (N_4562,In_1708,In_2558);
and U4563 (N_4563,In_505,In_676);
xor U4564 (N_4564,In_2532,In_432);
and U4565 (N_4565,In_508,In_2650);
nand U4566 (N_4566,In_534,In_1682);
and U4567 (N_4567,In_2181,In_1243);
and U4568 (N_4568,In_2382,In_2557);
xor U4569 (N_4569,In_1867,In_2092);
nand U4570 (N_4570,In_2355,In_233);
or U4571 (N_4571,In_2090,In_1014);
or U4572 (N_4572,In_1148,In_2501);
and U4573 (N_4573,In_2289,In_2413);
xnor U4574 (N_4574,In_2183,In_76);
xnor U4575 (N_4575,In_1836,In_1084);
xnor U4576 (N_4576,In_2607,In_1538);
or U4577 (N_4577,In_2246,In_1212);
or U4578 (N_4578,In_851,In_558);
and U4579 (N_4579,In_136,In_2212);
nand U4580 (N_4580,In_612,In_2105);
nor U4581 (N_4581,In_2498,In_702);
nand U4582 (N_4582,In_73,In_256);
or U4583 (N_4583,In_2640,In_2769);
nand U4584 (N_4584,In_1304,In_949);
nor U4585 (N_4585,In_2417,In_2227);
nand U4586 (N_4586,In_2113,In_1657);
nor U4587 (N_4587,In_2150,In_2800);
nor U4588 (N_4588,In_540,In_2901);
and U4589 (N_4589,In_566,In_1553);
nand U4590 (N_4590,In_345,In_2041);
xnor U4591 (N_4591,In_2142,In_468);
and U4592 (N_4592,In_457,In_487);
or U4593 (N_4593,In_980,In_1048);
nand U4594 (N_4594,In_2305,In_1170);
nor U4595 (N_4595,In_718,In_2560);
and U4596 (N_4596,In_1190,In_481);
or U4597 (N_4597,In_827,In_2773);
and U4598 (N_4598,In_1640,In_1895);
xnor U4599 (N_4599,In_514,In_1963);
or U4600 (N_4600,In_1395,In_2146);
and U4601 (N_4601,In_188,In_2283);
xnor U4602 (N_4602,In_428,In_628);
xor U4603 (N_4603,In_52,In_2433);
and U4604 (N_4604,In_1138,In_2860);
nand U4605 (N_4605,In_246,In_1243);
nand U4606 (N_4606,In_279,In_2348);
nor U4607 (N_4607,In_1872,In_1410);
nand U4608 (N_4608,In_2953,In_994);
and U4609 (N_4609,In_847,In_253);
or U4610 (N_4610,In_580,In_565);
or U4611 (N_4611,In_2961,In_867);
nor U4612 (N_4612,In_2081,In_716);
xor U4613 (N_4613,In_1303,In_642);
nand U4614 (N_4614,In_389,In_2148);
nand U4615 (N_4615,In_1537,In_2085);
or U4616 (N_4616,In_2811,In_969);
nor U4617 (N_4617,In_2464,In_788);
and U4618 (N_4618,In_1843,In_1484);
nand U4619 (N_4619,In_434,In_1541);
nor U4620 (N_4620,In_2460,In_2297);
nand U4621 (N_4621,In_2318,In_13);
and U4622 (N_4622,In_1754,In_2767);
nand U4623 (N_4623,In_1600,In_2008);
xnor U4624 (N_4624,In_2689,In_2149);
nor U4625 (N_4625,In_2932,In_2935);
xor U4626 (N_4626,In_624,In_2689);
nor U4627 (N_4627,In_144,In_872);
nand U4628 (N_4628,In_228,In_1201);
nand U4629 (N_4629,In_57,In_2421);
and U4630 (N_4630,In_1176,In_1906);
and U4631 (N_4631,In_195,In_1815);
nand U4632 (N_4632,In_2878,In_148);
nor U4633 (N_4633,In_303,In_2008);
nor U4634 (N_4634,In_1420,In_1668);
and U4635 (N_4635,In_2456,In_2403);
and U4636 (N_4636,In_1224,In_2717);
and U4637 (N_4637,In_1908,In_183);
nor U4638 (N_4638,In_2285,In_879);
nand U4639 (N_4639,In_1648,In_2311);
or U4640 (N_4640,In_2740,In_903);
xnor U4641 (N_4641,In_1415,In_408);
and U4642 (N_4642,In_1272,In_773);
xor U4643 (N_4643,In_2014,In_2980);
nand U4644 (N_4644,In_2078,In_2067);
nand U4645 (N_4645,In_839,In_1691);
nand U4646 (N_4646,In_1820,In_1634);
and U4647 (N_4647,In_2382,In_1491);
xor U4648 (N_4648,In_2403,In_1130);
xor U4649 (N_4649,In_272,In_630);
nand U4650 (N_4650,In_2703,In_2477);
nand U4651 (N_4651,In_437,In_648);
nand U4652 (N_4652,In_1179,In_2505);
nor U4653 (N_4653,In_1829,In_1868);
xnor U4654 (N_4654,In_1943,In_1356);
nor U4655 (N_4655,In_2985,In_2502);
nand U4656 (N_4656,In_2081,In_2658);
and U4657 (N_4657,In_2965,In_2770);
nand U4658 (N_4658,In_91,In_2720);
nor U4659 (N_4659,In_1665,In_80);
and U4660 (N_4660,In_2232,In_2322);
and U4661 (N_4661,In_817,In_1237);
and U4662 (N_4662,In_2677,In_1730);
nand U4663 (N_4663,In_1679,In_326);
xor U4664 (N_4664,In_2952,In_226);
nand U4665 (N_4665,In_2900,In_1287);
xnor U4666 (N_4666,In_354,In_1539);
or U4667 (N_4667,In_2188,In_1714);
and U4668 (N_4668,In_237,In_2153);
nand U4669 (N_4669,In_165,In_2966);
xor U4670 (N_4670,In_2682,In_2629);
or U4671 (N_4671,In_1106,In_257);
nand U4672 (N_4672,In_1544,In_2056);
and U4673 (N_4673,In_2471,In_2934);
and U4674 (N_4674,In_766,In_870);
and U4675 (N_4675,In_1174,In_2674);
nand U4676 (N_4676,In_2160,In_27);
and U4677 (N_4677,In_1211,In_825);
and U4678 (N_4678,In_788,In_455);
nand U4679 (N_4679,In_79,In_2266);
nor U4680 (N_4680,In_105,In_1768);
xnor U4681 (N_4681,In_150,In_2139);
or U4682 (N_4682,In_1793,In_2701);
nor U4683 (N_4683,In_1024,In_2239);
nand U4684 (N_4684,In_2534,In_2424);
nand U4685 (N_4685,In_888,In_2527);
nor U4686 (N_4686,In_187,In_2635);
xor U4687 (N_4687,In_2012,In_364);
or U4688 (N_4688,In_2673,In_1103);
nand U4689 (N_4689,In_664,In_1721);
and U4690 (N_4690,In_2965,In_2766);
xor U4691 (N_4691,In_1558,In_2863);
and U4692 (N_4692,In_2429,In_2896);
or U4693 (N_4693,In_2057,In_2556);
nor U4694 (N_4694,In_2621,In_663);
or U4695 (N_4695,In_1902,In_2680);
xor U4696 (N_4696,In_1826,In_1820);
nand U4697 (N_4697,In_2513,In_2559);
xnor U4698 (N_4698,In_2176,In_1895);
nor U4699 (N_4699,In_2023,In_189);
nand U4700 (N_4700,In_2111,In_2838);
xor U4701 (N_4701,In_1529,In_425);
and U4702 (N_4702,In_1402,In_2007);
nor U4703 (N_4703,In_2625,In_1802);
xor U4704 (N_4704,In_217,In_785);
or U4705 (N_4705,In_1301,In_2528);
and U4706 (N_4706,In_1204,In_280);
nor U4707 (N_4707,In_2381,In_2071);
and U4708 (N_4708,In_2580,In_2535);
nor U4709 (N_4709,In_176,In_596);
nand U4710 (N_4710,In_2475,In_2739);
xnor U4711 (N_4711,In_356,In_2561);
nand U4712 (N_4712,In_501,In_1792);
and U4713 (N_4713,In_274,In_100);
nor U4714 (N_4714,In_2703,In_848);
xnor U4715 (N_4715,In_1075,In_897);
nor U4716 (N_4716,In_1937,In_194);
and U4717 (N_4717,In_1005,In_2639);
and U4718 (N_4718,In_1375,In_536);
nand U4719 (N_4719,In_2519,In_2557);
nand U4720 (N_4720,In_768,In_1854);
and U4721 (N_4721,In_1736,In_335);
and U4722 (N_4722,In_834,In_820);
nor U4723 (N_4723,In_1916,In_1922);
xnor U4724 (N_4724,In_2982,In_1634);
xor U4725 (N_4725,In_413,In_520);
nor U4726 (N_4726,In_1002,In_681);
or U4727 (N_4727,In_673,In_629);
nand U4728 (N_4728,In_661,In_323);
or U4729 (N_4729,In_184,In_2831);
or U4730 (N_4730,In_1620,In_28);
nor U4731 (N_4731,In_2958,In_259);
xor U4732 (N_4732,In_1079,In_949);
or U4733 (N_4733,In_888,In_1854);
and U4734 (N_4734,In_1559,In_399);
or U4735 (N_4735,In_367,In_170);
or U4736 (N_4736,In_1963,In_2806);
or U4737 (N_4737,In_2587,In_1473);
and U4738 (N_4738,In_1938,In_1081);
nor U4739 (N_4739,In_1011,In_1198);
and U4740 (N_4740,In_2288,In_2076);
and U4741 (N_4741,In_2844,In_2747);
xor U4742 (N_4742,In_1355,In_2855);
xor U4743 (N_4743,In_2263,In_2010);
nand U4744 (N_4744,In_508,In_449);
nor U4745 (N_4745,In_2684,In_1749);
xnor U4746 (N_4746,In_1303,In_657);
nand U4747 (N_4747,In_457,In_674);
nor U4748 (N_4748,In_1112,In_2421);
xnor U4749 (N_4749,In_2527,In_1587);
nor U4750 (N_4750,In_2,In_147);
nand U4751 (N_4751,In_2774,In_1366);
or U4752 (N_4752,In_548,In_844);
or U4753 (N_4753,In_2456,In_2777);
and U4754 (N_4754,In_887,In_1104);
xor U4755 (N_4755,In_1901,In_1801);
nand U4756 (N_4756,In_331,In_1631);
and U4757 (N_4757,In_1526,In_1904);
nor U4758 (N_4758,In_173,In_2173);
and U4759 (N_4759,In_2389,In_189);
nand U4760 (N_4760,In_535,In_658);
nor U4761 (N_4761,In_1183,In_2168);
or U4762 (N_4762,In_1447,In_2429);
and U4763 (N_4763,In_322,In_2535);
or U4764 (N_4764,In_2833,In_964);
or U4765 (N_4765,In_1214,In_633);
nand U4766 (N_4766,In_2536,In_2408);
and U4767 (N_4767,In_89,In_997);
and U4768 (N_4768,In_2833,In_2134);
and U4769 (N_4769,In_862,In_2086);
or U4770 (N_4770,In_769,In_1166);
nor U4771 (N_4771,In_1796,In_98);
nor U4772 (N_4772,In_1013,In_137);
xor U4773 (N_4773,In_1382,In_1627);
nand U4774 (N_4774,In_698,In_904);
nand U4775 (N_4775,In_1381,In_142);
and U4776 (N_4776,In_2373,In_189);
nor U4777 (N_4777,In_437,In_1259);
and U4778 (N_4778,In_1290,In_1234);
nand U4779 (N_4779,In_1272,In_2635);
nor U4780 (N_4780,In_440,In_2647);
nand U4781 (N_4781,In_25,In_172);
xnor U4782 (N_4782,In_589,In_114);
nor U4783 (N_4783,In_984,In_1903);
nor U4784 (N_4784,In_2479,In_1086);
nor U4785 (N_4785,In_2387,In_2051);
or U4786 (N_4786,In_2894,In_889);
and U4787 (N_4787,In_1770,In_872);
nor U4788 (N_4788,In_2022,In_1230);
xnor U4789 (N_4789,In_1346,In_2278);
or U4790 (N_4790,In_1622,In_444);
nor U4791 (N_4791,In_2431,In_1819);
xnor U4792 (N_4792,In_895,In_2186);
and U4793 (N_4793,In_1243,In_1914);
or U4794 (N_4794,In_1168,In_1536);
or U4795 (N_4795,In_2029,In_2537);
xnor U4796 (N_4796,In_2730,In_288);
nor U4797 (N_4797,In_1557,In_464);
xnor U4798 (N_4798,In_1687,In_2812);
or U4799 (N_4799,In_2306,In_2000);
nor U4800 (N_4800,In_384,In_648);
nor U4801 (N_4801,In_2038,In_2354);
and U4802 (N_4802,In_2451,In_1902);
xor U4803 (N_4803,In_2598,In_1953);
and U4804 (N_4804,In_1557,In_2662);
nor U4805 (N_4805,In_1790,In_2282);
and U4806 (N_4806,In_371,In_497);
nand U4807 (N_4807,In_1990,In_837);
and U4808 (N_4808,In_2660,In_2819);
nand U4809 (N_4809,In_986,In_1858);
or U4810 (N_4810,In_2237,In_2102);
or U4811 (N_4811,In_2055,In_628);
xor U4812 (N_4812,In_951,In_157);
nand U4813 (N_4813,In_670,In_1103);
and U4814 (N_4814,In_1071,In_2307);
or U4815 (N_4815,In_1879,In_1856);
xnor U4816 (N_4816,In_271,In_480);
or U4817 (N_4817,In_2484,In_2837);
nor U4818 (N_4818,In_902,In_2363);
nand U4819 (N_4819,In_132,In_695);
or U4820 (N_4820,In_260,In_134);
nand U4821 (N_4821,In_2422,In_713);
or U4822 (N_4822,In_2030,In_2298);
and U4823 (N_4823,In_2187,In_970);
or U4824 (N_4824,In_1826,In_1586);
nor U4825 (N_4825,In_365,In_2363);
nand U4826 (N_4826,In_1748,In_2445);
nand U4827 (N_4827,In_381,In_393);
xnor U4828 (N_4828,In_2089,In_1215);
nand U4829 (N_4829,In_1301,In_1610);
and U4830 (N_4830,In_286,In_418);
or U4831 (N_4831,In_2746,In_2153);
nand U4832 (N_4832,In_1511,In_1737);
xnor U4833 (N_4833,In_910,In_833);
nand U4834 (N_4834,In_1222,In_2900);
and U4835 (N_4835,In_2124,In_588);
nor U4836 (N_4836,In_238,In_1196);
nor U4837 (N_4837,In_334,In_2564);
nor U4838 (N_4838,In_1201,In_1782);
xor U4839 (N_4839,In_220,In_839);
nor U4840 (N_4840,In_1753,In_13);
nand U4841 (N_4841,In_2351,In_2486);
xnor U4842 (N_4842,In_108,In_2745);
nor U4843 (N_4843,In_977,In_1366);
and U4844 (N_4844,In_2195,In_2898);
nand U4845 (N_4845,In_2136,In_1540);
nor U4846 (N_4846,In_304,In_2105);
nor U4847 (N_4847,In_1039,In_2890);
and U4848 (N_4848,In_1328,In_2905);
and U4849 (N_4849,In_2353,In_2289);
nor U4850 (N_4850,In_748,In_953);
or U4851 (N_4851,In_2328,In_1054);
nand U4852 (N_4852,In_2909,In_260);
or U4853 (N_4853,In_253,In_2816);
or U4854 (N_4854,In_526,In_407);
or U4855 (N_4855,In_2025,In_950);
nor U4856 (N_4856,In_2969,In_2856);
or U4857 (N_4857,In_2000,In_244);
nor U4858 (N_4858,In_1936,In_2849);
nor U4859 (N_4859,In_194,In_732);
nor U4860 (N_4860,In_2058,In_1058);
and U4861 (N_4861,In_191,In_756);
and U4862 (N_4862,In_2234,In_1435);
nand U4863 (N_4863,In_2816,In_2923);
xor U4864 (N_4864,In_2032,In_1892);
and U4865 (N_4865,In_1810,In_433);
or U4866 (N_4866,In_699,In_2039);
or U4867 (N_4867,In_1368,In_1407);
and U4868 (N_4868,In_941,In_1884);
xor U4869 (N_4869,In_1548,In_1857);
or U4870 (N_4870,In_2691,In_133);
nand U4871 (N_4871,In_868,In_74);
nor U4872 (N_4872,In_1114,In_2083);
or U4873 (N_4873,In_904,In_636);
and U4874 (N_4874,In_2183,In_1954);
xor U4875 (N_4875,In_1445,In_2843);
or U4876 (N_4876,In_131,In_241);
nand U4877 (N_4877,In_2490,In_1194);
nand U4878 (N_4878,In_1108,In_254);
or U4879 (N_4879,In_481,In_1801);
xor U4880 (N_4880,In_1484,In_2835);
nand U4881 (N_4881,In_2881,In_528);
nor U4882 (N_4882,In_1199,In_1157);
or U4883 (N_4883,In_1600,In_2235);
and U4884 (N_4884,In_1132,In_923);
and U4885 (N_4885,In_2372,In_1307);
or U4886 (N_4886,In_2978,In_95);
xor U4887 (N_4887,In_1375,In_1045);
nor U4888 (N_4888,In_1361,In_1653);
nand U4889 (N_4889,In_2837,In_410);
or U4890 (N_4890,In_863,In_2441);
and U4891 (N_4891,In_1368,In_2885);
nand U4892 (N_4892,In_1287,In_1952);
xnor U4893 (N_4893,In_378,In_1839);
nand U4894 (N_4894,In_1537,In_1491);
nand U4895 (N_4895,In_662,In_281);
nand U4896 (N_4896,In_2619,In_2604);
nor U4897 (N_4897,In_358,In_2040);
and U4898 (N_4898,In_996,In_628);
nor U4899 (N_4899,In_1491,In_904);
and U4900 (N_4900,In_2893,In_2571);
nor U4901 (N_4901,In_1506,In_468);
nand U4902 (N_4902,In_638,In_2676);
xor U4903 (N_4903,In_2462,In_1903);
nor U4904 (N_4904,In_860,In_2219);
and U4905 (N_4905,In_2048,In_206);
and U4906 (N_4906,In_1098,In_2891);
xor U4907 (N_4907,In_625,In_1599);
and U4908 (N_4908,In_892,In_2729);
xnor U4909 (N_4909,In_2862,In_2849);
and U4910 (N_4910,In_710,In_2899);
and U4911 (N_4911,In_783,In_2588);
xor U4912 (N_4912,In_2123,In_2540);
xor U4913 (N_4913,In_1688,In_2249);
or U4914 (N_4914,In_1017,In_2698);
or U4915 (N_4915,In_2963,In_2876);
and U4916 (N_4916,In_1114,In_2517);
nor U4917 (N_4917,In_1913,In_968);
nand U4918 (N_4918,In_944,In_2023);
and U4919 (N_4919,In_2185,In_313);
or U4920 (N_4920,In_422,In_2527);
xor U4921 (N_4921,In_1588,In_513);
and U4922 (N_4922,In_2573,In_735);
nand U4923 (N_4923,In_2679,In_458);
or U4924 (N_4924,In_1726,In_2521);
and U4925 (N_4925,In_1068,In_2001);
nor U4926 (N_4926,In_275,In_1016);
nor U4927 (N_4927,In_763,In_94);
nand U4928 (N_4928,In_900,In_1060);
nand U4929 (N_4929,In_1756,In_1894);
xnor U4930 (N_4930,In_1035,In_1163);
nor U4931 (N_4931,In_1375,In_388);
or U4932 (N_4932,In_2768,In_227);
or U4933 (N_4933,In_2770,In_1172);
xor U4934 (N_4934,In_1539,In_2291);
or U4935 (N_4935,In_629,In_1132);
xor U4936 (N_4936,In_2238,In_2184);
nor U4937 (N_4937,In_121,In_514);
nand U4938 (N_4938,In_257,In_1478);
nor U4939 (N_4939,In_2170,In_146);
and U4940 (N_4940,In_1136,In_669);
and U4941 (N_4941,In_2325,In_2897);
xor U4942 (N_4942,In_2004,In_415);
nor U4943 (N_4943,In_2517,In_1825);
nand U4944 (N_4944,In_718,In_2896);
xor U4945 (N_4945,In_39,In_2161);
xnor U4946 (N_4946,In_289,In_506);
nand U4947 (N_4947,In_543,In_1258);
and U4948 (N_4948,In_307,In_2203);
nor U4949 (N_4949,In_2489,In_2933);
or U4950 (N_4950,In_1361,In_1937);
and U4951 (N_4951,In_339,In_2111);
nor U4952 (N_4952,In_967,In_380);
nor U4953 (N_4953,In_1227,In_2971);
and U4954 (N_4954,In_816,In_2336);
or U4955 (N_4955,In_305,In_2866);
or U4956 (N_4956,In_1554,In_1054);
or U4957 (N_4957,In_1413,In_931);
and U4958 (N_4958,In_1574,In_394);
or U4959 (N_4959,In_1803,In_2610);
nand U4960 (N_4960,In_409,In_660);
nor U4961 (N_4961,In_875,In_2938);
and U4962 (N_4962,In_2534,In_2433);
nor U4963 (N_4963,In_1014,In_409);
nand U4964 (N_4964,In_1667,In_1807);
nand U4965 (N_4965,In_681,In_689);
or U4966 (N_4966,In_2053,In_1374);
xor U4967 (N_4967,In_2134,In_2682);
or U4968 (N_4968,In_818,In_98);
xnor U4969 (N_4969,In_1534,In_1461);
or U4970 (N_4970,In_861,In_1695);
nand U4971 (N_4971,In_2696,In_1472);
nand U4972 (N_4972,In_2960,In_2082);
xor U4973 (N_4973,In_1346,In_1603);
or U4974 (N_4974,In_1059,In_1185);
and U4975 (N_4975,In_1484,In_775);
nand U4976 (N_4976,In_1879,In_2849);
or U4977 (N_4977,In_83,In_1000);
and U4978 (N_4978,In_843,In_2181);
nand U4979 (N_4979,In_1227,In_2408);
and U4980 (N_4980,In_1221,In_683);
nor U4981 (N_4981,In_483,In_2048);
nor U4982 (N_4982,In_939,In_2298);
nand U4983 (N_4983,In_774,In_1468);
and U4984 (N_4984,In_73,In_328);
xnor U4985 (N_4985,In_798,In_554);
or U4986 (N_4986,In_2009,In_2279);
nor U4987 (N_4987,In_543,In_555);
xnor U4988 (N_4988,In_764,In_940);
or U4989 (N_4989,In_1214,In_1341);
nand U4990 (N_4990,In_415,In_2955);
xnor U4991 (N_4991,In_396,In_48);
and U4992 (N_4992,In_2898,In_1592);
and U4993 (N_4993,In_431,In_2746);
and U4994 (N_4994,In_886,In_2491);
and U4995 (N_4995,In_372,In_141);
nor U4996 (N_4996,In_2517,In_831);
xnor U4997 (N_4997,In_2300,In_2852);
nor U4998 (N_4998,In_1639,In_772);
or U4999 (N_4999,In_144,In_361);
and U5000 (N_5000,In_1143,In_2892);
or U5001 (N_5001,In_765,In_2057);
nor U5002 (N_5002,In_226,In_1967);
nand U5003 (N_5003,In_2824,In_2639);
or U5004 (N_5004,In_2820,In_2238);
nor U5005 (N_5005,In_621,In_934);
nor U5006 (N_5006,In_374,In_1267);
nor U5007 (N_5007,In_2150,In_2786);
and U5008 (N_5008,In_1846,In_2769);
or U5009 (N_5009,In_2909,In_2932);
xnor U5010 (N_5010,In_2489,In_897);
nand U5011 (N_5011,In_781,In_1094);
nand U5012 (N_5012,In_110,In_71);
nor U5013 (N_5013,In_1722,In_1884);
nor U5014 (N_5014,In_425,In_2610);
nor U5015 (N_5015,In_2963,In_1876);
nand U5016 (N_5016,In_2234,In_1675);
nor U5017 (N_5017,In_938,In_2519);
nor U5018 (N_5018,In_2117,In_330);
and U5019 (N_5019,In_1124,In_2990);
nand U5020 (N_5020,In_299,In_377);
or U5021 (N_5021,In_1671,In_1326);
nand U5022 (N_5022,In_2988,In_770);
xor U5023 (N_5023,In_692,In_2067);
nor U5024 (N_5024,In_2720,In_687);
nor U5025 (N_5025,In_2081,In_2787);
or U5026 (N_5026,In_809,In_1115);
and U5027 (N_5027,In_2169,In_2004);
xor U5028 (N_5028,In_2208,In_159);
or U5029 (N_5029,In_984,In_431);
nand U5030 (N_5030,In_1966,In_1046);
or U5031 (N_5031,In_2273,In_558);
xor U5032 (N_5032,In_888,In_1847);
xnor U5033 (N_5033,In_2475,In_484);
nand U5034 (N_5034,In_146,In_1094);
nand U5035 (N_5035,In_423,In_278);
xor U5036 (N_5036,In_1443,In_2751);
nor U5037 (N_5037,In_1627,In_1208);
and U5038 (N_5038,In_2334,In_584);
and U5039 (N_5039,In_2899,In_859);
nand U5040 (N_5040,In_2824,In_43);
nand U5041 (N_5041,In_1877,In_1505);
or U5042 (N_5042,In_1199,In_2457);
xor U5043 (N_5043,In_396,In_163);
or U5044 (N_5044,In_499,In_2669);
nor U5045 (N_5045,In_2984,In_414);
xnor U5046 (N_5046,In_1722,In_2386);
and U5047 (N_5047,In_2879,In_569);
or U5048 (N_5048,In_908,In_2988);
nor U5049 (N_5049,In_144,In_2638);
or U5050 (N_5050,In_872,In_2067);
nor U5051 (N_5051,In_146,In_9);
or U5052 (N_5052,In_2808,In_854);
nor U5053 (N_5053,In_990,In_906);
nand U5054 (N_5054,In_2872,In_196);
and U5055 (N_5055,In_1100,In_772);
nor U5056 (N_5056,In_631,In_2178);
or U5057 (N_5057,In_1968,In_2325);
or U5058 (N_5058,In_2574,In_2170);
xor U5059 (N_5059,In_1703,In_2322);
nor U5060 (N_5060,In_1173,In_1470);
nand U5061 (N_5061,In_2225,In_2308);
nor U5062 (N_5062,In_1148,In_1433);
and U5063 (N_5063,In_1170,In_197);
xor U5064 (N_5064,In_1350,In_390);
xnor U5065 (N_5065,In_1619,In_2230);
nor U5066 (N_5066,In_1471,In_1802);
or U5067 (N_5067,In_2429,In_1948);
xnor U5068 (N_5068,In_2471,In_904);
xnor U5069 (N_5069,In_14,In_1893);
xor U5070 (N_5070,In_2274,In_681);
or U5071 (N_5071,In_2669,In_2792);
nor U5072 (N_5072,In_2358,In_828);
nor U5073 (N_5073,In_1582,In_2951);
xnor U5074 (N_5074,In_2833,In_2513);
or U5075 (N_5075,In_83,In_1479);
nor U5076 (N_5076,In_527,In_2074);
nand U5077 (N_5077,In_2429,In_582);
nand U5078 (N_5078,In_2293,In_1019);
and U5079 (N_5079,In_1792,In_2005);
and U5080 (N_5080,In_2022,In_234);
xnor U5081 (N_5081,In_1973,In_1220);
and U5082 (N_5082,In_162,In_335);
xor U5083 (N_5083,In_251,In_651);
nor U5084 (N_5084,In_2329,In_814);
xnor U5085 (N_5085,In_2189,In_1123);
and U5086 (N_5086,In_1069,In_2067);
or U5087 (N_5087,In_2505,In_1721);
xnor U5088 (N_5088,In_2434,In_1327);
xor U5089 (N_5089,In_292,In_221);
and U5090 (N_5090,In_2298,In_2623);
nand U5091 (N_5091,In_1041,In_1108);
xnor U5092 (N_5092,In_1662,In_1311);
xor U5093 (N_5093,In_618,In_2822);
and U5094 (N_5094,In_1105,In_1539);
or U5095 (N_5095,In_871,In_0);
nand U5096 (N_5096,In_609,In_387);
or U5097 (N_5097,In_583,In_1950);
xnor U5098 (N_5098,In_1020,In_615);
nor U5099 (N_5099,In_215,In_2550);
xor U5100 (N_5100,In_1033,In_2296);
nand U5101 (N_5101,In_1852,In_1949);
xnor U5102 (N_5102,In_2907,In_811);
nand U5103 (N_5103,In_1924,In_807);
nand U5104 (N_5104,In_1280,In_1937);
and U5105 (N_5105,In_1409,In_1517);
nand U5106 (N_5106,In_2628,In_779);
or U5107 (N_5107,In_1140,In_1880);
and U5108 (N_5108,In_2253,In_2842);
nand U5109 (N_5109,In_1317,In_264);
and U5110 (N_5110,In_2193,In_2867);
and U5111 (N_5111,In_1090,In_2913);
and U5112 (N_5112,In_999,In_1224);
and U5113 (N_5113,In_181,In_1798);
nor U5114 (N_5114,In_2308,In_455);
and U5115 (N_5115,In_2088,In_650);
and U5116 (N_5116,In_2863,In_2850);
nor U5117 (N_5117,In_1193,In_16);
and U5118 (N_5118,In_1183,In_1132);
nand U5119 (N_5119,In_1294,In_1474);
or U5120 (N_5120,In_1178,In_364);
or U5121 (N_5121,In_417,In_1994);
xnor U5122 (N_5122,In_564,In_742);
nand U5123 (N_5123,In_665,In_1079);
or U5124 (N_5124,In_1517,In_2941);
xor U5125 (N_5125,In_1052,In_546);
and U5126 (N_5126,In_2623,In_229);
or U5127 (N_5127,In_2997,In_106);
nand U5128 (N_5128,In_1201,In_1440);
or U5129 (N_5129,In_2062,In_2501);
or U5130 (N_5130,In_2315,In_2679);
xnor U5131 (N_5131,In_553,In_338);
nor U5132 (N_5132,In_2974,In_604);
or U5133 (N_5133,In_1780,In_1504);
or U5134 (N_5134,In_2418,In_1948);
nand U5135 (N_5135,In_1214,In_1508);
and U5136 (N_5136,In_2572,In_1064);
nand U5137 (N_5137,In_2668,In_2856);
nor U5138 (N_5138,In_2826,In_1025);
xnor U5139 (N_5139,In_427,In_1771);
and U5140 (N_5140,In_2411,In_2035);
nand U5141 (N_5141,In_2991,In_674);
xor U5142 (N_5142,In_1313,In_4);
nor U5143 (N_5143,In_810,In_926);
or U5144 (N_5144,In_1606,In_336);
or U5145 (N_5145,In_527,In_2554);
nand U5146 (N_5146,In_2041,In_134);
xnor U5147 (N_5147,In_267,In_2138);
nand U5148 (N_5148,In_1339,In_875);
and U5149 (N_5149,In_288,In_2022);
xnor U5150 (N_5150,In_416,In_2352);
or U5151 (N_5151,In_273,In_2051);
or U5152 (N_5152,In_2490,In_2094);
and U5153 (N_5153,In_1618,In_255);
and U5154 (N_5154,In_1690,In_384);
xnor U5155 (N_5155,In_1449,In_2778);
xnor U5156 (N_5156,In_2014,In_932);
nand U5157 (N_5157,In_958,In_2291);
nor U5158 (N_5158,In_2768,In_1555);
nor U5159 (N_5159,In_1617,In_1296);
nand U5160 (N_5160,In_1395,In_2352);
or U5161 (N_5161,In_2550,In_698);
nor U5162 (N_5162,In_95,In_1055);
nand U5163 (N_5163,In_1719,In_1190);
nor U5164 (N_5164,In_2752,In_1253);
and U5165 (N_5165,In_1410,In_2750);
nand U5166 (N_5166,In_420,In_1344);
xor U5167 (N_5167,In_2620,In_1578);
or U5168 (N_5168,In_1808,In_2616);
xnor U5169 (N_5169,In_2490,In_2903);
nand U5170 (N_5170,In_1968,In_1899);
and U5171 (N_5171,In_2385,In_1443);
nand U5172 (N_5172,In_2213,In_649);
xor U5173 (N_5173,In_2783,In_2045);
nor U5174 (N_5174,In_2153,In_2779);
or U5175 (N_5175,In_2659,In_493);
or U5176 (N_5176,In_2784,In_2393);
or U5177 (N_5177,In_2763,In_2556);
xor U5178 (N_5178,In_2906,In_2444);
xor U5179 (N_5179,In_1578,In_1901);
and U5180 (N_5180,In_2971,In_1065);
and U5181 (N_5181,In_937,In_1129);
and U5182 (N_5182,In_963,In_2632);
or U5183 (N_5183,In_2067,In_1749);
xnor U5184 (N_5184,In_2896,In_1039);
and U5185 (N_5185,In_2379,In_209);
and U5186 (N_5186,In_1033,In_1213);
and U5187 (N_5187,In_2710,In_1095);
xor U5188 (N_5188,In_12,In_2355);
nand U5189 (N_5189,In_1725,In_278);
nor U5190 (N_5190,In_2112,In_1547);
or U5191 (N_5191,In_630,In_2232);
and U5192 (N_5192,In_2399,In_1013);
nand U5193 (N_5193,In_1461,In_2789);
and U5194 (N_5194,In_2361,In_114);
and U5195 (N_5195,In_781,In_416);
and U5196 (N_5196,In_2775,In_226);
or U5197 (N_5197,In_2532,In_192);
and U5198 (N_5198,In_2647,In_930);
nor U5199 (N_5199,In_2691,In_1349);
nor U5200 (N_5200,In_1458,In_1487);
nand U5201 (N_5201,In_1991,In_2218);
nand U5202 (N_5202,In_2758,In_1231);
or U5203 (N_5203,In_1455,In_1366);
nor U5204 (N_5204,In_2331,In_2352);
xor U5205 (N_5205,In_2849,In_139);
xnor U5206 (N_5206,In_2762,In_2778);
and U5207 (N_5207,In_1948,In_2214);
xnor U5208 (N_5208,In_2308,In_1894);
nor U5209 (N_5209,In_2832,In_2567);
nand U5210 (N_5210,In_2301,In_1425);
xor U5211 (N_5211,In_861,In_2602);
nand U5212 (N_5212,In_2098,In_2941);
xnor U5213 (N_5213,In_90,In_1036);
nor U5214 (N_5214,In_2807,In_1079);
nor U5215 (N_5215,In_1025,In_273);
or U5216 (N_5216,In_2193,In_2732);
or U5217 (N_5217,In_304,In_125);
or U5218 (N_5218,In_770,In_2282);
nand U5219 (N_5219,In_964,In_1236);
xor U5220 (N_5220,In_936,In_2508);
or U5221 (N_5221,In_2785,In_508);
nand U5222 (N_5222,In_1207,In_1855);
and U5223 (N_5223,In_990,In_2583);
nor U5224 (N_5224,In_736,In_1125);
xnor U5225 (N_5225,In_1797,In_760);
or U5226 (N_5226,In_2749,In_1645);
nand U5227 (N_5227,In_32,In_1888);
xnor U5228 (N_5228,In_2713,In_402);
xnor U5229 (N_5229,In_1935,In_1674);
and U5230 (N_5230,In_2174,In_589);
or U5231 (N_5231,In_2484,In_2758);
nor U5232 (N_5232,In_2987,In_1621);
or U5233 (N_5233,In_471,In_309);
and U5234 (N_5234,In_32,In_776);
nor U5235 (N_5235,In_744,In_237);
or U5236 (N_5236,In_2867,In_1848);
nor U5237 (N_5237,In_908,In_2683);
and U5238 (N_5238,In_1921,In_2502);
and U5239 (N_5239,In_955,In_946);
nand U5240 (N_5240,In_2751,In_520);
nand U5241 (N_5241,In_239,In_47);
nor U5242 (N_5242,In_2947,In_2424);
and U5243 (N_5243,In_441,In_985);
or U5244 (N_5244,In_488,In_1872);
or U5245 (N_5245,In_1509,In_57);
xnor U5246 (N_5246,In_1181,In_2103);
xnor U5247 (N_5247,In_1383,In_979);
xor U5248 (N_5248,In_2527,In_265);
and U5249 (N_5249,In_2418,In_1906);
nor U5250 (N_5250,In_2566,In_1029);
nor U5251 (N_5251,In_1618,In_1773);
and U5252 (N_5252,In_2102,In_1979);
nand U5253 (N_5253,In_2806,In_695);
nand U5254 (N_5254,In_547,In_2527);
and U5255 (N_5255,In_1717,In_984);
or U5256 (N_5256,In_1031,In_2278);
nand U5257 (N_5257,In_2686,In_791);
nor U5258 (N_5258,In_2941,In_1029);
and U5259 (N_5259,In_1696,In_67);
or U5260 (N_5260,In_960,In_2694);
nor U5261 (N_5261,In_1880,In_58);
nand U5262 (N_5262,In_700,In_2834);
xor U5263 (N_5263,In_434,In_2151);
or U5264 (N_5264,In_1333,In_2400);
nor U5265 (N_5265,In_558,In_419);
xor U5266 (N_5266,In_882,In_614);
nor U5267 (N_5267,In_1363,In_826);
or U5268 (N_5268,In_816,In_168);
nand U5269 (N_5269,In_1363,In_866);
or U5270 (N_5270,In_880,In_1187);
and U5271 (N_5271,In_1007,In_931);
xor U5272 (N_5272,In_2051,In_602);
nand U5273 (N_5273,In_216,In_777);
nor U5274 (N_5274,In_1984,In_2847);
and U5275 (N_5275,In_653,In_341);
or U5276 (N_5276,In_1728,In_1779);
or U5277 (N_5277,In_788,In_439);
xor U5278 (N_5278,In_1680,In_1328);
xor U5279 (N_5279,In_1231,In_935);
xor U5280 (N_5280,In_2169,In_2566);
and U5281 (N_5281,In_1342,In_2202);
or U5282 (N_5282,In_1368,In_1145);
and U5283 (N_5283,In_2608,In_2176);
nand U5284 (N_5284,In_1148,In_977);
xnor U5285 (N_5285,In_1509,In_1587);
and U5286 (N_5286,In_1814,In_2175);
xor U5287 (N_5287,In_1103,In_2323);
nand U5288 (N_5288,In_1338,In_2794);
or U5289 (N_5289,In_909,In_760);
nand U5290 (N_5290,In_719,In_2407);
nand U5291 (N_5291,In_1060,In_579);
xnor U5292 (N_5292,In_806,In_242);
and U5293 (N_5293,In_1487,In_2685);
nand U5294 (N_5294,In_1903,In_71);
nor U5295 (N_5295,In_958,In_1308);
xor U5296 (N_5296,In_2821,In_1678);
or U5297 (N_5297,In_224,In_1161);
nand U5298 (N_5298,In_349,In_252);
nand U5299 (N_5299,In_718,In_1608);
nand U5300 (N_5300,In_2855,In_915);
and U5301 (N_5301,In_1143,In_1779);
nor U5302 (N_5302,In_1078,In_960);
nand U5303 (N_5303,In_1819,In_383);
and U5304 (N_5304,In_1370,In_2106);
xor U5305 (N_5305,In_82,In_1240);
xnor U5306 (N_5306,In_177,In_2842);
or U5307 (N_5307,In_2930,In_69);
xnor U5308 (N_5308,In_1455,In_2899);
or U5309 (N_5309,In_526,In_759);
nand U5310 (N_5310,In_1517,In_818);
or U5311 (N_5311,In_716,In_1598);
xnor U5312 (N_5312,In_858,In_1199);
or U5313 (N_5313,In_2672,In_1050);
nand U5314 (N_5314,In_1099,In_770);
xnor U5315 (N_5315,In_60,In_2116);
or U5316 (N_5316,In_148,In_809);
nor U5317 (N_5317,In_1438,In_2449);
nand U5318 (N_5318,In_2026,In_2882);
nor U5319 (N_5319,In_68,In_1699);
nand U5320 (N_5320,In_2669,In_1064);
and U5321 (N_5321,In_1725,In_2779);
or U5322 (N_5322,In_1102,In_1104);
nand U5323 (N_5323,In_1483,In_351);
and U5324 (N_5324,In_1128,In_2079);
nand U5325 (N_5325,In_1525,In_2132);
and U5326 (N_5326,In_967,In_1412);
or U5327 (N_5327,In_1751,In_2363);
xnor U5328 (N_5328,In_2917,In_1485);
and U5329 (N_5329,In_939,In_1745);
or U5330 (N_5330,In_1060,In_526);
xnor U5331 (N_5331,In_388,In_1194);
nand U5332 (N_5332,In_1813,In_576);
nand U5333 (N_5333,In_950,In_333);
nand U5334 (N_5334,In_1695,In_294);
xnor U5335 (N_5335,In_172,In_1540);
nor U5336 (N_5336,In_1906,In_836);
xor U5337 (N_5337,In_1829,In_1618);
nor U5338 (N_5338,In_773,In_1274);
nand U5339 (N_5339,In_1128,In_2382);
xor U5340 (N_5340,In_2557,In_2295);
nor U5341 (N_5341,In_1438,In_137);
nand U5342 (N_5342,In_2158,In_1950);
nor U5343 (N_5343,In_776,In_955);
nor U5344 (N_5344,In_274,In_2911);
nand U5345 (N_5345,In_2678,In_1115);
or U5346 (N_5346,In_2271,In_2001);
nand U5347 (N_5347,In_507,In_1500);
nand U5348 (N_5348,In_748,In_743);
nor U5349 (N_5349,In_784,In_410);
nor U5350 (N_5350,In_1528,In_2550);
xnor U5351 (N_5351,In_2850,In_560);
nand U5352 (N_5352,In_2580,In_233);
nor U5353 (N_5353,In_213,In_795);
nor U5354 (N_5354,In_63,In_1875);
and U5355 (N_5355,In_2198,In_2434);
nor U5356 (N_5356,In_960,In_311);
and U5357 (N_5357,In_1822,In_1759);
nand U5358 (N_5358,In_2098,In_633);
and U5359 (N_5359,In_2746,In_1563);
and U5360 (N_5360,In_275,In_675);
and U5361 (N_5361,In_552,In_2613);
and U5362 (N_5362,In_623,In_2997);
nand U5363 (N_5363,In_62,In_1606);
nor U5364 (N_5364,In_2364,In_167);
nor U5365 (N_5365,In_975,In_1646);
xnor U5366 (N_5366,In_858,In_2478);
xnor U5367 (N_5367,In_1226,In_2761);
and U5368 (N_5368,In_887,In_86);
nor U5369 (N_5369,In_1927,In_322);
nand U5370 (N_5370,In_888,In_1359);
nand U5371 (N_5371,In_2115,In_131);
nand U5372 (N_5372,In_469,In_1191);
or U5373 (N_5373,In_1414,In_2896);
nand U5374 (N_5374,In_1524,In_376);
xor U5375 (N_5375,In_2007,In_1601);
nand U5376 (N_5376,In_1346,In_1282);
nor U5377 (N_5377,In_1142,In_651);
or U5378 (N_5378,In_2625,In_646);
nand U5379 (N_5379,In_1685,In_2777);
nor U5380 (N_5380,In_425,In_2713);
and U5381 (N_5381,In_1210,In_2501);
or U5382 (N_5382,In_1770,In_2850);
and U5383 (N_5383,In_1983,In_1352);
xnor U5384 (N_5384,In_2168,In_875);
or U5385 (N_5385,In_490,In_2259);
xnor U5386 (N_5386,In_2140,In_1155);
or U5387 (N_5387,In_2917,In_393);
nor U5388 (N_5388,In_1759,In_2177);
xor U5389 (N_5389,In_594,In_48);
and U5390 (N_5390,In_2661,In_698);
xor U5391 (N_5391,In_1173,In_1163);
or U5392 (N_5392,In_702,In_2773);
xnor U5393 (N_5393,In_877,In_2399);
or U5394 (N_5394,In_1981,In_573);
xnor U5395 (N_5395,In_1994,In_635);
nand U5396 (N_5396,In_1924,In_7);
nor U5397 (N_5397,In_1827,In_165);
xor U5398 (N_5398,In_1513,In_145);
xnor U5399 (N_5399,In_1488,In_1723);
nor U5400 (N_5400,In_2325,In_2889);
nand U5401 (N_5401,In_1892,In_591);
and U5402 (N_5402,In_1468,In_400);
and U5403 (N_5403,In_241,In_2137);
xnor U5404 (N_5404,In_902,In_1973);
xor U5405 (N_5405,In_2648,In_2689);
xnor U5406 (N_5406,In_1743,In_1380);
xnor U5407 (N_5407,In_154,In_245);
and U5408 (N_5408,In_130,In_561);
and U5409 (N_5409,In_1606,In_772);
nand U5410 (N_5410,In_1906,In_2931);
nor U5411 (N_5411,In_1930,In_1046);
nor U5412 (N_5412,In_803,In_2920);
nand U5413 (N_5413,In_1072,In_2780);
and U5414 (N_5414,In_1294,In_2010);
nor U5415 (N_5415,In_670,In_2860);
or U5416 (N_5416,In_1104,In_919);
nand U5417 (N_5417,In_1791,In_80);
or U5418 (N_5418,In_2439,In_1923);
and U5419 (N_5419,In_912,In_181);
nand U5420 (N_5420,In_1968,In_1833);
or U5421 (N_5421,In_2191,In_2433);
or U5422 (N_5422,In_2015,In_2613);
nor U5423 (N_5423,In_425,In_2954);
nand U5424 (N_5424,In_947,In_762);
and U5425 (N_5425,In_2126,In_1349);
or U5426 (N_5426,In_2625,In_1752);
nand U5427 (N_5427,In_1209,In_1846);
nand U5428 (N_5428,In_9,In_113);
and U5429 (N_5429,In_2116,In_1716);
nor U5430 (N_5430,In_2879,In_1763);
nor U5431 (N_5431,In_1055,In_2234);
nand U5432 (N_5432,In_2041,In_2606);
and U5433 (N_5433,In_1308,In_2688);
nor U5434 (N_5434,In_1350,In_2214);
nand U5435 (N_5435,In_2135,In_2477);
and U5436 (N_5436,In_513,In_2545);
or U5437 (N_5437,In_1279,In_1578);
nor U5438 (N_5438,In_2550,In_1483);
or U5439 (N_5439,In_986,In_2091);
or U5440 (N_5440,In_1725,In_1416);
nand U5441 (N_5441,In_1655,In_458);
nor U5442 (N_5442,In_2618,In_156);
xnor U5443 (N_5443,In_1313,In_2063);
and U5444 (N_5444,In_2885,In_457);
nor U5445 (N_5445,In_802,In_204);
xnor U5446 (N_5446,In_2358,In_113);
or U5447 (N_5447,In_2270,In_1981);
and U5448 (N_5448,In_1915,In_2705);
or U5449 (N_5449,In_2949,In_1278);
or U5450 (N_5450,In_1982,In_2533);
nand U5451 (N_5451,In_1250,In_2064);
nor U5452 (N_5452,In_944,In_1576);
nand U5453 (N_5453,In_1686,In_2384);
or U5454 (N_5454,In_842,In_2033);
or U5455 (N_5455,In_1974,In_332);
or U5456 (N_5456,In_408,In_2270);
and U5457 (N_5457,In_1951,In_81);
nand U5458 (N_5458,In_230,In_2663);
xnor U5459 (N_5459,In_2293,In_979);
xnor U5460 (N_5460,In_1878,In_1793);
xnor U5461 (N_5461,In_155,In_2596);
and U5462 (N_5462,In_2210,In_2441);
nor U5463 (N_5463,In_2399,In_2433);
xnor U5464 (N_5464,In_1185,In_2110);
nor U5465 (N_5465,In_1079,In_1118);
xor U5466 (N_5466,In_962,In_1606);
or U5467 (N_5467,In_407,In_2537);
xnor U5468 (N_5468,In_2780,In_196);
or U5469 (N_5469,In_1056,In_2586);
nand U5470 (N_5470,In_1635,In_1759);
and U5471 (N_5471,In_2770,In_76);
nand U5472 (N_5472,In_1623,In_2341);
xor U5473 (N_5473,In_2463,In_1302);
nand U5474 (N_5474,In_1557,In_225);
nand U5475 (N_5475,In_2295,In_1764);
or U5476 (N_5476,In_1075,In_2832);
and U5477 (N_5477,In_1684,In_2266);
or U5478 (N_5478,In_482,In_1229);
xnor U5479 (N_5479,In_2350,In_1638);
and U5480 (N_5480,In_2609,In_964);
and U5481 (N_5481,In_1445,In_2991);
or U5482 (N_5482,In_1460,In_384);
nor U5483 (N_5483,In_1758,In_1690);
and U5484 (N_5484,In_501,In_2365);
nand U5485 (N_5485,In_2167,In_1170);
xnor U5486 (N_5486,In_2088,In_2882);
nand U5487 (N_5487,In_885,In_1295);
and U5488 (N_5488,In_36,In_2177);
nand U5489 (N_5489,In_2676,In_2513);
nor U5490 (N_5490,In_65,In_1831);
or U5491 (N_5491,In_1991,In_1305);
nand U5492 (N_5492,In_2196,In_2081);
or U5493 (N_5493,In_1898,In_2099);
or U5494 (N_5494,In_1567,In_396);
xnor U5495 (N_5495,In_1682,In_2707);
xnor U5496 (N_5496,In_2569,In_1687);
xnor U5497 (N_5497,In_1180,In_1115);
or U5498 (N_5498,In_1648,In_1696);
or U5499 (N_5499,In_610,In_1878);
nor U5500 (N_5500,In_2659,In_2481);
nand U5501 (N_5501,In_884,In_1329);
nand U5502 (N_5502,In_1587,In_2605);
or U5503 (N_5503,In_146,In_1069);
nand U5504 (N_5504,In_432,In_2894);
or U5505 (N_5505,In_536,In_2247);
xnor U5506 (N_5506,In_1337,In_1253);
xor U5507 (N_5507,In_513,In_16);
nor U5508 (N_5508,In_1272,In_2626);
and U5509 (N_5509,In_982,In_2670);
xor U5510 (N_5510,In_2838,In_2348);
and U5511 (N_5511,In_2243,In_242);
nand U5512 (N_5512,In_1796,In_386);
nand U5513 (N_5513,In_1723,In_565);
xor U5514 (N_5514,In_1471,In_992);
and U5515 (N_5515,In_1048,In_1407);
xnor U5516 (N_5516,In_2323,In_359);
xor U5517 (N_5517,In_430,In_1445);
nor U5518 (N_5518,In_2381,In_870);
nor U5519 (N_5519,In_1260,In_880);
nand U5520 (N_5520,In_1342,In_2699);
xor U5521 (N_5521,In_2059,In_1865);
nor U5522 (N_5522,In_1311,In_1051);
and U5523 (N_5523,In_1269,In_1507);
nand U5524 (N_5524,In_607,In_1965);
nand U5525 (N_5525,In_2519,In_2299);
nor U5526 (N_5526,In_2937,In_79);
nand U5527 (N_5527,In_137,In_818);
nand U5528 (N_5528,In_1222,In_2127);
or U5529 (N_5529,In_1107,In_1793);
or U5530 (N_5530,In_937,In_180);
or U5531 (N_5531,In_555,In_2515);
nor U5532 (N_5532,In_1095,In_2576);
nand U5533 (N_5533,In_745,In_574);
and U5534 (N_5534,In_2644,In_1811);
nand U5535 (N_5535,In_504,In_700);
or U5536 (N_5536,In_458,In_785);
nor U5537 (N_5537,In_58,In_2056);
and U5538 (N_5538,In_2399,In_1265);
xnor U5539 (N_5539,In_950,In_1446);
xnor U5540 (N_5540,In_2441,In_2443);
xor U5541 (N_5541,In_1872,In_1753);
xnor U5542 (N_5542,In_577,In_1042);
or U5543 (N_5543,In_1899,In_2328);
xnor U5544 (N_5544,In_1766,In_1928);
nor U5545 (N_5545,In_2778,In_2975);
nand U5546 (N_5546,In_2639,In_2163);
nor U5547 (N_5547,In_2122,In_2656);
and U5548 (N_5548,In_2769,In_1344);
or U5549 (N_5549,In_2866,In_2466);
nor U5550 (N_5550,In_435,In_2926);
or U5551 (N_5551,In_1172,In_842);
xnor U5552 (N_5552,In_253,In_2754);
xnor U5553 (N_5553,In_1183,In_315);
xnor U5554 (N_5554,In_2788,In_1124);
nand U5555 (N_5555,In_1137,In_813);
or U5556 (N_5556,In_1968,In_22);
nand U5557 (N_5557,In_1726,In_1417);
or U5558 (N_5558,In_787,In_478);
nand U5559 (N_5559,In_1544,In_2967);
and U5560 (N_5560,In_1467,In_266);
nor U5561 (N_5561,In_1658,In_2543);
nor U5562 (N_5562,In_1566,In_976);
and U5563 (N_5563,In_216,In_2006);
or U5564 (N_5564,In_155,In_1184);
xor U5565 (N_5565,In_84,In_2013);
nand U5566 (N_5566,In_81,In_2141);
nand U5567 (N_5567,In_1933,In_1356);
nand U5568 (N_5568,In_1154,In_1199);
nand U5569 (N_5569,In_2400,In_182);
nand U5570 (N_5570,In_1668,In_172);
nand U5571 (N_5571,In_366,In_339);
xor U5572 (N_5572,In_152,In_1145);
nand U5573 (N_5573,In_2441,In_1867);
nand U5574 (N_5574,In_839,In_2914);
nand U5575 (N_5575,In_2293,In_1586);
and U5576 (N_5576,In_1218,In_2179);
nor U5577 (N_5577,In_1955,In_1221);
nand U5578 (N_5578,In_1800,In_2072);
nor U5579 (N_5579,In_2752,In_1046);
or U5580 (N_5580,In_1461,In_1939);
nor U5581 (N_5581,In_1381,In_2831);
or U5582 (N_5582,In_767,In_594);
nor U5583 (N_5583,In_752,In_1503);
nand U5584 (N_5584,In_1154,In_1616);
or U5585 (N_5585,In_2250,In_2393);
nor U5586 (N_5586,In_1743,In_1213);
or U5587 (N_5587,In_2307,In_2672);
nor U5588 (N_5588,In_1335,In_733);
nor U5589 (N_5589,In_1983,In_92);
xnor U5590 (N_5590,In_2030,In_2788);
or U5591 (N_5591,In_920,In_1808);
nand U5592 (N_5592,In_2342,In_2244);
and U5593 (N_5593,In_1783,In_1194);
nor U5594 (N_5594,In_1964,In_1182);
nor U5595 (N_5595,In_185,In_419);
nor U5596 (N_5596,In_2194,In_2561);
nand U5597 (N_5597,In_739,In_2073);
xor U5598 (N_5598,In_737,In_305);
nor U5599 (N_5599,In_1677,In_1334);
nand U5600 (N_5600,In_160,In_1941);
or U5601 (N_5601,In_2786,In_1747);
and U5602 (N_5602,In_1541,In_1307);
or U5603 (N_5603,In_800,In_2187);
and U5604 (N_5604,In_1073,In_1872);
or U5605 (N_5605,In_2086,In_166);
xnor U5606 (N_5606,In_455,In_602);
or U5607 (N_5607,In_1179,In_230);
nand U5608 (N_5608,In_1369,In_1322);
xor U5609 (N_5609,In_840,In_1516);
nand U5610 (N_5610,In_2791,In_2216);
or U5611 (N_5611,In_479,In_2635);
or U5612 (N_5612,In_2222,In_278);
or U5613 (N_5613,In_1112,In_965);
xor U5614 (N_5614,In_834,In_2345);
or U5615 (N_5615,In_1160,In_1384);
and U5616 (N_5616,In_129,In_2893);
or U5617 (N_5617,In_2406,In_307);
xor U5618 (N_5618,In_865,In_2669);
nand U5619 (N_5619,In_777,In_599);
xnor U5620 (N_5620,In_780,In_2267);
and U5621 (N_5621,In_1014,In_1272);
xor U5622 (N_5622,In_1604,In_928);
nor U5623 (N_5623,In_1886,In_1809);
or U5624 (N_5624,In_2384,In_2618);
xor U5625 (N_5625,In_560,In_1164);
xnor U5626 (N_5626,In_876,In_1811);
and U5627 (N_5627,In_1425,In_1083);
nand U5628 (N_5628,In_2258,In_673);
nor U5629 (N_5629,In_2249,In_1985);
nand U5630 (N_5630,In_1058,In_1174);
xnor U5631 (N_5631,In_2108,In_1333);
or U5632 (N_5632,In_1778,In_50);
nor U5633 (N_5633,In_1564,In_493);
xnor U5634 (N_5634,In_2823,In_2247);
xor U5635 (N_5635,In_675,In_1446);
nand U5636 (N_5636,In_1551,In_683);
xor U5637 (N_5637,In_2799,In_1410);
and U5638 (N_5638,In_349,In_2795);
and U5639 (N_5639,In_1271,In_2666);
or U5640 (N_5640,In_682,In_1102);
and U5641 (N_5641,In_278,In_1517);
and U5642 (N_5642,In_2804,In_1392);
nor U5643 (N_5643,In_2329,In_454);
xnor U5644 (N_5644,In_2469,In_941);
nand U5645 (N_5645,In_2968,In_1740);
nor U5646 (N_5646,In_190,In_2362);
or U5647 (N_5647,In_1261,In_880);
xor U5648 (N_5648,In_2186,In_312);
or U5649 (N_5649,In_2445,In_105);
nand U5650 (N_5650,In_2214,In_1496);
nor U5651 (N_5651,In_1284,In_2147);
nand U5652 (N_5652,In_2925,In_1196);
and U5653 (N_5653,In_539,In_835);
nor U5654 (N_5654,In_1572,In_2276);
nor U5655 (N_5655,In_1768,In_2415);
or U5656 (N_5656,In_245,In_62);
or U5657 (N_5657,In_1034,In_1581);
or U5658 (N_5658,In_1034,In_2799);
or U5659 (N_5659,In_1292,In_2860);
and U5660 (N_5660,In_2040,In_2217);
and U5661 (N_5661,In_2132,In_1997);
nor U5662 (N_5662,In_276,In_2082);
or U5663 (N_5663,In_42,In_2047);
xnor U5664 (N_5664,In_2388,In_2653);
xnor U5665 (N_5665,In_2944,In_1416);
nand U5666 (N_5666,In_76,In_2435);
nor U5667 (N_5667,In_2588,In_2740);
or U5668 (N_5668,In_2659,In_1731);
and U5669 (N_5669,In_1636,In_2687);
nor U5670 (N_5670,In_1821,In_2935);
or U5671 (N_5671,In_398,In_1951);
and U5672 (N_5672,In_2849,In_1535);
xor U5673 (N_5673,In_1686,In_707);
and U5674 (N_5674,In_655,In_893);
and U5675 (N_5675,In_1068,In_994);
xor U5676 (N_5676,In_2722,In_993);
xnor U5677 (N_5677,In_793,In_1727);
or U5678 (N_5678,In_1372,In_2681);
nor U5679 (N_5679,In_1236,In_2662);
and U5680 (N_5680,In_2280,In_734);
or U5681 (N_5681,In_2732,In_1968);
xor U5682 (N_5682,In_1625,In_1307);
xor U5683 (N_5683,In_1402,In_2112);
nor U5684 (N_5684,In_1001,In_99);
and U5685 (N_5685,In_18,In_790);
nand U5686 (N_5686,In_1517,In_510);
nand U5687 (N_5687,In_626,In_1965);
nor U5688 (N_5688,In_2017,In_1325);
or U5689 (N_5689,In_821,In_2730);
nor U5690 (N_5690,In_1819,In_1447);
and U5691 (N_5691,In_340,In_1877);
nor U5692 (N_5692,In_2423,In_2303);
nor U5693 (N_5693,In_2666,In_1131);
nand U5694 (N_5694,In_1622,In_562);
and U5695 (N_5695,In_1086,In_2249);
and U5696 (N_5696,In_2193,In_1676);
nor U5697 (N_5697,In_2247,In_2067);
and U5698 (N_5698,In_1041,In_1520);
and U5699 (N_5699,In_1815,In_1805);
and U5700 (N_5700,In_510,In_1689);
nor U5701 (N_5701,In_445,In_115);
nand U5702 (N_5702,In_1149,In_2027);
and U5703 (N_5703,In_745,In_1116);
nand U5704 (N_5704,In_616,In_2498);
nand U5705 (N_5705,In_959,In_479);
or U5706 (N_5706,In_810,In_1691);
xor U5707 (N_5707,In_1600,In_1766);
and U5708 (N_5708,In_2884,In_1858);
xor U5709 (N_5709,In_220,In_1483);
nand U5710 (N_5710,In_2480,In_1022);
xnor U5711 (N_5711,In_1394,In_1806);
nand U5712 (N_5712,In_102,In_351);
or U5713 (N_5713,In_2969,In_408);
or U5714 (N_5714,In_1644,In_2315);
or U5715 (N_5715,In_2004,In_2072);
and U5716 (N_5716,In_527,In_1087);
xnor U5717 (N_5717,In_2238,In_1867);
nand U5718 (N_5718,In_717,In_2111);
or U5719 (N_5719,In_516,In_2352);
and U5720 (N_5720,In_1572,In_2529);
or U5721 (N_5721,In_1024,In_1719);
nor U5722 (N_5722,In_2611,In_878);
and U5723 (N_5723,In_2923,In_514);
xnor U5724 (N_5724,In_815,In_2113);
nand U5725 (N_5725,In_1010,In_2441);
nor U5726 (N_5726,In_768,In_18);
and U5727 (N_5727,In_1411,In_924);
and U5728 (N_5728,In_2155,In_2097);
or U5729 (N_5729,In_2049,In_790);
nand U5730 (N_5730,In_2433,In_2053);
nor U5731 (N_5731,In_1578,In_597);
xnor U5732 (N_5732,In_1043,In_408);
or U5733 (N_5733,In_1393,In_1354);
nand U5734 (N_5734,In_1688,In_897);
or U5735 (N_5735,In_136,In_2892);
xnor U5736 (N_5736,In_1907,In_2877);
or U5737 (N_5737,In_548,In_1479);
nand U5738 (N_5738,In_1362,In_2142);
nand U5739 (N_5739,In_1006,In_991);
nor U5740 (N_5740,In_2310,In_2807);
and U5741 (N_5741,In_1384,In_1033);
nand U5742 (N_5742,In_2554,In_2375);
nor U5743 (N_5743,In_2833,In_2334);
nand U5744 (N_5744,In_2232,In_1216);
nor U5745 (N_5745,In_2994,In_699);
nand U5746 (N_5746,In_2508,In_2407);
nor U5747 (N_5747,In_1611,In_119);
nand U5748 (N_5748,In_1172,In_81);
or U5749 (N_5749,In_1854,In_2589);
nor U5750 (N_5750,In_367,In_802);
xor U5751 (N_5751,In_1865,In_2153);
and U5752 (N_5752,In_2550,In_100);
nor U5753 (N_5753,In_2792,In_833);
nor U5754 (N_5754,In_342,In_1339);
nand U5755 (N_5755,In_2182,In_374);
nor U5756 (N_5756,In_2701,In_1425);
nand U5757 (N_5757,In_2294,In_1736);
nand U5758 (N_5758,In_2340,In_2157);
or U5759 (N_5759,In_2541,In_1920);
nor U5760 (N_5760,In_216,In_1052);
nor U5761 (N_5761,In_1554,In_677);
xor U5762 (N_5762,In_2646,In_1604);
nor U5763 (N_5763,In_993,In_1157);
xor U5764 (N_5764,In_1587,In_179);
or U5765 (N_5765,In_2020,In_359);
xor U5766 (N_5766,In_1455,In_2356);
nor U5767 (N_5767,In_294,In_1755);
nor U5768 (N_5768,In_2615,In_2014);
or U5769 (N_5769,In_2912,In_707);
xnor U5770 (N_5770,In_1591,In_628);
nor U5771 (N_5771,In_2292,In_1693);
nor U5772 (N_5772,In_976,In_768);
nand U5773 (N_5773,In_106,In_2515);
or U5774 (N_5774,In_624,In_2932);
or U5775 (N_5775,In_203,In_2015);
and U5776 (N_5776,In_1493,In_1348);
nor U5777 (N_5777,In_655,In_1302);
or U5778 (N_5778,In_398,In_1930);
and U5779 (N_5779,In_1896,In_1169);
nand U5780 (N_5780,In_2511,In_2720);
xnor U5781 (N_5781,In_1912,In_2670);
and U5782 (N_5782,In_179,In_31);
and U5783 (N_5783,In_2945,In_526);
nand U5784 (N_5784,In_1885,In_1448);
or U5785 (N_5785,In_180,In_1712);
or U5786 (N_5786,In_723,In_1786);
nor U5787 (N_5787,In_2031,In_87);
or U5788 (N_5788,In_1033,In_2548);
or U5789 (N_5789,In_1475,In_17);
nand U5790 (N_5790,In_165,In_2589);
xor U5791 (N_5791,In_2273,In_1171);
nor U5792 (N_5792,In_1657,In_2573);
xor U5793 (N_5793,In_737,In_1268);
nand U5794 (N_5794,In_1671,In_1216);
nand U5795 (N_5795,In_1720,In_831);
or U5796 (N_5796,In_2967,In_1486);
or U5797 (N_5797,In_1916,In_309);
or U5798 (N_5798,In_2172,In_1696);
nor U5799 (N_5799,In_1551,In_1581);
and U5800 (N_5800,In_1538,In_2479);
nor U5801 (N_5801,In_1531,In_303);
or U5802 (N_5802,In_2454,In_2709);
and U5803 (N_5803,In_687,In_466);
and U5804 (N_5804,In_2672,In_392);
or U5805 (N_5805,In_650,In_1466);
nand U5806 (N_5806,In_1173,In_2024);
or U5807 (N_5807,In_665,In_1963);
or U5808 (N_5808,In_2527,In_1217);
nand U5809 (N_5809,In_1531,In_1029);
nand U5810 (N_5810,In_921,In_1835);
xnor U5811 (N_5811,In_1770,In_691);
and U5812 (N_5812,In_1729,In_2657);
or U5813 (N_5813,In_1469,In_2969);
or U5814 (N_5814,In_436,In_619);
nor U5815 (N_5815,In_1350,In_2512);
nand U5816 (N_5816,In_1147,In_1019);
or U5817 (N_5817,In_232,In_1526);
nor U5818 (N_5818,In_2000,In_181);
and U5819 (N_5819,In_1538,In_982);
xor U5820 (N_5820,In_800,In_348);
or U5821 (N_5821,In_2209,In_2674);
or U5822 (N_5822,In_1932,In_981);
or U5823 (N_5823,In_1898,In_1272);
and U5824 (N_5824,In_2379,In_456);
nand U5825 (N_5825,In_2592,In_2949);
nor U5826 (N_5826,In_1906,In_703);
xnor U5827 (N_5827,In_1826,In_1156);
xor U5828 (N_5828,In_1813,In_2453);
nor U5829 (N_5829,In_1994,In_1359);
or U5830 (N_5830,In_2875,In_110);
nor U5831 (N_5831,In_317,In_1730);
nor U5832 (N_5832,In_2748,In_2865);
nor U5833 (N_5833,In_2056,In_2997);
xor U5834 (N_5834,In_2029,In_1633);
nand U5835 (N_5835,In_1095,In_1927);
and U5836 (N_5836,In_1415,In_503);
nor U5837 (N_5837,In_1545,In_163);
nand U5838 (N_5838,In_2020,In_2285);
and U5839 (N_5839,In_2027,In_2474);
xnor U5840 (N_5840,In_1701,In_2112);
xor U5841 (N_5841,In_851,In_2344);
nor U5842 (N_5842,In_2916,In_1630);
xnor U5843 (N_5843,In_2336,In_929);
nor U5844 (N_5844,In_2907,In_1769);
xnor U5845 (N_5845,In_500,In_579);
nor U5846 (N_5846,In_2954,In_118);
nor U5847 (N_5847,In_1621,In_1120);
xnor U5848 (N_5848,In_2085,In_1645);
or U5849 (N_5849,In_1355,In_146);
nand U5850 (N_5850,In_713,In_2878);
nor U5851 (N_5851,In_39,In_497);
nand U5852 (N_5852,In_264,In_62);
and U5853 (N_5853,In_809,In_2190);
xor U5854 (N_5854,In_1815,In_276);
and U5855 (N_5855,In_574,In_2634);
nand U5856 (N_5856,In_2118,In_2541);
xnor U5857 (N_5857,In_1807,In_2318);
xor U5858 (N_5858,In_776,In_2165);
nor U5859 (N_5859,In_1176,In_2748);
nand U5860 (N_5860,In_2121,In_2553);
or U5861 (N_5861,In_1263,In_2636);
and U5862 (N_5862,In_2341,In_479);
xor U5863 (N_5863,In_725,In_963);
nand U5864 (N_5864,In_343,In_2632);
or U5865 (N_5865,In_2833,In_2304);
nor U5866 (N_5866,In_1762,In_490);
nor U5867 (N_5867,In_960,In_2149);
or U5868 (N_5868,In_360,In_1841);
nand U5869 (N_5869,In_565,In_2435);
nand U5870 (N_5870,In_2179,In_94);
xor U5871 (N_5871,In_2648,In_2198);
xnor U5872 (N_5872,In_2654,In_2970);
nor U5873 (N_5873,In_1494,In_2322);
nand U5874 (N_5874,In_805,In_290);
nand U5875 (N_5875,In_1750,In_1381);
nor U5876 (N_5876,In_788,In_1626);
and U5877 (N_5877,In_911,In_1406);
nor U5878 (N_5878,In_141,In_2044);
or U5879 (N_5879,In_1282,In_759);
and U5880 (N_5880,In_610,In_269);
nand U5881 (N_5881,In_1047,In_1009);
xor U5882 (N_5882,In_2216,In_655);
nand U5883 (N_5883,In_621,In_1767);
and U5884 (N_5884,In_116,In_2115);
or U5885 (N_5885,In_554,In_1252);
nand U5886 (N_5886,In_1697,In_1194);
xnor U5887 (N_5887,In_25,In_399);
or U5888 (N_5888,In_2465,In_2851);
nor U5889 (N_5889,In_2450,In_675);
nor U5890 (N_5890,In_985,In_555);
xnor U5891 (N_5891,In_573,In_451);
and U5892 (N_5892,In_926,In_266);
and U5893 (N_5893,In_528,In_1273);
or U5894 (N_5894,In_847,In_421);
xor U5895 (N_5895,In_2667,In_2757);
nand U5896 (N_5896,In_576,In_1439);
or U5897 (N_5897,In_1286,In_2060);
nor U5898 (N_5898,In_2758,In_362);
nand U5899 (N_5899,In_2250,In_1358);
xnor U5900 (N_5900,In_1634,In_182);
or U5901 (N_5901,In_2147,In_1064);
and U5902 (N_5902,In_1706,In_2193);
xor U5903 (N_5903,In_1172,In_1070);
xnor U5904 (N_5904,In_2559,In_629);
and U5905 (N_5905,In_2671,In_902);
nand U5906 (N_5906,In_1697,In_1420);
or U5907 (N_5907,In_779,In_455);
or U5908 (N_5908,In_946,In_2697);
and U5909 (N_5909,In_1947,In_2412);
or U5910 (N_5910,In_2238,In_915);
xor U5911 (N_5911,In_240,In_728);
nand U5912 (N_5912,In_421,In_148);
or U5913 (N_5913,In_1787,In_2023);
and U5914 (N_5914,In_1314,In_957);
xor U5915 (N_5915,In_1662,In_2973);
nor U5916 (N_5916,In_2084,In_2871);
xnor U5917 (N_5917,In_747,In_1481);
xnor U5918 (N_5918,In_1138,In_2517);
or U5919 (N_5919,In_1281,In_2728);
and U5920 (N_5920,In_1040,In_217);
or U5921 (N_5921,In_1581,In_844);
or U5922 (N_5922,In_2507,In_1547);
nor U5923 (N_5923,In_1323,In_2811);
xnor U5924 (N_5924,In_1526,In_1212);
and U5925 (N_5925,In_1601,In_2199);
and U5926 (N_5926,In_1726,In_404);
nor U5927 (N_5927,In_2858,In_2311);
nor U5928 (N_5928,In_1496,In_2678);
xor U5929 (N_5929,In_2201,In_2262);
or U5930 (N_5930,In_767,In_1041);
xnor U5931 (N_5931,In_1218,In_659);
nand U5932 (N_5932,In_2178,In_2367);
xnor U5933 (N_5933,In_877,In_1501);
nand U5934 (N_5934,In_451,In_624);
nor U5935 (N_5935,In_2667,In_2911);
xor U5936 (N_5936,In_262,In_2504);
nor U5937 (N_5937,In_2228,In_2954);
xnor U5938 (N_5938,In_1831,In_2618);
nor U5939 (N_5939,In_1088,In_527);
or U5940 (N_5940,In_2067,In_438);
nor U5941 (N_5941,In_1148,In_2167);
or U5942 (N_5942,In_2920,In_2035);
or U5943 (N_5943,In_708,In_1893);
and U5944 (N_5944,In_1986,In_2524);
nor U5945 (N_5945,In_2160,In_1052);
and U5946 (N_5946,In_1206,In_99);
nor U5947 (N_5947,In_2677,In_541);
xnor U5948 (N_5948,In_1655,In_1951);
nand U5949 (N_5949,In_1125,In_1349);
or U5950 (N_5950,In_1511,In_1345);
or U5951 (N_5951,In_2257,In_1281);
and U5952 (N_5952,In_1939,In_2610);
or U5953 (N_5953,In_2376,In_2173);
and U5954 (N_5954,In_1921,In_2427);
or U5955 (N_5955,In_2245,In_1461);
and U5956 (N_5956,In_290,In_672);
xor U5957 (N_5957,In_2130,In_1801);
nor U5958 (N_5958,In_587,In_2158);
nand U5959 (N_5959,In_2427,In_2946);
nand U5960 (N_5960,In_2276,In_1742);
or U5961 (N_5961,In_2158,In_2209);
and U5962 (N_5962,In_439,In_2138);
xor U5963 (N_5963,In_1806,In_1443);
xnor U5964 (N_5964,In_1769,In_2969);
and U5965 (N_5965,In_780,In_1372);
and U5966 (N_5966,In_1049,In_1886);
xor U5967 (N_5967,In_1134,In_1693);
or U5968 (N_5968,In_585,In_2758);
or U5969 (N_5969,In_574,In_2862);
nand U5970 (N_5970,In_106,In_2750);
and U5971 (N_5971,In_220,In_1790);
nand U5972 (N_5972,In_474,In_536);
and U5973 (N_5973,In_2609,In_2547);
and U5974 (N_5974,In_2740,In_950);
nand U5975 (N_5975,In_462,In_1164);
or U5976 (N_5976,In_1804,In_2406);
and U5977 (N_5977,In_1239,In_274);
and U5978 (N_5978,In_2919,In_384);
xnor U5979 (N_5979,In_2009,In_2733);
and U5980 (N_5980,In_2269,In_2005);
nand U5981 (N_5981,In_2488,In_2127);
or U5982 (N_5982,In_2453,In_648);
and U5983 (N_5983,In_1208,In_750);
xnor U5984 (N_5984,In_2759,In_1491);
and U5985 (N_5985,In_1598,In_101);
and U5986 (N_5986,In_1489,In_2574);
xnor U5987 (N_5987,In_2012,In_2852);
and U5988 (N_5988,In_2535,In_1342);
nand U5989 (N_5989,In_142,In_374);
xnor U5990 (N_5990,In_1919,In_2683);
nand U5991 (N_5991,In_2926,In_2326);
xnor U5992 (N_5992,In_2194,In_2032);
nor U5993 (N_5993,In_2619,In_1832);
nand U5994 (N_5994,In_1571,In_1062);
and U5995 (N_5995,In_2930,In_1925);
and U5996 (N_5996,In_1745,In_39);
or U5997 (N_5997,In_1658,In_2426);
and U5998 (N_5998,In_1826,In_231);
xor U5999 (N_5999,In_618,In_2792);
nor U6000 (N_6000,N_3694,N_2420);
nand U6001 (N_6001,N_1484,N_1341);
xnor U6002 (N_6002,N_1034,N_2228);
and U6003 (N_6003,N_1771,N_5402);
or U6004 (N_6004,N_4717,N_1903);
and U6005 (N_6005,N_1051,N_5894);
nor U6006 (N_6006,N_3081,N_2829);
nand U6007 (N_6007,N_4426,N_5395);
nor U6008 (N_6008,N_5887,N_2950);
and U6009 (N_6009,N_5265,N_4449);
nor U6010 (N_6010,N_5058,N_604);
xor U6011 (N_6011,N_952,N_639);
nand U6012 (N_6012,N_546,N_4036);
and U6013 (N_6013,N_1743,N_1878);
or U6014 (N_6014,N_3069,N_5637);
nand U6015 (N_6015,N_5740,N_2538);
and U6016 (N_6016,N_2512,N_3155);
and U6017 (N_6017,N_2004,N_4512);
and U6018 (N_6018,N_2428,N_3433);
nor U6019 (N_6019,N_2828,N_3643);
nand U6020 (N_6020,N_1798,N_4593);
or U6021 (N_6021,N_3921,N_4021);
and U6022 (N_6022,N_4911,N_3903);
or U6023 (N_6023,N_2199,N_3278);
nand U6024 (N_6024,N_3158,N_5112);
nor U6025 (N_6025,N_1014,N_192);
nor U6026 (N_6026,N_2594,N_2333);
nor U6027 (N_6027,N_5591,N_4012);
nor U6028 (N_6028,N_5042,N_4925);
or U6029 (N_6029,N_4746,N_3480);
nand U6030 (N_6030,N_5577,N_5775);
nand U6031 (N_6031,N_3030,N_818);
nand U6032 (N_6032,N_5700,N_4136);
and U6033 (N_6033,N_1809,N_2182);
nand U6034 (N_6034,N_3211,N_2591);
or U6035 (N_6035,N_3885,N_1176);
nand U6036 (N_6036,N_1331,N_4781);
nand U6037 (N_6037,N_2093,N_108);
or U6038 (N_6038,N_2364,N_4747);
nor U6039 (N_6039,N_5054,N_3843);
xnor U6040 (N_6040,N_3373,N_2602);
and U6041 (N_6041,N_419,N_1238);
and U6042 (N_6042,N_599,N_4713);
or U6043 (N_6043,N_5869,N_3127);
or U6044 (N_6044,N_418,N_4066);
xnor U6045 (N_6045,N_4608,N_3640);
nand U6046 (N_6046,N_4260,N_4529);
xor U6047 (N_6047,N_3840,N_3235);
or U6048 (N_6048,N_2571,N_2500);
nor U6049 (N_6049,N_5067,N_718);
nand U6050 (N_6050,N_2378,N_5852);
or U6051 (N_6051,N_822,N_1711);
xor U6052 (N_6052,N_3826,N_3602);
or U6053 (N_6053,N_1542,N_4722);
or U6054 (N_6054,N_3482,N_466);
nor U6055 (N_6055,N_2892,N_2032);
and U6056 (N_6056,N_4607,N_4114);
and U6057 (N_6057,N_669,N_5842);
nand U6058 (N_6058,N_1588,N_4708);
nor U6059 (N_6059,N_4896,N_4987);
or U6060 (N_6060,N_1157,N_3493);
and U6061 (N_6061,N_4615,N_452);
nand U6062 (N_6062,N_3120,N_139);
xnor U6063 (N_6063,N_980,N_1500);
xnor U6064 (N_6064,N_2643,N_4381);
or U6065 (N_6065,N_2907,N_40);
or U6066 (N_6066,N_2389,N_2120);
xor U6067 (N_6067,N_5335,N_699);
and U6068 (N_6068,N_371,N_2537);
nor U6069 (N_6069,N_1643,N_3291);
nand U6070 (N_6070,N_1653,N_4955);
nor U6071 (N_6071,N_5711,N_1892);
nand U6072 (N_6072,N_5464,N_2121);
xor U6073 (N_6073,N_4478,N_5032);
or U6074 (N_6074,N_4379,N_3626);
nor U6075 (N_6075,N_2436,N_4199);
xor U6076 (N_6076,N_310,N_5443);
nor U6077 (N_6077,N_3085,N_4762);
or U6078 (N_6078,N_4077,N_3404);
xnor U6079 (N_6079,N_3345,N_1082);
nor U6080 (N_6080,N_2175,N_4365);
nand U6081 (N_6081,N_4447,N_2999);
or U6082 (N_6082,N_3586,N_1921);
nor U6083 (N_6083,N_5837,N_709);
xnor U6084 (N_6084,N_2686,N_1391);
nand U6085 (N_6085,N_4366,N_3340);
nand U6086 (N_6086,N_412,N_2454);
nand U6087 (N_6087,N_5545,N_3572);
and U6088 (N_6088,N_107,N_3598);
nand U6089 (N_6089,N_4001,N_919);
and U6090 (N_6090,N_1307,N_2007);
nand U6091 (N_6091,N_4750,N_5612);
or U6092 (N_6092,N_1881,N_2746);
nand U6093 (N_6093,N_1482,N_413);
and U6094 (N_6094,N_5474,N_905);
or U6095 (N_6095,N_1069,N_3607);
and U6096 (N_6096,N_2026,N_491);
or U6097 (N_6097,N_1877,N_4929);
xor U6098 (N_6098,N_3204,N_2691);
xnor U6099 (N_6099,N_5087,N_4953);
nand U6100 (N_6100,N_702,N_5455);
or U6101 (N_6101,N_5777,N_3567);
and U6102 (N_6102,N_667,N_5975);
nand U6103 (N_6103,N_5841,N_5004);
and U6104 (N_6104,N_5799,N_5863);
and U6105 (N_6105,N_1362,N_2078);
xnor U6106 (N_6106,N_4129,N_4749);
or U6107 (N_6107,N_3017,N_2809);
and U6108 (N_6108,N_2158,N_1366);
and U6109 (N_6109,N_1987,N_1181);
and U6110 (N_6110,N_1053,N_1824);
nand U6111 (N_6111,N_5028,N_5206);
nand U6112 (N_6112,N_4906,N_3799);
nand U6113 (N_6113,N_42,N_740);
nand U6114 (N_6114,N_5737,N_1980);
or U6115 (N_6115,N_1978,N_5086);
nand U6116 (N_6116,N_605,N_1477);
or U6117 (N_6117,N_3000,N_1611);
and U6118 (N_6118,N_2190,N_4035);
nand U6119 (N_6119,N_2902,N_5245);
xnor U6120 (N_6120,N_14,N_3983);
xnor U6121 (N_6121,N_5131,N_2622);
nand U6122 (N_6122,N_1173,N_525);
nor U6123 (N_6123,N_2122,N_927);
nand U6124 (N_6124,N_370,N_4157);
and U6125 (N_6125,N_1690,N_2989);
or U6126 (N_6126,N_893,N_2468);
xnor U6127 (N_6127,N_1520,N_2363);
nand U6128 (N_6128,N_3776,N_4999);
nor U6129 (N_6129,N_202,N_3363);
nand U6130 (N_6130,N_4345,N_1349);
xor U6131 (N_6131,N_2849,N_463);
xor U6132 (N_6132,N_2943,N_4627);
and U6133 (N_6133,N_2618,N_2976);
and U6134 (N_6134,N_4149,N_4881);
xnor U6135 (N_6135,N_5676,N_5160);
and U6136 (N_6136,N_858,N_39);
nand U6137 (N_6137,N_1074,N_1540);
or U6138 (N_6138,N_4595,N_424);
nand U6139 (N_6139,N_159,N_4234);
xnor U6140 (N_6140,N_3312,N_1419);
nand U6141 (N_6141,N_5696,N_3320);
or U6142 (N_6142,N_1452,N_1265);
and U6143 (N_6143,N_4638,N_2164);
xnor U6144 (N_6144,N_813,N_403);
and U6145 (N_6145,N_5638,N_201);
and U6146 (N_6146,N_844,N_3819);
nand U6147 (N_6147,N_2337,N_5582);
nor U6148 (N_6148,N_4489,N_5651);
nand U6149 (N_6149,N_5529,N_5091);
or U6150 (N_6150,N_2697,N_2955);
nand U6151 (N_6151,N_1488,N_4903);
xor U6152 (N_6152,N_5022,N_2108);
or U6153 (N_6153,N_4098,N_3899);
xnor U6154 (N_6154,N_5300,N_5462);
nor U6155 (N_6155,N_544,N_5166);
or U6156 (N_6156,N_646,N_666);
or U6157 (N_6157,N_5321,N_4954);
and U6158 (N_6158,N_3760,N_2520);
nor U6159 (N_6159,N_4993,N_1188);
nand U6160 (N_6160,N_1775,N_157);
xnor U6161 (N_6161,N_5213,N_2814);
xnor U6162 (N_6162,N_2782,N_2394);
xor U6163 (N_6163,N_2321,N_5161);
nand U6164 (N_6164,N_2718,N_2716);
and U6165 (N_6165,N_2959,N_4828);
or U6166 (N_6166,N_4838,N_3835);
or U6167 (N_6167,N_3464,N_260);
and U6168 (N_6168,N_404,N_4554);
nor U6169 (N_6169,N_3279,N_3657);
xnor U6170 (N_6170,N_2731,N_2467);
nand U6171 (N_6171,N_5681,N_1544);
or U6172 (N_6172,N_712,N_4634);
xor U6173 (N_6173,N_2284,N_5619);
nand U6174 (N_6174,N_3653,N_1782);
xnor U6175 (N_6175,N_2864,N_5103);
and U6176 (N_6176,N_5795,N_5523);
or U6177 (N_6177,N_715,N_4885);
nand U6178 (N_6178,N_2605,N_2566);
xnor U6179 (N_6179,N_5480,N_2906);
or U6180 (N_6180,N_1143,N_488);
nand U6181 (N_6181,N_5561,N_4832);
and U6182 (N_6182,N_4636,N_5275);
xor U6183 (N_6183,N_3967,N_321);
and U6184 (N_6184,N_2752,N_5648);
or U6185 (N_6185,N_5401,N_4570);
nor U6186 (N_6186,N_1807,N_3829);
nand U6187 (N_6187,N_3578,N_5950);
or U6188 (N_6188,N_4960,N_4267);
xor U6189 (N_6189,N_4637,N_4068);
nor U6190 (N_6190,N_3744,N_975);
xnor U6191 (N_6191,N_5602,N_5763);
and U6192 (N_6192,N_129,N_868);
nand U6193 (N_6193,N_5753,N_4591);
nor U6194 (N_6194,N_3224,N_2744);
or U6195 (N_6195,N_2370,N_1663);
nor U6196 (N_6196,N_1167,N_3896);
nand U6197 (N_6197,N_135,N_1140);
nand U6198 (N_6198,N_5196,N_3528);
nor U6199 (N_6199,N_5437,N_4093);
or U6200 (N_6200,N_3001,N_2134);
or U6201 (N_6201,N_1744,N_3725);
and U6202 (N_6202,N_2625,N_4702);
nor U6203 (N_6203,N_3227,N_5885);
nor U6204 (N_6204,N_5834,N_5491);
nand U6205 (N_6205,N_802,N_2637);
xor U6206 (N_6206,N_4550,N_196);
nor U6207 (N_6207,N_4204,N_5949);
nand U6208 (N_6208,N_5666,N_278);
nor U6209 (N_6209,N_5438,N_5726);
nand U6210 (N_6210,N_1885,N_1563);
or U6211 (N_6211,N_656,N_4673);
and U6212 (N_6212,N_4401,N_3588);
nor U6213 (N_6213,N_3272,N_4775);
and U6214 (N_6214,N_1584,N_85);
nand U6215 (N_6215,N_3113,N_865);
or U6216 (N_6216,N_1989,N_2017);
or U6217 (N_6217,N_5027,N_811);
xor U6218 (N_6218,N_2434,N_4894);
or U6219 (N_6219,N_5796,N_2859);
and U6220 (N_6220,N_3396,N_4486);
xnor U6221 (N_6221,N_3476,N_2322);
and U6222 (N_6222,N_216,N_791);
xor U6223 (N_6223,N_1535,N_4241);
xor U6224 (N_6224,N_1360,N_90);
nand U6225 (N_6225,N_2210,N_62);
and U6226 (N_6226,N_970,N_5282);
xnor U6227 (N_6227,N_1624,N_1429);
nand U6228 (N_6228,N_3497,N_757);
xnor U6229 (N_6229,N_4000,N_4109);
xnor U6230 (N_6230,N_5544,N_5051);
nand U6231 (N_6231,N_2187,N_5844);
xor U6232 (N_6232,N_4210,N_2636);
and U6233 (N_6233,N_672,N_1379);
or U6234 (N_6234,N_3703,N_1061);
nor U6235 (N_6235,N_5147,N_5074);
or U6236 (N_6236,N_4473,N_3511);
nor U6237 (N_6237,N_4252,N_1505);
nor U6238 (N_6238,N_1297,N_5426);
nor U6239 (N_6239,N_5383,N_214);
xnor U6240 (N_6240,N_5185,N_5993);
and U6241 (N_6241,N_1043,N_4986);
nand U6242 (N_6242,N_3326,N_5351);
xor U6243 (N_6243,N_953,N_4823);
or U6244 (N_6244,N_2711,N_2839);
and U6245 (N_6245,N_737,N_1134);
nor U6246 (N_6246,N_2086,N_1722);
nor U6247 (N_6247,N_4744,N_1154);
and U6248 (N_6248,N_3372,N_2990);
nor U6249 (N_6249,N_3564,N_3397);
xnor U6250 (N_6250,N_2232,N_3797);
and U6251 (N_6251,N_2801,N_1677);
or U6252 (N_6252,N_3939,N_2014);
and U6253 (N_6253,N_4502,N_631);
xnor U6254 (N_6254,N_3745,N_978);
nor U6255 (N_6255,N_2547,N_1840);
nand U6256 (N_6256,N_5452,N_624);
and U6257 (N_6257,N_17,N_5492);
nor U6258 (N_6258,N_3680,N_711);
xor U6259 (N_6259,N_478,N_2088);
xnor U6260 (N_6260,N_5212,N_5498);
nand U6261 (N_6261,N_1103,N_4235);
or U6262 (N_6262,N_1764,N_206);
nand U6263 (N_6263,N_2802,N_5382);
nand U6264 (N_6264,N_272,N_5291);
xnor U6265 (N_6265,N_3946,N_4850);
nor U6266 (N_6266,N_1747,N_685);
and U6267 (N_6267,N_1511,N_4096);
nor U6268 (N_6268,N_3595,N_5961);
nor U6269 (N_6269,N_2267,N_227);
and U6270 (N_6270,N_183,N_365);
nand U6271 (N_6271,N_5013,N_955);
nand U6272 (N_6272,N_134,N_3505);
nor U6273 (N_6273,N_32,N_1669);
and U6274 (N_6274,N_5466,N_3398);
and U6275 (N_6275,N_3594,N_2162);
xor U6276 (N_6276,N_1376,N_326);
nor U6277 (N_6277,N_1905,N_5623);
nor U6278 (N_6278,N_723,N_901);
and U6279 (N_6279,N_4596,N_4263);
nand U6280 (N_6280,N_1417,N_2981);
or U6281 (N_6281,N_2488,N_4054);
or U6282 (N_6282,N_2576,N_1587);
xor U6283 (N_6283,N_4322,N_1378);
nand U6284 (N_6284,N_1739,N_5226);
nand U6285 (N_6285,N_1047,N_5862);
xnor U6286 (N_6286,N_3018,N_2805);
nand U6287 (N_6287,N_2312,N_2854);
nand U6288 (N_6288,N_826,N_5757);
xor U6289 (N_6289,N_998,N_5344);
and U6290 (N_6290,N_3804,N_4980);
xnor U6291 (N_6291,N_3263,N_854);
xnor U6292 (N_6292,N_512,N_1673);
and U6293 (N_6293,N_1105,N_843);
or U6294 (N_6294,N_5827,N_3850);
xor U6295 (N_6295,N_4847,N_4045);
and U6296 (N_6296,N_3977,N_835);
or U6297 (N_6297,N_3293,N_3292);
xor U6298 (N_6298,N_5512,N_575);
nor U6299 (N_6299,N_2174,N_3376);
nand U6300 (N_6300,N_5909,N_4148);
and U6301 (N_6301,N_2235,N_2180);
nor U6302 (N_6302,N_751,N_891);
or U6303 (N_6303,N_2393,N_4070);
xor U6304 (N_6304,N_4217,N_2114);
and U6305 (N_6305,N_3642,N_4534);
xor U6306 (N_6306,N_388,N_4058);
nand U6307 (N_6307,N_379,N_5428);
nor U6308 (N_6308,N_1699,N_5152);
nor U6309 (N_6309,N_5297,N_2001);
or U6310 (N_6310,N_4282,N_204);
and U6311 (N_6311,N_3683,N_1342);
or U6312 (N_6312,N_1182,N_3662);
and U6313 (N_6313,N_450,N_1800);
nor U6314 (N_6314,N_965,N_2964);
xnor U6315 (N_6315,N_1750,N_3690);
nand U6316 (N_6316,N_810,N_4716);
or U6317 (N_6317,N_3328,N_2740);
nand U6318 (N_6318,N_3050,N_290);
nand U6319 (N_6319,N_4536,N_4853);
nor U6320 (N_6320,N_1121,N_341);
xor U6321 (N_6321,N_4358,N_5957);
nor U6322 (N_6322,N_1539,N_89);
xnor U6323 (N_6323,N_5323,N_2720);
and U6324 (N_6324,N_3408,N_849);
xnor U6325 (N_6325,N_997,N_3086);
and U6326 (N_6326,N_1942,N_4569);
nor U6327 (N_6327,N_3118,N_427);
and U6328 (N_6328,N_4458,N_1597);
and U6329 (N_6329,N_1671,N_5843);
nand U6330 (N_6330,N_837,N_1760);
nor U6331 (N_6331,N_572,N_4089);
or U6332 (N_6332,N_1835,N_3230);
or U6333 (N_6333,N_4804,N_87);
nor U6334 (N_6334,N_4546,N_3632);
nor U6335 (N_6335,N_4496,N_877);
xnor U6336 (N_6336,N_4887,N_4539);
nor U6337 (N_6337,N_2067,N_4373);
and U6338 (N_6338,N_2830,N_4579);
xor U6339 (N_6339,N_2734,N_1296);
nor U6340 (N_6340,N_5913,N_3252);
xor U6341 (N_6341,N_3304,N_3898);
and U6342 (N_6342,N_2094,N_5072);
xor U6343 (N_6343,N_4545,N_1612);
nor U6344 (N_6344,N_3091,N_2459);
nand U6345 (N_6345,N_1943,N_446);
nor U6346 (N_6346,N_5195,N_3627);
nor U6347 (N_6347,N_3608,N_2935);
or U6348 (N_6348,N_5219,N_5965);
nand U6349 (N_6349,N_3707,N_212);
xnor U6350 (N_6350,N_1028,N_120);
nand U6351 (N_6351,N_1318,N_2497);
and U6352 (N_6352,N_3238,N_5202);
nor U6353 (N_6353,N_2745,N_2784);
nand U6354 (N_6354,N_4471,N_732);
nor U6355 (N_6355,N_4726,N_3256);
or U6356 (N_6356,N_4396,N_1995);
nand U6357 (N_6357,N_189,N_2865);
nor U6358 (N_6358,N_4564,N_547);
nand U6359 (N_6359,N_539,N_651);
xnor U6360 (N_6360,N_229,N_762);
nand U6361 (N_6361,N_4086,N_1490);
xor U6362 (N_6362,N_3167,N_2646);
and U6363 (N_6363,N_3334,N_2918);
xor U6364 (N_6364,N_5530,N_4841);
nor U6365 (N_6365,N_1434,N_435);
xor U6366 (N_6366,N_5399,N_155);
xor U6367 (N_6367,N_5257,N_4101);
xor U6368 (N_6368,N_951,N_2550);
and U6369 (N_6369,N_3992,N_5723);
and U6370 (N_6370,N_367,N_4150);
and U6371 (N_6371,N_4017,N_2823);
or U6372 (N_6372,N_4005,N_5653);
nand U6373 (N_6373,N_4644,N_608);
or U6374 (N_6374,N_5481,N_1623);
xor U6375 (N_6375,N_1091,N_5560);
and U6376 (N_6376,N_3868,N_3625);
xor U6377 (N_6377,N_5709,N_2714);
xnor U6378 (N_6378,N_708,N_1449);
nor U6379 (N_6379,N_5668,N_4811);
xor U6380 (N_6380,N_3569,N_2041);
xnor U6381 (N_6381,N_5050,N_1215);
nand U6382 (N_6382,N_5210,N_49);
nand U6383 (N_6383,N_1426,N_4650);
nand U6384 (N_6384,N_3777,N_495);
and U6385 (N_6385,N_4308,N_5915);
xnor U6386 (N_6386,N_5998,N_96);
and U6387 (N_6387,N_1644,N_5814);
nor U6388 (N_6388,N_4629,N_3308);
xor U6389 (N_6389,N_629,N_4418);
or U6390 (N_6390,N_841,N_5857);
xnor U6391 (N_6391,N_2925,N_582);
nand U6392 (N_6392,N_5979,N_4932);
nor U6393 (N_6393,N_4177,N_1194);
and U6394 (N_6394,N_1872,N_3310);
or U6395 (N_6395,N_765,N_5083);
nand U6396 (N_6396,N_344,N_1235);
nand U6397 (N_6397,N_1518,N_678);
nor U6398 (N_6398,N_508,N_5270);
nand U6399 (N_6399,N_5,N_3469);
and U6400 (N_6400,N_613,N_320);
nor U6401 (N_6401,N_5108,N_4113);
nor U6402 (N_6402,N_132,N_4494);
or U6403 (N_6403,N_2432,N_3971);
and U6404 (N_6404,N_2177,N_3111);
or U6405 (N_6405,N_3575,N_4665);
nand U6406 (N_6406,N_3581,N_5819);
nand U6407 (N_6407,N_84,N_1066);
or U6408 (N_6408,N_5449,N_163);
nor U6409 (N_6409,N_5927,N_2581);
or U6410 (N_6410,N_1803,N_2460);
and U6411 (N_6411,N_1357,N_3888);
and U6412 (N_6412,N_956,N_4472);
nand U6413 (N_6413,N_5920,N_1811);
xnor U6414 (N_6414,N_4586,N_5527);
nand U6415 (N_6415,N_5342,N_1551);
xor U6416 (N_6416,N_5044,N_3474);
xnor U6417 (N_6417,N_3920,N_3590);
nor U6418 (N_6418,N_3901,N_1383);
nor U6419 (N_6419,N_4508,N_1894);
and U6420 (N_6420,N_1621,N_1769);
and U6421 (N_6421,N_5370,N_1245);
xor U6422 (N_6422,N_3160,N_4110);
and U6423 (N_6423,N_3786,N_3002);
and U6424 (N_6424,N_5865,N_5465);
xnor U6425 (N_6425,N_3428,N_4950);
and U6426 (N_6426,N_2970,N_2635);
xor U6427 (N_6427,N_1461,N_298);
xor U6428 (N_6428,N_2501,N_3574);
and U6429 (N_6429,N_332,N_1422);
nor U6430 (N_6430,N_2624,N_2916);
xnor U6431 (N_6431,N_4069,N_2649);
xnor U6432 (N_6432,N_426,N_2910);
nor U6433 (N_6433,N_2045,N_4480);
and U6434 (N_6434,N_2040,N_1600);
or U6435 (N_6435,N_864,N_4800);
and U6436 (N_6436,N_4354,N_941);
nor U6437 (N_6437,N_2774,N_5043);
or U6438 (N_6438,N_3644,N_372);
and U6439 (N_6439,N_3671,N_1988);
nand U6440 (N_6440,N_1294,N_1441);
nor U6441 (N_6441,N_3218,N_1467);
nand U6442 (N_6442,N_1970,N_2796);
and U6443 (N_6443,N_1938,N_4930);
xor U6444 (N_6444,N_207,N_3861);
xnor U6445 (N_6445,N_3822,N_4727);
nand U6446 (N_6446,N_1709,N_4905);
nor U6447 (N_6447,N_1952,N_2962);
nor U6448 (N_6448,N_1423,N_4976);
nor U6449 (N_6449,N_3101,N_3226);
or U6450 (N_6450,N_434,N_4742);
nand U6451 (N_6451,N_3930,N_4316);
nand U6452 (N_6452,N_3651,N_3195);
and U6453 (N_6453,N_4334,N_2867);
nand U6454 (N_6454,N_2360,N_1468);
and U6455 (N_6455,N_1607,N_4524);
nand U6456 (N_6456,N_2266,N_306);
or U6457 (N_6457,N_432,N_37);
nand U6458 (N_6458,N_1851,N_3628);
or U6459 (N_6459,N_1256,N_2129);
nand U6460 (N_6460,N_3852,N_4798);
xnor U6461 (N_6461,N_5659,N_4886);
nand U6462 (N_6462,N_3098,N_4948);
nand U6463 (N_6463,N_4180,N_219);
and U6464 (N_6464,N_4594,N_2848);
nand U6465 (N_6465,N_579,N_663);
xor U6466 (N_6466,N_3999,N_1343);
xor U6467 (N_6467,N_1841,N_926);
or U6468 (N_6468,N_3989,N_3210);
or U6469 (N_6469,N_5625,N_1398);
and U6470 (N_6470,N_4051,N_805);
xor U6471 (N_6471,N_1073,N_4511);
xor U6472 (N_6472,N_5790,N_5117);
and U6473 (N_6473,N_4112,N_2191);
nand U6474 (N_6474,N_2403,N_5055);
nand U6475 (N_6475,N_4801,N_1957);
or U6476 (N_6476,N_5926,N_2879);
and U6477 (N_6477,N_1560,N_2518);
nor U6478 (N_6478,N_2342,N_1257);
or U6479 (N_6479,N_2837,N_3301);
nand U6480 (N_6480,N_2166,N_774);
xor U6481 (N_6481,N_5372,N_81);
and U6482 (N_6482,N_312,N_3802);
or U6483 (N_6483,N_4181,N_2928);
nor U6484 (N_6484,N_691,N_2738);
nor U6485 (N_6485,N_5888,N_5431);
xnor U6486 (N_6486,N_1680,N_3121);
nor U6487 (N_6487,N_3996,N_755);
and U6488 (N_6488,N_5507,N_4002);
nand U6489 (N_6489,N_1479,N_4154);
xor U6490 (N_6490,N_5876,N_1583);
nor U6491 (N_6491,N_645,N_2804);
nand U6492 (N_6492,N_442,N_3457);
nor U6493 (N_6493,N_971,N_4679);
or U6494 (N_6494,N_1593,N_3157);
nand U6495 (N_6495,N_2749,N_2392);
or U6496 (N_6496,N_2070,N_2299);
and U6497 (N_6497,N_172,N_5252);
xor U6498 (N_6498,N_3109,N_3488);
nand U6499 (N_6499,N_5253,N_5231);
nor U6500 (N_6500,N_4141,N_1276);
nor U6501 (N_6501,N_4146,N_4668);
xor U6502 (N_6502,N_3693,N_1395);
nand U6503 (N_6503,N_2669,N_1273);
nand U6504 (N_6504,N_4973,N_1688);
nor U6505 (N_6505,N_5100,N_2504);
nor U6506 (N_6506,N_5164,N_1558);
xor U6507 (N_6507,N_1730,N_1548);
nand U6508 (N_6508,N_3470,N_4132);
xnor U6509 (N_6509,N_676,N_4863);
nor U6510 (N_6510,N_540,N_2851);
xor U6511 (N_6511,N_3990,N_2878);
xnor U6512 (N_6512,N_4691,N_3944);
or U6513 (N_6513,N_4734,N_5520);
xor U6514 (N_6514,N_2983,N_1541);
xnor U6515 (N_6515,N_2797,N_1497);
nor U6516 (N_6516,N_4940,N_4764);
and U6517 (N_6517,N_3265,N_748);
xnor U6518 (N_6518,N_1932,N_1605);
xor U6519 (N_6519,N_989,N_1387);
or U6520 (N_6520,N_3274,N_4900);
or U6521 (N_6521,N_3054,N_5378);
nor U6522 (N_6522,N_3533,N_364);
or U6523 (N_6523,N_5848,N_2477);
nor U6524 (N_6524,N_3443,N_5482);
and U6525 (N_6525,N_4319,N_914);
or U6526 (N_6526,N_4908,N_2441);
and U6527 (N_6527,N_2795,N_2640);
and U6528 (N_6528,N_5243,N_1574);
xnor U6529 (N_6529,N_5047,N_2221);
xor U6530 (N_6530,N_1032,N_3833);
and U6531 (N_6531,N_4558,N_2709);
nor U6532 (N_6532,N_68,N_3911);
nor U6533 (N_6533,N_3231,N_2381);
xor U6534 (N_6534,N_5207,N_280);
xor U6535 (N_6535,N_4504,N_1818);
xor U6536 (N_6536,N_655,N_345);
or U6537 (N_6537,N_186,N_5644);
or U6538 (N_6538,N_4528,N_343);
nor U6539 (N_6539,N_2808,N_5607);
and U6540 (N_6540,N_720,N_2841);
or U6541 (N_6541,N_3629,N_3161);
or U6542 (N_6542,N_363,N_4698);
nand U6543 (N_6543,N_2681,N_1340);
nand U6544 (N_6544,N_5643,N_611);
nand U6545 (N_6545,N_2552,N_182);
and U6546 (N_6546,N_1676,N_5568);
or U6547 (N_6547,N_2077,N_3589);
and U6548 (N_6548,N_5393,N_2974);
and U6549 (N_6549,N_5296,N_3392);
or U6550 (N_6550,N_5828,N_1136);
and U6551 (N_6551,N_1088,N_3515);
and U6552 (N_6552,N_309,N_4193);
or U6553 (N_6553,N_814,N_2260);
nor U6554 (N_6554,N_4272,N_2551);
nor U6555 (N_6555,N_2025,N_4221);
nand U6556 (N_6556,N_5256,N_1755);
nand U6557 (N_6557,N_1191,N_559);
xor U6558 (N_6558,N_3236,N_1691);
or U6559 (N_6559,N_1347,N_4025);
nand U6560 (N_6560,N_634,N_4654);
xnor U6561 (N_6561,N_2762,N_5605);
and U6562 (N_6562,N_4337,N_5025);
nor U6563 (N_6563,N_2011,N_5276);
or U6564 (N_6564,N_1393,N_4794);
and U6565 (N_6565,N_2218,N_4359);
xnor U6566 (N_6566,N_2812,N_7);
nor U6567 (N_6567,N_4300,N_3796);
nand U6568 (N_6568,N_2245,N_2055);
nor U6569 (N_6569,N_4162,N_3724);
nor U6570 (N_6570,N_2354,N_5580);
and U6571 (N_6571,N_1396,N_98);
and U6572 (N_6572,N_3431,N_1063);
xor U6573 (N_6573,N_5407,N_3325);
and U6574 (N_6574,N_5182,N_3981);
nor U6575 (N_6575,N_3343,N_3893);
xnor U6576 (N_6576,N_3547,N_5944);
xnor U6577 (N_6577,N_683,N_588);
and U6578 (N_6578,N_1271,N_3424);
nor U6579 (N_6579,N_541,N_5771);
or U6580 (N_6580,N_2031,N_3924);
and U6581 (N_6581,N_5632,N_1965);
and U6582 (N_6582,N_5034,N_845);
nand U6583 (N_6583,N_2680,N_1266);
nand U6584 (N_6584,N_475,N_430);
nor U6585 (N_6585,N_601,N_177);
and U6586 (N_6586,N_4422,N_5184);
nor U6587 (N_6587,N_3689,N_4575);
nand U6588 (N_6588,N_1984,N_4063);
nand U6589 (N_6589,N_5290,N_284);
xnor U6590 (N_6590,N_2807,N_1089);
nand U6591 (N_6591,N_5171,N_197);
and U6592 (N_6592,N_4055,N_2728);
and U6593 (N_6593,N_3454,N_5614);
nor U6594 (N_6594,N_10,N_5945);
nor U6595 (N_6595,N_3878,N_5596);
and U6596 (N_6596,N_750,N_246);
xnor U6597 (N_6597,N_1062,N_4161);
or U6598 (N_6598,N_27,N_5473);
nor U6599 (N_6599,N_2700,N_620);
and U6600 (N_6600,N_4821,N_2582);
nand U6601 (N_6601,N_273,N_438);
and U6602 (N_6602,N_5155,N_2308);
and U6603 (N_6603,N_4187,N_1139);
or U6604 (N_6604,N_773,N_5722);
and U6605 (N_6605,N_5490,N_770);
or U6606 (N_6606,N_1906,N_1437);
xor U6607 (N_6607,N_3400,N_3234);
and U6608 (N_6608,N_5127,N_3082);
xor U6609 (N_6609,N_3406,N_4190);
and U6610 (N_6610,N_5135,N_516);
xnor U6611 (N_6611,N_3532,N_4395);
xnor U6612 (N_6612,N_5220,N_243);
nor U6613 (N_6613,N_1007,N_2937);
or U6614 (N_6614,N_2010,N_5536);
nand U6615 (N_6615,N_3556,N_4640);
and U6616 (N_6616,N_5145,N_4375);
and U6617 (N_6617,N_347,N_2279);
and U6618 (N_6618,N_5002,N_2695);
nor U6619 (N_6619,N_406,N_4901);
nor U6620 (N_6620,N_5172,N_504);
nor U6621 (N_6621,N_4686,N_4265);
or U6622 (N_6622,N_4630,N_3700);
or U6623 (N_6623,N_5514,N_706);
nor U6624 (N_6624,N_4347,N_1483);
nor U6625 (N_6625,N_4125,N_4139);
or U6626 (N_6626,N_2447,N_3175);
and U6627 (N_6627,N_2269,N_224);
or U6628 (N_6628,N_5254,N_3246);
xnor U6629 (N_6629,N_2301,N_242);
and U6630 (N_6630,N_1832,N_2319);
nand U6631 (N_6631,N_3947,N_4415);
nor U6632 (N_6632,N_311,N_383);
nand U6633 (N_6633,N_109,N_3257);
nor U6634 (N_6634,N_5376,N_5062);
xnor U6635 (N_6635,N_522,N_2502);
nand U6636 (N_6636,N_920,N_5504);
xnor U6637 (N_6637,N_2490,N_1058);
nor U6638 (N_6638,N_2346,N_2671);
nand U6639 (N_6639,N_1741,N_1622);
nand U6640 (N_6640,N_2553,N_5148);
xor U6641 (N_6641,N_5805,N_5080);
nor U6642 (N_6642,N_1478,N_105);
nor U6643 (N_6643,N_3019,N_1164);
xor U6644 (N_6644,N_5078,N_1386);
or U6645 (N_6645,N_902,N_1227);
and U6646 (N_6646,N_5867,N_1305);
or U6647 (N_6647,N_2147,N_2374);
and U6648 (N_6648,N_2226,N_4444);
xor U6649 (N_6649,N_3333,N_1631);
nand U6650 (N_6650,N_162,N_5762);
nor U6651 (N_6651,N_191,N_117);
and U6652 (N_6652,N_592,N_2656);
nor U6653 (N_6653,N_5756,N_1269);
and U6654 (N_6654,N_3052,N_3154);
nor U6655 (N_6655,N_4197,N_5884);
xor U6656 (N_6656,N_5664,N_2250);
or U6657 (N_6657,N_2450,N_851);
xor U6658 (N_6658,N_2398,N_5629);
xnor U6659 (N_6659,N_4917,N_333);
nand U6660 (N_6660,N_3664,N_1039);
xor U6661 (N_6661,N_5636,N_1234);
xor U6662 (N_6662,N_4933,N_3207);
xnor U6663 (N_6663,N_898,N_4555);
nand U6664 (N_6664,N_5031,N_3688);
or U6665 (N_6665,N_855,N_4544);
xor U6666 (N_6666,N_1609,N_1858);
nand U6667 (N_6667,N_4192,N_2466);
and U6668 (N_6668,N_5405,N_2288);
or U6669 (N_6669,N_4548,N_2647);
nand U6670 (N_6670,N_946,N_4244);
and U6671 (N_6671,N_3039,N_2155);
or U6672 (N_6672,N_1094,N_5368);
xnor U6673 (N_6673,N_529,N_5224);
and U6674 (N_6674,N_2135,N_1174);
or U6675 (N_6675,N_464,N_3785);
nor U6676 (N_6676,N_665,N_4921);
or U6677 (N_6677,N_2663,N_4085);
or U6678 (N_6678,N_384,N_4131);
nor U6679 (N_6679,N_5941,N_4844);
xor U6680 (N_6680,N_535,N_4809);
nand U6681 (N_6681,N_3666,N_5816);
or U6682 (N_6682,N_3582,N_4541);
nor U6683 (N_6683,N_3116,N_1247);
nor U6684 (N_6684,N_2715,N_1175);
xnor U6685 (N_6685,N_238,N_2326);
nand U6686 (N_6686,N_4784,N_3997);
and U6687 (N_6687,N_5144,N_894);
xor U6688 (N_6688,N_4947,N_5860);
or U6689 (N_6689,N_2452,N_1944);
xor U6690 (N_6690,N_2404,N_3960);
xor U6691 (N_6691,N_1568,N_2690);
or U6692 (N_6692,N_1410,N_5448);
xnor U6693 (N_6693,N_3201,N_1120);
nand U6694 (N_6694,N_3133,N_5997);
xnor U6695 (N_6695,N_3812,N_1403);
nor U6696 (N_6696,N_1493,N_4432);
nand U6697 (N_6697,N_3374,N_1746);
nor U6698 (N_6698,N_1369,N_5484);
and U6699 (N_6699,N_1902,N_3251);
or U6700 (N_6700,N_747,N_4475);
or U6701 (N_6701,N_1927,N_5248);
nand U6702 (N_6702,N_4023,N_3290);
nor U6703 (N_6703,N_5905,N_1237);
xnor U6704 (N_6704,N_3726,N_4352);
nand U6705 (N_6705,N_3163,N_2820);
xor U6706 (N_6706,N_4611,N_5594);
nor U6707 (N_6707,N_4700,N_151);
nor U6708 (N_6708,N_5146,N_4883);
or U6709 (N_6709,N_5119,N_1689);
nand U6710 (N_6710,N_1487,N_3803);
nor U6711 (N_6711,N_1804,N_1029);
nand U6712 (N_6712,N_4563,N_1124);
or U6713 (N_6713,N_1327,N_1843);
nor U6714 (N_6714,N_4525,N_3919);
nand U6715 (N_6715,N_106,N_2385);
or U6716 (N_6716,N_3148,N_1371);
xnor U6717 (N_6717,N_3991,N_1315);
nor U6718 (N_6718,N_5573,N_3727);
xnor U6719 (N_6719,N_5906,N_2881);
xor U6720 (N_6720,N_4424,N_1190);
nor U6721 (N_6721,N_3490,N_4019);
nor U6722 (N_6722,N_3636,N_3093);
and U6723 (N_6723,N_5020,N_187);
and U6724 (N_6724,N_2819,N_1280);
nor U6725 (N_6725,N_5794,N_1815);
and U6726 (N_6726,N_2924,N_4984);
and U6727 (N_6727,N_2058,N_746);
and U6728 (N_6728,N_119,N_3356);
or U6729 (N_6729,N_4018,N_4041);
xnor U6730 (N_6730,N_5608,N_543);
and U6731 (N_6731,N_1724,N_3702);
nand U6732 (N_6732,N_1131,N_71);
xor U6733 (N_6733,N_3461,N_5921);
nand U6734 (N_6734,N_492,N_1821);
or U6735 (N_6735,N_1599,N_4346);
nor U6736 (N_6736,N_3954,N_1165);
nand U6737 (N_6737,N_3275,N_2331);
xnor U6738 (N_6738,N_2383,N_3513);
xnor U6739 (N_6739,N_2198,N_2028);
or U6740 (N_6740,N_3871,N_848);
nor U6741 (N_6741,N_5557,N_3437);
nor U6742 (N_6742,N_2654,N_5343);
or U6743 (N_6743,N_5606,N_5970);
nand U6744 (N_6744,N_834,N_2462);
or U6745 (N_6745,N_1005,N_3305);
or U6746 (N_6746,N_5255,N_5311);
nor U6747 (N_6747,N_2813,N_4416);
xor U6748 (N_6748,N_1569,N_1056);
or U6749 (N_6749,N_410,N_3269);
xnor U6750 (N_6750,N_3593,N_5239);
or U6751 (N_6751,N_3141,N_2673);
or U6752 (N_6752,N_2118,N_1313);
nand U6753 (N_6753,N_257,N_1533);
xor U6754 (N_6754,N_4878,N_4559);
xnor U6755 (N_6755,N_2237,N_1635);
xnor U6756 (N_6756,N_1968,N_4459);
or U6757 (N_6757,N_250,N_5413);
xor U6758 (N_6758,N_3545,N_4463);
nand U6759 (N_6759,N_3144,N_4922);
nand U6760 (N_6760,N_2020,N_1633);
xnor U6761 (N_6761,N_5558,N_857);
or U6762 (N_6762,N_1382,N_5990);
xnor U6763 (N_6763,N_5735,N_1831);
and U6764 (N_6764,N_3667,N_3353);
xor U6765 (N_6765,N_3912,N_4816);
or U6766 (N_6766,N_1592,N_407);
nand U6767 (N_6767,N_3809,N_5710);
nand U6768 (N_6768,N_2052,N_1998);
xor U6769 (N_6769,N_3907,N_2059);
and U6770 (N_6770,N_2305,N_1793);
and U6771 (N_6771,N_1132,N_1863);
and U6772 (N_6772,N_3639,N_4335);
or U6773 (N_6773,N_536,N_274);
nor U6774 (N_6774,N_1374,N_929);
and U6775 (N_6775,N_5379,N_2991);
xnor U6776 (N_6776,N_5126,N_2101);
or U6777 (N_6777,N_5053,N_4882);
and U6778 (N_6778,N_1966,N_4507);
xor U6779 (N_6779,N_5924,N_1756);
and U6780 (N_6780,N_4230,N_1654);
nor U6781 (N_6781,N_3173,N_2192);
nor U6782 (N_6782,N_5242,N_721);
nor U6783 (N_6783,N_3341,N_4088);
nand U6784 (N_6784,N_2081,N_1767);
xor U6785 (N_6785,N_5380,N_2524);
or U6786 (N_6786,N_550,N_5856);
and U6787 (N_6787,N_357,N_3951);
xor U6788 (N_6788,N_5953,N_4423);
xnor U6789 (N_6789,N_5702,N_2144);
nor U6790 (N_6790,N_3894,N_1640);
nor U6791 (N_6791,N_2195,N_1214);
and U6792 (N_6792,N_76,N_2123);
nor U6793 (N_6793,N_3685,N_5692);
or U6794 (N_6794,N_2194,N_268);
xor U6795 (N_6795,N_4027,N_3439);
nand U6796 (N_6796,N_1158,N_4344);
xnor U6797 (N_6797,N_2604,N_3969);
and U6798 (N_6798,N_4164,N_2735);
nand U6799 (N_6799,N_127,N_5937);
xor U6800 (N_6800,N_619,N_5015);
nand U6801 (N_6801,N_4755,N_2229);
or U6802 (N_6802,N_5262,N_5665);
nand U6803 (N_6803,N_5630,N_291);
or U6804 (N_6804,N_5441,N_5987);
or U6805 (N_6805,N_573,N_4287);
nand U6806 (N_6806,N_628,N_4712);
nor U6807 (N_6807,N_3135,N_3350);
xnor U6808 (N_6808,N_3701,N_1142);
nor U6809 (N_6809,N_3696,N_2903);
or U6810 (N_6810,N_4339,N_1536);
nor U6811 (N_6811,N_1753,N_3014);
or U6812 (N_6812,N_1228,N_874);
or U6813 (N_6813,N_756,N_3458);
xor U6814 (N_6814,N_3959,N_4967);
xor U6815 (N_6815,N_4420,N_3949);
or U6816 (N_6816,N_5197,N_939);
xor U6817 (N_6817,N_1248,N_145);
xor U6818 (N_6818,N_3330,N_4376);
and U6819 (N_6819,N_5488,N_4870);
and U6820 (N_6820,N_5132,N_2292);
nor U6821 (N_6821,N_3865,N_2685);
and U6822 (N_6822,N_5759,N_4050);
and U6823 (N_6823,N_3394,N_1686);
or U6824 (N_6824,N_5459,N_2980);
xnor U6825 (N_6825,N_3015,N_3913);
and U6826 (N_6826,N_4602,N_3782);
nor U6827 (N_6827,N_3046,N_2540);
xor U6828 (N_6828,N_1162,N_3805);
and U6829 (N_6829,N_2127,N_3332);
and U6830 (N_6830,N_2968,N_3020);
and U6831 (N_6831,N_1900,N_4783);
or U6832 (N_6832,N_3447,N_3087);
or U6833 (N_6833,N_2297,N_4851);
nand U6834 (N_6834,N_1213,N_861);
nand U6835 (N_6835,N_967,N_5917);
or U6836 (N_6836,N_465,N_1736);
nor U6837 (N_6837,N_1529,N_693);
and U6838 (N_6838,N_8,N_4033);
nor U6839 (N_6839,N_1264,N_5030);
nor U6840 (N_6840,N_5598,N_3004);
xnor U6841 (N_6841,N_1790,N_5285);
or U6842 (N_6842,N_1346,N_3565);
or U6843 (N_6843,N_2773,N_4046);
xnor U6844 (N_6844,N_22,N_4212);
or U6845 (N_6845,N_5981,N_4099);
nand U6846 (N_6846,N_4171,N_661);
xnor U6847 (N_6847,N_1920,N_2136);
xor U6848 (N_6848,N_480,N_292);
nor U6849 (N_6849,N_1822,N_2658);
nand U6850 (N_6850,N_3277,N_754);
or U6851 (N_6851,N_5548,N_3056);
xnor U6852 (N_6852,N_1370,N_3710);
and U6853 (N_6853,N_589,N_2151);
nor U6854 (N_6854,N_4409,N_4935);
nand U6855 (N_6855,N_5279,N_313);
nand U6856 (N_6856,N_376,N_1030);
or U6857 (N_6857,N_3749,N_1337);
nand U6858 (N_6858,N_780,N_517);
xnor U6859 (N_6859,N_5287,N_3478);
or U6860 (N_6860,N_2203,N_4467);
nor U6861 (N_6861,N_4704,N_790);
and U6862 (N_6862,N_977,N_5295);
nor U6863 (N_6863,N_4834,N_2469);
or U6864 (N_6864,N_3143,N_648);
and U6865 (N_6865,N_3635,N_5367);
nor U6866 (N_6866,N_4350,N_4384);
nand U6867 (N_6867,N_3285,N_1727);
xnor U6868 (N_6868,N_799,N_884);
or U6869 (N_6869,N_3510,N_4981);
nand U6870 (N_6870,N_4329,N_484);
xnor U6871 (N_6871,N_4091,N_4623);
nand U6872 (N_6872,N_1985,N_3873);
and U6873 (N_6873,N_3389,N_5324);
and U6874 (N_6874,N_5371,N_5106);
or U6875 (N_6875,N_981,N_4793);
nand U6876 (N_6876,N_5928,N_3390);
or U6877 (N_6877,N_5859,N_1556);
nand U6878 (N_6878,N_1586,N_3237);
xnor U6879 (N_6879,N_5505,N_2701);
xnor U6880 (N_6880,N_4692,N_5559);
or U6881 (N_6881,N_950,N_3460);
or U6882 (N_6882,N_1415,N_4185);
or U6883 (N_6883,N_3808,N_4578);
and U6884 (N_6884,N_4934,N_846);
xor U6885 (N_6885,N_3783,N_1169);
and U6886 (N_6886,N_3180,N_4299);
nand U6887 (N_6887,N_1949,N_5453);
or U6888 (N_6888,N_5118,N_2002);
nand U6889 (N_6889,N_5313,N_1123);
xor U6890 (N_6890,N_1458,N_5011);
nor U6891 (N_6891,N_4661,N_3849);
and U6892 (N_6892,N_2565,N_28);
xnor U6893 (N_6893,N_5306,N_1525);
nor U6894 (N_6894,N_3945,N_4748);
xor U6895 (N_6895,N_4861,N_4703);
nand U6896 (N_6896,N_3676,N_3193);
nand U6897 (N_6897,N_5180,N_2433);
nor U6898 (N_6898,N_2515,N_5353);
xnor U6899 (N_6899,N_819,N_2688);
xor U6900 (N_6900,N_5697,N_33);
nand U6901 (N_6901,N_1151,N_3441);
and U6902 (N_6902,N_3806,N_4102);
xor U6903 (N_6903,N_391,N_1786);
or U6904 (N_6904,N_4044,N_4505);
or U6905 (N_6905,N_1060,N_1373);
nand U6906 (N_6906,N_2184,N_3770);
and U6907 (N_6907,N_2575,N_4670);
and U6908 (N_6908,N_5988,N_4448);
nand U6909 (N_6909,N_3976,N_3298);
xnor U6910 (N_6910,N_5318,N_932);
and U6911 (N_6911,N_2000,N_2756);
nand U6912 (N_6912,N_1381,N_5736);
or U6913 (N_6913,N_3993,N_3295);
nand U6914 (N_6914,N_4008,N_4868);
and U6915 (N_6915,N_797,N_2092);
or U6916 (N_6916,N_4765,N_474);
xnor U6917 (N_6917,N_4877,N_3970);
nand U6918 (N_6918,N_111,N_374);
nand U6919 (N_6919,N_5792,N_4233);
nor U6920 (N_6920,N_5177,N_5130);
nand U6921 (N_6921,N_2897,N_1931);
or U6922 (N_6922,N_2787,N_1726);
xnor U6923 (N_6923,N_3243,N_5817);
nor U6924 (N_6924,N_4520,N_4842);
or U6925 (N_6925,N_4992,N_2815);
xnor U6926 (N_6926,N_431,N_3254);
xor U6927 (N_6927,N_2069,N_2904);
or U6928 (N_6928,N_5976,N_5916);
nor U6929 (N_6929,N_2416,N_3479);
nand U6930 (N_6930,N_3886,N_19);
and U6931 (N_6931,N_4482,N_514);
xnor U6932 (N_6932,N_4588,N_1773);
nor U6933 (N_6933,N_2706,N_5932);
and U6934 (N_6934,N_1416,N_4247);
xor U6935 (N_6935,N_3232,N_2475);
nor U6936 (N_6936,N_2751,N_428);
nand U6937 (N_6937,N_266,N_4506);
nor U6938 (N_6938,N_4413,N_3641);
and U6939 (N_6939,N_471,N_4919);
nand U6940 (N_6940,N_2523,N_3974);
and U6941 (N_6941,N_2258,N_1647);
or U6942 (N_6942,N_4587,N_1645);
nor U6943 (N_6943,N_299,N_5543);
and U6944 (N_6944,N_179,N_4278);
xnor U6945 (N_6945,N_1552,N_3891);
nor U6946 (N_6946,N_5853,N_3445);
and U6947 (N_6947,N_5713,N_3294);
and U6948 (N_6948,N_5535,N_1002);
nand U6949 (N_6949,N_3213,N_4731);
or U6950 (N_6950,N_4431,N_1001);
xnor U6951 (N_6951,N_282,N_4296);
nand U6952 (N_6952,N_5186,N_1935);
or U6953 (N_6953,N_5124,N_2639);
or U6954 (N_6954,N_788,N_1819);
nand U6955 (N_6955,N_3,N_3619);
or U6956 (N_6956,N_3452,N_3877);
and U6957 (N_6957,N_181,N_5889);
nand U6958 (N_6958,N_1361,N_4360);
and U6959 (N_6959,N_5301,N_5524);
or U6960 (N_6960,N_502,N_4990);
or U6961 (N_6961,N_5811,N_534);
xor U6962 (N_6962,N_3916,N_3652);
or U6963 (N_6963,N_5908,N_2097);
or U6964 (N_6964,N_1896,N_3526);
nor U6965 (N_6965,N_3712,N_1933);
or U6966 (N_6966,N_4092,N_1765);
nor U6967 (N_6967,N_2675,N_3247);
xnor U6968 (N_6968,N_3048,N_5501);
or U6969 (N_6969,N_1895,N_387);
or U6970 (N_6970,N_346,N_4501);
or U6971 (N_6971,N_3863,N_1777);
nand U6972 (N_6972,N_2281,N_3314);
or U6973 (N_6973,N_248,N_1016);
nand U6974 (N_6974,N_2536,N_2038);
or U6975 (N_6975,N_1448,N_3355);
or U6976 (N_6976,N_703,N_4374);
or U6977 (N_6977,N_1823,N_616);
and U6978 (N_6978,N_1099,N_2457);
nor U6979 (N_6979,N_2479,N_4206);
or U6980 (N_6980,N_15,N_1608);
or U6981 (N_6981,N_4167,N_767);
nor U6982 (N_6982,N_3761,N_2684);
xor U6983 (N_6983,N_991,N_2778);
nand U6984 (N_6984,N_4915,N_3453);
nand U6985 (N_6985,N_5509,N_377);
nor U6986 (N_6986,N_5866,N_3206);
and U6987 (N_6987,N_1734,N_5541);
xnor U6988 (N_6988,N_3242,N_4743);
and U6989 (N_6989,N_5634,N_5883);
xnor U6990 (N_6990,N_1206,N_2651);
xnor U6991 (N_6991,N_5707,N_342);
and U6992 (N_6992,N_3691,N_2592);
xnor U6993 (N_6993,N_3631,N_2899);
and U6994 (N_6994,N_4658,N_4037);
nor U6995 (N_6995,N_1384,N_2057);
nand U6996 (N_6996,N_3540,N_3152);
or U6997 (N_6997,N_2366,N_5423);
nand U6998 (N_6998,N_5363,N_1639);
nand U6999 (N_6999,N_3620,N_3303);
nand U7000 (N_7000,N_2016,N_1236);
and U7001 (N_7001,N_5992,N_713);
nand U7002 (N_7002,N_3367,N_775);
and U7003 (N_7003,N_1826,N_4294);
nand U7004 (N_7004,N_5581,N_5549);
nand U7005 (N_7005,N_2614,N_5832);
or U7006 (N_7006,N_3336,N_524);
or U7007 (N_7007,N_5690,N_2660);
xnor U7008 (N_7008,N_1083,N_3740);
nand U7009 (N_7009,N_25,N_3713);
or U7010 (N_7010,N_5375,N_4551);
and U7011 (N_7011,N_300,N_1211);
nand U7012 (N_7012,N_1116,N_1085);
nand U7013 (N_7013,N_5955,N_5475);
and U7014 (N_7014,N_1646,N_5181);
or U7015 (N_7015,N_244,N_2425);
and U7016 (N_7016,N_2541,N_5179);
or U7017 (N_7017,N_2543,N_3695);
and U7018 (N_7018,N_185,N_2397);
or U7019 (N_7019,N_256,N_890);
nor U7020 (N_7020,N_580,N_5683);
and U7021 (N_7021,N_2361,N_3042);
nand U7022 (N_7022,N_5427,N_895);
nand U7023 (N_7023,N_287,N_5283);
nand U7024 (N_7024,N_5892,N_5628);
nand U7025 (N_7025,N_617,N_2984);
nor U7026 (N_7026,N_5486,N_553);
or U7027 (N_7027,N_2233,N_2167);
nand U7028 (N_7028,N_742,N_3649);
nand U7029 (N_7029,N_2933,N_2884);
nor U7030 (N_7030,N_2539,N_3522);
nand U7031 (N_7031,N_1138,N_3472);
and U7032 (N_7032,N_2988,N_4530);
xnor U7033 (N_7033,N_1781,N_2343);
or U7034 (N_7034,N_1615,N_4094);
nand U7035 (N_7035,N_1650,N_1930);
nor U7036 (N_7036,N_133,N_889);
nand U7037 (N_7037,N_3834,N_2969);
nand U7038 (N_7038,N_1290,N_2883);
nor U7039 (N_7039,N_5478,N_451);
nand U7040 (N_7040,N_4671,N_2472);
nor U7041 (N_7041,N_684,N_4684);
nand U7042 (N_7042,N_445,N_1862);
nor U7043 (N_7043,N_551,N_5204);
nor U7044 (N_7044,N_5056,N_4270);
and U7045 (N_7045,N_2476,N_4242);
and U7046 (N_7046,N_1339,N_828);
or U7047 (N_7047,N_4257,N_1719);
or U7048 (N_7048,N_4951,N_3253);
nand U7049 (N_7049,N_1735,N_5728);
and U7050 (N_7050,N_5645,N_1670);
xnor U7051 (N_7051,N_3194,N_2833);
nand U7052 (N_7052,N_759,N_2873);
xor U7053 (N_7053,N_4519,N_1674);
xnor U7054 (N_7054,N_3316,N_3698);
and U7055 (N_7055,N_4393,N_549);
and U7056 (N_7056,N_983,N_4961);
and U7057 (N_7057,N_2717,N_3500);
xnor U7058 (N_7058,N_225,N_2986);
xnor U7059 (N_7059,N_5506,N_5134);
nand U7060 (N_7060,N_1528,N_2781);
nor U7061 (N_7061,N_5656,N_2323);
nor U7062 (N_7062,N_4483,N_1522);
nand U7063 (N_7063,N_4064,N_4836);
and U7064 (N_7064,N_5818,N_4237);
xor U7065 (N_7065,N_1792,N_2800);
or U7066 (N_7066,N_1745,N_3520);
nand U7067 (N_7067,N_3699,N_2113);
or U7068 (N_7068,N_4616,N_2197);
xor U7069 (N_7069,N_3844,N_5374);
xor U7070 (N_7070,N_2672,N_3149);
nand U7071 (N_7071,N_4778,N_1104);
and U7072 (N_7072,N_938,N_1401);
xor U7073 (N_7073,N_4581,N_1702);
nor U7074 (N_7074,N_3432,N_984);
xnor U7075 (N_7075,N_1694,N_2951);
and U7076 (N_7076,N_1150,N_1006);
or U7077 (N_7077,N_4009,N_1003);
nand U7078 (N_7078,N_5396,N_2875);
xnor U7079 (N_7079,N_2265,N_3645);
nand U7080 (N_7080,N_5729,N_4403);
xor U7081 (N_7081,N_3823,N_38);
or U7082 (N_7082,N_3248,N_4470);
xnor U7083 (N_7083,N_2613,N_355);
nor U7084 (N_7084,N_1554,N_1993);
and U7085 (N_7085,N_4398,N_2036);
or U7086 (N_7086,N_5649,N_3708);
nand U7087 (N_7087,N_5304,N_3658);
nor U7088 (N_7088,N_1317,N_2857);
xnor U7089 (N_7089,N_5140,N_12);
xnor U7090 (N_7090,N_5654,N_2451);
nand U7091 (N_7091,N_4182,N_3596);
nor U7092 (N_7092,N_5218,N_5515);
xor U7093 (N_7093,N_1144,N_303);
and U7094 (N_7094,N_5354,N_1928);
nand U7095 (N_7095,N_1742,N_2722);
and U7096 (N_7096,N_1424,N_2303);
or U7097 (N_7097,N_2478,N_964);
nor U7098 (N_7098,N_2246,N_2238);
or U7099 (N_7099,N_4057,N_2156);
nand U7100 (N_7100,N_228,N_761);
xor U7101 (N_7101,N_5989,N_3379);
or U7102 (N_7102,N_2609,N_210);
nand U7103 (N_7103,N_1117,N_1776);
or U7104 (N_7104,N_2494,N_2170);
nor U7105 (N_7105,N_3338,N_5247);
nand U7106 (N_7106,N_4683,N_4610);
or U7107 (N_7107,N_2621,N_5007);
and U7108 (N_7108,N_1080,N_4107);
nand U7109 (N_7109,N_1084,N_2082);
or U7110 (N_7110,N_917,N_3918);
and U7111 (N_7111,N_36,N_1035);
or U7112 (N_7112,N_621,N_3347);
nor U7113 (N_7113,N_1801,N_4752);
nor U7114 (N_7114,N_4956,N_2409);
and U7115 (N_7115,N_86,N_2567);
and U7116 (N_7116,N_5599,N_2561);
and U7117 (N_7117,N_4258,N_4072);
xor U7118 (N_7118,N_5123,N_1126);
and U7119 (N_7119,N_5229,N_2583);
or U7120 (N_7120,N_5178,N_4277);
nand U7121 (N_7121,N_3722,N_1071);
nor U7122 (N_7122,N_5173,N_5154);
nor U7123 (N_7123,N_4907,N_2514);
or U7124 (N_7124,N_590,N_752);
or U7125 (N_7125,N_2091,N_3068);
nand U7126 (N_7126,N_3872,N_3359);
and U7127 (N_7127,N_530,N_2464);
nor U7128 (N_7128,N_1678,N_2661);
nor U7129 (N_7129,N_4290,N_1738);
and U7130 (N_7130,N_2139,N_1708);
and U7131 (N_7131,N_5751,N_3321);
or U7132 (N_7132,N_1816,N_1698);
or U7133 (N_7133,N_3875,N_2730);
and U7134 (N_7134,N_907,N_4385);
nand U7135 (N_7135,N_3729,N_3499);
xor U7136 (N_7136,N_2146,N_5163);
and U7137 (N_7137,N_2949,N_3060);
or U7138 (N_7138,N_3647,N_5570);
or U7139 (N_7139,N_5810,N_5661);
nand U7140 (N_7140,N_3383,N_3450);
nand U7141 (N_7141,N_2033,N_368);
nand U7142 (N_7142,N_4271,N_3309);
or U7143 (N_7143,N_758,N_1289);
xnor U7144 (N_7144,N_4584,N_1642);
or U7145 (N_7145,N_3781,N_262);
xor U7146 (N_7146,N_2678,N_460);
nor U7147 (N_7147,N_2842,N_275);
nand U7148 (N_7148,N_3825,N_4855);
and U7149 (N_7149,N_5674,N_2803);
xor U7150 (N_7150,N_2627,N_2076);
or U7151 (N_7151,N_1618,N_3673);
nor U7152 (N_7152,N_2005,N_4513);
nor U7153 (N_7153,N_2564,N_1682);
nand U7154 (N_7154,N_3754,N_121);
nand U7155 (N_7155,N_5433,N_3853);
nand U7156 (N_7156,N_2901,N_265);
and U7157 (N_7157,N_5734,N_5355);
nand U7158 (N_7158,N_1000,N_4229);
nor U7159 (N_7159,N_921,N_2793);
or U7160 (N_7160,N_4295,N_3342);
nor U7161 (N_7161,N_4013,N_803);
or U7162 (N_7162,N_5101,N_1077);
nor U7163 (N_7163,N_3585,N_4537);
xor U7164 (N_7164,N_509,N_2577);
nor U7165 (N_7165,N_787,N_2825);
and U7166 (N_7166,N_4205,N_1033);
xor U7167 (N_7167,N_4479,N_5384);
nand U7168 (N_7168,N_4942,N_4323);
xor U7169 (N_7169,N_1018,N_5494);
nand U7170 (N_7170,N_5199,N_118);
or U7171 (N_7171,N_1353,N_3646);
and U7172 (N_7172,N_3705,N_3172);
nand U7173 (N_7173,N_4872,N_2080);
and U7174 (N_7174,N_2652,N_173);
nor U7175 (N_7175,N_596,N_3388);
or U7176 (N_7176,N_3876,N_220);
and U7177 (N_7177,N_91,N_2677);
xnor U7178 (N_7178,N_3190,N_3882);
xnor U7179 (N_7179,N_5183,N_5209);
xnor U7180 (N_7180,N_729,N_4941);
nand U7181 (N_7181,N_3063,N_4059);
or U7182 (N_7182,N_5176,N_4298);
xor U7183 (N_7183,N_5369,N_2181);
nor U7184 (N_7184,N_1871,N_4566);
nand U7185 (N_7185,N_2948,N_5483);
xnor U7186 (N_7186,N_5442,N_1453);
nand U7187 (N_7187,N_4147,N_4666);
nor U7188 (N_7188,N_1913,N_2542);
xnor U7189 (N_7189,N_1012,N_3361);
or U7190 (N_7190,N_4808,N_2957);
nand U7191 (N_7191,N_4152,N_3051);
nand U7192 (N_7192,N_4590,N_5238);
nand U7193 (N_7193,N_4095,N_2426);
and U7194 (N_7194,N_2597,N_176);
or U7195 (N_7195,N_2131,N_1665);
nand U7196 (N_7196,N_485,N_2315);
nor U7197 (N_7197,N_5571,N_2347);
xnor U7198 (N_7198,N_4667,N_153);
xor U7199 (N_7199,N_5831,N_5225);
xnor U7200 (N_7200,N_4994,N_3958);
or U7201 (N_7201,N_1967,N_2317);
nand U7202 (N_7202,N_3968,N_381);
or U7203 (N_7203,N_4952,N_4445);
or U7204 (N_7204,N_2048,N_1321);
and U7205 (N_7205,N_4711,N_2225);
nand U7206 (N_7206,N_4677,N_1049);
or U7207 (N_7207,N_211,N_5289);
nor U7208 (N_7208,N_5260,N_5675);
and U7209 (N_7209,N_4526,N_50);
xor U7210 (N_7210,N_1595,N_771);
nand U7211 (N_7211,N_1013,N_511);
nand U7212 (N_7212,N_4910,N_4500);
nor U7213 (N_7213,N_4965,N_673);
and U7214 (N_7214,N_1023,N_4481);
and U7215 (N_7215,N_2588,N_1582);
or U7216 (N_7216,N_2049,N_99);
nor U7217 (N_7217,N_2148,N_2444);
or U7218 (N_7218,N_2391,N_2532);
or U7219 (N_7219,N_1975,N_4343);
nand U7220 (N_7220,N_658,N_4759);
nor U7221 (N_7221,N_3131,N_4892);
nand U7222 (N_7222,N_4963,N_2725);
or U7223 (N_7223,N_1911,N_5440);
xnor U7224 (N_7224,N_633,N_1196);
xor U7225 (N_7225,N_5552,N_5574);
and U7226 (N_7226,N_2446,N_193);
nand U7227 (N_7227,N_1789,N_5995);
nor U7228 (N_7228,N_3255,N_93);
or U7229 (N_7229,N_501,N_2256);
nor U7230 (N_7230,N_4394,N_5156);
or U7231 (N_7231,N_5686,N_4307);
xor U7232 (N_7232,N_5104,N_4318);
nand U7233 (N_7233,N_2159,N_1220);
xnor U7234 (N_7234,N_792,N_4995);
nand U7235 (N_7235,N_3956,N_1855);
xnor U7236 (N_7236,N_1634,N_1209);
nand U7237 (N_7237,N_5138,N_1355);
nor U7238 (N_7238,N_5627,N_302);
nor U7239 (N_7239,N_1992,N_4829);
xor U7240 (N_7240,N_1481,N_2125);
nand U7241 (N_7241,N_1783,N_555);
nand U7242 (N_7242,N_5361,N_3487);
or U7243 (N_7243,N_4406,N_1976);
or U7244 (N_7244,N_1904,N_1352);
xnor U7245 (N_7245,N_1508,N_5566);
or U7246 (N_7246,N_5601,N_821);
nand U7247 (N_7247,N_1017,N_1707);
and U7248 (N_7248,N_473,N_2065);
xnor U7249 (N_7249,N_2362,N_3792);
or U7250 (N_7250,N_4867,N_2596);
or U7251 (N_7251,N_1876,N_3186);
nor U7252 (N_7252,N_1304,N_3217);
or U7253 (N_7253,N_4254,N_1774);
nor U7254 (N_7254,N_677,N_2388);
nor U7255 (N_7255,N_1036,N_2373);
nor U7256 (N_7256,N_5791,N_4410);
and U7257 (N_7257,N_1356,N_696);
or U7258 (N_7258,N_5068,N_4839);
xor U7259 (N_7259,N_2761,N_1649);
xor U7260 (N_7260,N_4657,N_4460);
nand U7261 (N_7261,N_3759,N_650);
nor U7262 (N_7262,N_1156,N_2295);
nor U7263 (N_7263,N_2176,N_4642);
xor U7264 (N_7264,N_3249,N_1394);
or U7265 (N_7265,N_1368,N_2019);
xnor U7266 (N_7266,N_871,N_2336);
or U7267 (N_7267,N_3634,N_1205);
nor U7268 (N_7268,N_5116,N_5693);
nor U7269 (N_7269,N_2758,N_5415);
xnor U7270 (N_7270,N_3033,N_2780);
and U7271 (N_7271,N_2742,N_5359);
nand U7272 (N_7272,N_94,N_3827);
nor U7273 (N_7273,N_3108,N_627);
and U7274 (N_7274,N_911,N_741);
or U7275 (N_7275,N_2790,N_4739);
nand U7276 (N_7276,N_4718,N_5776);
nand U7277 (N_7277,N_5564,N_4010);
and U7278 (N_7278,N_700,N_3606);
and U7279 (N_7279,N_3711,N_123);
and U7280 (N_7280,N_966,N_745);
and U7281 (N_7281,N_3420,N_1986);
nor U7282 (N_7282,N_1641,N_3370);
nor U7283 (N_7283,N_13,N_2966);
nor U7284 (N_7284,N_1808,N_1664);
xor U7285 (N_7285,N_5040,N_258);
nand U7286 (N_7286,N_1572,N_1480);
and U7287 (N_7287,N_3209,N_5610);
xnor U7288 (N_7288,N_5767,N_1281);
and U7289 (N_7289,N_2645,N_1936);
and U7290 (N_7290,N_4517,N_587);
or U7291 (N_7291,N_3998,N_499);
or U7292 (N_7292,N_1748,N_2289);
nand U7293 (N_7293,N_4220,N_4356);
and U7294 (N_7294,N_2753,N_241);
nand U7295 (N_7295,N_4835,N_5546);
xor U7296 (N_7296,N_5667,N_830);
or U7297 (N_7297,N_2068,N_5230);
nand U7298 (N_7298,N_4291,N_1875);
or U7299 (N_7299,N_3718,N_1098);
or U7300 (N_7300,N_1910,N_3964);
or U7301 (N_7301,N_763,N_5967);
nor U7302 (N_7302,N_4061,N_5633);
or U7303 (N_7303,N_3734,N_362);
xor U7304 (N_7304,N_1723,N_307);
nor U7305 (N_7305,N_606,N_3925);
and U7306 (N_7306,N_1977,N_4516);
nor U7307 (N_7307,N_4490,N_5583);
xnor U7308 (N_7308,N_2965,N_5983);
and U7309 (N_7309,N_1462,N_527);
nor U7310 (N_7310,N_4664,N_4632);
nor U7311 (N_7311,N_4435,N_5615);
nand U7312 (N_7312,N_1922,N_4705);
or U7313 (N_7313,N_4633,N_5244);
xnor U7314 (N_7314,N_1223,N_2708);
xnor U7315 (N_7315,N_5797,N_3171);
nor U7316 (N_7316,N_1579,N_2201);
xnor U7317 (N_7317,N_5386,N_20);
and U7318 (N_7318,N_2832,N_3276);
nand U7319 (N_7319,N_2710,N_5175);
or U7320 (N_7320,N_3534,N_3007);
xor U7321 (N_7321,N_1951,N_5966);
xor U7322 (N_7322,N_5167,N_456);
nor U7323 (N_7323,N_180,N_5963);
nand U7324 (N_7324,N_786,N_5931);
xor U7325 (N_7325,N_3531,N_1788);
or U7326 (N_7326,N_1882,N_4341);
and U7327 (N_7327,N_4208,N_3409);
xor U7328 (N_7328,N_1867,N_5059);
nor U7329 (N_7329,N_3386,N_5362);
nand U7330 (N_7330,N_2024,N_2693);
nand U7331 (N_7331,N_4860,N_9);
nand U7332 (N_7332,N_2886,N_1596);
and U7333 (N_7333,N_3731,N_2324);
xnor U7334 (N_7334,N_4645,N_1994);
nand U7335 (N_7335,N_3552,N_4796);
and U7336 (N_7336,N_4970,N_3810);
xor U7337 (N_7337,N_2850,N_2713);
or U7338 (N_7338,N_4327,N_3610);
xor U7339 (N_7339,N_4246,N_3436);
xor U7340 (N_7340,N_1163,N_3289);
xor U7341 (N_7341,N_3337,N_3752);
xor U7342 (N_7342,N_1839,N_92);
nand U7343 (N_7343,N_2798,N_3008);
or U7344 (N_7344,N_1054,N_2183);
nor U7345 (N_7345,N_3509,N_4014);
xnor U7346 (N_7346,N_5715,N_4437);
and U7347 (N_7347,N_1404,N_4378);
or U7348 (N_7348,N_4909,N_3142);
xnor U7349 (N_7349,N_1491,N_990);
and U7350 (N_7350,N_4771,N_1795);
and U7351 (N_7351,N_1177,N_4803);
nor U7352 (N_7352,N_3948,N_2483);
and U7353 (N_7353,N_4231,N_1246);
xor U7354 (N_7354,N_281,N_3661);
and U7355 (N_7355,N_2775,N_5404);
or U7356 (N_7356,N_195,N_2545);
xor U7357 (N_7357,N_3767,N_3842);
nor U7358 (N_7358,N_4111,N_3978);
nand U7359 (N_7359,N_3504,N_3973);
nand U7360 (N_7360,N_5708,N_142);
xnor U7361 (N_7361,N_2549,N_5269);
xor U7362 (N_7362,N_4407,N_1295);
xor U7363 (N_7363,N_5800,N_4888);
nor U7364 (N_7364,N_4730,N_5277);
and U7365 (N_7365,N_1186,N_1109);
or U7366 (N_7366,N_72,N_1761);
xnor U7367 (N_7367,N_1359,N_4622);
and U7368 (N_7368,N_1038,N_215);
or U7369 (N_7369,N_5340,N_4143);
xor U7370 (N_7370,N_3943,N_2572);
nor U7371 (N_7371,N_1961,N_2574);
nand U7372 (N_7372,N_3465,N_1718);
nor U7373 (N_7373,N_2145,N_4135);
nor U7374 (N_7374,N_5678,N_75);
nor U7375 (N_7375,N_796,N_1218);
nor U7376 (N_7376,N_5076,N_2507);
nor U7377 (N_7377,N_1791,N_3660);
or U7378 (N_7378,N_2435,N_5250);
nor U7379 (N_7379,N_2862,N_2401);
nor U7380 (N_7380,N_5094,N_4108);
or U7381 (N_7381,N_4123,N_4292);
or U7382 (N_7382,N_4695,N_2188);
nor U7383 (N_7383,N_5540,N_3442);
or U7384 (N_7384,N_4787,N_1137);
nand U7385 (N_7385,N_3119,N_128);
nand U7386 (N_7386,N_5412,N_5162);
or U7387 (N_7387,N_4715,N_4776);
xor U7388 (N_7388,N_3554,N_3423);
or U7389 (N_7389,N_5746,N_2569);
nor U7390 (N_7390,N_3319,N_3013);
and U7391 (N_7391,N_4462,N_1329);
or U7392 (N_7392,N_794,N_2022);
nand U7393 (N_7393,N_3828,N_3550);
and U7394 (N_7394,N_141,N_4547);
and U7395 (N_7395,N_578,N_29);
and U7396 (N_7396,N_1149,N_3736);
or U7397 (N_7397,N_169,N_2358);
nand U7398 (N_7398,N_839,N_3200);
and U7399 (N_7399,N_3174,N_2495);
nor U7400 (N_7400,N_531,N_863);
and U7401 (N_7401,N_5964,N_2766);
xnor U7402 (N_7402,N_2641,N_4399);
nor U7403 (N_7403,N_3468,N_1476);
and U7404 (N_7404,N_4815,N_2719);
nand U7405 (N_7405,N_1658,N_1258);
or U7406 (N_7406,N_4372,N_657);
xor U7407 (N_7407,N_4652,N_2509);
nor U7408 (N_7408,N_5721,N_1759);
or U7409 (N_7409,N_5165,N_5725);
nand U7410 (N_7410,N_3241,N_283);
and U7411 (N_7411,N_5741,N_1075);
or U7412 (N_7412,N_4160,N_4978);
or U7413 (N_7413,N_3037,N_4846);
xor U7414 (N_7414,N_4213,N_3270);
nand U7415 (N_7415,N_1996,N_670);
or U7416 (N_7416,N_3456,N_2816);
and U7417 (N_7417,N_1559,N_329);
nor U7418 (N_7418,N_2975,N_3922);
and U7419 (N_7419,N_1865,N_2106);
and U7420 (N_7420,N_359,N_1312);
nand U7421 (N_7421,N_5538,N_2075);
nand U7422 (N_7422,N_3721,N_5485);
or U7423 (N_7423,N_2298,N_171);
nor U7424 (N_7424,N_2341,N_5936);
or U7425 (N_7425,N_5893,N_2936);
xor U7426 (N_7426,N_3917,N_487);
xor U7427 (N_7427,N_4791,N_5211);
nand U7428 (N_7428,N_3306,N_1888);
xor U7429 (N_7429,N_801,N_5233);
xor U7430 (N_7430,N_2573,N_3214);
xnor U7431 (N_7431,N_3491,N_4284);
and U7432 (N_7432,N_4364,N_679);
xor U7433 (N_7433,N_1616,N_5803);
or U7434 (N_7434,N_2215,N_4618);
xnor U7435 (N_7435,N_5513,N_4324);
and U7436 (N_7436,N_944,N_1601);
and U7437 (N_7437,N_5572,N_441);
nor U7438 (N_7438,N_5333,N_2599);
nand U7439 (N_7439,N_2440,N_528);
nand U7440 (N_7440,N_2234,N_5221);
nand U7441 (N_7441,N_5553,N_1856);
nand U7442 (N_7442,N_5136,N_47);
nand U7443 (N_7443,N_5411,N_972);
nor U7444 (N_7444,N_3324,N_3393);
or U7445 (N_7445,N_462,N_1550);
xor U7446 (N_7446,N_3859,N_591);
and U7447 (N_7447,N_251,N_5929);
nand U7448 (N_7448,N_4488,N_1580);
or U7449 (N_7449,N_3107,N_5235);
nor U7450 (N_7450,N_4538,N_925);
nor U7451 (N_7451,N_2768,N_3609);
or U7452 (N_7452,N_903,N_2443);
or U7453 (N_7453,N_3259,N_3208);
or U7454 (N_7454,N_1050,N_1561);
nand U7455 (N_7455,N_5088,N_4363);
nand U7456 (N_7456,N_2415,N_5516);
and U7457 (N_7457,N_5621,N_5739);
nand U7458 (N_7458,N_4738,N_3281);
or U7459 (N_7459,N_4194,N_1231);
or U7460 (N_7460,N_4688,N_960);
and U7461 (N_7461,N_2448,N_5201);
and U7462 (N_7462,N_3103,N_3484);
nand U7463 (N_7463,N_3980,N_1543);
or U7464 (N_7464,N_5139,N_1907);
xor U7465 (N_7465,N_2811,N_5510);
nor U7466 (N_7466,N_4795,N_56);
xor U7467 (N_7467,N_4672,N_2286);
and U7468 (N_7468,N_695,N_3928);
or U7469 (N_7469,N_3092,N_3335);
or U7470 (N_7470,N_5849,N_5397);
nor U7471 (N_7471,N_3323,N_3145);
nor U7472 (N_7472,N_1446,N_2168);
or U7473 (N_7473,N_2586,N_5349);
xor U7474 (N_7474,N_5315,N_5406);
nand U7475 (N_7475,N_2021,N_940);
and U7476 (N_7476,N_4142,N_3381);
xor U7477 (N_7477,N_5037,N_3544);
or U7478 (N_7478,N_766,N_3720);
or U7479 (N_7479,N_3223,N_2626);
nor U7480 (N_7480,N_1239,N_3414);
and U7481 (N_7481,N_2294,N_3587);
nor U7482 (N_7482,N_493,N_3790);
or U7483 (N_7483,N_65,N_4227);
nand U7484 (N_7484,N_3123,N_305);
nand U7485 (N_7485,N_1857,N_490);
or U7486 (N_7486,N_3879,N_4);
xor U7487 (N_7487,N_565,N_4613);
and U7488 (N_7488,N_1948,N_853);
or U7489 (N_7489,N_3763,N_2193);
xor U7490 (N_7490,N_1233,N_4939);
or U7491 (N_7491,N_2513,N_533);
nand U7492 (N_7492,N_5292,N_1268);
xor U7493 (N_7493,N_5190,N_3029);
nor U7494 (N_7494,N_5903,N_5684);
or U7495 (N_7495,N_5350,N_548);
and U7496 (N_7496,N_570,N_566);
nand U7497 (N_7497,N_5730,N_2390);
nor U7498 (N_7498,N_568,N_2043);
nor U7499 (N_7499,N_4331,N_640);
and U7500 (N_7500,N_812,N_4653);
nand U7501 (N_7501,N_1732,N_2855);
xor U7502 (N_7502,N_3811,N_2);
or U7503 (N_7503,N_3027,N_2277);
and U7504 (N_7504,N_3963,N_3937);
xor U7505 (N_7505,N_690,N_2116);
xnor U7506 (N_7506,N_1626,N_395);
xor U7507 (N_7507,N_3940,N_1715);
nor U7508 (N_7508,N_1172,N_5899);
xor U7509 (N_7509,N_199,N_170);
nor U7510 (N_7510,N_3025,N_203);
nand U7511 (N_7511,N_4071,N_916);
nor U7512 (N_7512,N_2821,N_2178);
and U7513 (N_7513,N_644,N_1187);
nor U7514 (N_7514,N_3038,N_3614);
or U7515 (N_7515,N_178,N_1199);
nand U7516 (N_7516,N_366,N_2889);
xor U7517 (N_7517,N_5603,N_3102);
nand U7518 (N_7518,N_4159,N_3089);
nor U7519 (N_7519,N_749,N_3527);
xor U7520 (N_7520,N_101,N_1010);
or U7521 (N_7521,N_2089,N_3074);
nor U7522 (N_7522,N_4020,N_3670);
or U7523 (N_7523,N_4320,N_3225);
nor U7524 (N_7524,N_2655,N_987);
xor U7525 (N_7525,N_66,N_3215);
nor U7526 (N_7526,N_2169,N_1443);
nand U7527 (N_7527,N_3136,N_5589);
and U7528 (N_7528,N_3789,N_1869);
xor U7529 (N_7529,N_2268,N_4565);
and U7530 (N_7530,N_5534,N_4920);
nor U7531 (N_7531,N_995,N_5467);
nor U7532 (N_7532,N_5897,N_1320);
nor U7533 (N_7533,N_5555,N_714);
nand U7534 (N_7534,N_494,N_3122);
or U7535 (N_7535,N_301,N_3909);
and U7536 (N_7536,N_5281,N_2117);
or U7537 (N_7537,N_4189,N_4388);
nand U7538 (N_7538,N_3405,N_3164);
and U7539 (N_7539,N_1260,N_697);
nand U7540 (N_7540,N_5084,N_4626);
xor U7541 (N_7541,N_1093,N_5489);
nor U7542 (N_7542,N_4158,N_61);
and U7543 (N_7543,N_560,N_5105);
xnor U7544 (N_7544,N_3296,N_5016);
nor U7545 (N_7545,N_1589,N_1240);
and U7546 (N_7546,N_671,N_779);
or U7547 (N_7547,N_1884,N_3860);
xnor U7548 (N_7548,N_2978,N_4503);
nand U7549 (N_7549,N_2531,N_1721);
nand U7550 (N_7550,N_5750,N_2430);
nor U7551 (N_7551,N_3869,N_1011);
nand U7552 (N_7552,N_4256,N_3403);
and U7553 (N_7553,N_4305,N_707);
or U7554 (N_7554,N_358,N_1243);
and U7555 (N_7555,N_4309,N_5023);
nand U7556 (N_7556,N_4377,N_4266);
nor U7557 (N_7557,N_78,N_915);
xnor U7558 (N_7558,N_4011,N_2449);
nand U7559 (N_7559,N_1717,N_140);
and U7560 (N_7560,N_3322,N_1145);
or U7561 (N_7561,N_4532,N_662);
or U7562 (N_7562,N_5408,N_146);
and U7563 (N_7563,N_5309,N_5346);
nor U7564 (N_7564,N_4880,N_1625);
nor U7565 (N_7565,N_686,N_5337);
xor U7566 (N_7566,N_1969,N_1797);
xnor U7567 (N_7567,N_2402,N_4259);
xnor U7568 (N_7568,N_2200,N_585);
or U7569 (N_7569,N_4015,N_2662);
xnor U7570 (N_7570,N_294,N_5823);
nor U7571 (N_7571,N_4572,N_3273);
and U7572 (N_7572,N_1272,N_985);
nand U7573 (N_7573,N_3591,N_5003);
xnor U7574 (N_7574,N_1713,N_3915);
and U7575 (N_7575,N_4155,N_3150);
xnor U7576 (N_7576,N_4179,N_5948);
xor U7577 (N_7577,N_4103,N_3010);
nor U7578 (N_7578,N_3090,N_4425);
and U7579 (N_7579,N_4301,N_3222);
and U7580 (N_7580,N_5214,N_4082);
and U7581 (N_7581,N_5882,N_5822);
and U7582 (N_7582,N_2384,N_1805);
nor U7583 (N_7583,N_5064,N_2880);
nor U7584 (N_7584,N_4871,N_5500);
and U7585 (N_7585,N_1322,N_4773);
or U7586 (N_7586,N_1330,N_397);
or U7587 (N_7587,N_1566,N_154);
xor U7588 (N_7588,N_5241,N_3023);
nand U7589 (N_7589,N_420,N_2750);
xor U7590 (N_7590,N_5251,N_4042);
or U7591 (N_7591,N_885,N_5345);
nand U7592 (N_7592,N_2694,N_545);
or U7593 (N_7593,N_3012,N_5261);
nor U7594 (N_7594,N_3753,N_1081);
nor U7595 (N_7595,N_369,N_2940);
nor U7596 (N_7596,N_21,N_3934);
nor U7597 (N_7597,N_4603,N_4549);
nor U7598 (N_7598,N_2861,N_1555);
nor U7599 (N_7599,N_4574,N_2006);
nand U7600 (N_7600,N_1842,N_1954);
nand U7601 (N_7601,N_4405,N_3529);
nand U7602 (N_7602,N_5809,N_1250);
nand U7603 (N_7603,N_5322,N_4105);
and U7604 (N_7604,N_4186,N_4962);
and U7605 (N_7605,N_2418,N_5738);
and U7606 (N_7606,N_4355,N_4251);
xnor U7607 (N_7607,N_1710,N_3088);
and U7608 (N_7608,N_3395,N_5626);
nor U7609 (N_7609,N_3675,N_500);
nor U7610 (N_7610,N_3714,N_4191);
nor U7611 (N_7611,N_5874,N_3035);
and U7612 (N_7612,N_2836,N_2570);
nor U7613 (N_7613,N_2484,N_5508);
or U7614 (N_7614,N_5620,N_5747);
xnor U7615 (N_7615,N_5789,N_4196);
nor U7616 (N_7616,N_1064,N_3816);
and U7617 (N_7617,N_2413,N_77);
nor U7618 (N_7618,N_5419,N_3772);
nor U7619 (N_7619,N_1704,N_778);
xnor U7620 (N_7620,N_402,N_2739);
xnor U7621 (N_7621,N_4195,N_1402);
xor U7622 (N_7622,N_2727,N_4281);
and U7623 (N_7623,N_5807,N_5018);
nor U7624 (N_7624,N_1463,N_3730);
or U7625 (N_7625,N_2698,N_2109);
nor U7626 (N_7626,N_4810,N_2616);
or U7627 (N_7627,N_125,N_2163);
nor U7628 (N_7628,N_5781,N_4279);
or U7629 (N_7629,N_5128,N_4770);
and U7630 (N_7630,N_815,N_5855);
nor U7631 (N_7631,N_724,N_5940);
xor U7632 (N_7632,N_4362,N_3952);
or U7633 (N_7633,N_1926,N_5778);
nand U7634 (N_7634,N_3360,N_4843);
and U7635 (N_7635,N_1118,N_3159);
nand U7636 (N_7636,N_337,N_2095);
and U7637 (N_7637,N_324,N_1425);
nor U7638 (N_7638,N_4223,N_2209);
or U7639 (N_7639,N_4926,N_2262);
or U7640 (N_7640,N_5720,N_164);
xnor U7641 (N_7641,N_5802,N_4789);
nor U7642 (N_7642,N_3284,N_1833);
and U7643 (N_7643,N_3016,N_4165);
or U7644 (N_7644,N_2921,N_897);
xor U7645 (N_7645,N_4515,N_3140);
and U7646 (N_7646,N_4173,N_5373);
or U7647 (N_7647,N_3570,N_5060);
and U7648 (N_7648,N_5595,N_3080);
and U7649 (N_7649,N_1292,N_2945);
and U7650 (N_7650,N_1847,N_390);
or U7651 (N_7651,N_4659,N_2528);
and U7652 (N_7652,N_2785,N_1189);
nand U7653 (N_7653,N_1358,N_1291);
nor U7654 (N_7654,N_4869,N_1799);
xor U7655 (N_7655,N_1323,N_1242);
nand U7656 (N_7656,N_694,N_1806);
and U7657 (N_7657,N_3768,N_1311);
and U7658 (N_7658,N_3205,N_4411);
xor U7659 (N_7659,N_785,N_4336);
and U7660 (N_7660,N_992,N_4214);
or U7661 (N_7661,N_3099,N_1565);
and U7662 (N_7662,N_3655,N_3266);
or U7663 (N_7663,N_4561,N_5717);
xnor U7664 (N_7664,N_3057,N_5813);
xnor U7665 (N_7665,N_5743,N_3352);
or U7666 (N_7666,N_820,N_1879);
nor U7667 (N_7667,N_4120,N_4440);
and U7668 (N_7668,N_3523,N_3475);
nand U7669 (N_7669,N_5232,N_385);
nor U7670 (N_7670,N_2230,N_2799);
nand U7671 (N_7671,N_1046,N_598);
and U7672 (N_7672,N_26,N_5925);
xor U7673 (N_7673,N_5310,N_1850);
or U7674 (N_7674,N_1499,N_4720);
nand U7675 (N_7675,N_2707,N_593);
xor U7676 (N_7676,N_5672,N_1814);
or U7677 (N_7677,N_5900,N_781);
or U7678 (N_7678,N_4466,N_1309);
and U7679 (N_7679,N_3501,N_5472);
nor U7680 (N_7680,N_5463,N_1515);
and U7681 (N_7681,N_4732,N_5646);
and U7682 (N_7682,N_2207,N_806);
or U7683 (N_7683,N_5435,N_2891);
nand U7684 (N_7684,N_3553,N_4328);
nor U7685 (N_7685,N_3369,N_860);
xnor U7686 (N_7686,N_1284,N_235);
xor U7687 (N_7687,N_3577,N_928);
nor U7688 (N_7688,N_3611,N_3817);
nor U7689 (N_7689,N_1100,N_615);
or U7690 (N_7690,N_5497,N_2141);
and U7691 (N_7691,N_31,N_44);
nand U7692 (N_7692,N_1629,N_577);
or U7693 (N_7693,N_354,N_2379);
xor U7694 (N_7694,N_583,N_722);
and U7695 (N_7695,N_5021,N_731);
xnor U7696 (N_7696,N_3422,N_2126);
or U7697 (N_7697,N_5079,N_4736);
nand U7698 (N_7698,N_2789,N_2792);
and U7699 (N_7699,N_1553,N_862);
or U7700 (N_7700,N_174,N_3538);
nand U7701 (N_7701,N_1009,N_1990);
or U7702 (N_7702,N_339,N_2767);
nor U7703 (N_7703,N_2757,N_3315);
and U7704 (N_7704,N_232,N_2034);
nand U7705 (N_7705,N_5327,N_892);
nand U7706 (N_7706,N_3600,N_1893);
nor U7707 (N_7707,N_5592,N_5445);
or U7708 (N_7708,N_733,N_4006);
nor U7709 (N_7709,N_1602,N_3933);
nor U7710 (N_7710,N_213,N_1286);
nand U7711 (N_7711,N_3723,N_4404);
xor U7712 (N_7712,N_3984,N_5271);
nand U7713 (N_7713,N_4635,N_3787);
and U7714 (N_7714,N_4567,N_5798);
or U7715 (N_7715,N_2650,N_2365);
or U7716 (N_7716,N_3979,N_1212);
xnor U7717 (N_7717,N_2060,N_3613);
and U7718 (N_7718,N_866,N_1168);
or U7719 (N_7719,N_2102,N_4262);
nand U7720 (N_7720,N_5687,N_1106);
xor U7721 (N_7721,N_467,N_3181);
nand U7722 (N_7722,N_340,N_209);
nor U7723 (N_7723,N_698,N_3384);
or U7724 (N_7724,N_4476,N_1203);
xor U7725 (N_7725,N_1846,N_4255);
or U7726 (N_7726,N_3349,N_3794);
or U7727 (N_7727,N_564,N_5460);
xor U7728 (N_7728,N_4813,N_5352);
xnor U7729 (N_7729,N_2224,N_5840);
nor U7730 (N_7730,N_1241,N_5575);
or U7731 (N_7731,N_5773,N_2791);
nand U7732 (N_7732,N_2417,N_850);
and U7733 (N_7733,N_3516,N_1472);
nor U7734 (N_7734,N_743,N_288);
nor U7735 (N_7735,N_2283,N_5216);
xor U7736 (N_7736,N_5385,N_408);
xnor U7737 (N_7737,N_5149,N_2827);
and U7738 (N_7738,N_4606,N_3339);
and U7739 (N_7739,N_4540,N_2871);
and U7740 (N_7740,N_4118,N_2754);
nor U7741 (N_7741,N_1766,N_3495);
nor U7742 (N_7742,N_4218,N_804);
and U7743 (N_7743,N_2482,N_4453);
nor U7744 (N_7744,N_1700,N_5045);
nor U7745 (N_7745,N_730,N_4419);
or U7746 (N_7746,N_1714,N_5319);
nor U7747 (N_7747,N_5820,N_4709);
xnor U7748 (N_7748,N_3261,N_4387);
and U7749 (N_7749,N_4958,N_3287);
xnor U7750 (N_7750,N_2247,N_4971);
xor U7751 (N_7751,N_5339,N_270);
xnor U7752 (N_7752,N_1421,N_808);
and U7753 (N_7753,N_649,N_3883);
or U7754 (N_7754,N_1812,N_4455);
nand U7755 (N_7755,N_126,N_3502);
nand U7756 (N_7756,N_4004,N_2979);
and U7757 (N_7757,N_3233,N_5240);
or U7758 (N_7758,N_5487,N_3049);
xor U7759 (N_7759,N_437,N_968);
and U7760 (N_7760,N_1184,N_3858);
or U7761 (N_7761,N_904,N_1119);
or U7762 (N_7762,N_2438,N_3346);
nor U7763 (N_7763,N_360,N_5933);
nor U7764 (N_7764,N_2771,N_2960);
and U7765 (N_7765,N_5205,N_3449);
xor U7766 (N_7766,N_4655,N_1377);
or U7767 (N_7767,N_2222,N_4441);
or U7768 (N_7768,N_5768,N_497);
xor U7769 (N_7769,N_1153,N_1274);
xor U7770 (N_7770,N_4414,N_5985);
or U7771 (N_7771,N_261,N_5511);
xor U7772 (N_7772,N_144,N_35);
and U7773 (N_7773,N_586,N_2644);
and U7774 (N_7774,N_769,N_231);
or U7775 (N_7775,N_5203,N_4029);
and U7776 (N_7776,N_2869,N_3375);
nand U7777 (N_7777,N_1632,N_3535);
and U7778 (N_7778,N_2270,N_3366);
nand U7779 (N_7779,N_3605,N_5133);
or U7780 (N_7780,N_4264,N_1473);
and U7781 (N_7781,N_2611,N_3542);
nand U7782 (N_7782,N_4209,N_1701);
or U7783 (N_7783,N_2185,N_3961);
xnor U7784 (N_7784,N_2682,N_5360);
nor U7785 (N_7785,N_389,N_4777);
or U7786 (N_7786,N_744,N_2794);
and U7787 (N_7787,N_3448,N_1447);
and U7788 (N_7788,N_1613,N_4115);
nor U7789 (N_7789,N_3077,N_5565);
nand U7790 (N_7790,N_3440,N_4078);
and U7791 (N_7791,N_1779,N_2271);
or U7792 (N_7792,N_3774,N_2558);
nand U7793 (N_7793,N_5670,N_3895);
xnor U7794 (N_7794,N_600,N_4891);
and U7795 (N_7795,N_24,N_5479);
nand U7796 (N_7796,N_296,N_2987);
and U7797 (N_7797,N_4542,N_3592);
and U7798 (N_7798,N_635,N_5249);
nand U7799 (N_7799,N_3942,N_3139);
nand U7800 (N_7800,N_3854,N_147);
nor U7801 (N_7801,N_5652,N_5121);
nor U7802 (N_7802,N_3836,N_2926);
xor U7803 (N_7803,N_4966,N_3932);
or U7804 (N_7804,N_2977,N_2400);
xor U7805 (N_7805,N_2481,N_1859);
nor U7806 (N_7806,N_873,N_2263);
or U7807 (N_7807,N_1537,N_5258);
and U7808 (N_7808,N_3179,N_5780);
nand U7809 (N_7809,N_1414,N_3053);
xnor U7810 (N_7810,N_5977,N_4576);
nand U7811 (N_7811,N_350,N_5999);
nand U7812 (N_7812,N_4852,N_5518);
or U7813 (N_7813,N_2264,N_1627);
xor U7814 (N_7814,N_3117,N_3507);
nor U7815 (N_7815,N_2526,N_5208);
xnor U7816 (N_7816,N_5143,N_1436);
nor U7817 (N_7817,N_4216,N_2580);
xnor U7818 (N_7818,N_1412,N_4685);
nand U7819 (N_7819,N_2562,N_5760);
xnor U7820 (N_7820,N_1070,N_3659);
xnor U7821 (N_7821,N_4946,N_5660);
or U7822 (N_7822,N_2304,N_3573);
or U7823 (N_7823,N_205,N_1042);
or U7824 (N_7824,N_4040,N_3156);
xnor U7825 (N_7825,N_2171,N_5115);
xnor U7826 (N_7826,N_315,N_4321);
or U7827 (N_7827,N_4600,N_4601);
nor U7828 (N_7828,N_3096,N_1510);
nor U7829 (N_7829,N_4369,N_3650);
and U7830 (N_7830,N_2412,N_4562);
nor U7831 (N_7831,N_3489,N_2952);
xor U7832 (N_7832,N_5698,N_3418);
or U7833 (N_7833,N_349,N_4067);
and U7834 (N_7834,N_2293,N_5845);
nand U7835 (N_7835,N_5089,N_5703);
nor U7836 (N_7836,N_3061,N_1506);
or U7837 (N_7837,N_5526,N_3421);
xnor U7838 (N_7838,N_4849,N_5640);
nand U7839 (N_7839,N_396,N_5302);
nand U7840 (N_7840,N_4938,N_503);
nand U7841 (N_7841,N_4766,N_1498);
and U7842 (N_7842,N_3021,N_4026);
and U7843 (N_7843,N_4779,N_3755);
nand U7844 (N_7844,N_3153,N_4268);
xnor U7845 (N_7845,N_2885,N_4175);
or U7846 (N_7846,N_2852,N_561);
or U7847 (N_7847,N_2212,N_416);
nor U7848 (N_7848,N_5305,N_2763);
or U7849 (N_7849,N_1277,N_43);
xor U7850 (N_7850,N_5868,N_5410);
and U7851 (N_7851,N_5096,N_3758);
or U7852 (N_7852,N_1364,N_3764);
or U7853 (N_7853,N_1166,N_3906);
nand U7854 (N_7854,N_5328,N_1785);
nand U7855 (N_7855,N_382,N_1301);
xnor U7856 (N_7856,N_5057,N_1545);
and U7857 (N_7857,N_1041,N_1887);
nor U7858 (N_7858,N_1338,N_1652);
and U7859 (N_7859,N_5871,N_2930);
xnor U7860 (N_7860,N_2350,N_2130);
and U7861 (N_7861,N_4465,N_3183);
and U7862 (N_7862,N_353,N_945);
and U7863 (N_7863,N_1659,N_5409);
nor U7864 (N_7864,N_1464,N_411);
and U7865 (N_7865,N_3633,N_4391);
and U7866 (N_7866,N_3219,N_352);
nand U7867 (N_7867,N_3557,N_3382);
xnor U7868 (N_7868,N_5954,N_2474);
xor U7869 (N_7869,N_2320,N_1024);
and U7870 (N_7870,N_2257,N_2073);
xnor U7871 (N_7871,N_1591,N_2824);
and U7872 (N_7872,N_4817,N_2670);
nand U7873 (N_7873,N_1097,N_254);
nor U7874 (N_7874,N_4893,N_562);
and U7875 (N_7875,N_2629,N_827);
nor U7876 (N_7876,N_4556,N_3684);
xnor U7877 (N_7877,N_334,N_2150);
or U7878 (N_7878,N_2339,N_3434);
nor U7879 (N_7879,N_4390,N_3746);
nand U7880 (N_7880,N_4521,N_5320);
or U7881 (N_7881,N_1962,N_5597);
or U7882 (N_7882,N_1411,N_3073);
and U7883 (N_7883,N_4049,N_4707);
nand U7884 (N_7884,N_373,N_236);
and U7885 (N_7885,N_1813,N_5877);
nor U7886 (N_7886,N_5312,N_4697);
nor U7887 (N_7887,N_4820,N_4913);
and U7888 (N_7888,N_1431,N_4681);
nand U7889 (N_7889,N_5471,N_175);
xor U7890 (N_7890,N_5338,N_4275);
or U7891 (N_7891,N_2726,N_1022);
and U7892 (N_7892,N_2872,N_882);
nor U7893 (N_7893,N_1898,N_4977);
nand U7894 (N_7894,N_3881,N_2487);
xnor U7895 (N_7895,N_1924,N_289);
xor U7896 (N_7896,N_5298,N_2584);
nor U7897 (N_7897,N_4172,N_1668);
xor U7898 (N_7898,N_4097,N_5706);
nand U7899 (N_7899,N_5008,N_2630);
nor U7900 (N_7900,N_2202,N_1185);
nor U7901 (N_7901,N_789,N_1044);
or U7902 (N_7902,N_3410,N_3814);
or U7903 (N_7903,N_1861,N_532);
xor U7904 (N_7904,N_5019,N_4687);
nor U7905 (N_7905,N_4646,N_2160);
and U7906 (N_7906,N_1200,N_5677);
or U7907 (N_7907,N_5585,N_1562);
and U7908 (N_7908,N_5830,N_483);
nor U7909 (N_7909,N_738,N_2332);
nand U7910 (N_7910,N_4582,N_2915);
or U7911 (N_7911,N_5958,N_130);
and U7912 (N_7912,N_3638,N_4126);
or U7913 (N_7913,N_3756,N_4454);
or U7914 (N_7914,N_1332,N_1864);
nand U7915 (N_7915,N_1817,N_5073);
or U7916 (N_7916,N_82,N_982);
xnor U7917 (N_7917,N_831,N_3856);
nor U7918 (N_7918,N_5752,N_2486);
or U7919 (N_7919,N_5719,N_2705);
nor U7920 (N_7920,N_1514,N_3624);
and U7921 (N_7921,N_1941,N_3059);
or U7922 (N_7922,N_948,N_486);
xnor U7923 (N_7923,N_3617,N_1263);
xor U7924 (N_7924,N_5584,N_3704);
and U7925 (N_7925,N_1772,N_4285);
xor U7926 (N_7926,N_2835,N_1883);
nor U7927 (N_7927,N_5038,N_705);
xor U7928 (N_7928,N_5895,N_4274);
xor U7929 (N_7929,N_4760,N_5563);
and U7930 (N_7930,N_1095,N_2689);
and U7931 (N_7931,N_4303,N_996);
or U7932 (N_7932,N_1160,N_4724);
xor U7933 (N_7933,N_1844,N_1737);
or U7934 (N_7934,N_1259,N_4116);
nor U7935 (N_7935,N_1045,N_3062);
or U7936 (N_7936,N_5192,N_3045);
and U7937 (N_7937,N_3097,N_5429);
xor U7938 (N_7938,N_1086,N_1983);
nor U7939 (N_7939,N_664,N_1179);
nor U7940 (N_7940,N_3094,N_3815);
nand U7941 (N_7941,N_3348,N_1465);
xor U7942 (N_7942,N_5701,N_4899);
and U7943 (N_7943,N_3560,N_4837);
nand U7944 (N_7944,N_4857,N_3715);
nand U7945 (N_7945,N_3066,N_4349);
nor U7946 (N_7946,N_5962,N_1606);
nand U7947 (N_7947,N_681,N_1796);
xnor U7948 (N_7948,N_5129,N_3686);
xor U7949 (N_7949,N_2329,N_5851);
nor U7950 (N_7950,N_1527,N_4799);
and U7951 (N_7951,N_2783,N_4293);
or U7952 (N_7952,N_4130,N_4756);
nand U7953 (N_7953,N_625,N_3044);
nand U7954 (N_7954,N_249,N_1107);
or U7955 (N_7955,N_1603,N_1178);
and U7956 (N_7956,N_2585,N_1389);
nor U7957 (N_7957,N_3604,N_3864);
xor U7958 (N_7958,N_198,N_1278);
and U7959 (N_7959,N_1725,N_5081);
or U7960 (N_7960,N_3583,N_3832);
nor U7961 (N_7961,N_5984,N_768);
nor U7962 (N_7962,N_2997,N_3798);
xor U7963 (N_7963,N_5151,N_4531);
xnor U7964 (N_7964,N_4436,N_2993);
or U7965 (N_7965,N_3561,N_3239);
xor U7966 (N_7966,N_1729,N_2755);
xor U7967 (N_7967,N_4151,N_2368);
and U7968 (N_7968,N_5228,N_3733);
and U7969 (N_7969,N_2142,N_692);
nor U7970 (N_7970,N_3318,N_1221);
nand U7971 (N_7971,N_4585,N_3112);
nor U7972 (N_7972,N_102,N_4080);
and U7973 (N_7973,N_1201,N_5215);
and U7974 (N_7974,N_5217,N_4560);
and U7975 (N_7975,N_2325,N_1667);
and U7976 (N_7976,N_3471,N_4812);
and U7977 (N_7977,N_4056,N_3669);
nand U7978 (N_7978,N_5194,N_5808);
or U7979 (N_7979,N_4927,N_1891);
nand U7980 (N_7980,N_5266,N_906);
nor U7981 (N_7981,N_3009,N_1655);
or U7982 (N_7982,N_1945,N_2544);
nand U7983 (N_7983,N_5918,N_4314);
nand U7984 (N_7984,N_3926,N_682);
nand U7985 (N_7985,N_1693,N_3070);
and U7986 (N_7986,N_2657,N_1110);
nor U7987 (N_7987,N_4827,N_896);
and U7988 (N_7988,N_4641,N_3548);
or U7989 (N_7989,N_1076,N_4232);
or U7990 (N_7990,N_1501,N_2510);
xor U7991 (N_7991,N_3769,N_1432);
nor U7992 (N_7992,N_481,N_1026);
nand U7993 (N_7993,N_2818,N_1567);
nand U7994 (N_7994,N_5617,N_5994);
xnor U7995 (N_7995,N_727,N_507);
and U7996 (N_7996,N_5754,N_5838);
nand U7997 (N_7997,N_1255,N_5650);
nand U7998 (N_7998,N_4451,N_2074);
and U7999 (N_7999,N_1751,N_30);
or U8000 (N_8000,N_2923,N_4249);
or U8001 (N_8001,N_4138,N_3818);
and U8002 (N_8002,N_2140,N_2946);
nand U8003 (N_8003,N_3184,N_5444);
nor U8004 (N_8004,N_2071,N_5934);
and U8005 (N_8005,N_636,N_1219);
nor U8006 (N_8006,N_4484,N_3297);
xnor U8007 (N_8007,N_468,N_5432);
nor U8008 (N_8008,N_5689,N_735);
and U8009 (N_8009,N_1934,N_2153);
and U8010 (N_8010,N_4034,N_1025);
and U8011 (N_8011,N_1275,N_2003);
or U8012 (N_8012,N_2723,N_2344);
or U8013 (N_8013,N_1912,N_4797);
and U8014 (N_8014,N_2274,N_80);
nand U8015 (N_8015,N_4198,N_4914);
nor U8016 (N_8016,N_1254,N_3189);
nand U8017 (N_8017,N_3067,N_1991);
xnor U8018 (N_8018,N_4073,N_1614);
and U8019 (N_8019,N_2888,N_3679);
and U8020 (N_8020,N_3536,N_2863);
or U8021 (N_8021,N_3884,N_4889);
and U8022 (N_8022,N_1577,N_870);
nor U8023 (N_8023,N_3084,N_726);
nor U8024 (N_8024,N_4226,N_5935);
nor U8025 (N_8025,N_2530,N_4121);
and U8026 (N_8026,N_5293,N_2208);
and U8027 (N_8027,N_3987,N_3887);
xor U8028 (N_8028,N_247,N_4074);
nor U8029 (N_8029,N_3962,N_5969);
or U8030 (N_8030,N_4219,N_4580);
and U8031 (N_8031,N_190,N_515);
xor U8032 (N_8032,N_1456,N_1040);
or U8033 (N_8033,N_2306,N_4782);
and U8034 (N_8034,N_4383,N_4573);
nor U8035 (N_8035,N_2860,N_4053);
and U8036 (N_8036,N_46,N_5854);
nand U8037 (N_8037,N_3965,N_1890);
nor U8038 (N_8038,N_5416,N_4522);
xor U8039 (N_8039,N_5846,N_2369);
or U8040 (N_8040,N_659,N_2115);
nor U8041 (N_8041,N_4153,N_2213);
nand U8042 (N_8042,N_5785,N_5336);
and U8043 (N_8043,N_4802,N_3988);
nor U8044 (N_8044,N_3576,N_4427);
or U8045 (N_8045,N_1651,N_680);
nor U8046 (N_8046,N_1310,N_158);
nand U8047 (N_8047,N_1438,N_5639);
nor U8048 (N_8048,N_4332,N_4371);
nor U8049 (N_8049,N_2340,N_1048);
and U8050 (N_8050,N_4597,N_0);
xnor U8051 (N_8051,N_5436,N_3034);
or U8052 (N_8052,N_5914,N_3518);
xnor U8053 (N_8053,N_223,N_3820);
nand U8054 (N_8054,N_4163,N_4450);
and U8055 (N_8055,N_5673,N_1252);
nor U8056 (N_8056,N_974,N_4996);
nor U8057 (N_8057,N_2914,N_2023);
xor U8058 (N_8058,N_277,N_725);
or U8059 (N_8059,N_4733,N_2152);
or U8060 (N_8060,N_1564,N_3368);
xnor U8061 (N_8061,N_5875,N_3391);
xnor U8062 (N_8062,N_3824,N_479);
nor U8063 (N_8063,N_2377,N_5029);
nand U8064 (N_8064,N_4243,N_1141);
nor U8065 (N_8065,N_5539,N_2535);
nand U8066 (N_8066,N_739,N_936);
nand U8067 (N_8067,N_5980,N_2900);
xnor U8068 (N_8068,N_5090,N_5388);
nand U8069 (N_8069,N_859,N_1695);
nand U8070 (N_8070,N_783,N_1146);
nand U8071 (N_8071,N_1974,N_688);
xnor U8072 (N_8072,N_986,N_1457);
nand U8073 (N_8073,N_1516,N_2066);
nor U8074 (N_8074,N_4592,N_736);
xor U8075 (N_8075,N_2030,N_3568);
xnor U8076 (N_8076,N_4117,N_829);
xor U8077 (N_8077,N_5114,N_4819);
nor U8078 (N_8078,N_4024,N_2012);
and U8079 (N_8079,N_3599,N_1749);
or U8080 (N_8080,N_5956,N_3838);
nor U8081 (N_8081,N_2603,N_3079);
and U8082 (N_8082,N_4128,N_1208);
and U8083 (N_8083,N_5246,N_4786);
xnor U8084 (N_8084,N_2046,N_2998);
xnor U8085 (N_8085,N_5272,N_883);
and U8086 (N_8086,N_1666,N_1392);
nor U8087 (N_8087,N_2096,N_1108);
xor U8088 (N_8088,N_5691,N_3889);
xnor U8089 (N_8089,N_1997,N_5907);
nand U8090 (N_8090,N_3897,N_5006);
nor U8091 (N_8091,N_5826,N_3485);
nand U8092 (N_8092,N_4048,N_2104);
and U8093 (N_8093,N_852,N_1960);
xnor U8094 (N_8094,N_2098,N_2721);
nor U8095 (N_8095,N_1820,N_610);
nand U8096 (N_8096,N_1021,N_4464);
nand U8097 (N_8097,N_603,N_2353);
and U8098 (N_8098,N_2610,N_4493);
xor U8099 (N_8099,N_3751,N_4499);
nor U8100 (N_8100,N_5622,N_5041);
nand U8101 (N_8101,N_887,N_526);
and U8102 (N_8102,N_1152,N_4699);
and U8103 (N_8103,N_1485,N_2674);
xor U8104 (N_8104,N_5390,N_1226);
xnor U8105 (N_8105,N_1455,N_4693);
and U8106 (N_8106,N_958,N_1619);
and U8107 (N_8107,N_1115,N_2335);
or U8108 (N_8108,N_1037,N_4043);
or U8109 (N_8109,N_5724,N_2593);
and U8110 (N_8110,N_5824,N_1314);
nand U8111 (N_8111,N_1787,N_1656);
or U8112 (N_8112,N_2110,N_976);
or U8113 (N_8113,N_3429,N_5960);
xnor U8114 (N_8114,N_2994,N_3459);
nand U8115 (N_8115,N_2919,N_5439);
or U8116 (N_8116,N_3985,N_4943);
xor U8117 (N_8117,N_4245,N_3530);
nor U8118 (N_8118,N_4477,N_1418);
or U8119 (N_8119,N_1784,N_3765);
and U8120 (N_8120,N_4865,N_3648);
or U8121 (N_8121,N_5593,N_2309);
or U8122 (N_8122,N_3857,N_2042);
and U8123 (N_8123,N_5387,N_2769);
nor U8124 (N_8124,N_993,N_2300);
nor U8125 (N_8125,N_4315,N_3357);
or U8126 (N_8126,N_295,N_5716);
xor U8127 (N_8127,N_4280,N_4382);
nand U8128 (N_8128,N_5731,N_3258);
nor U8129 (N_8129,N_1880,N_937);
nand U8130 (N_8130,N_2620,N_1836);
nand U8131 (N_8131,N_2411,N_4710);
nand U8132 (N_8132,N_1363,N_1754);
xnor U8133 (N_8133,N_4675,N_3435);
xnor U8134 (N_8134,N_4757,N_4215);
nor U8135 (N_8135,N_5417,N_1752);
nand U8136 (N_8136,N_581,N_1408);
nand U8137 (N_8137,N_3477,N_5447);
nor U8138 (N_8138,N_1571,N_4495);
and U8139 (N_8139,N_4945,N_5111);
nand U8140 (N_8140,N_3124,N_1914);
or U8141 (N_8141,N_5764,N_2856);
nor U8142 (N_8142,N_1148,N_3047);
nand U8143 (N_8143,N_400,N_3839);
nand U8144 (N_8144,N_5930,N_5609);
and U8145 (N_8145,N_4380,N_2231);
and U8146 (N_8146,N_5525,N_351);
or U8147 (N_8147,N_652,N_1092);
xnor U8148 (N_8148,N_1526,N_5836);
nand U8149 (N_8149,N_5198,N_1794);
or U8150 (N_8150,N_1768,N_994);
and U8151 (N_8151,N_2044,N_3455);
and U8152 (N_8152,N_152,N_2788);
nand U8153 (N_8153,N_1399,N_807);
and U8154 (N_8154,N_165,N_4625);
or U8155 (N_8155,N_809,N_793);
xnor U8156 (N_8156,N_3005,N_4188);
nor U8157 (N_8157,N_3975,N_5009);
xor U8158 (N_8158,N_3271,N_4304);
xnor U8159 (N_8159,N_54,N_2938);
nand U8160 (N_8160,N_245,N_4313);
and U8161 (N_8161,N_3831,N_2186);
xor U8162 (N_8162,N_1763,N_5528);
and U8163 (N_8163,N_1630,N_5077);
xnor U8164 (N_8164,N_4106,N_2429);
xor U8165 (N_8165,N_1524,N_2051);
nor U8166 (N_8166,N_3192,N_1445);
or U8167 (N_8167,N_2747,N_5263);
and U8168 (N_8168,N_2359,N_2822);
xnor U8169 (N_8169,N_4170,N_3735);
xnor U8170 (N_8170,N_4353,N_1958);
xnor U8171 (N_8171,N_2521,N_5102);
xnor U8172 (N_8172,N_2729,N_439);
nand U8173 (N_8173,N_642,N_3317);
nor U8174 (N_8174,N_16,N_776);
nand U8175 (N_8175,N_3927,N_2316);
or U8176 (N_8176,N_2737,N_1492);
nor U8177 (N_8177,N_5578,N_4474);
nand U8178 (N_8178,N_136,N_5567);
nand U8179 (N_8179,N_3780,N_4725);
xor U8180 (N_8180,N_2062,N_4224);
and U8181 (N_8181,N_3566,N_909);
or U8182 (N_8182,N_1575,N_2387);
and U8183 (N_8183,N_1637,N_2431);
nor U8184 (N_8184,N_4964,N_5682);
nand U8185 (N_8185,N_3151,N_5531);
and U8186 (N_8186,N_52,N_2522);
nor U8187 (N_8187,N_1728,N_1059);
xnor U8188 (N_8188,N_3597,N_1953);
or U8189 (N_8189,N_4461,N_5533);
nand U8190 (N_8190,N_2668,N_4729);
nor U8191 (N_8191,N_2357,N_4498);
and U8192 (N_8192,N_5450,N_4535);
nor U8193 (N_8193,N_3674,N_1638);
xor U8194 (N_8194,N_3416,N_2458);
nor U8195 (N_8195,N_1762,N_1170);
or U8196 (N_8196,N_2050,N_3494);
nor U8197 (N_8197,N_3240,N_5274);
nand U8198 (N_8198,N_4302,N_4518);
or U8199 (N_8199,N_2679,N_3380);
xor U8200 (N_8200,N_3800,N_2664);
nor U8201 (N_8201,N_5150,N_230);
and U8202 (N_8202,N_5005,N_3739);
or U8203 (N_8203,N_3365,N_3036);
and U8204 (N_8204,N_2958,N_1517);
and U8205 (N_8205,N_4589,N_1681);
or U8206 (N_8206,N_3687,N_3040);
and U8207 (N_8207,N_5325,N_1874);
or U8208 (N_8208,N_2770,N_2554);
nor U8209 (N_8209,N_2408,N_2874);
nand U8210 (N_8210,N_1229,N_409);
or U8211 (N_8211,N_5458,N_131);
nand U8212 (N_8212,N_959,N_2847);
or U8213 (N_8213,N_1475,N_3904);
xor U8214 (N_8214,N_1111,N_4452);
nand U8215 (N_8215,N_3549,N_609);
xnor U8216 (N_8216,N_2318,N_1778);
and U8217 (N_8217,N_3170,N_459);
and U8218 (N_8218,N_161,N_2810);
nand U8219 (N_8219,N_880,N_5280);
xor U8220 (N_8220,N_3244,N_5588);
xnor U8221 (N_8221,N_5461,N_3169);
xor U8222 (N_8222,N_4047,N_1222);
xor U8223 (N_8223,N_4624,N_1090);
nor U8224 (N_8224,N_5569,N_4228);
nor U8225 (N_8225,N_1,N_293);
xnor U8226 (N_8226,N_5381,N_1316);
nand U8227 (N_8227,N_2061,N_2029);
nor U8228 (N_8228,N_2252,N_3900);
nor U8229 (N_8229,N_847,N_4979);
or U8230 (N_8230,N_1590,N_23);
nand U8231 (N_8231,N_1067,N_660);
and U8232 (N_8232,N_5493,N_5157);
nor U8233 (N_8233,N_208,N_1253);
and U8234 (N_8234,N_704,N_1244);
xnor U8235 (N_8235,N_1078,N_4997);
xor U8236 (N_8236,N_5267,N_5662);
nor U8237 (N_8237,N_3498,N_637);
and U8238 (N_8238,N_3692,N_3846);
or U8239 (N_8239,N_267,N_5922);
nor U8240 (N_8240,N_1413,N_4297);
or U8241 (N_8241,N_1854,N_2617);
nor U8242 (N_8242,N_4417,N_1956);
nor U8243 (N_8243,N_3795,N_3697);
xnor U8244 (N_8244,N_4647,N_2275);
or U8245 (N_8245,N_2876,N_5153);
and U8246 (N_8246,N_3931,N_2615);
and U8247 (N_8247,N_3413,N_4428);
or U8248 (N_8248,N_824,N_4333);
or U8249 (N_8249,N_4609,N_2944);
nand U8250 (N_8250,N_4571,N_1101);
or U8251 (N_8251,N_4807,N_4568);
and U8252 (N_8252,N_4351,N_607);
nor U8253 (N_8253,N_947,N_4848);
nor U8254 (N_8254,N_5317,N_910);
or U8255 (N_8255,N_5804,N_5744);
or U8256 (N_8256,N_597,N_3737);
or U8257 (N_8257,N_5358,N_3982);
or U8258 (N_8258,N_3612,N_1509);
or U8259 (N_8259,N_5733,N_4833);
and U8260 (N_8260,N_5870,N_4936);
nand U8261 (N_8261,N_5742,N_3953);
nor U8262 (N_8262,N_79,N_1354);
and U8263 (N_8263,N_4944,N_5669);
or U8264 (N_8264,N_2712,N_3579);
and U8265 (N_8265,N_4830,N_2882);
nor U8266 (N_8266,N_1512,N_255);
nand U8267 (N_8267,N_5616,N_1696);
or U8268 (N_8268,N_1684,N_4998);
xor U8269 (N_8269,N_4169,N_4858);
or U8270 (N_8270,N_2196,N_5454);
or U8271 (N_8271,N_4875,N_2261);
nor U8272 (N_8272,N_2696,N_338);
nand U8273 (N_8273,N_618,N_2255);
and U8274 (N_8274,N_3065,N_2917);
and U8275 (N_8275,N_3654,N_348);
nand U8276 (N_8276,N_2227,N_318);
nor U8277 (N_8277,N_3462,N_4694);
nor U8278 (N_8278,N_3717,N_2189);
and U8279 (N_8279,N_4818,N_510);
xnor U8280 (N_8280,N_1008,N_5923);
nor U8281 (N_8281,N_3503,N_5904);
nand U8282 (N_8282,N_3986,N_253);
xor U8283 (N_8283,N_4119,N_2054);
nor U8284 (N_8284,N_5705,N_5391);
xnor U8285 (N_8285,N_2683,N_935);
xnor U8286 (N_8286,N_5968,N_222);
nand U8287 (N_8287,N_5890,N_5365);
nor U8288 (N_8288,N_4038,N_1336);
nor U8289 (N_8289,N_3972,N_2334);
nand U8290 (N_8290,N_5704,N_1127);
xnor U8291 (N_8291,N_1570,N_3677);
xnor U8292 (N_8292,N_3430,N_1731);
or U8293 (N_8293,N_2595,N_327);
or U8294 (N_8294,N_1503,N_4864);
nand U8295 (N_8295,N_594,N_5097);
and U8296 (N_8296,N_2405,N_840);
or U8297 (N_8297,N_1471,N_2064);
nand U8298 (N_8298,N_5784,N_5052);
nor U8299 (N_8299,N_58,N_2772);
xor U8300 (N_8300,N_2039,N_2546);
nor U8301 (N_8301,N_5268,N_2338);
or U8302 (N_8302,N_3411,N_5779);
or U8303 (N_8303,N_2013,N_1192);
xnor U8304 (N_8304,N_876,N_1113);
nand U8305 (N_8305,N_4446,N_496);
and U8306 (N_8306,N_2248,N_2018);
nand U8307 (N_8307,N_2776,N_4543);
xnor U8308 (N_8308,N_4326,N_2898);
nand U8309 (N_8309,N_457,N_1450);
nor U8310 (N_8310,N_5886,N_2492);
and U8311 (N_8311,N_2465,N_2380);
and U8312 (N_8312,N_2699,N_5519);
or U8313 (N_8313,N_5476,N_4261);
and U8314 (N_8314,N_942,N_5307);
and U8315 (N_8315,N_4826,N_687);
xnor U8316 (N_8316,N_4780,N_5137);
nand U8317 (N_8317,N_4792,N_122);
or U8318 (N_8318,N_4225,N_4491);
xor U8319 (N_8319,N_5422,N_2273);
nor U8320 (N_8320,N_5847,N_2422);
nand U8321 (N_8321,N_399,N_4822);
nand U8322 (N_8322,N_881,N_361);
nor U8323 (N_8323,N_961,N_4806);
nor U8324 (N_8324,N_5839,N_328);
or U8325 (N_8325,N_869,N_1908);
xnor U8326 (N_8326,N_923,N_4342);
and U8327 (N_8327,N_1125,N_5070);
and U8328 (N_8328,N_1004,N_67);
nand U8329 (N_8329,N_3064,N_5774);
xor U8330 (N_8330,N_2157,N_5663);
nand U8331 (N_8331,N_5159,N_4184);
nand U8332 (N_8332,N_5576,N_5222);
and U8333 (N_8333,N_1578,N_5191);
and U8334 (N_8334,N_1513,N_2272);
nand U8335 (N_8335,N_2840,N_3847);
xnor U8336 (N_8336,N_719,N_2133);
and U8337 (N_8337,N_5035,N_2517);
xor U8338 (N_8338,N_4104,N_5765);
and U8339 (N_8339,N_2214,N_563);
xor U8340 (N_8340,N_1810,N_912);
nand U8341 (N_8341,N_1679,N_2838);
nand U8342 (N_8342,N_1939,N_2456);
xnor U8343 (N_8343,N_5699,N_5046);
nor U8344 (N_8344,N_440,N_97);
xor U8345 (N_8345,N_5451,N_4492);
xor U8346 (N_8346,N_4912,N_1129);
nor U8347 (N_8347,N_2471,N_5793);
and U8348 (N_8348,N_1433,N_148);
nand U8349 (N_8349,N_3137,N_2985);
nor U8350 (N_8350,N_4236,N_4533);
nor U8351 (N_8351,N_2606,N_234);
and U8352 (N_8352,N_3486,N_3813);
xnor U8353 (N_8353,N_5082,N_3307);
or U8354 (N_8354,N_2493,N_1868);
and U8355 (N_8355,N_924,N_4972);
nand U8356 (N_8356,N_3866,N_2499);
and U8357 (N_8357,N_4754,N_2251);
and U8358 (N_8358,N_1112,N_2971);
or U8359 (N_8359,N_2601,N_1466);
or U8360 (N_8360,N_5330,N_4988);
and U8361 (N_8361,N_5801,N_1547);
or U8362 (N_8362,N_4991,N_675);
nand U8363 (N_8363,N_4824,N_436);
nand U8364 (N_8364,N_4456,N_2834);
and U8365 (N_8365,N_1283,N_3438);
nand U8366 (N_8366,N_2470,N_1852);
and U8367 (N_8367,N_4989,N_4421);
nand U8368 (N_8368,N_1225,N_5912);
and U8369 (N_8369,N_3407,N_4032);
nor U8370 (N_8370,N_2579,N_2896);
or U8371 (N_8371,N_2327,N_1494);
xor U8372 (N_8372,N_5758,N_5604);
or U8373 (N_8373,N_264,N_3031);
or U8374 (N_8374,N_4721,N_5316);
nand U8375 (N_8375,N_314,N_5000);
nor U8376 (N_8376,N_1202,N_2330);
and U8377 (N_8377,N_2619,N_4310);
nor U8378 (N_8378,N_4340,N_3264);
xnor U8379 (N_8379,N_1576,N_4552);
xor U8380 (N_8380,N_1889,N_1720);
or U8381 (N_8381,N_3463,N_1486);
xor U8382 (N_8382,N_2423,N_3425);
and U8383 (N_8383,N_2703,N_4238);
nor U8384 (N_8384,N_934,N_5049);
nor U8385 (N_8385,N_3663,N_3032);
xor U8386 (N_8386,N_5939,N_2149);
nor U8387 (N_8387,N_2633,N_5189);
or U8388 (N_8388,N_734,N_5107);
and U8389 (N_8389,N_574,N_2439);
xnor U8390 (N_8390,N_3559,N_3147);
and U8391 (N_8391,N_2953,N_4617);
xor U8392 (N_8392,N_95,N_2399);
nand U8393 (N_8393,N_2578,N_2236);
xnor U8394 (N_8394,N_1230,N_4497);
nor U8395 (N_8395,N_4240,N_115);
xnor U8396 (N_8396,N_2954,N_5187);
or U8397 (N_8397,N_3378,N_2290);
xnor U8398 (N_8398,N_5398,N_2866);
nand U8399 (N_8399,N_194,N_630);
and U8400 (N_8400,N_4723,N_1770);
nand U8401 (N_8401,N_3784,N_2759);
and U8402 (N_8402,N_5036,N_1697);
xor U8403 (N_8403,N_2659,N_1155);
nor U8404 (N_8404,N_63,N_1557);
or U8405 (N_8405,N_2967,N_4614);
or U8406 (N_8406,N_5113,N_4134);
and U8407 (N_8407,N_4392,N_2455);
nand U8408 (N_8408,N_4649,N_5873);
or U8409 (N_8409,N_5748,N_3615);
or U8410 (N_8410,N_4651,N_2372);
nand U8411 (N_8411,N_405,N_421);
nand U8412 (N_8412,N_888,N_5783);
nand U8413 (N_8413,N_5551,N_1837);
nand U8414 (N_8414,N_401,N_3742);
nor U8415 (N_8415,N_1325,N_3220);
nor U8416 (N_8416,N_3880,N_4959);
and U8417 (N_8417,N_3202,N_2278);
and U8418 (N_8418,N_3466,N_1052);
or U8419 (N_8419,N_1308,N_4283);
and U8420 (N_8420,N_5554,N_4662);
xor U8421 (N_8421,N_2376,N_1390);
nor U8422 (N_8422,N_1886,N_2211);
and U8423 (N_8423,N_949,N_5348);
and U8424 (N_8424,N_322,N_1128);
nand U8425 (N_8425,N_4457,N_425);
and U8426 (N_8426,N_1937,N_4931);
and U8427 (N_8427,N_3914,N_5069);
nor U8428 (N_8428,N_3892,N_1780);
xnor U8429 (N_8429,N_4902,N_999);
nand U8430 (N_8430,N_3177,N_3995);
nor U8431 (N_8431,N_378,N_2786);
xor U8432 (N_8432,N_513,N_5065);
and U8433 (N_8433,N_3245,N_2890);
xor U8434 (N_8434,N_5532,N_5770);
nand U8435 (N_8435,N_2367,N_1267);
xor U8436 (N_8436,N_5403,N_1180);
nor U8437 (N_8437,N_4276,N_4289);
xor U8438 (N_8438,N_2419,N_2107);
nor U8439 (N_8439,N_1733,N_4741);
nor U8440 (N_8440,N_1530,N_5264);
and U8441 (N_8441,N_5308,N_542);
nor U8442 (N_8442,N_2243,N_962);
or U8443 (N_8443,N_4663,N_1620);
or U8444 (N_8444,N_5694,N_4348);
or U8445 (N_8445,N_330,N_5978);
or U8446 (N_8446,N_3250,N_5158);
or U8447 (N_8447,N_2932,N_3537);
nand U8448 (N_8448,N_5782,N_2920);
or U8449 (N_8449,N_5695,N_5109);
nor U8450 (N_8450,N_482,N_3288);
nand U8451 (N_8451,N_2053,N_4674);
or U8452 (N_8452,N_1604,N_4772);
xor U8453 (N_8453,N_1999,N_3845);
nor U8454 (N_8454,N_2445,N_279);
and U8455 (N_8455,N_4317,N_3451);
xor U8456 (N_8456,N_782,N_5749);
or U8457 (N_8457,N_1270,N_2887);
nor U8458 (N_8458,N_2628,N_3546);
and U8459 (N_8459,N_18,N_2241);
nand U8460 (N_8460,N_1848,N_3580);
nand U8461 (N_8461,N_1685,N_5389);
xor U8462 (N_8462,N_51,N_2172);
nor U8463 (N_8463,N_4957,N_3910);
nand U8464 (N_8464,N_2424,N_4621);
and U8465 (N_8465,N_5227,N_1197);
xor U8466 (N_8466,N_3743,N_5430);
nand U8467 (N_8467,N_1802,N_1288);
xnor U8468 (N_8468,N_443,N_5341);
or U8469 (N_8469,N_233,N_3966);
nand U8470 (N_8470,N_124,N_4311);
nand U8471 (N_8471,N_1829,N_2511);
nand U8472 (N_8472,N_1657,N_4140);
and U8473 (N_8473,N_5896,N_5688);
nand U8474 (N_8474,N_3260,N_5745);
nor U8475 (N_8475,N_5392,N_1302);
xnor U8476 (N_8476,N_3387,N_137);
nor U8477 (N_8477,N_2733,N_316);
nor U8478 (N_8478,N_168,N_2259);
and U8479 (N_8479,N_3283,N_2047);
or U8480 (N_8480,N_4469,N_1918);
or U8481 (N_8481,N_3716,N_2587);
xnor U8482 (N_8482,N_3571,N_506);
or U8483 (N_8483,N_1282,N_4740);
xor U8484 (N_8484,N_2648,N_4485);
nor U8485 (N_8485,N_5891,N_4643);
xor U8486 (N_8486,N_5169,N_3385);
and U8487 (N_8487,N_5223,N_2913);
nand U8488 (N_8488,N_2244,N_2631);
nor U8489 (N_8489,N_5986,N_2736);
nor U8490 (N_8490,N_647,N_1232);
xnor U8491 (N_8491,N_4897,N_2912);
or U8492 (N_8492,N_3011,N_3006);
or U8493 (N_8493,N_4003,N_4983);
nand U8494 (N_8494,N_4557,N_4753);
xnor U8495 (N_8495,N_2083,N_5878);
or U8496 (N_8496,N_4639,N_856);
xor U8497 (N_8497,N_4176,N_4361);
or U8498 (N_8498,N_1982,N_1015);
nor U8499 (N_8499,N_83,N_2506);
nand U8500 (N_8500,N_2760,N_5099);
xor U8501 (N_8501,N_5942,N_4751);
nand U8502 (N_8502,N_4924,N_518);
and U8503 (N_8503,N_470,N_1333);
xor U8504 (N_8504,N_5039,N_602);
xnor U8505 (N_8505,N_3741,N_5366);
or U8506 (N_8506,N_3747,N_239);
xnor U8507 (N_8507,N_5825,N_5938);
and U8508 (N_8508,N_3003,N_1319);
or U8509 (N_8509,N_3905,N_913);
xor U8510 (N_8510,N_1683,N_3855);
xnor U8511 (N_8511,N_5001,N_3415);
xnor U8512 (N_8512,N_489,N_5329);
nand U8513 (N_8513,N_4831,N_143);
nand U8514 (N_8514,N_3198,N_2015);
xor U8515 (N_8515,N_1950,N_4763);
xor U8516 (N_8516,N_70,N_4714);
nand U8517 (N_8517,N_2927,N_2692);
nor U8518 (N_8518,N_1427,N_5418);
xnor U8519 (N_8519,N_3128,N_1020);
and U8520 (N_8520,N_3327,N_2406);
nand U8521 (N_8521,N_3519,N_3444);
xnor U8522 (N_8522,N_5170,N_5611);
nand U8523 (N_8523,N_1055,N_2138);
and U8524 (N_8524,N_3630,N_2556);
nand U8525 (N_8525,N_1675,N_252);
nor U8526 (N_8526,N_5974,N_2557);
nand U8527 (N_8527,N_5085,N_4680);
nor U8528 (N_8528,N_5787,N_641);
nor U8529 (N_8529,N_1873,N_2179);
and U8530 (N_8530,N_1133,N_3362);
xor U8531 (N_8531,N_5286,N_3417);
xnor U8532 (N_8532,N_1198,N_957);
xor U8533 (N_8533,N_5522,N_1407);
xnor U8534 (N_8534,N_4269,N_5499);
or U8535 (N_8535,N_5495,N_2276);
nor U8536 (N_8536,N_2533,N_4825);
and U8537 (N_8537,N_4030,N_1495);
nor U8538 (N_8538,N_4873,N_1287);
or U8539 (N_8539,N_59,N_4222);
xor U8540 (N_8540,N_1870,N_5947);
nand U8541 (N_8541,N_795,N_3182);
nand U8542 (N_8542,N_5237,N_4918);
nor U8543 (N_8543,N_2503,N_5788);
xor U8544 (N_8544,N_3058,N_4923);
and U8545 (N_8545,N_1705,N_5658);
or U8546 (N_8546,N_3311,N_3601);
nor U8547 (N_8547,N_3525,N_138);
and U8548 (N_8548,N_3132,N_2427);
nand U8549 (N_8549,N_2702,N_3957);
nand U8550 (N_8550,N_1740,N_1400);
or U8551 (N_8551,N_5590,N_2216);
or U8552 (N_8552,N_2908,N_1546);
and U8553 (N_8553,N_375,N_4075);
nand U8554 (N_8554,N_3280,N_3508);
nand U8555 (N_8555,N_4876,N_4250);
nor U8556 (N_8556,N_569,N_5910);
nor U8557 (N_8557,N_3185,N_2704);
nand U8558 (N_8558,N_2895,N_4402);
and U8559 (N_8559,N_4916,N_5093);
or U8560 (N_8560,N_5712,N_5959);
nor U8561 (N_8561,N_556,N_4735);
or U8562 (N_8562,N_4678,N_5517);
and U8563 (N_8563,N_2972,N_3126);
and U8564 (N_8564,N_5727,N_2516);
and U8565 (N_8565,N_3867,N_4370);
nor U8566 (N_8566,N_3766,N_1217);
nand U8567 (N_8567,N_4200,N_1757);
nor U8568 (N_8568,N_2128,N_1375);
and U8569 (N_8569,N_1195,N_3771);
xor U8570 (N_8570,N_2410,N_710);
and U8571 (N_8571,N_1306,N_3072);
nor U8572 (N_8572,N_4975,N_286);
nor U8573 (N_8573,N_2351,N_1830);
and U8574 (N_8574,N_1435,N_2173);
or U8575 (N_8575,N_943,N_3071);
or U8576 (N_8576,N_1594,N_933);
and U8577 (N_8577,N_963,N_2382);
nor U8578 (N_8578,N_114,N_1706);
or U8579 (N_8579,N_2519,N_5469);
nand U8580 (N_8580,N_816,N_2732);
nand U8581 (N_8581,N_2505,N_3637);
and U8582 (N_8582,N_3779,N_1581);
or U8583 (N_8583,N_777,N_3055);
nand U8584 (N_8584,N_3481,N_4144);
nor U8585 (N_8585,N_4468,N_1979);
nand U8586 (N_8586,N_160,N_4273);
xor U8587 (N_8587,N_167,N_2942);
xor U8588 (N_8588,N_5812,N_3623);
nor U8589 (N_8589,N_5542,N_557);
nand U8590 (N_8590,N_3216,N_4442);
and U8591 (N_8591,N_4487,N_2590);
or U8592 (N_8592,N_2105,N_417);
xnor U8593 (N_8593,N_2206,N_3329);
nand U8594 (N_8594,N_2817,N_1057);
nor U8595 (N_8595,N_1648,N_2111);
nor U8596 (N_8596,N_433,N_5872);
nand U8597 (N_8597,N_1161,N_4408);
nand U8598 (N_8598,N_5880,N_5174);
xor U8599 (N_8599,N_1971,N_595);
or U8600 (N_8600,N_4201,N_5685);
or U8601 (N_8601,N_4790,N_4122);
nor U8602 (N_8602,N_5982,N_336);
and U8603 (N_8603,N_2992,N_3130);
and U8604 (N_8604,N_269,N_2480);
and U8605 (N_8605,N_4007,N_4937);
nand U8606 (N_8606,N_5951,N_3168);
nor U8607 (N_8607,N_1860,N_2396);
or U8608 (N_8608,N_5911,N_4137);
and U8609 (N_8609,N_4330,N_4599);
xnor U8610 (N_8610,N_4060,N_414);
or U8611 (N_8611,N_3187,N_3083);
nor U8612 (N_8612,N_571,N_1334);
nor U8613 (N_8613,N_1940,N_5420);
nor U8614 (N_8614,N_1716,N_455);
nor U8615 (N_8615,N_3166,N_5635);
xor U8616 (N_8616,N_4127,N_5017);
or U8617 (N_8617,N_5503,N_931);
nand U8618 (N_8618,N_930,N_701);
xnor U8619 (N_8619,N_4856,N_2608);
and U8620 (N_8620,N_74,N_1849);
xnor U8621 (N_8621,N_1406,N_1687);
nand U8622 (N_8622,N_5303,N_3228);
xnor U8623 (N_8623,N_1328,N_3793);
nor U8624 (N_8624,N_2905,N_1496);
and U8625 (N_8625,N_4862,N_753);
nor U8626 (N_8626,N_4982,N_4676);
nand U8627 (N_8627,N_5434,N_3399);
and U8628 (N_8628,N_2843,N_3125);
and U8629 (N_8629,N_3106,N_2407);
nor U8630 (N_8630,N_1430,N_1923);
xnor U8631 (N_8631,N_3178,N_5647);
and U8632 (N_8632,N_3162,N_3221);
nor U8633 (N_8633,N_5347,N_5864);
or U8634 (N_8634,N_5421,N_1183);
xnor U8635 (N_8635,N_5110,N_5772);
nand U8636 (N_8636,N_4124,N_1147);
and U8637 (N_8637,N_2600,N_5946);
or U8638 (N_8638,N_4514,N_5881);
xnor U8639 (N_8639,N_2084,N_1636);
or U8640 (N_8640,N_3512,N_5470);
and U8641 (N_8641,N_2009,N_88);
and U8642 (N_8642,N_5718,N_4669);
and U8643 (N_8643,N_3146,N_3196);
nand U8644 (N_8644,N_654,N_1420);
xnor U8645 (N_8645,N_1925,N_2072);
nor U8646 (N_8646,N_5273,N_3514);
xnor U8647 (N_8647,N_2612,N_2027);
or U8648 (N_8648,N_3419,N_5294);
or U8649 (N_8649,N_1345,N_5357);
and U8650 (N_8650,N_69,N_3732);
nand U8651 (N_8651,N_1428,N_1866);
or U8652 (N_8652,N_392,N_878);
and U8653 (N_8653,N_1838,N_3268);
xor U8654 (N_8654,N_5996,N_2894);
nand U8655 (N_8655,N_505,N_2285);
or U8656 (N_8656,N_4577,N_922);
nor U8657 (N_8657,N_1065,N_716);
xnor U8658 (N_8658,N_2463,N_3543);
xor U8659 (N_8659,N_1523,N_2687);
nor U8660 (N_8660,N_3801,N_4412);
or U8661 (N_8661,N_4660,N_653);
and U8662 (N_8662,N_1442,N_2356);
or U8663 (N_8663,N_2846,N_4083);
nor U8664 (N_8664,N_2355,N_217);
nand U8665 (N_8665,N_3267,N_2560);
and U8666 (N_8666,N_3446,N_4788);
or U8667 (N_8667,N_3022,N_1972);
nor U8668 (N_8668,N_5714,N_5010);
xnor U8669 (N_8669,N_477,N_623);
xnor U8670 (N_8670,N_3563,N_918);
nor U8671 (N_8671,N_5456,N_4133);
or U8672 (N_8672,N_4400,N_969);
and U8673 (N_8673,N_4386,N_5193);
nor U8674 (N_8674,N_5377,N_4737);
xnor U8675 (N_8675,N_3026,N_1853);
nand U8676 (N_8676,N_4874,N_73);
xnor U8677 (N_8677,N_103,N_3300);
and U8678 (N_8678,N_4062,N_3672);
or U8679 (N_8679,N_3762,N_325);
nor U8680 (N_8680,N_3791,N_1072);
nand U8681 (N_8681,N_100,N_2205);
nor U8682 (N_8682,N_3024,N_2642);
nor U8683 (N_8683,N_1303,N_1204);
nor U8684 (N_8684,N_297,N_2844);
xor U8685 (N_8685,N_5850,N_2934);
or U8686 (N_8686,N_2947,N_4814);
and U8687 (N_8687,N_5631,N_5973);
nor U8688 (N_8688,N_2995,N_2870);
xnor U8689 (N_8689,N_5236,N_3134);
nand U8690 (N_8690,N_1385,N_1521);
nand U8691 (N_8691,N_836,N_4985);
xor U8692 (N_8692,N_2143,N_5364);
and U8693 (N_8693,N_2085,N_2666);
and U8694 (N_8694,N_5446,N_3483);
xor U8695 (N_8695,N_3841,N_2568);
or U8696 (N_8696,N_4974,N_1027);
nor U8697 (N_8697,N_1703,N_4898);
nor U8698 (N_8698,N_2806,N_2877);
xnor U8699 (N_8699,N_800,N_4367);
nand U8700 (N_8700,N_772,N_454);
and U8701 (N_8701,N_323,N_1262);
and U8702 (N_8702,N_2165,N_448);
nor U8703 (N_8703,N_1917,N_1224);
nand U8704 (N_8704,N_3551,N_674);
nand U8705 (N_8705,N_5278,N_2137);
and U8706 (N_8706,N_2124,N_3656);
or U8707 (N_8707,N_5642,N_2035);
xnor U8708 (N_8708,N_2868,N_1135);
nor U8709 (N_8709,N_5898,N_200);
nand U8710 (N_8710,N_833,N_1031);
nand U8711 (N_8711,N_1712,N_2748);
nor U8712 (N_8712,N_2099,N_2307);
xor U8713 (N_8713,N_5063,N_4031);
nand U8714 (N_8714,N_2223,N_188);
nor U8715 (N_8715,N_3165,N_1507);
and U8716 (N_8716,N_1828,N_2008);
xnor U8717 (N_8717,N_2154,N_3426);
and U8718 (N_8718,N_5556,N_519);
and U8719 (N_8719,N_2242,N_1963);
and U8720 (N_8720,N_4949,N_3994);
or U8721 (N_8721,N_5288,N_4758);
nor U8722 (N_8722,N_5972,N_5879);
or U8723 (N_8723,N_2453,N_5624);
or U8724 (N_8724,N_5971,N_4656);
and U8725 (N_8725,N_1122,N_1909);
nor U8726 (N_8726,N_4076,N_2473);
nand U8727 (N_8727,N_3539,N_60);
or U8728 (N_8728,N_1279,N_3358);
xnor U8729 (N_8729,N_3830,N_4719);
nand U8730 (N_8730,N_2352,N_3955);
nor U8731 (N_8731,N_4928,N_1897);
or U8732 (N_8732,N_1946,N_3757);
nor U8733 (N_8733,N_4628,N_447);
nor U8734 (N_8734,N_1397,N_2653);
and U8735 (N_8735,N_4397,N_1834);
nor U8736 (N_8736,N_817,N_304);
xnor U8737 (N_8737,N_4429,N_842);
xor U8738 (N_8738,N_3212,N_1845);
or U8739 (N_8739,N_2254,N_55);
or U8740 (N_8740,N_2395,N_3229);
or U8741 (N_8741,N_4065,N_1573);
and U8742 (N_8742,N_3936,N_2853);
nand U8743 (N_8743,N_3908,N_5332);
xor U8744 (N_8744,N_1380,N_5901);
and U8745 (N_8745,N_2328,N_3188);
nor U8746 (N_8746,N_4443,N_3821);
and U8747 (N_8747,N_5012,N_3496);
nor U8748 (N_8748,N_5477,N_4312);
nand U8749 (N_8749,N_4696,N_2220);
and U8750 (N_8750,N_2489,N_1532);
nand U8751 (N_8751,N_668,N_2996);
and U8752 (N_8752,N_2929,N_449);
xor U8753 (N_8753,N_2253,N_4168);
nor U8754 (N_8754,N_614,N_2314);
nor U8755 (N_8755,N_2559,N_5188);
nor U8756 (N_8756,N_1114,N_784);
and U8757 (N_8757,N_1102,N_4604);
and U8758 (N_8758,N_3678,N_5943);
xnor U8759 (N_8759,N_2375,N_5200);
nor U8760 (N_8760,N_2941,N_1973);
nand U8761 (N_8761,N_2291,N_6);
nand U8762 (N_8762,N_48,N_2310);
nor U8763 (N_8763,N_3043,N_764);
nor U8764 (N_8764,N_552,N_4879);
or U8765 (N_8765,N_104,N_2132);
nor U8766 (N_8766,N_150,N_899);
nor U8767 (N_8767,N_5014,N_1350);
nor U8768 (N_8768,N_988,N_5496);
or U8769 (N_8769,N_875,N_3282);
nor U8770 (N_8770,N_113,N_5141);
xor U8771 (N_8771,N_5120,N_2982);
nand U8772 (N_8772,N_1298,N_1519);
xor U8773 (N_8773,N_335,N_2741);
nand U8774 (N_8774,N_5786,N_584);
nand U8775 (N_8775,N_4166,N_1538);
nor U8776 (N_8776,N_319,N_760);
or U8777 (N_8777,N_3095,N_5618);
or U8778 (N_8778,N_3105,N_4859);
xor U8779 (N_8779,N_1585,N_3728);
nor U8780 (N_8780,N_3377,N_3197);
xor U8781 (N_8781,N_461,N_4648);
xor U8782 (N_8782,N_2634,N_4805);
nand U8783 (N_8783,N_1617,N_2607);
or U8784 (N_8784,N_4840,N_4203);
or U8785 (N_8785,N_2632,N_308);
or U8786 (N_8786,N_4598,N_3555);
nand U8787 (N_8787,N_386,N_4174);
or U8788 (N_8788,N_5835,N_2765);
xor U8789 (N_8789,N_3351,N_2087);
nor U8790 (N_8790,N_2103,N_1068);
or U8791 (N_8791,N_5537,N_1299);
xor U8792 (N_8792,N_259,N_3299);
nor U8793 (N_8793,N_5680,N_4631);
nand U8794 (N_8794,N_3706,N_5122);
nand U8795 (N_8795,N_4761,N_3199);
or U8796 (N_8796,N_3807,N_1130);
and U8797 (N_8797,N_4248,N_3603);
and U8798 (N_8798,N_271,N_2529);
nor U8799 (N_8799,N_184,N_5457);
nand U8800 (N_8800,N_1171,N_2638);
xor U8801 (N_8801,N_3709,N_1335);
or U8802 (N_8802,N_4338,N_3354);
and U8803 (N_8803,N_1439,N_638);
nand U8804 (N_8804,N_832,N_4286);
and U8805 (N_8805,N_1981,N_3748);
nor U8806 (N_8806,N_689,N_2724);
xnor U8807 (N_8807,N_429,N_3402);
nand U8808 (N_8808,N_458,N_2963);
nand U8809 (N_8809,N_3902,N_2442);
and U8810 (N_8810,N_1758,N_4028);
and U8811 (N_8811,N_3870,N_4969);
and U8812 (N_8812,N_3114,N_1899);
xnor U8813 (N_8813,N_398,N_2973);
nand U8814 (N_8814,N_285,N_1285);
nand U8815 (N_8815,N_4084,N_112);
or U8816 (N_8816,N_2219,N_149);
xnor U8817 (N_8817,N_2777,N_2525);
or U8818 (N_8818,N_4583,N_4968);
nor U8819 (N_8819,N_1489,N_1451);
nand U8820 (N_8820,N_1692,N_1598);
xnor U8821 (N_8821,N_4178,N_2302);
or U8822 (N_8822,N_4619,N_4890);
xor U8823 (N_8823,N_2345,N_1964);
xor U8824 (N_8824,N_2667,N_3621);
and U8825 (N_8825,N_1628,N_2421);
xor U8826 (N_8826,N_3506,N_476);
or U8827 (N_8827,N_1470,N_2485);
or U8828 (N_8828,N_5550,N_4081);
xor U8829 (N_8829,N_908,N_1672);
nor U8830 (N_8830,N_867,N_3100);
nor U8831 (N_8831,N_469,N_5033);
nor U8832 (N_8832,N_879,N_5579);
nor U8833 (N_8833,N_4767,N_2496);
nor U8834 (N_8834,N_2461,N_472);
or U8835 (N_8835,N_4523,N_5331);
nor U8836 (N_8836,N_954,N_5547);
xnor U8837 (N_8837,N_1827,N_3401);
or U8838 (N_8838,N_4202,N_1929);
nor U8839 (N_8839,N_3524,N_2598);
and U8840 (N_8840,N_2090,N_4306);
nor U8841 (N_8841,N_3302,N_3622);
nor U8842 (N_8842,N_226,N_5414);
nand U8843 (N_8843,N_3191,N_1549);
xor U8844 (N_8844,N_626,N_1096);
xor U8845 (N_8845,N_4389,N_1661);
or U8846 (N_8846,N_523,N_3041);
and U8847 (N_8847,N_1919,N_394);
or U8848 (N_8848,N_422,N_4207);
and U8849 (N_8849,N_4439,N_823);
nand U8850 (N_8850,N_567,N_2498);
or U8851 (N_8851,N_838,N_34);
nor U8852 (N_8852,N_1372,N_1531);
nand U8853 (N_8853,N_5761,N_166);
and U8854 (N_8854,N_3129,N_3890);
nand U8855 (N_8855,N_331,N_3541);
or U8856 (N_8856,N_3331,N_2665);
nand U8857 (N_8857,N_1440,N_3750);
xor U8858 (N_8858,N_5991,N_1019);
and U8859 (N_8859,N_5168,N_3562);
and U8860 (N_8860,N_5755,N_5657);
or U8861 (N_8861,N_3874,N_116);
nor U8862 (N_8862,N_5326,N_5092);
nand U8863 (N_8863,N_2239,N_45);
nor U8864 (N_8864,N_3104,N_4866);
and U8865 (N_8865,N_1079,N_2623);
and U8866 (N_8866,N_3203,N_5425);
xnor U8867 (N_8867,N_4253,N_5356);
nand U8868 (N_8868,N_5821,N_3558);
or U8869 (N_8869,N_2282,N_521);
nor U8870 (N_8870,N_2743,N_5125);
nor U8871 (N_8871,N_3618,N_2563);
nand U8872 (N_8872,N_5586,N_3778);
xor U8873 (N_8873,N_4689,N_5732);
nand U8874 (N_8874,N_53,N_2287);
or U8875 (N_8875,N_5815,N_1351);
nor U8876 (N_8876,N_4854,N_4052);
and U8877 (N_8877,N_4100,N_4434);
nand U8878 (N_8878,N_1454,N_4239);
xnor U8879 (N_8879,N_2249,N_4087);
or U8880 (N_8880,N_3078,N_1293);
or U8881 (N_8881,N_717,N_632);
and U8882 (N_8882,N_57,N_2063);
or U8883 (N_8883,N_5424,N_5259);
nor U8884 (N_8884,N_5024,N_1460);
or U8885 (N_8885,N_2961,N_3682);
nand U8886 (N_8886,N_4527,N_5314);
or U8887 (N_8887,N_1087,N_3492);
nor U8888 (N_8888,N_1660,N_5048);
or U8889 (N_8889,N_3935,N_2555);
nand U8890 (N_8890,N_4745,N_5071);
or U8891 (N_8891,N_4768,N_444);
or U8892 (N_8892,N_4438,N_3584);
xnor U8893 (N_8893,N_2437,N_1444);
and U8894 (N_8894,N_156,N_4509);
xor U8895 (N_8895,N_380,N_4904);
or U8896 (N_8896,N_3427,N_2348);
xnor U8897 (N_8897,N_5098,N_5613);
or U8898 (N_8898,N_1344,N_2313);
or U8899 (N_8899,N_554,N_3364);
or U8900 (N_8900,N_537,N_3941);
xor U8901 (N_8901,N_4701,N_979);
nand U8902 (N_8902,N_4016,N_1474);
nand U8903 (N_8903,N_3938,N_1261);
xor U8904 (N_8904,N_1405,N_5061);
nor U8905 (N_8905,N_237,N_356);
and U8906 (N_8906,N_4612,N_4211);
or U8907 (N_8907,N_2764,N_5679);
and U8908 (N_8908,N_1959,N_1348);
nand U8909 (N_8909,N_2204,N_5468);
xnor U8910 (N_8910,N_218,N_558);
xor U8911 (N_8911,N_4079,N_498);
and U8912 (N_8912,N_1159,N_4145);
nand U8913 (N_8913,N_221,N_872);
nor U8914 (N_8914,N_1388,N_5587);
nor U8915 (N_8915,N_3923,N_3738);
xor U8916 (N_8916,N_5600,N_3719);
xor U8917 (N_8917,N_3517,N_1662);
and U8918 (N_8918,N_622,N_1249);
or U8919 (N_8919,N_5066,N_5394);
and U8920 (N_8920,N_5284,N_612);
and U8921 (N_8921,N_728,N_3028);
nor U8922 (N_8922,N_2280,N_2956);
xnor U8923 (N_8923,N_5234,N_798);
xor U8924 (N_8924,N_276,N_2508);
nand U8925 (N_8925,N_110,N_3075);
nand U8926 (N_8926,N_3848,N_3851);
nand U8927 (N_8927,N_2037,N_5806);
or U8928 (N_8928,N_2079,N_4156);
nor U8929 (N_8929,N_3110,N_1193);
or U8930 (N_8930,N_3138,N_393);
nor U8931 (N_8931,N_5142,N_2100);
nand U8932 (N_8932,N_1409,N_2845);
and U8933 (N_8933,N_5861,N_4769);
nor U8934 (N_8934,N_2349,N_1469);
xnor U8935 (N_8935,N_3467,N_3668);
xor U8936 (N_8936,N_4605,N_5829);
nand U8937 (N_8937,N_900,N_2161);
and U8938 (N_8938,N_5521,N_3313);
nand U8939 (N_8939,N_2056,N_3176);
nor U8940 (N_8940,N_973,N_1326);
nand U8941 (N_8941,N_1207,N_1504);
and U8942 (N_8942,N_1365,N_4325);
and U8943 (N_8943,N_4845,N_4774);
and U8944 (N_8944,N_1915,N_2119);
nor U8945 (N_8945,N_5655,N_1502);
xor U8946 (N_8946,N_5952,N_3950);
and U8947 (N_8947,N_3262,N_3775);
nand U8948 (N_8948,N_4430,N_5026);
or U8949 (N_8949,N_1610,N_1901);
nand U8950 (N_8950,N_1216,N_520);
or U8951 (N_8951,N_4288,N_3862);
or U8952 (N_8952,N_2911,N_3837);
or U8953 (N_8953,N_3788,N_263);
xor U8954 (N_8954,N_2240,N_1367);
and U8955 (N_8955,N_5858,N_1300);
xnor U8956 (N_8956,N_4895,N_4682);
nor U8957 (N_8957,N_4433,N_2534);
or U8958 (N_8958,N_3521,N_3665);
or U8959 (N_8959,N_1324,N_2858);
and U8960 (N_8960,N_3286,N_1459);
nor U8961 (N_8961,N_5299,N_5502);
and U8962 (N_8962,N_4357,N_2676);
xor U8963 (N_8963,N_4620,N_2939);
or U8964 (N_8964,N_4690,N_4553);
xor U8965 (N_8965,N_2922,N_2779);
nand U8966 (N_8966,N_1534,N_4728);
xnor U8967 (N_8967,N_4706,N_2217);
and U8968 (N_8968,N_5833,N_3616);
nand U8969 (N_8969,N_5919,N_5641);
xnor U8970 (N_8970,N_643,N_576);
nor U8971 (N_8971,N_453,N_41);
xnor U8972 (N_8972,N_3076,N_2491);
nand U8973 (N_8973,N_3115,N_5334);
or U8974 (N_8974,N_240,N_4884);
nand U8975 (N_8975,N_5400,N_2548);
nor U8976 (N_8976,N_4510,N_4039);
and U8977 (N_8977,N_4368,N_4090);
nand U8978 (N_8978,N_2826,N_2296);
or U8979 (N_8979,N_3773,N_2414);
nor U8980 (N_8980,N_2112,N_2909);
nand U8981 (N_8981,N_5095,N_5902);
and U8982 (N_8982,N_2589,N_2527);
and U8983 (N_8983,N_415,N_3473);
xnor U8984 (N_8984,N_3344,N_4785);
xnor U8985 (N_8985,N_3929,N_423);
nand U8986 (N_8986,N_5562,N_4022);
or U8987 (N_8987,N_4183,N_1947);
nor U8988 (N_8988,N_886,N_64);
nand U8989 (N_8989,N_5769,N_11);
xnor U8990 (N_8990,N_2371,N_2386);
nor U8991 (N_8991,N_2931,N_538);
nor U8992 (N_8992,N_2893,N_2311);
or U8993 (N_8993,N_3681,N_3371);
and U8994 (N_8994,N_317,N_1955);
nor U8995 (N_8995,N_5075,N_1210);
and U8996 (N_8996,N_3412,N_2831);
xnor U8997 (N_8997,N_5766,N_1916);
xor U8998 (N_8998,N_1825,N_1251);
and U8999 (N_8999,N_825,N_5671);
xnor U9000 (N_9000,N_962,N_4491);
nand U9001 (N_9001,N_691,N_4585);
or U9002 (N_9002,N_90,N_936);
or U9003 (N_9003,N_5607,N_3789);
nor U9004 (N_9004,N_4053,N_4403);
nor U9005 (N_9005,N_2367,N_1372);
or U9006 (N_9006,N_2096,N_5375);
or U9007 (N_9007,N_4595,N_5200);
nor U9008 (N_9008,N_2424,N_1175);
and U9009 (N_9009,N_3621,N_506);
nand U9010 (N_9010,N_2854,N_5304);
and U9011 (N_9011,N_2304,N_4589);
xor U9012 (N_9012,N_4098,N_5694);
nand U9013 (N_9013,N_4447,N_2777);
or U9014 (N_9014,N_5056,N_4868);
or U9015 (N_9015,N_2427,N_1809);
nor U9016 (N_9016,N_2032,N_1955);
and U9017 (N_9017,N_2964,N_2147);
xor U9018 (N_9018,N_324,N_1449);
nand U9019 (N_9019,N_4645,N_3101);
xor U9020 (N_9020,N_1719,N_1700);
nor U9021 (N_9021,N_4370,N_5733);
nand U9022 (N_9022,N_21,N_1779);
xor U9023 (N_9023,N_4740,N_3482);
xnor U9024 (N_9024,N_1585,N_4783);
nand U9025 (N_9025,N_416,N_586);
nor U9026 (N_9026,N_1158,N_3339);
nor U9027 (N_9027,N_1976,N_5646);
xnor U9028 (N_9028,N_1118,N_5978);
xor U9029 (N_9029,N_2524,N_225);
nand U9030 (N_9030,N_2001,N_5266);
and U9031 (N_9031,N_3720,N_5413);
xor U9032 (N_9032,N_5109,N_2985);
nor U9033 (N_9033,N_3838,N_1094);
xnor U9034 (N_9034,N_3964,N_2709);
and U9035 (N_9035,N_5295,N_1286);
nor U9036 (N_9036,N_1943,N_923);
nand U9037 (N_9037,N_2567,N_4792);
nand U9038 (N_9038,N_5165,N_2939);
and U9039 (N_9039,N_4702,N_4198);
xnor U9040 (N_9040,N_56,N_4783);
or U9041 (N_9041,N_2522,N_334);
nand U9042 (N_9042,N_1201,N_3795);
and U9043 (N_9043,N_82,N_2869);
and U9044 (N_9044,N_2677,N_2786);
nand U9045 (N_9045,N_4132,N_658);
xnor U9046 (N_9046,N_3134,N_2152);
or U9047 (N_9047,N_2207,N_801);
or U9048 (N_9048,N_5262,N_1044);
nor U9049 (N_9049,N_3629,N_1609);
nand U9050 (N_9050,N_2123,N_5789);
nor U9051 (N_9051,N_4067,N_3386);
xor U9052 (N_9052,N_4950,N_722);
or U9053 (N_9053,N_419,N_594);
nand U9054 (N_9054,N_297,N_2434);
nand U9055 (N_9055,N_2600,N_5467);
nand U9056 (N_9056,N_4656,N_1957);
xor U9057 (N_9057,N_2555,N_1326);
nor U9058 (N_9058,N_2767,N_2050);
nor U9059 (N_9059,N_5508,N_318);
nand U9060 (N_9060,N_2802,N_4813);
xor U9061 (N_9061,N_3935,N_4779);
nor U9062 (N_9062,N_5804,N_1766);
nor U9063 (N_9063,N_3507,N_2607);
or U9064 (N_9064,N_187,N_4253);
xnor U9065 (N_9065,N_1117,N_5274);
xnor U9066 (N_9066,N_5424,N_3610);
xnor U9067 (N_9067,N_4370,N_5399);
nand U9068 (N_9068,N_3170,N_1442);
nor U9069 (N_9069,N_939,N_2255);
xor U9070 (N_9070,N_1680,N_163);
nor U9071 (N_9071,N_205,N_4371);
nand U9072 (N_9072,N_2976,N_4443);
nor U9073 (N_9073,N_429,N_3280);
nor U9074 (N_9074,N_2809,N_680);
or U9075 (N_9075,N_4347,N_1568);
or U9076 (N_9076,N_3772,N_3146);
nor U9077 (N_9077,N_2765,N_3183);
or U9078 (N_9078,N_2360,N_3032);
or U9079 (N_9079,N_240,N_4410);
nor U9080 (N_9080,N_4418,N_4063);
and U9081 (N_9081,N_4103,N_3885);
xnor U9082 (N_9082,N_1314,N_1428);
and U9083 (N_9083,N_4292,N_5989);
nand U9084 (N_9084,N_4008,N_1157);
nor U9085 (N_9085,N_5070,N_1817);
xor U9086 (N_9086,N_1361,N_886);
xnor U9087 (N_9087,N_1576,N_5155);
nand U9088 (N_9088,N_5936,N_4922);
and U9089 (N_9089,N_4138,N_4804);
and U9090 (N_9090,N_5589,N_2145);
nor U9091 (N_9091,N_5739,N_3797);
nor U9092 (N_9092,N_5094,N_1112);
or U9093 (N_9093,N_65,N_1733);
nor U9094 (N_9094,N_1134,N_3425);
and U9095 (N_9095,N_1480,N_5290);
nor U9096 (N_9096,N_344,N_1155);
or U9097 (N_9097,N_3001,N_3547);
nor U9098 (N_9098,N_2910,N_4755);
and U9099 (N_9099,N_1942,N_1562);
nor U9100 (N_9100,N_1762,N_184);
nor U9101 (N_9101,N_1393,N_1094);
nor U9102 (N_9102,N_4667,N_5497);
or U9103 (N_9103,N_2442,N_5240);
and U9104 (N_9104,N_4083,N_1938);
nand U9105 (N_9105,N_1194,N_4575);
nor U9106 (N_9106,N_5874,N_3449);
nand U9107 (N_9107,N_4906,N_5260);
or U9108 (N_9108,N_5633,N_4430);
nand U9109 (N_9109,N_4192,N_562);
or U9110 (N_9110,N_5420,N_4491);
and U9111 (N_9111,N_3325,N_1624);
nor U9112 (N_9112,N_1916,N_5722);
nand U9113 (N_9113,N_2713,N_5937);
and U9114 (N_9114,N_3850,N_4189);
nor U9115 (N_9115,N_5442,N_3431);
nor U9116 (N_9116,N_4750,N_890);
and U9117 (N_9117,N_2761,N_4696);
nor U9118 (N_9118,N_3927,N_190);
and U9119 (N_9119,N_674,N_5240);
nand U9120 (N_9120,N_3357,N_4833);
or U9121 (N_9121,N_4889,N_2523);
nand U9122 (N_9122,N_5244,N_5684);
and U9123 (N_9123,N_471,N_5838);
or U9124 (N_9124,N_804,N_1772);
and U9125 (N_9125,N_4143,N_3684);
nor U9126 (N_9126,N_1703,N_3972);
or U9127 (N_9127,N_2512,N_2116);
nor U9128 (N_9128,N_711,N_5252);
or U9129 (N_9129,N_4654,N_2011);
nand U9130 (N_9130,N_5908,N_2155);
xnor U9131 (N_9131,N_5966,N_3766);
or U9132 (N_9132,N_1323,N_4390);
or U9133 (N_9133,N_1282,N_435);
and U9134 (N_9134,N_4024,N_755);
nand U9135 (N_9135,N_505,N_1441);
nor U9136 (N_9136,N_5150,N_5971);
or U9137 (N_9137,N_5065,N_5398);
nand U9138 (N_9138,N_3294,N_3681);
nand U9139 (N_9139,N_5066,N_5270);
nand U9140 (N_9140,N_2723,N_2497);
or U9141 (N_9141,N_5230,N_4723);
nor U9142 (N_9142,N_2962,N_699);
and U9143 (N_9143,N_2666,N_2681);
nor U9144 (N_9144,N_5925,N_3072);
or U9145 (N_9145,N_5753,N_2896);
or U9146 (N_9146,N_2950,N_1748);
xnor U9147 (N_9147,N_851,N_603);
or U9148 (N_9148,N_4026,N_3574);
nand U9149 (N_9149,N_3879,N_905);
and U9150 (N_9150,N_1916,N_4590);
xnor U9151 (N_9151,N_3090,N_887);
and U9152 (N_9152,N_2120,N_735);
or U9153 (N_9153,N_1731,N_3368);
nand U9154 (N_9154,N_3020,N_1788);
and U9155 (N_9155,N_4309,N_28);
nor U9156 (N_9156,N_2544,N_4684);
nor U9157 (N_9157,N_1531,N_3061);
xnor U9158 (N_9158,N_4214,N_729);
nor U9159 (N_9159,N_4125,N_299);
xnor U9160 (N_9160,N_1578,N_3647);
xnor U9161 (N_9161,N_1726,N_3519);
and U9162 (N_9162,N_5826,N_3983);
nor U9163 (N_9163,N_3949,N_2974);
and U9164 (N_9164,N_5668,N_5738);
or U9165 (N_9165,N_5269,N_2778);
and U9166 (N_9166,N_1117,N_5187);
nand U9167 (N_9167,N_3157,N_5453);
nor U9168 (N_9168,N_5348,N_501);
and U9169 (N_9169,N_5615,N_1644);
nor U9170 (N_9170,N_281,N_3540);
and U9171 (N_9171,N_1845,N_4450);
and U9172 (N_9172,N_5568,N_3362);
nor U9173 (N_9173,N_2835,N_474);
and U9174 (N_9174,N_1863,N_2907);
or U9175 (N_9175,N_2998,N_4853);
xor U9176 (N_9176,N_4287,N_2847);
or U9177 (N_9177,N_1616,N_1102);
nor U9178 (N_9178,N_4076,N_1340);
nor U9179 (N_9179,N_1457,N_4342);
or U9180 (N_9180,N_5760,N_1143);
xnor U9181 (N_9181,N_363,N_808);
and U9182 (N_9182,N_5945,N_825);
and U9183 (N_9183,N_4400,N_4928);
nor U9184 (N_9184,N_5700,N_3305);
nand U9185 (N_9185,N_1925,N_1850);
or U9186 (N_9186,N_3770,N_2475);
and U9187 (N_9187,N_3916,N_5838);
and U9188 (N_9188,N_1776,N_4833);
or U9189 (N_9189,N_197,N_1166);
nor U9190 (N_9190,N_3701,N_4428);
and U9191 (N_9191,N_1612,N_1950);
or U9192 (N_9192,N_4812,N_572);
xor U9193 (N_9193,N_5587,N_4370);
or U9194 (N_9194,N_2122,N_5699);
or U9195 (N_9195,N_4743,N_326);
or U9196 (N_9196,N_806,N_4370);
nor U9197 (N_9197,N_3874,N_633);
and U9198 (N_9198,N_5410,N_5857);
or U9199 (N_9199,N_4747,N_3354);
or U9200 (N_9200,N_984,N_5288);
nand U9201 (N_9201,N_4792,N_5370);
nand U9202 (N_9202,N_3706,N_5493);
or U9203 (N_9203,N_341,N_671);
and U9204 (N_9204,N_2567,N_930);
or U9205 (N_9205,N_2844,N_5766);
or U9206 (N_9206,N_5420,N_5824);
nor U9207 (N_9207,N_2434,N_2301);
or U9208 (N_9208,N_5913,N_1185);
and U9209 (N_9209,N_1756,N_5832);
and U9210 (N_9210,N_3667,N_476);
and U9211 (N_9211,N_2866,N_4469);
xor U9212 (N_9212,N_2366,N_2359);
nand U9213 (N_9213,N_458,N_3080);
nand U9214 (N_9214,N_4375,N_5788);
nand U9215 (N_9215,N_3650,N_1086);
or U9216 (N_9216,N_4983,N_5413);
and U9217 (N_9217,N_3566,N_4215);
xor U9218 (N_9218,N_2937,N_4704);
xnor U9219 (N_9219,N_2262,N_5720);
and U9220 (N_9220,N_5623,N_2804);
or U9221 (N_9221,N_5287,N_3590);
and U9222 (N_9222,N_2716,N_1360);
xor U9223 (N_9223,N_5437,N_4927);
or U9224 (N_9224,N_79,N_2857);
or U9225 (N_9225,N_5461,N_1575);
nand U9226 (N_9226,N_709,N_5585);
nor U9227 (N_9227,N_4997,N_4981);
nor U9228 (N_9228,N_1013,N_3194);
and U9229 (N_9229,N_4909,N_5186);
xnor U9230 (N_9230,N_5037,N_4295);
xor U9231 (N_9231,N_2148,N_260);
or U9232 (N_9232,N_262,N_5084);
xor U9233 (N_9233,N_4266,N_400);
or U9234 (N_9234,N_1710,N_133);
nand U9235 (N_9235,N_1719,N_3834);
nor U9236 (N_9236,N_5540,N_370);
or U9237 (N_9237,N_5764,N_2654);
and U9238 (N_9238,N_201,N_2469);
nand U9239 (N_9239,N_2561,N_2595);
xor U9240 (N_9240,N_1156,N_4101);
nor U9241 (N_9241,N_2046,N_3056);
nand U9242 (N_9242,N_4312,N_5860);
xor U9243 (N_9243,N_5348,N_3945);
xnor U9244 (N_9244,N_1066,N_2442);
xor U9245 (N_9245,N_2294,N_704);
or U9246 (N_9246,N_4324,N_637);
or U9247 (N_9247,N_1036,N_3187);
and U9248 (N_9248,N_3332,N_2362);
nor U9249 (N_9249,N_3186,N_2572);
nor U9250 (N_9250,N_1032,N_683);
nand U9251 (N_9251,N_1781,N_2837);
nor U9252 (N_9252,N_3968,N_4388);
or U9253 (N_9253,N_31,N_2129);
and U9254 (N_9254,N_3604,N_2829);
xnor U9255 (N_9255,N_1764,N_5959);
nor U9256 (N_9256,N_2488,N_1787);
or U9257 (N_9257,N_3519,N_1903);
nor U9258 (N_9258,N_2008,N_4546);
xor U9259 (N_9259,N_1368,N_3806);
or U9260 (N_9260,N_3715,N_1842);
xnor U9261 (N_9261,N_3852,N_3415);
or U9262 (N_9262,N_884,N_5421);
and U9263 (N_9263,N_4773,N_3648);
and U9264 (N_9264,N_3508,N_3662);
nor U9265 (N_9265,N_5734,N_101);
nand U9266 (N_9266,N_1590,N_4787);
nor U9267 (N_9267,N_3145,N_2590);
nand U9268 (N_9268,N_690,N_2265);
nand U9269 (N_9269,N_3225,N_5907);
nor U9270 (N_9270,N_5962,N_1319);
nand U9271 (N_9271,N_218,N_5586);
xor U9272 (N_9272,N_319,N_227);
nor U9273 (N_9273,N_3526,N_2852);
nand U9274 (N_9274,N_764,N_4629);
nor U9275 (N_9275,N_2965,N_1527);
or U9276 (N_9276,N_355,N_4289);
and U9277 (N_9277,N_5953,N_2917);
xor U9278 (N_9278,N_1823,N_3653);
nand U9279 (N_9279,N_5473,N_412);
or U9280 (N_9280,N_3246,N_833);
or U9281 (N_9281,N_5093,N_2120);
nand U9282 (N_9282,N_1658,N_5189);
nand U9283 (N_9283,N_1883,N_525);
and U9284 (N_9284,N_2947,N_4474);
nand U9285 (N_9285,N_1408,N_193);
or U9286 (N_9286,N_5376,N_2305);
nor U9287 (N_9287,N_909,N_1836);
nor U9288 (N_9288,N_1756,N_5250);
nor U9289 (N_9289,N_2244,N_2492);
xnor U9290 (N_9290,N_4393,N_5967);
nor U9291 (N_9291,N_5822,N_3984);
and U9292 (N_9292,N_2921,N_4937);
xor U9293 (N_9293,N_888,N_705);
or U9294 (N_9294,N_5547,N_5900);
nand U9295 (N_9295,N_4892,N_189);
nand U9296 (N_9296,N_5033,N_4310);
and U9297 (N_9297,N_200,N_1568);
or U9298 (N_9298,N_1527,N_740);
nand U9299 (N_9299,N_3000,N_1325);
xor U9300 (N_9300,N_3620,N_4411);
or U9301 (N_9301,N_860,N_5399);
nand U9302 (N_9302,N_4006,N_1556);
xnor U9303 (N_9303,N_4520,N_3073);
nand U9304 (N_9304,N_2541,N_3927);
nand U9305 (N_9305,N_4540,N_225);
xor U9306 (N_9306,N_4500,N_1279);
or U9307 (N_9307,N_1003,N_4459);
or U9308 (N_9308,N_5289,N_1607);
and U9309 (N_9309,N_1558,N_5318);
or U9310 (N_9310,N_887,N_5172);
or U9311 (N_9311,N_3147,N_1774);
or U9312 (N_9312,N_1547,N_2989);
and U9313 (N_9313,N_5058,N_5531);
and U9314 (N_9314,N_3937,N_2239);
xnor U9315 (N_9315,N_4793,N_1561);
nand U9316 (N_9316,N_499,N_500);
xnor U9317 (N_9317,N_5306,N_2);
nand U9318 (N_9318,N_4934,N_5843);
or U9319 (N_9319,N_4896,N_514);
nand U9320 (N_9320,N_4544,N_3511);
xor U9321 (N_9321,N_3618,N_4210);
nor U9322 (N_9322,N_5551,N_3399);
nor U9323 (N_9323,N_5941,N_4076);
or U9324 (N_9324,N_4816,N_2505);
xnor U9325 (N_9325,N_4643,N_3532);
and U9326 (N_9326,N_1155,N_4977);
xor U9327 (N_9327,N_674,N_3947);
nand U9328 (N_9328,N_5331,N_5240);
nand U9329 (N_9329,N_5314,N_3769);
nand U9330 (N_9330,N_2972,N_494);
xor U9331 (N_9331,N_2805,N_3632);
xnor U9332 (N_9332,N_2282,N_3043);
and U9333 (N_9333,N_3660,N_5488);
or U9334 (N_9334,N_1109,N_5058);
nand U9335 (N_9335,N_4544,N_1472);
nor U9336 (N_9336,N_4675,N_2334);
or U9337 (N_9337,N_5181,N_2902);
nand U9338 (N_9338,N_2665,N_1282);
xnor U9339 (N_9339,N_2725,N_5423);
and U9340 (N_9340,N_1109,N_5486);
nand U9341 (N_9341,N_5671,N_386);
nand U9342 (N_9342,N_181,N_3128);
and U9343 (N_9343,N_225,N_1998);
and U9344 (N_9344,N_5041,N_5799);
nand U9345 (N_9345,N_3820,N_5650);
nor U9346 (N_9346,N_2667,N_5257);
nor U9347 (N_9347,N_4289,N_568);
nor U9348 (N_9348,N_4304,N_3280);
nand U9349 (N_9349,N_2404,N_3997);
nor U9350 (N_9350,N_5868,N_274);
xnor U9351 (N_9351,N_3581,N_2288);
nor U9352 (N_9352,N_1103,N_4416);
nor U9353 (N_9353,N_1347,N_4449);
and U9354 (N_9354,N_916,N_1827);
nand U9355 (N_9355,N_2319,N_4690);
or U9356 (N_9356,N_261,N_288);
or U9357 (N_9357,N_3023,N_2631);
nand U9358 (N_9358,N_1697,N_5084);
nor U9359 (N_9359,N_2545,N_265);
nor U9360 (N_9360,N_5608,N_1615);
xor U9361 (N_9361,N_1991,N_3047);
xnor U9362 (N_9362,N_4852,N_4201);
xnor U9363 (N_9363,N_5782,N_3825);
nand U9364 (N_9364,N_5998,N_1398);
and U9365 (N_9365,N_2058,N_391);
nand U9366 (N_9366,N_1497,N_5684);
xnor U9367 (N_9367,N_2176,N_3864);
and U9368 (N_9368,N_2624,N_2256);
or U9369 (N_9369,N_3341,N_4281);
nor U9370 (N_9370,N_4250,N_645);
or U9371 (N_9371,N_2960,N_4076);
xor U9372 (N_9372,N_604,N_1144);
and U9373 (N_9373,N_3201,N_1626);
and U9374 (N_9374,N_296,N_5265);
xor U9375 (N_9375,N_2149,N_1489);
xor U9376 (N_9376,N_79,N_5187);
xor U9377 (N_9377,N_3242,N_3451);
nand U9378 (N_9378,N_2720,N_5920);
or U9379 (N_9379,N_3521,N_2511);
nand U9380 (N_9380,N_1233,N_5739);
and U9381 (N_9381,N_797,N_5628);
nand U9382 (N_9382,N_1331,N_2133);
nand U9383 (N_9383,N_1292,N_2199);
nor U9384 (N_9384,N_3281,N_4213);
and U9385 (N_9385,N_4966,N_1283);
or U9386 (N_9386,N_1010,N_3704);
nand U9387 (N_9387,N_1931,N_655);
nand U9388 (N_9388,N_4503,N_224);
nor U9389 (N_9389,N_5428,N_309);
xnor U9390 (N_9390,N_1278,N_2905);
nand U9391 (N_9391,N_4135,N_672);
nor U9392 (N_9392,N_1696,N_3056);
or U9393 (N_9393,N_2831,N_4478);
or U9394 (N_9394,N_3769,N_887);
nand U9395 (N_9395,N_1965,N_3232);
or U9396 (N_9396,N_3003,N_3060);
nand U9397 (N_9397,N_4866,N_2081);
and U9398 (N_9398,N_2527,N_4222);
or U9399 (N_9399,N_2070,N_1113);
nor U9400 (N_9400,N_5305,N_5774);
nor U9401 (N_9401,N_806,N_1710);
nor U9402 (N_9402,N_3159,N_3484);
and U9403 (N_9403,N_2077,N_1254);
or U9404 (N_9404,N_2505,N_2951);
xor U9405 (N_9405,N_1083,N_2891);
or U9406 (N_9406,N_4500,N_5715);
or U9407 (N_9407,N_2773,N_3638);
and U9408 (N_9408,N_2613,N_5680);
xor U9409 (N_9409,N_1252,N_3660);
xnor U9410 (N_9410,N_2888,N_1350);
nor U9411 (N_9411,N_1926,N_2027);
nand U9412 (N_9412,N_4865,N_5895);
and U9413 (N_9413,N_2387,N_2778);
or U9414 (N_9414,N_4162,N_5524);
and U9415 (N_9415,N_397,N_644);
xnor U9416 (N_9416,N_1527,N_2495);
or U9417 (N_9417,N_1177,N_4732);
xnor U9418 (N_9418,N_5493,N_2410);
nor U9419 (N_9419,N_595,N_1186);
or U9420 (N_9420,N_5874,N_3292);
nor U9421 (N_9421,N_2314,N_4869);
nand U9422 (N_9422,N_43,N_5138);
nor U9423 (N_9423,N_4521,N_45);
nor U9424 (N_9424,N_269,N_3689);
and U9425 (N_9425,N_955,N_4142);
xnor U9426 (N_9426,N_2949,N_5807);
xnor U9427 (N_9427,N_369,N_2592);
or U9428 (N_9428,N_3750,N_5320);
nand U9429 (N_9429,N_1780,N_701);
and U9430 (N_9430,N_2700,N_2088);
xor U9431 (N_9431,N_4757,N_1118);
xnor U9432 (N_9432,N_5167,N_212);
and U9433 (N_9433,N_1337,N_1132);
nand U9434 (N_9434,N_450,N_1898);
nor U9435 (N_9435,N_2381,N_4087);
xor U9436 (N_9436,N_5031,N_4788);
xnor U9437 (N_9437,N_1368,N_176);
xor U9438 (N_9438,N_4830,N_5038);
and U9439 (N_9439,N_706,N_2795);
nor U9440 (N_9440,N_3285,N_2383);
xnor U9441 (N_9441,N_633,N_2435);
and U9442 (N_9442,N_731,N_1581);
or U9443 (N_9443,N_35,N_3346);
or U9444 (N_9444,N_989,N_3141);
nand U9445 (N_9445,N_5036,N_1093);
and U9446 (N_9446,N_1736,N_5881);
nand U9447 (N_9447,N_195,N_4024);
nor U9448 (N_9448,N_1204,N_4946);
nand U9449 (N_9449,N_4666,N_5349);
nor U9450 (N_9450,N_4072,N_5774);
and U9451 (N_9451,N_4073,N_5504);
and U9452 (N_9452,N_2510,N_1521);
nand U9453 (N_9453,N_1725,N_3639);
or U9454 (N_9454,N_4638,N_5113);
or U9455 (N_9455,N_1399,N_1648);
nor U9456 (N_9456,N_2828,N_4315);
nand U9457 (N_9457,N_5320,N_3021);
or U9458 (N_9458,N_4795,N_4083);
nor U9459 (N_9459,N_3253,N_5994);
nor U9460 (N_9460,N_3875,N_5047);
xor U9461 (N_9461,N_544,N_3510);
or U9462 (N_9462,N_989,N_5653);
xor U9463 (N_9463,N_5690,N_5741);
nand U9464 (N_9464,N_4212,N_5985);
or U9465 (N_9465,N_3283,N_274);
or U9466 (N_9466,N_3891,N_1599);
xor U9467 (N_9467,N_4703,N_248);
nand U9468 (N_9468,N_3716,N_2544);
xor U9469 (N_9469,N_625,N_5900);
nor U9470 (N_9470,N_2060,N_2209);
xor U9471 (N_9471,N_2364,N_2975);
nand U9472 (N_9472,N_106,N_726);
or U9473 (N_9473,N_1469,N_3641);
xnor U9474 (N_9474,N_2371,N_3461);
nor U9475 (N_9475,N_3631,N_170);
nor U9476 (N_9476,N_4841,N_5583);
nand U9477 (N_9477,N_1189,N_2399);
nand U9478 (N_9478,N_1212,N_2161);
nor U9479 (N_9479,N_306,N_3333);
nor U9480 (N_9480,N_2800,N_3581);
nand U9481 (N_9481,N_5209,N_5187);
nor U9482 (N_9482,N_5929,N_1599);
and U9483 (N_9483,N_3010,N_2789);
or U9484 (N_9484,N_1672,N_1329);
xnor U9485 (N_9485,N_1695,N_1379);
or U9486 (N_9486,N_4136,N_2535);
or U9487 (N_9487,N_5591,N_1343);
nor U9488 (N_9488,N_4032,N_1100);
nor U9489 (N_9489,N_4780,N_2664);
or U9490 (N_9490,N_5569,N_1333);
nor U9491 (N_9491,N_5040,N_3602);
nor U9492 (N_9492,N_5209,N_4570);
or U9493 (N_9493,N_1913,N_1872);
nand U9494 (N_9494,N_660,N_2857);
xor U9495 (N_9495,N_62,N_261);
and U9496 (N_9496,N_3898,N_2263);
xor U9497 (N_9497,N_2574,N_3291);
xor U9498 (N_9498,N_305,N_3639);
or U9499 (N_9499,N_665,N_5961);
xnor U9500 (N_9500,N_3785,N_760);
nor U9501 (N_9501,N_2272,N_5795);
and U9502 (N_9502,N_1965,N_4041);
nand U9503 (N_9503,N_1425,N_4324);
xor U9504 (N_9504,N_5096,N_806);
nor U9505 (N_9505,N_3668,N_5208);
or U9506 (N_9506,N_2366,N_370);
xnor U9507 (N_9507,N_3132,N_3619);
or U9508 (N_9508,N_198,N_461);
nand U9509 (N_9509,N_2863,N_299);
nand U9510 (N_9510,N_3728,N_867);
nand U9511 (N_9511,N_4331,N_2511);
and U9512 (N_9512,N_4382,N_2256);
or U9513 (N_9513,N_4820,N_650);
nand U9514 (N_9514,N_4697,N_5030);
xor U9515 (N_9515,N_740,N_4965);
nand U9516 (N_9516,N_2198,N_1340);
nand U9517 (N_9517,N_930,N_4948);
or U9518 (N_9518,N_4987,N_187);
and U9519 (N_9519,N_3667,N_4561);
xnor U9520 (N_9520,N_3806,N_2965);
nor U9521 (N_9521,N_3482,N_2541);
nand U9522 (N_9522,N_4523,N_2732);
or U9523 (N_9523,N_486,N_2056);
and U9524 (N_9524,N_2919,N_4929);
xor U9525 (N_9525,N_5321,N_5988);
and U9526 (N_9526,N_3372,N_1921);
xnor U9527 (N_9527,N_5633,N_1861);
or U9528 (N_9528,N_5915,N_1436);
xnor U9529 (N_9529,N_1331,N_1026);
xor U9530 (N_9530,N_2249,N_4073);
nand U9531 (N_9531,N_5955,N_1597);
and U9532 (N_9532,N_3762,N_2341);
nor U9533 (N_9533,N_1773,N_3692);
nor U9534 (N_9534,N_3563,N_5652);
or U9535 (N_9535,N_5275,N_387);
xor U9536 (N_9536,N_4220,N_5174);
nor U9537 (N_9537,N_5225,N_1344);
and U9538 (N_9538,N_4507,N_1988);
and U9539 (N_9539,N_342,N_5083);
xnor U9540 (N_9540,N_4234,N_2497);
and U9541 (N_9541,N_2119,N_3333);
and U9542 (N_9542,N_5255,N_2667);
or U9543 (N_9543,N_2153,N_910);
nand U9544 (N_9544,N_2440,N_4249);
or U9545 (N_9545,N_5232,N_1128);
or U9546 (N_9546,N_3588,N_2689);
nor U9547 (N_9547,N_704,N_4026);
and U9548 (N_9548,N_5883,N_2060);
xor U9549 (N_9549,N_1322,N_915);
nand U9550 (N_9550,N_3443,N_1975);
nand U9551 (N_9551,N_1424,N_3433);
nand U9552 (N_9552,N_5078,N_5148);
or U9553 (N_9553,N_4692,N_3417);
nand U9554 (N_9554,N_2033,N_4370);
or U9555 (N_9555,N_5845,N_2839);
nand U9556 (N_9556,N_1667,N_3735);
and U9557 (N_9557,N_37,N_5892);
nor U9558 (N_9558,N_1045,N_3645);
nor U9559 (N_9559,N_5026,N_2394);
or U9560 (N_9560,N_4681,N_2624);
nor U9561 (N_9561,N_5145,N_380);
nor U9562 (N_9562,N_4890,N_5381);
and U9563 (N_9563,N_3295,N_4789);
or U9564 (N_9564,N_3022,N_5658);
and U9565 (N_9565,N_2488,N_3384);
and U9566 (N_9566,N_1917,N_681);
nand U9567 (N_9567,N_5734,N_2773);
and U9568 (N_9568,N_3349,N_5417);
and U9569 (N_9569,N_5040,N_5847);
nor U9570 (N_9570,N_4536,N_393);
nand U9571 (N_9571,N_4930,N_445);
and U9572 (N_9572,N_1355,N_5050);
nor U9573 (N_9573,N_188,N_3378);
xor U9574 (N_9574,N_1948,N_5671);
nand U9575 (N_9575,N_5906,N_2138);
or U9576 (N_9576,N_2983,N_75);
or U9577 (N_9577,N_4991,N_4589);
nand U9578 (N_9578,N_1817,N_1763);
nand U9579 (N_9579,N_1843,N_3077);
and U9580 (N_9580,N_5979,N_1529);
nand U9581 (N_9581,N_5223,N_2674);
nor U9582 (N_9582,N_3218,N_2530);
xnor U9583 (N_9583,N_3471,N_135);
xnor U9584 (N_9584,N_1889,N_879);
and U9585 (N_9585,N_2062,N_2627);
nand U9586 (N_9586,N_2144,N_637);
or U9587 (N_9587,N_4689,N_898);
or U9588 (N_9588,N_4738,N_4038);
nor U9589 (N_9589,N_5044,N_3571);
nand U9590 (N_9590,N_5475,N_5374);
and U9591 (N_9591,N_3053,N_499);
xnor U9592 (N_9592,N_1218,N_1304);
nand U9593 (N_9593,N_5454,N_853);
or U9594 (N_9594,N_3748,N_4127);
or U9595 (N_9595,N_5759,N_2421);
or U9596 (N_9596,N_5148,N_5109);
and U9597 (N_9597,N_573,N_3434);
or U9598 (N_9598,N_16,N_2226);
xnor U9599 (N_9599,N_3043,N_821);
and U9600 (N_9600,N_1827,N_3492);
and U9601 (N_9601,N_1511,N_1428);
nor U9602 (N_9602,N_4652,N_3822);
nand U9603 (N_9603,N_82,N_2852);
nand U9604 (N_9604,N_541,N_2162);
xnor U9605 (N_9605,N_3309,N_3230);
nand U9606 (N_9606,N_761,N_5076);
and U9607 (N_9607,N_308,N_5151);
and U9608 (N_9608,N_3,N_823);
xor U9609 (N_9609,N_627,N_4819);
nand U9610 (N_9610,N_2728,N_3971);
xnor U9611 (N_9611,N_3798,N_329);
nor U9612 (N_9612,N_2896,N_4999);
and U9613 (N_9613,N_863,N_5372);
or U9614 (N_9614,N_3123,N_2201);
or U9615 (N_9615,N_4114,N_4965);
xor U9616 (N_9616,N_2552,N_2823);
and U9617 (N_9617,N_4310,N_3835);
and U9618 (N_9618,N_4586,N_5356);
and U9619 (N_9619,N_3636,N_443);
and U9620 (N_9620,N_5480,N_4286);
and U9621 (N_9621,N_3090,N_1891);
and U9622 (N_9622,N_4167,N_111);
or U9623 (N_9623,N_2561,N_1565);
xnor U9624 (N_9624,N_5700,N_1931);
nor U9625 (N_9625,N_797,N_1240);
xor U9626 (N_9626,N_483,N_3676);
and U9627 (N_9627,N_1218,N_4750);
xor U9628 (N_9628,N_602,N_1351);
nand U9629 (N_9629,N_1138,N_1359);
nor U9630 (N_9630,N_4607,N_3549);
nand U9631 (N_9631,N_4847,N_3170);
nor U9632 (N_9632,N_2941,N_4209);
nand U9633 (N_9633,N_4593,N_4035);
xor U9634 (N_9634,N_1753,N_1086);
xnor U9635 (N_9635,N_5088,N_1270);
xnor U9636 (N_9636,N_1729,N_2166);
or U9637 (N_9637,N_1401,N_3305);
nand U9638 (N_9638,N_5596,N_1269);
and U9639 (N_9639,N_2068,N_1505);
or U9640 (N_9640,N_3760,N_5106);
xnor U9641 (N_9641,N_794,N_1086);
nand U9642 (N_9642,N_4165,N_4462);
or U9643 (N_9643,N_4020,N_4273);
nor U9644 (N_9644,N_1297,N_4884);
and U9645 (N_9645,N_2264,N_5709);
nand U9646 (N_9646,N_5432,N_3208);
and U9647 (N_9647,N_4018,N_5658);
xor U9648 (N_9648,N_4840,N_3990);
nand U9649 (N_9649,N_4794,N_942);
xnor U9650 (N_9650,N_4614,N_1769);
or U9651 (N_9651,N_3089,N_4380);
and U9652 (N_9652,N_387,N_4195);
nor U9653 (N_9653,N_3048,N_5146);
or U9654 (N_9654,N_5325,N_1380);
nand U9655 (N_9655,N_1762,N_208);
nand U9656 (N_9656,N_3764,N_2836);
nand U9657 (N_9657,N_972,N_2682);
or U9658 (N_9658,N_449,N_3925);
and U9659 (N_9659,N_5382,N_2247);
and U9660 (N_9660,N_3995,N_3702);
nand U9661 (N_9661,N_692,N_1966);
and U9662 (N_9662,N_2645,N_4807);
nor U9663 (N_9663,N_3967,N_4238);
or U9664 (N_9664,N_2554,N_5495);
or U9665 (N_9665,N_1054,N_4557);
nor U9666 (N_9666,N_1162,N_5662);
xnor U9667 (N_9667,N_5850,N_1062);
or U9668 (N_9668,N_3908,N_1122);
and U9669 (N_9669,N_3324,N_981);
xor U9670 (N_9670,N_4643,N_5033);
xnor U9671 (N_9671,N_5866,N_202);
nor U9672 (N_9672,N_66,N_3385);
or U9673 (N_9673,N_262,N_1654);
nor U9674 (N_9674,N_524,N_1600);
nand U9675 (N_9675,N_1083,N_5833);
nand U9676 (N_9676,N_1646,N_3472);
or U9677 (N_9677,N_570,N_5951);
nand U9678 (N_9678,N_3972,N_1309);
or U9679 (N_9679,N_3142,N_3951);
and U9680 (N_9680,N_300,N_1754);
nor U9681 (N_9681,N_1640,N_3251);
nand U9682 (N_9682,N_4109,N_3873);
nand U9683 (N_9683,N_3742,N_2441);
and U9684 (N_9684,N_338,N_238);
or U9685 (N_9685,N_593,N_1326);
nand U9686 (N_9686,N_5868,N_238);
or U9687 (N_9687,N_2372,N_2451);
xnor U9688 (N_9688,N_3857,N_2359);
nand U9689 (N_9689,N_736,N_5551);
xnor U9690 (N_9690,N_3826,N_3031);
xnor U9691 (N_9691,N_1037,N_3259);
nor U9692 (N_9692,N_5058,N_4487);
nand U9693 (N_9693,N_4731,N_3285);
xnor U9694 (N_9694,N_2917,N_4320);
or U9695 (N_9695,N_3823,N_5248);
xor U9696 (N_9696,N_5322,N_4330);
nor U9697 (N_9697,N_4778,N_5237);
xnor U9698 (N_9698,N_5339,N_927);
nor U9699 (N_9699,N_2692,N_384);
and U9700 (N_9700,N_4464,N_2074);
xnor U9701 (N_9701,N_5878,N_753);
nand U9702 (N_9702,N_1846,N_5797);
and U9703 (N_9703,N_959,N_1789);
and U9704 (N_9704,N_3801,N_253);
nand U9705 (N_9705,N_2289,N_599);
nor U9706 (N_9706,N_5496,N_330);
and U9707 (N_9707,N_2615,N_4202);
xor U9708 (N_9708,N_3497,N_269);
nor U9709 (N_9709,N_4377,N_2507);
or U9710 (N_9710,N_5209,N_422);
and U9711 (N_9711,N_4354,N_649);
or U9712 (N_9712,N_3216,N_978);
xor U9713 (N_9713,N_2276,N_2262);
and U9714 (N_9714,N_351,N_313);
nor U9715 (N_9715,N_4459,N_771);
nand U9716 (N_9716,N_271,N_4023);
xnor U9717 (N_9717,N_2653,N_2752);
and U9718 (N_9718,N_3054,N_2554);
nand U9719 (N_9719,N_777,N_1862);
xor U9720 (N_9720,N_275,N_1130);
and U9721 (N_9721,N_5235,N_1757);
nand U9722 (N_9722,N_810,N_723);
or U9723 (N_9723,N_2133,N_5137);
or U9724 (N_9724,N_5649,N_4038);
nand U9725 (N_9725,N_1155,N_993);
nor U9726 (N_9726,N_3226,N_870);
and U9727 (N_9727,N_1666,N_3445);
nor U9728 (N_9728,N_2164,N_4226);
nand U9729 (N_9729,N_1543,N_1358);
and U9730 (N_9730,N_499,N_2448);
or U9731 (N_9731,N_1215,N_5102);
or U9732 (N_9732,N_2161,N_5669);
and U9733 (N_9733,N_1039,N_486);
or U9734 (N_9734,N_1074,N_1141);
xnor U9735 (N_9735,N_4082,N_1107);
nand U9736 (N_9736,N_2434,N_3836);
and U9737 (N_9737,N_3931,N_5637);
and U9738 (N_9738,N_1450,N_4077);
nand U9739 (N_9739,N_5363,N_4834);
and U9740 (N_9740,N_2177,N_4683);
or U9741 (N_9741,N_4371,N_3325);
nor U9742 (N_9742,N_1305,N_3121);
or U9743 (N_9743,N_348,N_5825);
and U9744 (N_9744,N_4554,N_5564);
xnor U9745 (N_9745,N_5415,N_4477);
and U9746 (N_9746,N_5642,N_5992);
xor U9747 (N_9747,N_5350,N_1105);
nand U9748 (N_9748,N_1466,N_3963);
nor U9749 (N_9749,N_398,N_405);
nand U9750 (N_9750,N_5990,N_5994);
nand U9751 (N_9751,N_1437,N_5595);
nor U9752 (N_9752,N_5327,N_5943);
nor U9753 (N_9753,N_2573,N_761);
and U9754 (N_9754,N_2448,N_396);
nor U9755 (N_9755,N_4344,N_2468);
nand U9756 (N_9756,N_5260,N_499);
nand U9757 (N_9757,N_2228,N_1613);
and U9758 (N_9758,N_1267,N_3686);
or U9759 (N_9759,N_2114,N_1369);
nand U9760 (N_9760,N_5244,N_2628);
xor U9761 (N_9761,N_7,N_212);
xnor U9762 (N_9762,N_1327,N_5914);
or U9763 (N_9763,N_180,N_4151);
and U9764 (N_9764,N_569,N_5438);
nor U9765 (N_9765,N_1988,N_263);
xnor U9766 (N_9766,N_3448,N_5374);
xnor U9767 (N_9767,N_3353,N_2787);
or U9768 (N_9768,N_1175,N_4956);
and U9769 (N_9769,N_3211,N_4849);
nor U9770 (N_9770,N_4225,N_3977);
nand U9771 (N_9771,N_3539,N_2588);
nor U9772 (N_9772,N_3754,N_5373);
xnor U9773 (N_9773,N_5770,N_5098);
nor U9774 (N_9774,N_4380,N_5491);
xnor U9775 (N_9775,N_1354,N_1321);
nor U9776 (N_9776,N_2110,N_3178);
and U9777 (N_9777,N_5784,N_1464);
or U9778 (N_9778,N_4379,N_2577);
nand U9779 (N_9779,N_2602,N_1722);
or U9780 (N_9780,N_980,N_3077);
nand U9781 (N_9781,N_4268,N_5524);
nand U9782 (N_9782,N_3967,N_5188);
xnor U9783 (N_9783,N_5074,N_5865);
or U9784 (N_9784,N_4120,N_1030);
and U9785 (N_9785,N_149,N_4352);
xnor U9786 (N_9786,N_3241,N_4559);
xnor U9787 (N_9787,N_52,N_2897);
nand U9788 (N_9788,N_5370,N_5845);
xnor U9789 (N_9789,N_4484,N_1174);
nand U9790 (N_9790,N_1785,N_4201);
or U9791 (N_9791,N_2054,N_5493);
and U9792 (N_9792,N_3381,N_5595);
nor U9793 (N_9793,N_4995,N_1326);
xnor U9794 (N_9794,N_4879,N_3260);
and U9795 (N_9795,N_3712,N_1261);
nand U9796 (N_9796,N_3011,N_1538);
and U9797 (N_9797,N_5300,N_4942);
or U9798 (N_9798,N_5527,N_4101);
nand U9799 (N_9799,N_618,N_3149);
xnor U9800 (N_9800,N_3486,N_2484);
xor U9801 (N_9801,N_4977,N_771);
xnor U9802 (N_9802,N_1991,N_2022);
and U9803 (N_9803,N_4103,N_4612);
and U9804 (N_9804,N_4691,N_5247);
nand U9805 (N_9805,N_4919,N_2038);
and U9806 (N_9806,N_5785,N_3417);
xnor U9807 (N_9807,N_712,N_4029);
xor U9808 (N_9808,N_4058,N_5123);
and U9809 (N_9809,N_298,N_5831);
and U9810 (N_9810,N_5452,N_5026);
or U9811 (N_9811,N_4750,N_2857);
or U9812 (N_9812,N_2384,N_4633);
and U9813 (N_9813,N_3933,N_5456);
or U9814 (N_9814,N_2789,N_5105);
or U9815 (N_9815,N_305,N_5636);
xnor U9816 (N_9816,N_3388,N_3907);
or U9817 (N_9817,N_4763,N_1768);
and U9818 (N_9818,N_4974,N_2606);
and U9819 (N_9819,N_3111,N_3816);
or U9820 (N_9820,N_2719,N_4471);
nor U9821 (N_9821,N_469,N_4028);
nand U9822 (N_9822,N_2639,N_4684);
nor U9823 (N_9823,N_1790,N_4434);
or U9824 (N_9824,N_4447,N_275);
nor U9825 (N_9825,N_300,N_3039);
and U9826 (N_9826,N_2022,N_3304);
and U9827 (N_9827,N_919,N_1818);
nor U9828 (N_9828,N_723,N_3685);
nand U9829 (N_9829,N_2624,N_2155);
nor U9830 (N_9830,N_4340,N_4537);
and U9831 (N_9831,N_4288,N_2585);
and U9832 (N_9832,N_4027,N_1588);
or U9833 (N_9833,N_4935,N_3305);
nand U9834 (N_9834,N_5960,N_1837);
or U9835 (N_9835,N_4549,N_3968);
nor U9836 (N_9836,N_1058,N_4751);
and U9837 (N_9837,N_2526,N_2507);
and U9838 (N_9838,N_5286,N_5977);
nor U9839 (N_9839,N_4637,N_1703);
xnor U9840 (N_9840,N_1866,N_2648);
nor U9841 (N_9841,N_4056,N_5925);
nor U9842 (N_9842,N_1926,N_5802);
and U9843 (N_9843,N_1682,N_5658);
xnor U9844 (N_9844,N_1466,N_4308);
and U9845 (N_9845,N_4606,N_4830);
nand U9846 (N_9846,N_916,N_74);
or U9847 (N_9847,N_2823,N_331);
xnor U9848 (N_9848,N_1497,N_2257);
and U9849 (N_9849,N_5550,N_4817);
nand U9850 (N_9850,N_3708,N_4961);
nor U9851 (N_9851,N_1461,N_957);
nand U9852 (N_9852,N_4599,N_721);
xnor U9853 (N_9853,N_2541,N_4301);
or U9854 (N_9854,N_5196,N_4938);
nor U9855 (N_9855,N_2277,N_3719);
or U9856 (N_9856,N_3049,N_3395);
nand U9857 (N_9857,N_1971,N_3773);
and U9858 (N_9858,N_753,N_5626);
and U9859 (N_9859,N_1220,N_5789);
nor U9860 (N_9860,N_5969,N_2145);
nor U9861 (N_9861,N_4606,N_2088);
xnor U9862 (N_9862,N_4787,N_4896);
nand U9863 (N_9863,N_2001,N_120);
or U9864 (N_9864,N_5729,N_3821);
xor U9865 (N_9865,N_5596,N_322);
xor U9866 (N_9866,N_1165,N_3255);
or U9867 (N_9867,N_4137,N_3989);
and U9868 (N_9868,N_4257,N_5182);
and U9869 (N_9869,N_4554,N_156);
and U9870 (N_9870,N_2430,N_3245);
nand U9871 (N_9871,N_5039,N_4152);
and U9872 (N_9872,N_3582,N_5760);
and U9873 (N_9873,N_5759,N_4979);
nor U9874 (N_9874,N_5857,N_126);
xnor U9875 (N_9875,N_5391,N_2181);
nand U9876 (N_9876,N_2444,N_1922);
nand U9877 (N_9877,N_3823,N_2477);
nand U9878 (N_9878,N_84,N_1103);
xnor U9879 (N_9879,N_10,N_4131);
or U9880 (N_9880,N_5352,N_1387);
nor U9881 (N_9881,N_4306,N_2150);
xor U9882 (N_9882,N_4672,N_651);
or U9883 (N_9883,N_3169,N_3034);
nor U9884 (N_9884,N_1556,N_3045);
nand U9885 (N_9885,N_3987,N_4787);
and U9886 (N_9886,N_671,N_4978);
or U9887 (N_9887,N_5650,N_4698);
or U9888 (N_9888,N_2103,N_1570);
nor U9889 (N_9889,N_5071,N_2005);
nor U9890 (N_9890,N_2522,N_2808);
nor U9891 (N_9891,N_4199,N_3575);
nand U9892 (N_9892,N_1786,N_5310);
xnor U9893 (N_9893,N_4393,N_3770);
nor U9894 (N_9894,N_2855,N_3583);
nand U9895 (N_9895,N_3195,N_5575);
or U9896 (N_9896,N_2362,N_4798);
xor U9897 (N_9897,N_1496,N_3732);
xor U9898 (N_9898,N_4119,N_2026);
nor U9899 (N_9899,N_3955,N_755);
nor U9900 (N_9900,N_3925,N_2661);
or U9901 (N_9901,N_4656,N_3498);
or U9902 (N_9902,N_1242,N_4286);
xnor U9903 (N_9903,N_1334,N_4203);
xor U9904 (N_9904,N_5650,N_3627);
and U9905 (N_9905,N_2463,N_3026);
nand U9906 (N_9906,N_4007,N_1448);
and U9907 (N_9907,N_1150,N_1821);
or U9908 (N_9908,N_5060,N_2947);
nand U9909 (N_9909,N_3870,N_4869);
xor U9910 (N_9910,N_1437,N_3218);
xor U9911 (N_9911,N_1866,N_1369);
xnor U9912 (N_9912,N_4613,N_3430);
and U9913 (N_9913,N_3328,N_5355);
nor U9914 (N_9914,N_548,N_1926);
xnor U9915 (N_9915,N_5212,N_598);
nand U9916 (N_9916,N_2577,N_5713);
or U9917 (N_9917,N_4158,N_5925);
or U9918 (N_9918,N_4104,N_3404);
nor U9919 (N_9919,N_2567,N_726);
nand U9920 (N_9920,N_3390,N_2969);
xor U9921 (N_9921,N_360,N_5835);
nor U9922 (N_9922,N_1475,N_3571);
nor U9923 (N_9923,N_3383,N_524);
nor U9924 (N_9924,N_4315,N_5016);
nor U9925 (N_9925,N_974,N_4175);
nand U9926 (N_9926,N_374,N_534);
or U9927 (N_9927,N_5355,N_3406);
and U9928 (N_9928,N_1445,N_481);
or U9929 (N_9929,N_5984,N_3738);
or U9930 (N_9930,N_749,N_3483);
xnor U9931 (N_9931,N_5758,N_2353);
nand U9932 (N_9932,N_1953,N_4361);
or U9933 (N_9933,N_958,N_470);
or U9934 (N_9934,N_4927,N_1933);
or U9935 (N_9935,N_2430,N_5835);
and U9936 (N_9936,N_4570,N_3664);
or U9937 (N_9937,N_2714,N_5965);
nand U9938 (N_9938,N_5901,N_2401);
and U9939 (N_9939,N_1544,N_2223);
xor U9940 (N_9940,N_2041,N_4587);
xnor U9941 (N_9941,N_1835,N_2548);
or U9942 (N_9942,N_3141,N_4309);
nand U9943 (N_9943,N_2846,N_856);
and U9944 (N_9944,N_1172,N_5843);
nor U9945 (N_9945,N_1991,N_667);
or U9946 (N_9946,N_718,N_4445);
and U9947 (N_9947,N_3836,N_3037);
and U9948 (N_9948,N_1660,N_3280);
xor U9949 (N_9949,N_939,N_4317);
xnor U9950 (N_9950,N_203,N_817);
xnor U9951 (N_9951,N_4607,N_3811);
or U9952 (N_9952,N_5404,N_2394);
nor U9953 (N_9953,N_4694,N_4319);
nor U9954 (N_9954,N_3358,N_1620);
nand U9955 (N_9955,N_2032,N_4633);
nor U9956 (N_9956,N_1474,N_2493);
nand U9957 (N_9957,N_3764,N_2625);
nor U9958 (N_9958,N_4285,N_4282);
nand U9959 (N_9959,N_2110,N_1604);
nand U9960 (N_9960,N_3374,N_5173);
and U9961 (N_9961,N_1175,N_1017);
and U9962 (N_9962,N_3403,N_3833);
xor U9963 (N_9963,N_5267,N_218);
nor U9964 (N_9964,N_257,N_647);
nand U9965 (N_9965,N_4986,N_525);
nand U9966 (N_9966,N_3536,N_3074);
xnor U9967 (N_9967,N_5506,N_3919);
xor U9968 (N_9968,N_2065,N_281);
and U9969 (N_9969,N_5003,N_4673);
nor U9970 (N_9970,N_2844,N_3946);
nand U9971 (N_9971,N_2980,N_3616);
or U9972 (N_9972,N_2977,N_5885);
nor U9973 (N_9973,N_5307,N_298);
xor U9974 (N_9974,N_444,N_3095);
nor U9975 (N_9975,N_5355,N_338);
or U9976 (N_9976,N_479,N_2440);
or U9977 (N_9977,N_2583,N_2004);
nor U9978 (N_9978,N_20,N_292);
nor U9979 (N_9979,N_3570,N_1012);
nor U9980 (N_9980,N_5182,N_5628);
and U9981 (N_9981,N_2803,N_4547);
nor U9982 (N_9982,N_5527,N_3256);
and U9983 (N_9983,N_3410,N_2845);
or U9984 (N_9984,N_4848,N_292);
nor U9985 (N_9985,N_3282,N_2336);
or U9986 (N_9986,N_3015,N_5652);
nor U9987 (N_9987,N_2999,N_1135);
or U9988 (N_9988,N_2849,N_2480);
nand U9989 (N_9989,N_310,N_2442);
xnor U9990 (N_9990,N_5351,N_2918);
and U9991 (N_9991,N_3351,N_647);
nor U9992 (N_9992,N_448,N_4683);
nand U9993 (N_9993,N_1088,N_4269);
nand U9994 (N_9994,N_3376,N_1029);
nand U9995 (N_9995,N_2447,N_5532);
or U9996 (N_9996,N_5743,N_4770);
nor U9997 (N_9997,N_1295,N_975);
nor U9998 (N_9998,N_2466,N_5638);
and U9999 (N_9999,N_2400,N_3469);
or U10000 (N_10000,N_2348,N_247);
nor U10001 (N_10001,N_518,N_922);
or U10002 (N_10002,N_3353,N_2298);
and U10003 (N_10003,N_2726,N_4663);
or U10004 (N_10004,N_5259,N_786);
nand U10005 (N_10005,N_2776,N_5307);
nor U10006 (N_10006,N_5631,N_956);
nor U10007 (N_10007,N_5771,N_2305);
and U10008 (N_10008,N_2371,N_224);
nor U10009 (N_10009,N_3775,N_3480);
xnor U10010 (N_10010,N_2303,N_3139);
or U10011 (N_10011,N_3652,N_5776);
and U10012 (N_10012,N_4179,N_3161);
or U10013 (N_10013,N_5371,N_4009);
and U10014 (N_10014,N_1571,N_5649);
xnor U10015 (N_10015,N_1473,N_1110);
nand U10016 (N_10016,N_2606,N_462);
nand U10017 (N_10017,N_2421,N_1661);
xor U10018 (N_10018,N_593,N_4867);
or U10019 (N_10019,N_461,N_4893);
or U10020 (N_10020,N_3598,N_1013);
nor U10021 (N_10021,N_761,N_3800);
and U10022 (N_10022,N_5181,N_5028);
and U10023 (N_10023,N_1179,N_1349);
or U10024 (N_10024,N_4067,N_5199);
or U10025 (N_10025,N_1468,N_3994);
nand U10026 (N_10026,N_4903,N_5113);
nor U10027 (N_10027,N_4933,N_581);
xor U10028 (N_10028,N_3530,N_2243);
nor U10029 (N_10029,N_1978,N_1848);
nand U10030 (N_10030,N_2227,N_2842);
nor U10031 (N_10031,N_2371,N_279);
or U10032 (N_10032,N_3506,N_1162);
and U10033 (N_10033,N_2145,N_1894);
xnor U10034 (N_10034,N_1139,N_262);
nand U10035 (N_10035,N_4867,N_2317);
or U10036 (N_10036,N_5327,N_2707);
nand U10037 (N_10037,N_4403,N_1383);
and U10038 (N_10038,N_3438,N_306);
and U10039 (N_10039,N_5652,N_3842);
nand U10040 (N_10040,N_5588,N_3476);
nand U10041 (N_10041,N_2882,N_4264);
nand U10042 (N_10042,N_3946,N_4127);
xor U10043 (N_10043,N_1120,N_1844);
nand U10044 (N_10044,N_1634,N_1319);
nor U10045 (N_10045,N_3477,N_365);
or U10046 (N_10046,N_846,N_5571);
nand U10047 (N_10047,N_3906,N_4515);
nor U10048 (N_10048,N_734,N_5943);
nand U10049 (N_10049,N_3913,N_4732);
nor U10050 (N_10050,N_5410,N_5315);
and U10051 (N_10051,N_2762,N_1406);
or U10052 (N_10052,N_1979,N_5377);
and U10053 (N_10053,N_3481,N_1676);
nand U10054 (N_10054,N_3947,N_3787);
xor U10055 (N_10055,N_5898,N_1719);
or U10056 (N_10056,N_4508,N_3427);
nand U10057 (N_10057,N_2764,N_4344);
nand U10058 (N_10058,N_1693,N_295);
xor U10059 (N_10059,N_1560,N_428);
nor U10060 (N_10060,N_664,N_1352);
xor U10061 (N_10061,N_529,N_5481);
or U10062 (N_10062,N_224,N_1688);
and U10063 (N_10063,N_5502,N_2004);
and U10064 (N_10064,N_4210,N_5881);
xnor U10065 (N_10065,N_1643,N_3452);
xor U10066 (N_10066,N_5624,N_1349);
xor U10067 (N_10067,N_4091,N_307);
and U10068 (N_10068,N_5231,N_3556);
and U10069 (N_10069,N_276,N_3451);
nand U10070 (N_10070,N_2470,N_3775);
nand U10071 (N_10071,N_4330,N_5874);
nor U10072 (N_10072,N_1320,N_101);
nor U10073 (N_10073,N_2392,N_1773);
nand U10074 (N_10074,N_89,N_4779);
nand U10075 (N_10075,N_3463,N_3839);
or U10076 (N_10076,N_1618,N_1751);
xnor U10077 (N_10077,N_2233,N_1983);
or U10078 (N_10078,N_217,N_3284);
nand U10079 (N_10079,N_211,N_5939);
and U10080 (N_10080,N_2172,N_4954);
or U10081 (N_10081,N_227,N_1432);
nand U10082 (N_10082,N_3939,N_1593);
xnor U10083 (N_10083,N_5927,N_1549);
and U10084 (N_10084,N_2594,N_197);
nand U10085 (N_10085,N_5118,N_1806);
or U10086 (N_10086,N_3517,N_5718);
or U10087 (N_10087,N_3450,N_2683);
xnor U10088 (N_10088,N_5651,N_3371);
nor U10089 (N_10089,N_4837,N_2190);
xor U10090 (N_10090,N_3274,N_1951);
nor U10091 (N_10091,N_5978,N_3000);
nand U10092 (N_10092,N_3557,N_2730);
xor U10093 (N_10093,N_4939,N_2222);
and U10094 (N_10094,N_2377,N_5522);
xnor U10095 (N_10095,N_5239,N_3305);
xor U10096 (N_10096,N_1268,N_4278);
nand U10097 (N_10097,N_4340,N_5600);
nand U10098 (N_10098,N_5849,N_5933);
xor U10099 (N_10099,N_3930,N_713);
and U10100 (N_10100,N_3014,N_3524);
or U10101 (N_10101,N_3330,N_5454);
nor U10102 (N_10102,N_2041,N_2383);
nand U10103 (N_10103,N_4888,N_1457);
nor U10104 (N_10104,N_3301,N_4738);
and U10105 (N_10105,N_5131,N_2219);
nand U10106 (N_10106,N_852,N_4527);
nand U10107 (N_10107,N_1732,N_2809);
or U10108 (N_10108,N_5971,N_4902);
or U10109 (N_10109,N_7,N_4904);
and U10110 (N_10110,N_3097,N_4021);
xnor U10111 (N_10111,N_837,N_3338);
xnor U10112 (N_10112,N_263,N_3175);
xnor U10113 (N_10113,N_1660,N_2009);
and U10114 (N_10114,N_3391,N_3525);
nand U10115 (N_10115,N_1654,N_4933);
nor U10116 (N_10116,N_5240,N_2537);
and U10117 (N_10117,N_1287,N_2805);
and U10118 (N_10118,N_3170,N_1488);
and U10119 (N_10119,N_1606,N_5458);
and U10120 (N_10120,N_2248,N_5347);
nor U10121 (N_10121,N_2556,N_4749);
or U10122 (N_10122,N_3931,N_2759);
or U10123 (N_10123,N_5403,N_2776);
and U10124 (N_10124,N_5359,N_4014);
nand U10125 (N_10125,N_2798,N_2477);
xnor U10126 (N_10126,N_1338,N_3768);
xnor U10127 (N_10127,N_2132,N_1689);
and U10128 (N_10128,N_1168,N_5970);
nor U10129 (N_10129,N_1849,N_3318);
and U10130 (N_10130,N_1087,N_1419);
nand U10131 (N_10131,N_1066,N_5498);
xnor U10132 (N_10132,N_4388,N_1566);
and U10133 (N_10133,N_787,N_4493);
and U10134 (N_10134,N_3358,N_2169);
xnor U10135 (N_10135,N_2110,N_2557);
nor U10136 (N_10136,N_1406,N_5006);
or U10137 (N_10137,N_5249,N_1300);
or U10138 (N_10138,N_3076,N_1820);
nor U10139 (N_10139,N_5662,N_1746);
xor U10140 (N_10140,N_4128,N_4989);
nand U10141 (N_10141,N_2260,N_1805);
and U10142 (N_10142,N_1943,N_5608);
or U10143 (N_10143,N_5047,N_3242);
or U10144 (N_10144,N_583,N_2300);
nor U10145 (N_10145,N_5808,N_1957);
nor U10146 (N_10146,N_4950,N_5305);
and U10147 (N_10147,N_1394,N_2315);
nand U10148 (N_10148,N_4040,N_1985);
nor U10149 (N_10149,N_1735,N_5362);
and U10150 (N_10150,N_1956,N_4119);
nor U10151 (N_10151,N_961,N_3772);
xnor U10152 (N_10152,N_4415,N_4560);
xnor U10153 (N_10153,N_4063,N_767);
nand U10154 (N_10154,N_2946,N_1679);
and U10155 (N_10155,N_827,N_4539);
nand U10156 (N_10156,N_1649,N_4288);
or U10157 (N_10157,N_2896,N_3949);
and U10158 (N_10158,N_2971,N_2491);
nand U10159 (N_10159,N_1647,N_5282);
and U10160 (N_10160,N_910,N_2868);
and U10161 (N_10161,N_3966,N_4934);
xnor U10162 (N_10162,N_4928,N_4917);
and U10163 (N_10163,N_873,N_4377);
and U10164 (N_10164,N_2241,N_431);
nand U10165 (N_10165,N_5640,N_2764);
xor U10166 (N_10166,N_1785,N_822);
nand U10167 (N_10167,N_2317,N_1302);
and U10168 (N_10168,N_5221,N_2075);
or U10169 (N_10169,N_1654,N_2289);
or U10170 (N_10170,N_4089,N_968);
nor U10171 (N_10171,N_396,N_5354);
and U10172 (N_10172,N_5442,N_3148);
nor U10173 (N_10173,N_5931,N_527);
nand U10174 (N_10174,N_2586,N_4049);
and U10175 (N_10175,N_2905,N_5855);
or U10176 (N_10176,N_5742,N_4030);
nor U10177 (N_10177,N_4220,N_4816);
nand U10178 (N_10178,N_4653,N_5283);
and U10179 (N_10179,N_1782,N_302);
or U10180 (N_10180,N_5754,N_5054);
nor U10181 (N_10181,N_345,N_4808);
nand U10182 (N_10182,N_5599,N_2348);
or U10183 (N_10183,N_1006,N_4235);
and U10184 (N_10184,N_5280,N_3463);
and U10185 (N_10185,N_2696,N_2809);
or U10186 (N_10186,N_2023,N_1173);
nor U10187 (N_10187,N_442,N_1878);
and U10188 (N_10188,N_4292,N_4691);
and U10189 (N_10189,N_5045,N_5925);
nor U10190 (N_10190,N_3565,N_3239);
or U10191 (N_10191,N_5712,N_4107);
and U10192 (N_10192,N_4264,N_5333);
or U10193 (N_10193,N_2644,N_5691);
and U10194 (N_10194,N_3564,N_4794);
nand U10195 (N_10195,N_4735,N_1350);
nand U10196 (N_10196,N_802,N_1626);
xnor U10197 (N_10197,N_1629,N_969);
and U10198 (N_10198,N_2368,N_1202);
or U10199 (N_10199,N_5371,N_4891);
nand U10200 (N_10200,N_98,N_1537);
and U10201 (N_10201,N_2818,N_5340);
nand U10202 (N_10202,N_5381,N_2814);
nand U10203 (N_10203,N_440,N_3120);
nand U10204 (N_10204,N_1298,N_949);
xor U10205 (N_10205,N_4055,N_1116);
nor U10206 (N_10206,N_2485,N_5891);
and U10207 (N_10207,N_658,N_5433);
and U10208 (N_10208,N_5387,N_265);
xnor U10209 (N_10209,N_3571,N_5352);
nand U10210 (N_10210,N_4908,N_2900);
or U10211 (N_10211,N_5263,N_5519);
nand U10212 (N_10212,N_2406,N_1436);
or U10213 (N_10213,N_2131,N_5978);
nand U10214 (N_10214,N_236,N_3213);
xnor U10215 (N_10215,N_3751,N_3731);
nor U10216 (N_10216,N_1590,N_74);
or U10217 (N_10217,N_5839,N_5712);
nand U10218 (N_10218,N_5684,N_5224);
and U10219 (N_10219,N_771,N_1227);
xnor U10220 (N_10220,N_1284,N_1396);
nor U10221 (N_10221,N_2655,N_4499);
nand U10222 (N_10222,N_1642,N_455);
and U10223 (N_10223,N_2337,N_4325);
and U10224 (N_10224,N_5649,N_5499);
or U10225 (N_10225,N_2744,N_3112);
nand U10226 (N_10226,N_5039,N_3849);
nand U10227 (N_10227,N_4823,N_2120);
nor U10228 (N_10228,N_1388,N_3644);
and U10229 (N_10229,N_1718,N_3456);
xnor U10230 (N_10230,N_5275,N_4739);
nand U10231 (N_10231,N_3947,N_5466);
xnor U10232 (N_10232,N_5385,N_5432);
nor U10233 (N_10233,N_5949,N_4083);
and U10234 (N_10234,N_4848,N_3971);
nand U10235 (N_10235,N_1279,N_4186);
nand U10236 (N_10236,N_3938,N_4712);
and U10237 (N_10237,N_446,N_1561);
nor U10238 (N_10238,N_267,N_3016);
nor U10239 (N_10239,N_751,N_2991);
nand U10240 (N_10240,N_3335,N_5744);
and U10241 (N_10241,N_991,N_1691);
xnor U10242 (N_10242,N_3135,N_1438);
xor U10243 (N_10243,N_3252,N_2496);
xnor U10244 (N_10244,N_4628,N_5579);
nand U10245 (N_10245,N_2837,N_4919);
nor U10246 (N_10246,N_1669,N_5501);
and U10247 (N_10247,N_921,N_4512);
xor U10248 (N_10248,N_4345,N_5074);
nor U10249 (N_10249,N_5194,N_2594);
nor U10250 (N_10250,N_3239,N_4638);
nor U10251 (N_10251,N_1366,N_1042);
nor U10252 (N_10252,N_38,N_5541);
and U10253 (N_10253,N_5126,N_3951);
nand U10254 (N_10254,N_940,N_4349);
nand U10255 (N_10255,N_2356,N_1654);
or U10256 (N_10256,N_2958,N_3061);
nor U10257 (N_10257,N_996,N_3970);
and U10258 (N_10258,N_4756,N_4842);
or U10259 (N_10259,N_1071,N_5484);
nand U10260 (N_10260,N_2346,N_5505);
or U10261 (N_10261,N_5334,N_895);
nor U10262 (N_10262,N_4620,N_3305);
nand U10263 (N_10263,N_4145,N_2855);
and U10264 (N_10264,N_2474,N_3834);
nor U10265 (N_10265,N_3014,N_5093);
xor U10266 (N_10266,N_2668,N_4252);
xnor U10267 (N_10267,N_1351,N_352);
nand U10268 (N_10268,N_710,N_4897);
or U10269 (N_10269,N_4241,N_4110);
and U10270 (N_10270,N_82,N_1576);
nor U10271 (N_10271,N_2629,N_1297);
or U10272 (N_10272,N_2150,N_4895);
xor U10273 (N_10273,N_3822,N_4725);
or U10274 (N_10274,N_2106,N_5322);
or U10275 (N_10275,N_2571,N_5222);
nand U10276 (N_10276,N_3475,N_1698);
or U10277 (N_10277,N_5868,N_3304);
nor U10278 (N_10278,N_2846,N_5470);
nand U10279 (N_10279,N_8,N_2919);
nor U10280 (N_10280,N_3988,N_3168);
or U10281 (N_10281,N_4285,N_387);
xnor U10282 (N_10282,N_5198,N_4698);
xnor U10283 (N_10283,N_5595,N_361);
xor U10284 (N_10284,N_2502,N_4723);
and U10285 (N_10285,N_2614,N_2922);
nor U10286 (N_10286,N_595,N_1135);
xor U10287 (N_10287,N_1260,N_20);
nor U10288 (N_10288,N_385,N_4560);
or U10289 (N_10289,N_1146,N_2495);
nor U10290 (N_10290,N_111,N_236);
or U10291 (N_10291,N_1225,N_3528);
xor U10292 (N_10292,N_2790,N_4986);
xnor U10293 (N_10293,N_1947,N_5974);
and U10294 (N_10294,N_565,N_5530);
nor U10295 (N_10295,N_2562,N_4264);
or U10296 (N_10296,N_5729,N_2386);
or U10297 (N_10297,N_2400,N_4931);
nor U10298 (N_10298,N_541,N_4181);
nand U10299 (N_10299,N_1839,N_5475);
and U10300 (N_10300,N_2534,N_2207);
xnor U10301 (N_10301,N_4069,N_2514);
xor U10302 (N_10302,N_1391,N_170);
nand U10303 (N_10303,N_1098,N_2319);
nor U10304 (N_10304,N_5067,N_4143);
or U10305 (N_10305,N_1837,N_4016);
nand U10306 (N_10306,N_43,N_2619);
nor U10307 (N_10307,N_3568,N_3851);
nor U10308 (N_10308,N_521,N_5768);
xor U10309 (N_10309,N_5395,N_2132);
or U10310 (N_10310,N_2116,N_5101);
or U10311 (N_10311,N_3746,N_1731);
xnor U10312 (N_10312,N_4783,N_2990);
nor U10313 (N_10313,N_5651,N_1398);
nor U10314 (N_10314,N_5678,N_1361);
nor U10315 (N_10315,N_2292,N_4466);
nand U10316 (N_10316,N_3530,N_5278);
or U10317 (N_10317,N_1066,N_3276);
and U10318 (N_10318,N_2643,N_5557);
nand U10319 (N_10319,N_560,N_5388);
nor U10320 (N_10320,N_5203,N_1453);
nor U10321 (N_10321,N_139,N_204);
and U10322 (N_10322,N_1034,N_214);
nor U10323 (N_10323,N_1631,N_857);
or U10324 (N_10324,N_3830,N_2420);
nand U10325 (N_10325,N_1027,N_1644);
nand U10326 (N_10326,N_3111,N_2663);
and U10327 (N_10327,N_3790,N_5613);
nand U10328 (N_10328,N_421,N_4606);
nand U10329 (N_10329,N_4998,N_66);
xnor U10330 (N_10330,N_4106,N_2755);
xor U10331 (N_10331,N_4564,N_5651);
or U10332 (N_10332,N_9,N_3073);
xor U10333 (N_10333,N_4571,N_1622);
nand U10334 (N_10334,N_4441,N_3998);
or U10335 (N_10335,N_1831,N_2541);
nor U10336 (N_10336,N_5444,N_4112);
or U10337 (N_10337,N_3553,N_3405);
and U10338 (N_10338,N_4956,N_1660);
nor U10339 (N_10339,N_1464,N_4452);
xnor U10340 (N_10340,N_4415,N_1202);
nand U10341 (N_10341,N_5411,N_3270);
and U10342 (N_10342,N_1133,N_243);
and U10343 (N_10343,N_140,N_569);
nand U10344 (N_10344,N_2901,N_5881);
xnor U10345 (N_10345,N_213,N_5316);
xnor U10346 (N_10346,N_5981,N_2844);
and U10347 (N_10347,N_4950,N_5550);
and U10348 (N_10348,N_5513,N_945);
nor U10349 (N_10349,N_4599,N_4429);
or U10350 (N_10350,N_1267,N_1700);
xnor U10351 (N_10351,N_605,N_3663);
nor U10352 (N_10352,N_2360,N_2718);
xnor U10353 (N_10353,N_2451,N_2063);
nor U10354 (N_10354,N_4798,N_3037);
nor U10355 (N_10355,N_3208,N_1343);
nand U10356 (N_10356,N_1415,N_1256);
nor U10357 (N_10357,N_2694,N_424);
and U10358 (N_10358,N_1656,N_278);
nor U10359 (N_10359,N_1875,N_2328);
xor U10360 (N_10360,N_3117,N_47);
nand U10361 (N_10361,N_2332,N_2559);
nand U10362 (N_10362,N_4212,N_5043);
nand U10363 (N_10363,N_624,N_983);
nor U10364 (N_10364,N_2476,N_1528);
or U10365 (N_10365,N_385,N_3921);
nor U10366 (N_10366,N_3742,N_3924);
or U10367 (N_10367,N_4812,N_1412);
nand U10368 (N_10368,N_4616,N_2330);
xor U10369 (N_10369,N_4550,N_2184);
or U10370 (N_10370,N_2845,N_1532);
nand U10371 (N_10371,N_3287,N_2581);
nand U10372 (N_10372,N_3874,N_3818);
xor U10373 (N_10373,N_1437,N_3329);
nor U10374 (N_10374,N_4129,N_1881);
or U10375 (N_10375,N_3403,N_1191);
or U10376 (N_10376,N_3751,N_4460);
or U10377 (N_10377,N_3845,N_642);
xnor U10378 (N_10378,N_3702,N_5935);
and U10379 (N_10379,N_5764,N_5124);
or U10380 (N_10380,N_1497,N_4828);
nand U10381 (N_10381,N_848,N_2759);
and U10382 (N_10382,N_5896,N_1887);
nand U10383 (N_10383,N_2315,N_5541);
xnor U10384 (N_10384,N_2846,N_3941);
and U10385 (N_10385,N_5590,N_1711);
and U10386 (N_10386,N_301,N_2023);
and U10387 (N_10387,N_41,N_3384);
nand U10388 (N_10388,N_4782,N_3457);
xor U10389 (N_10389,N_2964,N_3915);
or U10390 (N_10390,N_4405,N_1826);
and U10391 (N_10391,N_978,N_1470);
and U10392 (N_10392,N_804,N_5402);
or U10393 (N_10393,N_1547,N_699);
or U10394 (N_10394,N_103,N_5757);
or U10395 (N_10395,N_4509,N_2390);
xnor U10396 (N_10396,N_975,N_4437);
xnor U10397 (N_10397,N_3366,N_1967);
and U10398 (N_10398,N_1549,N_2107);
and U10399 (N_10399,N_4460,N_135);
nor U10400 (N_10400,N_3595,N_3759);
nor U10401 (N_10401,N_3986,N_3669);
nand U10402 (N_10402,N_1215,N_1867);
nor U10403 (N_10403,N_1163,N_5899);
or U10404 (N_10404,N_736,N_641);
nor U10405 (N_10405,N_1579,N_2054);
nor U10406 (N_10406,N_5944,N_2035);
nor U10407 (N_10407,N_337,N_1439);
and U10408 (N_10408,N_5977,N_736);
xor U10409 (N_10409,N_4780,N_5625);
nor U10410 (N_10410,N_3202,N_878);
xnor U10411 (N_10411,N_5834,N_3320);
xor U10412 (N_10412,N_1656,N_646);
and U10413 (N_10413,N_19,N_5900);
xnor U10414 (N_10414,N_1493,N_3373);
nand U10415 (N_10415,N_38,N_5955);
and U10416 (N_10416,N_4733,N_1298);
xnor U10417 (N_10417,N_5697,N_169);
xor U10418 (N_10418,N_1438,N_292);
nand U10419 (N_10419,N_1376,N_374);
or U10420 (N_10420,N_3617,N_696);
and U10421 (N_10421,N_5976,N_2069);
xnor U10422 (N_10422,N_2209,N_1521);
nor U10423 (N_10423,N_2138,N_1935);
nand U10424 (N_10424,N_2296,N_1115);
or U10425 (N_10425,N_3934,N_188);
or U10426 (N_10426,N_4472,N_2265);
xnor U10427 (N_10427,N_3600,N_2054);
or U10428 (N_10428,N_3403,N_3813);
xor U10429 (N_10429,N_2298,N_3674);
nor U10430 (N_10430,N_1731,N_5214);
and U10431 (N_10431,N_2949,N_1945);
and U10432 (N_10432,N_4633,N_825);
and U10433 (N_10433,N_5837,N_4258);
xnor U10434 (N_10434,N_5916,N_5518);
nor U10435 (N_10435,N_4468,N_509);
xor U10436 (N_10436,N_2661,N_3018);
nand U10437 (N_10437,N_4411,N_4507);
nor U10438 (N_10438,N_3231,N_971);
and U10439 (N_10439,N_5181,N_5930);
nor U10440 (N_10440,N_1519,N_5218);
or U10441 (N_10441,N_2302,N_868);
or U10442 (N_10442,N_268,N_424);
xnor U10443 (N_10443,N_215,N_603);
nor U10444 (N_10444,N_3523,N_2073);
xnor U10445 (N_10445,N_113,N_5725);
or U10446 (N_10446,N_175,N_4992);
xor U10447 (N_10447,N_2583,N_3136);
xor U10448 (N_10448,N_3477,N_5151);
or U10449 (N_10449,N_5628,N_4929);
nand U10450 (N_10450,N_3029,N_533);
or U10451 (N_10451,N_5663,N_3240);
xor U10452 (N_10452,N_910,N_4787);
xnor U10453 (N_10453,N_2320,N_4988);
xnor U10454 (N_10454,N_3519,N_3599);
nor U10455 (N_10455,N_323,N_1226);
nand U10456 (N_10456,N_702,N_5940);
or U10457 (N_10457,N_907,N_183);
and U10458 (N_10458,N_4204,N_423);
and U10459 (N_10459,N_191,N_43);
nor U10460 (N_10460,N_486,N_1995);
and U10461 (N_10461,N_1517,N_3409);
or U10462 (N_10462,N_2706,N_1439);
nor U10463 (N_10463,N_3469,N_1292);
and U10464 (N_10464,N_4982,N_773);
nor U10465 (N_10465,N_5936,N_5210);
xnor U10466 (N_10466,N_2894,N_878);
nor U10467 (N_10467,N_255,N_4521);
or U10468 (N_10468,N_1242,N_2237);
or U10469 (N_10469,N_4672,N_3824);
xor U10470 (N_10470,N_5046,N_2819);
or U10471 (N_10471,N_1385,N_5855);
or U10472 (N_10472,N_5606,N_3903);
and U10473 (N_10473,N_5599,N_1049);
nor U10474 (N_10474,N_2828,N_5307);
nor U10475 (N_10475,N_4858,N_2014);
or U10476 (N_10476,N_2079,N_3354);
and U10477 (N_10477,N_1285,N_1799);
nor U10478 (N_10478,N_5158,N_1778);
nand U10479 (N_10479,N_2013,N_3003);
and U10480 (N_10480,N_619,N_3210);
nand U10481 (N_10481,N_1245,N_2925);
nand U10482 (N_10482,N_882,N_446);
nor U10483 (N_10483,N_973,N_753);
nand U10484 (N_10484,N_980,N_1964);
nor U10485 (N_10485,N_3278,N_4367);
xor U10486 (N_10486,N_4357,N_2398);
or U10487 (N_10487,N_584,N_3198);
nor U10488 (N_10488,N_1322,N_3551);
nor U10489 (N_10489,N_636,N_3830);
or U10490 (N_10490,N_5632,N_5271);
and U10491 (N_10491,N_2959,N_483);
nor U10492 (N_10492,N_3913,N_2879);
and U10493 (N_10493,N_1052,N_5829);
or U10494 (N_10494,N_4573,N_4844);
and U10495 (N_10495,N_5102,N_994);
nand U10496 (N_10496,N_2216,N_1148);
xor U10497 (N_10497,N_2998,N_5013);
nand U10498 (N_10498,N_3935,N_48);
xnor U10499 (N_10499,N_1090,N_3666);
nand U10500 (N_10500,N_409,N_3055);
nand U10501 (N_10501,N_3020,N_3610);
xnor U10502 (N_10502,N_2466,N_4158);
nand U10503 (N_10503,N_4586,N_5517);
and U10504 (N_10504,N_1650,N_5796);
and U10505 (N_10505,N_4229,N_1942);
nand U10506 (N_10506,N_2749,N_3141);
xor U10507 (N_10507,N_5038,N_1300);
or U10508 (N_10508,N_5713,N_4352);
and U10509 (N_10509,N_4481,N_1567);
nand U10510 (N_10510,N_5871,N_5311);
and U10511 (N_10511,N_5659,N_3463);
and U10512 (N_10512,N_979,N_1325);
nand U10513 (N_10513,N_5520,N_135);
nor U10514 (N_10514,N_4772,N_118);
nand U10515 (N_10515,N_1420,N_2578);
or U10516 (N_10516,N_5911,N_4177);
or U10517 (N_10517,N_3619,N_3914);
and U10518 (N_10518,N_3761,N_2033);
nor U10519 (N_10519,N_364,N_4574);
nor U10520 (N_10520,N_5534,N_1723);
and U10521 (N_10521,N_5264,N_2110);
nor U10522 (N_10522,N_5099,N_725);
nand U10523 (N_10523,N_4395,N_19);
nor U10524 (N_10524,N_4544,N_1788);
nor U10525 (N_10525,N_5460,N_3774);
nor U10526 (N_10526,N_5910,N_5628);
and U10527 (N_10527,N_5992,N_3606);
nor U10528 (N_10528,N_1738,N_2098);
nand U10529 (N_10529,N_3814,N_4235);
nand U10530 (N_10530,N_5242,N_906);
nor U10531 (N_10531,N_4473,N_5345);
nor U10532 (N_10532,N_3041,N_1882);
nor U10533 (N_10533,N_621,N_1801);
nor U10534 (N_10534,N_1216,N_1845);
nor U10535 (N_10535,N_749,N_3539);
nor U10536 (N_10536,N_4316,N_2368);
xor U10537 (N_10537,N_5281,N_4894);
nand U10538 (N_10538,N_3010,N_273);
or U10539 (N_10539,N_1080,N_869);
nor U10540 (N_10540,N_2799,N_3639);
or U10541 (N_10541,N_3138,N_2822);
nor U10542 (N_10542,N_961,N_2852);
xor U10543 (N_10543,N_4579,N_2613);
or U10544 (N_10544,N_5297,N_1099);
or U10545 (N_10545,N_430,N_193);
xor U10546 (N_10546,N_3818,N_2130);
and U10547 (N_10547,N_1230,N_729);
and U10548 (N_10548,N_4954,N_4958);
and U10549 (N_10549,N_1153,N_3876);
or U10550 (N_10550,N_1340,N_2909);
nor U10551 (N_10551,N_5055,N_3631);
nor U10552 (N_10552,N_2130,N_4983);
nand U10553 (N_10553,N_1900,N_2009);
xnor U10554 (N_10554,N_2686,N_258);
nor U10555 (N_10555,N_1802,N_2620);
xnor U10556 (N_10556,N_1441,N_3392);
nand U10557 (N_10557,N_4089,N_2891);
nor U10558 (N_10558,N_3534,N_3975);
or U10559 (N_10559,N_4071,N_1434);
nand U10560 (N_10560,N_3126,N_1207);
xor U10561 (N_10561,N_3927,N_5132);
nor U10562 (N_10562,N_2109,N_2424);
xnor U10563 (N_10563,N_4824,N_399);
nor U10564 (N_10564,N_137,N_1192);
nor U10565 (N_10565,N_1574,N_402);
or U10566 (N_10566,N_3666,N_5919);
or U10567 (N_10567,N_2355,N_4932);
and U10568 (N_10568,N_5751,N_2167);
nand U10569 (N_10569,N_2306,N_4972);
xnor U10570 (N_10570,N_3585,N_3492);
nor U10571 (N_10571,N_4221,N_1636);
and U10572 (N_10572,N_2554,N_724);
xnor U10573 (N_10573,N_865,N_4975);
or U10574 (N_10574,N_4639,N_3083);
nor U10575 (N_10575,N_891,N_3159);
or U10576 (N_10576,N_2576,N_5336);
or U10577 (N_10577,N_2663,N_310);
and U10578 (N_10578,N_871,N_18);
xor U10579 (N_10579,N_1021,N_4511);
and U10580 (N_10580,N_1737,N_3643);
nor U10581 (N_10581,N_441,N_3024);
nor U10582 (N_10582,N_2172,N_3995);
and U10583 (N_10583,N_3529,N_5468);
or U10584 (N_10584,N_4926,N_4517);
xnor U10585 (N_10585,N_521,N_5073);
nor U10586 (N_10586,N_1827,N_564);
xor U10587 (N_10587,N_5518,N_1965);
nand U10588 (N_10588,N_3004,N_5961);
xor U10589 (N_10589,N_2891,N_834);
or U10590 (N_10590,N_660,N_1372);
nor U10591 (N_10591,N_486,N_2447);
nor U10592 (N_10592,N_361,N_4869);
xnor U10593 (N_10593,N_2834,N_1398);
nand U10594 (N_10594,N_4649,N_5797);
nand U10595 (N_10595,N_4315,N_3938);
nor U10596 (N_10596,N_313,N_1821);
or U10597 (N_10597,N_4322,N_2207);
and U10598 (N_10598,N_4444,N_2798);
nor U10599 (N_10599,N_4957,N_4909);
or U10600 (N_10600,N_3569,N_4583);
or U10601 (N_10601,N_1453,N_656);
or U10602 (N_10602,N_5178,N_5210);
nor U10603 (N_10603,N_4399,N_38);
nor U10604 (N_10604,N_1626,N_237);
nor U10605 (N_10605,N_753,N_5938);
xor U10606 (N_10606,N_4057,N_3144);
nand U10607 (N_10607,N_2771,N_2071);
and U10608 (N_10608,N_1238,N_2140);
nor U10609 (N_10609,N_1529,N_1884);
and U10610 (N_10610,N_1873,N_144);
xnor U10611 (N_10611,N_2279,N_5553);
or U10612 (N_10612,N_3712,N_303);
nor U10613 (N_10613,N_4671,N_4248);
xor U10614 (N_10614,N_2766,N_3192);
xnor U10615 (N_10615,N_2739,N_3097);
and U10616 (N_10616,N_5506,N_4885);
or U10617 (N_10617,N_1224,N_4784);
and U10618 (N_10618,N_5271,N_3223);
nand U10619 (N_10619,N_2790,N_2385);
or U10620 (N_10620,N_1010,N_2157);
nor U10621 (N_10621,N_5572,N_2649);
or U10622 (N_10622,N_1681,N_315);
or U10623 (N_10623,N_5968,N_1677);
nor U10624 (N_10624,N_628,N_564);
and U10625 (N_10625,N_5269,N_743);
nor U10626 (N_10626,N_3751,N_876);
xnor U10627 (N_10627,N_5180,N_5845);
or U10628 (N_10628,N_4942,N_2310);
nand U10629 (N_10629,N_274,N_5924);
and U10630 (N_10630,N_5114,N_2221);
nor U10631 (N_10631,N_5290,N_969);
nor U10632 (N_10632,N_763,N_1241);
and U10633 (N_10633,N_4249,N_1152);
nor U10634 (N_10634,N_5122,N_1289);
and U10635 (N_10635,N_5190,N_3206);
and U10636 (N_10636,N_5225,N_1254);
xnor U10637 (N_10637,N_4176,N_5008);
nor U10638 (N_10638,N_3095,N_1944);
nand U10639 (N_10639,N_5982,N_5049);
and U10640 (N_10640,N_4022,N_218);
or U10641 (N_10641,N_2184,N_3001);
nor U10642 (N_10642,N_2117,N_2292);
nand U10643 (N_10643,N_472,N_2102);
nand U10644 (N_10644,N_4407,N_4960);
xnor U10645 (N_10645,N_1297,N_2390);
and U10646 (N_10646,N_3347,N_4633);
xnor U10647 (N_10647,N_5242,N_3169);
xor U10648 (N_10648,N_3346,N_5967);
nor U10649 (N_10649,N_5438,N_3326);
xor U10650 (N_10650,N_4045,N_1835);
nand U10651 (N_10651,N_3533,N_4857);
xnor U10652 (N_10652,N_1603,N_1767);
xnor U10653 (N_10653,N_3778,N_3884);
nor U10654 (N_10654,N_5966,N_3027);
nor U10655 (N_10655,N_1620,N_1458);
nand U10656 (N_10656,N_2009,N_3256);
nor U10657 (N_10657,N_277,N_5136);
or U10658 (N_10658,N_1504,N_1424);
nand U10659 (N_10659,N_957,N_5053);
xor U10660 (N_10660,N_1470,N_2027);
nor U10661 (N_10661,N_77,N_2098);
xnor U10662 (N_10662,N_1686,N_2980);
xor U10663 (N_10663,N_4842,N_2055);
nand U10664 (N_10664,N_3210,N_3737);
xnor U10665 (N_10665,N_1400,N_4846);
nand U10666 (N_10666,N_209,N_2419);
xor U10667 (N_10667,N_4454,N_5950);
xor U10668 (N_10668,N_5141,N_3850);
nor U10669 (N_10669,N_2044,N_725);
and U10670 (N_10670,N_3589,N_366);
nor U10671 (N_10671,N_4399,N_305);
or U10672 (N_10672,N_271,N_2626);
and U10673 (N_10673,N_2213,N_704);
xnor U10674 (N_10674,N_2801,N_112);
xnor U10675 (N_10675,N_5020,N_542);
nand U10676 (N_10676,N_2945,N_3381);
nor U10677 (N_10677,N_2175,N_1947);
and U10678 (N_10678,N_5207,N_4932);
or U10679 (N_10679,N_2272,N_3844);
nor U10680 (N_10680,N_2547,N_4863);
nand U10681 (N_10681,N_2490,N_3142);
xor U10682 (N_10682,N_5618,N_4004);
nor U10683 (N_10683,N_3988,N_4345);
or U10684 (N_10684,N_5061,N_1911);
and U10685 (N_10685,N_4176,N_1167);
or U10686 (N_10686,N_2856,N_3143);
xor U10687 (N_10687,N_1979,N_2796);
xor U10688 (N_10688,N_1658,N_5201);
nor U10689 (N_10689,N_2687,N_3257);
nor U10690 (N_10690,N_4941,N_641);
xor U10691 (N_10691,N_2592,N_4560);
and U10692 (N_10692,N_5321,N_1817);
and U10693 (N_10693,N_207,N_5998);
xnor U10694 (N_10694,N_4851,N_5468);
nor U10695 (N_10695,N_4918,N_5428);
nor U10696 (N_10696,N_4351,N_2025);
or U10697 (N_10697,N_3782,N_1000);
xor U10698 (N_10698,N_3695,N_1801);
and U10699 (N_10699,N_4405,N_1107);
and U10700 (N_10700,N_147,N_143);
nand U10701 (N_10701,N_243,N_2447);
and U10702 (N_10702,N_371,N_1178);
and U10703 (N_10703,N_2742,N_3814);
nand U10704 (N_10704,N_2311,N_1098);
or U10705 (N_10705,N_4703,N_1517);
or U10706 (N_10706,N_2539,N_4469);
nand U10707 (N_10707,N_5449,N_4601);
or U10708 (N_10708,N_1455,N_3245);
xnor U10709 (N_10709,N_326,N_3047);
nand U10710 (N_10710,N_2689,N_2001);
or U10711 (N_10711,N_5742,N_3193);
or U10712 (N_10712,N_3584,N_3802);
or U10713 (N_10713,N_5726,N_5327);
and U10714 (N_10714,N_3243,N_5882);
and U10715 (N_10715,N_1024,N_2958);
nand U10716 (N_10716,N_1943,N_622);
nand U10717 (N_10717,N_4264,N_2251);
xor U10718 (N_10718,N_4944,N_3835);
or U10719 (N_10719,N_262,N_72);
nor U10720 (N_10720,N_4243,N_2299);
nor U10721 (N_10721,N_1222,N_5953);
nor U10722 (N_10722,N_3674,N_278);
nand U10723 (N_10723,N_3411,N_2297);
nor U10724 (N_10724,N_3525,N_2311);
nor U10725 (N_10725,N_5288,N_5809);
or U10726 (N_10726,N_4634,N_1412);
and U10727 (N_10727,N_5378,N_3193);
nand U10728 (N_10728,N_5613,N_1522);
nor U10729 (N_10729,N_5048,N_2924);
nand U10730 (N_10730,N_1313,N_5461);
and U10731 (N_10731,N_5973,N_5410);
xor U10732 (N_10732,N_2039,N_1238);
nand U10733 (N_10733,N_5228,N_5995);
and U10734 (N_10734,N_2356,N_4691);
nor U10735 (N_10735,N_2225,N_3518);
nor U10736 (N_10736,N_3162,N_1913);
or U10737 (N_10737,N_3890,N_2897);
xnor U10738 (N_10738,N_4265,N_357);
nand U10739 (N_10739,N_1059,N_2918);
xnor U10740 (N_10740,N_1574,N_3088);
nor U10741 (N_10741,N_4941,N_1442);
nor U10742 (N_10742,N_3030,N_2467);
nor U10743 (N_10743,N_2444,N_3353);
xor U10744 (N_10744,N_850,N_2881);
nor U10745 (N_10745,N_5317,N_100);
nand U10746 (N_10746,N_3893,N_4308);
xnor U10747 (N_10747,N_5445,N_4189);
nand U10748 (N_10748,N_1131,N_5407);
nor U10749 (N_10749,N_5811,N_1408);
nor U10750 (N_10750,N_5892,N_432);
nor U10751 (N_10751,N_1241,N_409);
nand U10752 (N_10752,N_5366,N_2963);
and U10753 (N_10753,N_2455,N_5234);
or U10754 (N_10754,N_4625,N_4311);
nor U10755 (N_10755,N_3856,N_1405);
nor U10756 (N_10756,N_3447,N_4771);
xor U10757 (N_10757,N_5398,N_3312);
and U10758 (N_10758,N_3498,N_5551);
and U10759 (N_10759,N_208,N_1083);
nor U10760 (N_10760,N_2244,N_4957);
and U10761 (N_10761,N_4356,N_4110);
or U10762 (N_10762,N_94,N_1008);
nand U10763 (N_10763,N_3589,N_2547);
or U10764 (N_10764,N_3672,N_2569);
nor U10765 (N_10765,N_5105,N_2727);
or U10766 (N_10766,N_5570,N_5770);
xor U10767 (N_10767,N_4006,N_5357);
xor U10768 (N_10768,N_2968,N_1005);
and U10769 (N_10769,N_71,N_1856);
xor U10770 (N_10770,N_5987,N_3023);
nor U10771 (N_10771,N_1646,N_2754);
nand U10772 (N_10772,N_1005,N_4181);
nand U10773 (N_10773,N_1319,N_3872);
and U10774 (N_10774,N_2701,N_3056);
nand U10775 (N_10775,N_3521,N_386);
and U10776 (N_10776,N_5105,N_5345);
nand U10777 (N_10777,N_2351,N_636);
and U10778 (N_10778,N_2958,N_5975);
nand U10779 (N_10779,N_4944,N_2408);
nor U10780 (N_10780,N_4116,N_5571);
nor U10781 (N_10781,N_2228,N_457);
nand U10782 (N_10782,N_2550,N_2606);
nand U10783 (N_10783,N_1330,N_1083);
or U10784 (N_10784,N_495,N_5383);
nand U10785 (N_10785,N_3332,N_453);
xnor U10786 (N_10786,N_3759,N_5260);
nand U10787 (N_10787,N_5467,N_4672);
or U10788 (N_10788,N_3768,N_2370);
or U10789 (N_10789,N_5649,N_1776);
and U10790 (N_10790,N_4451,N_5860);
xor U10791 (N_10791,N_2460,N_2136);
xor U10792 (N_10792,N_3361,N_1933);
nand U10793 (N_10793,N_5441,N_2171);
nor U10794 (N_10794,N_583,N_5585);
nor U10795 (N_10795,N_1000,N_556);
nand U10796 (N_10796,N_4479,N_4494);
nor U10797 (N_10797,N_1472,N_3385);
or U10798 (N_10798,N_2327,N_5433);
nor U10799 (N_10799,N_2627,N_2452);
nor U10800 (N_10800,N_4620,N_685);
and U10801 (N_10801,N_799,N_2276);
nor U10802 (N_10802,N_2442,N_205);
or U10803 (N_10803,N_3452,N_716);
nor U10804 (N_10804,N_3696,N_2444);
and U10805 (N_10805,N_3859,N_118);
nand U10806 (N_10806,N_4779,N_525);
xnor U10807 (N_10807,N_1773,N_4606);
xnor U10808 (N_10808,N_2494,N_4481);
nand U10809 (N_10809,N_1681,N_1919);
nand U10810 (N_10810,N_203,N_4215);
xor U10811 (N_10811,N_1793,N_1028);
nand U10812 (N_10812,N_5137,N_5306);
xnor U10813 (N_10813,N_5090,N_2113);
nand U10814 (N_10814,N_2290,N_2047);
and U10815 (N_10815,N_603,N_3962);
or U10816 (N_10816,N_1159,N_2293);
xor U10817 (N_10817,N_3842,N_3055);
nand U10818 (N_10818,N_1405,N_5907);
nor U10819 (N_10819,N_2955,N_3311);
or U10820 (N_10820,N_2191,N_1778);
nand U10821 (N_10821,N_5150,N_1348);
or U10822 (N_10822,N_5003,N_1391);
or U10823 (N_10823,N_5693,N_2493);
or U10824 (N_10824,N_869,N_415);
or U10825 (N_10825,N_720,N_4861);
nor U10826 (N_10826,N_529,N_496);
and U10827 (N_10827,N_4651,N_3617);
xor U10828 (N_10828,N_2290,N_4914);
and U10829 (N_10829,N_5009,N_2313);
or U10830 (N_10830,N_5045,N_2371);
and U10831 (N_10831,N_3255,N_5060);
nand U10832 (N_10832,N_5213,N_979);
nand U10833 (N_10833,N_187,N_1963);
xnor U10834 (N_10834,N_1511,N_5157);
or U10835 (N_10835,N_4040,N_4849);
nor U10836 (N_10836,N_2001,N_1634);
or U10837 (N_10837,N_2142,N_3691);
or U10838 (N_10838,N_5896,N_3013);
nor U10839 (N_10839,N_5198,N_2235);
nand U10840 (N_10840,N_697,N_3312);
or U10841 (N_10841,N_2596,N_5248);
or U10842 (N_10842,N_2294,N_5052);
xnor U10843 (N_10843,N_5849,N_3130);
nor U10844 (N_10844,N_3913,N_118);
and U10845 (N_10845,N_2749,N_4301);
and U10846 (N_10846,N_763,N_3987);
and U10847 (N_10847,N_2074,N_2450);
or U10848 (N_10848,N_4088,N_228);
xnor U10849 (N_10849,N_5230,N_5206);
or U10850 (N_10850,N_1286,N_2368);
nor U10851 (N_10851,N_354,N_5634);
and U10852 (N_10852,N_3075,N_1225);
nand U10853 (N_10853,N_1618,N_5246);
nor U10854 (N_10854,N_1781,N_3642);
nand U10855 (N_10855,N_1133,N_1326);
and U10856 (N_10856,N_1426,N_452);
or U10857 (N_10857,N_5731,N_1793);
xnor U10858 (N_10858,N_2547,N_5150);
and U10859 (N_10859,N_1819,N_4887);
or U10860 (N_10860,N_512,N_4743);
or U10861 (N_10861,N_1159,N_4468);
xor U10862 (N_10862,N_9,N_4602);
and U10863 (N_10863,N_1670,N_5404);
nand U10864 (N_10864,N_3520,N_3302);
nand U10865 (N_10865,N_4403,N_164);
nand U10866 (N_10866,N_939,N_2331);
and U10867 (N_10867,N_4270,N_4733);
and U10868 (N_10868,N_2715,N_4519);
nand U10869 (N_10869,N_2319,N_1360);
or U10870 (N_10870,N_968,N_3588);
or U10871 (N_10871,N_1088,N_2002);
or U10872 (N_10872,N_2508,N_3408);
or U10873 (N_10873,N_614,N_4020);
or U10874 (N_10874,N_70,N_5176);
and U10875 (N_10875,N_1104,N_1024);
and U10876 (N_10876,N_5432,N_3220);
nor U10877 (N_10877,N_3782,N_774);
and U10878 (N_10878,N_4759,N_2749);
or U10879 (N_10879,N_5631,N_1615);
nand U10880 (N_10880,N_4869,N_4147);
or U10881 (N_10881,N_1159,N_2546);
xor U10882 (N_10882,N_4391,N_430);
nand U10883 (N_10883,N_4001,N_1136);
and U10884 (N_10884,N_994,N_4728);
nand U10885 (N_10885,N_2775,N_2959);
or U10886 (N_10886,N_3833,N_1736);
xor U10887 (N_10887,N_1843,N_4554);
nor U10888 (N_10888,N_2743,N_5192);
or U10889 (N_10889,N_4761,N_3479);
nand U10890 (N_10890,N_2472,N_1284);
nor U10891 (N_10891,N_2709,N_5523);
xor U10892 (N_10892,N_5197,N_2165);
or U10893 (N_10893,N_3900,N_2696);
xnor U10894 (N_10894,N_3739,N_233);
and U10895 (N_10895,N_5366,N_5390);
nand U10896 (N_10896,N_3886,N_4498);
nand U10897 (N_10897,N_666,N_1225);
nand U10898 (N_10898,N_4020,N_4540);
nand U10899 (N_10899,N_3585,N_2217);
nor U10900 (N_10900,N_4010,N_245);
nand U10901 (N_10901,N_543,N_673);
or U10902 (N_10902,N_5942,N_4812);
and U10903 (N_10903,N_5951,N_42);
nand U10904 (N_10904,N_4554,N_4431);
xor U10905 (N_10905,N_294,N_2470);
and U10906 (N_10906,N_3732,N_5542);
nand U10907 (N_10907,N_5498,N_2644);
nor U10908 (N_10908,N_2881,N_2992);
xnor U10909 (N_10909,N_4720,N_4064);
or U10910 (N_10910,N_1039,N_3496);
nor U10911 (N_10911,N_4842,N_3478);
and U10912 (N_10912,N_1831,N_5271);
nor U10913 (N_10913,N_1821,N_3242);
or U10914 (N_10914,N_733,N_76);
nor U10915 (N_10915,N_2361,N_2876);
nor U10916 (N_10916,N_139,N_4299);
nor U10917 (N_10917,N_1136,N_4967);
or U10918 (N_10918,N_3553,N_1147);
nand U10919 (N_10919,N_2597,N_5064);
nand U10920 (N_10920,N_5141,N_2487);
nor U10921 (N_10921,N_5256,N_4696);
nor U10922 (N_10922,N_1565,N_1506);
nor U10923 (N_10923,N_4647,N_2846);
xor U10924 (N_10924,N_2135,N_3589);
or U10925 (N_10925,N_2099,N_5570);
xor U10926 (N_10926,N_3153,N_1959);
nand U10927 (N_10927,N_2215,N_1303);
or U10928 (N_10928,N_3228,N_3588);
nor U10929 (N_10929,N_5583,N_3313);
xnor U10930 (N_10930,N_5808,N_834);
or U10931 (N_10931,N_446,N_3352);
or U10932 (N_10932,N_1430,N_4592);
xor U10933 (N_10933,N_921,N_875);
xnor U10934 (N_10934,N_4834,N_1195);
or U10935 (N_10935,N_4439,N_3598);
nand U10936 (N_10936,N_5417,N_2985);
nor U10937 (N_10937,N_5258,N_1370);
nand U10938 (N_10938,N_4077,N_5522);
or U10939 (N_10939,N_855,N_5215);
and U10940 (N_10940,N_2979,N_3107);
nand U10941 (N_10941,N_2927,N_2860);
or U10942 (N_10942,N_2324,N_2399);
or U10943 (N_10943,N_496,N_4406);
and U10944 (N_10944,N_1746,N_272);
nor U10945 (N_10945,N_901,N_4594);
or U10946 (N_10946,N_5314,N_3181);
xor U10947 (N_10947,N_1629,N_834);
xor U10948 (N_10948,N_3658,N_4908);
nand U10949 (N_10949,N_3343,N_3487);
and U10950 (N_10950,N_1613,N_3573);
or U10951 (N_10951,N_5567,N_5107);
nor U10952 (N_10952,N_3409,N_5468);
xor U10953 (N_10953,N_2274,N_2065);
and U10954 (N_10954,N_156,N_3247);
or U10955 (N_10955,N_2998,N_3955);
xor U10956 (N_10956,N_2374,N_5819);
nor U10957 (N_10957,N_779,N_3474);
nand U10958 (N_10958,N_2603,N_2895);
and U10959 (N_10959,N_2126,N_4654);
xor U10960 (N_10960,N_2066,N_5769);
and U10961 (N_10961,N_4047,N_3077);
nor U10962 (N_10962,N_772,N_3479);
xor U10963 (N_10963,N_5455,N_3947);
nand U10964 (N_10964,N_968,N_2955);
nand U10965 (N_10965,N_3937,N_17);
and U10966 (N_10966,N_5008,N_1475);
or U10967 (N_10967,N_3148,N_4241);
xor U10968 (N_10968,N_1891,N_2156);
nand U10969 (N_10969,N_1664,N_1526);
xnor U10970 (N_10970,N_5388,N_4912);
xnor U10971 (N_10971,N_226,N_3766);
nor U10972 (N_10972,N_561,N_5237);
and U10973 (N_10973,N_4824,N_215);
xnor U10974 (N_10974,N_4304,N_3668);
or U10975 (N_10975,N_314,N_1405);
nand U10976 (N_10976,N_2107,N_2145);
or U10977 (N_10977,N_1194,N_4340);
nor U10978 (N_10978,N_2472,N_923);
nor U10979 (N_10979,N_5957,N_4123);
or U10980 (N_10980,N_1210,N_5162);
or U10981 (N_10981,N_994,N_5166);
and U10982 (N_10982,N_1235,N_1783);
nor U10983 (N_10983,N_4935,N_1523);
xnor U10984 (N_10984,N_197,N_5251);
nor U10985 (N_10985,N_5884,N_1878);
xor U10986 (N_10986,N_1957,N_5303);
nor U10987 (N_10987,N_1198,N_652);
xnor U10988 (N_10988,N_5767,N_2241);
nand U10989 (N_10989,N_951,N_2693);
nand U10990 (N_10990,N_3577,N_3713);
nor U10991 (N_10991,N_4717,N_2281);
and U10992 (N_10992,N_871,N_4498);
or U10993 (N_10993,N_844,N_4946);
and U10994 (N_10994,N_5580,N_4577);
nor U10995 (N_10995,N_3330,N_456);
nand U10996 (N_10996,N_4832,N_1956);
nor U10997 (N_10997,N_5286,N_4305);
xor U10998 (N_10998,N_1157,N_2838);
and U10999 (N_10999,N_748,N_4509);
or U11000 (N_11000,N_1806,N_3865);
or U11001 (N_11001,N_5830,N_4005);
and U11002 (N_11002,N_3632,N_2432);
and U11003 (N_11003,N_3907,N_1925);
or U11004 (N_11004,N_1030,N_2177);
nor U11005 (N_11005,N_4681,N_772);
or U11006 (N_11006,N_5646,N_3389);
and U11007 (N_11007,N_3731,N_1908);
and U11008 (N_11008,N_4293,N_635);
nand U11009 (N_11009,N_4885,N_698);
nor U11010 (N_11010,N_5142,N_1628);
xnor U11011 (N_11011,N_1253,N_3491);
nor U11012 (N_11012,N_1090,N_4731);
xnor U11013 (N_11013,N_5897,N_5031);
and U11014 (N_11014,N_5938,N_5162);
and U11015 (N_11015,N_1465,N_233);
or U11016 (N_11016,N_1351,N_4529);
and U11017 (N_11017,N_1515,N_1535);
nor U11018 (N_11018,N_2619,N_5610);
nand U11019 (N_11019,N_4892,N_1815);
or U11020 (N_11020,N_1077,N_3765);
nand U11021 (N_11021,N_5779,N_3904);
nand U11022 (N_11022,N_5717,N_676);
or U11023 (N_11023,N_5189,N_917);
and U11024 (N_11024,N_3400,N_4091);
xnor U11025 (N_11025,N_928,N_4505);
nand U11026 (N_11026,N_1746,N_2156);
xnor U11027 (N_11027,N_197,N_3775);
or U11028 (N_11028,N_5823,N_4385);
or U11029 (N_11029,N_1740,N_1770);
and U11030 (N_11030,N_5905,N_1365);
nand U11031 (N_11031,N_781,N_782);
xor U11032 (N_11032,N_5999,N_5894);
or U11033 (N_11033,N_5112,N_3844);
nor U11034 (N_11034,N_601,N_4013);
or U11035 (N_11035,N_408,N_2450);
or U11036 (N_11036,N_4002,N_1901);
xnor U11037 (N_11037,N_4714,N_5627);
and U11038 (N_11038,N_5190,N_1380);
or U11039 (N_11039,N_621,N_5740);
xor U11040 (N_11040,N_5552,N_4009);
and U11041 (N_11041,N_4926,N_2629);
xor U11042 (N_11042,N_4273,N_5564);
or U11043 (N_11043,N_936,N_5419);
xor U11044 (N_11044,N_221,N_4742);
nand U11045 (N_11045,N_2734,N_4704);
and U11046 (N_11046,N_3450,N_2804);
nand U11047 (N_11047,N_4955,N_4979);
xor U11048 (N_11048,N_4236,N_1830);
or U11049 (N_11049,N_5191,N_1642);
nor U11050 (N_11050,N_1764,N_271);
nand U11051 (N_11051,N_3757,N_2913);
nor U11052 (N_11052,N_863,N_5028);
nor U11053 (N_11053,N_2521,N_1203);
nand U11054 (N_11054,N_4818,N_2170);
or U11055 (N_11055,N_1229,N_1247);
nor U11056 (N_11056,N_2708,N_4164);
nand U11057 (N_11057,N_1069,N_573);
nor U11058 (N_11058,N_1700,N_4931);
nand U11059 (N_11059,N_1133,N_2118);
or U11060 (N_11060,N_129,N_3730);
or U11061 (N_11061,N_4881,N_5278);
and U11062 (N_11062,N_4995,N_1727);
or U11063 (N_11063,N_1277,N_1871);
xor U11064 (N_11064,N_4025,N_4352);
nor U11065 (N_11065,N_2407,N_1962);
nor U11066 (N_11066,N_586,N_4917);
and U11067 (N_11067,N_1963,N_3234);
and U11068 (N_11068,N_1788,N_5396);
and U11069 (N_11069,N_2802,N_5424);
and U11070 (N_11070,N_378,N_204);
xor U11071 (N_11071,N_1445,N_2649);
nor U11072 (N_11072,N_5747,N_2413);
xor U11073 (N_11073,N_2167,N_1909);
nor U11074 (N_11074,N_122,N_1424);
or U11075 (N_11075,N_3344,N_1831);
or U11076 (N_11076,N_903,N_3447);
and U11077 (N_11077,N_2572,N_3222);
xnor U11078 (N_11078,N_5395,N_1527);
or U11079 (N_11079,N_400,N_1560);
xnor U11080 (N_11080,N_1050,N_766);
nand U11081 (N_11081,N_2986,N_2374);
or U11082 (N_11082,N_5802,N_4592);
and U11083 (N_11083,N_3732,N_5086);
or U11084 (N_11084,N_2879,N_2371);
nor U11085 (N_11085,N_5600,N_195);
nand U11086 (N_11086,N_3908,N_5115);
nor U11087 (N_11087,N_4288,N_2840);
or U11088 (N_11088,N_4382,N_3006);
nand U11089 (N_11089,N_4478,N_4759);
xor U11090 (N_11090,N_4719,N_3776);
and U11091 (N_11091,N_247,N_580);
nor U11092 (N_11092,N_1510,N_2942);
and U11093 (N_11093,N_993,N_1540);
and U11094 (N_11094,N_5666,N_1819);
and U11095 (N_11095,N_5723,N_1474);
nor U11096 (N_11096,N_1555,N_5029);
nor U11097 (N_11097,N_3042,N_5274);
nor U11098 (N_11098,N_2580,N_4772);
nand U11099 (N_11099,N_257,N_2295);
and U11100 (N_11100,N_5802,N_2469);
nor U11101 (N_11101,N_5214,N_2920);
or U11102 (N_11102,N_1193,N_4221);
nor U11103 (N_11103,N_5397,N_3403);
nand U11104 (N_11104,N_5021,N_4776);
xnor U11105 (N_11105,N_5794,N_1342);
nand U11106 (N_11106,N_5090,N_5827);
nor U11107 (N_11107,N_5405,N_1098);
and U11108 (N_11108,N_4094,N_4743);
nor U11109 (N_11109,N_477,N_3914);
and U11110 (N_11110,N_1083,N_1832);
nor U11111 (N_11111,N_5220,N_4579);
xor U11112 (N_11112,N_5978,N_1912);
and U11113 (N_11113,N_4586,N_5718);
and U11114 (N_11114,N_2801,N_4170);
nand U11115 (N_11115,N_2020,N_10);
xnor U11116 (N_11116,N_4631,N_1444);
nor U11117 (N_11117,N_2472,N_5731);
nor U11118 (N_11118,N_5496,N_2093);
xor U11119 (N_11119,N_1116,N_2848);
or U11120 (N_11120,N_3452,N_3634);
or U11121 (N_11121,N_5057,N_525);
nand U11122 (N_11122,N_3944,N_5645);
xnor U11123 (N_11123,N_2915,N_3813);
and U11124 (N_11124,N_5466,N_4654);
nor U11125 (N_11125,N_651,N_3533);
nor U11126 (N_11126,N_3933,N_4152);
nor U11127 (N_11127,N_199,N_2978);
xnor U11128 (N_11128,N_3319,N_1503);
nor U11129 (N_11129,N_4871,N_2571);
or U11130 (N_11130,N_5706,N_1608);
nor U11131 (N_11131,N_4898,N_1037);
and U11132 (N_11132,N_2063,N_5080);
nor U11133 (N_11133,N_3281,N_4644);
and U11134 (N_11134,N_2063,N_2365);
and U11135 (N_11135,N_4512,N_3463);
xor U11136 (N_11136,N_4813,N_2741);
and U11137 (N_11137,N_2580,N_80);
nand U11138 (N_11138,N_618,N_1997);
nor U11139 (N_11139,N_2331,N_5986);
and U11140 (N_11140,N_3154,N_1236);
or U11141 (N_11141,N_501,N_2542);
xor U11142 (N_11142,N_3944,N_5227);
nor U11143 (N_11143,N_3231,N_2176);
nor U11144 (N_11144,N_4774,N_326);
and U11145 (N_11145,N_3227,N_4381);
nand U11146 (N_11146,N_2528,N_14);
or U11147 (N_11147,N_1649,N_5348);
nor U11148 (N_11148,N_951,N_945);
and U11149 (N_11149,N_3731,N_3865);
and U11150 (N_11150,N_1187,N_5081);
nand U11151 (N_11151,N_4409,N_748);
nand U11152 (N_11152,N_2072,N_3519);
nand U11153 (N_11153,N_2768,N_4823);
xor U11154 (N_11154,N_5464,N_3570);
xor U11155 (N_11155,N_4800,N_4140);
nor U11156 (N_11156,N_5380,N_5655);
or U11157 (N_11157,N_2093,N_1);
or U11158 (N_11158,N_145,N_1086);
nor U11159 (N_11159,N_3969,N_2259);
nand U11160 (N_11160,N_4585,N_3414);
nand U11161 (N_11161,N_2421,N_807);
and U11162 (N_11162,N_883,N_3147);
and U11163 (N_11163,N_4053,N_4457);
nand U11164 (N_11164,N_217,N_3110);
nor U11165 (N_11165,N_3803,N_2063);
and U11166 (N_11166,N_3835,N_5221);
nor U11167 (N_11167,N_513,N_751);
nor U11168 (N_11168,N_1484,N_5539);
nand U11169 (N_11169,N_2767,N_3548);
or U11170 (N_11170,N_1979,N_3651);
nor U11171 (N_11171,N_474,N_5425);
nand U11172 (N_11172,N_2231,N_2391);
or U11173 (N_11173,N_888,N_1919);
nor U11174 (N_11174,N_5913,N_3980);
xnor U11175 (N_11175,N_4535,N_4741);
and U11176 (N_11176,N_2382,N_3249);
nor U11177 (N_11177,N_4898,N_129);
nor U11178 (N_11178,N_4779,N_328);
nor U11179 (N_11179,N_159,N_548);
nand U11180 (N_11180,N_433,N_902);
and U11181 (N_11181,N_5480,N_3554);
or U11182 (N_11182,N_1943,N_1042);
nor U11183 (N_11183,N_4445,N_767);
and U11184 (N_11184,N_5301,N_4023);
nand U11185 (N_11185,N_1494,N_1480);
and U11186 (N_11186,N_3952,N_4374);
xor U11187 (N_11187,N_3463,N_55);
nand U11188 (N_11188,N_4554,N_4886);
xnor U11189 (N_11189,N_3806,N_5415);
and U11190 (N_11190,N_2073,N_2219);
or U11191 (N_11191,N_1412,N_4924);
xnor U11192 (N_11192,N_1200,N_1668);
xor U11193 (N_11193,N_4730,N_2737);
or U11194 (N_11194,N_4973,N_1571);
nor U11195 (N_11195,N_3090,N_3975);
nor U11196 (N_11196,N_487,N_2434);
and U11197 (N_11197,N_699,N_1328);
nor U11198 (N_11198,N_2736,N_5628);
nand U11199 (N_11199,N_1413,N_5537);
and U11200 (N_11200,N_4731,N_3262);
nand U11201 (N_11201,N_1074,N_5156);
nand U11202 (N_11202,N_5720,N_2270);
nor U11203 (N_11203,N_5759,N_5829);
and U11204 (N_11204,N_5488,N_2604);
or U11205 (N_11205,N_2739,N_326);
xnor U11206 (N_11206,N_1817,N_1907);
nand U11207 (N_11207,N_5014,N_2304);
or U11208 (N_11208,N_242,N_919);
nor U11209 (N_11209,N_1454,N_602);
nor U11210 (N_11210,N_2296,N_4090);
and U11211 (N_11211,N_3623,N_1497);
nor U11212 (N_11212,N_3840,N_1957);
or U11213 (N_11213,N_1096,N_776);
nor U11214 (N_11214,N_5536,N_3544);
nor U11215 (N_11215,N_134,N_5286);
nand U11216 (N_11216,N_2594,N_2123);
nor U11217 (N_11217,N_2042,N_1891);
nand U11218 (N_11218,N_3839,N_3649);
xnor U11219 (N_11219,N_20,N_3334);
xnor U11220 (N_11220,N_5908,N_4608);
xor U11221 (N_11221,N_2972,N_1118);
xnor U11222 (N_11222,N_3113,N_854);
xnor U11223 (N_11223,N_1861,N_3764);
nand U11224 (N_11224,N_5072,N_3460);
xor U11225 (N_11225,N_835,N_5282);
and U11226 (N_11226,N_5418,N_5528);
and U11227 (N_11227,N_5184,N_681);
and U11228 (N_11228,N_2606,N_3974);
nor U11229 (N_11229,N_4,N_1614);
nor U11230 (N_11230,N_2531,N_269);
and U11231 (N_11231,N_42,N_3093);
and U11232 (N_11232,N_1885,N_3743);
xor U11233 (N_11233,N_3665,N_1000);
nand U11234 (N_11234,N_2696,N_2129);
xnor U11235 (N_11235,N_2650,N_168);
or U11236 (N_11236,N_102,N_2239);
xnor U11237 (N_11237,N_2899,N_3195);
and U11238 (N_11238,N_4598,N_2659);
nand U11239 (N_11239,N_1999,N_391);
nor U11240 (N_11240,N_3314,N_1715);
or U11241 (N_11241,N_3776,N_1600);
nand U11242 (N_11242,N_3380,N_384);
and U11243 (N_11243,N_748,N_1972);
xnor U11244 (N_11244,N_5691,N_802);
and U11245 (N_11245,N_4089,N_2008);
or U11246 (N_11246,N_3852,N_2952);
or U11247 (N_11247,N_2078,N_2955);
nor U11248 (N_11248,N_2227,N_1258);
nand U11249 (N_11249,N_1311,N_5738);
or U11250 (N_11250,N_2690,N_2607);
or U11251 (N_11251,N_703,N_1239);
and U11252 (N_11252,N_1142,N_4848);
nand U11253 (N_11253,N_3990,N_4428);
or U11254 (N_11254,N_338,N_5379);
xor U11255 (N_11255,N_2777,N_857);
and U11256 (N_11256,N_1756,N_2351);
nor U11257 (N_11257,N_3770,N_5972);
or U11258 (N_11258,N_3322,N_5766);
nand U11259 (N_11259,N_5665,N_3575);
xnor U11260 (N_11260,N_9,N_4363);
nand U11261 (N_11261,N_2464,N_3597);
nand U11262 (N_11262,N_582,N_4162);
xor U11263 (N_11263,N_4620,N_5646);
or U11264 (N_11264,N_350,N_4582);
nand U11265 (N_11265,N_2300,N_854);
nor U11266 (N_11266,N_623,N_3149);
and U11267 (N_11267,N_4697,N_3753);
nand U11268 (N_11268,N_1403,N_1808);
and U11269 (N_11269,N_5852,N_5251);
and U11270 (N_11270,N_966,N_882);
nand U11271 (N_11271,N_2668,N_895);
nand U11272 (N_11272,N_5570,N_5745);
nand U11273 (N_11273,N_2204,N_2197);
xnor U11274 (N_11274,N_4153,N_1766);
or U11275 (N_11275,N_5975,N_939);
and U11276 (N_11276,N_5767,N_4995);
and U11277 (N_11277,N_2897,N_4410);
nand U11278 (N_11278,N_5522,N_5294);
and U11279 (N_11279,N_3044,N_1521);
nor U11280 (N_11280,N_5273,N_737);
xnor U11281 (N_11281,N_2724,N_4672);
or U11282 (N_11282,N_3192,N_5084);
nor U11283 (N_11283,N_2593,N_5390);
and U11284 (N_11284,N_2746,N_1597);
or U11285 (N_11285,N_4991,N_952);
and U11286 (N_11286,N_2409,N_2445);
and U11287 (N_11287,N_2366,N_3470);
nand U11288 (N_11288,N_3277,N_790);
or U11289 (N_11289,N_5227,N_972);
xor U11290 (N_11290,N_1778,N_5145);
or U11291 (N_11291,N_2479,N_906);
xor U11292 (N_11292,N_2513,N_2362);
xnor U11293 (N_11293,N_2984,N_1748);
nand U11294 (N_11294,N_48,N_5462);
and U11295 (N_11295,N_1398,N_2727);
or U11296 (N_11296,N_4516,N_981);
nor U11297 (N_11297,N_3589,N_5598);
and U11298 (N_11298,N_3813,N_1404);
or U11299 (N_11299,N_4426,N_2574);
nand U11300 (N_11300,N_4102,N_627);
or U11301 (N_11301,N_394,N_5846);
nor U11302 (N_11302,N_5796,N_3567);
and U11303 (N_11303,N_3473,N_1002);
nand U11304 (N_11304,N_3764,N_5472);
and U11305 (N_11305,N_1959,N_2468);
nor U11306 (N_11306,N_5935,N_1399);
xnor U11307 (N_11307,N_1614,N_1173);
xnor U11308 (N_11308,N_1641,N_1478);
nand U11309 (N_11309,N_1307,N_2930);
nor U11310 (N_11310,N_4171,N_1359);
xor U11311 (N_11311,N_5752,N_4048);
or U11312 (N_11312,N_937,N_2802);
nor U11313 (N_11313,N_1146,N_4435);
nand U11314 (N_11314,N_690,N_3241);
nor U11315 (N_11315,N_5601,N_2317);
nand U11316 (N_11316,N_435,N_1749);
or U11317 (N_11317,N_3285,N_528);
or U11318 (N_11318,N_907,N_280);
xor U11319 (N_11319,N_1073,N_1309);
nand U11320 (N_11320,N_1256,N_3212);
xor U11321 (N_11321,N_5362,N_298);
nand U11322 (N_11322,N_1840,N_4802);
and U11323 (N_11323,N_2624,N_4496);
nand U11324 (N_11324,N_2933,N_5526);
nand U11325 (N_11325,N_613,N_4100);
xor U11326 (N_11326,N_2781,N_5727);
and U11327 (N_11327,N_5966,N_1584);
xnor U11328 (N_11328,N_4988,N_1111);
and U11329 (N_11329,N_4753,N_653);
and U11330 (N_11330,N_1205,N_74);
nor U11331 (N_11331,N_5012,N_4867);
nand U11332 (N_11332,N_87,N_2027);
nand U11333 (N_11333,N_1712,N_4256);
or U11334 (N_11334,N_5430,N_785);
nor U11335 (N_11335,N_2845,N_4285);
nor U11336 (N_11336,N_327,N_3058);
and U11337 (N_11337,N_384,N_2329);
and U11338 (N_11338,N_4676,N_2858);
nand U11339 (N_11339,N_3518,N_4266);
nand U11340 (N_11340,N_461,N_2775);
and U11341 (N_11341,N_4606,N_2599);
or U11342 (N_11342,N_4305,N_5384);
nor U11343 (N_11343,N_2120,N_3056);
nand U11344 (N_11344,N_245,N_4698);
xnor U11345 (N_11345,N_3175,N_1646);
nand U11346 (N_11346,N_3916,N_2657);
nand U11347 (N_11347,N_3660,N_5324);
and U11348 (N_11348,N_5050,N_2481);
nand U11349 (N_11349,N_4219,N_3248);
xor U11350 (N_11350,N_3179,N_3951);
nand U11351 (N_11351,N_3985,N_1580);
and U11352 (N_11352,N_5940,N_1451);
nand U11353 (N_11353,N_1072,N_96);
and U11354 (N_11354,N_3403,N_2561);
and U11355 (N_11355,N_4860,N_5968);
xnor U11356 (N_11356,N_5457,N_317);
nor U11357 (N_11357,N_1948,N_2724);
and U11358 (N_11358,N_124,N_4310);
and U11359 (N_11359,N_1816,N_683);
xnor U11360 (N_11360,N_1913,N_2257);
xnor U11361 (N_11361,N_4722,N_1569);
or U11362 (N_11362,N_3116,N_3193);
or U11363 (N_11363,N_1175,N_2142);
and U11364 (N_11364,N_3941,N_5984);
nor U11365 (N_11365,N_3683,N_3718);
xnor U11366 (N_11366,N_5199,N_3740);
and U11367 (N_11367,N_4482,N_4901);
nor U11368 (N_11368,N_4371,N_4452);
nand U11369 (N_11369,N_217,N_3624);
nand U11370 (N_11370,N_5497,N_4126);
or U11371 (N_11371,N_831,N_851);
nand U11372 (N_11372,N_2843,N_2703);
xnor U11373 (N_11373,N_2207,N_2445);
nand U11374 (N_11374,N_1968,N_4591);
nand U11375 (N_11375,N_2301,N_5511);
nand U11376 (N_11376,N_2766,N_2227);
nand U11377 (N_11377,N_1931,N_1787);
nor U11378 (N_11378,N_309,N_893);
and U11379 (N_11379,N_2308,N_2949);
xor U11380 (N_11380,N_5324,N_1596);
xor U11381 (N_11381,N_5473,N_4686);
xnor U11382 (N_11382,N_1082,N_1657);
or U11383 (N_11383,N_2110,N_442);
nand U11384 (N_11384,N_311,N_1529);
or U11385 (N_11385,N_464,N_1374);
and U11386 (N_11386,N_4096,N_2386);
nor U11387 (N_11387,N_4971,N_4467);
xnor U11388 (N_11388,N_2504,N_3087);
nand U11389 (N_11389,N_2643,N_3597);
nand U11390 (N_11390,N_5972,N_3584);
nor U11391 (N_11391,N_3618,N_2871);
nor U11392 (N_11392,N_2331,N_172);
xnor U11393 (N_11393,N_3787,N_2373);
or U11394 (N_11394,N_2439,N_5499);
and U11395 (N_11395,N_4680,N_2151);
or U11396 (N_11396,N_4384,N_2858);
xor U11397 (N_11397,N_865,N_2067);
xor U11398 (N_11398,N_3935,N_4315);
nor U11399 (N_11399,N_4690,N_563);
and U11400 (N_11400,N_594,N_2042);
nor U11401 (N_11401,N_624,N_2512);
or U11402 (N_11402,N_1650,N_2036);
xor U11403 (N_11403,N_2948,N_2681);
xnor U11404 (N_11404,N_2553,N_3127);
nand U11405 (N_11405,N_445,N_4171);
nor U11406 (N_11406,N_3939,N_5645);
xor U11407 (N_11407,N_1962,N_1755);
nor U11408 (N_11408,N_4095,N_882);
nor U11409 (N_11409,N_1430,N_1198);
nand U11410 (N_11410,N_3897,N_3160);
or U11411 (N_11411,N_1784,N_5106);
or U11412 (N_11412,N_2219,N_5877);
nor U11413 (N_11413,N_733,N_1094);
or U11414 (N_11414,N_1899,N_4873);
xnor U11415 (N_11415,N_3208,N_2065);
nand U11416 (N_11416,N_2796,N_2992);
nand U11417 (N_11417,N_204,N_4883);
nor U11418 (N_11418,N_5674,N_1643);
xnor U11419 (N_11419,N_1230,N_386);
or U11420 (N_11420,N_2954,N_5606);
or U11421 (N_11421,N_2353,N_5049);
nor U11422 (N_11422,N_1401,N_1304);
and U11423 (N_11423,N_1894,N_2696);
nand U11424 (N_11424,N_5199,N_3822);
nor U11425 (N_11425,N_2688,N_956);
and U11426 (N_11426,N_1,N_3018);
xnor U11427 (N_11427,N_917,N_221);
xor U11428 (N_11428,N_5568,N_4689);
and U11429 (N_11429,N_4401,N_1577);
xnor U11430 (N_11430,N_5561,N_4863);
nor U11431 (N_11431,N_66,N_3563);
or U11432 (N_11432,N_2757,N_3261);
nand U11433 (N_11433,N_5699,N_5856);
nand U11434 (N_11434,N_3955,N_1704);
nand U11435 (N_11435,N_3203,N_3061);
and U11436 (N_11436,N_1962,N_1520);
or U11437 (N_11437,N_4670,N_5861);
nor U11438 (N_11438,N_5460,N_57);
nor U11439 (N_11439,N_647,N_1018);
nor U11440 (N_11440,N_1949,N_5321);
and U11441 (N_11441,N_155,N_1152);
and U11442 (N_11442,N_2535,N_1393);
or U11443 (N_11443,N_3909,N_5694);
nand U11444 (N_11444,N_2484,N_4665);
or U11445 (N_11445,N_4797,N_3922);
xnor U11446 (N_11446,N_1372,N_5250);
nor U11447 (N_11447,N_281,N_1853);
nor U11448 (N_11448,N_2336,N_64);
or U11449 (N_11449,N_4064,N_4349);
xnor U11450 (N_11450,N_2800,N_4876);
xnor U11451 (N_11451,N_2275,N_5487);
and U11452 (N_11452,N_2125,N_533);
and U11453 (N_11453,N_1842,N_4798);
nor U11454 (N_11454,N_5638,N_1707);
nor U11455 (N_11455,N_2017,N_1860);
nand U11456 (N_11456,N_2135,N_5434);
xnor U11457 (N_11457,N_2174,N_5791);
nor U11458 (N_11458,N_1048,N_3617);
nor U11459 (N_11459,N_3605,N_5191);
nor U11460 (N_11460,N_2199,N_5693);
and U11461 (N_11461,N_1363,N_1436);
xnor U11462 (N_11462,N_1867,N_5581);
xor U11463 (N_11463,N_888,N_2205);
nand U11464 (N_11464,N_1621,N_4217);
nand U11465 (N_11465,N_5236,N_1183);
and U11466 (N_11466,N_2215,N_464);
or U11467 (N_11467,N_2538,N_5012);
or U11468 (N_11468,N_3222,N_5453);
xor U11469 (N_11469,N_1560,N_815);
xor U11470 (N_11470,N_2411,N_3078);
nand U11471 (N_11471,N_295,N_2282);
and U11472 (N_11472,N_1905,N_5131);
xnor U11473 (N_11473,N_5011,N_5066);
nor U11474 (N_11474,N_4303,N_1388);
xnor U11475 (N_11475,N_5251,N_1333);
or U11476 (N_11476,N_3159,N_5044);
xnor U11477 (N_11477,N_3624,N_2752);
nand U11478 (N_11478,N_4414,N_1891);
nand U11479 (N_11479,N_5855,N_1746);
nand U11480 (N_11480,N_5094,N_5302);
nand U11481 (N_11481,N_3057,N_964);
xor U11482 (N_11482,N_4830,N_4731);
xor U11483 (N_11483,N_405,N_2757);
nor U11484 (N_11484,N_1274,N_1189);
and U11485 (N_11485,N_2181,N_3603);
or U11486 (N_11486,N_2949,N_1387);
xnor U11487 (N_11487,N_93,N_1970);
nand U11488 (N_11488,N_5761,N_5891);
nor U11489 (N_11489,N_4191,N_4836);
or U11490 (N_11490,N_1459,N_4612);
nor U11491 (N_11491,N_460,N_1331);
xor U11492 (N_11492,N_5244,N_4555);
nor U11493 (N_11493,N_96,N_2508);
xnor U11494 (N_11494,N_3095,N_4240);
and U11495 (N_11495,N_4406,N_1530);
nand U11496 (N_11496,N_56,N_1016);
nor U11497 (N_11497,N_5982,N_4526);
xnor U11498 (N_11498,N_5757,N_5475);
and U11499 (N_11499,N_4797,N_3310);
and U11500 (N_11500,N_993,N_5318);
xor U11501 (N_11501,N_5997,N_655);
nand U11502 (N_11502,N_1852,N_1380);
nand U11503 (N_11503,N_47,N_4036);
nand U11504 (N_11504,N_421,N_1090);
and U11505 (N_11505,N_2105,N_883);
nor U11506 (N_11506,N_837,N_5437);
nand U11507 (N_11507,N_752,N_3909);
xnor U11508 (N_11508,N_2973,N_1852);
and U11509 (N_11509,N_792,N_4982);
nor U11510 (N_11510,N_2033,N_3735);
or U11511 (N_11511,N_1468,N_5308);
or U11512 (N_11512,N_4513,N_3444);
or U11513 (N_11513,N_5276,N_1799);
or U11514 (N_11514,N_4277,N_449);
and U11515 (N_11515,N_5092,N_5235);
or U11516 (N_11516,N_983,N_1839);
nand U11517 (N_11517,N_2237,N_3614);
and U11518 (N_11518,N_4839,N_2460);
nor U11519 (N_11519,N_2292,N_386);
or U11520 (N_11520,N_1003,N_5554);
nand U11521 (N_11521,N_3497,N_4746);
or U11522 (N_11522,N_1799,N_4072);
xnor U11523 (N_11523,N_5401,N_2396);
nor U11524 (N_11524,N_5169,N_2679);
and U11525 (N_11525,N_5,N_499);
and U11526 (N_11526,N_946,N_2788);
and U11527 (N_11527,N_1974,N_5325);
or U11528 (N_11528,N_3726,N_4726);
and U11529 (N_11529,N_4587,N_2351);
xor U11530 (N_11530,N_2394,N_945);
or U11531 (N_11531,N_4505,N_21);
and U11532 (N_11532,N_2140,N_1411);
nand U11533 (N_11533,N_286,N_242);
xnor U11534 (N_11534,N_1176,N_4271);
nand U11535 (N_11535,N_1637,N_3464);
or U11536 (N_11536,N_1865,N_3165);
and U11537 (N_11537,N_3320,N_5441);
and U11538 (N_11538,N_3838,N_477);
and U11539 (N_11539,N_120,N_1852);
nor U11540 (N_11540,N_1852,N_1478);
nand U11541 (N_11541,N_1819,N_5378);
and U11542 (N_11542,N_2382,N_5526);
nand U11543 (N_11543,N_353,N_866);
xnor U11544 (N_11544,N_4499,N_4548);
or U11545 (N_11545,N_3791,N_2865);
or U11546 (N_11546,N_5677,N_2827);
nor U11547 (N_11547,N_1888,N_4700);
or U11548 (N_11548,N_2940,N_1649);
nand U11549 (N_11549,N_4033,N_2069);
and U11550 (N_11550,N_4040,N_4506);
nor U11551 (N_11551,N_998,N_3071);
nand U11552 (N_11552,N_3709,N_3617);
and U11553 (N_11553,N_1695,N_2109);
nor U11554 (N_11554,N_4092,N_925);
xnor U11555 (N_11555,N_2472,N_5547);
or U11556 (N_11556,N_1838,N_5779);
or U11557 (N_11557,N_1596,N_4502);
nand U11558 (N_11558,N_4892,N_4033);
nand U11559 (N_11559,N_1074,N_1152);
nand U11560 (N_11560,N_190,N_2696);
xor U11561 (N_11561,N_5069,N_5908);
nand U11562 (N_11562,N_291,N_4781);
or U11563 (N_11563,N_5437,N_1088);
or U11564 (N_11564,N_3635,N_434);
or U11565 (N_11565,N_1016,N_5374);
xnor U11566 (N_11566,N_5660,N_2906);
and U11567 (N_11567,N_1964,N_4963);
nor U11568 (N_11568,N_3267,N_3634);
or U11569 (N_11569,N_3699,N_5604);
and U11570 (N_11570,N_3884,N_70);
nor U11571 (N_11571,N_5461,N_2231);
nand U11572 (N_11572,N_5645,N_4319);
or U11573 (N_11573,N_2634,N_5454);
or U11574 (N_11574,N_2470,N_4295);
nor U11575 (N_11575,N_4260,N_494);
nand U11576 (N_11576,N_3423,N_4444);
xor U11577 (N_11577,N_4139,N_0);
nor U11578 (N_11578,N_4621,N_5597);
and U11579 (N_11579,N_2846,N_4600);
and U11580 (N_11580,N_1803,N_2191);
or U11581 (N_11581,N_3678,N_2369);
nand U11582 (N_11582,N_3903,N_3327);
or U11583 (N_11583,N_703,N_4190);
nor U11584 (N_11584,N_2878,N_4146);
or U11585 (N_11585,N_3390,N_1894);
nor U11586 (N_11586,N_2498,N_3484);
and U11587 (N_11587,N_502,N_2098);
or U11588 (N_11588,N_4197,N_5148);
and U11589 (N_11589,N_954,N_2514);
nor U11590 (N_11590,N_530,N_2532);
nand U11591 (N_11591,N_2863,N_5939);
xnor U11592 (N_11592,N_3967,N_2269);
and U11593 (N_11593,N_2662,N_3328);
nand U11594 (N_11594,N_1213,N_923);
and U11595 (N_11595,N_350,N_5090);
nand U11596 (N_11596,N_5431,N_2586);
nor U11597 (N_11597,N_4965,N_4168);
nand U11598 (N_11598,N_3677,N_4754);
or U11599 (N_11599,N_1133,N_1369);
xnor U11600 (N_11600,N_2556,N_5966);
and U11601 (N_11601,N_3315,N_4943);
xor U11602 (N_11602,N_4393,N_5719);
nor U11603 (N_11603,N_2005,N_1772);
or U11604 (N_11604,N_311,N_5366);
nand U11605 (N_11605,N_3687,N_4866);
xor U11606 (N_11606,N_5473,N_1687);
nand U11607 (N_11607,N_3006,N_4084);
xnor U11608 (N_11608,N_3272,N_2766);
xnor U11609 (N_11609,N_331,N_2282);
xnor U11610 (N_11610,N_4832,N_5821);
xor U11611 (N_11611,N_2313,N_5857);
nand U11612 (N_11612,N_5665,N_5263);
and U11613 (N_11613,N_3891,N_4784);
xor U11614 (N_11614,N_3321,N_4318);
nor U11615 (N_11615,N_4061,N_5958);
nand U11616 (N_11616,N_826,N_5597);
or U11617 (N_11617,N_2558,N_1115);
or U11618 (N_11618,N_4530,N_1227);
nand U11619 (N_11619,N_1019,N_2401);
nand U11620 (N_11620,N_3881,N_612);
nand U11621 (N_11621,N_3294,N_3529);
nor U11622 (N_11622,N_1307,N_3377);
xnor U11623 (N_11623,N_1907,N_2731);
nand U11624 (N_11624,N_1577,N_1089);
nand U11625 (N_11625,N_1223,N_1652);
xor U11626 (N_11626,N_4825,N_3862);
nand U11627 (N_11627,N_1295,N_5791);
or U11628 (N_11628,N_5643,N_1070);
or U11629 (N_11629,N_3264,N_3215);
or U11630 (N_11630,N_1196,N_2906);
nand U11631 (N_11631,N_3973,N_3775);
xnor U11632 (N_11632,N_3836,N_5724);
or U11633 (N_11633,N_3545,N_2217);
nor U11634 (N_11634,N_818,N_23);
nand U11635 (N_11635,N_144,N_4715);
and U11636 (N_11636,N_4332,N_5374);
and U11637 (N_11637,N_4185,N_49);
and U11638 (N_11638,N_4187,N_5821);
nor U11639 (N_11639,N_5678,N_5413);
and U11640 (N_11640,N_874,N_5590);
nor U11641 (N_11641,N_4724,N_3022);
nand U11642 (N_11642,N_183,N_652);
and U11643 (N_11643,N_3032,N_2608);
and U11644 (N_11644,N_769,N_3339);
and U11645 (N_11645,N_3603,N_616);
nand U11646 (N_11646,N_5630,N_5758);
nand U11647 (N_11647,N_1611,N_4408);
nand U11648 (N_11648,N_2534,N_5823);
nor U11649 (N_11649,N_1144,N_5647);
nand U11650 (N_11650,N_5222,N_1801);
nand U11651 (N_11651,N_5057,N_3585);
nor U11652 (N_11652,N_5309,N_4788);
nand U11653 (N_11653,N_3284,N_698);
or U11654 (N_11654,N_4767,N_5123);
xnor U11655 (N_11655,N_2865,N_1902);
nor U11656 (N_11656,N_4297,N_3343);
and U11657 (N_11657,N_2772,N_2775);
nor U11658 (N_11658,N_4375,N_613);
or U11659 (N_11659,N_3476,N_2983);
xor U11660 (N_11660,N_3043,N_431);
and U11661 (N_11661,N_5287,N_4806);
nor U11662 (N_11662,N_1412,N_3557);
nor U11663 (N_11663,N_5575,N_4205);
nand U11664 (N_11664,N_5919,N_456);
xnor U11665 (N_11665,N_755,N_4887);
nor U11666 (N_11666,N_813,N_1267);
nor U11667 (N_11667,N_171,N_94);
nand U11668 (N_11668,N_5478,N_63);
xor U11669 (N_11669,N_5952,N_839);
nor U11670 (N_11670,N_5847,N_582);
nand U11671 (N_11671,N_4271,N_135);
or U11672 (N_11672,N_2377,N_869);
and U11673 (N_11673,N_3468,N_5093);
nor U11674 (N_11674,N_1859,N_1975);
nor U11675 (N_11675,N_4419,N_4575);
nand U11676 (N_11676,N_1146,N_3319);
or U11677 (N_11677,N_4679,N_1115);
and U11678 (N_11678,N_5317,N_4779);
nor U11679 (N_11679,N_2264,N_4468);
or U11680 (N_11680,N_4993,N_402);
xor U11681 (N_11681,N_3223,N_4717);
xor U11682 (N_11682,N_956,N_170);
xnor U11683 (N_11683,N_208,N_4262);
nand U11684 (N_11684,N_5165,N_4539);
or U11685 (N_11685,N_2377,N_1141);
and U11686 (N_11686,N_3403,N_5763);
nand U11687 (N_11687,N_2793,N_5193);
nand U11688 (N_11688,N_2865,N_2720);
xnor U11689 (N_11689,N_27,N_1195);
nand U11690 (N_11690,N_5830,N_974);
and U11691 (N_11691,N_5173,N_1372);
xor U11692 (N_11692,N_2129,N_3054);
xor U11693 (N_11693,N_3489,N_3272);
nand U11694 (N_11694,N_4660,N_18);
nand U11695 (N_11695,N_5781,N_657);
xnor U11696 (N_11696,N_5762,N_3258);
nand U11697 (N_11697,N_2556,N_4617);
nor U11698 (N_11698,N_4367,N_1004);
or U11699 (N_11699,N_2505,N_3122);
nor U11700 (N_11700,N_4159,N_5804);
and U11701 (N_11701,N_5339,N_1304);
or U11702 (N_11702,N_3384,N_4661);
nor U11703 (N_11703,N_712,N_2593);
and U11704 (N_11704,N_2007,N_1265);
and U11705 (N_11705,N_951,N_4656);
and U11706 (N_11706,N_561,N_3630);
nand U11707 (N_11707,N_3601,N_2059);
and U11708 (N_11708,N_2032,N_1859);
and U11709 (N_11709,N_2651,N_2599);
nand U11710 (N_11710,N_3282,N_2980);
and U11711 (N_11711,N_3342,N_4194);
xnor U11712 (N_11712,N_2050,N_1666);
nand U11713 (N_11713,N_1331,N_5765);
xor U11714 (N_11714,N_3913,N_3299);
nor U11715 (N_11715,N_4850,N_5304);
and U11716 (N_11716,N_1923,N_1544);
xnor U11717 (N_11717,N_3693,N_2152);
nor U11718 (N_11718,N_1851,N_1596);
nor U11719 (N_11719,N_4964,N_3905);
xor U11720 (N_11720,N_5463,N_5752);
or U11721 (N_11721,N_4550,N_2021);
and U11722 (N_11722,N_3790,N_5794);
nor U11723 (N_11723,N_4825,N_3789);
nor U11724 (N_11724,N_2580,N_4537);
xnor U11725 (N_11725,N_4932,N_1359);
or U11726 (N_11726,N_2334,N_3583);
or U11727 (N_11727,N_4083,N_234);
or U11728 (N_11728,N_5969,N_724);
or U11729 (N_11729,N_582,N_4095);
nand U11730 (N_11730,N_3062,N_33);
or U11731 (N_11731,N_1252,N_4209);
and U11732 (N_11732,N_3058,N_757);
xnor U11733 (N_11733,N_4729,N_3890);
xor U11734 (N_11734,N_407,N_4027);
nand U11735 (N_11735,N_4825,N_2590);
nand U11736 (N_11736,N_5724,N_3961);
nor U11737 (N_11737,N_3505,N_5826);
nor U11738 (N_11738,N_2471,N_3649);
or U11739 (N_11739,N_2477,N_3569);
xnor U11740 (N_11740,N_4333,N_897);
xnor U11741 (N_11741,N_4108,N_5894);
nand U11742 (N_11742,N_1442,N_3485);
nor U11743 (N_11743,N_3982,N_2771);
xor U11744 (N_11744,N_3708,N_3355);
nand U11745 (N_11745,N_4625,N_1149);
or U11746 (N_11746,N_280,N_5001);
and U11747 (N_11747,N_3661,N_2117);
nor U11748 (N_11748,N_967,N_2362);
xnor U11749 (N_11749,N_544,N_2280);
and U11750 (N_11750,N_4348,N_2782);
nand U11751 (N_11751,N_1327,N_3029);
nand U11752 (N_11752,N_2463,N_2921);
xor U11753 (N_11753,N_2601,N_2551);
xor U11754 (N_11754,N_3531,N_3720);
nand U11755 (N_11755,N_1508,N_3672);
nor U11756 (N_11756,N_5449,N_3219);
nand U11757 (N_11757,N_1995,N_258);
xnor U11758 (N_11758,N_2478,N_2451);
nor U11759 (N_11759,N_3287,N_2789);
xnor U11760 (N_11760,N_2216,N_1914);
nand U11761 (N_11761,N_4187,N_1231);
nor U11762 (N_11762,N_2224,N_3367);
nand U11763 (N_11763,N_4470,N_393);
and U11764 (N_11764,N_3559,N_2895);
nand U11765 (N_11765,N_3051,N_1417);
xnor U11766 (N_11766,N_826,N_2889);
nand U11767 (N_11767,N_3953,N_1602);
xnor U11768 (N_11768,N_1869,N_2239);
and U11769 (N_11769,N_3463,N_3319);
nand U11770 (N_11770,N_2935,N_5982);
nor U11771 (N_11771,N_4681,N_1444);
nand U11772 (N_11772,N_2693,N_4804);
nand U11773 (N_11773,N_3897,N_2786);
xnor U11774 (N_11774,N_3000,N_3685);
xor U11775 (N_11775,N_4977,N_3874);
nor U11776 (N_11776,N_3700,N_3040);
nor U11777 (N_11777,N_2396,N_3972);
nor U11778 (N_11778,N_2251,N_3487);
xor U11779 (N_11779,N_166,N_1138);
nor U11780 (N_11780,N_4359,N_5552);
xor U11781 (N_11781,N_5763,N_3047);
and U11782 (N_11782,N_2864,N_5273);
or U11783 (N_11783,N_4855,N_4255);
and U11784 (N_11784,N_809,N_2382);
or U11785 (N_11785,N_3232,N_2957);
nand U11786 (N_11786,N_2443,N_222);
or U11787 (N_11787,N_1526,N_2535);
or U11788 (N_11788,N_4477,N_2593);
nand U11789 (N_11789,N_2550,N_3397);
xnor U11790 (N_11790,N_2029,N_3419);
nand U11791 (N_11791,N_345,N_782);
and U11792 (N_11792,N_2057,N_5484);
and U11793 (N_11793,N_4164,N_4500);
or U11794 (N_11794,N_465,N_4574);
and U11795 (N_11795,N_2609,N_1784);
xnor U11796 (N_11796,N_5560,N_4685);
nand U11797 (N_11797,N_4131,N_5551);
nand U11798 (N_11798,N_3947,N_2518);
nor U11799 (N_11799,N_2615,N_4845);
and U11800 (N_11800,N_5178,N_2109);
xor U11801 (N_11801,N_3065,N_1706);
nor U11802 (N_11802,N_2635,N_4112);
xnor U11803 (N_11803,N_2498,N_1322);
and U11804 (N_11804,N_3144,N_2577);
nand U11805 (N_11805,N_2350,N_2711);
or U11806 (N_11806,N_792,N_1582);
or U11807 (N_11807,N_5527,N_3554);
and U11808 (N_11808,N_3338,N_4356);
nand U11809 (N_11809,N_2989,N_4674);
and U11810 (N_11810,N_2599,N_5634);
nor U11811 (N_11811,N_1064,N_5340);
and U11812 (N_11812,N_418,N_1374);
nor U11813 (N_11813,N_1556,N_1806);
xor U11814 (N_11814,N_4322,N_1190);
or U11815 (N_11815,N_5967,N_2592);
or U11816 (N_11816,N_1118,N_2190);
nand U11817 (N_11817,N_3388,N_5502);
nor U11818 (N_11818,N_5436,N_3674);
xor U11819 (N_11819,N_247,N_265);
xnor U11820 (N_11820,N_2598,N_653);
nor U11821 (N_11821,N_769,N_2213);
xnor U11822 (N_11822,N_2440,N_4551);
or U11823 (N_11823,N_4041,N_4862);
and U11824 (N_11824,N_4020,N_5404);
nor U11825 (N_11825,N_2050,N_2322);
nand U11826 (N_11826,N_3418,N_3792);
nand U11827 (N_11827,N_2305,N_2458);
and U11828 (N_11828,N_3229,N_280);
or U11829 (N_11829,N_3690,N_2338);
and U11830 (N_11830,N_1227,N_4950);
xor U11831 (N_11831,N_5219,N_5674);
or U11832 (N_11832,N_1499,N_2920);
and U11833 (N_11833,N_5144,N_5384);
and U11834 (N_11834,N_1132,N_2182);
and U11835 (N_11835,N_2539,N_5930);
and U11836 (N_11836,N_830,N_1728);
nand U11837 (N_11837,N_4148,N_815);
nor U11838 (N_11838,N_2984,N_2269);
nand U11839 (N_11839,N_1260,N_5395);
or U11840 (N_11840,N_2841,N_5656);
xnor U11841 (N_11841,N_774,N_4780);
nor U11842 (N_11842,N_4214,N_1411);
or U11843 (N_11843,N_4313,N_3726);
nor U11844 (N_11844,N_311,N_3902);
and U11845 (N_11845,N_4922,N_2177);
xnor U11846 (N_11846,N_1528,N_83);
xnor U11847 (N_11847,N_1811,N_4856);
nor U11848 (N_11848,N_2050,N_4246);
or U11849 (N_11849,N_3093,N_3249);
nor U11850 (N_11850,N_3468,N_701);
xnor U11851 (N_11851,N_2194,N_704);
nand U11852 (N_11852,N_1831,N_2272);
nor U11853 (N_11853,N_699,N_5098);
nor U11854 (N_11854,N_2671,N_3496);
and U11855 (N_11855,N_4633,N_3288);
and U11856 (N_11856,N_2844,N_3129);
xnor U11857 (N_11857,N_5449,N_4382);
nor U11858 (N_11858,N_4052,N_3303);
xnor U11859 (N_11859,N_4676,N_1034);
nand U11860 (N_11860,N_4403,N_351);
and U11861 (N_11861,N_4001,N_948);
xnor U11862 (N_11862,N_1869,N_5296);
or U11863 (N_11863,N_2492,N_5630);
and U11864 (N_11864,N_2025,N_1181);
nand U11865 (N_11865,N_5248,N_1558);
and U11866 (N_11866,N_1484,N_3169);
xor U11867 (N_11867,N_1327,N_675);
and U11868 (N_11868,N_3719,N_370);
nand U11869 (N_11869,N_4757,N_5270);
or U11870 (N_11870,N_2394,N_4698);
xnor U11871 (N_11871,N_1341,N_5714);
and U11872 (N_11872,N_3662,N_4302);
or U11873 (N_11873,N_5091,N_3543);
and U11874 (N_11874,N_3283,N_1350);
nor U11875 (N_11875,N_844,N_3181);
and U11876 (N_11876,N_3161,N_4768);
nor U11877 (N_11877,N_5339,N_2050);
and U11878 (N_11878,N_5797,N_753);
and U11879 (N_11879,N_4265,N_1266);
nand U11880 (N_11880,N_1085,N_2414);
and U11881 (N_11881,N_5620,N_782);
xor U11882 (N_11882,N_1621,N_3591);
and U11883 (N_11883,N_399,N_1384);
or U11884 (N_11884,N_751,N_3233);
or U11885 (N_11885,N_3803,N_5211);
xnor U11886 (N_11886,N_1492,N_4416);
and U11887 (N_11887,N_2700,N_4725);
and U11888 (N_11888,N_1159,N_5318);
and U11889 (N_11889,N_5704,N_2911);
xor U11890 (N_11890,N_5034,N_3924);
nand U11891 (N_11891,N_2386,N_2127);
and U11892 (N_11892,N_269,N_1797);
nand U11893 (N_11893,N_3334,N_1815);
and U11894 (N_11894,N_3788,N_848);
and U11895 (N_11895,N_4625,N_1257);
nor U11896 (N_11896,N_5402,N_3956);
nor U11897 (N_11897,N_4129,N_5714);
nand U11898 (N_11898,N_2349,N_1079);
nor U11899 (N_11899,N_3807,N_5747);
nand U11900 (N_11900,N_2278,N_5961);
nand U11901 (N_11901,N_1468,N_2867);
or U11902 (N_11902,N_3319,N_4644);
xor U11903 (N_11903,N_5855,N_3849);
and U11904 (N_11904,N_1653,N_3036);
nor U11905 (N_11905,N_1493,N_5126);
and U11906 (N_11906,N_5561,N_1117);
xor U11907 (N_11907,N_3241,N_2822);
xnor U11908 (N_11908,N_1385,N_2917);
and U11909 (N_11909,N_3512,N_2698);
or U11910 (N_11910,N_313,N_1489);
xor U11911 (N_11911,N_2030,N_1958);
or U11912 (N_11912,N_236,N_2534);
nor U11913 (N_11913,N_2948,N_5323);
nand U11914 (N_11914,N_2913,N_765);
nor U11915 (N_11915,N_1030,N_1467);
xor U11916 (N_11916,N_4902,N_2979);
nand U11917 (N_11917,N_5784,N_1676);
xor U11918 (N_11918,N_2570,N_3108);
nor U11919 (N_11919,N_1554,N_2421);
xor U11920 (N_11920,N_4834,N_2277);
xnor U11921 (N_11921,N_34,N_1243);
nand U11922 (N_11922,N_1148,N_3400);
nor U11923 (N_11923,N_4006,N_469);
nor U11924 (N_11924,N_1211,N_336);
nand U11925 (N_11925,N_5507,N_4192);
and U11926 (N_11926,N_2027,N_706);
and U11927 (N_11927,N_2485,N_4181);
nand U11928 (N_11928,N_512,N_703);
nor U11929 (N_11929,N_3022,N_5895);
nand U11930 (N_11930,N_5033,N_706);
and U11931 (N_11931,N_4353,N_4303);
nand U11932 (N_11932,N_4220,N_5807);
nand U11933 (N_11933,N_1024,N_2927);
or U11934 (N_11934,N_4274,N_184);
and U11935 (N_11935,N_5555,N_1873);
xor U11936 (N_11936,N_429,N_2084);
nor U11937 (N_11937,N_2689,N_1937);
and U11938 (N_11938,N_4821,N_45);
or U11939 (N_11939,N_5754,N_3677);
or U11940 (N_11940,N_102,N_3198);
or U11941 (N_11941,N_2178,N_5141);
and U11942 (N_11942,N_5691,N_5342);
or U11943 (N_11943,N_4035,N_4148);
and U11944 (N_11944,N_1244,N_4120);
xor U11945 (N_11945,N_319,N_1603);
and U11946 (N_11946,N_557,N_3328);
or U11947 (N_11947,N_2583,N_2563);
or U11948 (N_11948,N_2845,N_1345);
nand U11949 (N_11949,N_314,N_2678);
and U11950 (N_11950,N_5741,N_944);
xnor U11951 (N_11951,N_4261,N_4179);
nand U11952 (N_11952,N_1489,N_1464);
nor U11953 (N_11953,N_4808,N_5306);
nand U11954 (N_11954,N_1397,N_1899);
nor U11955 (N_11955,N_3718,N_959);
nand U11956 (N_11956,N_4609,N_2903);
xnor U11957 (N_11957,N_2030,N_2051);
or U11958 (N_11958,N_916,N_2835);
and U11959 (N_11959,N_3737,N_2137);
or U11960 (N_11960,N_5240,N_244);
xnor U11961 (N_11961,N_3808,N_5136);
or U11962 (N_11962,N_1191,N_4489);
nor U11963 (N_11963,N_5797,N_2176);
xor U11964 (N_11964,N_4926,N_2744);
nand U11965 (N_11965,N_1022,N_1718);
and U11966 (N_11966,N_2236,N_4662);
and U11967 (N_11967,N_1717,N_3183);
and U11968 (N_11968,N_3111,N_4198);
and U11969 (N_11969,N_1284,N_1365);
and U11970 (N_11970,N_4272,N_3973);
and U11971 (N_11971,N_3665,N_264);
nor U11972 (N_11972,N_2178,N_1691);
nand U11973 (N_11973,N_2106,N_1834);
and U11974 (N_11974,N_2930,N_3349);
and U11975 (N_11975,N_2028,N_4511);
xnor U11976 (N_11976,N_1825,N_4654);
and U11977 (N_11977,N_4979,N_2064);
xnor U11978 (N_11978,N_1191,N_5449);
or U11979 (N_11979,N_2833,N_4750);
or U11980 (N_11980,N_643,N_5661);
and U11981 (N_11981,N_273,N_3616);
nand U11982 (N_11982,N_5021,N_4721);
nor U11983 (N_11983,N_2353,N_3394);
and U11984 (N_11984,N_1973,N_1036);
xor U11985 (N_11985,N_2128,N_2916);
xor U11986 (N_11986,N_5012,N_733);
nor U11987 (N_11987,N_5011,N_4060);
nand U11988 (N_11988,N_1893,N_2106);
or U11989 (N_11989,N_2553,N_5074);
nor U11990 (N_11990,N_5621,N_5841);
nor U11991 (N_11991,N_2165,N_1955);
and U11992 (N_11992,N_5123,N_3561);
nor U11993 (N_11993,N_4013,N_1840);
xnor U11994 (N_11994,N_1731,N_2247);
xnor U11995 (N_11995,N_3380,N_1452);
nor U11996 (N_11996,N_5133,N_4665);
xor U11997 (N_11997,N_5307,N_1845);
nand U11998 (N_11998,N_3329,N_2674);
nor U11999 (N_11999,N_3625,N_4253);
nor U12000 (N_12000,N_9413,N_10047);
or U12001 (N_12001,N_6487,N_8490);
and U12002 (N_12002,N_7252,N_7320);
nor U12003 (N_12003,N_6167,N_11898);
nor U12004 (N_12004,N_11896,N_10495);
nor U12005 (N_12005,N_8838,N_11755);
and U12006 (N_12006,N_11719,N_11078);
xnor U12007 (N_12007,N_6283,N_11351);
nand U12008 (N_12008,N_10486,N_8286);
or U12009 (N_12009,N_7866,N_10348);
xnor U12010 (N_12010,N_7739,N_10819);
and U12011 (N_12011,N_7631,N_11260);
nand U12012 (N_12012,N_10343,N_11090);
or U12013 (N_12013,N_8377,N_10867);
nand U12014 (N_12014,N_10533,N_10192);
nand U12015 (N_12015,N_8319,N_6844);
or U12016 (N_12016,N_6701,N_10532);
xnor U12017 (N_12017,N_11235,N_11271);
xnor U12018 (N_12018,N_10810,N_6675);
nor U12019 (N_12019,N_9041,N_10604);
xnor U12020 (N_12020,N_6045,N_11190);
xor U12021 (N_12021,N_9404,N_11628);
or U12022 (N_12022,N_8106,N_11737);
or U12023 (N_12023,N_10124,N_10457);
nand U12024 (N_12024,N_9808,N_9957);
or U12025 (N_12025,N_11830,N_8924);
or U12026 (N_12026,N_9474,N_7239);
and U12027 (N_12027,N_6777,N_10657);
and U12028 (N_12028,N_9981,N_6307);
and U12029 (N_12029,N_10676,N_10099);
nand U12030 (N_12030,N_7568,N_7813);
nand U12031 (N_12031,N_10323,N_8040);
and U12032 (N_12032,N_7695,N_8442);
or U12033 (N_12033,N_6639,N_10718);
or U12034 (N_12034,N_8791,N_10918);
xnor U12035 (N_12035,N_9691,N_7335);
nor U12036 (N_12036,N_11786,N_11670);
or U12037 (N_12037,N_11988,N_10686);
or U12038 (N_12038,N_8648,N_10145);
nor U12039 (N_12039,N_11503,N_6989);
or U12040 (N_12040,N_11335,N_6747);
and U12041 (N_12041,N_6704,N_11552);
nor U12042 (N_12042,N_7597,N_8145);
xor U12043 (N_12043,N_7845,N_11821);
nor U12044 (N_12044,N_10159,N_8095);
nand U12045 (N_12045,N_9435,N_7445);
nand U12046 (N_12046,N_9279,N_7843);
nor U12047 (N_12047,N_6243,N_7170);
xor U12048 (N_12048,N_6696,N_6149);
or U12049 (N_12049,N_9677,N_7562);
and U12050 (N_12050,N_10366,N_8684);
xor U12051 (N_12051,N_7666,N_10120);
and U12052 (N_12052,N_10302,N_8797);
nand U12053 (N_12053,N_6444,N_11339);
and U12054 (N_12054,N_11826,N_6629);
or U12055 (N_12055,N_6948,N_10611);
nand U12056 (N_12056,N_10266,N_7167);
or U12057 (N_12057,N_11342,N_11903);
xnor U12058 (N_12058,N_8203,N_10478);
nor U12059 (N_12059,N_8258,N_6859);
nand U12060 (N_12060,N_11321,N_6199);
or U12061 (N_12061,N_9222,N_6402);
and U12062 (N_12062,N_6568,N_11020);
and U12063 (N_12063,N_9735,N_9513);
nand U12064 (N_12064,N_8772,N_7582);
or U12065 (N_12065,N_8630,N_7925);
or U12066 (N_12066,N_10947,N_11879);
nor U12067 (N_12067,N_11519,N_6168);
or U12068 (N_12068,N_8977,N_7990);
nand U12069 (N_12069,N_6713,N_7140);
xor U12070 (N_12070,N_10267,N_8333);
and U12071 (N_12071,N_7796,N_10950);
or U12072 (N_12072,N_8875,N_10948);
nand U12073 (N_12073,N_9718,N_10025);
nand U12074 (N_12074,N_6066,N_9436);
nand U12075 (N_12075,N_7916,N_11138);
nor U12076 (N_12076,N_10783,N_8813);
nor U12077 (N_12077,N_11851,N_9809);
or U12078 (N_12078,N_7962,N_8491);
or U12079 (N_12079,N_9382,N_8248);
xnor U12080 (N_12080,N_9768,N_11077);
nor U12081 (N_12081,N_10751,N_10815);
nand U12082 (N_12082,N_7852,N_7256);
and U12083 (N_12083,N_9873,N_11238);
xnor U12084 (N_12084,N_6228,N_10733);
xnor U12085 (N_12085,N_7920,N_10095);
and U12086 (N_12086,N_9673,N_10014);
nor U12087 (N_12087,N_7393,N_10545);
or U12088 (N_12088,N_8588,N_9487);
and U12089 (N_12089,N_9063,N_8998);
and U12090 (N_12090,N_11493,N_7757);
xnor U12091 (N_12091,N_6262,N_7483);
nand U12092 (N_12092,N_6575,N_9180);
nor U12093 (N_12093,N_10363,N_8762);
nor U12094 (N_12094,N_11840,N_8346);
xnor U12095 (N_12095,N_8614,N_7657);
xnor U12096 (N_12096,N_8511,N_11564);
nor U12097 (N_12097,N_6273,N_8800);
xnor U12098 (N_12098,N_11931,N_6560);
nand U12099 (N_12099,N_10537,N_10771);
nand U12100 (N_12100,N_7537,N_10445);
xor U12101 (N_12101,N_11723,N_8887);
or U12102 (N_12102,N_10905,N_6317);
nor U12103 (N_12103,N_11734,N_11150);
and U12104 (N_12104,N_8079,N_10572);
and U12105 (N_12105,N_6294,N_6740);
nand U12106 (N_12106,N_6947,N_7605);
nand U12107 (N_12107,N_7086,N_8602);
or U12108 (N_12108,N_10193,N_6897);
nor U12109 (N_12109,N_7290,N_10297);
or U12110 (N_12110,N_10487,N_6014);
or U12111 (N_12111,N_7197,N_9420);
and U12112 (N_12112,N_10855,N_10602);
nand U12113 (N_12113,N_8433,N_6248);
nor U12114 (N_12114,N_8649,N_9045);
and U12115 (N_12115,N_10491,N_11421);
nor U12116 (N_12116,N_11115,N_11960);
nor U12117 (N_12117,N_8489,N_10433);
nand U12118 (N_12118,N_7669,N_10835);
xor U12119 (N_12119,N_6174,N_10869);
xnor U12120 (N_12120,N_10494,N_11206);
xor U12121 (N_12121,N_6375,N_9592);
xnor U12122 (N_12122,N_6710,N_7204);
nand U12123 (N_12123,N_7224,N_7255);
xnor U12124 (N_12124,N_7128,N_8350);
nor U12125 (N_12125,N_7487,N_8352);
xor U12126 (N_12126,N_10345,N_9363);
xnor U12127 (N_12127,N_10017,N_10434);
nor U12128 (N_12128,N_11964,N_8856);
and U12129 (N_12129,N_7242,N_10121);
nand U12130 (N_12130,N_6417,N_10992);
and U12131 (N_12131,N_6870,N_7060);
xor U12132 (N_12132,N_8805,N_11127);
nand U12133 (N_12133,N_9203,N_11810);
nor U12134 (N_12134,N_7534,N_11071);
nand U12135 (N_12135,N_7720,N_7803);
nand U12136 (N_12136,N_8179,N_7510);
and U12137 (N_12137,N_9772,N_11914);
or U12138 (N_12138,N_11789,N_6043);
or U12139 (N_12139,N_6949,N_6345);
nand U12140 (N_12140,N_8228,N_9937);
or U12141 (N_12141,N_10253,N_8906);
and U12142 (N_12142,N_10032,N_7194);
nor U12143 (N_12143,N_11806,N_6546);
nand U12144 (N_12144,N_11853,N_11758);
and U12145 (N_12145,N_11813,N_6628);
nand U12146 (N_12146,N_7158,N_9411);
nand U12147 (N_12147,N_7323,N_9167);
and U12148 (N_12148,N_9200,N_7182);
nand U12149 (N_12149,N_7650,N_6792);
nand U12150 (N_12150,N_11736,N_6006);
or U12151 (N_12151,N_9270,N_7165);
nor U12152 (N_12152,N_10796,N_11153);
or U12153 (N_12153,N_8781,N_10091);
nor U12154 (N_12154,N_10483,N_6428);
or U12155 (N_12155,N_10560,N_7930);
or U12156 (N_12156,N_11200,N_8664);
or U12157 (N_12157,N_7895,N_10829);
xnor U12158 (N_12158,N_9428,N_11614);
and U12159 (N_12159,N_10632,N_11319);
nand U12160 (N_12160,N_9509,N_6980);
or U12161 (N_12161,N_11543,N_9380);
xor U12162 (N_12162,N_10268,N_8445);
nand U12163 (N_12163,N_7377,N_8240);
xnor U12164 (N_12164,N_11066,N_7826);
or U12165 (N_12165,N_8940,N_8195);
nand U12166 (N_12166,N_10142,N_10339);
xor U12167 (N_12167,N_9520,N_6434);
nor U12168 (N_12168,N_8970,N_7765);
nand U12169 (N_12169,N_6690,N_6994);
nand U12170 (N_12170,N_8871,N_7183);
nand U12171 (N_12171,N_10010,N_7791);
nand U12172 (N_12172,N_8972,N_7294);
nor U12173 (N_12173,N_8413,N_8733);
xor U12174 (N_12174,N_7509,N_11795);
nor U12175 (N_12175,N_10277,N_10135);
nor U12176 (N_12176,N_6440,N_10655);
or U12177 (N_12177,N_10938,N_6898);
or U12178 (N_12178,N_9986,N_9666);
xnor U12179 (N_12179,N_8361,N_10084);
nor U12180 (N_12180,N_7269,N_7913);
xor U12181 (N_12181,N_9726,N_6706);
nand U12182 (N_12182,N_6500,N_11815);
xnor U12183 (N_12183,N_9778,N_7091);
nand U12184 (N_12184,N_8168,N_10830);
xor U12185 (N_12185,N_8674,N_11094);
or U12186 (N_12186,N_9060,N_6462);
and U12187 (N_12187,N_8042,N_8638);
and U12188 (N_12188,N_11373,N_6025);
and U12189 (N_12189,N_11763,N_9886);
nand U12190 (N_12190,N_11465,N_11022);
nor U12191 (N_12191,N_10667,N_6902);
and U12192 (N_12192,N_6037,N_9439);
or U12193 (N_12193,N_10175,N_6674);
nand U12194 (N_12194,N_8290,N_6321);
nand U12195 (N_12195,N_9869,N_7907);
nor U12196 (N_12196,N_8349,N_7071);
nand U12197 (N_12197,N_9066,N_11188);
xnor U12198 (N_12198,N_9745,N_6324);
nor U12199 (N_12199,N_11175,N_7953);
and U12200 (N_12200,N_10238,N_7786);
nor U12201 (N_12201,N_10214,N_7363);
or U12202 (N_12202,N_8927,N_9202);
nor U12203 (N_12203,N_7237,N_8533);
or U12204 (N_12204,N_11247,N_11143);
and U12205 (N_12205,N_11113,N_9996);
and U12206 (N_12206,N_9843,N_11461);
nand U12207 (N_12207,N_8916,N_6769);
nor U12208 (N_12208,N_7019,N_10720);
and U12209 (N_12209,N_8971,N_11298);
or U12210 (N_12210,N_8129,N_10273);
nand U12211 (N_12211,N_10332,N_6825);
xor U12212 (N_12212,N_6064,N_8153);
and U12213 (N_12213,N_9391,N_11360);
nand U12214 (N_12214,N_6123,N_6745);
nand U12215 (N_12215,N_6954,N_6178);
and U12216 (N_12216,N_6193,N_7297);
and U12217 (N_12217,N_10616,N_6935);
nand U12218 (N_12218,N_10984,N_9348);
nand U12219 (N_12219,N_11831,N_8462);
nor U12220 (N_12220,N_10850,N_11386);
and U12221 (N_12221,N_11192,N_8735);
and U12222 (N_12222,N_6712,N_9695);
xor U12223 (N_12223,N_6315,N_9959);
and U12224 (N_12224,N_8915,N_10104);
nand U12225 (N_12225,N_9774,N_9727);
nand U12226 (N_12226,N_6351,N_7641);
nand U12227 (N_12227,N_10558,N_7589);
and U12228 (N_12228,N_6197,N_10516);
and U12229 (N_12229,N_6737,N_6219);
and U12230 (N_12230,N_11366,N_6565);
or U12231 (N_12231,N_8383,N_10407);
and U12232 (N_12232,N_10702,N_8751);
nand U12233 (N_12233,N_6079,N_9241);
xnor U12234 (N_12234,N_6015,N_8356);
nor U12235 (N_12235,N_9795,N_6000);
nor U12236 (N_12236,N_8303,N_8789);
xnor U12237 (N_12237,N_7917,N_11654);
and U12238 (N_12238,N_8102,N_7577);
or U12239 (N_12239,N_7213,N_10936);
xor U12240 (N_12240,N_9507,N_8635);
or U12241 (N_12241,N_8398,N_8298);
nand U12242 (N_12242,N_8773,N_11476);
and U12243 (N_12243,N_10841,N_11820);
and U12244 (N_12244,N_10391,N_10524);
nor U12245 (N_12245,N_7690,N_9237);
or U12246 (N_12246,N_9175,N_10708);
and U12247 (N_12247,N_11932,N_9033);
xor U12248 (N_12248,N_10717,N_8914);
xnor U12249 (N_12249,N_11054,N_8718);
nor U12250 (N_12250,N_8764,N_10644);
and U12251 (N_12251,N_10534,N_7730);
or U12252 (N_12252,N_10319,N_10557);
xor U12253 (N_12253,N_10417,N_6403);
xnor U12254 (N_12254,N_9582,N_10400);
xnor U12255 (N_12255,N_8200,N_7939);
or U12256 (N_12256,N_10776,N_11578);
nand U12257 (N_12257,N_9909,N_9248);
or U12258 (N_12258,N_9193,N_8339);
nand U12259 (N_12259,N_9883,N_10744);
nand U12260 (N_12260,N_7463,N_7176);
or U12261 (N_12261,N_8320,N_7570);
or U12262 (N_12262,N_6218,N_8645);
nor U12263 (N_12263,N_11495,N_9417);
nand U12264 (N_12264,N_6781,N_9295);
xor U12265 (N_12265,N_10249,N_6888);
or U12266 (N_12266,N_9186,N_10974);
nor U12267 (N_12267,N_9668,N_7051);
or U12268 (N_12268,N_8341,N_6975);
nor U12269 (N_12269,N_6304,N_8204);
nand U12270 (N_12270,N_11527,N_8162);
and U12271 (N_12271,N_7877,N_11929);
xnor U12272 (N_12272,N_11742,N_7081);
nor U12273 (N_12273,N_11207,N_10995);
and U12274 (N_12274,N_8394,N_9120);
and U12275 (N_12275,N_6453,N_9553);
xor U12276 (N_12276,N_8231,N_6636);
and U12277 (N_12277,N_7688,N_6343);
xor U12278 (N_12278,N_6528,N_9347);
and U12279 (N_12279,N_10186,N_10797);
nand U12280 (N_12280,N_10031,N_9081);
xor U12281 (N_12281,N_9438,N_9729);
nor U12282 (N_12282,N_9731,N_7890);
xor U12283 (N_12283,N_10668,N_6072);
or U12284 (N_12284,N_6973,N_9263);
and U12285 (N_12285,N_10619,N_6320);
nand U12286 (N_12286,N_7685,N_6976);
xor U12287 (N_12287,N_10853,N_8725);
xnor U12288 (N_12288,N_6939,N_7614);
xor U12289 (N_12289,N_7681,N_6067);
or U12290 (N_12290,N_10975,N_7879);
nand U12291 (N_12291,N_9770,N_11909);
and U12292 (N_12292,N_7623,N_11318);
nor U12293 (N_12293,N_9521,N_6758);
or U12294 (N_12294,N_6081,N_11458);
xnor U12295 (N_12295,N_7417,N_10581);
nand U12296 (N_12296,N_9050,N_9112);
and U12297 (N_12297,N_10097,N_10069);
and U12298 (N_12298,N_6438,N_8568);
and U12299 (N_12299,N_10052,N_10139);
nand U12300 (N_12300,N_9458,N_11405);
xnor U12301 (N_12301,N_9523,N_10264);
and U12302 (N_12302,N_10048,N_10168);
nand U12303 (N_12303,N_8532,N_9389);
or U12304 (N_12304,N_6786,N_6926);
nand U12305 (N_12305,N_9094,N_8090);
or U12306 (N_12306,N_11715,N_9003);
and U12307 (N_12307,N_9540,N_6799);
xnor U12308 (N_12308,N_7817,N_11456);
nand U12309 (N_12309,N_9123,N_11656);
nor U12310 (N_12310,N_7531,N_9586);
and U12311 (N_12311,N_8613,N_7659);
and U12312 (N_12312,N_8175,N_6141);
nand U12313 (N_12313,N_6863,N_10228);
nor U12314 (N_12314,N_8721,N_6279);
xnor U12315 (N_12315,N_9035,N_8870);
xor U12316 (N_12316,N_7202,N_8246);
nor U12317 (N_12317,N_8889,N_8880);
xnor U12318 (N_12318,N_11973,N_8712);
xnor U12319 (N_12319,N_6454,N_9701);
nand U12320 (N_12320,N_10926,N_6288);
and U12321 (N_12321,N_11477,N_10247);
or U12322 (N_12322,N_11357,N_6614);
or U12323 (N_12323,N_8318,N_9785);
or U12324 (N_12324,N_6676,N_11387);
and U12325 (N_12325,N_8708,N_7760);
nand U12326 (N_12326,N_10555,N_7234);
nand U12327 (N_12327,N_9629,N_6012);
nor U12328 (N_12328,N_9385,N_10358);
nand U12329 (N_12329,N_11509,N_11391);
nand U12330 (N_12330,N_9676,N_11327);
nor U12331 (N_12331,N_8601,N_9792);
nand U12332 (N_12332,N_7017,N_7085);
nor U12333 (N_12333,N_11496,N_10456);
nand U12334 (N_12334,N_8795,N_7538);
or U12335 (N_12335,N_6915,N_7119);
or U12336 (N_12336,N_9303,N_11487);
nand U12337 (N_12337,N_10996,N_7495);
xnor U12338 (N_12338,N_6780,N_7686);
xnor U12339 (N_12339,N_6641,N_9495);
or U12340 (N_12340,N_6734,N_7196);
nand U12341 (N_12341,N_8355,N_7478);
nor U12342 (N_12342,N_9921,N_7310);
nor U12343 (N_12343,N_9512,N_10226);
and U12344 (N_12344,N_8653,N_9848);
nand U12345 (N_12345,N_10133,N_6765);
nor U12346 (N_12346,N_7099,N_6435);
or U12347 (N_12347,N_9034,N_7228);
or U12348 (N_12348,N_8798,N_7160);
nor U12349 (N_12349,N_10146,N_8405);
xnor U12350 (N_12350,N_11145,N_6291);
or U12351 (N_12351,N_8218,N_6512);
nand U12352 (N_12352,N_10563,N_9433);
nor U12353 (N_12353,N_7192,N_8408);
or U12354 (N_12354,N_10500,N_8873);
nand U12355 (N_12355,N_11292,N_7475);
or U12356 (N_12356,N_11839,N_9658);
nor U12357 (N_12357,N_11035,N_8211);
and U12358 (N_12358,N_6689,N_10707);
and U12359 (N_12359,N_9920,N_8714);
or U12360 (N_12360,N_9854,N_10106);
and U12361 (N_12361,N_8858,N_11924);
xor U12362 (N_12362,N_11764,N_9758);
and U12363 (N_12363,N_10162,N_9434);
nand U12364 (N_12364,N_11144,N_9409);
or U12365 (N_12365,N_11595,N_10399);
or U12366 (N_12366,N_11666,N_9269);
and U12367 (N_12367,N_10397,N_11384);
and U12368 (N_12368,N_9675,N_8606);
nor U12369 (N_12369,N_11655,N_11286);
or U12370 (N_12370,N_11513,N_9122);
nor U12371 (N_12371,N_7752,N_6480);
nand U12372 (N_12372,N_6984,N_6756);
nor U12373 (N_12373,N_6388,N_8809);
or U12374 (N_12374,N_6760,N_7807);
nor U12375 (N_12375,N_9752,N_7714);
nor U12376 (N_12376,N_7231,N_7494);
nor U12377 (N_12377,N_7079,N_6937);
nor U12378 (N_12378,N_9682,N_8487);
nor U12379 (N_12379,N_7087,N_10489);
nor U12380 (N_12380,N_7387,N_11007);
nor U12381 (N_12381,N_10326,N_11678);
xor U12382 (N_12382,N_6159,N_10592);
and U12383 (N_12383,N_9925,N_10933);
nand U12384 (N_12384,N_7117,N_11662);
or U12385 (N_12385,N_9178,N_7512);
and U12386 (N_12386,N_8522,N_8549);
nor U12387 (N_12387,N_8159,N_11307);
xor U12388 (N_12388,N_9543,N_11852);
or U12389 (N_12389,N_9723,N_11289);
xor U12390 (N_12390,N_6295,N_9220);
or U12391 (N_12391,N_7472,N_7676);
and U12392 (N_12392,N_11548,N_7347);
xnor U12393 (N_12393,N_7958,N_11951);
nor U12394 (N_12394,N_10254,N_11334);
nand U12395 (N_12395,N_6257,N_11180);
nand U12396 (N_12396,N_9659,N_8437);
nor U12397 (N_12397,N_8205,N_10617);
nor U12398 (N_12398,N_11096,N_6941);
nor U12399 (N_12399,N_11123,N_8284);
and U12400 (N_12400,N_9335,N_10077);
nand U12401 (N_12401,N_6795,N_9575);
and U12402 (N_12402,N_8595,N_6856);
nor U12403 (N_12403,N_8883,N_10654);
and U12404 (N_12404,N_9650,N_9631);
xor U12405 (N_12405,N_8172,N_7084);
nor U12406 (N_12406,N_6789,N_9860);
xnor U12407 (N_12407,N_6415,N_6549);
and U12408 (N_12408,N_10394,N_7761);
nand U12409 (N_12409,N_8103,N_11752);
nand U12410 (N_12410,N_8086,N_6269);
nor U12411 (N_12411,N_10136,N_8982);
xnor U12412 (N_12412,N_8265,N_9005);
nor U12413 (N_12413,N_6996,N_7013);
or U12414 (N_12414,N_6196,N_10356);
nor U12415 (N_12415,N_11234,N_11488);
and U12416 (N_12416,N_7222,N_8446);
nor U12417 (N_12417,N_6865,N_8860);
nor U12418 (N_12418,N_6718,N_6604);
nor U12419 (N_12419,N_6068,N_7299);
nand U12420 (N_12420,N_8990,N_9845);
nand U12421 (N_12421,N_10743,N_10012);
xor U12422 (N_12422,N_11051,N_11198);
nor U12423 (N_12423,N_6717,N_11316);
xnor U12424 (N_12424,N_6313,N_6903);
nor U12425 (N_12425,N_11404,N_11649);
and U12426 (N_12426,N_10740,N_11520);
xnor U12427 (N_12427,N_7704,N_11184);
nand U12428 (N_12428,N_11599,N_8697);
xnor U12429 (N_12429,N_8119,N_10252);
and U12430 (N_12430,N_8569,N_9661);
nand U12431 (N_12431,N_7578,N_11379);
nor U12432 (N_12432,N_10941,N_7642);
nor U12433 (N_12433,N_9155,N_9781);
xnor U12434 (N_12434,N_9058,N_6494);
xor U12435 (N_12435,N_7089,N_7069);
xor U12436 (N_12436,N_7558,N_11221);
xnor U12437 (N_12437,N_11858,N_7726);
xnor U12438 (N_12438,N_6848,N_10503);
and U12439 (N_12439,N_10325,N_7206);
nand U12440 (N_12440,N_8308,N_9036);
nor U12441 (N_12441,N_6818,N_8957);
xnor U12442 (N_12442,N_11709,N_10894);
xnor U12443 (N_12443,N_7652,N_9206);
xor U12444 (N_12444,N_6801,N_8903);
xnor U12445 (N_12445,N_10837,N_6490);
and U12446 (N_12446,N_10351,N_9622);
or U12447 (N_12447,N_10535,N_8967);
xor U12448 (N_12448,N_8024,N_11032);
and U12449 (N_12449,N_7661,N_11486);
nor U12450 (N_12450,N_9462,N_10210);
nor U12451 (N_12451,N_7932,N_7973);
nor U12452 (N_12452,N_7049,N_8615);
xnor U12453 (N_12453,N_11783,N_11243);
nor U12454 (N_12454,N_8215,N_6110);
and U12455 (N_12455,N_9480,N_9009);
xor U12456 (N_12456,N_9977,N_11120);
or U12457 (N_12457,N_10785,N_6693);
xnor U12458 (N_12458,N_11972,N_9106);
xnor U12459 (N_12459,N_10647,N_10150);
nor U12460 (N_12460,N_9634,N_6601);
nand U12461 (N_12461,N_9604,N_10123);
nand U12462 (N_12462,N_11510,N_9266);
nand U12463 (N_12463,N_7812,N_8104);
nor U12464 (N_12464,N_10362,N_10767);
xor U12465 (N_12465,N_8301,N_11660);
xor U12466 (N_12466,N_10514,N_9093);
xnor U12467 (N_12467,N_9281,N_11099);
xor U12468 (N_12468,N_7104,N_8699);
xnor U12469 (N_12469,N_7448,N_7198);
and U12470 (N_12470,N_7126,N_6680);
or U12471 (N_12471,N_9580,N_7763);
xor U12472 (N_12472,N_10396,N_10704);
nor U12473 (N_12473,N_9061,N_7378);
and U12474 (N_12474,N_10416,N_7798);
xnor U12475 (N_12475,N_6504,N_9097);
nand U12476 (N_12476,N_10736,N_8075);
xor U12477 (N_12477,N_11639,N_6593);
nor U12478 (N_12478,N_11952,N_8707);
nor U12479 (N_12479,N_10278,N_6100);
or U12480 (N_12480,N_11607,N_11374);
nand U12481 (N_12481,N_8894,N_7970);
nor U12482 (N_12482,N_8156,N_10927);
nor U12483 (N_12483,N_10270,N_10115);
nand U12484 (N_12484,N_11470,N_10475);
xnor U12485 (N_12485,N_11833,N_8582);
nand U12486 (N_12486,N_11001,N_11888);
nand U12487 (N_12487,N_9847,N_9457);
nor U12488 (N_12488,N_10335,N_6626);
xnor U12489 (N_12489,N_9762,N_10481);
and U12490 (N_12490,N_10479,N_10909);
or U12491 (N_12491,N_10364,N_6239);
and U12492 (N_12492,N_8477,N_6361);
xnor U12493 (N_12493,N_11257,N_8315);
nor U12494 (N_12494,N_10515,N_10287);
nand U12495 (N_12495,N_6331,N_8192);
or U12496 (N_12496,N_9573,N_6927);
xnor U12497 (N_12497,N_8942,N_6905);
and U12498 (N_12498,N_10626,N_6923);
or U12499 (N_12499,N_6842,N_6586);
nor U12500 (N_12500,N_8661,N_11163);
or U12501 (N_12501,N_10111,N_9316);
or U12502 (N_12502,N_11686,N_7241);
or U12503 (N_12503,N_6702,N_10113);
xor U12504 (N_12504,N_6344,N_7712);
nand U12505 (N_12505,N_7395,N_9092);
nor U12506 (N_12506,N_6893,N_6305);
nor U12507 (N_12507,N_11098,N_8249);
nor U12508 (N_12508,N_9953,N_8815);
nor U12509 (N_12509,N_7179,N_7557);
or U12510 (N_12510,N_9223,N_8263);
or U12511 (N_12511,N_6040,N_11895);
nor U12512 (N_12512,N_7508,N_9779);
nand U12513 (N_12513,N_11516,N_6506);
nor U12514 (N_12514,N_7032,N_8585);
and U12515 (N_12515,N_8583,N_10056);
or U12516 (N_12516,N_7217,N_11962);
nor U12517 (N_12517,N_9326,N_7426);
or U12518 (N_12518,N_8807,N_11353);
xor U12519 (N_12519,N_6249,N_7358);
nand U12520 (N_12520,N_10890,N_7599);
and U12521 (N_12521,N_7208,N_10468);
nand U12522 (N_12522,N_7602,N_8694);
and U12523 (N_12523,N_8482,N_7571);
or U12524 (N_12524,N_9288,N_8986);
xnor U12525 (N_12525,N_6314,N_7880);
and U12526 (N_12526,N_9199,N_8229);
nand U12527 (N_12527,N_7556,N_7579);
and U12528 (N_12528,N_6325,N_8015);
nand U12529 (N_12529,N_8780,N_9246);
nand U12530 (N_12530,N_8828,N_7264);
nand U12531 (N_12531,N_7754,N_10805);
xor U12532 (N_12532,N_11563,N_11355);
xor U12533 (N_12533,N_7014,N_8814);
nand U12534 (N_12534,N_11086,N_9133);
and U12535 (N_12535,N_6406,N_7995);
or U12536 (N_12536,N_6545,N_9642);
and U12537 (N_12537,N_6194,N_11602);
or U12538 (N_12538,N_9587,N_9109);
xor U12539 (N_12539,N_7595,N_9214);
nand U12540 (N_12540,N_11919,N_9500);
nor U12541 (N_12541,N_7643,N_11799);
xnor U12542 (N_12542,N_11976,N_7368);
and U12543 (N_12543,N_11729,N_9032);
nand U12544 (N_12544,N_7365,N_7526);
or U12545 (N_12545,N_8586,N_8461);
xnor U12546 (N_12546,N_8336,N_11793);
xor U12547 (N_12547,N_10912,N_8472);
xor U12548 (N_12548,N_8151,N_7078);
nor U12549 (N_12549,N_7729,N_6052);
xnor U12550 (N_12550,N_9697,N_6211);
nor U12551 (N_12551,N_7164,N_9684);
or U12552 (N_12552,N_6475,N_10379);
nand U12553 (N_12553,N_7040,N_8335);
and U12554 (N_12554,N_10485,N_7043);
and U12555 (N_12555,N_11092,N_10161);
nor U12556 (N_12556,N_11659,N_6379);
nor U12557 (N_12557,N_9049,N_10715);
and U12558 (N_12558,N_10692,N_10221);
or U12559 (N_12559,N_6468,N_7784);
nand U12560 (N_12560,N_7677,N_7804);
and U12561 (N_12561,N_10036,N_10672);
nor U12562 (N_12562,N_6121,N_7076);
nor U12563 (N_12563,N_10887,N_9317);
xnor U12564 (N_12564,N_9482,N_6093);
nand U12565 (N_12565,N_10251,N_7027);
nor U12566 (N_12566,N_8304,N_8907);
nor U12567 (N_12567,N_7507,N_11166);
xor U12568 (N_12568,N_8074,N_11440);
xor U12569 (N_12569,N_11721,N_9796);
or U12570 (N_12570,N_7163,N_9278);
xnor U12571 (N_12571,N_8251,N_7471);
xor U12572 (N_12572,N_6882,N_10999);
nand U12573 (N_12573,N_10143,N_10051);
nand U12574 (N_12574,N_7864,N_11756);
nor U12575 (N_12575,N_10066,N_8963);
and U12576 (N_12576,N_8801,N_8219);
xor U12577 (N_12577,N_11154,N_8239);
xnor U12578 (N_12578,N_7540,N_10004);
or U12579 (N_12579,N_10447,N_10127);
nand U12580 (N_12580,N_8732,N_8953);
xnor U12581 (N_12581,N_7731,N_7909);
nor U12582 (N_12582,N_6499,N_7572);
and U12583 (N_12583,N_7357,N_7893);
nand U12584 (N_12584,N_10641,N_10615);
nor U12585 (N_12585,N_9182,N_6441);
nor U12586 (N_12586,N_7074,N_10937);
nor U12587 (N_12587,N_6097,N_8245);
or U12588 (N_12588,N_6967,N_6522);
and U12589 (N_12589,N_10299,N_10005);
nand U12590 (N_12590,N_8622,N_8403);
and U12591 (N_12591,N_10295,N_7173);
nand U12592 (N_12592,N_7713,N_9381);
or U12593 (N_12593,N_9447,N_11525);
and U12594 (N_12594,N_6311,N_8786);
and U12595 (N_12595,N_6505,N_9027);
or U12596 (N_12596,N_11164,N_10750);
or U12597 (N_12597,N_8518,N_11957);
nand U12598 (N_12598,N_11226,N_9862);
nand U12599 (N_12599,N_7783,N_10690);
nand U12600 (N_12600,N_11224,N_8382);
nand U12601 (N_12601,N_7671,N_6991);
or U12602 (N_12602,N_8765,N_7191);
nor U12603 (N_12603,N_9361,N_8509);
nand U12604 (N_12604,N_8317,N_11645);
nor U12605 (N_12605,N_6683,N_7746);
xor U12606 (N_12606,N_9185,N_8665);
xnor U12607 (N_12607,N_10752,N_10645);
xor U12608 (N_12608,N_9351,N_7102);
nand U12609 (N_12609,N_10068,N_10454);
nor U12610 (N_12610,N_7574,N_8539);
nand U12611 (N_12611,N_7115,N_7833);
nand U12612 (N_12612,N_11518,N_11553);
nor U12613 (N_12613,N_11982,N_7585);
nand U12614 (N_12614,N_7200,N_11778);
nor U12615 (N_12615,N_10280,N_8763);
or U12616 (N_12616,N_6833,N_7298);
or U12617 (N_12617,N_11565,N_10341);
nor U12618 (N_12618,N_6556,N_6547);
or U12619 (N_12619,N_9952,N_7892);
or U12620 (N_12620,N_8851,N_8096);
and U12621 (N_12621,N_7952,N_6038);
nor U12622 (N_12622,N_9903,N_6117);
xor U12623 (N_12623,N_7042,N_11848);
nor U12624 (N_12624,N_11522,N_10211);
and U12625 (N_12625,N_8076,N_9431);
nand U12626 (N_12626,N_9424,N_9557);
nor U12627 (N_12627,N_10714,N_10412);
and U12628 (N_12628,N_8223,N_11274);
or U12629 (N_12629,N_8748,N_10824);
or U12630 (N_12630,N_9354,N_8479);
nand U12631 (N_12631,N_11610,N_11978);
nor U12632 (N_12632,N_8425,N_6296);
or U12633 (N_12633,N_10816,N_9046);
or U12634 (N_12634,N_8234,N_7919);
nor U12635 (N_12635,N_10034,N_11255);
or U12636 (N_12636,N_8407,N_9709);
xor U12637 (N_12637,N_10223,N_9606);
nand U12638 (N_12638,N_6360,N_8527);
nor U12639 (N_12639,N_11170,N_9946);
and U12640 (N_12640,N_6474,N_7246);
nor U12641 (N_12641,N_11288,N_10795);
nand U12642 (N_12642,N_9824,N_9990);
xnor U12643 (N_12643,N_6771,N_7878);
xnor U12644 (N_12644,N_8334,N_8073);
and U12645 (N_12645,N_10309,N_10862);
xnor U12646 (N_12646,N_9565,N_6207);
nor U12647 (N_12647,N_10016,N_6112);
nor U12648 (N_12648,N_11886,N_8418);
or U12649 (N_12649,N_7143,N_10782);
xnor U12650 (N_12650,N_7157,N_7185);
xnor U12651 (N_12651,N_6150,N_6383);
nor U12652 (N_12652,N_9352,N_7349);
or U12653 (N_12653,N_8170,N_6019);
xor U12654 (N_12654,N_7797,N_7535);
xnor U12655 (N_12655,N_10474,N_11883);
and U12656 (N_12656,N_7756,N_6192);
nand U12657 (N_12657,N_7831,N_11884);
nand U12658 (N_12658,N_6059,N_10122);
and U12659 (N_12659,N_7905,N_10562);
xor U12660 (N_12660,N_9116,N_11768);
xor U12661 (N_12661,N_6534,N_6312);
or U12662 (N_12662,N_11068,N_9449);
or U12663 (N_12663,N_9670,N_7061);
nor U12664 (N_12664,N_8655,N_11530);
xor U12665 (N_12665,N_9755,N_7984);
nor U12666 (N_12666,N_11483,N_10803);
nor U12667 (N_12667,N_9628,N_6722);
nor U12668 (N_12668,N_8143,N_8570);
nand U12669 (N_12669,N_9224,N_6819);
xnor U12670 (N_12670,N_8166,N_11393);
xnor U12671 (N_12671,N_9426,N_9712);
nand U12672 (N_12672,N_8078,N_10990);
nand U12673 (N_12673,N_9329,N_9441);
nor U12674 (N_12674,N_8577,N_9932);
nand U12675 (N_12675,N_10711,N_9008);
xor U12676 (N_12676,N_7247,N_7521);
or U12677 (N_12677,N_10605,N_7401);
nor U12678 (N_12678,N_7132,N_6686);
and U12679 (N_12679,N_7964,N_7147);
xnor U12680 (N_12680,N_10942,N_9819);
nor U12681 (N_12681,N_7549,N_8935);
nand U12682 (N_12682,N_11017,N_10245);
nor U12683 (N_12683,N_8089,N_10152);
or U12684 (N_12684,N_10958,N_6763);
nor U12685 (N_12685,N_6585,N_11936);
or U12686 (N_12686,N_11236,N_8130);
nand U12687 (N_12687,N_10291,N_11993);
nor U12688 (N_12688,N_7004,N_11312);
nor U12689 (N_12689,N_7388,N_11638);
nand U12690 (N_12690,N_8904,N_10141);
or U12691 (N_12691,N_8590,N_6826);
or U12692 (N_12692,N_10039,N_7697);
nor U12693 (N_12693,N_10140,N_10373);
nor U12694 (N_12694,N_9325,N_6143);
nand U12695 (N_12695,N_8125,N_11983);
xor U12696 (N_12696,N_8531,N_11691);
or U12697 (N_12697,N_8464,N_6655);
or U12698 (N_12698,N_9085,N_10438);
nand U12699 (N_12699,N_9310,N_9473);
and U12700 (N_12700,N_10614,N_9219);
nand U12701 (N_12701,N_9338,N_8850);
xor U12702 (N_12702,N_7453,N_7929);
or U12703 (N_12703,N_7664,N_11524);
and U12704 (N_12704,N_11861,N_10449);
and U12705 (N_12705,N_6009,N_6581);
nand U12706 (N_12706,N_9825,N_7046);
and U12707 (N_12707,N_10892,N_11211);
and U12708 (N_12708,N_6552,N_9962);
xnor U12709 (N_12709,N_11843,N_6945);
and U12710 (N_12710,N_7050,N_10257);
or U12711 (N_12711,N_11774,N_9465);
nor U12712 (N_12712,N_11997,N_7141);
xor U12713 (N_12713,N_10808,N_8560);
nand U12714 (N_12714,N_11572,N_9827);
nor U12715 (N_12715,N_8727,N_9941);
or U12716 (N_12716,N_7819,N_10721);
nor U12717 (N_12717,N_9072,N_6004);
xor U12718 (N_12718,N_9961,N_6963);
or U12719 (N_12719,N_10344,N_9970);
or U12720 (N_12720,N_7258,N_10908);
and U12721 (N_12721,N_9013,N_10109);
xor U12722 (N_12722,N_8022,N_9599);
and U12723 (N_12723,N_7300,N_10380);
and U12724 (N_12724,N_11121,N_8965);
nor U12725 (N_12725,N_10801,N_9312);
and U12726 (N_12726,N_10336,N_11232);
xnor U12727 (N_12727,N_7301,N_6472);
nor U12728 (N_12728,N_10110,N_9368);
or U12729 (N_12729,N_7774,N_10684);
nand U12730 (N_12730,N_8656,N_9196);
or U12731 (N_12731,N_7956,N_9802);
nor U12732 (N_12732,N_10746,N_11508);
or U12733 (N_12733,N_10506,N_11859);
nor U12734 (N_12734,N_11279,N_6607);
and U12735 (N_12735,N_8756,N_11208);
nor U12736 (N_12736,N_10989,N_6368);
nor U12737 (N_12737,N_11004,N_10346);
nor U12738 (N_12738,N_8138,N_6238);
xnor U12739 (N_12739,N_8663,N_7470);
and U12740 (N_12740,N_11055,N_10768);
nand U12741 (N_12741,N_11060,N_10849);
and U12742 (N_12742,N_11336,N_10747);
nand U12743 (N_12743,N_8703,N_7021);
or U12744 (N_12744,N_8537,N_10105);
xnor U12745 (N_12745,N_10664,N_7809);
xnor U12746 (N_12746,N_7721,N_10998);
and U12747 (N_12747,N_9100,N_11812);
nand U12748 (N_12748,N_9715,N_8344);
nor U12749 (N_12749,N_8591,N_11281);
or U12750 (N_12750,N_7354,N_10547);
or U12751 (N_12751,N_10969,N_7856);
or U12752 (N_12752,N_11220,N_8270);
and U12753 (N_12753,N_11775,N_9488);
nor U12754 (N_12754,N_6750,N_8559);
or U12755 (N_12755,N_7172,N_6334);
xor U12756 (N_12756,N_6377,N_6850);
and U12757 (N_12757,N_9313,N_8794);
nand U12758 (N_12758,N_11681,N_6061);
and U12759 (N_12759,N_6214,N_11966);
or U12760 (N_12760,N_10821,N_6483);
xor U12761 (N_12761,N_9387,N_10265);
or U12762 (N_12762,N_7541,N_9605);
nand U12763 (N_12763,N_7719,N_9950);
nor U12764 (N_12764,N_8724,N_8475);
nand U12765 (N_12765,N_8989,N_9154);
nor U12766 (N_12766,N_11642,N_10167);
or U12767 (N_12767,N_7443,N_10035);
nand U12768 (N_12768,N_7260,N_9885);
xor U12769 (N_12769,N_11773,N_9780);
nand U12770 (N_12770,N_9829,N_9588);
nor U12771 (N_12771,N_7122,N_8799);
or U12772 (N_12772,N_9552,N_9922);
or U12773 (N_12773,N_8679,N_9442);
or U12774 (N_12774,N_6743,N_7897);
or U12775 (N_12775,N_8323,N_10383);
and U12776 (N_12776,N_6142,N_10101);
nor U12777 (N_12777,N_7997,N_11634);
xnor U12778 (N_12778,N_8621,N_8137);
nor U12779 (N_12779,N_8342,N_8572);
and U12780 (N_12780,N_8702,N_9602);
or U12781 (N_12781,N_6988,N_10972);
nand U12782 (N_12782,N_9468,N_11028);
nor U12783 (N_12783,N_6635,N_8267);
or U12784 (N_12784,N_6306,N_9832);
xnor U12785 (N_12785,N_7983,N_10838);
nand U12786 (N_12786,N_10184,N_11481);
xor U12787 (N_12787,N_7352,N_10112);
nand U12788 (N_12788,N_6862,N_11986);
nand U12789 (N_12789,N_11651,N_9235);
nand U12790 (N_12790,N_8521,N_8278);
nor U12791 (N_12791,N_6620,N_6050);
and U12792 (N_12792,N_9451,N_6060);
or U12793 (N_12793,N_6978,N_6153);
or U12794 (N_12794,N_10931,N_9463);
and U12795 (N_12795,N_8092,N_8080);
or U12796 (N_12796,N_9026,N_6492);
nand U12797 (N_12797,N_10330,N_7612);
nor U12798 (N_12798,N_6764,N_10386);
nand U12799 (N_12799,N_7386,N_6757);
nand U12800 (N_12800,N_7111,N_6102);
xnor U12801 (N_12801,N_11676,N_6424);
xnor U12802 (N_12802,N_11471,N_10842);
nor U12803 (N_12803,N_6564,N_6362);
nor U12804 (N_12804,N_9807,N_11928);
xnor U12805 (N_12805,N_7454,N_9838);
nor U12806 (N_12806,N_8910,N_6527);
and U12807 (N_12807,N_7918,N_11245);
nand U12808 (N_12808,N_6230,N_11354);
and U12809 (N_12809,N_6866,N_11575);
and U12810 (N_12810,N_9088,N_10589);
or U12811 (N_12811,N_6503,N_6420);
or U12812 (N_12812,N_11213,N_11744);
xnor U12813 (N_12813,N_9861,N_8181);
and U12814 (N_12814,N_8576,N_6754);
nor U12815 (N_12815,N_10866,N_10156);
or U12816 (N_12816,N_6521,N_11864);
and U12817 (N_12817,N_11125,N_8366);
xor U12818 (N_12818,N_8247,N_6465);
or U12819 (N_12819,N_9078,N_11269);
and U12820 (N_12820,N_8608,N_10597);
or U12821 (N_12821,N_11942,N_10965);
nor U12822 (N_12822,N_6516,N_8208);
and U12823 (N_12823,N_11772,N_9654);
or U12824 (N_12824,N_8255,N_8534);
nor U12825 (N_12825,N_6698,N_10467);
or U12826 (N_12826,N_6971,N_11058);
nand U12827 (N_12827,N_11801,N_10024);
nor U12828 (N_12828,N_7211,N_8455);
xor U12829 (N_12829,N_11796,N_9669);
xor U12830 (N_12830,N_10760,N_9344);
xor U12831 (N_12831,N_10847,N_10452);
and U12832 (N_12832,N_10194,N_8643);
nor U12833 (N_12833,N_9461,N_11911);
nor U12834 (N_12834,N_9083,N_8438);
nand U12835 (N_12835,N_11403,N_11700);
nand U12836 (N_12836,N_9390,N_8639);
or U12837 (N_12837,N_11368,N_7616);
nor U12838 (N_12838,N_11383,N_7942);
xor U12839 (N_12839,N_6401,N_7134);
xnor U12840 (N_12840,N_10300,N_8014);
nor U12841 (N_12841,N_6553,N_10274);
nand U12842 (N_12842,N_7658,N_6633);
and U12843 (N_12843,N_9362,N_11937);
xnor U12844 (N_12844,N_10536,N_9498);
nor U12845 (N_12845,N_10565,N_8347);
and U12846 (N_12846,N_7883,N_10612);
or U12847 (N_12847,N_7284,N_6161);
and U12848 (N_12848,N_7699,N_9662);
nand U12849 (N_12849,N_9965,N_6887);
nand U12850 (N_12850,N_9623,N_10823);
and U12851 (N_12851,N_8612,N_9080);
nor U12852 (N_12852,N_10575,N_9818);
nand U12853 (N_12853,N_11418,N_11116);
xor U12854 (N_12854,N_8983,N_10019);
and U12855 (N_12855,N_6255,N_11024);
or U12856 (N_12856,N_11067,N_10825);
nand U12857 (N_12857,N_7072,N_6128);
xor U12858 (N_12858,N_7188,N_8381);
nor U12859 (N_12859,N_10579,N_11583);
and U12860 (N_12860,N_7293,N_9874);
and U12861 (N_12861,N_10778,N_11713);
nor U12862 (N_12862,N_8510,N_11922);
nand U12863 (N_12863,N_8419,N_11076);
nor U12864 (N_12864,N_6309,N_11427);
nand U12865 (N_12865,N_11420,N_7758);
nand U12866 (N_12866,N_9077,N_8071);
nor U12867 (N_12867,N_9407,N_11794);
nand U12868 (N_12868,N_11601,N_11474);
or U12869 (N_12869,N_7493,N_8111);
or U12870 (N_12870,N_11956,N_7914);
or U12871 (N_12871,N_9126,N_8026);
nand U12872 (N_12872,N_6723,N_7904);
xnor U12873 (N_12873,N_7055,N_10582);
nor U12874 (N_12874,N_10868,N_9503);
nor U12875 (N_12875,N_7092,N_11472);
nand U12876 (N_12876,N_11406,N_7679);
and U12877 (N_12877,N_11149,N_10773);
nor U12878 (N_12878,N_6920,N_8755);
or U12879 (N_12879,N_7840,N_11129);
and U12880 (N_12880,N_10789,N_7317);
and U12881 (N_12881,N_11101,N_10218);
xnor U12882 (N_12882,N_8607,N_11008);
or U12883 (N_12883,N_7684,N_11473);
nor U12884 (N_12884,N_11265,N_6667);
nand U12885 (N_12885,N_9191,N_6386);
and U12886 (N_12886,N_10698,N_6571);
nor U12887 (N_12887,N_8671,N_7244);
or U12888 (N_12888,N_7646,N_8161);
or U12889 (N_12889,N_6918,N_9741);
and U12890 (N_12890,N_6959,N_8806);
nand U12891 (N_12891,N_8465,N_7101);
nand U12892 (N_12892,N_11434,N_9105);
and U12893 (N_12893,N_9589,N_10256);
xor U12894 (N_12894,N_10508,N_10919);
xnor U12895 (N_12895,N_6520,N_6094);
nor U12896 (N_12896,N_7832,N_7825);
or U12897 (N_12897,N_6719,N_9851);
xor U12898 (N_12898,N_7701,N_6855);
xor U12899 (N_12899,N_9867,N_10981);
and U12900 (N_12900,N_7171,N_10725);
xnor U12901 (N_12901,N_8264,N_6154);
nand U12902 (N_12902,N_7584,N_7432);
nand U12903 (N_12903,N_8163,N_7938);
nor U12904 (N_12904,N_6048,N_10375);
and U12905 (N_12905,N_6661,N_8144);
xor U12906 (N_12906,N_9618,N_6814);
and U12907 (N_12907,N_10876,N_9403);
and U12908 (N_12908,N_10081,N_10497);
xnor U12909 (N_12909,N_6032,N_8775);
nor U12910 (N_12910,N_10504,N_11372);
nand U12911 (N_12911,N_9973,N_9803);
xnor U12912 (N_12912,N_11542,N_7901);
xor U12913 (N_12913,N_11285,N_10730);
nor U12914 (N_12914,N_8077,N_7346);
or U12915 (N_12915,N_10628,N_9747);
xnor U12916 (N_12916,N_10443,N_10670);
or U12917 (N_12917,N_7402,N_8057);
xnor U12918 (N_12918,N_11679,N_10759);
xnor U12919 (N_12919,N_11210,N_9262);
nand U12920 (N_12920,N_9732,N_10809);
and U12921 (N_12921,N_8326,N_11606);
or U12922 (N_12922,N_11053,N_7353);
or U12923 (N_12923,N_7109,N_7860);
nor U12924 (N_12924,N_7898,N_10551);
nand U12925 (N_12925,N_6797,N_6342);
xor U12926 (N_12926,N_7336,N_9452);
or U12927 (N_12927,N_8514,N_8984);
nor U12928 (N_12928,N_7727,N_10473);
nand U12929 (N_12929,N_6970,N_11506);
xnor U12930 (N_12930,N_9665,N_10624);
nand U12931 (N_12931,N_9070,N_11485);
or U12932 (N_12932,N_11370,N_7668);
xor U12933 (N_12933,N_8720,N_8793);
nor U12934 (N_12934,N_7343,N_9405);
nor U12935 (N_12935,N_6244,N_7106);
or U12936 (N_12936,N_8139,N_9388);
or U12937 (N_12937,N_6846,N_11498);
nand U12938 (N_12938,N_10880,N_8579);
or U12939 (N_12939,N_10329,N_8578);
and U12940 (N_12940,N_8981,N_6467);
or U12941 (N_12941,N_6548,N_8865);
xnor U12942 (N_12942,N_6894,N_6353);
and U12943 (N_12943,N_10951,N_10129);
and U12944 (N_12944,N_9919,N_11422);
or U12945 (N_12945,N_11781,N_11484);
xor U12946 (N_12946,N_6922,N_11112);
nor U12947 (N_12947,N_7936,N_10205);
nor U12948 (N_12948,N_9340,N_8668);
or U12949 (N_12949,N_11571,N_9467);
or U12950 (N_12950,N_6685,N_11865);
nand U12951 (N_12951,N_11777,N_6803);
nand U12952 (N_12952,N_11376,N_10523);
nor U12953 (N_12953,N_9484,N_9892);
and U12954 (N_12954,N_7982,N_9739);
nand U12955 (N_12955,N_9043,N_9637);
nand U12956 (N_12956,N_10595,N_7513);
and U12957 (N_12957,N_9232,N_11015);
xor U12958 (N_12958,N_6625,N_10543);
and U12959 (N_12959,N_9690,N_11672);
and U12960 (N_12960,N_7482,N_6359);
xnor U12961 (N_12961,N_11938,N_6241);
or U12962 (N_12962,N_10419,N_10409);
and U12963 (N_12963,N_6397,N_7024);
and U12964 (N_12964,N_10864,N_9397);
xor U12965 (N_12965,N_9485,N_10923);
nor U12966 (N_12966,N_9517,N_11267);
and U12967 (N_12967,N_6134,N_9555);
or U12968 (N_12968,N_6027,N_8742);
nand U12969 (N_12969,N_6749,N_9656);
nor U12970 (N_12970,N_11531,N_7044);
nor U12971 (N_12971,N_6103,N_7836);
xnor U12972 (N_12972,N_10891,N_6381);
or U12973 (N_12973,N_9804,N_6457);
or U12974 (N_12974,N_9794,N_6695);
or U12975 (N_12975,N_10554,N_9835);
xor U12976 (N_12976,N_8810,N_11069);
nor U12977 (N_12977,N_9483,N_8776);
or U12978 (N_12978,N_7527,N_8241);
nand U12979 (N_12979,N_11974,N_9124);
or U12980 (N_12980,N_10086,N_9603);
nand U12981 (N_12981,N_10359,N_9640);
nor U12982 (N_12982,N_11916,N_7573);
and U12983 (N_12983,N_7665,N_7861);
nor U12984 (N_12984,N_9813,N_11541);
or U12985 (N_12985,N_7332,N_7077);
or U12986 (N_12986,N_8099,N_11557);
nor U12987 (N_12987,N_6113,N_9936);
and U12988 (N_12988,N_8027,N_10243);
nor U12989 (N_12989,N_9938,N_7617);
or U12990 (N_12990,N_11687,N_6299);
nor U12991 (N_12991,N_9059,N_8058);
nand U12992 (N_12992,N_11556,N_6065);
or U12993 (N_12993,N_9496,N_9298);
or U12994 (N_12994,N_10064,N_8140);
nor U12995 (N_12995,N_7530,N_6806);
or U12996 (N_12996,N_6562,N_6222);
and U12997 (N_12997,N_11367,N_10328);
xnor U12998 (N_12998,N_6597,N_8698);
nor U12999 (N_12999,N_8224,N_9734);
xnor U13000 (N_13000,N_7660,N_10573);
nand U13001 (N_13001,N_10822,N_10527);
or U13002 (N_13002,N_7663,N_9300);
xnor U13003 (N_13003,N_9799,N_7292);
xor U13004 (N_13004,N_10442,N_6173);
nor U13005 (N_13005,N_10685,N_10630);
and U13006 (N_13006,N_7476,N_7609);
xor U13007 (N_13007,N_11902,N_11176);
and U13008 (N_13008,N_11996,N_11399);
xnor U13009 (N_13009,N_9836,N_8184);
nand U13010 (N_13010,N_7435,N_9189);
nand U13011 (N_13011,N_11169,N_11749);
and U13012 (N_13012,N_6682,N_8833);
or U13013 (N_13013,N_6804,N_11648);
and U13014 (N_13014,N_7456,N_9140);
and U13015 (N_13015,N_11673,N_9700);
nand U13016 (N_13016,N_7948,N_10202);
and U13017 (N_13017,N_7429,N_11653);
nor U13018 (N_13018,N_11239,N_6648);
xor U13019 (N_13019,N_9896,N_11080);
xor U13020 (N_13020,N_8123,N_11537);
nor U13021 (N_13021,N_8540,N_7219);
or U13022 (N_13022,N_10215,N_10428);
or U13023 (N_13023,N_8017,N_9187);
xor U13024 (N_13024,N_7458,N_9525);
nand U13025 (N_13025,N_11534,N_11097);
nor U13026 (N_13026,N_7127,N_7177);
and U13027 (N_13027,N_9791,N_7156);
and U13028 (N_13028,N_11479,N_6473);
xor U13029 (N_13029,N_10896,N_6580);
xnor U13030 (N_13030,N_6152,N_7142);
nor U13031 (N_13031,N_6773,N_11680);
xnor U13032 (N_13032,N_8046,N_10067);
xor U13033 (N_13033,N_10065,N_6543);
nand U13034 (N_13034,N_6638,N_10057);
nand U13035 (N_13035,N_7415,N_6827);
or U13036 (N_13036,N_10466,N_11428);
nor U13037 (N_13037,N_6140,N_11019);
nand U13038 (N_13038,N_6466,N_8938);
or U13039 (N_13039,N_7976,N_10455);
xor U13040 (N_13040,N_9569,N_7865);
nand U13041 (N_13041,N_8843,N_7653);
xnor U13042 (N_13042,N_7138,N_8134);
nor U13043 (N_13043,N_7544,N_10281);
xnor U13044 (N_13044,N_7559,N_10944);
xnor U13045 (N_13045,N_6738,N_11913);
and U13046 (N_13046,N_10471,N_8529);
or U13047 (N_13047,N_8978,N_11394);
nor U13048 (N_13048,N_11738,N_11622);
or U13049 (N_13049,N_10945,N_11887);
nor U13050 (N_13050,N_11819,N_11401);
and U13051 (N_13051,N_10652,N_8666);
and U13052 (N_13052,N_10955,N_10415);
nor U13053 (N_13053,N_7307,N_7308);
or U13054 (N_13054,N_8669,N_11108);
and U13055 (N_13055,N_11718,N_6392);
nand U13056 (N_13056,N_9478,N_8019);
and U13057 (N_13057,N_7226,N_10877);
nand U13058 (N_13058,N_11788,N_6105);
nor U13059 (N_13059,N_11455,N_6874);
nor U13060 (N_13060,N_7963,N_8500);
nor U13061 (N_13061,N_11617,N_9118);
nand U13062 (N_13062,N_6419,N_6119);
xor U13063 (N_13063,N_9913,N_11855);
nor U13064 (N_13064,N_10322,N_9183);
nand U13065 (N_13065,N_11323,N_9148);
nand U13066 (N_13066,N_7862,N_9265);
and U13067 (N_13067,N_10669,N_6987);
xor U13068 (N_13068,N_11302,N_11923);
nand U13069 (N_13069,N_7547,N_7850);
nand U13070 (N_13070,N_6895,N_9236);
or U13071 (N_13071,N_10888,N_11760);
nor U13072 (N_13072,N_10635,N_7306);
and U13073 (N_13073,N_9590,N_10792);
and U13074 (N_13074,N_6099,N_8611);
and U13075 (N_13075,N_7946,N_9923);
and U13076 (N_13076,N_6884,N_9378);
or U13077 (N_13077,N_10586,N_8980);
or U13078 (N_13078,N_6767,N_6725);
nand U13079 (N_13079,N_7980,N_6221);
nor U13080 (N_13080,N_9502,N_9481);
nand U13081 (N_13081,N_6400,N_8513);
nor U13082 (N_13082,N_6421,N_9139);
nand U13083 (N_13083,N_11014,N_8603);
nand U13084 (N_13084,N_10385,N_7716);
xnor U13085 (N_13085,N_9044,N_9548);
nor U13086 (N_13086,N_8945,N_6774);
and U13087 (N_13087,N_10355,N_6182);
and U13088 (N_13088,N_11539,N_10646);
xor U13089 (N_13089,N_7431,N_7775);
nor U13090 (N_13090,N_11168,N_8506);
xor U13091 (N_13091,N_10190,N_9765);
nand U13092 (N_13092,N_11365,N_11824);
nand U13093 (N_13093,N_8493,N_10436);
and U13094 (N_13094,N_8760,N_10700);
and U13095 (N_13095,N_11725,N_6646);
nor U13096 (N_13096,N_9210,N_11002);
or U13097 (N_13097,N_8309,N_7610);
and U13098 (N_13098,N_6907,N_11597);
or U13099 (N_13099,N_6493,N_11940);
or U13100 (N_13100,N_7692,N_6446);
and U13101 (N_13101,N_9611,N_9989);
or U13102 (N_13102,N_10505,N_7220);
and U13103 (N_13103,N_11209,N_6618);
or U13104 (N_13104,N_9306,N_10781);
nor U13105 (N_13105,N_10472,N_11244);
and U13106 (N_13106,N_7921,N_10488);
nor U13107 (N_13107,N_8007,N_9115);
nor U13108 (N_13108,N_9788,N_10078);
and U13109 (N_13109,N_8034,N_6670);
or U13110 (N_13110,N_11204,N_9584);
and U13111 (N_13111,N_7680,N_7773);
nand U13112 (N_13112,N_8504,N_6972);
nand U13113 (N_13113,N_10418,N_7505);
or U13114 (N_13114,N_8360,N_9064);
nand U13115 (N_13115,N_7627,N_11959);
and U13116 (N_13116,N_8599,N_7249);
nor U13117 (N_13117,N_10643,N_7441);
or U13118 (N_13118,N_6356,N_10430);
or U13119 (N_13119,N_8397,N_8767);
xor U13120 (N_13120,N_6509,N_8640);
and U13121 (N_13121,N_9011,N_8696);
or U13122 (N_13122,N_8774,N_8485);
or U13123 (N_13123,N_6627,N_6212);
nand U13124 (N_13124,N_10591,N_10179);
and U13125 (N_13125,N_7545,N_8068);
nand U13126 (N_13126,N_10424,N_7702);
or U13127 (N_13127,N_7626,N_10649);
xor U13128 (N_13128,N_8142,N_9328);
xor U13129 (N_13129,N_8070,N_11711);
or U13130 (N_13130,N_7933,N_10765);
xor U13131 (N_13131,N_10603,N_11532);
or U13132 (N_13132,N_7047,N_11901);
and U13133 (N_13133,N_11490,N_6303);
or U13134 (N_13134,N_10900,N_7212);
xnor U13135 (N_13135,N_10878,N_8118);
nor U13136 (N_13136,N_6047,N_7131);
or U13137 (N_13137,N_7717,N_11880);
nand U13138 (N_13138,N_9107,N_9479);
nor U13139 (N_13139,N_10160,N_6308);
nor U13140 (N_13140,N_9578,N_9574);
nand U13141 (N_13141,N_7961,N_7436);
and U13142 (N_13142,N_9305,N_6501);
nand U13143 (N_13143,N_8362,N_6240);
or U13144 (N_13144,N_6912,N_8846);
xnor U13145 (N_13145,N_6458,N_9927);
and U13146 (N_13146,N_10333,N_11920);
xnor U13147 (N_13147,N_9868,N_6554);
and U13148 (N_13148,N_7724,N_8180);
xor U13149 (N_13149,N_11977,N_6280);
or U13150 (N_13150,N_7369,N_10741);
nand U13151 (N_13151,N_8758,N_10271);
and U13152 (N_13152,N_6267,N_6200);
or U13153 (N_13153,N_8757,N_10521);
nand U13154 (N_13154,N_10209,N_10834);
and U13155 (N_13155,N_7203,N_7947);
and U13156 (N_13156,N_10962,N_11732);
and U13157 (N_13157,N_7872,N_9145);
xnor U13158 (N_13158,N_10117,N_6209);
and U13159 (N_13159,N_6018,N_6974);
or U13160 (N_13160,N_7419,N_6617);
nor U13161 (N_13161,N_9272,N_10682);
and U13162 (N_13162,N_6281,N_8626);
or U13163 (N_13163,N_10079,N_10832);
or U13164 (N_13164,N_8384,N_9711);
or U13165 (N_13165,N_9814,N_7400);
or U13166 (N_13166,N_8188,N_8988);
xor U13167 (N_13167,N_11874,N_8690);
xor U13168 (N_13168,N_11197,N_11897);
or U13169 (N_13169,N_11671,N_9964);
or U13170 (N_13170,N_11105,N_8704);
and U13171 (N_13171,N_6017,N_7038);
nand U13172 (N_13172,N_7068,N_11603);
and U13173 (N_13173,N_6616,N_8770);
nor U13174 (N_13174,N_11863,N_10015);
nand U13175 (N_13175,N_11953,N_6266);
xnor U13176 (N_13176,N_10102,N_8277);
xnor U13177 (N_13177,N_6338,N_10098);
and U13178 (N_13178,N_7747,N_10609);
xor U13179 (N_13179,N_7186,N_11593);
xnor U13180 (N_13180,N_11029,N_11325);
nor U13181 (N_13181,N_7370,N_10413);
or U13182 (N_13182,N_6164,N_8565);
xor U13183 (N_13183,N_9114,N_8376);
or U13184 (N_13184,N_6258,N_6982);
nor U13185 (N_13185,N_11140,N_10151);
nor U13186 (N_13186,N_8723,N_9159);
nor U13187 (N_13187,N_6416,N_10458);
xor U13188 (N_13188,N_10826,N_9073);
and U13189 (N_13189,N_7869,N_6684);
nand U13190 (N_13190,N_10680,N_11780);
and U13191 (N_13191,N_9360,N_10662);
and U13192 (N_13192,N_11118,N_11413);
and U13193 (N_13193,N_10627,N_9894);
nand U13194 (N_13194,N_10530,N_9688);
xor U13195 (N_13195,N_8115,N_8059);
xnor U13196 (N_13196,N_8566,N_7935);
nor U13197 (N_13197,N_10203,N_11417);
or U13198 (N_13198,N_9099,N_6938);
and U13199 (N_13199,N_7945,N_9811);
xor U13200 (N_13200,N_6449,N_11841);
nor U13201 (N_13201,N_6076,N_7424);
nand U13202 (N_13202,N_6171,N_8434);
nor U13203 (N_13203,N_9893,N_8327);
or U13204 (N_13204,N_7145,N_10000);
nand U13205 (N_13205,N_7447,N_10683);
xor U13206 (N_13206,N_10082,N_6615);
or U13207 (N_13207,N_8731,N_7274);
nor U13208 (N_13208,N_7550,N_8966);
or U13209 (N_13209,N_6950,N_11300);
xor U13210 (N_13210,N_8849,N_11454);
xor U13211 (N_13211,N_9243,N_9514);
nand U13212 (N_13212,N_7967,N_7762);
or U13213 (N_13213,N_8868,N_11065);
and U13214 (N_13214,N_7251,N_11677);
or U13215 (N_13215,N_7858,N_7455);
and U13216 (N_13216,N_7708,N_11276);
nand U13217 (N_13217,N_6961,N_10119);
xnor U13218 (N_13218,N_11528,N_9440);
xor U13219 (N_13219,N_10671,N_7460);
or U13220 (N_13220,N_9400,N_11358);
and U13221 (N_13221,N_11397,N_11467);
and U13222 (N_13222,N_6390,N_10831);
nand U13223 (N_13223,N_7772,N_6511);
nand U13224 (N_13224,N_9510,N_6944);
xor U13225 (N_13225,N_11052,N_11179);
nor U13226 (N_13226,N_11705,N_6582);
nor U13227 (N_13227,N_8009,N_8973);
nand U13228 (N_13228,N_11227,N_9527);
or U13229 (N_13229,N_8836,N_10539);
and U13230 (N_13230,N_7054,N_11688);
nand U13231 (N_13231,N_6808,N_8209);
xnor U13232 (N_13232,N_11600,N_6830);
and U13233 (N_13233,N_7002,N_6073);
nand U13234 (N_13234,N_9601,N_10294);
and U13235 (N_13235,N_10593,N_11890);
nand U13236 (N_13236,N_6566,N_9750);
nor U13237 (N_13237,N_7123,N_10220);
xnor U13238 (N_13238,N_9163,N_6813);
nand U13239 (N_13239,N_8624,N_10470);
nand U13240 (N_13240,N_10902,N_10963);
xnor U13241 (N_13241,N_6858,N_8826);
xor U13242 (N_13242,N_9384,N_9916);
xnor U13243 (N_13243,N_6569,N_8652);
or U13244 (N_13244,N_7233,N_10087);
nand U13245 (N_13245,N_11507,N_10114);
xor U13246 (N_13246,N_7790,N_10960);
or U13247 (N_13247,N_10677,N_7854);
and U13248 (N_13248,N_7394,N_9972);
nand U13249 (N_13249,N_10286,N_10320);
nand U13250 (N_13250,N_9369,N_6775);
and U13251 (N_13251,N_11407,N_6933);
or U13252 (N_13252,N_11482,N_10094);
nand U13253 (N_13253,N_7227,N_9394);
nand U13254 (N_13254,N_11229,N_6316);
nor U13255 (N_13255,N_8882,N_9134);
or U13256 (N_13256,N_10724,N_10564);
nand U13257 (N_13257,N_7751,N_9707);
and U13258 (N_13258,N_10762,N_7275);
or U13259 (N_13259,N_8855,N_9231);
nand U13260 (N_13260,N_10705,N_6917);
and U13261 (N_13261,N_11566,N_8426);
nor U13262 (N_13262,N_11770,N_9294);
nand U13263 (N_13263,N_11588,N_9632);
or U13264 (N_13264,N_10836,N_6095);
or U13265 (N_13265,N_10206,N_11106);
nand U13266 (N_13266,N_8968,N_6175);
nand U13267 (N_13267,N_11081,N_9888);
and U13268 (N_13268,N_10283,N_6999);
or U13269 (N_13269,N_6310,N_9522);
nor U13270 (N_13270,N_9533,N_8928);
xnor U13271 (N_13271,N_7080,N_8396);
nor U13272 (N_13272,N_7362,N_7174);
nor U13273 (N_13273,N_7485,N_7968);
nor U13274 (N_13274,N_6605,N_6788);
xnor U13275 (N_13275,N_8400,N_9213);
xnor U13276 (N_13276,N_6908,N_6396);
and U13277 (N_13277,N_10924,N_10236);
xor U13278 (N_13278,N_9025,N_6930);
nand U13279 (N_13279,N_7863,N_11872);
xor U13280 (N_13280,N_10229,N_8985);
xnor U13281 (N_13281,N_7844,N_6998);
nand U13282 (N_13282,N_8332,N_8958);
xnor U13283 (N_13283,N_11460,N_8266);
and U13284 (N_13284,N_8152,N_10622);
xor U13285 (N_13285,N_6293,N_6237);
xnor U13286 (N_13286,N_11337,N_6382);
or U13287 (N_13287,N_8505,N_9817);
xnor U13288 (N_13288,N_8253,N_8338);
nand U13289 (N_13289,N_6371,N_11433);
nand U13290 (N_13290,N_6643,N_6236);
nor U13291 (N_13291,N_9143,N_7399);
nor U13292 (N_13292,N_11378,N_8117);
or U13293 (N_13293,N_10342,N_6125);
or U13294 (N_13294,N_11137,N_7450);
xor U13295 (N_13295,N_10577,N_9373);
and U13296 (N_13296,N_9410,N_11608);
and U13297 (N_13297,N_9040,N_10199);
xnor U13298 (N_13298,N_6653,N_11064);
and U13299 (N_13299,N_7474,N_8198);
and U13300 (N_13300,N_9349,N_7303);
and U13301 (N_13301,N_10568,N_10570);
xnor U13302 (N_13302,N_10580,N_8354);
nor U13303 (N_13303,N_11043,N_8325);
or U13304 (N_13304,N_7900,N_11377);
nor U13305 (N_13305,N_9857,N_10729);
and U13306 (N_13306,N_6668,N_7276);
and U13307 (N_13307,N_9858,N_9024);
nand U13308 (N_13308,N_9375,N_7302);
xor U13309 (N_13309,N_8313,N_11559);
xnor U13310 (N_13310,N_10421,N_9475);
xor U13311 (N_13311,N_7199,N_11620);
xor U13312 (N_13312,N_11963,N_9423);
or U13313 (N_13313,N_8715,N_8625);
nor U13314 (N_13314,N_10360,N_10874);
nand U13315 (N_13315,N_7805,N_6011);
and U13316 (N_13316,N_6800,N_6688);
and U13317 (N_13317,N_9399,N_6968);
and U13318 (N_13318,N_10255,N_7330);
xor U13319 (N_13319,N_11805,N_8257);
xor U13320 (N_13320,N_11605,N_9430);
or U13321 (N_13321,N_10757,N_7795);
or U13322 (N_13322,N_7500,N_6272);
xnor U13323 (N_13323,N_10096,N_8631);
or U13324 (N_13324,N_8554,N_7696);
xor U13325 (N_13325,N_9904,N_6678);
nand U13326 (N_13326,N_11930,N_6877);
xnor U13327 (N_13327,N_10710,N_11217);
nor U13328 (N_13328,N_10588,N_10688);
nand U13329 (N_13329,N_11158,N_9225);
nor U13330 (N_13330,N_7135,N_9350);
nor U13331 (N_13331,N_11720,N_7289);
or U13332 (N_13332,N_6921,N_11233);
or U13333 (N_13333,N_10235,N_8126);
xor U13334 (N_13334,N_10727,N_8154);
nor U13335 (N_13335,N_7787,N_6437);
and U13336 (N_13336,N_6111,N_9982);
nand U13337 (N_13337,N_11612,N_11845);
or U13338 (N_13338,N_7607,N_9875);
xor U13339 (N_13339,N_10377,N_8691);
or U13340 (N_13340,N_10922,N_10594);
xor U13341 (N_13341,N_8687,N_8629);
or U13342 (N_13342,N_11329,N_6587);
xor U13343 (N_13343,N_6158,N_9233);
or U13344 (N_13344,N_8881,N_9418);
nor U13345 (N_13345,N_6226,N_8944);
nand U13346 (N_13346,N_11650,N_9641);
and U13347 (N_13347,N_10973,N_9311);
and U13348 (N_13348,N_9646,N_11202);
or U13349 (N_13349,N_7328,N_9336);
nand U13350 (N_13350,N_6036,N_8832);
xnor U13351 (N_13351,N_6517,N_10917);
xor U13352 (N_13352,N_7533,N_6023);
xnor U13353 (N_13353,N_8388,N_9470);
xor U13354 (N_13354,N_9877,N_6958);
nor U13355 (N_13355,N_10772,N_6355);
nor U13356 (N_13356,N_9737,N_7151);
nand U13357 (N_13357,N_8272,N_6410);
nand U13358 (N_13358,N_8778,N_7759);
nor U13359 (N_13359,N_9551,N_7405);
or U13360 (N_13360,N_7788,N_11003);
and U13361 (N_13361,N_10787,N_9912);
nor U13362 (N_13362,N_10107,N_9188);
nand U13363 (N_13363,N_8562,N_8431);
and U13364 (N_13364,N_10860,N_6216);
xnor U13365 (N_13365,N_10147,N_9844);
or U13366 (N_13366,N_6576,N_9660);
or U13367 (N_13367,N_8340,N_11196);
nand U13368 (N_13368,N_10183,N_8358);
xnor U13369 (N_13369,N_11451,N_9062);
or U13370 (N_13370,N_7423,N_9374);
and U13371 (N_13371,N_6469,N_11423);
or U13372 (N_13372,N_8283,N_9766);
and U13373 (N_13373,N_11240,N_6407);
nor U13374 (N_13374,N_7187,N_11148);
xor U13375 (N_13375,N_7304,N_8069);
xor U13376 (N_13376,N_10578,N_7440);
nand U13377 (N_13377,N_10851,N_11133);
xnor U13378 (N_13378,N_7022,N_6092);
and U13379 (N_13379,N_7083,N_8536);
and U13380 (N_13380,N_11268,N_7503);
nand U13381 (N_13381,N_9607,N_7634);
and U13382 (N_13382,N_10437,N_6423);
nand U13383 (N_13383,N_10756,N_7238);
or U13384 (N_13384,N_6835,N_11430);
or U13385 (N_13385,N_8116,N_9345);
or U13386 (N_13386,N_10726,N_9172);
xnor U13387 (N_13387,N_7769,N_8227);
or U13388 (N_13388,N_11241,N_9131);
xor U13389 (N_13389,N_11110,N_10728);
nor U13390 (N_13390,N_8063,N_6832);
nor U13391 (N_13391,N_8563,N_6577);
nand U13392 (N_13392,N_7291,N_6083);
nor U13393 (N_13393,N_6610,N_10378);
and U13394 (N_13394,N_9974,N_10587);
nor U13395 (N_13395,N_7620,N_8293);
nand U13396 (N_13396,N_10435,N_8486);
xor U13397 (N_13397,N_8659,N_7749);
nor U13398 (N_13398,N_8201,N_11131);
or U13399 (N_13399,N_7285,N_9576);
xnor U13400 (N_13400,N_10420,N_9764);
nand U13401 (N_13401,N_11290,N_8925);
and U13402 (N_13402,N_10276,N_7601);
xnor U13403 (N_13403,N_8001,N_7821);
xnor U13404 (N_13404,N_7868,N_7345);
xor U13405 (N_13405,N_7418,N_7993);
xor U13406 (N_13406,N_11504,N_6843);
nand U13407 (N_13407,N_6838,N_10134);
and U13408 (N_13408,N_7159,N_11746);
nand U13409 (N_13409,N_9625,N_9396);
nand U13410 (N_13410,N_6770,N_9971);
nor U13411 (N_13411,N_8642,N_11219);
and U13412 (N_13412,N_6405,N_11615);
nor U13413 (N_13413,N_9958,N_7154);
nor U13414 (N_13414,N_6716,N_10246);
nand U13415 (N_13415,N_10561,N_8879);
nand U13416 (N_13416,N_6860,N_9985);
nor U13417 (N_13417,N_6742,N_9208);
and U13418 (N_13418,N_10148,N_11818);
xnor U13419 (N_13419,N_6731,N_8541);
and U13420 (N_13420,N_8052,N_8322);
xnor U13421 (N_13421,N_6666,N_9657);
nand U13422 (N_13422,N_9117,N_9082);
nand U13423 (N_13423,N_9721,N_6510);
xor U13424 (N_13424,N_8474,N_8160);
or U13425 (N_13425,N_8785,N_6246);
xnor U13426 (N_13426,N_10966,N_9157);
nor U13427 (N_13427,N_11178,N_7587);
or U13428 (N_13428,N_9506,N_11592);
nand U13429 (N_13429,N_9944,N_9006);
nand U13430 (N_13430,N_6482,N_10659);
nor U13431 (N_13431,N_10367,N_8406);
nor U13432 (N_13432,N_11272,N_7999);
xor U13433 (N_13433,N_8728,N_7613);
nor U13434 (N_13434,N_9501,N_11635);
nand U13435 (N_13435,N_8676,N_10063);
and U13436 (N_13436,N_9577,N_9166);
xnor U13437 (N_13437,N_10943,N_6489);
xor U13438 (N_13438,N_6129,N_11254);
xor U13439 (N_13439,N_9079,N_9786);
or U13440 (N_13440,N_9102,N_7662);
nor U13441 (N_13441,N_6259,N_11038);
and U13442 (N_13442,N_10062,N_9365);
xnor U13443 (N_13443,N_11452,N_10072);
and U13444 (N_13444,N_11561,N_6232);
nor U13445 (N_13445,N_9515,N_10085);
or U13446 (N_13446,N_7767,N_8066);
nor U13447 (N_13447,N_7120,N_10306);
and U13448 (N_13448,N_6347,N_10009);
or U13449 (N_13449,N_11449,N_9793);
or U13450 (N_13450,N_7647,N_7058);
xnor U13451 (N_13451,N_9194,N_8936);
or U13452 (N_13452,N_9330,N_8932);
xnor U13453 (N_13453,N_6679,N_10940);
and U13454 (N_13454,N_7954,N_10076);
xnor U13455 (N_13455,N_8498,N_11586);
and U13456 (N_13456,N_7827,N_9280);
or U13457 (N_13457,N_6491,N_9594);
nand U13458 (N_13458,N_8252,N_8538);
nand U13459 (N_13459,N_9445,N_11926);
xor U13460 (N_13460,N_10388,N_11667);
nor U13461 (N_13461,N_11787,N_6481);
xor U13462 (N_13462,N_8459,N_7281);
xor U13463 (N_13463,N_10314,N_8330);
xor U13464 (N_13464,N_6931,N_9645);
nand U13465 (N_13465,N_11311,N_11328);
nand U13466 (N_13466,N_8299,N_7490);
nand U13467 (N_13467,N_9192,N_8749);
nor U13468 (N_13468,N_7427,N_10406);
nand U13469 (N_13469,N_10980,N_7743);
and U13470 (N_13470,N_6540,N_8886);
nor U13471 (N_13471,N_6692,N_11250);
xor U13472 (N_13472,N_9719,N_10623);
or U13473 (N_13473,N_7315,N_11402);
or U13474 (N_13474,N_9581,N_6739);
or U13475 (N_13475,N_6138,N_10784);
and U13476 (N_13476,N_10244,N_6374);
and U13477 (N_13477,N_10224,N_7150);
or U13478 (N_13478,N_8039,N_6443);
nand U13479 (N_13479,N_11320,N_10103);
nor U13480 (N_13480,N_10634,N_10706);
xnor U13481 (N_13481,N_11139,N_6823);
nand U13482 (N_13482,N_7603,N_6077);
xor U13483 (N_13483,N_10820,N_7125);
and U13484 (N_13484,N_6028,N_7383);
nand U13485 (N_13485,N_8242,N_10863);
and U13486 (N_13486,N_10804,N_10207);
xnor U13487 (N_13487,N_6357,N_11616);
and U13488 (N_13488,N_7026,N_11545);
and U13489 (N_13489,N_11011,N_10289);
nand U13490 (N_13490,N_9174,N_6864);
and U13491 (N_13491,N_11844,N_7180);
or U13492 (N_13492,N_8515,N_10656);
nor U13493 (N_13493,N_8369,N_10090);
and U13494 (N_13494,N_11275,N_8544);
and U13495 (N_13495,N_10817,N_7023);
nor U13496 (N_13496,N_9086,N_7331);
nand U13497 (N_13497,N_11692,N_9532);
and U13498 (N_13498,N_11979,N_7656);
nand U13499 (N_13499,N_6234,N_7768);
nor U13500 (N_13500,N_9307,N_11927);
and U13501 (N_13501,N_8100,N_7576);
xnor U13502 (N_13502,N_9815,N_8345);
nor U13503 (N_13503,N_8392,N_11546);
nand U13504 (N_13504,N_8225,N_9529);
and U13505 (N_13505,N_6284,N_8374);
nor U13506 (N_13506,N_6319,N_10916);
nand U13507 (N_13507,N_11501,N_9620);
nor U13508 (N_13508,N_11703,N_8460);
xor U13509 (N_13509,N_9828,N_11750);
and U13510 (N_13510,N_6836,N_7687);
xnor U13511 (N_13511,N_7262,N_7981);
xnor U13512 (N_13512,N_9477,N_11900);
and U13513 (N_13513,N_6058,N_6828);
nor U13514 (N_13514,N_7839,N_9907);
nor U13515 (N_13515,N_7375,N_8021);
nand U13516 (N_13516,N_9037,N_6254);
xnor U13517 (N_13517,N_11034,N_7214);
or U13518 (N_13518,N_10376,N_11223);
nand U13519 (N_13519,N_7501,N_6418);
and U13520 (N_13520,N_7263,N_9190);
nand U13521 (N_13521,N_10748,N_11299);
xor U13522 (N_13522,N_7273,N_6365);
or U13523 (N_13523,N_8093,N_11689);
or U13524 (N_13524,N_10858,N_8885);
and U13525 (N_13525,N_8912,N_8738);
nand U13526 (N_13526,N_10222,N_9897);
xor U13527 (N_13527,N_11296,N_7492);
nor U13528 (N_13528,N_10673,N_10128);
xor U13529 (N_13529,N_6393,N_11933);
or U13530 (N_13530,N_10233,N_10813);
or U13531 (N_13531,N_11364,N_7414);
xor U13532 (N_13532,N_11925,N_7899);
nand U13533 (N_13533,N_8516,N_6573);
xor U13534 (N_13534,N_8667,N_11104);
xor U13535 (N_13535,N_10324,N_11822);
and U13536 (N_13536,N_10350,N_7633);
or U13537 (N_13537,N_10365,N_7230);
or U13538 (N_13538,N_7923,N_6596);
nor U13539 (N_13539,N_8020,N_10404);
nand U13540 (N_13540,N_11294,N_6849);
xnor U13541 (N_13541,N_6910,N_6139);
nor U13542 (N_13542,N_8158,N_11722);
xnor U13543 (N_13543,N_9626,N_9608);
xnor U13544 (N_13544,N_8747,N_10665);
nor U13545 (N_13545,N_10189,N_9408);
xor U13546 (N_13546,N_6953,N_11584);
xor U13547 (N_13547,N_8641,N_7912);
and U13548 (N_13548,N_6651,N_7810);
xnor U13549 (N_13549,N_7703,N_6101);
or U13550 (N_13550,N_8900,N_11258);
nand U13551 (N_13551,N_8710,N_7888);
xnor U13552 (N_13552,N_7009,N_11194);
xor U13553 (N_13553,N_11808,N_9450);
and U13554 (N_13554,N_6082,N_6452);
xor U13555 (N_13555,N_9355,N_9299);
or U13556 (N_13556,N_8808,N_7979);
or U13557 (N_13557,N_7413,N_8650);
and U13558 (N_13558,N_10566,N_8852);
xnor U13559 (N_13559,N_6030,N_10542);
nand U13560 (N_13560,N_7321,N_8141);
nand U13561 (N_13561,N_8960,N_10987);
nand U13562 (N_13562,N_10198,N_7569);
nor U13563 (N_13563,N_11702,N_8276);
or U13564 (N_13564,N_10519,N_7523);
nor U13565 (N_13565,N_6594,N_10165);
or U13566 (N_13566,N_10620,N_10201);
xnor U13567 (N_13567,N_9722,N_9181);
or U13568 (N_13568,N_6075,N_6621);
nand U13569 (N_13569,N_8421,N_8468);
nor U13570 (N_13570,N_6033,N_9429);
nand U13571 (N_13571,N_8594,N_11693);
nor U13572 (N_13572,N_10529,N_7806);
xnor U13573 (N_13573,N_11724,N_8217);
or U13574 (N_13574,N_10675,N_8221);
nor U13575 (N_13575,N_8677,N_11816);
xnor U13576 (N_13576,N_6256,N_9002);
nor U13577 (N_13577,N_10790,N_8053);
and U13578 (N_13578,N_8709,N_11426);
nand U13579 (N_13579,N_7225,N_10621);
xnor U13580 (N_13580,N_7011,N_11776);
nand U13581 (N_13581,N_10870,N_9884);
nor U13582 (N_13582,N_9271,N_6513);
or U13583 (N_13583,N_7555,N_11893);
and U13584 (N_13584,N_8232,N_7254);
nand U13585 (N_13585,N_11270,N_11550);
nand U13586 (N_13586,N_6869,N_11381);
and U13587 (N_13587,N_8872,N_7041);
nor U13588 (N_13588,N_9069,N_9693);
xnor U13589 (N_13589,N_11266,N_6876);
or U13590 (N_13590,N_10272,N_6965);
nand U13591 (N_13591,N_6455,N_7232);
or U13592 (N_13592,N_9170,N_6591);
or U13593 (N_13593,N_7489,N_10935);
nand U13594 (N_13594,N_8550,N_8273);
and U13595 (N_13595,N_8292,N_11046);
nand U13596 (N_13596,N_11867,N_8888);
nor U13597 (N_13597,N_7886,N_8646);
nand U13598 (N_13598,N_8926,N_8399);
and U13599 (N_13599,N_10292,N_10775);
nand U13600 (N_13600,N_8441,N_6691);
nor U13601 (N_13601,N_10493,N_10232);
xnor U13602 (N_13602,N_8771,N_11526);
nand U13603 (N_13603,N_10239,N_7563);
and U13604 (N_13604,N_9493,N_11762);
xor U13605 (N_13605,N_11710,N_10049);
or U13606 (N_13606,N_6551,N_10054);
or U13607 (N_13607,N_7139,N_6451);
and U13608 (N_13608,N_11551,N_6929);
nand U13609 (N_13609,N_9983,N_6051);
nor U13610 (N_13610,N_8526,N_9751);
or U13611 (N_13611,N_7457,N_7020);
xnor U13612 (N_13612,N_11647,N_6519);
nand U13613 (N_13613,N_7670,N_6471);
and U13614 (N_13614,N_10991,N_8113);
nand U13615 (N_13615,N_10703,N_11280);
and U13616 (N_13616,N_6224,N_11657);
and U13617 (N_13617,N_9627,N_9110);
and U13618 (N_13618,N_7367,N_7728);
and U13619 (N_13619,N_6409,N_8108);
nand U13620 (N_13620,N_6533,N_8782);
or U13621 (N_13621,N_8467,N_7278);
xnor U13622 (N_13622,N_9000,N_6340);
xnor U13623 (N_13623,N_11012,N_9004);
xor U13624 (N_13624,N_10045,N_6861);
nand U13625 (N_13625,N_7965,N_6964);
xnor U13626 (N_13626,N_8890,N_7645);
or U13627 (N_13627,N_9259,N_6821);
and U13628 (N_13628,N_11934,N_6078);
and U13629 (N_13629,N_9419,N_9536);
xor U13630 (N_13630,N_10310,N_6290);
and U13631 (N_13631,N_7629,N_7341);
nand U13632 (N_13632,N_8443,N_9144);
and U13633 (N_13633,N_6508,N_8124);
nor U13634 (N_13634,N_8812,N_8135);
nand U13635 (N_13635,N_11135,N_7753);
or U13636 (N_13636,N_6496,N_6364);
or U13637 (N_13637,N_8996,N_11915);
or U13638 (N_13638,N_10964,N_6346);
xnor U13639 (N_13639,N_6007,N_9898);
nor U13640 (N_13640,N_8994,N_6847);
xnor U13641 (N_13641,N_9988,N_8357);
or U13642 (N_13642,N_8274,N_6350);
nand U13643 (N_13643,N_10055,N_9872);
nand U13644 (N_13644,N_10011,N_9619);
nand U13645 (N_13645,N_10638,N_6275);
and U13646 (N_13646,N_10182,N_8032);
nand U13647 (N_13647,N_11087,N_11517);
and U13648 (N_13648,N_7407,N_9852);
or U13649 (N_13649,N_6372,N_8692);
nand U13650 (N_13650,N_11348,N_11074);
and U13651 (N_13651,N_8784,N_6126);
nand U13652 (N_13652,N_11905,N_10033);
nor U13653 (N_13653,N_10956,N_11860);
nand U13654 (N_13654,N_7064,N_11346);
xnor U13655 (N_13655,N_9769,N_6039);
nand U13656 (N_13656,N_8197,N_8587);
nand U13657 (N_13657,N_11248,N_10003);
nand U13658 (N_13658,N_10260,N_11716);
nand U13659 (N_13659,N_11277,N_9249);
xor U13660 (N_13660,N_9379,N_11569);
nand U13661 (N_13661,N_8939,N_10131);
xnor U13662 (N_13662,N_11646,N_7095);
and U13663 (N_13663,N_8351,N_9570);
or U13664 (N_13664,N_9679,N_9165);
or U13665 (N_13665,N_11424,N_8524);
nand U13666 (N_13666,N_8683,N_7885);
xnor U13667 (N_13667,N_9469,N_8088);
nand U13668 (N_13668,N_8122,N_6463);
nand U13669 (N_13669,N_8827,N_7288);
and U13670 (N_13670,N_6247,N_7412);
or U13671 (N_13671,N_11664,N_7625);
and U13672 (N_13672,N_8567,N_8373);
nor U13673 (N_13673,N_6376,N_7166);
xor U13674 (N_13674,N_8736,N_8296);
xnor U13675 (N_13675,N_10023,N_6118);
and U13676 (N_13676,N_6906,N_6395);
or U13677 (N_13677,N_7012,N_11573);
nand U13678 (N_13678,N_7305,N_7144);
or U13679 (N_13679,N_9184,N_9047);
and U13680 (N_13680,N_7511,N_10625);
and U13681 (N_13681,N_9296,N_6328);
xor U13682 (N_13682,N_10216,N_8060);
or U13683 (N_13683,N_11189,N_7744);
nor U13684 (N_13684,N_6195,N_9969);
or U13685 (N_13685,N_11049,N_9993);
nand U13686 (N_13686,N_9290,N_9882);
and U13687 (N_13687,N_6608,N_7908);
nand U13688 (N_13688,N_6871,N_8657);
xnor U13689 (N_13689,N_6201,N_6301);
and U13690 (N_13690,N_7467,N_6652);
nor U13691 (N_13691,N_7422,N_11324);
xor U13692 (N_13692,N_9138,N_6264);
nand U13693 (N_13693,N_10929,N_6091);
xor U13694 (N_13694,N_8364,N_8555);
xnor U13695 (N_13695,N_10932,N_10092);
xnor U13696 (N_13696,N_11457,N_11637);
or U13697 (N_13697,N_7894,N_8136);
or U13698 (N_13698,N_7830,N_6708);
nor U13699 (N_13699,N_11023,N_10059);
nor U13700 (N_13700,N_8525,N_6147);
nor U13701 (N_13701,N_6535,N_9239);
nor U13702 (N_13702,N_9459,N_8528);
nand U13703 (N_13703,N_8743,N_11251);
nor U13704 (N_13704,N_8818,N_9358);
nand U13705 (N_13705,N_7735,N_11871);
nor U13706 (N_13706,N_11308,N_11694);
xnor U13707 (N_13707,N_6223,N_6867);
xnor U13708 (N_13708,N_11031,N_8453);
and U13709 (N_13709,N_6645,N_9976);
nand U13710 (N_13710,N_9849,N_9929);
and U13711 (N_13711,N_9486,N_7103);
nor U13712 (N_13712,N_8681,N_11151);
and U13713 (N_13713,N_11811,N_7837);
and U13714 (N_13714,N_6599,N_11846);
nor U13715 (N_13715,N_9720,N_9051);
xnor U13716 (N_13716,N_11500,N_6348);
nor U13717 (N_13717,N_7667,N_11441);
xor U13718 (N_13718,N_7915,N_11155);
nand U13719 (N_13719,N_7469,N_10510);
nand U13720 (N_13720,N_11585,N_11013);
nand U13721 (N_13721,N_6526,N_6940);
nor U13722 (N_13722,N_8386,N_11574);
nand U13723 (N_13723,N_11278,N_9850);
xnor U13724 (N_13724,N_8816,N_10002);
nand U13725 (N_13725,N_9371,N_9644);
or U13726 (N_13726,N_8920,N_9975);
nor U13727 (N_13727,N_6180,N_10780);
xnor U13728 (N_13728,N_11868,N_10811);
nor U13729 (N_13729,N_6538,N_7789);
and U13730 (N_13730,N_7245,N_6188);
xor U13731 (N_13731,N_8114,N_10550);
xor U13732 (N_13732,N_11771,N_8271);
nand U13733 (N_13733,N_11939,N_9103);
xnor U13734 (N_13734,N_7333,N_11704);
and U13735 (N_13735,N_7121,N_10195);
and U13736 (N_13736,N_7161,N_8680);
nor U13737 (N_13737,N_11825,N_7229);
and U13738 (N_13738,N_7529,N_8859);
nor U13739 (N_13739,N_7005,N_11136);
nand U13740 (N_13740,N_11117,N_9948);
and U13741 (N_13741,N_6845,N_10618);
nand U13742 (N_13742,N_10839,N_7449);
or U13743 (N_13743,N_9489,N_7287);
nand U13744 (N_13744,N_9810,N_10788);
and U13745 (N_13745,N_10953,N_9664);
or U13746 (N_13746,N_8956,N_11344);
nor U13747 (N_13747,N_9260,N_6839);
nor U13748 (N_13748,N_8261,N_6016);
xor U13749 (N_13749,N_7223,N_9910);
xnor U13750 (N_13750,N_10732,N_6426);
or U13751 (N_13751,N_8167,N_8164);
nor U13752 (N_13752,N_9617,N_10660);
xnor U13753 (N_13753,N_11613,N_7479);
xnor U13754 (N_13754,N_9453,N_9749);
or U13755 (N_13755,N_6450,N_6932);
nand U13756 (N_13756,N_11514,N_7356);
nor U13757 (N_13757,N_10498,N_6840);
xnor U13758 (N_13758,N_11249,N_10217);
nand U13759 (N_13759,N_11847,N_8147);
or U13760 (N_13760,N_10116,N_10861);
nand U13761 (N_13761,N_10541,N_7499);
nand U13762 (N_13762,N_11618,N_11446);
and U13763 (N_13763,N_8236,N_9615);
or U13764 (N_13764,N_8685,N_10381);
xor U13765 (N_13765,N_9740,N_9169);
nor U13766 (N_13766,N_7590,N_10075);
nand U13767 (N_13767,N_11726,N_8189);
and U13768 (N_13768,N_11480,N_9286);
xor U13769 (N_13769,N_10712,N_11494);
xor U13770 (N_13770,N_6202,N_9613);
or U13771 (N_13771,N_6186,N_8701);
nor U13772 (N_13772,N_8481,N_6986);
and U13773 (N_13773,N_8307,N_7018);
or U13774 (N_13774,N_9671,N_10689);
xnor U13775 (N_13775,N_9984,N_6879);
and U13776 (N_13776,N_8084,N_8424);
and U13777 (N_13777,N_11669,N_9926);
and U13778 (N_13778,N_9879,N_8370);
nor U13779 (N_13779,N_8269,N_9833);
xnor U13780 (N_13780,N_11643,N_8964);
and U13781 (N_13781,N_8133,N_9648);
nand U13782 (N_13782,N_8575,N_6837);
xnor U13783 (N_13783,N_10701,N_11877);
xor U13784 (N_13784,N_9773,N_9742);
and U13785 (N_13785,N_6544,N_7162);
or U13786 (N_13786,N_11797,N_9994);
nand U13787 (N_13787,N_11730,N_9490);
or U13788 (N_13788,N_8802,N_7950);
xnor U13789 (N_13789,N_10774,N_11878);
nand U13790 (N_13790,N_7824,N_11382);
nand U13791 (N_13791,N_10482,N_7070);
nand U13792 (N_13792,N_8722,N_8501);
or U13793 (N_13793,N_6514,N_10469);
and U13794 (N_13794,N_7926,N_9425);
or U13795 (N_13795,N_9716,N_9319);
nor U13796 (N_13796,N_11757,N_8911);
and U13797 (N_13797,N_9526,N_11971);
and U13798 (N_13798,N_9902,N_11958);
nor U13799 (N_13799,N_10163,N_11955);
and U13800 (N_13800,N_6021,N_7190);
xnor U13801 (N_13801,N_11994,N_6969);
nor U13802 (N_13802,N_10507,N_6776);
nand U13803 (N_13803,N_10307,N_11954);
or U13804 (N_13804,N_8331,N_8581);
xnor U13805 (N_13805,N_8329,N_6460);
nor U13806 (N_13806,N_11668,N_9173);
nand U13807 (N_13807,N_8584,N_11326);
xnor U13808 (N_13808,N_7110,N_6327);
and U13809 (N_13809,N_10423,N_11091);
nor U13810 (N_13810,N_10694,N_6951);
and U13811 (N_13811,N_8548,N_8746);
and U13812 (N_13812,N_7736,N_10875);
xnor U13813 (N_13813,N_9616,N_11283);
or U13814 (N_13814,N_9084,N_9754);
nand U13815 (N_13815,N_8574,N_9544);
xnor U13816 (N_13816,N_10312,N_10786);
xnor U13817 (N_13817,N_9558,N_11975);
xnor U13818 (N_13818,N_10050,N_8237);
nor U13819 (N_13819,N_11409,N_8185);
and U13820 (N_13820,N_9763,N_11904);
and U13821 (N_13821,N_8155,N_10108);
nor U13822 (N_13822,N_10770,N_7974);
nor U13823 (N_13823,N_9748,N_6598);
and U13824 (N_13824,N_7741,N_10321);
nor U13825 (N_13825,N_11063,N_10484);
nand U13826 (N_13826,N_6411,N_8847);
nand U13827 (N_13827,N_7057,N_10882);
nand U13828 (N_13828,N_11885,N_6160);
or U13829 (N_13829,N_11491,N_8390);
and U13830 (N_13830,N_8634,N_11443);
and U13831 (N_13831,N_8067,N_9519);
nor U13832 (N_13832,N_6369,N_7215);
nor U13833 (N_13833,N_7785,N_7691);
nand U13834 (N_13834,N_8711,N_7364);
and U13835 (N_13835,N_6824,N_7801);
nand U13836 (N_13836,N_9856,N_9101);
xor U13837 (N_13837,N_7594,N_8753);
nand U13838 (N_13838,N_9152,N_7052);
xnor U13839 (N_13839,N_10637,N_6387);
or U13840 (N_13840,N_11644,N_11804);
or U13841 (N_13841,N_11102,N_8109);
or U13842 (N_13842,N_6005,N_6518);
or U13843 (N_13843,N_11580,N_11701);
and U13844 (N_13844,N_8931,N_9010);
and U13845 (N_13845,N_10970,N_8547);
xnor U13846 (N_13846,N_8213,N_6955);
xor U13847 (N_13847,N_9609,N_7028);
and U13848 (N_13848,N_9643,N_11621);
xnor U13849 (N_13849,N_6282,N_9706);
and U13850 (N_13850,N_9261,N_10856);
nor U13851 (N_13851,N_9571,N_7279);
and U13852 (N_13852,N_8312,N_9258);
nor U13853 (N_13853,N_7566,N_10827);
or U13854 (N_13854,N_9372,N_10185);
nor U13855 (N_13855,N_11918,N_8450);
or U13856 (N_13856,N_10390,N_11315);
and U13857 (N_13857,N_9111,N_8456);
nand U13858 (N_13858,N_10293,N_9153);
or U13859 (N_13859,N_7514,N_8395);
and U13860 (N_13860,N_8825,N_8359);
and U13861 (N_13861,N_9113,N_7874);
nor U13862 (N_13862,N_9367,N_8535);
nor U13863 (N_13863,N_10426,N_10696);
nand U13864 (N_13864,N_10118,N_7520);
xnor U13865 (N_13865,N_7742,N_9287);
xnor U13866 (N_13866,N_7949,N_7522);
xnor U13867 (N_13867,N_10170,N_8787);
or U13868 (N_13868,N_6053,N_10949);
nor U13869 (N_13869,N_10137,N_6339);
nand U13870 (N_13870,N_6358,N_10242);
xnor U13871 (N_13871,N_9614,N_7815);
xor U13872 (N_13872,N_8853,N_8941);
and U13873 (N_13873,N_9960,N_10879);
xor U13874 (N_13874,N_10608,N_7847);
xor U13875 (N_13875,N_10425,N_8788);
or U13876 (N_13876,N_11558,N_11889);
or U13877 (N_13877,N_10843,N_6658);
nand U13878 (N_13878,N_6890,N_7257);
or U13879 (N_13879,N_10806,N_9499);
and U13880 (N_13880,N_7348,N_10132);
nand U13881 (N_13881,N_10800,N_6330);
nand U13882 (N_13882,N_10977,N_8451);
nand U13883 (N_13883,N_7035,N_6729);
nand U13884 (N_13884,N_9432,N_8592);
nand U13885 (N_13885,N_6574,N_8492);
and U13886 (N_13886,N_7351,N_6478);
and U13887 (N_13887,N_11989,N_10269);
nor U13888 (N_13888,N_10046,N_11981);
and U13889 (N_13889,N_10978,N_7725);
xnor U13890 (N_13890,N_11156,N_11948);
nor U13891 (N_13891,N_8416,N_7093);
nor U13892 (N_13892,N_6089,N_9250);
xnor U13893 (N_13893,N_10930,N_6637);
nor U13894 (N_13894,N_11147,N_11623);
or U13895 (N_13895,N_8233,N_8083);
nand U13896 (N_13896,N_8128,N_9635);
xor U13897 (N_13897,N_7265,N_9251);
xor U13898 (N_13898,N_8297,N_9663);
nor U13899 (N_13899,N_11463,N_6525);
and U13900 (N_13900,N_8754,N_7608);
nand U13901 (N_13901,N_6412,N_9537);
nor U13902 (N_13902,N_7486,N_11761);
and U13903 (N_13903,N_6289,N_8512);
nand U13904 (N_13904,N_6135,N_11731);
xnor U13905 (N_13905,N_11626,N_7943);
or U13906 (N_13906,N_7818,N_6131);
nor U13907 (N_13907,N_6752,N_7842);
nand U13908 (N_13908,N_11906,N_11395);
nand U13909 (N_13909,N_9156,N_9630);
nor U13910 (N_13910,N_8120,N_6145);
or U13911 (N_13911,N_9672,N_8779);
or U13912 (N_13912,N_10304,N_10340);
nor U13913 (N_13913,N_8132,N_6579);
nor U13914 (N_13914,N_7124,N_6523);
nor U13915 (N_13915,N_6120,N_10173);
xor U13916 (N_13916,N_9730,N_8254);
nor U13917 (N_13917,N_9738,N_7851);
nand U13918 (N_13918,N_10737,N_6671);
nand U13919 (N_13919,N_10763,N_6260);
xnor U13920 (N_13920,N_11753,N_8484);
xnor U13921 (N_13921,N_10154,N_7480);
nor U13922 (N_13922,N_11631,N_10845);
nor U13923 (N_13923,N_9911,N_6936);
and U13924 (N_13924,N_7873,N_10007);
and U13925 (N_13925,N_11432,N_11568);
nand U13926 (N_13926,N_8444,N_6829);
nor U13927 (N_13927,N_11468,N_6515);
or U13928 (N_13928,N_10798,N_9364);
and U13929 (N_13929,N_9942,N_6705);
nand U13930 (N_13930,N_11228,N_11589);
nor U13931 (N_13931,N_9252,N_7814);
nor U13932 (N_13932,N_9530,N_11714);
and U13933 (N_13933,N_10709,N_8610);
xor U13934 (N_13934,N_7955,N_7337);
xnor U13935 (N_13935,N_6146,N_11293);
xnor U13936 (N_13936,N_8617,N_10496);
xnor U13937 (N_13937,N_7136,N_6287);
xor U13938 (N_13938,N_11287,N_7261);
nor U13939 (N_13939,N_11591,N_6176);
nand U13940 (N_13940,N_11685,N_7406);
nand U13941 (N_13941,N_11005,N_8428);
xnor U13942 (N_13942,N_8105,N_8930);
or U13943 (N_13943,N_9179,N_7361);
and U13944 (N_13944,N_7396,N_7887);
and U13945 (N_13945,N_10749,N_6349);
nor U13946 (N_13946,N_9001,N_8558);
nor U13947 (N_13947,N_8379,N_9997);
nor U13948 (N_13948,N_6956,N_6669);
and U13949 (N_13949,N_7404,N_9398);
nand U13950 (N_13950,N_9314,N_10401);
and U13951 (N_13951,N_10432,N_9508);
and U13952 (N_13952,N_10571,N_7381);
and U13953 (N_13953,N_8627,N_10848);
and U13954 (N_13954,N_7560,N_9471);
and U13955 (N_13955,N_6561,N_6220);
or U13956 (N_13956,N_7334,N_9289);
and U13957 (N_13957,N_11416,N_10176);
xnor U13958 (N_13958,N_10285,N_7000);
or U13959 (N_13959,N_8604,N_7779);
nor U13960 (N_13960,N_10463,N_10080);
and U13961 (N_13961,N_6644,N_6529);
xor U13962 (N_13962,N_7452,N_6210);
xor U13963 (N_13963,N_7169,N_8081);
or U13964 (N_13964,N_6235,N_7636);
and U13965 (N_13965,N_8037,N_9029);
or U13966 (N_13966,N_9161,N_8923);
and U13967 (N_13967,N_9065,N_6285);
or U13968 (N_13968,N_7654,N_9460);
and U13969 (N_13969,N_11218,N_7705);
or U13970 (N_13970,N_11000,N_11611);
and U13971 (N_13971,N_10208,N_7253);
nor U13972 (N_13972,N_8605,N_8372);
xnor U13973 (N_13973,N_11191,N_6798);
or U13974 (N_13974,N_10044,N_9421);
and U13975 (N_13975,N_7420,N_11511);
nor U13976 (N_13976,N_8543,N_10731);
nand U13977 (N_13977,N_7296,N_7621);
xnor U13978 (N_13978,N_6507,N_9076);
xnor U13979 (N_13979,N_8545,N_6919);
nand U13980 (N_13980,N_8520,N_8171);
xor U13981 (N_13981,N_7794,N_8216);
nor U13982 (N_13982,N_7416,N_6157);
nand U13983 (N_13983,N_9209,N_11295);
xnor U13984 (N_13984,N_8997,N_8962);
nand U13985 (N_13985,N_8422,N_10699);
or U13986 (N_13986,N_8741,N_10599);
and U13987 (N_13987,N_10812,N_11809);
nand U13988 (N_13988,N_10889,N_11547);
xnor U13989 (N_13989,N_9863,N_6793);
xor U13990 (N_13990,N_10262,N_10444);
and U13991 (N_13991,N_10071,N_11748);
xor U13992 (N_13992,N_6962,N_7678);
xnor U13993 (N_13993,N_6603,N_8974);
nor U13994 (N_13994,N_11740,N_7216);
nand U13995 (N_13995,N_7380,N_6892);
nand U13996 (N_13996,N_11842,N_8979);
nor U13997 (N_13997,N_8222,N_8937);
nand U13998 (N_13998,N_7316,N_8282);
and U13999 (N_13999,N_10296,N_9121);
and U14000 (N_14000,N_7740,N_11562);
and U14001 (N_14001,N_10501,N_10946);
xor U14002 (N_14002,N_8817,N_6130);
and U14003 (N_14003,N_6497,N_6276);
xor U14004 (N_14004,N_11632,N_10596);
xor U14005 (N_14005,N_6127,N_7870);
xor U14006 (N_14006,N_7649,N_10040);
and U14007 (N_14007,N_6532,N_10653);
and U14008 (N_14008,N_11187,N_7986);
nand U14009 (N_14009,N_9275,N_9798);
and U14010 (N_14010,N_10857,N_8717);
nor U14011 (N_14011,N_11385,N_6189);
nor U14012 (N_14012,N_7994,N_6085);
xnor U14013 (N_14013,N_6900,N_6647);
nor U14014 (N_14014,N_10191,N_11536);
or U14015 (N_14015,N_6448,N_10305);
nand U14016 (N_14016,N_11980,N_10779);
or U14017 (N_14017,N_11103,N_11088);
or U14018 (N_14018,N_6657,N_9564);
xnor U14019 (N_14019,N_9545,N_10093);
nor U14020 (N_14020,N_7442,N_6762);
and U14021 (N_14021,N_10687,N_6204);
and U14022 (N_14022,N_9091,N_10584);
nor U14023 (N_14023,N_6292,N_10462);
xor U14024 (N_14024,N_9406,N_6029);
or U14025 (N_14025,N_8530,N_8975);
and U14026 (N_14026,N_6373,N_8713);
nand U14027 (N_14027,N_11837,N_8874);
nand U14028 (N_14028,N_9991,N_8633);
xor U14029 (N_14029,N_10606,N_11006);
nand U14030 (N_14030,N_9333,N_8288);
and U14031 (N_14031,N_6274,N_8783);
and U14032 (N_14032,N_6104,N_10499);
xor U14033 (N_14033,N_7410,N_10648);
nor U14034 (N_14034,N_10284,N_7428);
nor U14035 (N_14035,N_6539,N_10865);
xnor U14036 (N_14036,N_6071,N_11380);
and U14037 (N_14037,N_9633,N_11392);
or U14038 (N_14038,N_10574,N_10001);
nand U14039 (N_14039,N_10723,N_7446);
nor U14040 (N_14040,N_7823,N_9315);
or U14041 (N_14041,N_7672,N_10427);
nand U14042 (N_14042,N_11698,N_11998);
or U14043 (N_14043,N_11222,N_6170);
and U14044 (N_14044,N_7834,N_6389);
xor U14045 (N_14045,N_8919,N_8632);
nor U14046 (N_14046,N_11869,N_6761);
or U14047 (N_14047,N_11947,N_10225);
xor U14048 (N_14048,N_9127,N_10298);
xor U14049 (N_14049,N_8470,N_8768);
or U14050 (N_14050,N_7209,N_6297);
and U14051 (N_14051,N_7066,N_6229);
nand U14052 (N_14052,N_6109,N_11173);
nand U14053 (N_14053,N_10459,N_6502);
or U14054 (N_14054,N_9149,N_7564);
and U14055 (N_14055,N_8673,N_7941);
and U14056 (N_14056,N_10556,N_11263);
or U14057 (N_14057,N_7637,N_9554);
or U14058 (N_14058,N_6759,N_6181);
or U14059 (N_14059,N_6624,N_8415);
nand U14060 (N_14060,N_11039,N_7606);
xnor U14061 (N_14061,N_8146,N_7340);
or U14062 (N_14062,N_11442,N_9119);
nor U14063 (N_14063,N_7506,N_7409);
nor U14064 (N_14064,N_11172,N_11683);
nor U14065 (N_14065,N_11567,N_11555);
nor U14066 (N_14066,N_7462,N_11985);
and U14067 (N_14067,N_8306,N_11193);
nor U14068 (N_14068,N_6263,N_9221);
xnor U14069 (N_14069,N_11044,N_10317);
nor U14070 (N_14070,N_6687,N_10735);
nand U14071 (N_14071,N_11059,N_9356);
nand U14072 (N_14072,N_10352,N_8183);
or U14073 (N_14073,N_6031,N_8495);
and U14074 (N_14074,N_8777,N_6208);
and U14075 (N_14075,N_9840,N_9455);
and U14076 (N_14076,N_9841,N_7045);
xor U14077 (N_14077,N_11436,N_11640);
and U14078 (N_14078,N_10439,N_9071);
and U14079 (N_14079,N_11747,N_11363);
and U14080 (N_14080,N_7133,N_7360);
and U14081 (N_14081,N_8662,N_9392);
xor U14082 (N_14082,N_11047,N_10275);
nand U14083 (N_14083,N_6277,N_8285);
xor U14084 (N_14084,N_11917,N_9518);
and U14085 (N_14085,N_11630,N_7966);
nand U14086 (N_14086,N_7698,N_8766);
or U14087 (N_14087,N_10353,N_6398);
and U14088 (N_14088,N_7114,N_8678);
and U14089 (N_14089,N_10240,N_7397);
nand U14090 (N_14090,N_10448,N_9089);
nor U14091 (N_14091,N_6026,N_7992);
nand U14092 (N_14092,N_8861,N_7398);
and U14093 (N_14093,N_6868,N_7770);
nor U14094 (N_14094,N_8044,N_8497);
nand U14095 (N_14095,N_10384,N_10794);
and U14096 (N_14096,N_6794,N_10522);
and U14097 (N_14097,N_6476,N_7711);
and U14098 (N_14098,N_8822,N_10465);
or U14099 (N_14099,N_9579,N_10088);
nand U14100 (N_14100,N_7755,N_6187);
xor U14101 (N_14101,N_11264,N_10337);
nor U14102 (N_14102,N_10569,N_8471);
and U14103 (N_14103,N_8571,N_9652);
and U14104 (N_14104,N_9098,N_10197);
xor U14105 (N_14105,N_6746,N_7855);
xnor U14106 (N_14106,N_6979,N_10212);
xor U14107 (N_14107,N_10476,N_11696);
and U14108 (N_14108,N_6834,N_8169);
nand U14109 (N_14109,N_11894,N_11652);
xor U14110 (N_14110,N_9142,N_11016);
and U14111 (N_14111,N_7853,N_6252);
xnor U14112 (N_14112,N_8841,N_9777);
or U14113 (N_14113,N_8848,N_6010);
nand U14114 (N_14114,N_7771,N_10642);
nor U14115 (N_14115,N_10089,N_9562);
nand U14116 (N_14116,N_6572,N_6673);
nand U14117 (N_14117,N_11134,N_6151);
nor U14118 (N_14118,N_6802,N_10026);
nor U14119 (N_14119,N_6155,N_8804);
or U14120 (N_14120,N_9542,N_8003);
xor U14121 (N_14121,N_9456,N_11706);
or U14122 (N_14122,N_10029,N_9572);
and U14123 (N_14123,N_8404,N_7596);
nor U14124 (N_14124,N_8235,N_9934);
and U14125 (N_14125,N_8517,N_11352);
nand U14126 (N_14126,N_6592,N_8734);
nor U14127 (N_14127,N_7430,N_11782);
or U14128 (N_14128,N_7155,N_8025);
xnor U14129 (N_14129,N_9687,N_11162);
nor U14130 (N_14130,N_11743,N_10477);
nand U14131 (N_14131,N_10369,N_11850);
xor U14132 (N_14132,N_11041,N_7978);
and U14133 (N_14133,N_6990,N_8287);
nor U14134 (N_14134,N_10576,N_9128);
or U14135 (N_14135,N_8842,N_8913);
or U14136 (N_14136,N_7996,N_8933);
nor U14137 (N_14137,N_6677,N_7542);
and U14138 (N_14138,N_8644,N_6041);
xnor U14139 (N_14139,N_7548,N_10158);
nor U14140 (N_14140,N_6883,N_10988);
or U14141 (N_14141,N_9561,N_11590);
and U14142 (N_14142,N_9359,N_10899);
xor U14143 (N_14143,N_8097,N_10308);
and U14144 (N_14144,N_6811,N_7910);
nand U14145 (N_14145,N_10451,N_6730);
or U14146 (N_14146,N_11314,N_6302);
xnor U14147 (N_14147,N_9012,N_11921);
or U14148 (N_14148,N_9683,N_8207);
nor U14149 (N_14149,N_6634,N_11690);
nor U14150 (N_14150,N_9195,N_7776);
nor U14151 (N_14151,N_9337,N_8314);
xnor U14152 (N_14152,N_7745,N_7849);
nor U14153 (N_14153,N_6217,N_9414);
xor U14154 (N_14154,N_11056,N_11009);
and U14155 (N_14155,N_9992,N_11073);
nand U14156 (N_14156,N_7648,N_8243);
xnor U14157 (N_14157,N_11832,N_6942);
nor U14158 (N_14158,N_6070,N_9234);
xor U14159 (N_14159,N_6995,N_10713);
nand U14160 (N_14160,N_10153,N_11183);
xnor U14161 (N_14161,N_9056,N_9725);
xor U14162 (N_14162,N_11107,N_7700);
or U14163 (N_14163,N_7149,N_7985);
and U14164 (N_14164,N_8199,N_9621);
nor U14165 (N_14165,N_8854,N_9443);
or U14166 (N_14166,N_11663,N_9401);
and U14167 (N_14167,N_6909,N_9201);
or U14168 (N_14168,N_11411,N_8149);
xor U14169 (N_14169,N_7434,N_6384);
xor U14170 (N_14170,N_6570,N_7766);
and U14171 (N_14171,N_11658,N_8556);
and U14172 (N_14172,N_6946,N_9437);
and U14173 (N_14173,N_8033,N_10886);
and U14174 (N_14174,N_7733,N_8054);
nand U14175 (N_14175,N_6385,N_9274);
and U14176 (N_14176,N_8820,N_10074);
or U14177 (N_14177,N_10997,N_8647);
nand U14178 (N_14178,N_9125,N_8739);
and U14179 (N_14179,N_8600,N_9901);
xnor U14180 (N_14180,N_10758,N_11177);
nor U14181 (N_14181,N_8176,N_8995);
or U14182 (N_14182,N_6672,N_9253);
nor U14183 (N_14183,N_6697,N_7384);
or U14184 (N_14184,N_8065,N_11036);
nand U14185 (N_14185,N_11849,N_6096);
nor U14186 (N_14186,N_11182,N_7619);
nand U14187 (N_14187,N_6477,N_11464);
and U14188 (N_14188,N_9205,N_8250);
nor U14189 (N_14189,N_11026,N_11345);
and U14190 (N_14190,N_6132,N_6751);
nor U14191 (N_14191,N_11502,N_7693);
or U14192 (N_14192,N_10559,N_8256);
nor U14193 (N_14193,N_8311,N_8934);
xnor U14194 (N_14194,N_8829,N_9743);
nor U14195 (N_14195,N_8908,N_9412);
and U14196 (N_14196,N_9304,N_8877);
nor U14197 (N_14197,N_10349,N_10058);
xnor U14198 (N_14198,N_9935,N_11836);
or U14199 (N_14199,N_8483,N_6602);
and U14200 (N_14200,N_9284,N_9756);
xor U14201 (N_14201,N_11215,N_7075);
or U14202 (N_14202,N_9297,N_7922);
nor U14203 (N_14203,N_8230,N_8922);
and U14204 (N_14204,N_11075,N_11027);
nor U14205 (N_14205,N_8463,N_10169);
or U14206 (N_14206,N_10259,N_10263);
nor U14207 (N_14207,N_9998,N_7673);
xor U14208 (N_14208,N_9472,N_8609);
xnor U14209 (N_14209,N_10517,N_8946);
nand U14210 (N_14210,N_11400,N_8302);
nor U14211 (N_14211,N_11021,N_8268);
nand U14212 (N_14212,N_10041,N_9822);
and U14213 (N_14213,N_6659,N_8353);
nand U14214 (N_14214,N_6589,N_8598);
xnor U14215 (N_14215,N_10155,N_7977);
nand U14216 (N_14216,N_8480,N_9268);
or U14217 (N_14217,N_10525,N_9273);
xnor U14218 (N_14218,N_7709,N_7312);
and U14219 (N_14219,N_8043,N_7322);
xnor U14220 (N_14220,N_7444,N_11025);
xor U14221 (N_14221,N_7638,N_6886);
and U14222 (N_14222,N_10492,N_9535);
nor U14223 (N_14223,N_6464,N_9095);
and U14224 (N_14224,N_7567,N_7146);
or U14225 (N_14225,N_8186,N_6563);
and U14226 (N_14226,N_8087,N_9839);
xnor U14227 (N_14227,N_8623,N_8447);
nand U14228 (N_14228,N_8182,N_10290);
and U14229 (N_14229,N_7175,N_7059);
and U14230 (N_14230,N_10745,N_9511);
nand U14231 (N_14231,N_6107,N_7517);
and U14232 (N_14232,N_10911,N_11827);
and U14233 (N_14233,N_10083,N_8030);
and U14234 (N_14234,N_7178,N_6715);
and U14235 (N_14235,N_9596,N_10531);
nand U14236 (N_14236,N_10164,N_7924);
nor U14237 (N_14237,N_7867,N_8730);
and U14238 (N_14238,N_9393,N_9556);
and U14239 (N_14239,N_10716,N_7113);
nand U14240 (N_14240,N_11453,N_9395);
xor U14241 (N_14241,N_7359,N_6583);
xor U14242 (N_14242,N_8503,N_6873);
and U14243 (N_14243,N_8375,N_6456);
nand U14244 (N_14244,N_8947,N_9038);
xnor U14245 (N_14245,N_10833,N_8867);
and U14246 (N_14246,N_6271,N_11961);
nor U14247 (N_14247,N_7622,N_7944);
xor U14248 (N_14248,N_10983,N_11203);
nor U14249 (N_14249,N_6370,N_9383);
or U14250 (N_14250,N_11216,N_10446);
and U14251 (N_14251,N_9736,N_7090);
nand U14252 (N_14252,N_9151,N_10674);
or U14253 (N_14253,N_9074,N_7588);
or U14254 (N_14254,N_11444,N_9229);
xnor U14255 (N_14255,N_7439,N_9708);
nand U14256 (N_14256,N_9054,N_6785);
nand U14257 (N_14257,N_6784,N_9956);
or U14258 (N_14258,N_11410,N_9940);
nand U14259 (N_14259,N_8148,N_6250);
nor U14260 (N_14260,N_9782,N_7615);
xnor U14261 (N_14261,N_8427,N_9160);
or U14262 (N_14262,N_7640,N_7100);
xnor U14263 (N_14263,N_9945,N_10241);
or U14264 (N_14264,N_8385,N_11291);
nor U14265 (N_14265,N_7875,N_8055);
xnor U14266 (N_14266,N_6611,N_8193);
nor U14267 (N_14267,N_8196,N_9550);
or U14268 (N_14268,N_8452,N_11388);
and U14269 (N_14269,N_11990,N_7201);
or U14270 (N_14270,N_9686,N_8029);
nor U14271 (N_14271,N_10347,N_10846);
xor U14272 (N_14272,N_6878,N_8893);
xnor U14273 (N_14273,N_7311,N_8244);
or U14274 (N_14274,N_10982,N_10513);
nor U14275 (N_14275,N_10871,N_8343);
or U14276 (N_14276,N_6642,N_6872);
nand U14277 (N_14277,N_11492,N_11305);
nor U14278 (N_14278,N_6650,N_11594);
nand U14279 (N_14279,N_8457,N_7778);
and U14280 (N_14280,N_9292,N_8295);
and U14281 (N_14281,N_8740,N_10414);
nand U14282 (N_14282,N_9999,N_10691);
or U14283 (N_14283,N_9446,N_10610);
and U14284 (N_14284,N_6046,N_10313);
nor U14285 (N_14285,N_8454,N_9022);
nor U14286 (N_14286,N_9042,N_7718);
xor U14287 (N_14287,N_8909,N_6852);
nand U14288 (N_14288,N_6664,N_7148);
or U14289 (N_14289,N_11082,N_8206);
xor U14290 (N_14290,N_11875,N_6184);
xor U14291 (N_14291,N_7438,N_6992);
nor U14292 (N_14292,N_6470,N_11231);
or U14293 (N_14293,N_10231,N_8523);
or U14294 (N_14294,N_8987,N_11935);
nor U14295 (N_14295,N_10181,N_10681);
xnor U14296 (N_14296,N_8064,N_8036);
or U14297 (N_14297,N_6726,N_8839);
or U14298 (N_14298,N_7067,N_9415);
or U14299 (N_14299,N_10818,N_8672);
and U14300 (N_14300,N_9343,N_9837);
nand U14301 (N_14301,N_8619,N_6524);
or U14302 (N_14302,N_9339,N_11322);
xnor U14303 (N_14303,N_11304,N_10020);
and U14304 (N_14304,N_10008,N_6783);
or U14305 (N_14305,N_6013,N_11045);
or U14306 (N_14306,N_8056,N_8593);
xor U14307 (N_14307,N_7750,N_9954);
nand U14308 (N_14308,N_11070,N_11870);
nor U14309 (N_14309,N_7266,N_9023);
nand U14310 (N_14310,N_7411,N_7971);
and U14311 (N_14311,N_7195,N_6022);
nand U14312 (N_14312,N_6997,N_7611);
nor U14313 (N_14313,N_7036,N_10441);
or U14314 (N_14314,N_8473,N_11817);
nor U14315 (N_14315,N_6728,N_6815);
or U14316 (N_14316,N_7882,N_10073);
nand U14317 (N_14317,N_7820,N_6367);
nor U14318 (N_14318,N_7927,N_7016);
and U14319 (N_14319,N_9866,N_6914);
xnor U14320 (N_14320,N_8367,N_10985);
xor U14321 (N_14321,N_10598,N_11061);
xor U14322 (N_14322,N_8401,N_8969);
or U14323 (N_14323,N_9876,N_11448);
and U14324 (N_14324,N_10440,N_11083);
xor U14325 (N_14325,N_6049,N_10230);
xnor U14326 (N_14326,N_9980,N_8596);
nand U14327 (N_14327,N_9806,N_6714);
and U14328 (N_14328,N_6268,N_11338);
nor U14329 (N_14329,N_10187,N_10881);
or U14330 (N_14330,N_6363,N_11359);
or U14331 (N_14331,N_10053,N_8597);
xor U14332 (N_14332,N_10639,N_9464);
or U14333 (N_14333,N_11538,N_8693);
or U14334 (N_14334,N_6609,N_9318);
and U14335 (N_14335,N_9880,N_8884);
or U14336 (N_14336,N_6215,N_6205);
xor U14337 (N_14337,N_11800,N_11587);
nor U14338 (N_14338,N_6557,N_8507);
nand U14339 (N_14339,N_6056,N_10027);
xor U14340 (N_14340,N_10398,N_10546);
nor U14341 (N_14341,N_9647,N_6394);
and U14342 (N_14342,N_7857,N_10915);
or U14343 (N_14343,N_7433,N_11161);
or U14344 (N_14344,N_6810,N_6787);
nand U14345 (N_14345,N_8897,N_8085);
xnor U14346 (N_14346,N_9821,N_10450);
xnor U14347 (N_14347,N_9497,N_6322);
nor U14348 (N_14348,N_11766,N_6001);
nand U14349 (N_14349,N_7382,N_6433);
nand U14350 (N_14350,N_7286,N_9057);
nor U14351 (N_14351,N_8458,N_11999);
and U14352 (N_14352,N_9775,N_9491);
xor U14353 (N_14353,N_11945,N_6768);
nand U14354 (N_14354,N_6790,N_8557);
xnor U14355 (N_14355,N_10613,N_11030);
nand U14356 (N_14356,N_8220,N_7129);
and U14357 (N_14357,N_6326,N_6588);
nor U14358 (N_14358,N_9021,N_7271);
and U14359 (N_14359,N_10548,N_11253);
nor U14360 (N_14360,N_7391,N_9639);
and U14361 (N_14361,N_6251,N_6558);
nand U14362 (N_14362,N_9245,N_7053);
nor U14363 (N_14363,N_11050,N_11751);
nor U14364 (N_14364,N_11598,N_10968);
or U14365 (N_14365,N_6265,N_6183);
and U14366 (N_14366,N_9674,N_9494);
xnor U14367 (N_14367,N_11033,N_8902);
nor U14368 (N_14368,N_7777,N_8502);
nand U14369 (N_14369,N_9016,N_9087);
xor U14370 (N_14370,N_8864,N_9256);
nor U14371 (N_14371,N_9597,N_6166);
nand U14372 (N_14372,N_8921,N_6817);
nor U14373 (N_14373,N_9826,N_7516);
nor U14374 (N_14374,N_7221,N_8127);
nand U14375 (N_14375,N_10722,N_10334);
nand U14376 (N_14376,N_8469,N_6088);
and U14377 (N_14377,N_11261,N_9505);
xnor U14378 (N_14378,N_9207,N_11111);
nor U14379 (N_14379,N_9678,N_11549);
and U14380 (N_14380,N_7062,N_8830);
nor U14381 (N_14381,N_7318,N_9244);
xor U14382 (N_14382,N_8752,N_11784);
nand U14383 (N_14383,N_10885,N_11984);
and U14384 (N_14384,N_6116,N_11497);
nand U14385 (N_14385,N_7793,N_9283);
nand U14386 (N_14386,N_10739,N_10967);
nand U14387 (N_14387,N_9789,N_11408);
xor U14388 (N_14388,N_9377,N_6924);
and U14389 (N_14389,N_7235,N_11636);
xor U14390 (N_14390,N_11072,N_9162);
nor U14391 (N_14391,N_6925,N_8013);
nand U14392 (N_14392,N_11085,N_7707);
nor U14393 (N_14393,N_11560,N_8368);
and U14394 (N_14394,N_6816,N_8991);
and U14395 (N_14395,N_7811,N_7889);
xnor U14396 (N_14396,N_11284,N_7959);
nor U14397 (N_14397,N_11230,N_11362);
nand U14398 (N_14398,N_9217,N_6699);
xnor U14399 (N_14399,N_9327,N_9831);
and U14400 (N_14400,N_9370,N_10460);
and U14401 (N_14401,N_7344,N_6901);
and U14402 (N_14402,N_9031,N_8387);
nand U14403 (N_14403,N_6977,N_11807);
nor U14404 (N_14404,N_6960,N_7624);
or U14405 (N_14405,N_6854,N_9908);
or U14406 (N_14406,N_11435,N_11741);
nor U14407 (N_14407,N_9137,N_9805);
nand U14408 (N_14408,N_10769,N_8824);
xnor U14409 (N_14409,N_11625,N_9541);
xnor U14410 (N_14410,N_7025,N_11447);
nor U14411 (N_14411,N_10755,N_8091);
or U14412 (N_14412,N_6559,N_7385);
xor U14413 (N_14413,N_7504,N_8177);
and U14414 (N_14414,N_7940,N_9899);
nor U14415 (N_14415,N_8992,N_7991);
nand U14416 (N_14416,N_8006,N_9864);
nor U14417 (N_14417,N_7591,N_10234);
and U14418 (N_14418,N_10961,N_10248);
and U14419 (N_14419,N_6020,N_9342);
nor U14420 (N_14420,N_8686,N_7554);
and U14421 (N_14421,N_10840,N_6479);
and U14422 (N_14422,N_8294,N_11899);
or U14423 (N_14423,N_9129,N_7338);
and U14424 (N_14424,N_6665,N_9889);
nor U14425 (N_14425,N_11330,N_6206);
xnor U14426 (N_14426,N_8082,N_6853);
nand U14427 (N_14427,N_11431,N_7031);
and U14428 (N_14428,N_9048,N_9015);
nor U14429 (N_14429,N_8955,N_10678);
xnor U14430 (N_14430,N_8279,N_6885);
nor U14431 (N_14431,N_6035,N_6709);
or U14432 (N_14432,N_10793,N_11124);
xor U14433 (N_14433,N_6225,N_11037);
nand U14434 (N_14434,N_8620,N_6733);
xor U14435 (N_14435,N_6172,N_9783);
or U14436 (N_14436,N_10393,N_7210);
nand U14437 (N_14437,N_8654,N_8305);
nand U14438 (N_14438,N_10422,N_10898);
and U14439 (N_14439,N_9759,N_8051);
and U14440 (N_14440,N_9978,N_7639);
or U14441 (N_14441,N_8391,N_8834);
or U14442 (N_14442,N_9132,N_6425);
and U14443 (N_14443,N_7007,N_10018);
and U14444 (N_14444,N_6431,N_11332);
and U14445 (N_14445,N_6542,N_7706);
or U14446 (N_14446,N_8837,N_7118);
nor U14447 (N_14447,N_11199,N_7268);
nand U14448 (N_14448,N_11995,N_10939);
and U14449 (N_14449,N_8905,N_9842);
nand U14450 (N_14450,N_11475,N_7543);
or U14451 (N_14451,N_8675,N_9681);
nor U14452 (N_14452,N_11699,N_7243);
xor U14453 (N_14453,N_6904,N_9476);
nand U14454 (N_14454,N_8993,N_11505);
or U14455 (N_14455,N_9744,N_11499);
and U14456 (N_14456,N_8348,N_8552);
or U14457 (N_14457,N_6242,N_9067);
and U14458 (N_14458,N_9014,N_9853);
nor U14459 (N_14459,N_7628,N_9218);
xor U14460 (N_14460,N_11128,N_11912);
xor U14461 (N_14461,N_9293,N_11707);
xor U14462 (N_14462,N_8901,N_8035);
xnor U14463 (N_14463,N_6981,N_8737);
xor U14464 (N_14464,N_10138,N_10920);
or U14465 (N_14465,N_6122,N_8796);
and U14466 (N_14466,N_7309,N_11739);
and U14467 (N_14467,N_11866,N_9865);
nand U14468 (N_14468,N_10828,N_11369);
xnor U14469 (N_14469,N_11641,N_9353);
nor U14470 (N_14470,N_9538,N_8371);
nand U14471 (N_14471,N_8430,N_8041);
nor U14472 (N_14472,N_6136,N_11349);
nand U14473 (N_14473,N_7604,N_9704);
nand U14474 (N_14474,N_8745,N_7030);
or U14475 (N_14475,N_9583,N_9733);
nand U14476 (N_14476,N_11126,N_11142);
and U14477 (N_14477,N_8951,N_11438);
xnor U14478 (N_14478,N_11674,N_6841);
or U14479 (N_14479,N_7267,N_9531);
nand U14480 (N_14480,N_10600,N_6550);
or U14481 (N_14481,N_11462,N_9694);
nand U14482 (N_14482,N_9341,N_6329);
nor U14483 (N_14483,N_9593,N_10526);
or U14484 (N_14484,N_7951,N_10994);
nand U14485 (N_14485,N_9146,N_7451);
and U14486 (N_14486,N_10157,N_7934);
xor U14487 (N_14487,N_7600,N_9917);
xor U14488 (N_14488,N_9823,N_10021);
xor U14489 (N_14489,N_10979,N_6851);
or U14490 (N_14490,N_11907,N_10601);
xor U14491 (N_14491,N_11512,N_11987);
nand U14492 (N_14492,N_11759,N_6681);
nor U14493 (N_14493,N_10403,N_7010);
nand U14494 (N_14494,N_6148,N_7632);
xnor U14495 (N_14495,N_6555,N_7006);
or U14496 (N_14496,N_7593,N_6766);
xor U14497 (N_14497,N_10006,N_6318);
xnor U14498 (N_14498,N_9448,N_6404);
or U14499 (N_14499,N_11084,N_11414);
xor U14500 (N_14500,N_9052,N_8729);
and U14501 (N_14501,N_8048,N_7313);
nor U14502 (N_14502,N_6632,N_7350);
or U14503 (N_14503,N_7319,N_11186);
nor U14504 (N_14504,N_8429,N_11157);
or U14505 (N_14505,N_6231,N_9702);
nand U14506 (N_14506,N_10100,N_6857);
or U14507 (N_14507,N_9638,N_9979);
and U14508 (N_14508,N_6899,N_9549);
or U14509 (N_14509,N_11396,N_11132);
and U14510 (N_14510,N_9068,N_7034);
xnor U14511 (N_14511,N_11282,N_11237);
xor U14512 (N_14512,N_11876,N_11828);
or U14513 (N_14513,N_11968,N_8280);
nand U14514 (N_14514,N_7911,N_10288);
and U14515 (N_14515,N_11576,N_8262);
nand U14516 (N_14516,N_11596,N_6034);
xor U14517 (N_14517,N_7738,N_11415);
xor U14518 (N_14518,N_7082,N_11469);
nand U14519 (N_14519,N_10227,N_7581);
or U14520 (N_14520,N_6809,N_7859);
or U14521 (N_14521,N_9915,N_11018);
nor U14522 (N_14522,N_6772,N_10957);
or U14523 (N_14523,N_9321,N_7546);
or U14524 (N_14524,N_10282,N_8047);
nand U14525 (N_14525,N_11629,N_11301);
nor U14526 (N_14526,N_10402,N_10070);
and U14527 (N_14527,N_7722,N_6732);
xnor U14528 (N_14528,N_11201,N_7366);
or U14529 (N_14529,N_8412,N_10766);
or U14530 (N_14530,N_8011,N_9812);
nand U14531 (N_14531,N_8863,N_10200);
or U14532 (N_14532,N_9655,N_10061);
and U14533 (N_14533,N_7314,N_7389);
and U14534 (N_14534,N_6881,N_7326);
and U14535 (N_14535,N_8695,N_7207);
or U14536 (N_14536,N_9963,N_11882);
and U14537 (N_14537,N_10361,N_8898);
or U14538 (N_14538,N_10852,N_11042);
and U14539 (N_14539,N_7748,N_9696);
nor U14540 (N_14540,N_11970,N_10697);
xnor U14541 (N_14541,N_7461,N_10042);
xnor U14542 (N_14542,N_6442,N_9334);
xor U14543 (N_14543,N_6084,N_9331);
nor U14544 (N_14544,N_7329,N_9136);
and U14545 (N_14545,N_9951,N_9680);
nand U14546 (N_14546,N_6298,N_9566);
nor U14547 (N_14547,N_9914,N_8499);
or U14548 (N_14548,N_11089,N_9255);
xor U14549 (N_14549,N_7181,N_8016);
xnor U14550 (N_14550,N_8744,N_10178);
and U14551 (N_14551,N_10907,N_8682);
and U14552 (N_14552,N_11122,N_7655);
and U14553 (N_14553,N_8949,N_6332);
and U14554 (N_14554,N_11350,N_11181);
nand U14555 (N_14555,N_6055,N_7800);
nor U14556 (N_14556,N_10043,N_8488);
xnor U14557 (N_14557,N_6952,N_11262);
or U14558 (N_14558,N_8202,N_9881);
or U14559 (N_14559,N_11633,N_7193);
or U14560 (N_14560,N_10196,N_11834);
nor U14561 (N_14561,N_10893,N_9020);
nor U14562 (N_14562,N_10650,N_9150);
xnor U14563 (N_14563,N_9918,N_10844);
or U14564 (N_14564,N_11225,N_8999);
nand U14565 (N_14565,N_10897,N_11246);
xnor U14566 (N_14566,N_11950,N_6630);
xnor U14567 (N_14567,N_10540,N_6530);
nand U14568 (N_14568,N_8496,N_9924);
and U14569 (N_14569,N_6485,N_9211);
and U14570 (N_14570,N_9257,N_11791);
xor U14571 (N_14571,N_7987,N_11733);
or U14572 (N_14572,N_6619,N_10237);
nor U14573 (N_14573,N_10382,N_6623);
or U14574 (N_14574,N_11891,N_11390);
or U14575 (N_14575,N_8112,N_9787);
nand U14576 (N_14576,N_10872,N_11765);
xor U14577 (N_14577,N_6612,N_8670);
nor U14578 (N_14578,N_9090,N_7502);
and U14579 (N_14579,N_11944,N_8705);
and U14580 (N_14580,N_10301,N_7033);
nor U14581 (N_14581,N_11943,N_8478);
xnor U14582 (N_14582,N_6337,N_6622);
and U14583 (N_14583,N_6399,N_10976);
xor U14584 (N_14584,N_10631,N_6169);
xnor U14585 (N_14585,N_9890,N_7835);
and U14586 (N_14586,N_11767,N_11969);
or U14587 (N_14587,N_11838,N_9240);
or U14588 (N_14588,N_6943,N_7583);
xor U14589 (N_14589,N_7130,N_11356);
or U14590 (N_14590,N_9177,N_9230);
xnor U14591 (N_14591,N_6115,N_6163);
xor U14592 (N_14592,N_7379,N_11665);
nand U14593 (N_14593,N_10354,N_7989);
or U14594 (N_14594,N_9547,N_9939);
xor U14595 (N_14595,N_8045,N_7466);
nand U14596 (N_14596,N_9995,N_10144);
or U14597 (N_14597,N_10213,N_11754);
xnor U14598 (N_14598,N_8018,N_11459);
or U14599 (N_14599,N_11297,N_9017);
or U14600 (N_14600,N_9197,N_9376);
nor U14601 (N_14601,N_8061,N_11450);
nand U14602 (N_14602,N_9104,N_6831);
nor U14603 (N_14603,N_9346,N_6162);
and U14604 (N_14604,N_6323,N_6727);
and U14605 (N_14605,N_8289,N_10884);
xor U14606 (N_14606,N_10125,N_8324);
or U14607 (N_14607,N_10585,N_11371);
xor U14608 (N_14608,N_11814,N_6537);
and U14609 (N_14609,N_11908,N_10553);
xnor U14610 (N_14610,N_7168,N_11873);
or U14611 (N_14611,N_7723,N_10607);
xnor U14612 (N_14612,N_7484,N_10461);
nor U14613 (N_14613,N_8651,N_9776);
xor U14614 (N_14614,N_10316,N_9176);
and U14615 (N_14615,N_8636,N_8178);
nand U14616 (N_14616,N_6429,N_9028);
xnor U14617 (N_14617,N_7373,N_7342);
xor U14618 (N_14618,N_6779,N_10279);
and U14619 (N_14619,N_8561,N_10060);
and U14620 (N_14620,N_11695,N_10959);
or U14621 (N_14621,N_7528,N_6445);
xnor U14622 (N_14622,N_9933,N_6889);
nand U14623 (N_14623,N_9585,N_11159);
nand U14624 (N_14624,N_6227,N_11437);
nor U14625 (N_14625,N_11361,N_10453);
or U14626 (N_14626,N_9228,N_6631);
nand U14627 (N_14627,N_7107,N_8238);
and U14628 (N_14628,N_6791,N_9324);
and U14629 (N_14629,N_6536,N_6432);
xnor U14630 (N_14630,N_6335,N_7881);
or U14631 (N_14631,N_8943,N_10738);
nor U14632 (N_14632,N_6042,N_11048);
xor U14633 (N_14633,N_8157,N_11109);
nor U14634 (N_14634,N_8564,N_8363);
nand U14635 (N_14635,N_8716,N_6720);
and U14636 (N_14636,N_6600,N_6245);
xor U14637 (N_14637,N_6934,N_8573);
nor U14638 (N_14638,N_8260,N_7592);
xor U14639 (N_14639,N_8300,N_7029);
nand U14640 (N_14640,N_7552,N_9267);
or U14641 (N_14641,N_10480,N_9492);
xnor U14642 (N_14642,N_8023,N_6098);
nor U14643 (N_14643,N_6408,N_8402);
and U14644 (N_14644,N_11303,N_11252);
xnor U14645 (N_14645,N_8212,N_6261);
xnor U14646 (N_14646,N_7651,N_10331);
xor U14647 (N_14647,N_8658,N_9689);
xnor U14648 (N_14648,N_10552,N_8190);
and U14649 (N_14649,N_10799,N_7003);
xor U14650 (N_14650,N_9830,N_11195);
or U14651 (N_14651,N_7598,N_6179);
or U14652 (N_14652,N_6983,N_11521);
and U14653 (N_14653,N_8004,N_11057);
or U14654 (N_14654,N_7848,N_6002);
nand U14655 (N_14655,N_11881,N_11343);
and U14656 (N_14656,N_10395,N_11727);
nand U14657 (N_14657,N_6782,N_9698);
or U14658 (N_14658,N_11167,N_11627);
xnor U14659 (N_14659,N_9820,N_10126);
nor U14660 (N_14660,N_9967,N_9504);
or U14661 (N_14661,N_7969,N_8918);
xor U14662 (N_14662,N_8466,N_7732);
xnor U14663 (N_14663,N_10802,N_11992);
nor U14664 (N_14664,N_7488,N_11862);
xor U14665 (N_14665,N_10661,N_11835);
nor U14666 (N_14666,N_7575,N_6270);
or U14667 (N_14667,N_8173,N_11310);
or U14668 (N_14668,N_7098,N_8420);
and U14669 (N_14669,N_9285,N_7822);
nor U14670 (N_14670,N_10429,N_11609);
xor U14671 (N_14671,N_7782,N_7001);
or U14672 (N_14672,N_11604,N_10651);
and U14673 (N_14673,N_9987,N_11792);
nor U14674 (N_14674,N_8948,N_11735);
or U14675 (N_14675,N_7498,N_10518);
nor U14676 (N_14676,N_7372,N_11010);
nand U14677 (N_14677,N_6106,N_10666);
or U14678 (N_14678,N_7871,N_7218);
nor U14679 (N_14679,N_9667,N_9264);
or U14680 (N_14680,N_7998,N_8803);
nand U14681 (N_14681,N_8440,N_8380);
and U14682 (N_14682,N_7931,N_7536);
nor U14683 (N_14683,N_7425,N_8439);
nor U14684 (N_14684,N_9422,N_6057);
or U14685 (N_14685,N_8821,N_11892);
nor U14686 (N_14686,N_7618,N_7105);
nand U14687 (N_14687,N_6796,N_6378);
and U14688 (N_14688,N_7829,N_7802);
nand U14689 (N_14689,N_8835,N_7630);
nor U14690 (N_14690,N_9928,N_11062);
xor U14691 (N_14691,N_11745,N_9797);
nor U14692 (N_14692,N_10528,N_9610);
or U14693 (N_14693,N_9516,N_9870);
and U14694 (N_14694,N_7960,N_7780);
xor U14695 (N_14695,N_9427,N_8072);
or U14696 (N_14696,N_6203,N_9171);
and U14697 (N_14697,N_7816,N_6703);
nand U14698 (N_14698,N_8553,N_9955);
nand U14699 (N_14699,N_10791,N_9947);
or U14700 (N_14700,N_11333,N_11675);
nor U14701 (N_14701,N_8811,N_8291);
and U14702 (N_14702,N_10411,N_10464);
and U14703 (N_14703,N_7097,N_10873);
or U14704 (N_14704,N_8840,N_7282);
and U14705 (N_14705,N_6352,N_8857);
nor U14706 (N_14706,N_9968,N_6436);
nand U14707 (N_14707,N_8976,N_6366);
nand U14708 (N_14708,N_10633,N_6165);
or U14709 (N_14709,N_6062,N_10405);
and U14710 (N_14710,N_8542,N_10520);
and U14711 (N_14711,N_6133,N_8436);
or U14712 (N_14712,N_9108,N_9247);
nor U14713 (N_14713,N_8750,N_9767);
or U14714 (N_14714,N_7792,N_9007);
or U14715 (N_14715,N_10629,N_6567);
or U14716 (N_14716,N_9216,N_11331);
nand U14717 (N_14717,N_6913,N_7694);
nor U14718 (N_14718,N_7248,N_6660);
or U14719 (N_14719,N_11515,N_6753);
or U14720 (N_14720,N_9624,N_9949);
nand U14721 (N_14721,N_8845,N_9444);
and U14722 (N_14722,N_11466,N_10327);
nand U14723 (N_14723,N_9055,N_11214);
nand U14724 (N_14724,N_7799,N_9096);
and U14725 (N_14725,N_8891,N_10172);
xor U14726 (N_14726,N_8411,N_8726);
nor U14727 (N_14727,N_7828,N_6233);
nor U14728 (N_14728,N_9141,N_11790);
and U14729 (N_14729,N_7565,N_11445);
nand U14730 (N_14730,N_7896,N_9567);
nor U14731 (N_14731,N_8917,N_9703);
or U14732 (N_14732,N_10371,N_11212);
and U14733 (N_14733,N_9276,N_10037);
nor U14734 (N_14734,N_6812,N_11119);
and U14735 (N_14735,N_11717,N_7841);
nand U14736 (N_14736,N_6531,N_6461);
nor U14737 (N_14737,N_9039,N_8449);
xor U14738 (N_14738,N_11398,N_7403);
and U14739 (N_14739,N_10204,N_11273);
xnor U14740 (N_14740,N_6177,N_11165);
nor U14741 (N_14741,N_6300,N_9717);
xor U14742 (N_14742,N_10590,N_6087);
or U14743 (N_14743,N_10509,N_9800);
nand U14744 (N_14744,N_11523,N_6654);
or U14745 (N_14745,N_10734,N_7891);
xnor U14746 (N_14746,N_9728,N_9559);
or U14747 (N_14747,N_10913,N_11205);
xor U14748 (N_14748,N_6003,N_7975);
or U14749 (N_14749,N_8432,N_6198);
or U14750 (N_14750,N_7496,N_8961);
and U14751 (N_14751,N_6966,N_9568);
and U14752 (N_14752,N_10028,N_10357);
nand U14753 (N_14753,N_10925,N_6191);
or U14754 (N_14754,N_8761,N_7465);
and U14755 (N_14755,N_11256,N_8028);
xnor U14756 (N_14756,N_10318,N_6391);
nand U14757 (N_14757,N_8008,N_9277);
xnor U14758 (N_14758,N_7481,N_7421);
nand U14759 (N_14759,N_7437,N_6736);
nand U14760 (N_14760,N_11306,N_10431);
xor U14761 (N_14761,N_11798,N_8389);
xor U14762 (N_14762,N_8121,N_9846);
or U14763 (N_14763,N_7048,N_11489);
or U14764 (N_14764,N_11712,N_11529);
nor U14765 (N_14765,N_10022,N_11540);
and U14766 (N_14766,N_11697,N_7715);
xnor U14767 (N_14767,N_8310,N_8628);
and U14768 (N_14768,N_8062,N_10303);
nand U14769 (N_14769,N_8688,N_11439);
and U14770 (N_14770,N_9402,N_9713);
nor U14771 (N_14771,N_8689,N_9600);
nor U14772 (N_14772,N_9147,N_9598);
or U14773 (N_14773,N_6024,N_7152);
nor U14774 (N_14774,N_9018,N_8226);
nor U14775 (N_14775,N_9649,N_7519);
xnor U14776 (N_14776,N_11544,N_9168);
nand U14777 (N_14777,N_7189,N_6114);
and U14778 (N_14778,N_8519,N_11854);
or U14779 (N_14779,N_6778,N_8494);
xor U14780 (N_14780,N_7270,N_8895);
nor U14781 (N_14781,N_7539,N_6896);
nand U14782 (N_14782,N_8150,N_10695);
xnor U14783 (N_14783,N_9323,N_9560);
or U14784 (N_14784,N_9322,N_7272);
xnor U14785 (N_14785,N_9878,N_6595);
nand U14786 (N_14786,N_8050,N_7580);
or U14787 (N_14787,N_9636,N_9320);
xor U14788 (N_14788,N_7838,N_11823);
and U14789 (N_14789,N_11100,N_6090);
xnor U14790 (N_14790,N_10934,N_6498);
or U14791 (N_14791,N_9943,N_7957);
nand U14792 (N_14792,N_8866,N_11965);
xnor U14793 (N_14793,N_6054,N_6253);
and U14794 (N_14794,N_7586,N_9332);
xor U14795 (N_14795,N_9905,N_9790);
nand U14796 (N_14796,N_10177,N_10693);
nor U14797 (N_14797,N_11802,N_7553);
and U14798 (N_14798,N_9164,N_8409);
xnor U14799 (N_14799,N_11412,N_6086);
nand U14800 (N_14800,N_10408,N_11130);
or U14801 (N_14801,N_11146,N_6447);
or U14802 (N_14802,N_7153,N_8094);
nand U14803 (N_14803,N_11581,N_10901);
xnor U14804 (N_14804,N_9242,N_6662);
or U14805 (N_14805,N_6486,N_7644);
and U14806 (N_14806,N_8844,N_7682);
xor U14807 (N_14807,N_11317,N_6578);
nand U14808 (N_14808,N_11341,N_6822);
nor U14809 (N_14809,N_9466,N_8210);
and U14810 (N_14810,N_7339,N_8892);
nand U14811 (N_14811,N_10640,N_7675);
and U14812 (N_14812,N_10410,N_10954);
xor U14813 (N_14813,N_6640,N_6916);
xnor U14814 (N_14814,N_6656,N_9710);
and U14815 (N_14815,N_11949,N_8010);
nand U14816 (N_14816,N_8719,N_10921);
xnor U14817 (N_14817,N_11779,N_6993);
and U14818 (N_14818,N_6336,N_9761);
or U14819 (N_14819,N_9282,N_7390);
nor U14820 (N_14820,N_10502,N_10311);
nor U14821 (N_14821,N_7903,N_10374);
xor U14822 (N_14822,N_10149,N_11340);
nand U14823 (N_14823,N_6380,N_6880);
nor U14824 (N_14824,N_9534,N_8414);
and U14825 (N_14825,N_8869,N_10904);
nand U14826 (N_14826,N_9135,N_7988);
nor U14827 (N_14827,N_7184,N_9855);
and U14828 (N_14828,N_8618,N_8012);
xor U14829 (N_14829,N_10777,N_8862);
xnor U14830 (N_14830,N_8337,N_7277);
or U14831 (N_14831,N_8959,N_8546);
and U14832 (N_14832,N_7972,N_9930);
nand U14833 (N_14833,N_11079,N_7689);
nor U14834 (N_14834,N_10338,N_6124);
xnor U14835 (N_14835,N_7518,N_11478);
and U14836 (N_14836,N_8819,N_7236);
nand U14837 (N_14837,N_11577,N_7112);
nand U14838 (N_14838,N_10030,N_6063);
or U14839 (N_14839,N_8000,N_10854);
or U14840 (N_14840,N_7525,N_7906);
nor U14841 (N_14841,N_9714,N_8107);
or U14842 (N_14842,N_9887,N_9834);
or U14843 (N_14843,N_6606,N_10013);
nor U14844 (N_14844,N_11682,N_6484);
nor U14845 (N_14845,N_9366,N_11829);
or U14846 (N_14846,N_7280,N_9528);
xor U14847 (N_14847,N_7515,N_6649);
or U14848 (N_14848,N_6985,N_10906);
nor U14849 (N_14849,N_8410,N_8954);
and U14850 (N_14850,N_7295,N_11728);
nor U14851 (N_14851,N_9539,N_8423);
xor U14852 (N_14852,N_7491,N_9030);
nor U14853 (N_14853,N_8899,N_9075);
nor U14854 (N_14854,N_7683,N_7473);
xor U14855 (N_14855,N_11708,N_11160);
nand U14856 (N_14856,N_10753,N_11114);
and U14857 (N_14857,N_11856,N_9416);
or U14858 (N_14858,N_8876,N_8038);
nand U14859 (N_14859,N_7561,N_7374);
xor U14860 (N_14860,N_7551,N_6590);
nor U14861 (N_14861,N_10130,N_8831);
nand U14862 (N_14862,N_9357,N_7764);
or U14863 (N_14863,N_8448,N_10392);
nand U14864 (N_14864,N_11242,N_6724);
or U14865 (N_14865,N_8706,N_11661);
nand U14866 (N_14866,N_6721,N_9692);
nor U14867 (N_14867,N_8580,N_8759);
and U14868 (N_14868,N_10807,N_9019);
or U14869 (N_14869,N_9705,N_6488);
or U14870 (N_14870,N_10986,N_7408);
and U14871 (N_14871,N_7902,N_7056);
or U14872 (N_14872,N_9308,N_9895);
or U14873 (N_14873,N_7808,N_8194);
and U14874 (N_14874,N_10490,N_9226);
xor U14875 (N_14875,N_8950,N_11419);
xnor U14876 (N_14876,N_11535,N_6354);
or U14877 (N_14877,N_10389,N_11185);
or U14878 (N_14878,N_10549,N_8878);
nand U14879 (N_14879,N_10914,N_9612);
xnor U14880 (N_14880,N_10174,N_9198);
nand U14881 (N_14881,N_8049,N_10636);
and U14882 (N_14882,N_9215,N_11857);
or U14883 (N_14883,N_6427,N_9816);
or U14884 (N_14884,N_8187,N_11684);
xnor U14885 (N_14885,N_7327,N_11991);
nor U14886 (N_14886,N_10719,N_6430);
nand U14887 (N_14887,N_7108,N_11967);
xnor U14888 (N_14888,N_7635,N_10658);
and U14889 (N_14889,N_9130,N_9871);
nor U14890 (N_14890,N_8131,N_8551);
and U14891 (N_14891,N_10258,N_11579);
nand U14892 (N_14892,N_8435,N_11429);
or U14893 (N_14893,N_10219,N_7734);
and U14894 (N_14894,N_7532,N_6137);
xor U14895 (N_14895,N_6744,N_8790);
and U14896 (N_14896,N_7477,N_8101);
or U14897 (N_14897,N_9302,N_9651);
nand U14898 (N_14898,N_11785,N_10895);
or U14899 (N_14899,N_10370,N_6875);
nor U14900 (N_14900,N_7468,N_10261);
xnor U14901 (N_14901,N_6694,N_7065);
or U14902 (N_14902,N_9771,N_7283);
nor U14903 (N_14903,N_10859,N_7459);
nand U14904 (N_14904,N_9254,N_7781);
nor U14905 (N_14905,N_9301,N_6707);
nor U14906 (N_14906,N_7205,N_7392);
and U14907 (N_14907,N_11313,N_8616);
xor U14908 (N_14908,N_9746,N_8660);
nand U14909 (N_14909,N_8328,N_6044);
xor U14910 (N_14910,N_6278,N_6190);
nor U14911 (N_14911,N_9454,N_10910);
nor U14912 (N_14912,N_11095,N_9653);
xnor U14913 (N_14913,N_6069,N_11141);
nand U14914 (N_14914,N_9546,N_8637);
nand U14915 (N_14915,N_6459,N_10742);
or U14916 (N_14916,N_9753,N_6495);
nor U14917 (N_14917,N_7063,N_8365);
and U14918 (N_14918,N_10250,N_10372);
or U14919 (N_14919,N_7876,N_9386);
nor U14920 (N_14920,N_7846,N_7464);
nor U14921 (N_14921,N_7737,N_8589);
and U14922 (N_14922,N_6741,N_9760);
xnor U14923 (N_14923,N_8792,N_8031);
nand U14924 (N_14924,N_9291,N_6185);
or U14925 (N_14925,N_9757,N_6080);
or U14926 (N_14926,N_9801,N_8393);
or U14927 (N_14927,N_11941,N_11769);
xor U14928 (N_14928,N_11152,N_6807);
nand U14929 (N_14929,N_8417,N_10567);
or U14930 (N_14930,N_10814,N_11582);
nor U14931 (N_14931,N_6911,N_11309);
nand U14932 (N_14932,N_9204,N_7250);
xnor U14933 (N_14933,N_10993,N_10315);
xnor U14934 (N_14934,N_10171,N_11040);
nand U14935 (N_14935,N_9859,N_10538);
or U14936 (N_14936,N_8823,N_11347);
nand U14937 (N_14937,N_10544,N_6613);
or U14938 (N_14938,N_10754,N_8316);
or U14939 (N_14939,N_8005,N_7094);
xnor U14940 (N_14940,N_11570,N_7325);
or U14941 (N_14941,N_9966,N_6755);
nor U14942 (N_14942,N_9053,N_11375);
and U14943 (N_14943,N_6663,N_11093);
or U14944 (N_14944,N_6820,N_9309);
nand U14945 (N_14945,N_8098,N_9784);
xor U14946 (N_14946,N_6008,N_10764);
xor U14947 (N_14947,N_8281,N_6413);
and U14948 (N_14948,N_9891,N_8508);
nor U14949 (N_14949,N_7039,N_8259);
nand U14950 (N_14950,N_11259,N_8952);
nand U14951 (N_14951,N_6735,N_7497);
nor U14952 (N_14952,N_11803,N_8110);
xnor U14953 (N_14953,N_9238,N_6341);
and U14954 (N_14954,N_9900,N_6074);
nand U14955 (N_14955,N_11533,N_11946);
and U14956 (N_14956,N_9158,N_7710);
nor U14957 (N_14957,N_11554,N_6928);
xor U14958 (N_14958,N_9227,N_10663);
or U14959 (N_14959,N_8002,N_9591);
and U14960 (N_14960,N_7008,N_7937);
nand U14961 (N_14961,N_10903,N_6156);
nor U14962 (N_14962,N_7073,N_9724);
and U14963 (N_14963,N_8378,N_8476);
or U14964 (N_14964,N_6584,N_7674);
and U14965 (N_14965,N_10512,N_7371);
and U14966 (N_14966,N_8191,N_11171);
nand U14967 (N_14967,N_10188,N_10511);
nor U14968 (N_14968,N_8700,N_9563);
nor U14969 (N_14969,N_10679,N_6108);
and U14970 (N_14970,N_10166,N_8214);
nand U14971 (N_14971,N_6805,N_7015);
xnor U14972 (N_14972,N_7088,N_6439);
xor U14973 (N_14973,N_8769,N_8165);
xnor U14974 (N_14974,N_8929,N_9906);
nand U14975 (N_14975,N_6333,N_6213);
nor U14976 (N_14976,N_6286,N_9595);
nand U14977 (N_14977,N_6748,N_8321);
nor U14978 (N_14978,N_10883,N_7524);
nor U14979 (N_14979,N_7116,N_7137);
and U14980 (N_14980,N_6957,N_10180);
nor U14981 (N_14981,N_9699,N_11174);
nand U14982 (N_14982,N_11619,N_9524);
and U14983 (N_14983,N_9931,N_11389);
and U14984 (N_14984,N_7355,N_8896);
or U14985 (N_14985,N_9212,N_6422);
or U14986 (N_14986,N_6700,N_10368);
or U14987 (N_14987,N_8275,N_10387);
and U14988 (N_14988,N_7240,N_10761);
xor U14989 (N_14989,N_7324,N_10583);
nand U14990 (N_14990,N_6541,N_7376);
nand U14991 (N_14991,N_9685,N_11624);
nand U14992 (N_14992,N_7259,N_6711);
or U14993 (N_14993,N_10928,N_6414);
nand U14994 (N_14994,N_7037,N_10952);
nor U14995 (N_14995,N_10971,N_7928);
nand U14996 (N_14996,N_6891,N_7884);
or U14997 (N_14997,N_8174,N_11910);
xnor U14998 (N_14998,N_10038,N_7096);
nand U14999 (N_14999,N_11425,N_6144);
nand U15000 (N_15000,N_6896,N_6752);
and U15001 (N_15001,N_8618,N_11037);
or U15002 (N_15002,N_11398,N_11856);
or U15003 (N_15003,N_11643,N_11439);
xnor U15004 (N_15004,N_9145,N_7589);
nand U15005 (N_15005,N_7244,N_6288);
or U15006 (N_15006,N_6748,N_9175);
or U15007 (N_15007,N_6787,N_11315);
xnor U15008 (N_15008,N_6820,N_10811);
nand U15009 (N_15009,N_10929,N_10274);
nand U15010 (N_15010,N_9883,N_10513);
xor U15011 (N_15011,N_10186,N_8098);
and U15012 (N_15012,N_7721,N_9737);
and U15013 (N_15013,N_7535,N_11400);
nand U15014 (N_15014,N_7946,N_7181);
nor U15015 (N_15015,N_8633,N_9330);
xnor U15016 (N_15016,N_9964,N_9461);
and U15017 (N_15017,N_11032,N_8713);
nor U15018 (N_15018,N_9150,N_8359);
nor U15019 (N_15019,N_9400,N_11303);
nor U15020 (N_15020,N_10141,N_11818);
xnor U15021 (N_15021,N_11353,N_8422);
or U15022 (N_15022,N_10806,N_7591);
nor U15023 (N_15023,N_11056,N_8638);
and U15024 (N_15024,N_9313,N_8563);
or U15025 (N_15025,N_10999,N_9962);
nand U15026 (N_15026,N_10716,N_9878);
nor U15027 (N_15027,N_9169,N_11036);
nor U15028 (N_15028,N_11113,N_11856);
xnor U15029 (N_15029,N_8788,N_8944);
nor U15030 (N_15030,N_6155,N_6158);
nand U15031 (N_15031,N_8856,N_8219);
nand U15032 (N_15032,N_7779,N_11505);
or U15033 (N_15033,N_6510,N_10783);
xor U15034 (N_15034,N_8497,N_11967);
nand U15035 (N_15035,N_11043,N_6342);
xor U15036 (N_15036,N_9827,N_6817);
nand U15037 (N_15037,N_8081,N_9778);
nand U15038 (N_15038,N_11621,N_10518);
and U15039 (N_15039,N_8768,N_7410);
and U15040 (N_15040,N_10306,N_9885);
nor U15041 (N_15041,N_7547,N_7718);
or U15042 (N_15042,N_6606,N_9945);
or U15043 (N_15043,N_8326,N_9633);
nor U15044 (N_15044,N_11189,N_11216);
nand U15045 (N_15045,N_9583,N_6910);
xnor U15046 (N_15046,N_6726,N_11426);
nor U15047 (N_15047,N_10564,N_11091);
xnor U15048 (N_15048,N_10973,N_9265);
nor U15049 (N_15049,N_8075,N_9326);
xor U15050 (N_15050,N_10464,N_9634);
or U15051 (N_15051,N_6901,N_10942);
or U15052 (N_15052,N_8156,N_6976);
nor U15053 (N_15053,N_6387,N_6149);
xnor U15054 (N_15054,N_6979,N_10625);
or U15055 (N_15055,N_11220,N_6688);
xnor U15056 (N_15056,N_8458,N_7678);
xnor U15057 (N_15057,N_6397,N_6040);
xnor U15058 (N_15058,N_10233,N_8066);
nor U15059 (N_15059,N_6402,N_9198);
or U15060 (N_15060,N_8585,N_11992);
xnor U15061 (N_15061,N_7731,N_6075);
or U15062 (N_15062,N_10414,N_8044);
and U15063 (N_15063,N_6899,N_8955);
or U15064 (N_15064,N_7943,N_10885);
or U15065 (N_15065,N_10156,N_8874);
and U15066 (N_15066,N_6985,N_8544);
or U15067 (N_15067,N_9651,N_6346);
nand U15068 (N_15068,N_11212,N_11054);
nand U15069 (N_15069,N_7268,N_11418);
and U15070 (N_15070,N_7261,N_8449);
nand U15071 (N_15071,N_10325,N_7012);
xor U15072 (N_15072,N_11942,N_6962);
and U15073 (N_15073,N_11836,N_11377);
or U15074 (N_15074,N_7034,N_7888);
and U15075 (N_15075,N_10176,N_6502);
and U15076 (N_15076,N_7488,N_10861);
xnor U15077 (N_15077,N_8207,N_6227);
nand U15078 (N_15078,N_10123,N_9157);
and U15079 (N_15079,N_10565,N_9046);
and U15080 (N_15080,N_6165,N_11629);
xor U15081 (N_15081,N_9114,N_10330);
or U15082 (N_15082,N_11526,N_9838);
or U15083 (N_15083,N_7723,N_7262);
xor U15084 (N_15084,N_7728,N_7280);
nor U15085 (N_15085,N_11481,N_8725);
nor U15086 (N_15086,N_6555,N_11048);
and U15087 (N_15087,N_11864,N_10778);
nand U15088 (N_15088,N_11856,N_6939);
or U15089 (N_15089,N_11897,N_7584);
xnor U15090 (N_15090,N_7993,N_11917);
nand U15091 (N_15091,N_11632,N_11331);
and U15092 (N_15092,N_8521,N_9461);
nand U15093 (N_15093,N_8348,N_11453);
or U15094 (N_15094,N_9785,N_8655);
xnor U15095 (N_15095,N_11445,N_11750);
nand U15096 (N_15096,N_8782,N_8638);
nand U15097 (N_15097,N_11230,N_10213);
and U15098 (N_15098,N_8503,N_11626);
nor U15099 (N_15099,N_7281,N_11404);
and U15100 (N_15100,N_11537,N_7459);
or U15101 (N_15101,N_9267,N_8207);
and U15102 (N_15102,N_7095,N_7176);
xor U15103 (N_15103,N_6003,N_11668);
xor U15104 (N_15104,N_9048,N_7025);
nor U15105 (N_15105,N_8614,N_9957);
nand U15106 (N_15106,N_7016,N_10851);
nor U15107 (N_15107,N_8384,N_10936);
and U15108 (N_15108,N_6081,N_11306);
xnor U15109 (N_15109,N_10833,N_10478);
nand U15110 (N_15110,N_6826,N_11285);
or U15111 (N_15111,N_11695,N_6421);
nor U15112 (N_15112,N_6750,N_10036);
and U15113 (N_15113,N_10771,N_8601);
or U15114 (N_15114,N_6012,N_11692);
and U15115 (N_15115,N_11911,N_8584);
nor U15116 (N_15116,N_11837,N_10634);
nor U15117 (N_15117,N_10926,N_10729);
or U15118 (N_15118,N_6443,N_10522);
nor U15119 (N_15119,N_6176,N_8600);
and U15120 (N_15120,N_9718,N_10989);
xnor U15121 (N_15121,N_11308,N_6953);
nand U15122 (N_15122,N_9926,N_8042);
or U15123 (N_15123,N_10134,N_7936);
nor U15124 (N_15124,N_6261,N_7496);
nand U15125 (N_15125,N_7242,N_11507);
nor U15126 (N_15126,N_10663,N_11406);
or U15127 (N_15127,N_10141,N_11642);
xnor U15128 (N_15128,N_9909,N_7903);
xor U15129 (N_15129,N_7397,N_11767);
or U15130 (N_15130,N_10798,N_10212);
and U15131 (N_15131,N_8419,N_6000);
xor U15132 (N_15132,N_11587,N_10372);
nand U15133 (N_15133,N_6776,N_9951);
xor U15134 (N_15134,N_11448,N_10833);
nor U15135 (N_15135,N_6333,N_11431);
or U15136 (N_15136,N_9810,N_8633);
nand U15137 (N_15137,N_9717,N_10697);
xor U15138 (N_15138,N_6124,N_11138);
xnor U15139 (N_15139,N_10292,N_7582);
nor U15140 (N_15140,N_11722,N_9572);
nand U15141 (N_15141,N_11464,N_8394);
xnor U15142 (N_15142,N_10785,N_10220);
nand U15143 (N_15143,N_8476,N_8143);
xor U15144 (N_15144,N_11955,N_6528);
xor U15145 (N_15145,N_7543,N_7162);
nand U15146 (N_15146,N_11609,N_11960);
or U15147 (N_15147,N_11809,N_8387);
and U15148 (N_15148,N_10815,N_8948);
or U15149 (N_15149,N_9979,N_11024);
nand U15150 (N_15150,N_8325,N_9847);
nor U15151 (N_15151,N_8385,N_8889);
xnor U15152 (N_15152,N_7316,N_11082);
and U15153 (N_15153,N_11135,N_10825);
and U15154 (N_15154,N_11518,N_10779);
and U15155 (N_15155,N_7816,N_10657);
and U15156 (N_15156,N_11705,N_9109);
nor U15157 (N_15157,N_10410,N_6909);
nand U15158 (N_15158,N_7807,N_10167);
xnor U15159 (N_15159,N_10514,N_9401);
nor U15160 (N_15160,N_11082,N_9156);
or U15161 (N_15161,N_8573,N_8922);
nor U15162 (N_15162,N_9732,N_8801);
nor U15163 (N_15163,N_6388,N_6245);
nor U15164 (N_15164,N_10901,N_10113);
and U15165 (N_15165,N_9896,N_8474);
xnor U15166 (N_15166,N_10880,N_9740);
and U15167 (N_15167,N_7328,N_10340);
nor U15168 (N_15168,N_9487,N_8628);
nand U15169 (N_15169,N_7052,N_8348);
nand U15170 (N_15170,N_11417,N_8642);
nand U15171 (N_15171,N_8227,N_6510);
or U15172 (N_15172,N_8629,N_8884);
or U15173 (N_15173,N_9331,N_10399);
or U15174 (N_15174,N_9560,N_10118);
or U15175 (N_15175,N_11682,N_6974);
nand U15176 (N_15176,N_8876,N_6534);
or U15177 (N_15177,N_10184,N_11782);
nand U15178 (N_15178,N_7425,N_6549);
nand U15179 (N_15179,N_11817,N_10555);
nand U15180 (N_15180,N_7147,N_11190);
xor U15181 (N_15181,N_9366,N_8150);
and U15182 (N_15182,N_9584,N_6229);
and U15183 (N_15183,N_9527,N_11550);
nor U15184 (N_15184,N_8337,N_10654);
or U15185 (N_15185,N_6459,N_9698);
nor U15186 (N_15186,N_6196,N_11746);
nand U15187 (N_15187,N_10318,N_6971);
and U15188 (N_15188,N_11595,N_7798);
or U15189 (N_15189,N_10969,N_6677);
or U15190 (N_15190,N_10627,N_6469);
or U15191 (N_15191,N_10656,N_9416);
nor U15192 (N_15192,N_11598,N_8284);
nor U15193 (N_15193,N_8646,N_11876);
nor U15194 (N_15194,N_9722,N_11633);
nor U15195 (N_15195,N_9520,N_6575);
xnor U15196 (N_15196,N_9549,N_6011);
nand U15197 (N_15197,N_10044,N_8178);
nand U15198 (N_15198,N_7560,N_11545);
nor U15199 (N_15199,N_8526,N_11384);
nor U15200 (N_15200,N_8490,N_11198);
xnor U15201 (N_15201,N_6291,N_7326);
nand U15202 (N_15202,N_7987,N_8704);
and U15203 (N_15203,N_7644,N_8630);
nor U15204 (N_15204,N_6950,N_6681);
nor U15205 (N_15205,N_7216,N_10080);
or U15206 (N_15206,N_9012,N_11291);
xor U15207 (N_15207,N_10465,N_6293);
or U15208 (N_15208,N_8651,N_7038);
nor U15209 (N_15209,N_11696,N_7338);
or U15210 (N_15210,N_7262,N_8073);
and U15211 (N_15211,N_7150,N_11003);
xor U15212 (N_15212,N_8372,N_10527);
nand U15213 (N_15213,N_6037,N_11097);
xnor U15214 (N_15214,N_11682,N_10617);
or U15215 (N_15215,N_8592,N_7889);
nand U15216 (N_15216,N_7545,N_7147);
nor U15217 (N_15217,N_7447,N_6436);
and U15218 (N_15218,N_7282,N_11191);
nand U15219 (N_15219,N_11437,N_11883);
or U15220 (N_15220,N_8473,N_8823);
nor U15221 (N_15221,N_8903,N_9880);
xor U15222 (N_15222,N_9053,N_8328);
nand U15223 (N_15223,N_11207,N_7666);
nand U15224 (N_15224,N_10319,N_7704);
or U15225 (N_15225,N_7627,N_8195);
xor U15226 (N_15226,N_9232,N_11003);
nand U15227 (N_15227,N_6604,N_11880);
nor U15228 (N_15228,N_8248,N_9068);
xor U15229 (N_15229,N_9114,N_9315);
nand U15230 (N_15230,N_11862,N_6009);
xnor U15231 (N_15231,N_7854,N_11190);
xnor U15232 (N_15232,N_9452,N_10902);
nor U15233 (N_15233,N_6398,N_11959);
xnor U15234 (N_15234,N_6592,N_6334);
nor U15235 (N_15235,N_9517,N_9020);
xnor U15236 (N_15236,N_8086,N_7842);
or U15237 (N_15237,N_7116,N_10944);
and U15238 (N_15238,N_11102,N_9202);
nand U15239 (N_15239,N_6488,N_9134);
nor U15240 (N_15240,N_9274,N_11513);
nand U15241 (N_15241,N_11451,N_8707);
nand U15242 (N_15242,N_9291,N_7256);
xor U15243 (N_15243,N_6773,N_9069);
nor U15244 (N_15244,N_9408,N_10550);
nor U15245 (N_15245,N_8221,N_11157);
nor U15246 (N_15246,N_7683,N_8922);
xnor U15247 (N_15247,N_9831,N_6554);
xor U15248 (N_15248,N_8138,N_9500);
nor U15249 (N_15249,N_10373,N_7825);
nor U15250 (N_15250,N_7231,N_9450);
and U15251 (N_15251,N_11283,N_11159);
nand U15252 (N_15252,N_8965,N_11478);
or U15253 (N_15253,N_8476,N_8177);
nand U15254 (N_15254,N_10868,N_11726);
and U15255 (N_15255,N_10384,N_7719);
and U15256 (N_15256,N_10666,N_11400);
nand U15257 (N_15257,N_6762,N_9292);
nand U15258 (N_15258,N_7857,N_9037);
and U15259 (N_15259,N_7082,N_8102);
and U15260 (N_15260,N_9236,N_6447);
or U15261 (N_15261,N_6198,N_10451);
and U15262 (N_15262,N_11376,N_11945);
xnor U15263 (N_15263,N_7099,N_6552);
and U15264 (N_15264,N_6300,N_7374);
nand U15265 (N_15265,N_6787,N_9113);
or U15266 (N_15266,N_6318,N_11029);
nor U15267 (N_15267,N_10911,N_11132);
and U15268 (N_15268,N_10016,N_10053);
nor U15269 (N_15269,N_9530,N_9123);
nor U15270 (N_15270,N_8318,N_8957);
or U15271 (N_15271,N_7952,N_11762);
or U15272 (N_15272,N_8474,N_6033);
or U15273 (N_15273,N_9199,N_7452);
or U15274 (N_15274,N_8197,N_6425);
or U15275 (N_15275,N_9498,N_6921);
xnor U15276 (N_15276,N_7215,N_10547);
nand U15277 (N_15277,N_9549,N_8553);
nor U15278 (N_15278,N_9017,N_10591);
xor U15279 (N_15279,N_8661,N_9949);
or U15280 (N_15280,N_6574,N_9023);
xor U15281 (N_15281,N_7227,N_10429);
and U15282 (N_15282,N_9061,N_7557);
nand U15283 (N_15283,N_11705,N_7161);
nand U15284 (N_15284,N_8958,N_11291);
and U15285 (N_15285,N_11782,N_8767);
and U15286 (N_15286,N_9687,N_10445);
nor U15287 (N_15287,N_7446,N_8232);
and U15288 (N_15288,N_10761,N_9333);
nand U15289 (N_15289,N_6649,N_7955);
and U15290 (N_15290,N_9711,N_8474);
or U15291 (N_15291,N_8284,N_9267);
or U15292 (N_15292,N_6593,N_10785);
nor U15293 (N_15293,N_8840,N_10883);
nor U15294 (N_15294,N_8300,N_6815);
xnor U15295 (N_15295,N_8666,N_8064);
or U15296 (N_15296,N_11759,N_9885);
and U15297 (N_15297,N_8050,N_11953);
nor U15298 (N_15298,N_7213,N_11404);
and U15299 (N_15299,N_11347,N_8231);
and U15300 (N_15300,N_9954,N_10715);
or U15301 (N_15301,N_10323,N_6194);
xnor U15302 (N_15302,N_8984,N_11727);
or U15303 (N_15303,N_8532,N_7901);
nand U15304 (N_15304,N_6063,N_9742);
and U15305 (N_15305,N_9866,N_6024);
nand U15306 (N_15306,N_11835,N_7341);
or U15307 (N_15307,N_11552,N_6462);
nor U15308 (N_15308,N_10534,N_6723);
nor U15309 (N_15309,N_8665,N_7354);
or U15310 (N_15310,N_8004,N_8385);
xnor U15311 (N_15311,N_9015,N_8553);
xor U15312 (N_15312,N_10460,N_11046);
nor U15313 (N_15313,N_11044,N_7600);
or U15314 (N_15314,N_7989,N_7591);
nand U15315 (N_15315,N_8456,N_11406);
nor U15316 (N_15316,N_11442,N_11485);
nor U15317 (N_15317,N_6721,N_8355);
or U15318 (N_15318,N_9649,N_8791);
xnor U15319 (N_15319,N_8310,N_9930);
xnor U15320 (N_15320,N_10149,N_9662);
xor U15321 (N_15321,N_10042,N_8070);
nand U15322 (N_15322,N_7204,N_8620);
nand U15323 (N_15323,N_6319,N_6893);
nand U15324 (N_15324,N_9319,N_10389);
or U15325 (N_15325,N_10914,N_7369);
and U15326 (N_15326,N_9710,N_11841);
and U15327 (N_15327,N_11775,N_6366);
xor U15328 (N_15328,N_8861,N_6838);
nand U15329 (N_15329,N_7893,N_10008);
xnor U15330 (N_15330,N_7730,N_7289);
nand U15331 (N_15331,N_11771,N_11993);
nand U15332 (N_15332,N_7014,N_8330);
xor U15333 (N_15333,N_6587,N_9143);
and U15334 (N_15334,N_9131,N_9386);
nand U15335 (N_15335,N_8492,N_10390);
xnor U15336 (N_15336,N_10530,N_10022);
nor U15337 (N_15337,N_6560,N_7560);
nor U15338 (N_15338,N_7368,N_8850);
nor U15339 (N_15339,N_7627,N_7753);
or U15340 (N_15340,N_11394,N_10899);
nor U15341 (N_15341,N_6743,N_10960);
nor U15342 (N_15342,N_9605,N_11238);
nand U15343 (N_15343,N_10118,N_8493);
nor U15344 (N_15344,N_7017,N_7891);
or U15345 (N_15345,N_6980,N_10150);
nor U15346 (N_15346,N_8039,N_6890);
xor U15347 (N_15347,N_10511,N_9859);
nand U15348 (N_15348,N_7114,N_7686);
nor U15349 (N_15349,N_9058,N_9623);
xor U15350 (N_15350,N_7091,N_11425);
or U15351 (N_15351,N_7178,N_7122);
nor U15352 (N_15352,N_7122,N_10282);
nand U15353 (N_15353,N_8809,N_6765);
nor U15354 (N_15354,N_10750,N_11266);
nor U15355 (N_15355,N_9664,N_6788);
or U15356 (N_15356,N_9860,N_7600);
nand U15357 (N_15357,N_11554,N_6786);
and U15358 (N_15358,N_11252,N_10020);
or U15359 (N_15359,N_11900,N_10232);
or U15360 (N_15360,N_11909,N_6010);
nor U15361 (N_15361,N_10155,N_11521);
nor U15362 (N_15362,N_6299,N_9704);
nand U15363 (N_15363,N_7392,N_11823);
or U15364 (N_15364,N_6126,N_8719);
nor U15365 (N_15365,N_7820,N_6988);
or U15366 (N_15366,N_6197,N_7259);
nor U15367 (N_15367,N_7749,N_10514);
or U15368 (N_15368,N_8596,N_10951);
or U15369 (N_15369,N_8691,N_8853);
nor U15370 (N_15370,N_6972,N_8478);
nor U15371 (N_15371,N_6103,N_9246);
and U15372 (N_15372,N_8592,N_9787);
and U15373 (N_15373,N_11423,N_8874);
or U15374 (N_15374,N_7302,N_10383);
and U15375 (N_15375,N_6953,N_10217);
nand U15376 (N_15376,N_7342,N_11468);
xor U15377 (N_15377,N_9770,N_7845);
nor U15378 (N_15378,N_8039,N_9406);
nor U15379 (N_15379,N_7153,N_10655);
and U15380 (N_15380,N_7636,N_7694);
xnor U15381 (N_15381,N_9013,N_6756);
xor U15382 (N_15382,N_11295,N_7865);
nor U15383 (N_15383,N_8122,N_10917);
nor U15384 (N_15384,N_11116,N_11011);
and U15385 (N_15385,N_7913,N_6529);
nor U15386 (N_15386,N_9513,N_9372);
nand U15387 (N_15387,N_6460,N_10524);
xnor U15388 (N_15388,N_8743,N_7390);
nor U15389 (N_15389,N_6502,N_11926);
or U15390 (N_15390,N_10207,N_8922);
and U15391 (N_15391,N_10798,N_7722);
nand U15392 (N_15392,N_10688,N_11659);
or U15393 (N_15393,N_11332,N_10274);
xor U15394 (N_15394,N_8792,N_8193);
and U15395 (N_15395,N_8733,N_9143);
and U15396 (N_15396,N_10376,N_11590);
nor U15397 (N_15397,N_8732,N_10520);
nor U15398 (N_15398,N_10160,N_11220);
or U15399 (N_15399,N_11638,N_10492);
nand U15400 (N_15400,N_6312,N_8150);
xnor U15401 (N_15401,N_7752,N_9331);
nand U15402 (N_15402,N_6349,N_6594);
xor U15403 (N_15403,N_11842,N_7182);
and U15404 (N_15404,N_7472,N_11298);
or U15405 (N_15405,N_7678,N_9691);
nand U15406 (N_15406,N_8856,N_6869);
nor U15407 (N_15407,N_9921,N_6078);
xor U15408 (N_15408,N_8767,N_11781);
nor U15409 (N_15409,N_9577,N_10041);
and U15410 (N_15410,N_9862,N_7730);
nor U15411 (N_15411,N_10698,N_8232);
or U15412 (N_15412,N_6634,N_8477);
nor U15413 (N_15413,N_6849,N_9028);
nor U15414 (N_15414,N_9535,N_11515);
xor U15415 (N_15415,N_10494,N_11661);
nor U15416 (N_15416,N_6807,N_7981);
nand U15417 (N_15417,N_11029,N_10174);
or U15418 (N_15418,N_10377,N_11807);
xor U15419 (N_15419,N_11339,N_6362);
or U15420 (N_15420,N_8307,N_11281);
or U15421 (N_15421,N_6268,N_9664);
and U15422 (N_15422,N_8033,N_9059);
and U15423 (N_15423,N_6157,N_11133);
or U15424 (N_15424,N_8404,N_9931);
nor U15425 (N_15425,N_9657,N_9385);
and U15426 (N_15426,N_9302,N_10340);
or U15427 (N_15427,N_11412,N_11715);
or U15428 (N_15428,N_7751,N_7694);
nor U15429 (N_15429,N_9452,N_7952);
nor U15430 (N_15430,N_9401,N_8430);
nand U15431 (N_15431,N_9268,N_11631);
nor U15432 (N_15432,N_6854,N_7996);
nand U15433 (N_15433,N_6994,N_11994);
or U15434 (N_15434,N_8848,N_6590);
nand U15435 (N_15435,N_6795,N_7327);
and U15436 (N_15436,N_7953,N_6658);
or U15437 (N_15437,N_9152,N_6794);
and U15438 (N_15438,N_6248,N_9304);
or U15439 (N_15439,N_9001,N_9245);
xor U15440 (N_15440,N_11623,N_6158);
and U15441 (N_15441,N_8789,N_11155);
and U15442 (N_15442,N_9110,N_8986);
nand U15443 (N_15443,N_10185,N_11434);
and U15444 (N_15444,N_6534,N_8367);
nor U15445 (N_15445,N_11602,N_10905);
or U15446 (N_15446,N_7152,N_6980);
nor U15447 (N_15447,N_10236,N_11872);
nand U15448 (N_15448,N_8888,N_6216);
xor U15449 (N_15449,N_6643,N_6554);
xnor U15450 (N_15450,N_6717,N_11012);
nand U15451 (N_15451,N_8959,N_10890);
xnor U15452 (N_15452,N_6591,N_7712);
or U15453 (N_15453,N_8353,N_8730);
or U15454 (N_15454,N_10038,N_6575);
nand U15455 (N_15455,N_8512,N_9146);
or U15456 (N_15456,N_11812,N_8009);
xor U15457 (N_15457,N_8970,N_11343);
and U15458 (N_15458,N_6533,N_8275);
and U15459 (N_15459,N_6330,N_6831);
nand U15460 (N_15460,N_11335,N_7972);
and U15461 (N_15461,N_10295,N_7243);
and U15462 (N_15462,N_8777,N_11874);
xor U15463 (N_15463,N_7389,N_6337);
and U15464 (N_15464,N_8164,N_11317);
nor U15465 (N_15465,N_6647,N_9487);
nor U15466 (N_15466,N_6177,N_10946);
nor U15467 (N_15467,N_6713,N_6032);
xnor U15468 (N_15468,N_7194,N_7114);
xnor U15469 (N_15469,N_6576,N_9087);
xor U15470 (N_15470,N_9814,N_10919);
nor U15471 (N_15471,N_8858,N_8941);
nor U15472 (N_15472,N_10055,N_6861);
xor U15473 (N_15473,N_10918,N_8093);
and U15474 (N_15474,N_8297,N_9873);
or U15475 (N_15475,N_6579,N_11005);
xnor U15476 (N_15476,N_7827,N_8588);
xnor U15477 (N_15477,N_8845,N_11176);
or U15478 (N_15478,N_6386,N_11978);
xor U15479 (N_15479,N_9786,N_11241);
and U15480 (N_15480,N_9115,N_9836);
or U15481 (N_15481,N_6954,N_7682);
or U15482 (N_15482,N_8424,N_9328);
nand U15483 (N_15483,N_10765,N_7028);
xnor U15484 (N_15484,N_8994,N_10896);
nand U15485 (N_15485,N_9540,N_8249);
nand U15486 (N_15486,N_9006,N_10971);
nand U15487 (N_15487,N_6140,N_8507);
nand U15488 (N_15488,N_8759,N_11628);
or U15489 (N_15489,N_9244,N_11586);
or U15490 (N_15490,N_7824,N_8298);
or U15491 (N_15491,N_10573,N_10525);
nand U15492 (N_15492,N_8266,N_9845);
or U15493 (N_15493,N_10771,N_10734);
and U15494 (N_15494,N_11232,N_10813);
nand U15495 (N_15495,N_10055,N_10862);
xnor U15496 (N_15496,N_8167,N_10694);
or U15497 (N_15497,N_11252,N_11840);
or U15498 (N_15498,N_6786,N_9430);
nor U15499 (N_15499,N_10916,N_7291);
or U15500 (N_15500,N_9394,N_6262);
nor U15501 (N_15501,N_7541,N_7296);
nand U15502 (N_15502,N_11266,N_6562);
xnor U15503 (N_15503,N_7727,N_10046);
nor U15504 (N_15504,N_6617,N_10720);
nor U15505 (N_15505,N_10039,N_11842);
or U15506 (N_15506,N_6068,N_11577);
and U15507 (N_15507,N_7478,N_11858);
nor U15508 (N_15508,N_9266,N_9672);
or U15509 (N_15509,N_7805,N_11837);
or U15510 (N_15510,N_11469,N_10804);
or U15511 (N_15511,N_11081,N_11033);
xor U15512 (N_15512,N_10440,N_11044);
xor U15513 (N_15513,N_10504,N_6248);
and U15514 (N_15514,N_9873,N_7494);
xor U15515 (N_15515,N_6198,N_8823);
xor U15516 (N_15516,N_7900,N_8525);
and U15517 (N_15517,N_10972,N_7467);
or U15518 (N_15518,N_10734,N_7132);
or U15519 (N_15519,N_7535,N_11569);
or U15520 (N_15520,N_11577,N_7991);
and U15521 (N_15521,N_9260,N_9342);
nor U15522 (N_15522,N_7484,N_7107);
xnor U15523 (N_15523,N_9563,N_6224);
xor U15524 (N_15524,N_8841,N_6356);
and U15525 (N_15525,N_6456,N_7258);
nand U15526 (N_15526,N_11928,N_8490);
and U15527 (N_15527,N_8327,N_7241);
xor U15528 (N_15528,N_6535,N_9653);
or U15529 (N_15529,N_7600,N_10281);
nor U15530 (N_15530,N_11612,N_11332);
xor U15531 (N_15531,N_8032,N_9375);
nor U15532 (N_15532,N_10374,N_11607);
nor U15533 (N_15533,N_11032,N_8683);
or U15534 (N_15534,N_6740,N_8850);
or U15535 (N_15535,N_7006,N_11343);
nor U15536 (N_15536,N_11752,N_8742);
nand U15537 (N_15537,N_6858,N_7615);
nor U15538 (N_15538,N_8276,N_8049);
nor U15539 (N_15539,N_10420,N_6285);
and U15540 (N_15540,N_10707,N_10191);
nand U15541 (N_15541,N_11875,N_7994);
or U15542 (N_15542,N_9755,N_11887);
or U15543 (N_15543,N_8500,N_10942);
or U15544 (N_15544,N_11912,N_8654);
and U15545 (N_15545,N_9171,N_6724);
nand U15546 (N_15546,N_11604,N_11082);
xor U15547 (N_15547,N_6881,N_9237);
and U15548 (N_15548,N_9748,N_8212);
or U15549 (N_15549,N_7098,N_10227);
nor U15550 (N_15550,N_10976,N_6425);
xor U15551 (N_15551,N_11259,N_10475);
xnor U15552 (N_15552,N_10092,N_11900);
xor U15553 (N_15553,N_10758,N_9525);
xor U15554 (N_15554,N_6464,N_11653);
nand U15555 (N_15555,N_10565,N_10327);
or U15556 (N_15556,N_8753,N_6637);
nand U15557 (N_15557,N_11647,N_11346);
nand U15558 (N_15558,N_9981,N_9405);
or U15559 (N_15559,N_6020,N_8202);
xor U15560 (N_15560,N_8237,N_8794);
and U15561 (N_15561,N_6303,N_7938);
nor U15562 (N_15562,N_11524,N_10861);
or U15563 (N_15563,N_9133,N_10456);
nor U15564 (N_15564,N_6663,N_9276);
and U15565 (N_15565,N_11928,N_6264);
nor U15566 (N_15566,N_10790,N_9680);
or U15567 (N_15567,N_9224,N_8458);
or U15568 (N_15568,N_11564,N_7247);
or U15569 (N_15569,N_6672,N_7595);
xnor U15570 (N_15570,N_11984,N_8104);
or U15571 (N_15571,N_6329,N_11417);
or U15572 (N_15572,N_9896,N_9302);
nand U15573 (N_15573,N_6380,N_9169);
xnor U15574 (N_15574,N_8052,N_6608);
nor U15575 (N_15575,N_11108,N_6138);
or U15576 (N_15576,N_10111,N_9988);
nor U15577 (N_15577,N_10417,N_11956);
nand U15578 (N_15578,N_6121,N_7705);
xnor U15579 (N_15579,N_9728,N_10698);
or U15580 (N_15580,N_8291,N_8411);
nand U15581 (N_15581,N_8265,N_6126);
or U15582 (N_15582,N_6132,N_11167);
or U15583 (N_15583,N_9531,N_11228);
and U15584 (N_15584,N_7780,N_7947);
nor U15585 (N_15585,N_6337,N_10934);
or U15586 (N_15586,N_7920,N_7505);
or U15587 (N_15587,N_8114,N_10945);
nor U15588 (N_15588,N_11347,N_11600);
nor U15589 (N_15589,N_9909,N_11501);
xor U15590 (N_15590,N_6337,N_10268);
and U15591 (N_15591,N_8640,N_7786);
nor U15592 (N_15592,N_9001,N_9020);
and U15593 (N_15593,N_7922,N_7645);
xor U15594 (N_15594,N_8479,N_8829);
nand U15595 (N_15595,N_8294,N_7392);
nand U15596 (N_15596,N_10553,N_9240);
nor U15597 (N_15597,N_11313,N_9786);
nand U15598 (N_15598,N_9029,N_6986);
and U15599 (N_15599,N_11831,N_8119);
nand U15600 (N_15600,N_9297,N_6908);
and U15601 (N_15601,N_11363,N_6144);
xnor U15602 (N_15602,N_9399,N_6095);
and U15603 (N_15603,N_8458,N_8767);
nand U15604 (N_15604,N_11542,N_7911);
xnor U15605 (N_15605,N_11184,N_10191);
and U15606 (N_15606,N_10663,N_8093);
nor U15607 (N_15607,N_6912,N_7138);
nor U15608 (N_15608,N_8548,N_10761);
and U15609 (N_15609,N_11935,N_10670);
xnor U15610 (N_15610,N_10484,N_10334);
or U15611 (N_15611,N_6697,N_7915);
nor U15612 (N_15612,N_11030,N_6574);
and U15613 (N_15613,N_10387,N_9403);
or U15614 (N_15614,N_7487,N_7580);
and U15615 (N_15615,N_11278,N_7866);
nand U15616 (N_15616,N_10948,N_7457);
or U15617 (N_15617,N_10050,N_11481);
xnor U15618 (N_15618,N_7267,N_9195);
and U15619 (N_15619,N_8094,N_8788);
nand U15620 (N_15620,N_8945,N_10458);
nand U15621 (N_15621,N_9674,N_8939);
nand U15622 (N_15622,N_9802,N_7897);
nand U15623 (N_15623,N_11300,N_6214);
or U15624 (N_15624,N_6624,N_6420);
nand U15625 (N_15625,N_7237,N_9748);
or U15626 (N_15626,N_9572,N_10046);
or U15627 (N_15627,N_9539,N_10293);
xor U15628 (N_15628,N_6712,N_10811);
nand U15629 (N_15629,N_9514,N_7694);
and U15630 (N_15630,N_7938,N_9484);
nand U15631 (N_15631,N_9069,N_6870);
nand U15632 (N_15632,N_7973,N_8089);
nor U15633 (N_15633,N_7626,N_7028);
nand U15634 (N_15634,N_8171,N_10329);
and U15635 (N_15635,N_9565,N_11732);
and U15636 (N_15636,N_7365,N_7190);
nand U15637 (N_15637,N_9979,N_10583);
nor U15638 (N_15638,N_7142,N_11106);
or U15639 (N_15639,N_9635,N_8497);
and U15640 (N_15640,N_7458,N_11195);
nand U15641 (N_15641,N_9839,N_7584);
and U15642 (N_15642,N_11418,N_11740);
nand U15643 (N_15643,N_6848,N_9512);
xor U15644 (N_15644,N_11583,N_11179);
xor U15645 (N_15645,N_8372,N_9835);
nor U15646 (N_15646,N_10488,N_9516);
nor U15647 (N_15647,N_8003,N_7544);
nand U15648 (N_15648,N_9465,N_6219);
nor U15649 (N_15649,N_7441,N_10817);
nor U15650 (N_15650,N_9627,N_9964);
and U15651 (N_15651,N_10217,N_9739);
and U15652 (N_15652,N_10935,N_10716);
or U15653 (N_15653,N_10999,N_9629);
nor U15654 (N_15654,N_9339,N_6593);
and U15655 (N_15655,N_8483,N_6028);
xnor U15656 (N_15656,N_9386,N_7235);
nor U15657 (N_15657,N_7598,N_10918);
and U15658 (N_15658,N_10329,N_9470);
nand U15659 (N_15659,N_7290,N_8056);
nand U15660 (N_15660,N_8100,N_6835);
nand U15661 (N_15661,N_9244,N_6695);
or U15662 (N_15662,N_11426,N_6719);
nand U15663 (N_15663,N_7558,N_10031);
nor U15664 (N_15664,N_8641,N_6105);
and U15665 (N_15665,N_9015,N_9208);
nor U15666 (N_15666,N_9301,N_7556);
nor U15667 (N_15667,N_8557,N_6090);
and U15668 (N_15668,N_9029,N_10359);
and U15669 (N_15669,N_6934,N_7143);
and U15670 (N_15670,N_6719,N_8403);
xnor U15671 (N_15671,N_7685,N_8185);
and U15672 (N_15672,N_11470,N_8132);
xor U15673 (N_15673,N_9775,N_11288);
or U15674 (N_15674,N_10048,N_9611);
or U15675 (N_15675,N_11512,N_9408);
and U15676 (N_15676,N_6365,N_7175);
or U15677 (N_15677,N_10929,N_11783);
nand U15678 (N_15678,N_10987,N_7112);
nor U15679 (N_15679,N_10302,N_6500);
nand U15680 (N_15680,N_9759,N_8165);
nor U15681 (N_15681,N_11957,N_6398);
or U15682 (N_15682,N_6532,N_11537);
nor U15683 (N_15683,N_9685,N_6297);
xnor U15684 (N_15684,N_10639,N_7284);
nand U15685 (N_15685,N_6358,N_9781);
nor U15686 (N_15686,N_10204,N_10015);
nor U15687 (N_15687,N_7544,N_9459);
nand U15688 (N_15688,N_7289,N_9216);
and U15689 (N_15689,N_6321,N_11832);
and U15690 (N_15690,N_10769,N_8823);
or U15691 (N_15691,N_6340,N_11621);
nand U15692 (N_15692,N_11991,N_9281);
nor U15693 (N_15693,N_9957,N_9126);
nand U15694 (N_15694,N_8335,N_7618);
and U15695 (N_15695,N_7452,N_9591);
and U15696 (N_15696,N_9030,N_7676);
nand U15697 (N_15697,N_8687,N_7074);
nand U15698 (N_15698,N_11071,N_9917);
xnor U15699 (N_15699,N_6686,N_11935);
nor U15700 (N_15700,N_7498,N_8095);
or U15701 (N_15701,N_7342,N_8681);
xor U15702 (N_15702,N_10452,N_10803);
xor U15703 (N_15703,N_9400,N_9997);
nand U15704 (N_15704,N_8616,N_8697);
and U15705 (N_15705,N_7376,N_8325);
and U15706 (N_15706,N_11079,N_9074);
or U15707 (N_15707,N_9888,N_7682);
nand U15708 (N_15708,N_8420,N_6166);
nor U15709 (N_15709,N_9770,N_7863);
nand U15710 (N_15710,N_8229,N_6152);
and U15711 (N_15711,N_11993,N_10071);
nor U15712 (N_15712,N_9920,N_6084);
nand U15713 (N_15713,N_7673,N_10880);
xnor U15714 (N_15714,N_7955,N_10527);
and U15715 (N_15715,N_9807,N_9374);
or U15716 (N_15716,N_7553,N_11960);
or U15717 (N_15717,N_10092,N_7344);
or U15718 (N_15718,N_6012,N_11662);
or U15719 (N_15719,N_9466,N_6686);
and U15720 (N_15720,N_9529,N_8883);
and U15721 (N_15721,N_6854,N_7598);
nor U15722 (N_15722,N_9432,N_9568);
xor U15723 (N_15723,N_7906,N_11092);
xnor U15724 (N_15724,N_7371,N_7627);
and U15725 (N_15725,N_9815,N_6873);
or U15726 (N_15726,N_11337,N_11091);
nor U15727 (N_15727,N_8148,N_8070);
xor U15728 (N_15728,N_6069,N_11417);
nand U15729 (N_15729,N_7542,N_8049);
or U15730 (N_15730,N_8392,N_11641);
xnor U15731 (N_15731,N_9507,N_6086);
or U15732 (N_15732,N_8004,N_9815);
xor U15733 (N_15733,N_8238,N_11968);
nor U15734 (N_15734,N_7301,N_7989);
xor U15735 (N_15735,N_8989,N_7099);
xor U15736 (N_15736,N_10825,N_7565);
nand U15737 (N_15737,N_11184,N_6259);
nand U15738 (N_15738,N_10471,N_9500);
or U15739 (N_15739,N_6825,N_8824);
nand U15740 (N_15740,N_10197,N_10857);
and U15741 (N_15741,N_10876,N_10165);
nor U15742 (N_15742,N_6599,N_8391);
or U15743 (N_15743,N_9736,N_7366);
and U15744 (N_15744,N_9355,N_6957);
or U15745 (N_15745,N_8013,N_7361);
or U15746 (N_15746,N_8134,N_6543);
nand U15747 (N_15747,N_6221,N_9738);
nor U15748 (N_15748,N_6703,N_10760);
and U15749 (N_15749,N_6151,N_6907);
xnor U15750 (N_15750,N_6416,N_7367);
nor U15751 (N_15751,N_8513,N_9602);
xnor U15752 (N_15752,N_10622,N_6253);
nand U15753 (N_15753,N_10818,N_6075);
xor U15754 (N_15754,N_6570,N_9708);
or U15755 (N_15755,N_6578,N_9350);
and U15756 (N_15756,N_7543,N_9251);
or U15757 (N_15757,N_11817,N_9237);
nor U15758 (N_15758,N_9347,N_9469);
or U15759 (N_15759,N_6018,N_6123);
and U15760 (N_15760,N_10788,N_10139);
nand U15761 (N_15761,N_9050,N_7003);
xor U15762 (N_15762,N_8805,N_11579);
xor U15763 (N_15763,N_9169,N_6585);
nand U15764 (N_15764,N_6475,N_8566);
and U15765 (N_15765,N_6094,N_10112);
nor U15766 (N_15766,N_7995,N_7472);
or U15767 (N_15767,N_7458,N_9742);
nor U15768 (N_15768,N_7539,N_7088);
nand U15769 (N_15769,N_8138,N_11435);
and U15770 (N_15770,N_10343,N_10227);
xor U15771 (N_15771,N_8865,N_8653);
xnor U15772 (N_15772,N_6185,N_6816);
nor U15773 (N_15773,N_8612,N_6245);
and U15774 (N_15774,N_11858,N_7201);
and U15775 (N_15775,N_9813,N_6062);
xor U15776 (N_15776,N_7156,N_8532);
nand U15777 (N_15777,N_8922,N_6866);
nor U15778 (N_15778,N_10824,N_6703);
nand U15779 (N_15779,N_11678,N_6601);
nor U15780 (N_15780,N_6579,N_6545);
nor U15781 (N_15781,N_7947,N_11889);
xnor U15782 (N_15782,N_8200,N_6035);
and U15783 (N_15783,N_7448,N_6344);
and U15784 (N_15784,N_6360,N_11738);
nand U15785 (N_15785,N_8852,N_11602);
nor U15786 (N_15786,N_6413,N_7796);
nand U15787 (N_15787,N_8974,N_8714);
xnor U15788 (N_15788,N_8530,N_8613);
or U15789 (N_15789,N_6134,N_11963);
or U15790 (N_15790,N_8442,N_7615);
xor U15791 (N_15791,N_7305,N_10981);
and U15792 (N_15792,N_7652,N_9992);
nand U15793 (N_15793,N_10885,N_6319);
nand U15794 (N_15794,N_6085,N_8351);
and U15795 (N_15795,N_6037,N_10182);
nor U15796 (N_15796,N_6615,N_9266);
xnor U15797 (N_15797,N_10168,N_9656);
nor U15798 (N_15798,N_11109,N_6041);
xor U15799 (N_15799,N_8919,N_10062);
or U15800 (N_15800,N_7171,N_7625);
and U15801 (N_15801,N_9933,N_11952);
nand U15802 (N_15802,N_7905,N_6349);
nand U15803 (N_15803,N_8461,N_7668);
or U15804 (N_15804,N_8937,N_9776);
or U15805 (N_15805,N_8462,N_9870);
nand U15806 (N_15806,N_7854,N_8170);
nor U15807 (N_15807,N_11495,N_10247);
or U15808 (N_15808,N_9470,N_7886);
or U15809 (N_15809,N_11783,N_10596);
nor U15810 (N_15810,N_11910,N_6824);
or U15811 (N_15811,N_7464,N_11124);
xnor U15812 (N_15812,N_6645,N_8769);
nand U15813 (N_15813,N_8250,N_9911);
xor U15814 (N_15814,N_9272,N_6931);
nor U15815 (N_15815,N_7385,N_8031);
nand U15816 (N_15816,N_10093,N_7959);
or U15817 (N_15817,N_8083,N_11097);
or U15818 (N_15818,N_8705,N_7999);
and U15819 (N_15819,N_8422,N_6681);
and U15820 (N_15820,N_8743,N_7429);
xor U15821 (N_15821,N_7969,N_8361);
and U15822 (N_15822,N_8578,N_8409);
nand U15823 (N_15823,N_10285,N_6664);
or U15824 (N_15824,N_11387,N_10988);
nand U15825 (N_15825,N_11438,N_10983);
xnor U15826 (N_15826,N_7337,N_10521);
xnor U15827 (N_15827,N_10361,N_11085);
and U15828 (N_15828,N_7209,N_9406);
and U15829 (N_15829,N_7615,N_8772);
xnor U15830 (N_15830,N_8813,N_9270);
nor U15831 (N_15831,N_6891,N_7069);
xnor U15832 (N_15832,N_11543,N_10233);
xnor U15833 (N_15833,N_6722,N_8215);
or U15834 (N_15834,N_7740,N_6315);
xnor U15835 (N_15835,N_8954,N_8523);
and U15836 (N_15836,N_9530,N_10952);
or U15837 (N_15837,N_11855,N_6620);
or U15838 (N_15838,N_8405,N_8586);
nor U15839 (N_15839,N_7417,N_7860);
nor U15840 (N_15840,N_6944,N_6975);
nand U15841 (N_15841,N_9196,N_8645);
nor U15842 (N_15842,N_11687,N_7495);
and U15843 (N_15843,N_6730,N_11221);
and U15844 (N_15844,N_11510,N_8483);
xor U15845 (N_15845,N_8631,N_9748);
or U15846 (N_15846,N_6636,N_6286);
xor U15847 (N_15847,N_7134,N_6688);
nor U15848 (N_15848,N_6309,N_7406);
nor U15849 (N_15849,N_10551,N_9097);
and U15850 (N_15850,N_8591,N_10928);
nand U15851 (N_15851,N_8014,N_6646);
nor U15852 (N_15852,N_7938,N_10463);
xor U15853 (N_15853,N_8039,N_11294);
and U15854 (N_15854,N_11693,N_8182);
and U15855 (N_15855,N_8024,N_11100);
or U15856 (N_15856,N_11085,N_9248);
and U15857 (N_15857,N_9980,N_10898);
nand U15858 (N_15858,N_9826,N_6617);
or U15859 (N_15859,N_11778,N_11389);
xnor U15860 (N_15860,N_7431,N_8418);
xor U15861 (N_15861,N_6316,N_10249);
and U15862 (N_15862,N_7958,N_8090);
nand U15863 (N_15863,N_6814,N_7118);
or U15864 (N_15864,N_11603,N_8309);
nand U15865 (N_15865,N_7199,N_6148);
xnor U15866 (N_15866,N_6410,N_11107);
nor U15867 (N_15867,N_10360,N_8635);
and U15868 (N_15868,N_11122,N_8150);
and U15869 (N_15869,N_10140,N_9386);
or U15870 (N_15870,N_6088,N_10112);
xnor U15871 (N_15871,N_7713,N_8609);
or U15872 (N_15872,N_6322,N_8802);
nor U15873 (N_15873,N_8451,N_9578);
and U15874 (N_15874,N_8934,N_9055);
nor U15875 (N_15875,N_8164,N_7137);
xnor U15876 (N_15876,N_6304,N_10259);
xnor U15877 (N_15877,N_11383,N_7999);
and U15878 (N_15878,N_8475,N_7412);
or U15879 (N_15879,N_6919,N_11759);
nand U15880 (N_15880,N_6570,N_11209);
nor U15881 (N_15881,N_9008,N_10962);
or U15882 (N_15882,N_6848,N_6020);
nor U15883 (N_15883,N_10439,N_6196);
nor U15884 (N_15884,N_7178,N_9276);
xor U15885 (N_15885,N_7551,N_11240);
xor U15886 (N_15886,N_9427,N_9440);
or U15887 (N_15887,N_6661,N_9229);
and U15888 (N_15888,N_8761,N_9536);
or U15889 (N_15889,N_7459,N_9174);
nand U15890 (N_15890,N_10197,N_10749);
and U15891 (N_15891,N_6079,N_7826);
xnor U15892 (N_15892,N_9647,N_6200);
nor U15893 (N_15893,N_6738,N_10893);
xor U15894 (N_15894,N_9891,N_10025);
and U15895 (N_15895,N_11494,N_10991);
nor U15896 (N_15896,N_10232,N_6447);
nand U15897 (N_15897,N_7033,N_10865);
and U15898 (N_15898,N_10403,N_10963);
and U15899 (N_15899,N_8061,N_11732);
xnor U15900 (N_15900,N_9786,N_6611);
xnor U15901 (N_15901,N_6989,N_9844);
nand U15902 (N_15902,N_7401,N_7022);
xnor U15903 (N_15903,N_7342,N_7128);
nor U15904 (N_15904,N_9051,N_6143);
and U15905 (N_15905,N_10499,N_7360);
or U15906 (N_15906,N_7330,N_8875);
nand U15907 (N_15907,N_9772,N_8684);
xnor U15908 (N_15908,N_8650,N_8804);
nor U15909 (N_15909,N_11338,N_10116);
xnor U15910 (N_15910,N_8056,N_8119);
xnor U15911 (N_15911,N_11694,N_10826);
and U15912 (N_15912,N_7303,N_11215);
xor U15913 (N_15913,N_10490,N_11032);
or U15914 (N_15914,N_7314,N_9044);
or U15915 (N_15915,N_7305,N_8484);
nor U15916 (N_15916,N_9089,N_8749);
nand U15917 (N_15917,N_9727,N_10154);
and U15918 (N_15918,N_10548,N_11845);
xnor U15919 (N_15919,N_6055,N_11191);
nor U15920 (N_15920,N_6737,N_10749);
xor U15921 (N_15921,N_7229,N_9150);
or U15922 (N_15922,N_8365,N_11961);
and U15923 (N_15923,N_10390,N_9526);
xor U15924 (N_15924,N_6189,N_10061);
and U15925 (N_15925,N_10271,N_9442);
nor U15926 (N_15926,N_10004,N_6723);
nand U15927 (N_15927,N_7559,N_8891);
and U15928 (N_15928,N_6862,N_10043);
and U15929 (N_15929,N_9103,N_10183);
nor U15930 (N_15930,N_10226,N_10586);
xor U15931 (N_15931,N_10433,N_10924);
nand U15932 (N_15932,N_7822,N_9314);
and U15933 (N_15933,N_10383,N_8694);
xnor U15934 (N_15934,N_9727,N_6352);
nor U15935 (N_15935,N_6882,N_6875);
nor U15936 (N_15936,N_8949,N_8671);
or U15937 (N_15937,N_6201,N_8860);
nor U15938 (N_15938,N_10003,N_11122);
nor U15939 (N_15939,N_9978,N_11598);
nand U15940 (N_15940,N_9096,N_7322);
or U15941 (N_15941,N_10010,N_10242);
nand U15942 (N_15942,N_8697,N_8174);
nor U15943 (N_15943,N_7596,N_7631);
and U15944 (N_15944,N_6514,N_6168);
xor U15945 (N_15945,N_10200,N_6270);
or U15946 (N_15946,N_10458,N_11693);
and U15947 (N_15947,N_10434,N_11725);
nand U15948 (N_15948,N_9685,N_7320);
nand U15949 (N_15949,N_6949,N_7792);
and U15950 (N_15950,N_11082,N_9339);
nor U15951 (N_15951,N_9332,N_8449);
xor U15952 (N_15952,N_6864,N_10793);
nand U15953 (N_15953,N_6026,N_7411);
and U15954 (N_15954,N_9465,N_8922);
xor U15955 (N_15955,N_9683,N_9296);
xor U15956 (N_15956,N_8431,N_9443);
or U15957 (N_15957,N_9661,N_8697);
and U15958 (N_15958,N_8344,N_11904);
and U15959 (N_15959,N_8997,N_11676);
xnor U15960 (N_15960,N_11814,N_10205);
xor U15961 (N_15961,N_10240,N_11179);
xnor U15962 (N_15962,N_7676,N_9448);
or U15963 (N_15963,N_10024,N_10978);
nand U15964 (N_15964,N_9679,N_11809);
and U15965 (N_15965,N_6338,N_8831);
nor U15966 (N_15966,N_6312,N_9828);
xor U15967 (N_15967,N_6336,N_8796);
nand U15968 (N_15968,N_9754,N_6129);
xnor U15969 (N_15969,N_8810,N_7377);
nand U15970 (N_15970,N_6137,N_8029);
nand U15971 (N_15971,N_11123,N_10623);
nor U15972 (N_15972,N_6113,N_7414);
nand U15973 (N_15973,N_9087,N_6585);
and U15974 (N_15974,N_9132,N_8384);
or U15975 (N_15975,N_11065,N_6562);
or U15976 (N_15976,N_7112,N_8283);
nor U15977 (N_15977,N_8818,N_8534);
nand U15978 (N_15978,N_7925,N_10647);
and U15979 (N_15979,N_9482,N_9447);
xor U15980 (N_15980,N_11539,N_6356);
nand U15981 (N_15981,N_8466,N_7677);
or U15982 (N_15982,N_10169,N_11028);
nand U15983 (N_15983,N_10522,N_9438);
nand U15984 (N_15984,N_10812,N_11919);
nor U15985 (N_15985,N_8482,N_6778);
and U15986 (N_15986,N_9421,N_11011);
xor U15987 (N_15987,N_11731,N_7234);
or U15988 (N_15988,N_7554,N_11707);
or U15989 (N_15989,N_10369,N_7850);
nand U15990 (N_15990,N_7265,N_10533);
and U15991 (N_15991,N_8651,N_10964);
nand U15992 (N_15992,N_10634,N_8374);
nand U15993 (N_15993,N_9196,N_7297);
xnor U15994 (N_15994,N_7501,N_6489);
and U15995 (N_15995,N_6099,N_6019);
and U15996 (N_15996,N_6853,N_8759);
or U15997 (N_15997,N_8341,N_6845);
or U15998 (N_15998,N_8810,N_7894);
xnor U15999 (N_15999,N_6521,N_10485);
and U16000 (N_16000,N_9694,N_9356);
or U16001 (N_16001,N_10013,N_10168);
or U16002 (N_16002,N_10710,N_11750);
and U16003 (N_16003,N_7975,N_11669);
nor U16004 (N_16004,N_9773,N_10166);
or U16005 (N_16005,N_8877,N_6755);
nor U16006 (N_16006,N_9538,N_9356);
xor U16007 (N_16007,N_6433,N_6782);
or U16008 (N_16008,N_8626,N_10225);
and U16009 (N_16009,N_6944,N_6733);
or U16010 (N_16010,N_6480,N_7074);
or U16011 (N_16011,N_8433,N_9706);
nor U16012 (N_16012,N_8256,N_6274);
nor U16013 (N_16013,N_6347,N_11065);
or U16014 (N_16014,N_6469,N_11259);
nor U16015 (N_16015,N_9910,N_10481);
xnor U16016 (N_16016,N_10660,N_6216);
nand U16017 (N_16017,N_9509,N_8676);
or U16018 (N_16018,N_11398,N_8062);
or U16019 (N_16019,N_11069,N_7623);
nor U16020 (N_16020,N_8934,N_11109);
nand U16021 (N_16021,N_10667,N_11825);
and U16022 (N_16022,N_7268,N_8383);
nor U16023 (N_16023,N_11832,N_8810);
nor U16024 (N_16024,N_9751,N_11682);
nand U16025 (N_16025,N_7386,N_11099);
nand U16026 (N_16026,N_10161,N_8433);
nor U16027 (N_16027,N_7267,N_10240);
and U16028 (N_16028,N_7866,N_11367);
xnor U16029 (N_16029,N_10434,N_11968);
or U16030 (N_16030,N_7252,N_7084);
and U16031 (N_16031,N_9570,N_9509);
or U16032 (N_16032,N_8867,N_7684);
xnor U16033 (N_16033,N_9998,N_6059);
nor U16034 (N_16034,N_10773,N_11281);
or U16035 (N_16035,N_10402,N_9372);
nor U16036 (N_16036,N_8126,N_10548);
or U16037 (N_16037,N_9814,N_8767);
nor U16038 (N_16038,N_11662,N_11124);
or U16039 (N_16039,N_10472,N_10934);
xnor U16040 (N_16040,N_8046,N_7721);
xnor U16041 (N_16041,N_9780,N_6713);
xor U16042 (N_16042,N_8409,N_6876);
and U16043 (N_16043,N_10033,N_9125);
nor U16044 (N_16044,N_9466,N_10445);
nor U16045 (N_16045,N_11760,N_9003);
nand U16046 (N_16046,N_6246,N_8920);
and U16047 (N_16047,N_7332,N_10714);
xnor U16048 (N_16048,N_8718,N_7423);
xor U16049 (N_16049,N_8035,N_11569);
nor U16050 (N_16050,N_6911,N_7076);
xor U16051 (N_16051,N_7163,N_8848);
or U16052 (N_16052,N_6721,N_9225);
and U16053 (N_16053,N_11653,N_10143);
or U16054 (N_16054,N_11209,N_8283);
xor U16055 (N_16055,N_11120,N_6683);
and U16056 (N_16056,N_7771,N_7613);
nand U16057 (N_16057,N_8966,N_11931);
and U16058 (N_16058,N_10859,N_10395);
nor U16059 (N_16059,N_8519,N_10128);
xor U16060 (N_16060,N_10827,N_9301);
and U16061 (N_16061,N_9462,N_8602);
nand U16062 (N_16062,N_8286,N_8486);
xor U16063 (N_16063,N_11076,N_8376);
nor U16064 (N_16064,N_8767,N_10029);
and U16065 (N_16065,N_9866,N_8716);
nand U16066 (N_16066,N_9653,N_9415);
or U16067 (N_16067,N_9951,N_9308);
nor U16068 (N_16068,N_11311,N_8739);
nand U16069 (N_16069,N_9293,N_7293);
and U16070 (N_16070,N_11730,N_7561);
and U16071 (N_16071,N_8721,N_7583);
xnor U16072 (N_16072,N_9964,N_7837);
nand U16073 (N_16073,N_9428,N_9622);
or U16074 (N_16074,N_9930,N_7306);
or U16075 (N_16075,N_10169,N_6147);
xnor U16076 (N_16076,N_10123,N_10533);
nand U16077 (N_16077,N_9741,N_10088);
nand U16078 (N_16078,N_10010,N_8989);
nand U16079 (N_16079,N_11965,N_10733);
nand U16080 (N_16080,N_8439,N_11503);
nand U16081 (N_16081,N_8853,N_6117);
and U16082 (N_16082,N_6157,N_11186);
and U16083 (N_16083,N_11309,N_10343);
xor U16084 (N_16084,N_10745,N_9459);
and U16085 (N_16085,N_7173,N_9923);
nor U16086 (N_16086,N_8509,N_6780);
nor U16087 (N_16087,N_8486,N_8595);
nand U16088 (N_16088,N_6167,N_11583);
and U16089 (N_16089,N_11993,N_11542);
and U16090 (N_16090,N_9132,N_11406);
or U16091 (N_16091,N_9808,N_9519);
and U16092 (N_16092,N_10493,N_11514);
xnor U16093 (N_16093,N_10653,N_10536);
or U16094 (N_16094,N_7847,N_7262);
or U16095 (N_16095,N_8865,N_8516);
and U16096 (N_16096,N_10189,N_7529);
or U16097 (N_16097,N_6481,N_7187);
nand U16098 (N_16098,N_10144,N_11754);
and U16099 (N_16099,N_9290,N_11190);
or U16100 (N_16100,N_11553,N_9443);
nor U16101 (N_16101,N_8779,N_8528);
or U16102 (N_16102,N_9684,N_10146);
nor U16103 (N_16103,N_11448,N_8314);
or U16104 (N_16104,N_9216,N_10257);
or U16105 (N_16105,N_6909,N_8597);
xnor U16106 (N_16106,N_11813,N_11364);
nand U16107 (N_16107,N_9005,N_9560);
or U16108 (N_16108,N_10333,N_7275);
nor U16109 (N_16109,N_10244,N_8059);
xor U16110 (N_16110,N_10044,N_7761);
nand U16111 (N_16111,N_10529,N_11345);
nand U16112 (N_16112,N_10810,N_7787);
or U16113 (N_16113,N_11148,N_10470);
nor U16114 (N_16114,N_8646,N_11313);
and U16115 (N_16115,N_8619,N_11489);
or U16116 (N_16116,N_7451,N_11563);
nor U16117 (N_16117,N_8036,N_10967);
nor U16118 (N_16118,N_8970,N_8814);
xnor U16119 (N_16119,N_9800,N_10918);
nor U16120 (N_16120,N_9945,N_10936);
xor U16121 (N_16121,N_11282,N_9047);
xnor U16122 (N_16122,N_6124,N_8077);
nand U16123 (N_16123,N_7574,N_8951);
nor U16124 (N_16124,N_8430,N_7367);
nand U16125 (N_16125,N_7442,N_11834);
xnor U16126 (N_16126,N_10897,N_6769);
nand U16127 (N_16127,N_6907,N_10891);
nor U16128 (N_16128,N_9490,N_9694);
or U16129 (N_16129,N_6911,N_11323);
nor U16130 (N_16130,N_8637,N_7231);
or U16131 (N_16131,N_10944,N_8380);
nand U16132 (N_16132,N_9871,N_8488);
nand U16133 (N_16133,N_10000,N_6788);
or U16134 (N_16134,N_7784,N_9933);
and U16135 (N_16135,N_7691,N_6310);
or U16136 (N_16136,N_6398,N_7746);
xor U16137 (N_16137,N_9501,N_9013);
and U16138 (N_16138,N_9837,N_7263);
nor U16139 (N_16139,N_10063,N_6354);
xnor U16140 (N_16140,N_8709,N_6297);
nand U16141 (N_16141,N_6854,N_6841);
nand U16142 (N_16142,N_10943,N_6529);
nor U16143 (N_16143,N_9968,N_6973);
nor U16144 (N_16144,N_8143,N_10716);
xor U16145 (N_16145,N_7177,N_6204);
xor U16146 (N_16146,N_9407,N_10581);
or U16147 (N_16147,N_11720,N_6526);
nor U16148 (N_16148,N_7645,N_6181);
or U16149 (N_16149,N_8758,N_9821);
or U16150 (N_16150,N_8521,N_6066);
xor U16151 (N_16151,N_7223,N_6905);
and U16152 (N_16152,N_6705,N_8894);
nand U16153 (N_16153,N_7052,N_9325);
or U16154 (N_16154,N_7537,N_10435);
or U16155 (N_16155,N_10360,N_10070);
or U16156 (N_16156,N_6984,N_11830);
nand U16157 (N_16157,N_7511,N_8234);
nor U16158 (N_16158,N_9532,N_11148);
nand U16159 (N_16159,N_9201,N_10389);
or U16160 (N_16160,N_6310,N_8149);
or U16161 (N_16161,N_11544,N_8952);
or U16162 (N_16162,N_11232,N_11444);
and U16163 (N_16163,N_9412,N_7027);
or U16164 (N_16164,N_9853,N_11981);
and U16165 (N_16165,N_10597,N_8155);
nor U16166 (N_16166,N_7351,N_6878);
or U16167 (N_16167,N_11609,N_10831);
nand U16168 (N_16168,N_11678,N_8590);
nor U16169 (N_16169,N_6505,N_11113);
or U16170 (N_16170,N_7285,N_11458);
or U16171 (N_16171,N_11967,N_7973);
nand U16172 (N_16172,N_8448,N_10119);
nor U16173 (N_16173,N_11729,N_8459);
or U16174 (N_16174,N_7620,N_9911);
nand U16175 (N_16175,N_6702,N_9768);
xnor U16176 (N_16176,N_7465,N_11319);
and U16177 (N_16177,N_6192,N_10390);
nor U16178 (N_16178,N_11703,N_10806);
nand U16179 (N_16179,N_8742,N_10017);
and U16180 (N_16180,N_6561,N_11142);
nand U16181 (N_16181,N_10267,N_10765);
nand U16182 (N_16182,N_9291,N_8360);
nor U16183 (N_16183,N_11081,N_11644);
xor U16184 (N_16184,N_6956,N_8025);
and U16185 (N_16185,N_11725,N_11775);
and U16186 (N_16186,N_11677,N_8550);
or U16187 (N_16187,N_8905,N_9945);
or U16188 (N_16188,N_7676,N_8377);
nand U16189 (N_16189,N_11117,N_10376);
xor U16190 (N_16190,N_8676,N_7358);
or U16191 (N_16191,N_6290,N_9481);
nand U16192 (N_16192,N_6595,N_8393);
or U16193 (N_16193,N_7542,N_6890);
and U16194 (N_16194,N_11935,N_6091);
nor U16195 (N_16195,N_7393,N_10998);
nor U16196 (N_16196,N_7008,N_7500);
or U16197 (N_16197,N_6153,N_10602);
and U16198 (N_16198,N_9689,N_9625);
nor U16199 (N_16199,N_11008,N_8536);
or U16200 (N_16200,N_8203,N_7645);
xor U16201 (N_16201,N_10514,N_6843);
nand U16202 (N_16202,N_9393,N_8672);
and U16203 (N_16203,N_6666,N_10567);
or U16204 (N_16204,N_7764,N_7428);
nand U16205 (N_16205,N_10406,N_8529);
nand U16206 (N_16206,N_6920,N_6788);
xor U16207 (N_16207,N_11754,N_6089);
nor U16208 (N_16208,N_11889,N_9629);
and U16209 (N_16209,N_6762,N_9239);
nand U16210 (N_16210,N_10091,N_10981);
or U16211 (N_16211,N_6672,N_6943);
and U16212 (N_16212,N_10042,N_8387);
xor U16213 (N_16213,N_8245,N_11889);
or U16214 (N_16214,N_9549,N_6313);
xor U16215 (N_16215,N_8150,N_10458);
nor U16216 (N_16216,N_6250,N_10447);
xor U16217 (N_16217,N_11257,N_10575);
or U16218 (N_16218,N_8078,N_6491);
xor U16219 (N_16219,N_6260,N_10204);
xor U16220 (N_16220,N_9300,N_9041);
nor U16221 (N_16221,N_11308,N_10350);
nand U16222 (N_16222,N_8978,N_11088);
nor U16223 (N_16223,N_11265,N_11213);
and U16224 (N_16224,N_10165,N_7017);
xnor U16225 (N_16225,N_8242,N_7580);
nor U16226 (N_16226,N_11998,N_10385);
or U16227 (N_16227,N_11598,N_11835);
xor U16228 (N_16228,N_9129,N_9624);
or U16229 (N_16229,N_7339,N_9431);
and U16230 (N_16230,N_8914,N_7479);
nand U16231 (N_16231,N_10694,N_11795);
xor U16232 (N_16232,N_6295,N_10622);
nand U16233 (N_16233,N_10497,N_11988);
nand U16234 (N_16234,N_6634,N_6487);
xor U16235 (N_16235,N_11211,N_10252);
or U16236 (N_16236,N_10725,N_9920);
xor U16237 (N_16237,N_6121,N_8572);
nand U16238 (N_16238,N_6694,N_10147);
nor U16239 (N_16239,N_9889,N_10399);
xor U16240 (N_16240,N_8796,N_9704);
and U16241 (N_16241,N_11335,N_9124);
nor U16242 (N_16242,N_8703,N_9775);
nor U16243 (N_16243,N_10124,N_8355);
nor U16244 (N_16244,N_8654,N_9194);
nor U16245 (N_16245,N_8773,N_10893);
nor U16246 (N_16246,N_8005,N_6242);
xor U16247 (N_16247,N_6917,N_11435);
nand U16248 (N_16248,N_9824,N_11866);
nand U16249 (N_16249,N_7597,N_8084);
xnor U16250 (N_16250,N_9609,N_8095);
nor U16251 (N_16251,N_10116,N_6468);
or U16252 (N_16252,N_10715,N_9669);
or U16253 (N_16253,N_9671,N_6440);
xor U16254 (N_16254,N_10645,N_7637);
xnor U16255 (N_16255,N_8655,N_7676);
nor U16256 (N_16256,N_6817,N_11279);
nand U16257 (N_16257,N_7717,N_9916);
nor U16258 (N_16258,N_11797,N_11606);
xnor U16259 (N_16259,N_9273,N_6486);
xnor U16260 (N_16260,N_10059,N_8466);
nand U16261 (N_16261,N_8058,N_11301);
nor U16262 (N_16262,N_11258,N_8289);
xor U16263 (N_16263,N_9829,N_11092);
nor U16264 (N_16264,N_6565,N_8502);
and U16265 (N_16265,N_7350,N_9457);
and U16266 (N_16266,N_9840,N_10191);
and U16267 (N_16267,N_9688,N_8568);
or U16268 (N_16268,N_7884,N_10170);
and U16269 (N_16269,N_11696,N_10958);
nor U16270 (N_16270,N_6545,N_10655);
nor U16271 (N_16271,N_6445,N_10974);
nand U16272 (N_16272,N_6714,N_11340);
nor U16273 (N_16273,N_10734,N_7563);
or U16274 (N_16274,N_7859,N_11831);
and U16275 (N_16275,N_7615,N_6495);
and U16276 (N_16276,N_7562,N_10997);
nor U16277 (N_16277,N_10311,N_6033);
and U16278 (N_16278,N_8747,N_10730);
or U16279 (N_16279,N_10022,N_11019);
and U16280 (N_16280,N_9051,N_11963);
xor U16281 (N_16281,N_7103,N_8711);
nor U16282 (N_16282,N_10831,N_6778);
xnor U16283 (N_16283,N_7136,N_11032);
and U16284 (N_16284,N_9105,N_8274);
xor U16285 (N_16285,N_11982,N_7667);
nand U16286 (N_16286,N_9327,N_9332);
or U16287 (N_16287,N_9475,N_7470);
nand U16288 (N_16288,N_9118,N_6456);
and U16289 (N_16289,N_9761,N_9843);
or U16290 (N_16290,N_7185,N_7879);
xnor U16291 (N_16291,N_8838,N_9398);
nor U16292 (N_16292,N_11007,N_9262);
xor U16293 (N_16293,N_6322,N_6502);
nor U16294 (N_16294,N_9921,N_11875);
nand U16295 (N_16295,N_6367,N_8352);
and U16296 (N_16296,N_9420,N_6904);
nand U16297 (N_16297,N_9589,N_10932);
nand U16298 (N_16298,N_11072,N_8415);
nor U16299 (N_16299,N_10147,N_9137);
xnor U16300 (N_16300,N_9122,N_11071);
nor U16301 (N_16301,N_10332,N_8726);
xor U16302 (N_16302,N_11113,N_11441);
and U16303 (N_16303,N_8919,N_6343);
nor U16304 (N_16304,N_8063,N_9022);
or U16305 (N_16305,N_8160,N_7935);
xor U16306 (N_16306,N_10164,N_11862);
xor U16307 (N_16307,N_8739,N_7032);
or U16308 (N_16308,N_7031,N_11787);
and U16309 (N_16309,N_10141,N_7220);
nand U16310 (N_16310,N_11799,N_10373);
and U16311 (N_16311,N_6482,N_7450);
xor U16312 (N_16312,N_11862,N_6016);
xnor U16313 (N_16313,N_11965,N_9381);
nor U16314 (N_16314,N_10080,N_8885);
or U16315 (N_16315,N_10103,N_8383);
nand U16316 (N_16316,N_6610,N_9537);
nand U16317 (N_16317,N_8797,N_7155);
xnor U16318 (N_16318,N_6098,N_7995);
or U16319 (N_16319,N_7260,N_11512);
and U16320 (N_16320,N_8067,N_8869);
or U16321 (N_16321,N_6930,N_11094);
xnor U16322 (N_16322,N_10054,N_8468);
and U16323 (N_16323,N_9112,N_7208);
or U16324 (N_16324,N_7640,N_10127);
nor U16325 (N_16325,N_9041,N_10579);
nand U16326 (N_16326,N_11318,N_10596);
nand U16327 (N_16327,N_11010,N_9886);
nand U16328 (N_16328,N_6906,N_11017);
xor U16329 (N_16329,N_10040,N_10668);
nor U16330 (N_16330,N_7507,N_8557);
xor U16331 (N_16331,N_8206,N_11274);
nor U16332 (N_16332,N_10325,N_9605);
xor U16333 (N_16333,N_8997,N_8052);
xnor U16334 (N_16334,N_10894,N_7736);
or U16335 (N_16335,N_8591,N_6400);
or U16336 (N_16336,N_10734,N_11653);
or U16337 (N_16337,N_8941,N_10922);
nand U16338 (N_16338,N_10503,N_7914);
xnor U16339 (N_16339,N_10735,N_10337);
nor U16340 (N_16340,N_10176,N_8914);
or U16341 (N_16341,N_9237,N_9787);
and U16342 (N_16342,N_7032,N_8827);
xor U16343 (N_16343,N_8004,N_8125);
or U16344 (N_16344,N_9644,N_8297);
nand U16345 (N_16345,N_7885,N_7295);
nor U16346 (N_16346,N_9381,N_11418);
or U16347 (N_16347,N_10208,N_8536);
nor U16348 (N_16348,N_8478,N_11723);
xnor U16349 (N_16349,N_8103,N_10384);
and U16350 (N_16350,N_11867,N_10633);
xnor U16351 (N_16351,N_11654,N_6144);
or U16352 (N_16352,N_11101,N_10589);
or U16353 (N_16353,N_8696,N_10372);
xor U16354 (N_16354,N_7841,N_6404);
nand U16355 (N_16355,N_9257,N_8165);
nand U16356 (N_16356,N_10929,N_9913);
xor U16357 (N_16357,N_11134,N_7722);
or U16358 (N_16358,N_8191,N_11022);
or U16359 (N_16359,N_11444,N_7286);
nor U16360 (N_16360,N_7918,N_7725);
nor U16361 (N_16361,N_6729,N_8122);
nand U16362 (N_16362,N_8518,N_8142);
nor U16363 (N_16363,N_11770,N_9586);
and U16364 (N_16364,N_11555,N_7763);
xnor U16365 (N_16365,N_11728,N_10395);
nand U16366 (N_16366,N_7717,N_10252);
or U16367 (N_16367,N_10317,N_11633);
and U16368 (N_16368,N_6110,N_7221);
and U16369 (N_16369,N_8508,N_9226);
and U16370 (N_16370,N_11483,N_9213);
nand U16371 (N_16371,N_10689,N_10076);
nand U16372 (N_16372,N_9112,N_7687);
nand U16373 (N_16373,N_10686,N_9467);
or U16374 (N_16374,N_8724,N_10410);
or U16375 (N_16375,N_10718,N_9198);
nor U16376 (N_16376,N_9490,N_11264);
and U16377 (N_16377,N_10114,N_7879);
nor U16378 (N_16378,N_7965,N_8164);
nand U16379 (N_16379,N_10115,N_9463);
and U16380 (N_16380,N_7460,N_8547);
and U16381 (N_16381,N_9811,N_9262);
xor U16382 (N_16382,N_6572,N_11575);
nor U16383 (N_16383,N_8516,N_8791);
and U16384 (N_16384,N_6014,N_10456);
or U16385 (N_16385,N_8229,N_11168);
and U16386 (N_16386,N_7882,N_10039);
nand U16387 (N_16387,N_10912,N_9002);
nand U16388 (N_16388,N_10943,N_9248);
xnor U16389 (N_16389,N_6898,N_7700);
or U16390 (N_16390,N_6808,N_10051);
nor U16391 (N_16391,N_10955,N_7689);
nand U16392 (N_16392,N_10505,N_11707);
nor U16393 (N_16393,N_9998,N_9270);
xor U16394 (N_16394,N_11446,N_9775);
nand U16395 (N_16395,N_9718,N_10229);
nor U16396 (N_16396,N_11647,N_9815);
and U16397 (N_16397,N_9457,N_11290);
and U16398 (N_16398,N_8846,N_10089);
xor U16399 (N_16399,N_7504,N_11926);
nand U16400 (N_16400,N_6460,N_9984);
nor U16401 (N_16401,N_10021,N_9005);
xnor U16402 (N_16402,N_6463,N_8442);
nor U16403 (N_16403,N_8343,N_8073);
nor U16404 (N_16404,N_6529,N_9965);
xnor U16405 (N_16405,N_8908,N_11457);
and U16406 (N_16406,N_6317,N_11652);
and U16407 (N_16407,N_10717,N_7071);
and U16408 (N_16408,N_9680,N_11571);
nor U16409 (N_16409,N_10137,N_6264);
or U16410 (N_16410,N_6870,N_11366);
and U16411 (N_16411,N_6583,N_6438);
or U16412 (N_16412,N_11416,N_7499);
nand U16413 (N_16413,N_9073,N_7290);
or U16414 (N_16414,N_9236,N_8330);
nand U16415 (N_16415,N_9753,N_10557);
xnor U16416 (N_16416,N_9103,N_6241);
nor U16417 (N_16417,N_6780,N_9720);
xor U16418 (N_16418,N_11382,N_10672);
or U16419 (N_16419,N_8144,N_9306);
nor U16420 (N_16420,N_11260,N_6089);
nand U16421 (N_16421,N_6987,N_8740);
and U16422 (N_16422,N_8453,N_10933);
nor U16423 (N_16423,N_8881,N_10410);
and U16424 (N_16424,N_11979,N_8478);
nand U16425 (N_16425,N_7762,N_8921);
and U16426 (N_16426,N_11928,N_7806);
xor U16427 (N_16427,N_6656,N_9985);
or U16428 (N_16428,N_7862,N_8137);
and U16429 (N_16429,N_9421,N_6864);
nor U16430 (N_16430,N_6652,N_10955);
xor U16431 (N_16431,N_7534,N_9899);
xor U16432 (N_16432,N_11364,N_10188);
nor U16433 (N_16433,N_11974,N_9803);
nand U16434 (N_16434,N_7711,N_11345);
xnor U16435 (N_16435,N_6780,N_10535);
and U16436 (N_16436,N_8415,N_7879);
and U16437 (N_16437,N_11562,N_9897);
nand U16438 (N_16438,N_8672,N_10637);
and U16439 (N_16439,N_6103,N_10812);
nor U16440 (N_16440,N_11509,N_11596);
or U16441 (N_16441,N_6573,N_10058);
nand U16442 (N_16442,N_9528,N_11572);
nand U16443 (N_16443,N_9376,N_7027);
nand U16444 (N_16444,N_8036,N_7196);
xor U16445 (N_16445,N_11183,N_10048);
xor U16446 (N_16446,N_9057,N_8311);
nor U16447 (N_16447,N_7978,N_11942);
nand U16448 (N_16448,N_8592,N_10933);
nor U16449 (N_16449,N_10111,N_7160);
and U16450 (N_16450,N_6138,N_11188);
or U16451 (N_16451,N_7222,N_11156);
nor U16452 (N_16452,N_11681,N_6218);
and U16453 (N_16453,N_8019,N_8050);
and U16454 (N_16454,N_7083,N_6342);
xor U16455 (N_16455,N_9847,N_8984);
nand U16456 (N_16456,N_11058,N_11375);
nand U16457 (N_16457,N_11711,N_6468);
and U16458 (N_16458,N_11382,N_11825);
and U16459 (N_16459,N_7786,N_7562);
nand U16460 (N_16460,N_7621,N_6292);
and U16461 (N_16461,N_10906,N_7125);
and U16462 (N_16462,N_11238,N_10133);
nand U16463 (N_16463,N_10009,N_10692);
xnor U16464 (N_16464,N_10939,N_6709);
xor U16465 (N_16465,N_11899,N_11906);
and U16466 (N_16466,N_9845,N_9624);
xor U16467 (N_16467,N_8963,N_10460);
xor U16468 (N_16468,N_6067,N_8026);
and U16469 (N_16469,N_9823,N_9420);
xor U16470 (N_16470,N_10342,N_6251);
and U16471 (N_16471,N_10316,N_7185);
nor U16472 (N_16472,N_6885,N_10120);
and U16473 (N_16473,N_10327,N_6461);
nand U16474 (N_16474,N_11682,N_7646);
or U16475 (N_16475,N_7266,N_6959);
nand U16476 (N_16476,N_10851,N_6543);
or U16477 (N_16477,N_8602,N_9350);
and U16478 (N_16478,N_9669,N_6707);
or U16479 (N_16479,N_11738,N_11841);
and U16480 (N_16480,N_8004,N_10405);
nor U16481 (N_16481,N_9692,N_6932);
or U16482 (N_16482,N_6997,N_6382);
nand U16483 (N_16483,N_7265,N_8479);
and U16484 (N_16484,N_9517,N_10819);
nor U16485 (N_16485,N_9295,N_9657);
nor U16486 (N_16486,N_11562,N_11891);
xor U16487 (N_16487,N_9911,N_6498);
nor U16488 (N_16488,N_8434,N_9884);
xor U16489 (N_16489,N_9522,N_10174);
nand U16490 (N_16490,N_11177,N_9511);
nor U16491 (N_16491,N_6679,N_6287);
nor U16492 (N_16492,N_10298,N_11851);
and U16493 (N_16493,N_7326,N_8768);
nand U16494 (N_16494,N_11624,N_11667);
and U16495 (N_16495,N_8643,N_10318);
or U16496 (N_16496,N_8824,N_11168);
and U16497 (N_16497,N_7952,N_6786);
and U16498 (N_16498,N_8855,N_8215);
and U16499 (N_16499,N_10390,N_7807);
nor U16500 (N_16500,N_7357,N_7368);
or U16501 (N_16501,N_6840,N_6910);
and U16502 (N_16502,N_9379,N_10085);
nand U16503 (N_16503,N_8523,N_8870);
and U16504 (N_16504,N_8447,N_10842);
or U16505 (N_16505,N_6238,N_7924);
nand U16506 (N_16506,N_9539,N_10578);
and U16507 (N_16507,N_7368,N_8492);
and U16508 (N_16508,N_7078,N_10076);
nor U16509 (N_16509,N_11851,N_10891);
nand U16510 (N_16510,N_7842,N_7475);
and U16511 (N_16511,N_6939,N_9873);
nand U16512 (N_16512,N_6303,N_9391);
and U16513 (N_16513,N_8956,N_9942);
and U16514 (N_16514,N_9390,N_8807);
nand U16515 (N_16515,N_7139,N_10665);
xnor U16516 (N_16516,N_6697,N_9417);
xor U16517 (N_16517,N_6391,N_10106);
and U16518 (N_16518,N_7510,N_9110);
xor U16519 (N_16519,N_11253,N_7868);
or U16520 (N_16520,N_7704,N_10521);
nor U16521 (N_16521,N_10024,N_7231);
nand U16522 (N_16522,N_9268,N_9156);
nor U16523 (N_16523,N_11123,N_10607);
or U16524 (N_16524,N_7591,N_8973);
nor U16525 (N_16525,N_10157,N_9517);
nand U16526 (N_16526,N_7838,N_9971);
and U16527 (N_16527,N_11545,N_8068);
or U16528 (N_16528,N_6178,N_7212);
nor U16529 (N_16529,N_7246,N_10335);
nor U16530 (N_16530,N_6843,N_10751);
xnor U16531 (N_16531,N_9763,N_10649);
xnor U16532 (N_16532,N_11096,N_10736);
and U16533 (N_16533,N_11650,N_6319);
and U16534 (N_16534,N_8016,N_11214);
nor U16535 (N_16535,N_8068,N_9437);
xor U16536 (N_16536,N_11418,N_9415);
and U16537 (N_16537,N_7557,N_9369);
xnor U16538 (N_16538,N_9794,N_8381);
nand U16539 (N_16539,N_8820,N_11060);
and U16540 (N_16540,N_9888,N_8513);
xnor U16541 (N_16541,N_8758,N_8230);
or U16542 (N_16542,N_8682,N_8564);
nor U16543 (N_16543,N_11587,N_11471);
or U16544 (N_16544,N_7227,N_11400);
nand U16545 (N_16545,N_11998,N_8150);
xnor U16546 (N_16546,N_7930,N_11367);
nor U16547 (N_16547,N_9223,N_10758);
or U16548 (N_16548,N_11397,N_6609);
nand U16549 (N_16549,N_10683,N_9759);
and U16550 (N_16550,N_7050,N_11407);
nor U16551 (N_16551,N_11316,N_8622);
xor U16552 (N_16552,N_9949,N_9206);
and U16553 (N_16553,N_11625,N_9281);
nand U16554 (N_16554,N_6032,N_9057);
or U16555 (N_16555,N_7355,N_7572);
xor U16556 (N_16556,N_6459,N_6028);
xor U16557 (N_16557,N_11478,N_9827);
nor U16558 (N_16558,N_6210,N_10964);
nor U16559 (N_16559,N_9682,N_9832);
nor U16560 (N_16560,N_10042,N_10320);
xor U16561 (N_16561,N_6196,N_9846);
xnor U16562 (N_16562,N_9658,N_6446);
xor U16563 (N_16563,N_11559,N_8850);
or U16564 (N_16564,N_6896,N_7530);
nand U16565 (N_16565,N_9349,N_7257);
nand U16566 (N_16566,N_10670,N_8749);
or U16567 (N_16567,N_6394,N_8030);
nor U16568 (N_16568,N_9907,N_9033);
or U16569 (N_16569,N_9636,N_7980);
and U16570 (N_16570,N_6716,N_9034);
nor U16571 (N_16571,N_9175,N_11942);
nor U16572 (N_16572,N_9539,N_6121);
nor U16573 (N_16573,N_11304,N_11216);
or U16574 (N_16574,N_6662,N_6219);
nand U16575 (N_16575,N_11176,N_7581);
or U16576 (N_16576,N_11873,N_9887);
and U16577 (N_16577,N_9929,N_8500);
and U16578 (N_16578,N_9756,N_6963);
nor U16579 (N_16579,N_6652,N_9334);
and U16580 (N_16580,N_9620,N_8484);
and U16581 (N_16581,N_9464,N_9416);
nand U16582 (N_16582,N_6473,N_8142);
xor U16583 (N_16583,N_11969,N_9960);
xnor U16584 (N_16584,N_8317,N_6270);
or U16585 (N_16585,N_6217,N_10981);
and U16586 (N_16586,N_7140,N_10683);
nand U16587 (N_16587,N_10721,N_7339);
nor U16588 (N_16588,N_9323,N_9938);
or U16589 (N_16589,N_9968,N_11913);
nor U16590 (N_16590,N_9807,N_10310);
or U16591 (N_16591,N_8940,N_9631);
nor U16592 (N_16592,N_11707,N_11775);
nand U16593 (N_16593,N_6890,N_11189);
nand U16594 (N_16594,N_9188,N_7239);
nor U16595 (N_16595,N_6842,N_9262);
xor U16596 (N_16596,N_10011,N_8368);
nor U16597 (N_16597,N_7447,N_8316);
or U16598 (N_16598,N_8058,N_10698);
or U16599 (N_16599,N_8021,N_9445);
nand U16600 (N_16600,N_10084,N_6896);
xor U16601 (N_16601,N_11032,N_6151);
and U16602 (N_16602,N_8675,N_9341);
and U16603 (N_16603,N_9715,N_8929);
nor U16604 (N_16604,N_8773,N_11479);
nor U16605 (N_16605,N_8626,N_7967);
or U16606 (N_16606,N_7475,N_7396);
or U16607 (N_16607,N_11125,N_8961);
or U16608 (N_16608,N_6027,N_6140);
nor U16609 (N_16609,N_9928,N_9019);
xor U16610 (N_16610,N_7833,N_7584);
xor U16611 (N_16611,N_6252,N_9891);
nand U16612 (N_16612,N_10663,N_8913);
or U16613 (N_16613,N_9363,N_6139);
nor U16614 (N_16614,N_11173,N_11280);
xnor U16615 (N_16615,N_7505,N_6005);
xor U16616 (N_16616,N_6160,N_9098);
or U16617 (N_16617,N_11595,N_10984);
xor U16618 (N_16618,N_6657,N_7382);
and U16619 (N_16619,N_10264,N_11974);
or U16620 (N_16620,N_9803,N_11065);
and U16621 (N_16621,N_7406,N_10804);
nor U16622 (N_16622,N_10515,N_7241);
or U16623 (N_16623,N_7765,N_9226);
or U16624 (N_16624,N_11725,N_9494);
nor U16625 (N_16625,N_8296,N_6220);
nor U16626 (N_16626,N_8353,N_6295);
nand U16627 (N_16627,N_9398,N_8459);
nand U16628 (N_16628,N_7943,N_9646);
or U16629 (N_16629,N_11939,N_7737);
and U16630 (N_16630,N_6762,N_10056);
or U16631 (N_16631,N_9515,N_9421);
nand U16632 (N_16632,N_6676,N_7938);
nor U16633 (N_16633,N_10481,N_7480);
nand U16634 (N_16634,N_6612,N_10731);
and U16635 (N_16635,N_10636,N_10038);
and U16636 (N_16636,N_6260,N_8341);
nor U16637 (N_16637,N_7439,N_11650);
or U16638 (N_16638,N_7209,N_8093);
nor U16639 (N_16639,N_7085,N_10451);
nand U16640 (N_16640,N_7359,N_8779);
and U16641 (N_16641,N_10012,N_8076);
or U16642 (N_16642,N_8597,N_7182);
or U16643 (N_16643,N_6624,N_6475);
nand U16644 (N_16644,N_7957,N_11970);
nor U16645 (N_16645,N_6946,N_6650);
and U16646 (N_16646,N_7160,N_6092);
or U16647 (N_16647,N_8167,N_9868);
and U16648 (N_16648,N_6216,N_11729);
xor U16649 (N_16649,N_6410,N_7550);
nor U16650 (N_16650,N_10618,N_7326);
or U16651 (N_16651,N_10783,N_9014);
and U16652 (N_16652,N_7134,N_7925);
and U16653 (N_16653,N_11599,N_7144);
and U16654 (N_16654,N_9798,N_8836);
xnor U16655 (N_16655,N_10501,N_9598);
and U16656 (N_16656,N_7551,N_10468);
xor U16657 (N_16657,N_7778,N_8155);
and U16658 (N_16658,N_7761,N_9005);
nor U16659 (N_16659,N_10642,N_11787);
and U16660 (N_16660,N_10493,N_10782);
nor U16661 (N_16661,N_9321,N_9187);
xor U16662 (N_16662,N_6803,N_10151);
or U16663 (N_16663,N_6914,N_10963);
nor U16664 (N_16664,N_11773,N_8798);
nand U16665 (N_16665,N_7781,N_8248);
nor U16666 (N_16666,N_6872,N_11885);
nand U16667 (N_16667,N_6645,N_8568);
xnor U16668 (N_16668,N_9687,N_6138);
xor U16669 (N_16669,N_6775,N_8238);
and U16670 (N_16670,N_11358,N_9016);
nor U16671 (N_16671,N_7375,N_7853);
and U16672 (N_16672,N_8188,N_8838);
nand U16673 (N_16673,N_6928,N_11103);
nor U16674 (N_16674,N_8248,N_7736);
nand U16675 (N_16675,N_6260,N_9069);
xor U16676 (N_16676,N_8542,N_9517);
nand U16677 (N_16677,N_11290,N_7322);
xor U16678 (N_16678,N_7752,N_6540);
xnor U16679 (N_16679,N_8334,N_8011);
nand U16680 (N_16680,N_7676,N_9402);
nor U16681 (N_16681,N_7634,N_6697);
and U16682 (N_16682,N_8722,N_8295);
xnor U16683 (N_16683,N_8133,N_6515);
or U16684 (N_16684,N_10915,N_10923);
xor U16685 (N_16685,N_10291,N_9663);
and U16686 (N_16686,N_6981,N_8519);
or U16687 (N_16687,N_7997,N_7825);
nor U16688 (N_16688,N_10035,N_10451);
nand U16689 (N_16689,N_9146,N_10833);
and U16690 (N_16690,N_6604,N_8547);
or U16691 (N_16691,N_8770,N_9385);
xor U16692 (N_16692,N_8092,N_10572);
nand U16693 (N_16693,N_9936,N_11213);
or U16694 (N_16694,N_6070,N_7331);
and U16695 (N_16695,N_8880,N_11281);
and U16696 (N_16696,N_8113,N_10408);
nor U16697 (N_16697,N_11665,N_7731);
nor U16698 (N_16698,N_9035,N_8235);
or U16699 (N_16699,N_7815,N_8088);
or U16700 (N_16700,N_9060,N_10679);
nor U16701 (N_16701,N_11095,N_9602);
and U16702 (N_16702,N_8798,N_8455);
and U16703 (N_16703,N_6633,N_6827);
nand U16704 (N_16704,N_6589,N_10569);
and U16705 (N_16705,N_8037,N_10543);
or U16706 (N_16706,N_7395,N_11556);
nor U16707 (N_16707,N_8017,N_7902);
nor U16708 (N_16708,N_10348,N_7393);
nand U16709 (N_16709,N_8310,N_7297);
or U16710 (N_16710,N_11913,N_10781);
nor U16711 (N_16711,N_11309,N_11750);
nand U16712 (N_16712,N_7055,N_6076);
and U16713 (N_16713,N_6560,N_8803);
nand U16714 (N_16714,N_9006,N_9437);
nand U16715 (N_16715,N_9099,N_8922);
and U16716 (N_16716,N_8136,N_11888);
xnor U16717 (N_16717,N_9303,N_8485);
or U16718 (N_16718,N_7389,N_6488);
or U16719 (N_16719,N_7658,N_9579);
and U16720 (N_16720,N_7766,N_9008);
nor U16721 (N_16721,N_10044,N_9973);
nand U16722 (N_16722,N_6241,N_9390);
xor U16723 (N_16723,N_10386,N_9052);
nand U16724 (N_16724,N_7883,N_8267);
xor U16725 (N_16725,N_10299,N_11877);
xor U16726 (N_16726,N_9974,N_6030);
and U16727 (N_16727,N_8178,N_7384);
nor U16728 (N_16728,N_6058,N_6192);
nand U16729 (N_16729,N_9804,N_8149);
nand U16730 (N_16730,N_10729,N_11350);
nand U16731 (N_16731,N_8742,N_6312);
nor U16732 (N_16732,N_8156,N_8157);
nand U16733 (N_16733,N_11228,N_11604);
and U16734 (N_16734,N_10977,N_11661);
xor U16735 (N_16735,N_9016,N_7330);
or U16736 (N_16736,N_11016,N_9304);
or U16737 (N_16737,N_11618,N_11172);
nor U16738 (N_16738,N_9529,N_10796);
xnor U16739 (N_16739,N_6096,N_6474);
or U16740 (N_16740,N_7999,N_9631);
xnor U16741 (N_16741,N_8851,N_11291);
and U16742 (N_16742,N_9893,N_6574);
or U16743 (N_16743,N_6750,N_7158);
and U16744 (N_16744,N_8355,N_9362);
nand U16745 (N_16745,N_8288,N_8707);
or U16746 (N_16746,N_9053,N_6104);
xor U16747 (N_16747,N_6783,N_8849);
nand U16748 (N_16748,N_6504,N_7289);
or U16749 (N_16749,N_6937,N_10007);
nor U16750 (N_16750,N_7804,N_9887);
nor U16751 (N_16751,N_7933,N_8128);
nor U16752 (N_16752,N_9849,N_7097);
or U16753 (N_16753,N_8910,N_8987);
xnor U16754 (N_16754,N_7922,N_11411);
xnor U16755 (N_16755,N_9485,N_8155);
and U16756 (N_16756,N_6466,N_9293);
or U16757 (N_16757,N_8056,N_9161);
or U16758 (N_16758,N_11298,N_8798);
nand U16759 (N_16759,N_9858,N_9793);
or U16760 (N_16760,N_11489,N_11381);
nor U16761 (N_16761,N_6046,N_11244);
nor U16762 (N_16762,N_11367,N_10636);
and U16763 (N_16763,N_7992,N_9233);
or U16764 (N_16764,N_11249,N_9554);
and U16765 (N_16765,N_10746,N_11959);
nor U16766 (N_16766,N_8952,N_6962);
xnor U16767 (N_16767,N_11421,N_11163);
and U16768 (N_16768,N_11760,N_8943);
xnor U16769 (N_16769,N_6467,N_10669);
nand U16770 (N_16770,N_6185,N_8136);
or U16771 (N_16771,N_7097,N_9807);
nor U16772 (N_16772,N_10872,N_10052);
nor U16773 (N_16773,N_8078,N_10350);
and U16774 (N_16774,N_7157,N_9043);
nor U16775 (N_16775,N_8062,N_7521);
xor U16776 (N_16776,N_7658,N_9943);
or U16777 (N_16777,N_11594,N_7417);
xor U16778 (N_16778,N_8931,N_7096);
nand U16779 (N_16779,N_7030,N_10596);
nor U16780 (N_16780,N_7827,N_9551);
or U16781 (N_16781,N_11515,N_9793);
nand U16782 (N_16782,N_9533,N_11365);
nand U16783 (N_16783,N_6823,N_8554);
nand U16784 (N_16784,N_8382,N_8383);
or U16785 (N_16785,N_8317,N_9223);
and U16786 (N_16786,N_9146,N_7738);
or U16787 (N_16787,N_9047,N_11829);
and U16788 (N_16788,N_8108,N_11386);
and U16789 (N_16789,N_6825,N_10140);
and U16790 (N_16790,N_9787,N_6871);
or U16791 (N_16791,N_10922,N_10973);
and U16792 (N_16792,N_8764,N_7419);
and U16793 (N_16793,N_6976,N_6196);
or U16794 (N_16794,N_10862,N_8250);
and U16795 (N_16795,N_10383,N_10914);
or U16796 (N_16796,N_10407,N_11275);
nand U16797 (N_16797,N_8897,N_9498);
xnor U16798 (N_16798,N_7275,N_10426);
or U16799 (N_16799,N_10389,N_11987);
and U16800 (N_16800,N_8178,N_8479);
and U16801 (N_16801,N_7201,N_7709);
nand U16802 (N_16802,N_11894,N_6514);
and U16803 (N_16803,N_6324,N_8226);
and U16804 (N_16804,N_7053,N_7233);
and U16805 (N_16805,N_10933,N_10536);
nor U16806 (N_16806,N_11893,N_7177);
and U16807 (N_16807,N_6518,N_7834);
nor U16808 (N_16808,N_7911,N_7255);
xnor U16809 (N_16809,N_9050,N_6718);
nand U16810 (N_16810,N_8251,N_10902);
or U16811 (N_16811,N_9788,N_11973);
nor U16812 (N_16812,N_11240,N_9028);
and U16813 (N_16813,N_7003,N_6566);
nor U16814 (N_16814,N_6922,N_11117);
and U16815 (N_16815,N_9325,N_10572);
nor U16816 (N_16816,N_6956,N_7955);
nor U16817 (N_16817,N_11566,N_10557);
xnor U16818 (N_16818,N_11933,N_10785);
or U16819 (N_16819,N_6030,N_10145);
nand U16820 (N_16820,N_8986,N_6364);
nand U16821 (N_16821,N_11449,N_7740);
or U16822 (N_16822,N_11118,N_11746);
nor U16823 (N_16823,N_9769,N_7764);
nor U16824 (N_16824,N_10795,N_8836);
xor U16825 (N_16825,N_6693,N_6191);
nor U16826 (N_16826,N_7814,N_7238);
and U16827 (N_16827,N_7938,N_7931);
xnor U16828 (N_16828,N_7208,N_9081);
and U16829 (N_16829,N_11887,N_9358);
nor U16830 (N_16830,N_10213,N_9288);
nand U16831 (N_16831,N_8701,N_11717);
and U16832 (N_16832,N_8724,N_7837);
nand U16833 (N_16833,N_6270,N_10964);
or U16834 (N_16834,N_11634,N_8857);
or U16835 (N_16835,N_6781,N_11266);
nor U16836 (N_16836,N_7436,N_11768);
or U16837 (N_16837,N_6320,N_7210);
nand U16838 (N_16838,N_7196,N_9437);
xor U16839 (N_16839,N_9462,N_9507);
xnor U16840 (N_16840,N_7170,N_11553);
nor U16841 (N_16841,N_11340,N_9136);
nor U16842 (N_16842,N_9161,N_10295);
nor U16843 (N_16843,N_11835,N_7770);
or U16844 (N_16844,N_6436,N_8289);
or U16845 (N_16845,N_7955,N_8693);
or U16846 (N_16846,N_11654,N_8412);
and U16847 (N_16847,N_10738,N_6919);
xor U16848 (N_16848,N_8628,N_10790);
xor U16849 (N_16849,N_6249,N_6485);
nand U16850 (N_16850,N_11956,N_9488);
nand U16851 (N_16851,N_6323,N_7254);
xor U16852 (N_16852,N_7800,N_7483);
xor U16853 (N_16853,N_10257,N_10277);
nand U16854 (N_16854,N_6749,N_10074);
xnor U16855 (N_16855,N_10909,N_6174);
nor U16856 (N_16856,N_9225,N_7988);
nor U16857 (N_16857,N_11659,N_8260);
or U16858 (N_16858,N_6523,N_8016);
or U16859 (N_16859,N_9239,N_6889);
xor U16860 (N_16860,N_7165,N_7609);
xor U16861 (N_16861,N_9509,N_7706);
nor U16862 (N_16862,N_6535,N_11577);
or U16863 (N_16863,N_6399,N_8753);
or U16864 (N_16864,N_10630,N_8364);
xor U16865 (N_16865,N_9408,N_8201);
and U16866 (N_16866,N_6457,N_8995);
nor U16867 (N_16867,N_8579,N_11642);
or U16868 (N_16868,N_11114,N_11586);
xnor U16869 (N_16869,N_6562,N_10580);
nand U16870 (N_16870,N_9562,N_9383);
nand U16871 (N_16871,N_7264,N_9716);
nor U16872 (N_16872,N_10151,N_11234);
and U16873 (N_16873,N_10358,N_10506);
nand U16874 (N_16874,N_7849,N_10438);
xor U16875 (N_16875,N_8777,N_6572);
xnor U16876 (N_16876,N_9529,N_9510);
nand U16877 (N_16877,N_9916,N_11588);
nand U16878 (N_16878,N_11679,N_10159);
nand U16879 (N_16879,N_6357,N_11799);
and U16880 (N_16880,N_10762,N_8964);
or U16881 (N_16881,N_7188,N_8966);
and U16882 (N_16882,N_7939,N_9821);
xor U16883 (N_16883,N_9935,N_11655);
and U16884 (N_16884,N_9291,N_6099);
nor U16885 (N_16885,N_8145,N_10666);
or U16886 (N_16886,N_10718,N_11345);
and U16887 (N_16887,N_10419,N_8956);
nor U16888 (N_16888,N_8573,N_6546);
or U16889 (N_16889,N_9552,N_9592);
nand U16890 (N_16890,N_8707,N_11404);
or U16891 (N_16891,N_9531,N_11270);
nor U16892 (N_16892,N_6870,N_7845);
and U16893 (N_16893,N_9913,N_7859);
nor U16894 (N_16894,N_9610,N_7082);
nand U16895 (N_16895,N_6433,N_10929);
nand U16896 (N_16896,N_7751,N_7000);
nor U16897 (N_16897,N_10134,N_8230);
nor U16898 (N_16898,N_8775,N_6242);
or U16899 (N_16899,N_9722,N_10887);
nand U16900 (N_16900,N_9074,N_8398);
nor U16901 (N_16901,N_9282,N_9186);
and U16902 (N_16902,N_11755,N_6983);
nand U16903 (N_16903,N_7605,N_8964);
nor U16904 (N_16904,N_10838,N_9849);
and U16905 (N_16905,N_6276,N_11254);
nor U16906 (N_16906,N_10592,N_10231);
xor U16907 (N_16907,N_9930,N_8210);
or U16908 (N_16908,N_9410,N_8631);
and U16909 (N_16909,N_10910,N_7721);
or U16910 (N_16910,N_10950,N_6167);
xor U16911 (N_16911,N_9457,N_11537);
nand U16912 (N_16912,N_6761,N_6022);
nand U16913 (N_16913,N_11826,N_10093);
nor U16914 (N_16914,N_10173,N_10795);
xnor U16915 (N_16915,N_9395,N_7685);
xnor U16916 (N_16916,N_10062,N_10474);
and U16917 (N_16917,N_10130,N_9825);
xnor U16918 (N_16918,N_10397,N_7040);
and U16919 (N_16919,N_10828,N_7246);
and U16920 (N_16920,N_6105,N_7718);
or U16921 (N_16921,N_11780,N_8518);
or U16922 (N_16922,N_8358,N_9371);
nor U16923 (N_16923,N_11057,N_9896);
and U16924 (N_16924,N_11482,N_6688);
nor U16925 (N_16925,N_10239,N_6748);
xnor U16926 (N_16926,N_9490,N_6555);
xor U16927 (N_16927,N_8220,N_11744);
and U16928 (N_16928,N_10056,N_8219);
nor U16929 (N_16929,N_9493,N_7061);
and U16930 (N_16930,N_10292,N_10867);
and U16931 (N_16931,N_9925,N_8504);
nor U16932 (N_16932,N_10122,N_11409);
and U16933 (N_16933,N_11990,N_7121);
nor U16934 (N_16934,N_8605,N_7810);
nor U16935 (N_16935,N_9988,N_6445);
or U16936 (N_16936,N_9108,N_6664);
nor U16937 (N_16937,N_10084,N_8300);
nand U16938 (N_16938,N_8440,N_7307);
and U16939 (N_16939,N_10678,N_7590);
or U16940 (N_16940,N_9681,N_10231);
nand U16941 (N_16941,N_8753,N_6169);
nand U16942 (N_16942,N_6833,N_10563);
and U16943 (N_16943,N_11596,N_9655);
or U16944 (N_16944,N_9538,N_10703);
or U16945 (N_16945,N_7606,N_9137);
and U16946 (N_16946,N_11945,N_11776);
xnor U16947 (N_16947,N_10045,N_9978);
xor U16948 (N_16948,N_11904,N_8612);
and U16949 (N_16949,N_6213,N_9519);
or U16950 (N_16950,N_7966,N_8106);
xnor U16951 (N_16951,N_6139,N_7785);
xnor U16952 (N_16952,N_7410,N_7007);
nor U16953 (N_16953,N_7405,N_9155);
nor U16954 (N_16954,N_7545,N_7729);
or U16955 (N_16955,N_8162,N_6484);
and U16956 (N_16956,N_6636,N_6075);
nor U16957 (N_16957,N_8472,N_6937);
or U16958 (N_16958,N_9241,N_6731);
xnor U16959 (N_16959,N_11799,N_6006);
and U16960 (N_16960,N_8322,N_9252);
and U16961 (N_16961,N_7127,N_8885);
nor U16962 (N_16962,N_11984,N_7142);
xor U16963 (N_16963,N_6355,N_7098);
nand U16964 (N_16964,N_6217,N_10948);
nand U16965 (N_16965,N_9386,N_9798);
xor U16966 (N_16966,N_7865,N_11265);
nor U16967 (N_16967,N_6531,N_8469);
and U16968 (N_16968,N_9405,N_7613);
nand U16969 (N_16969,N_10009,N_9294);
and U16970 (N_16970,N_10362,N_11116);
or U16971 (N_16971,N_8324,N_7716);
nor U16972 (N_16972,N_6579,N_9536);
nand U16973 (N_16973,N_11162,N_9312);
nor U16974 (N_16974,N_10372,N_9224);
or U16975 (N_16975,N_8732,N_6338);
and U16976 (N_16976,N_8479,N_8271);
or U16977 (N_16977,N_7781,N_11654);
xor U16978 (N_16978,N_11397,N_7676);
and U16979 (N_16979,N_6732,N_6248);
nand U16980 (N_16980,N_10776,N_11298);
or U16981 (N_16981,N_7080,N_8163);
or U16982 (N_16982,N_7129,N_7016);
or U16983 (N_16983,N_8722,N_9544);
and U16984 (N_16984,N_9852,N_6315);
xor U16985 (N_16985,N_8140,N_10965);
and U16986 (N_16986,N_10824,N_10292);
and U16987 (N_16987,N_10499,N_8504);
xor U16988 (N_16988,N_7882,N_6973);
and U16989 (N_16989,N_10720,N_9064);
or U16990 (N_16990,N_8081,N_9551);
or U16991 (N_16991,N_10978,N_9345);
xnor U16992 (N_16992,N_9922,N_7796);
and U16993 (N_16993,N_11339,N_7022);
xnor U16994 (N_16994,N_7043,N_8247);
or U16995 (N_16995,N_10100,N_6272);
or U16996 (N_16996,N_8886,N_10678);
nor U16997 (N_16997,N_6222,N_6613);
and U16998 (N_16998,N_10763,N_10767);
nand U16999 (N_16999,N_8839,N_9902);
or U17000 (N_17000,N_11415,N_11617);
or U17001 (N_17001,N_11544,N_6838);
or U17002 (N_17002,N_9474,N_6489);
xnor U17003 (N_17003,N_11682,N_7481);
nor U17004 (N_17004,N_10179,N_7491);
nor U17005 (N_17005,N_6175,N_8792);
xnor U17006 (N_17006,N_10371,N_8312);
nor U17007 (N_17007,N_10090,N_10042);
or U17008 (N_17008,N_10256,N_7805);
xnor U17009 (N_17009,N_7451,N_11475);
and U17010 (N_17010,N_10565,N_8414);
nor U17011 (N_17011,N_8252,N_10916);
nor U17012 (N_17012,N_10754,N_10098);
nand U17013 (N_17013,N_10344,N_6919);
and U17014 (N_17014,N_11900,N_11653);
xnor U17015 (N_17015,N_7367,N_10129);
xor U17016 (N_17016,N_7095,N_7730);
nand U17017 (N_17017,N_9009,N_7704);
nor U17018 (N_17018,N_9230,N_7152);
and U17019 (N_17019,N_8431,N_6982);
nand U17020 (N_17020,N_8529,N_10275);
xor U17021 (N_17021,N_8725,N_9553);
or U17022 (N_17022,N_11170,N_11525);
nand U17023 (N_17023,N_8329,N_11408);
or U17024 (N_17024,N_11380,N_11411);
xnor U17025 (N_17025,N_11736,N_8785);
xnor U17026 (N_17026,N_11623,N_10681);
nand U17027 (N_17027,N_9513,N_7331);
and U17028 (N_17028,N_10717,N_6047);
or U17029 (N_17029,N_7702,N_8704);
or U17030 (N_17030,N_8502,N_9646);
or U17031 (N_17031,N_7102,N_8083);
xnor U17032 (N_17032,N_6876,N_8634);
nand U17033 (N_17033,N_9468,N_6379);
xnor U17034 (N_17034,N_8108,N_11755);
nor U17035 (N_17035,N_10257,N_8470);
nor U17036 (N_17036,N_8106,N_10627);
or U17037 (N_17037,N_8431,N_8028);
and U17038 (N_17038,N_8185,N_10897);
or U17039 (N_17039,N_9874,N_6962);
or U17040 (N_17040,N_11494,N_9821);
and U17041 (N_17041,N_7025,N_11402);
nor U17042 (N_17042,N_6814,N_8315);
nand U17043 (N_17043,N_11320,N_9702);
and U17044 (N_17044,N_11884,N_9705);
nand U17045 (N_17045,N_8056,N_6072);
nor U17046 (N_17046,N_9652,N_6105);
nor U17047 (N_17047,N_7657,N_8850);
nor U17048 (N_17048,N_8259,N_9161);
xor U17049 (N_17049,N_8575,N_9050);
nor U17050 (N_17050,N_6431,N_7796);
nor U17051 (N_17051,N_11159,N_6596);
or U17052 (N_17052,N_10856,N_11293);
or U17053 (N_17053,N_11411,N_10438);
xor U17054 (N_17054,N_11768,N_10206);
nand U17055 (N_17055,N_7875,N_9427);
or U17056 (N_17056,N_6742,N_7573);
or U17057 (N_17057,N_11953,N_6031);
nor U17058 (N_17058,N_7562,N_9833);
nand U17059 (N_17059,N_6362,N_9677);
or U17060 (N_17060,N_7795,N_8197);
nand U17061 (N_17061,N_6615,N_6382);
nand U17062 (N_17062,N_9680,N_6705);
or U17063 (N_17063,N_10742,N_10912);
and U17064 (N_17064,N_8003,N_8271);
and U17065 (N_17065,N_9638,N_11398);
nor U17066 (N_17066,N_9249,N_6950);
or U17067 (N_17067,N_11326,N_7480);
and U17068 (N_17068,N_10650,N_11680);
and U17069 (N_17069,N_6292,N_7289);
nor U17070 (N_17070,N_7410,N_10543);
and U17071 (N_17071,N_11795,N_6528);
or U17072 (N_17072,N_9575,N_8305);
or U17073 (N_17073,N_10487,N_8760);
nor U17074 (N_17074,N_9084,N_10513);
and U17075 (N_17075,N_11998,N_9917);
nand U17076 (N_17076,N_9790,N_6586);
and U17077 (N_17077,N_11522,N_11178);
and U17078 (N_17078,N_11393,N_7184);
or U17079 (N_17079,N_11292,N_7892);
nor U17080 (N_17080,N_11869,N_8552);
xnor U17081 (N_17081,N_9785,N_6279);
or U17082 (N_17082,N_9606,N_9131);
xnor U17083 (N_17083,N_7622,N_8647);
xor U17084 (N_17084,N_7932,N_9292);
or U17085 (N_17085,N_10927,N_6391);
xor U17086 (N_17086,N_11649,N_9930);
nand U17087 (N_17087,N_9428,N_7318);
nor U17088 (N_17088,N_7740,N_6396);
and U17089 (N_17089,N_10811,N_6753);
or U17090 (N_17090,N_10875,N_9629);
nor U17091 (N_17091,N_9206,N_6139);
or U17092 (N_17092,N_6489,N_7419);
or U17093 (N_17093,N_10327,N_9459);
nand U17094 (N_17094,N_10521,N_7119);
nand U17095 (N_17095,N_6398,N_8903);
and U17096 (N_17096,N_9338,N_11392);
or U17097 (N_17097,N_6586,N_9516);
nor U17098 (N_17098,N_9312,N_9118);
xnor U17099 (N_17099,N_10472,N_11725);
nor U17100 (N_17100,N_11581,N_6166);
xnor U17101 (N_17101,N_6636,N_7829);
or U17102 (N_17102,N_6739,N_8965);
and U17103 (N_17103,N_10705,N_9700);
nor U17104 (N_17104,N_7037,N_11703);
nand U17105 (N_17105,N_9893,N_11191);
and U17106 (N_17106,N_9634,N_11820);
nand U17107 (N_17107,N_8985,N_7612);
nand U17108 (N_17108,N_6658,N_11531);
and U17109 (N_17109,N_10783,N_8588);
and U17110 (N_17110,N_10901,N_8963);
nand U17111 (N_17111,N_7826,N_11463);
and U17112 (N_17112,N_9274,N_11489);
nor U17113 (N_17113,N_7098,N_7761);
xnor U17114 (N_17114,N_6944,N_10680);
nand U17115 (N_17115,N_7350,N_10860);
xor U17116 (N_17116,N_9464,N_7504);
or U17117 (N_17117,N_10329,N_10080);
xor U17118 (N_17118,N_10079,N_10434);
and U17119 (N_17119,N_11084,N_8221);
nand U17120 (N_17120,N_8953,N_7377);
nand U17121 (N_17121,N_10745,N_11976);
xnor U17122 (N_17122,N_7611,N_8629);
xor U17123 (N_17123,N_9081,N_6608);
nand U17124 (N_17124,N_7718,N_10825);
nand U17125 (N_17125,N_11783,N_11892);
nor U17126 (N_17126,N_11607,N_10712);
nand U17127 (N_17127,N_6427,N_9146);
xnor U17128 (N_17128,N_11620,N_7942);
xnor U17129 (N_17129,N_10183,N_9527);
nor U17130 (N_17130,N_11037,N_6811);
or U17131 (N_17131,N_8593,N_10300);
xnor U17132 (N_17132,N_11412,N_8940);
nand U17133 (N_17133,N_8095,N_10825);
or U17134 (N_17134,N_10232,N_8889);
or U17135 (N_17135,N_7071,N_7304);
xor U17136 (N_17136,N_7855,N_8495);
xnor U17137 (N_17137,N_7128,N_6960);
and U17138 (N_17138,N_11954,N_7062);
nand U17139 (N_17139,N_6488,N_6702);
or U17140 (N_17140,N_6345,N_8535);
xnor U17141 (N_17141,N_9641,N_6230);
or U17142 (N_17142,N_9135,N_11984);
and U17143 (N_17143,N_11950,N_8007);
nor U17144 (N_17144,N_11486,N_7846);
nand U17145 (N_17145,N_10005,N_8860);
nand U17146 (N_17146,N_6716,N_11243);
nor U17147 (N_17147,N_10936,N_10702);
xnor U17148 (N_17148,N_7435,N_6356);
nor U17149 (N_17149,N_7801,N_7476);
nor U17150 (N_17150,N_10575,N_6439);
xor U17151 (N_17151,N_10379,N_8967);
and U17152 (N_17152,N_6399,N_6009);
nor U17153 (N_17153,N_6652,N_9090);
nand U17154 (N_17154,N_11727,N_11554);
nor U17155 (N_17155,N_8560,N_9101);
nor U17156 (N_17156,N_10227,N_6159);
nand U17157 (N_17157,N_6497,N_9184);
and U17158 (N_17158,N_8348,N_7761);
or U17159 (N_17159,N_11999,N_8000);
or U17160 (N_17160,N_9132,N_7843);
xnor U17161 (N_17161,N_7404,N_11396);
nand U17162 (N_17162,N_7117,N_6716);
nor U17163 (N_17163,N_9317,N_6191);
and U17164 (N_17164,N_8096,N_11680);
or U17165 (N_17165,N_8860,N_6242);
and U17166 (N_17166,N_7558,N_6115);
and U17167 (N_17167,N_7813,N_10299);
or U17168 (N_17168,N_8793,N_11959);
xnor U17169 (N_17169,N_10184,N_9180);
xor U17170 (N_17170,N_6285,N_11638);
xor U17171 (N_17171,N_10499,N_10566);
nor U17172 (N_17172,N_10180,N_6888);
or U17173 (N_17173,N_9273,N_10158);
and U17174 (N_17174,N_6733,N_10882);
and U17175 (N_17175,N_8194,N_10345);
and U17176 (N_17176,N_10079,N_10287);
nor U17177 (N_17177,N_9822,N_8206);
nand U17178 (N_17178,N_7800,N_7790);
and U17179 (N_17179,N_7417,N_11877);
nand U17180 (N_17180,N_6267,N_10148);
nand U17181 (N_17181,N_6625,N_10291);
xor U17182 (N_17182,N_10929,N_10410);
or U17183 (N_17183,N_6039,N_8848);
xor U17184 (N_17184,N_7815,N_11290);
nand U17185 (N_17185,N_7201,N_7309);
xnor U17186 (N_17186,N_6625,N_10250);
or U17187 (N_17187,N_11676,N_8278);
xnor U17188 (N_17188,N_9072,N_7096);
xor U17189 (N_17189,N_9069,N_6115);
and U17190 (N_17190,N_11004,N_10436);
nand U17191 (N_17191,N_11065,N_6884);
nor U17192 (N_17192,N_8267,N_6521);
nor U17193 (N_17193,N_8884,N_11726);
and U17194 (N_17194,N_9076,N_7569);
xnor U17195 (N_17195,N_7381,N_9354);
nand U17196 (N_17196,N_10083,N_11869);
nor U17197 (N_17197,N_8833,N_6251);
nor U17198 (N_17198,N_9383,N_7323);
xor U17199 (N_17199,N_10829,N_7713);
nor U17200 (N_17200,N_11139,N_10498);
nand U17201 (N_17201,N_11692,N_7080);
or U17202 (N_17202,N_7944,N_7031);
or U17203 (N_17203,N_9546,N_9616);
nor U17204 (N_17204,N_8683,N_9380);
and U17205 (N_17205,N_7223,N_10338);
xnor U17206 (N_17206,N_10124,N_10427);
and U17207 (N_17207,N_6415,N_7039);
or U17208 (N_17208,N_8867,N_6919);
or U17209 (N_17209,N_10365,N_7027);
or U17210 (N_17210,N_9972,N_6747);
or U17211 (N_17211,N_6841,N_6443);
xor U17212 (N_17212,N_10171,N_7715);
xor U17213 (N_17213,N_6808,N_7110);
nor U17214 (N_17214,N_6053,N_6037);
and U17215 (N_17215,N_9076,N_8869);
and U17216 (N_17216,N_7473,N_11991);
and U17217 (N_17217,N_10164,N_10060);
nor U17218 (N_17218,N_9525,N_8102);
and U17219 (N_17219,N_10432,N_6788);
and U17220 (N_17220,N_10749,N_9252);
or U17221 (N_17221,N_6124,N_10458);
xor U17222 (N_17222,N_9227,N_6536);
or U17223 (N_17223,N_6650,N_6320);
or U17224 (N_17224,N_7749,N_9150);
nor U17225 (N_17225,N_10265,N_8304);
nand U17226 (N_17226,N_6510,N_7362);
and U17227 (N_17227,N_11806,N_10772);
nor U17228 (N_17228,N_8687,N_11436);
nor U17229 (N_17229,N_9313,N_9553);
nor U17230 (N_17230,N_11217,N_6693);
or U17231 (N_17231,N_7333,N_10596);
nor U17232 (N_17232,N_8527,N_6676);
or U17233 (N_17233,N_10163,N_6676);
or U17234 (N_17234,N_7070,N_10913);
and U17235 (N_17235,N_6948,N_9861);
and U17236 (N_17236,N_9448,N_6036);
nor U17237 (N_17237,N_9579,N_10845);
and U17238 (N_17238,N_7848,N_9338);
xnor U17239 (N_17239,N_7169,N_11611);
xnor U17240 (N_17240,N_8792,N_9577);
xor U17241 (N_17241,N_10887,N_11621);
or U17242 (N_17242,N_9822,N_11924);
or U17243 (N_17243,N_10423,N_6002);
nor U17244 (N_17244,N_11461,N_6528);
nor U17245 (N_17245,N_11751,N_10554);
or U17246 (N_17246,N_6196,N_7461);
or U17247 (N_17247,N_7019,N_9718);
xnor U17248 (N_17248,N_6350,N_6128);
nand U17249 (N_17249,N_8041,N_6118);
xor U17250 (N_17250,N_8750,N_11269);
nand U17251 (N_17251,N_8102,N_8516);
nand U17252 (N_17252,N_9592,N_11084);
nor U17253 (N_17253,N_7495,N_9895);
xnor U17254 (N_17254,N_9049,N_11781);
nand U17255 (N_17255,N_8554,N_7213);
nand U17256 (N_17256,N_7879,N_11905);
nand U17257 (N_17257,N_8569,N_7061);
or U17258 (N_17258,N_11253,N_6405);
or U17259 (N_17259,N_11683,N_11439);
and U17260 (N_17260,N_6973,N_7639);
and U17261 (N_17261,N_6763,N_9927);
xor U17262 (N_17262,N_10749,N_10556);
nor U17263 (N_17263,N_10231,N_10992);
xor U17264 (N_17264,N_11019,N_9898);
or U17265 (N_17265,N_7503,N_7774);
nor U17266 (N_17266,N_9416,N_6200);
xor U17267 (N_17267,N_10201,N_11697);
xor U17268 (N_17268,N_6539,N_11700);
or U17269 (N_17269,N_10571,N_6294);
nand U17270 (N_17270,N_11869,N_9059);
and U17271 (N_17271,N_8512,N_10280);
nor U17272 (N_17272,N_10091,N_11664);
xor U17273 (N_17273,N_9623,N_6453);
xnor U17274 (N_17274,N_9611,N_10986);
or U17275 (N_17275,N_7551,N_6039);
or U17276 (N_17276,N_10923,N_8229);
xor U17277 (N_17277,N_6950,N_9250);
nand U17278 (N_17278,N_8220,N_8769);
nor U17279 (N_17279,N_7687,N_6458);
xnor U17280 (N_17280,N_9626,N_6688);
nand U17281 (N_17281,N_11804,N_6702);
nor U17282 (N_17282,N_11153,N_7758);
xor U17283 (N_17283,N_6325,N_8303);
nand U17284 (N_17284,N_7312,N_9547);
nor U17285 (N_17285,N_10154,N_7676);
and U17286 (N_17286,N_9582,N_9876);
and U17287 (N_17287,N_7786,N_11252);
xnor U17288 (N_17288,N_10086,N_9469);
or U17289 (N_17289,N_6419,N_8161);
nor U17290 (N_17290,N_9091,N_11833);
or U17291 (N_17291,N_7117,N_6547);
or U17292 (N_17292,N_9006,N_11097);
and U17293 (N_17293,N_8992,N_7597);
xor U17294 (N_17294,N_9296,N_10364);
and U17295 (N_17295,N_6689,N_11459);
nor U17296 (N_17296,N_9346,N_6923);
xor U17297 (N_17297,N_6409,N_10388);
xnor U17298 (N_17298,N_11159,N_7636);
nand U17299 (N_17299,N_7251,N_10050);
or U17300 (N_17300,N_8766,N_7495);
nand U17301 (N_17301,N_10362,N_11587);
nand U17302 (N_17302,N_11639,N_6313);
xnor U17303 (N_17303,N_8849,N_11851);
nand U17304 (N_17304,N_9691,N_6789);
xor U17305 (N_17305,N_7088,N_9322);
nand U17306 (N_17306,N_7284,N_8605);
nand U17307 (N_17307,N_8273,N_6214);
nor U17308 (N_17308,N_7849,N_10746);
xor U17309 (N_17309,N_9766,N_9504);
nand U17310 (N_17310,N_10147,N_9277);
or U17311 (N_17311,N_7930,N_10334);
nand U17312 (N_17312,N_6017,N_9961);
or U17313 (N_17313,N_8402,N_7863);
nand U17314 (N_17314,N_7292,N_8224);
nand U17315 (N_17315,N_6508,N_8545);
and U17316 (N_17316,N_9815,N_8230);
xnor U17317 (N_17317,N_9288,N_11008);
xnor U17318 (N_17318,N_6788,N_7350);
and U17319 (N_17319,N_7817,N_8884);
nor U17320 (N_17320,N_10548,N_11957);
or U17321 (N_17321,N_9660,N_11751);
and U17322 (N_17322,N_8149,N_8484);
nand U17323 (N_17323,N_7024,N_9429);
nor U17324 (N_17324,N_9123,N_9848);
xnor U17325 (N_17325,N_11644,N_8951);
and U17326 (N_17326,N_9376,N_9745);
nor U17327 (N_17327,N_9937,N_11525);
xnor U17328 (N_17328,N_11455,N_10890);
or U17329 (N_17329,N_9543,N_11992);
xor U17330 (N_17330,N_8382,N_10110);
and U17331 (N_17331,N_10449,N_8830);
and U17332 (N_17332,N_11275,N_10361);
xnor U17333 (N_17333,N_8010,N_11614);
or U17334 (N_17334,N_11015,N_10412);
or U17335 (N_17335,N_6391,N_6268);
nand U17336 (N_17336,N_11368,N_8860);
and U17337 (N_17337,N_7810,N_9351);
nor U17338 (N_17338,N_6536,N_8642);
nor U17339 (N_17339,N_11952,N_10681);
xor U17340 (N_17340,N_10640,N_8900);
nor U17341 (N_17341,N_8070,N_10586);
nor U17342 (N_17342,N_8416,N_6207);
nor U17343 (N_17343,N_7734,N_7014);
nor U17344 (N_17344,N_7274,N_9037);
and U17345 (N_17345,N_10176,N_8637);
nand U17346 (N_17346,N_11320,N_8947);
nor U17347 (N_17347,N_9860,N_11343);
and U17348 (N_17348,N_9215,N_9406);
and U17349 (N_17349,N_6924,N_6312);
or U17350 (N_17350,N_7280,N_9544);
or U17351 (N_17351,N_7212,N_10982);
or U17352 (N_17352,N_9966,N_7454);
or U17353 (N_17353,N_7890,N_10516);
nand U17354 (N_17354,N_8640,N_7822);
nor U17355 (N_17355,N_10286,N_6459);
and U17356 (N_17356,N_8224,N_10472);
nand U17357 (N_17357,N_10643,N_9325);
and U17358 (N_17358,N_7123,N_9873);
nor U17359 (N_17359,N_10909,N_8513);
xnor U17360 (N_17360,N_9540,N_11390);
or U17361 (N_17361,N_11068,N_8991);
xor U17362 (N_17362,N_10005,N_11026);
nor U17363 (N_17363,N_8338,N_9228);
or U17364 (N_17364,N_9264,N_8620);
or U17365 (N_17365,N_6067,N_10511);
xnor U17366 (N_17366,N_10075,N_7305);
xnor U17367 (N_17367,N_8000,N_6779);
and U17368 (N_17368,N_9830,N_8560);
and U17369 (N_17369,N_9102,N_9475);
nor U17370 (N_17370,N_9193,N_7568);
or U17371 (N_17371,N_11404,N_8237);
nor U17372 (N_17372,N_11400,N_10551);
and U17373 (N_17373,N_8911,N_6722);
xnor U17374 (N_17374,N_8703,N_6473);
or U17375 (N_17375,N_11941,N_11282);
or U17376 (N_17376,N_6224,N_6102);
or U17377 (N_17377,N_11050,N_8312);
nand U17378 (N_17378,N_6762,N_10215);
or U17379 (N_17379,N_6862,N_9986);
and U17380 (N_17380,N_7252,N_9628);
xor U17381 (N_17381,N_6392,N_10633);
nor U17382 (N_17382,N_7232,N_10465);
nand U17383 (N_17383,N_8129,N_11204);
xor U17384 (N_17384,N_6290,N_7665);
xnor U17385 (N_17385,N_7375,N_9448);
xnor U17386 (N_17386,N_7672,N_10817);
xor U17387 (N_17387,N_7133,N_11901);
or U17388 (N_17388,N_9104,N_8546);
nand U17389 (N_17389,N_7600,N_11703);
or U17390 (N_17390,N_11096,N_8028);
xor U17391 (N_17391,N_8704,N_6111);
and U17392 (N_17392,N_11575,N_6389);
xnor U17393 (N_17393,N_9277,N_10709);
nor U17394 (N_17394,N_6385,N_9215);
nand U17395 (N_17395,N_8252,N_8354);
xor U17396 (N_17396,N_9078,N_7476);
nand U17397 (N_17397,N_9413,N_6407);
xnor U17398 (N_17398,N_10857,N_9509);
nand U17399 (N_17399,N_6668,N_8173);
nor U17400 (N_17400,N_7800,N_8388);
nor U17401 (N_17401,N_11280,N_6475);
xor U17402 (N_17402,N_10795,N_8339);
xor U17403 (N_17403,N_10065,N_6061);
or U17404 (N_17404,N_9392,N_10634);
or U17405 (N_17405,N_9334,N_10695);
and U17406 (N_17406,N_8849,N_7988);
nand U17407 (N_17407,N_11726,N_8252);
nand U17408 (N_17408,N_11773,N_10096);
xor U17409 (N_17409,N_9741,N_10150);
nor U17410 (N_17410,N_6786,N_10780);
nand U17411 (N_17411,N_10708,N_7494);
xnor U17412 (N_17412,N_10772,N_9096);
nor U17413 (N_17413,N_7517,N_7806);
xor U17414 (N_17414,N_11973,N_10333);
xor U17415 (N_17415,N_8665,N_11844);
xor U17416 (N_17416,N_10576,N_11878);
nor U17417 (N_17417,N_10303,N_10572);
nor U17418 (N_17418,N_9752,N_8520);
nor U17419 (N_17419,N_7521,N_10712);
xor U17420 (N_17420,N_10585,N_9200);
nor U17421 (N_17421,N_11155,N_11590);
nand U17422 (N_17422,N_7465,N_6630);
nor U17423 (N_17423,N_9317,N_9127);
and U17424 (N_17424,N_7108,N_10458);
nand U17425 (N_17425,N_10623,N_7847);
xor U17426 (N_17426,N_10979,N_7055);
nand U17427 (N_17427,N_6970,N_9608);
xnor U17428 (N_17428,N_10537,N_7913);
nor U17429 (N_17429,N_7720,N_9113);
nand U17430 (N_17430,N_10689,N_7655);
xnor U17431 (N_17431,N_7389,N_7699);
nor U17432 (N_17432,N_10813,N_10784);
and U17433 (N_17433,N_11188,N_10715);
nor U17434 (N_17434,N_10532,N_6246);
nand U17435 (N_17435,N_9429,N_6923);
or U17436 (N_17436,N_10366,N_6096);
and U17437 (N_17437,N_7323,N_11597);
and U17438 (N_17438,N_11921,N_6284);
and U17439 (N_17439,N_11262,N_7376);
or U17440 (N_17440,N_8974,N_6135);
nor U17441 (N_17441,N_11096,N_7064);
xor U17442 (N_17442,N_7094,N_9859);
xor U17443 (N_17443,N_10952,N_11464);
nor U17444 (N_17444,N_6012,N_6164);
nor U17445 (N_17445,N_7646,N_10053);
xor U17446 (N_17446,N_6518,N_9034);
and U17447 (N_17447,N_6396,N_8816);
nand U17448 (N_17448,N_7760,N_8501);
xor U17449 (N_17449,N_9358,N_11538);
and U17450 (N_17450,N_10392,N_10396);
and U17451 (N_17451,N_9803,N_11249);
and U17452 (N_17452,N_6138,N_11446);
nand U17453 (N_17453,N_11999,N_9114);
or U17454 (N_17454,N_6619,N_8235);
or U17455 (N_17455,N_9250,N_7059);
xnor U17456 (N_17456,N_8216,N_10102);
xor U17457 (N_17457,N_11067,N_8441);
nor U17458 (N_17458,N_10447,N_11513);
nand U17459 (N_17459,N_6593,N_10613);
xnor U17460 (N_17460,N_9222,N_9657);
or U17461 (N_17461,N_9777,N_7234);
nand U17462 (N_17462,N_10253,N_11610);
and U17463 (N_17463,N_10633,N_11799);
xnor U17464 (N_17464,N_7761,N_10130);
nor U17465 (N_17465,N_11024,N_8999);
nor U17466 (N_17466,N_10186,N_9357);
xor U17467 (N_17467,N_9468,N_7658);
or U17468 (N_17468,N_11041,N_8607);
or U17469 (N_17469,N_6329,N_11429);
nand U17470 (N_17470,N_6932,N_6856);
xor U17471 (N_17471,N_11212,N_8640);
nor U17472 (N_17472,N_7895,N_7786);
xor U17473 (N_17473,N_11748,N_7087);
nand U17474 (N_17474,N_9939,N_11939);
nand U17475 (N_17475,N_8875,N_6823);
xnor U17476 (N_17476,N_11344,N_8759);
xnor U17477 (N_17477,N_10985,N_10932);
nand U17478 (N_17478,N_7089,N_6006);
and U17479 (N_17479,N_9267,N_7260);
or U17480 (N_17480,N_9476,N_7183);
nor U17481 (N_17481,N_8845,N_10204);
or U17482 (N_17482,N_11205,N_10488);
and U17483 (N_17483,N_7210,N_7426);
nand U17484 (N_17484,N_11157,N_11610);
or U17485 (N_17485,N_9996,N_11214);
and U17486 (N_17486,N_11199,N_9707);
or U17487 (N_17487,N_8838,N_7594);
or U17488 (N_17488,N_11271,N_7785);
nand U17489 (N_17489,N_8864,N_11726);
and U17490 (N_17490,N_6951,N_8893);
or U17491 (N_17491,N_8147,N_11807);
xor U17492 (N_17492,N_10367,N_6603);
xnor U17493 (N_17493,N_8617,N_6665);
nor U17494 (N_17494,N_8073,N_11592);
xor U17495 (N_17495,N_11123,N_7675);
xor U17496 (N_17496,N_10479,N_7791);
xnor U17497 (N_17497,N_6006,N_9444);
and U17498 (N_17498,N_9616,N_7568);
nand U17499 (N_17499,N_11043,N_6340);
xnor U17500 (N_17500,N_8719,N_9568);
nor U17501 (N_17501,N_8207,N_7613);
xnor U17502 (N_17502,N_8143,N_9753);
and U17503 (N_17503,N_9106,N_10894);
xnor U17504 (N_17504,N_8513,N_6828);
nand U17505 (N_17505,N_6934,N_10369);
or U17506 (N_17506,N_11780,N_8741);
or U17507 (N_17507,N_7696,N_8519);
or U17508 (N_17508,N_11298,N_6859);
and U17509 (N_17509,N_6976,N_6949);
nor U17510 (N_17510,N_7199,N_6027);
nor U17511 (N_17511,N_6664,N_11850);
nor U17512 (N_17512,N_6065,N_11060);
nand U17513 (N_17513,N_10892,N_6027);
nor U17514 (N_17514,N_6739,N_7334);
nand U17515 (N_17515,N_8031,N_11387);
nand U17516 (N_17516,N_6833,N_10448);
or U17517 (N_17517,N_6199,N_6870);
xor U17518 (N_17518,N_9352,N_10243);
or U17519 (N_17519,N_10619,N_6718);
and U17520 (N_17520,N_11434,N_10030);
or U17521 (N_17521,N_11471,N_9440);
nand U17522 (N_17522,N_8363,N_8907);
nor U17523 (N_17523,N_11416,N_8849);
or U17524 (N_17524,N_8978,N_6599);
nor U17525 (N_17525,N_8268,N_9563);
nor U17526 (N_17526,N_6327,N_8276);
or U17527 (N_17527,N_7595,N_9519);
nor U17528 (N_17528,N_10478,N_9195);
xnor U17529 (N_17529,N_9461,N_8030);
or U17530 (N_17530,N_7450,N_9298);
nand U17531 (N_17531,N_7612,N_7108);
and U17532 (N_17532,N_8800,N_11082);
or U17533 (N_17533,N_10648,N_8073);
xnor U17534 (N_17534,N_6323,N_7659);
nand U17535 (N_17535,N_11679,N_7136);
nand U17536 (N_17536,N_10262,N_9965);
nor U17537 (N_17537,N_7066,N_8579);
or U17538 (N_17538,N_7965,N_9878);
nor U17539 (N_17539,N_7169,N_6909);
and U17540 (N_17540,N_11034,N_11027);
xor U17541 (N_17541,N_7343,N_6568);
or U17542 (N_17542,N_10618,N_11311);
and U17543 (N_17543,N_11830,N_7974);
nor U17544 (N_17544,N_7940,N_6728);
and U17545 (N_17545,N_11273,N_8813);
nor U17546 (N_17546,N_6276,N_6880);
and U17547 (N_17547,N_6067,N_6659);
and U17548 (N_17548,N_9778,N_11969);
or U17549 (N_17549,N_11492,N_7784);
and U17550 (N_17550,N_11927,N_10936);
nor U17551 (N_17551,N_9739,N_6534);
nor U17552 (N_17552,N_6842,N_9673);
xor U17553 (N_17553,N_7215,N_11800);
xor U17554 (N_17554,N_8204,N_7077);
xnor U17555 (N_17555,N_10391,N_9700);
nor U17556 (N_17556,N_8630,N_9870);
xor U17557 (N_17557,N_8479,N_9297);
or U17558 (N_17558,N_7932,N_7409);
nand U17559 (N_17559,N_7518,N_7334);
nor U17560 (N_17560,N_6154,N_10885);
and U17561 (N_17561,N_6003,N_11098);
nor U17562 (N_17562,N_6405,N_10442);
and U17563 (N_17563,N_10669,N_8971);
nor U17564 (N_17564,N_8944,N_10660);
and U17565 (N_17565,N_7557,N_8772);
and U17566 (N_17566,N_8708,N_9276);
and U17567 (N_17567,N_6380,N_9102);
or U17568 (N_17568,N_9723,N_8021);
xor U17569 (N_17569,N_11892,N_11916);
xor U17570 (N_17570,N_9110,N_6119);
xor U17571 (N_17571,N_10650,N_11760);
nand U17572 (N_17572,N_6091,N_7994);
xor U17573 (N_17573,N_6597,N_6648);
nand U17574 (N_17574,N_9818,N_6237);
or U17575 (N_17575,N_9354,N_6049);
xnor U17576 (N_17576,N_10795,N_6114);
nand U17577 (N_17577,N_9219,N_11928);
and U17578 (N_17578,N_10955,N_9496);
and U17579 (N_17579,N_8890,N_9480);
nand U17580 (N_17580,N_8786,N_11700);
xnor U17581 (N_17581,N_11215,N_10591);
nand U17582 (N_17582,N_8073,N_10436);
or U17583 (N_17583,N_9112,N_6931);
nor U17584 (N_17584,N_8563,N_7852);
xor U17585 (N_17585,N_11598,N_9041);
and U17586 (N_17586,N_11913,N_11187);
nor U17587 (N_17587,N_8578,N_7446);
nor U17588 (N_17588,N_8204,N_8146);
nor U17589 (N_17589,N_11782,N_8704);
nand U17590 (N_17590,N_9481,N_9084);
and U17591 (N_17591,N_11236,N_6624);
xor U17592 (N_17592,N_9711,N_8143);
xor U17593 (N_17593,N_10713,N_8455);
and U17594 (N_17594,N_10809,N_6377);
and U17595 (N_17595,N_9653,N_11029);
nor U17596 (N_17596,N_10709,N_6037);
or U17597 (N_17597,N_9806,N_7769);
nand U17598 (N_17598,N_9652,N_11963);
nand U17599 (N_17599,N_6941,N_9450);
or U17600 (N_17600,N_7715,N_6023);
and U17601 (N_17601,N_7899,N_8031);
xnor U17602 (N_17602,N_7640,N_7886);
and U17603 (N_17603,N_11901,N_9106);
xor U17604 (N_17604,N_6731,N_9791);
xor U17605 (N_17605,N_10388,N_8442);
xnor U17606 (N_17606,N_7777,N_11673);
and U17607 (N_17607,N_11217,N_11902);
or U17608 (N_17608,N_9127,N_11196);
xor U17609 (N_17609,N_6555,N_10366);
nand U17610 (N_17610,N_10137,N_10643);
and U17611 (N_17611,N_7553,N_8559);
xor U17612 (N_17612,N_6633,N_8030);
and U17613 (N_17613,N_6679,N_6857);
nand U17614 (N_17614,N_6510,N_10520);
nand U17615 (N_17615,N_7320,N_8978);
nor U17616 (N_17616,N_8694,N_10165);
nand U17617 (N_17617,N_9187,N_7460);
nor U17618 (N_17618,N_10272,N_11066);
xor U17619 (N_17619,N_10530,N_10550);
nor U17620 (N_17620,N_6261,N_6899);
or U17621 (N_17621,N_11124,N_7907);
nand U17622 (N_17622,N_10835,N_8953);
xnor U17623 (N_17623,N_10413,N_6785);
nand U17624 (N_17624,N_6769,N_11759);
or U17625 (N_17625,N_8776,N_10816);
and U17626 (N_17626,N_7629,N_6392);
and U17627 (N_17627,N_9180,N_11509);
nand U17628 (N_17628,N_11193,N_8276);
nand U17629 (N_17629,N_11310,N_10590);
nor U17630 (N_17630,N_7954,N_7489);
and U17631 (N_17631,N_8208,N_6279);
or U17632 (N_17632,N_10331,N_10212);
xor U17633 (N_17633,N_9661,N_10684);
or U17634 (N_17634,N_9308,N_6467);
and U17635 (N_17635,N_8844,N_7897);
nor U17636 (N_17636,N_10337,N_10204);
nor U17637 (N_17637,N_8480,N_7562);
and U17638 (N_17638,N_8577,N_11830);
and U17639 (N_17639,N_7614,N_9136);
nand U17640 (N_17640,N_10611,N_7052);
nand U17641 (N_17641,N_9952,N_9459);
and U17642 (N_17642,N_11319,N_7757);
or U17643 (N_17643,N_6899,N_7733);
and U17644 (N_17644,N_6550,N_6146);
or U17645 (N_17645,N_9425,N_6307);
nor U17646 (N_17646,N_10628,N_7418);
xnor U17647 (N_17647,N_7966,N_9393);
nor U17648 (N_17648,N_7287,N_9849);
and U17649 (N_17649,N_9370,N_10386);
xnor U17650 (N_17650,N_9523,N_9834);
nor U17651 (N_17651,N_9025,N_6584);
or U17652 (N_17652,N_11533,N_9201);
or U17653 (N_17653,N_7730,N_9816);
xor U17654 (N_17654,N_6252,N_7086);
xnor U17655 (N_17655,N_7461,N_10778);
nand U17656 (N_17656,N_6650,N_9768);
nand U17657 (N_17657,N_8966,N_11936);
and U17658 (N_17658,N_10930,N_10727);
nor U17659 (N_17659,N_11295,N_7180);
and U17660 (N_17660,N_6896,N_11840);
nor U17661 (N_17661,N_6211,N_9425);
xnor U17662 (N_17662,N_9796,N_6272);
xor U17663 (N_17663,N_10275,N_11402);
and U17664 (N_17664,N_11814,N_10155);
and U17665 (N_17665,N_6832,N_9570);
xnor U17666 (N_17666,N_9615,N_11754);
nand U17667 (N_17667,N_7984,N_10480);
nor U17668 (N_17668,N_10999,N_10902);
nor U17669 (N_17669,N_6885,N_11777);
or U17670 (N_17670,N_8195,N_8892);
nor U17671 (N_17671,N_6970,N_8386);
and U17672 (N_17672,N_6978,N_6177);
nor U17673 (N_17673,N_7567,N_11181);
xnor U17674 (N_17674,N_7447,N_11145);
or U17675 (N_17675,N_6483,N_6886);
xor U17676 (N_17676,N_6425,N_9593);
nand U17677 (N_17677,N_10569,N_9115);
or U17678 (N_17678,N_7550,N_11331);
xnor U17679 (N_17679,N_8346,N_6891);
xor U17680 (N_17680,N_8917,N_9710);
and U17681 (N_17681,N_10620,N_11152);
or U17682 (N_17682,N_11792,N_10511);
nand U17683 (N_17683,N_11449,N_8577);
nor U17684 (N_17684,N_7176,N_7989);
and U17685 (N_17685,N_11679,N_7802);
and U17686 (N_17686,N_6225,N_6802);
or U17687 (N_17687,N_10659,N_7012);
and U17688 (N_17688,N_10923,N_9097);
or U17689 (N_17689,N_6684,N_6627);
nor U17690 (N_17690,N_8263,N_8767);
nand U17691 (N_17691,N_10571,N_10151);
and U17692 (N_17692,N_10848,N_7528);
or U17693 (N_17693,N_10408,N_8915);
and U17694 (N_17694,N_6723,N_11195);
nor U17695 (N_17695,N_8463,N_11503);
nor U17696 (N_17696,N_6621,N_7870);
nor U17697 (N_17697,N_7388,N_6754);
and U17698 (N_17698,N_8150,N_6854);
nor U17699 (N_17699,N_8395,N_10634);
and U17700 (N_17700,N_8055,N_9441);
or U17701 (N_17701,N_6077,N_6860);
and U17702 (N_17702,N_6862,N_8609);
and U17703 (N_17703,N_6283,N_8484);
nor U17704 (N_17704,N_10513,N_10501);
and U17705 (N_17705,N_7864,N_9428);
or U17706 (N_17706,N_8228,N_9540);
and U17707 (N_17707,N_8400,N_9667);
nand U17708 (N_17708,N_7346,N_7997);
nor U17709 (N_17709,N_10558,N_8950);
or U17710 (N_17710,N_9146,N_11852);
nand U17711 (N_17711,N_11977,N_11663);
and U17712 (N_17712,N_11093,N_6277);
or U17713 (N_17713,N_9376,N_10258);
nand U17714 (N_17714,N_11263,N_9258);
and U17715 (N_17715,N_10281,N_10683);
and U17716 (N_17716,N_11292,N_10261);
nor U17717 (N_17717,N_6643,N_11750);
and U17718 (N_17718,N_11390,N_9934);
or U17719 (N_17719,N_11319,N_9833);
xor U17720 (N_17720,N_9774,N_7393);
and U17721 (N_17721,N_11112,N_6468);
and U17722 (N_17722,N_10137,N_6018);
nor U17723 (N_17723,N_6648,N_9971);
or U17724 (N_17724,N_8841,N_10529);
or U17725 (N_17725,N_7554,N_11205);
and U17726 (N_17726,N_10574,N_6096);
and U17727 (N_17727,N_9754,N_7057);
nand U17728 (N_17728,N_8799,N_7002);
nand U17729 (N_17729,N_9939,N_7736);
nor U17730 (N_17730,N_11586,N_9186);
or U17731 (N_17731,N_9098,N_11987);
nor U17732 (N_17732,N_6671,N_6878);
xnor U17733 (N_17733,N_11668,N_9076);
nand U17734 (N_17734,N_11686,N_9852);
nor U17735 (N_17735,N_6046,N_9385);
or U17736 (N_17736,N_10414,N_6231);
nand U17737 (N_17737,N_11468,N_9290);
nand U17738 (N_17738,N_9167,N_11746);
or U17739 (N_17739,N_9994,N_6900);
and U17740 (N_17740,N_7330,N_8470);
xor U17741 (N_17741,N_10015,N_10989);
and U17742 (N_17742,N_11589,N_9067);
nand U17743 (N_17743,N_9946,N_7132);
nor U17744 (N_17744,N_8252,N_10062);
nor U17745 (N_17745,N_8833,N_8152);
and U17746 (N_17746,N_11895,N_10692);
or U17747 (N_17747,N_10092,N_6605);
nor U17748 (N_17748,N_10504,N_9300);
nor U17749 (N_17749,N_10896,N_10248);
or U17750 (N_17750,N_6862,N_9589);
nor U17751 (N_17751,N_8960,N_11715);
nand U17752 (N_17752,N_8694,N_10289);
or U17753 (N_17753,N_8988,N_7631);
xor U17754 (N_17754,N_10532,N_9131);
nor U17755 (N_17755,N_7120,N_8605);
xnor U17756 (N_17756,N_11253,N_8424);
or U17757 (N_17757,N_6468,N_8453);
xnor U17758 (N_17758,N_10286,N_7037);
nand U17759 (N_17759,N_9830,N_7472);
or U17760 (N_17760,N_9451,N_6474);
nor U17761 (N_17761,N_11985,N_10608);
nor U17762 (N_17762,N_6736,N_8401);
and U17763 (N_17763,N_9253,N_7015);
nand U17764 (N_17764,N_10941,N_7196);
xor U17765 (N_17765,N_6751,N_7478);
xnor U17766 (N_17766,N_11591,N_7011);
nand U17767 (N_17767,N_11194,N_8548);
or U17768 (N_17768,N_8867,N_11063);
and U17769 (N_17769,N_10197,N_7571);
xor U17770 (N_17770,N_11828,N_11647);
and U17771 (N_17771,N_7945,N_10694);
or U17772 (N_17772,N_10479,N_8501);
nand U17773 (N_17773,N_8792,N_9644);
and U17774 (N_17774,N_9910,N_9670);
and U17775 (N_17775,N_11469,N_11765);
nand U17776 (N_17776,N_10517,N_7366);
and U17777 (N_17777,N_11219,N_9499);
xor U17778 (N_17778,N_9573,N_11327);
nand U17779 (N_17779,N_8241,N_6336);
or U17780 (N_17780,N_8193,N_6522);
or U17781 (N_17781,N_6443,N_10995);
nand U17782 (N_17782,N_7814,N_9168);
or U17783 (N_17783,N_7097,N_6929);
nand U17784 (N_17784,N_9867,N_10069);
and U17785 (N_17785,N_8791,N_9816);
nor U17786 (N_17786,N_11097,N_8541);
and U17787 (N_17787,N_11614,N_10176);
and U17788 (N_17788,N_11115,N_9941);
nand U17789 (N_17789,N_9444,N_9293);
or U17790 (N_17790,N_8852,N_11922);
nor U17791 (N_17791,N_9242,N_11931);
xor U17792 (N_17792,N_7995,N_7612);
and U17793 (N_17793,N_7343,N_6796);
nand U17794 (N_17794,N_11032,N_6050);
nand U17795 (N_17795,N_8926,N_11894);
and U17796 (N_17796,N_7833,N_11328);
or U17797 (N_17797,N_9604,N_8266);
nand U17798 (N_17798,N_9887,N_9228);
and U17799 (N_17799,N_9075,N_10380);
nor U17800 (N_17800,N_7166,N_11327);
nand U17801 (N_17801,N_11714,N_9817);
xor U17802 (N_17802,N_9687,N_6526);
nor U17803 (N_17803,N_11759,N_8749);
nand U17804 (N_17804,N_9158,N_10115);
nor U17805 (N_17805,N_11727,N_10813);
nor U17806 (N_17806,N_8490,N_8570);
nand U17807 (N_17807,N_6394,N_7957);
nor U17808 (N_17808,N_10901,N_7696);
nor U17809 (N_17809,N_7984,N_8020);
nor U17810 (N_17810,N_8717,N_9419);
xor U17811 (N_17811,N_9901,N_11062);
xnor U17812 (N_17812,N_9839,N_6128);
or U17813 (N_17813,N_8640,N_9341);
or U17814 (N_17814,N_8131,N_6386);
nand U17815 (N_17815,N_9442,N_6886);
nand U17816 (N_17816,N_11864,N_11477);
xor U17817 (N_17817,N_6637,N_8653);
nand U17818 (N_17818,N_6793,N_6730);
and U17819 (N_17819,N_9934,N_6473);
nor U17820 (N_17820,N_7141,N_9139);
nand U17821 (N_17821,N_8354,N_11749);
nand U17822 (N_17822,N_10184,N_11200);
or U17823 (N_17823,N_7493,N_11452);
nor U17824 (N_17824,N_7258,N_7461);
xor U17825 (N_17825,N_7379,N_6042);
and U17826 (N_17826,N_7618,N_11167);
nor U17827 (N_17827,N_6161,N_6656);
nand U17828 (N_17828,N_9508,N_10779);
nand U17829 (N_17829,N_7862,N_7790);
or U17830 (N_17830,N_10392,N_8680);
or U17831 (N_17831,N_7542,N_7242);
nor U17832 (N_17832,N_9577,N_9206);
nor U17833 (N_17833,N_9770,N_10310);
xor U17834 (N_17834,N_10965,N_8593);
nand U17835 (N_17835,N_10179,N_9468);
nor U17836 (N_17836,N_8267,N_11333);
or U17837 (N_17837,N_10268,N_8990);
nor U17838 (N_17838,N_8350,N_7642);
nand U17839 (N_17839,N_7557,N_8951);
or U17840 (N_17840,N_8100,N_10777);
nand U17841 (N_17841,N_7898,N_11335);
xor U17842 (N_17842,N_7939,N_10997);
nand U17843 (N_17843,N_8566,N_6587);
and U17844 (N_17844,N_6141,N_10717);
xor U17845 (N_17845,N_11685,N_7103);
and U17846 (N_17846,N_11310,N_8381);
xor U17847 (N_17847,N_6609,N_8959);
or U17848 (N_17848,N_6785,N_9348);
nand U17849 (N_17849,N_6722,N_9243);
and U17850 (N_17850,N_7257,N_10317);
and U17851 (N_17851,N_6306,N_8973);
nand U17852 (N_17852,N_11018,N_9159);
and U17853 (N_17853,N_6953,N_9398);
nand U17854 (N_17854,N_10307,N_10807);
nor U17855 (N_17855,N_9726,N_6179);
and U17856 (N_17856,N_11811,N_8325);
and U17857 (N_17857,N_7581,N_11421);
or U17858 (N_17858,N_6968,N_7904);
nor U17859 (N_17859,N_10645,N_10978);
or U17860 (N_17860,N_7106,N_8462);
or U17861 (N_17861,N_10127,N_8217);
xnor U17862 (N_17862,N_10576,N_9361);
xor U17863 (N_17863,N_11927,N_11867);
and U17864 (N_17864,N_9685,N_6633);
nand U17865 (N_17865,N_11393,N_10950);
nor U17866 (N_17866,N_10026,N_7866);
or U17867 (N_17867,N_10343,N_9206);
and U17868 (N_17868,N_9583,N_8355);
and U17869 (N_17869,N_7461,N_10891);
nor U17870 (N_17870,N_11911,N_11341);
or U17871 (N_17871,N_9621,N_11626);
and U17872 (N_17872,N_7186,N_11073);
or U17873 (N_17873,N_7778,N_6941);
or U17874 (N_17874,N_11425,N_10022);
or U17875 (N_17875,N_9035,N_8179);
nor U17876 (N_17876,N_11799,N_9397);
nand U17877 (N_17877,N_9923,N_10918);
or U17878 (N_17878,N_10882,N_10074);
nand U17879 (N_17879,N_10216,N_10401);
and U17880 (N_17880,N_10532,N_8827);
xor U17881 (N_17881,N_9557,N_10553);
and U17882 (N_17882,N_8849,N_7729);
nand U17883 (N_17883,N_11766,N_10645);
nor U17884 (N_17884,N_9645,N_7687);
nor U17885 (N_17885,N_9219,N_7673);
nand U17886 (N_17886,N_11091,N_9884);
nand U17887 (N_17887,N_10691,N_11925);
or U17888 (N_17888,N_6259,N_9272);
xnor U17889 (N_17889,N_11414,N_8420);
nor U17890 (N_17890,N_9229,N_11198);
nor U17891 (N_17891,N_9282,N_10989);
nor U17892 (N_17892,N_10275,N_7832);
or U17893 (N_17893,N_9532,N_8065);
nor U17894 (N_17894,N_7427,N_7663);
or U17895 (N_17895,N_9807,N_6897);
nor U17896 (N_17896,N_11620,N_8513);
or U17897 (N_17897,N_11383,N_6043);
or U17898 (N_17898,N_6745,N_10058);
and U17899 (N_17899,N_8267,N_11109);
or U17900 (N_17900,N_6678,N_9074);
and U17901 (N_17901,N_6978,N_9411);
xnor U17902 (N_17902,N_6102,N_11473);
nor U17903 (N_17903,N_8600,N_7186);
or U17904 (N_17904,N_11165,N_7600);
and U17905 (N_17905,N_10742,N_11189);
or U17906 (N_17906,N_8022,N_9702);
and U17907 (N_17907,N_8258,N_9176);
nor U17908 (N_17908,N_8725,N_10410);
nand U17909 (N_17909,N_9250,N_6480);
nand U17910 (N_17910,N_10029,N_6674);
and U17911 (N_17911,N_8133,N_8345);
nand U17912 (N_17912,N_9321,N_7380);
or U17913 (N_17913,N_6014,N_9547);
and U17914 (N_17914,N_9038,N_6627);
xor U17915 (N_17915,N_7293,N_8401);
nand U17916 (N_17916,N_7110,N_7590);
xor U17917 (N_17917,N_10992,N_11713);
or U17918 (N_17918,N_11245,N_6496);
nor U17919 (N_17919,N_7205,N_6612);
nor U17920 (N_17920,N_6127,N_10615);
and U17921 (N_17921,N_9138,N_10277);
nand U17922 (N_17922,N_8259,N_8807);
xor U17923 (N_17923,N_10525,N_9549);
and U17924 (N_17924,N_6011,N_8898);
nor U17925 (N_17925,N_7666,N_10188);
nand U17926 (N_17926,N_10789,N_10224);
nand U17927 (N_17927,N_6076,N_10237);
xor U17928 (N_17928,N_10414,N_7612);
xor U17929 (N_17929,N_9703,N_10059);
and U17930 (N_17930,N_9815,N_11949);
nor U17931 (N_17931,N_6038,N_8821);
or U17932 (N_17932,N_6418,N_11541);
nor U17933 (N_17933,N_9650,N_6740);
xnor U17934 (N_17934,N_7856,N_6274);
nand U17935 (N_17935,N_7346,N_7171);
nand U17936 (N_17936,N_6302,N_11769);
and U17937 (N_17937,N_9950,N_11574);
nor U17938 (N_17938,N_7750,N_10725);
or U17939 (N_17939,N_11865,N_7544);
or U17940 (N_17940,N_6874,N_9826);
or U17941 (N_17941,N_7127,N_9033);
and U17942 (N_17942,N_11782,N_8449);
and U17943 (N_17943,N_6595,N_11065);
xnor U17944 (N_17944,N_8880,N_9899);
or U17945 (N_17945,N_9325,N_9431);
nand U17946 (N_17946,N_6447,N_9759);
nor U17947 (N_17947,N_6171,N_7350);
nand U17948 (N_17948,N_10849,N_6918);
nor U17949 (N_17949,N_10539,N_10905);
nor U17950 (N_17950,N_9024,N_7813);
nor U17951 (N_17951,N_8656,N_10264);
nand U17952 (N_17952,N_10935,N_11353);
xor U17953 (N_17953,N_7298,N_6461);
nand U17954 (N_17954,N_8412,N_9956);
and U17955 (N_17955,N_7054,N_11894);
or U17956 (N_17956,N_10880,N_11965);
nand U17957 (N_17957,N_7237,N_8393);
nor U17958 (N_17958,N_10479,N_8423);
nor U17959 (N_17959,N_7663,N_9727);
xnor U17960 (N_17960,N_7133,N_10712);
nand U17961 (N_17961,N_11298,N_7933);
nor U17962 (N_17962,N_8017,N_7387);
and U17963 (N_17963,N_6473,N_6393);
or U17964 (N_17964,N_11218,N_7804);
or U17965 (N_17965,N_11145,N_8052);
xnor U17966 (N_17966,N_8965,N_7107);
nor U17967 (N_17967,N_7184,N_10649);
or U17968 (N_17968,N_9704,N_8961);
nand U17969 (N_17969,N_11835,N_6489);
xor U17970 (N_17970,N_9808,N_6986);
xnor U17971 (N_17971,N_6410,N_7149);
xnor U17972 (N_17972,N_7963,N_6449);
and U17973 (N_17973,N_6812,N_9985);
nand U17974 (N_17974,N_9681,N_8530);
and U17975 (N_17975,N_9064,N_11856);
nand U17976 (N_17976,N_9287,N_6901);
or U17977 (N_17977,N_6934,N_7157);
nor U17978 (N_17978,N_8719,N_11633);
and U17979 (N_17979,N_9491,N_6168);
xor U17980 (N_17980,N_10025,N_7204);
nand U17981 (N_17981,N_8623,N_7538);
or U17982 (N_17982,N_10309,N_7659);
xnor U17983 (N_17983,N_6421,N_6844);
nand U17984 (N_17984,N_6797,N_10655);
and U17985 (N_17985,N_9517,N_11758);
or U17986 (N_17986,N_7185,N_9288);
nor U17987 (N_17987,N_9886,N_8802);
nor U17988 (N_17988,N_10424,N_10990);
nand U17989 (N_17989,N_7757,N_8744);
nand U17990 (N_17990,N_8051,N_11497);
or U17991 (N_17991,N_7950,N_11087);
nor U17992 (N_17992,N_9472,N_7357);
and U17993 (N_17993,N_8242,N_10569);
xnor U17994 (N_17994,N_7361,N_8363);
nand U17995 (N_17995,N_10198,N_6916);
nor U17996 (N_17996,N_7356,N_10452);
nand U17997 (N_17997,N_9365,N_11750);
nand U17998 (N_17998,N_8147,N_7169);
and U17999 (N_17999,N_7500,N_11834);
and U18000 (N_18000,N_13309,N_14723);
nor U18001 (N_18001,N_16753,N_13161);
nand U18002 (N_18002,N_15777,N_15813);
or U18003 (N_18003,N_13609,N_16839);
nor U18004 (N_18004,N_13325,N_13747);
and U18005 (N_18005,N_17138,N_17975);
xnor U18006 (N_18006,N_15076,N_15241);
xor U18007 (N_18007,N_12058,N_16600);
or U18008 (N_18008,N_13103,N_16379);
nand U18009 (N_18009,N_17087,N_15832);
or U18010 (N_18010,N_12112,N_15977);
and U18011 (N_18011,N_17384,N_13199);
or U18012 (N_18012,N_17373,N_13176);
and U18013 (N_18013,N_13565,N_16250);
xor U18014 (N_18014,N_16328,N_15688);
nor U18015 (N_18015,N_16408,N_15510);
and U18016 (N_18016,N_15147,N_14730);
nand U18017 (N_18017,N_12697,N_13310);
nand U18018 (N_18018,N_17772,N_17552);
or U18019 (N_18019,N_16259,N_17357);
nand U18020 (N_18020,N_15600,N_17162);
or U18021 (N_18021,N_13919,N_12127);
xnor U18022 (N_18022,N_16254,N_12710);
and U18023 (N_18023,N_16874,N_15134);
nand U18024 (N_18024,N_16786,N_12348);
xnor U18025 (N_18025,N_13964,N_15718);
or U18026 (N_18026,N_13872,N_12769);
nor U18027 (N_18027,N_17962,N_12427);
nor U18028 (N_18028,N_13195,N_17313);
xor U18029 (N_18029,N_14878,N_14257);
nor U18030 (N_18030,N_14280,N_15377);
and U18031 (N_18031,N_17199,N_14591);
nand U18032 (N_18032,N_14958,N_13519);
nor U18033 (N_18033,N_17548,N_17059);
or U18034 (N_18034,N_15712,N_14446);
xnor U18035 (N_18035,N_14367,N_12502);
or U18036 (N_18036,N_16823,N_13480);
nand U18037 (N_18037,N_13462,N_12435);
nand U18038 (N_18038,N_12480,N_15272);
xor U18039 (N_18039,N_16351,N_12102);
nand U18040 (N_18040,N_17562,N_14140);
xor U18041 (N_18041,N_13220,N_16972);
nor U18042 (N_18042,N_15169,N_15914);
and U18043 (N_18043,N_12837,N_12218);
and U18044 (N_18044,N_15238,N_14255);
nor U18045 (N_18045,N_15925,N_15677);
nor U18046 (N_18046,N_16237,N_12096);
nor U18047 (N_18047,N_16426,N_13746);
or U18048 (N_18048,N_13253,N_16130);
nand U18049 (N_18049,N_14356,N_12984);
nor U18050 (N_18050,N_12315,N_16005);
or U18051 (N_18051,N_14177,N_15244);
xnor U18052 (N_18052,N_13643,N_13223);
nand U18053 (N_18053,N_13332,N_16196);
or U18054 (N_18054,N_14141,N_15975);
or U18055 (N_18055,N_12347,N_13236);
and U18056 (N_18056,N_17394,N_13046);
or U18057 (N_18057,N_17558,N_17420);
nand U18058 (N_18058,N_13007,N_17148);
and U18059 (N_18059,N_13151,N_14099);
xnor U18060 (N_18060,N_14284,N_15230);
nor U18061 (N_18061,N_14150,N_12303);
nand U18062 (N_18062,N_12660,N_14914);
nor U18063 (N_18063,N_12320,N_14756);
nor U18064 (N_18064,N_15397,N_16820);
or U18065 (N_18065,N_17710,N_16164);
and U18066 (N_18066,N_17591,N_16424);
nand U18067 (N_18067,N_15261,N_17079);
nand U18068 (N_18068,N_13686,N_16766);
nand U18069 (N_18069,N_13128,N_14176);
or U18070 (N_18070,N_13698,N_14139);
nor U18071 (N_18071,N_13755,N_17919);
and U18072 (N_18072,N_12706,N_17714);
and U18073 (N_18073,N_13976,N_16582);
and U18074 (N_18074,N_14473,N_15470);
xor U18075 (N_18075,N_16664,N_15066);
and U18076 (N_18076,N_14910,N_14221);
or U18077 (N_18077,N_17312,N_13264);
nand U18078 (N_18078,N_15254,N_16593);
nand U18079 (N_18079,N_15376,N_14035);
and U18080 (N_18080,N_12164,N_17198);
nor U18081 (N_18081,N_14364,N_14429);
nor U18082 (N_18082,N_12300,N_14934);
and U18083 (N_18083,N_15372,N_16634);
nor U18084 (N_18084,N_12605,N_16461);
nand U18085 (N_18085,N_17887,N_14037);
xor U18086 (N_18086,N_12270,N_17554);
and U18087 (N_18087,N_17435,N_17091);
or U18088 (N_18088,N_14091,N_16743);
nor U18089 (N_18089,N_15497,N_16904);
nand U18090 (N_18090,N_16622,N_15528);
nand U18091 (N_18091,N_15083,N_16098);
xnor U18092 (N_18092,N_16526,N_12634);
nand U18093 (N_18093,N_16176,N_16769);
or U18094 (N_18094,N_12225,N_13774);
and U18095 (N_18095,N_14541,N_15594);
xor U18096 (N_18096,N_14464,N_14128);
or U18097 (N_18097,N_17186,N_14351);
nor U18098 (N_18098,N_13918,N_17106);
and U18099 (N_18099,N_17544,N_15828);
xnor U18100 (N_18100,N_14931,N_13801);
nor U18101 (N_18101,N_15296,N_16261);
xor U18102 (N_18102,N_16594,N_12911);
and U18103 (N_18103,N_14537,N_14892);
or U18104 (N_18104,N_13868,N_16206);
nand U18105 (N_18105,N_16893,N_14854);
or U18106 (N_18106,N_13384,N_14437);
xnor U18107 (N_18107,N_17927,N_14234);
nand U18108 (N_18108,N_13299,N_15219);
nand U18109 (N_18109,N_15086,N_16875);
xnor U18110 (N_18110,N_16301,N_14462);
xnor U18111 (N_18111,N_16434,N_13379);
nor U18112 (N_18112,N_12784,N_14058);
nor U18113 (N_18113,N_12556,N_16761);
and U18114 (N_18114,N_13559,N_12592);
xor U18115 (N_18115,N_15571,N_15611);
or U18116 (N_18116,N_17187,N_16486);
or U18117 (N_18117,N_13394,N_12254);
nor U18118 (N_18118,N_12169,N_13461);
nand U18119 (N_18119,N_16018,N_16213);
or U18120 (N_18120,N_12123,N_14387);
and U18121 (N_18121,N_13181,N_12441);
xor U18122 (N_18122,N_12179,N_14592);
nand U18123 (N_18123,N_14186,N_13425);
or U18124 (N_18124,N_15865,N_14406);
nor U18125 (N_18125,N_17523,N_12230);
or U18126 (N_18126,N_13884,N_13557);
nand U18127 (N_18127,N_17350,N_14774);
and U18128 (N_18128,N_15052,N_17581);
nor U18129 (N_18129,N_13693,N_13427);
nor U18130 (N_18130,N_12758,N_15746);
nor U18131 (N_18131,N_17053,N_13039);
nand U18132 (N_18132,N_15609,N_12700);
or U18133 (N_18133,N_17702,N_12770);
nor U18134 (N_18134,N_12419,N_13776);
xnor U18135 (N_18135,N_17925,N_17612);
or U18136 (N_18136,N_15585,N_16479);
nor U18137 (N_18137,N_16722,N_17078);
or U18138 (N_18138,N_13120,N_14414);
or U18139 (N_18139,N_12155,N_15429);
xnor U18140 (N_18140,N_14922,N_13691);
nor U18141 (N_18141,N_15093,N_15969);
nor U18142 (N_18142,N_17092,N_15324);
and U18143 (N_18143,N_15620,N_15684);
xor U18144 (N_18144,N_14156,N_15519);
and U18145 (N_18145,N_14070,N_12606);
nand U18146 (N_18146,N_16077,N_12167);
xor U18147 (N_18147,N_15907,N_15649);
or U18148 (N_18148,N_14815,N_13994);
nand U18149 (N_18149,N_13647,N_15651);
nor U18150 (N_18150,N_14779,N_17922);
or U18151 (N_18151,N_14641,N_15686);
nor U18152 (N_18152,N_13378,N_12460);
nor U18153 (N_18153,N_17484,N_17587);
nand U18154 (N_18154,N_17039,N_13386);
xor U18155 (N_18155,N_13540,N_17153);
xor U18156 (N_18156,N_12530,N_13237);
nor U18157 (N_18157,N_17691,N_14456);
and U18158 (N_18158,N_13912,N_14836);
and U18159 (N_18159,N_16111,N_12628);
xor U18160 (N_18160,N_13988,N_15165);
nor U18161 (N_18161,N_12065,N_15517);
and U18162 (N_18162,N_14278,N_14082);
xor U18163 (N_18163,N_15741,N_15447);
xnor U18164 (N_18164,N_16986,N_12656);
and U18165 (N_18165,N_17391,N_16534);
xnor U18166 (N_18166,N_17040,N_15088);
or U18167 (N_18167,N_16861,N_13187);
nand U18168 (N_18168,N_12060,N_15970);
xnor U18169 (N_18169,N_14864,N_14845);
or U18170 (N_18170,N_13337,N_16046);
xnor U18171 (N_18171,N_15524,N_15862);
and U18172 (N_18172,N_12172,N_14321);
xor U18173 (N_18173,N_16420,N_16982);
xnor U18174 (N_18174,N_12386,N_12082);
nor U18175 (N_18175,N_12509,N_15009);
and U18176 (N_18176,N_12566,N_13257);
and U18177 (N_18177,N_17054,N_14108);
or U18178 (N_18178,N_17147,N_15680);
nor U18179 (N_18179,N_14515,N_13485);
nand U18180 (N_18180,N_12339,N_15547);
nand U18181 (N_18181,N_16455,N_17487);
nand U18182 (N_18182,N_17288,N_13247);
nor U18183 (N_18183,N_17004,N_17972);
and U18184 (N_18184,N_17959,N_16059);
or U18185 (N_18185,N_13629,N_16521);
or U18186 (N_18186,N_12901,N_17692);
xor U18187 (N_18187,N_15409,N_14149);
and U18188 (N_18188,N_12773,N_17620);
nor U18189 (N_18189,N_14699,N_16210);
or U18190 (N_18190,N_15352,N_17640);
nand U18191 (N_18191,N_14528,N_13662);
nand U18192 (N_18192,N_17322,N_16025);
or U18193 (N_18193,N_14790,N_13071);
nand U18194 (N_18194,N_14759,N_12174);
nand U18195 (N_18195,N_15877,N_16106);
and U18196 (N_18196,N_16207,N_17607);
nor U18197 (N_18197,N_12716,N_16884);
nand U18198 (N_18198,N_12830,N_15802);
nor U18199 (N_18199,N_16507,N_17434);
xor U18200 (N_18200,N_13501,N_15366);
and U18201 (N_18201,N_15455,N_12594);
nand U18202 (N_18202,N_15826,N_14214);
and U18203 (N_18203,N_15054,N_16191);
or U18204 (N_18204,N_14605,N_16710);
or U18205 (N_18205,N_14427,N_12229);
nand U18206 (N_18206,N_12908,N_14154);
and U18207 (N_18207,N_13751,N_12704);
and U18208 (N_18208,N_15252,N_16709);
and U18209 (N_18209,N_15889,N_14238);
xor U18210 (N_18210,N_14978,N_14152);
and U18211 (N_18211,N_12863,N_16173);
xor U18212 (N_18212,N_13213,N_15941);
and U18213 (N_18213,N_15520,N_14308);
nand U18214 (N_18214,N_15477,N_15583);
or U18215 (N_18215,N_12917,N_14867);
and U18216 (N_18216,N_17014,N_12681);
nor U18217 (N_18217,N_13465,N_12399);
xor U18218 (N_18218,N_12925,N_14106);
or U18219 (N_18219,N_14757,N_13757);
nor U18220 (N_18220,N_16219,N_16590);
nor U18221 (N_18221,N_16027,N_17169);
or U18222 (N_18222,N_17097,N_17404);
or U18223 (N_18223,N_12068,N_15807);
and U18224 (N_18224,N_14946,N_17285);
and U18225 (N_18225,N_15617,N_17117);
and U18226 (N_18226,N_12162,N_13363);
nor U18227 (N_18227,N_16319,N_17726);
and U18228 (N_18228,N_17760,N_17996);
xor U18229 (N_18229,N_13721,N_17084);
nor U18230 (N_18230,N_13252,N_17409);
and U18231 (N_18231,N_13082,N_14219);
xnor U18232 (N_18232,N_17622,N_14969);
nor U18233 (N_18233,N_15428,N_13466);
and U18234 (N_18234,N_17593,N_13273);
or U18235 (N_18235,N_14500,N_13162);
or U18236 (N_18236,N_12195,N_13869);
nor U18237 (N_18237,N_13612,N_17597);
and U18238 (N_18238,N_14374,N_13148);
or U18239 (N_18239,N_15494,N_15613);
xor U18240 (N_18240,N_17197,N_13726);
or U18241 (N_18241,N_14337,N_17496);
xnor U18242 (N_18242,N_14244,N_16711);
xnor U18243 (N_18243,N_12902,N_14434);
nand U18244 (N_18244,N_12540,N_14416);
nor U18245 (N_18245,N_16389,N_17795);
nor U18246 (N_18246,N_12821,N_12376);
xor U18247 (N_18247,N_16816,N_17706);
or U18248 (N_18248,N_14345,N_16555);
nor U18249 (N_18249,N_12274,N_16443);
xnor U18250 (N_18250,N_15345,N_17130);
nor U18251 (N_18251,N_15131,N_16810);
xnor U18252 (N_18252,N_14598,N_13914);
nor U18253 (N_18253,N_12576,N_17690);
or U18254 (N_18254,N_17570,N_14382);
xor U18255 (N_18255,N_16517,N_13944);
and U18256 (N_18256,N_17881,N_14460);
and U18257 (N_18257,N_14706,N_14372);
xnor U18258 (N_18258,N_12554,N_15559);
xnor U18259 (N_18259,N_16230,N_12783);
or U18260 (N_18260,N_14388,N_17224);
nor U18261 (N_18261,N_16955,N_17563);
nand U18262 (N_18262,N_14819,N_17712);
xor U18263 (N_18263,N_16684,N_15880);
nand U18264 (N_18264,N_17316,N_15876);
and U18265 (N_18265,N_16400,N_16264);
or U18266 (N_18266,N_16220,N_14005);
and U18267 (N_18267,N_14916,N_16843);
and U18268 (N_18268,N_17245,N_12688);
or U18269 (N_18269,N_15210,N_16050);
xnor U18270 (N_18270,N_16125,N_16960);
xor U18271 (N_18271,N_13591,N_13270);
xnor U18272 (N_18272,N_13929,N_14474);
nor U18273 (N_18273,N_15640,N_14135);
and U18274 (N_18274,N_12956,N_15312);
nand U18275 (N_18275,N_16421,N_14032);
xor U18276 (N_18276,N_17157,N_14334);
and U18277 (N_18277,N_15691,N_13837);
and U18278 (N_18278,N_17907,N_14668);
nand U18279 (N_18279,N_13268,N_15365);
nor U18280 (N_18280,N_13585,N_14237);
or U18281 (N_18281,N_17821,N_17880);
xor U18282 (N_18282,N_16951,N_17883);
nor U18283 (N_18283,N_15216,N_17750);
or U18284 (N_18284,N_15485,N_16789);
or U18285 (N_18285,N_13095,N_17836);
xor U18286 (N_18286,N_15708,N_17542);
nor U18287 (N_18287,N_17817,N_15607);
nand U18288 (N_18288,N_15417,N_13784);
or U18289 (N_18289,N_14253,N_12816);
xnor U18290 (N_18290,N_15323,N_16900);
nor U18291 (N_18291,N_14890,N_13375);
nand U18292 (N_18292,N_14943,N_16778);
xnor U18293 (N_18293,N_12786,N_15055);
xor U18294 (N_18294,N_16509,N_13149);
and U18295 (N_18295,N_17291,N_12792);
or U18296 (N_18296,N_13677,N_14875);
or U18297 (N_18297,N_13496,N_12472);
nor U18298 (N_18298,N_17095,N_15687);
and U18299 (N_18299,N_15157,N_13642);
and U18300 (N_18300,N_13418,N_16211);
xnor U18301 (N_18301,N_15382,N_13548);
xor U18302 (N_18302,N_12817,N_13844);
and U18303 (N_18303,N_17891,N_14195);
nor U18304 (N_18304,N_12527,N_16163);
nand U18305 (N_18305,N_15259,N_13750);
nand U18306 (N_18306,N_17223,N_17843);
or U18307 (N_18307,N_15139,N_16638);
or U18308 (N_18308,N_15848,N_12845);
or U18309 (N_18309,N_17276,N_15505);
nand U18310 (N_18310,N_12044,N_13981);
xnor U18311 (N_18311,N_16263,N_14459);
xnor U18312 (N_18312,N_16290,N_14550);
xnor U18313 (N_18313,N_12775,N_17976);
nor U18314 (N_18314,N_12856,N_17734);
nand U18315 (N_18315,N_16796,N_15019);
and U18316 (N_18316,N_12782,N_14069);
xnor U18317 (N_18317,N_17512,N_15732);
xor U18318 (N_18318,N_17708,N_13835);
nand U18319 (N_18319,N_17851,N_15881);
and U18320 (N_18320,N_14590,N_16599);
nand U18321 (N_18321,N_13690,N_17740);
nor U18322 (N_18322,N_17306,N_14493);
and U18323 (N_18323,N_17897,N_12820);
and U18324 (N_18324,N_17433,N_14595);
or U18325 (N_18325,N_12090,N_13954);
or U18326 (N_18326,N_17145,N_16682);
or U18327 (N_18327,N_17266,N_12354);
nand U18328 (N_18328,N_14695,N_13739);
nor U18329 (N_18329,N_13152,N_12343);
and U18330 (N_18330,N_12426,N_14711);
xnor U18331 (N_18331,N_17093,N_14942);
and U18332 (N_18332,N_12057,N_16536);
and U18333 (N_18333,N_13536,N_17535);
nor U18334 (N_18334,N_13985,N_16656);
nor U18335 (N_18335,N_16569,N_16645);
nand U18336 (N_18336,N_12880,N_17564);
nand U18337 (N_18337,N_17522,N_13001);
nor U18338 (N_18338,N_15422,N_17924);
nand U18339 (N_18339,N_13772,N_13968);
xnor U18340 (N_18340,N_12698,N_13804);
or U18341 (N_18341,N_16744,N_12212);
nand U18342 (N_18342,N_16723,N_15383);
or U18343 (N_18343,N_16775,N_17906);
nor U18344 (N_18344,N_16431,N_13081);
or U18345 (N_18345,N_15328,N_15648);
or U18346 (N_18346,N_15722,N_13275);
and U18347 (N_18347,N_13850,N_12895);
and U18348 (N_18348,N_17381,N_15435);
nand U18349 (N_18349,N_16931,N_15836);
nor U18350 (N_18350,N_15883,N_14556);
or U18351 (N_18351,N_13493,N_12744);
or U18352 (N_18352,N_12754,N_12317);
nand U18353 (N_18353,N_16105,N_13699);
or U18354 (N_18354,N_15187,N_13949);
nand U18355 (N_18355,N_14750,N_12785);
and U18356 (N_18356,N_12379,N_16733);
and U18357 (N_18357,N_17617,N_17214);
nand U18358 (N_18358,N_17978,N_14807);
and U18359 (N_18359,N_17069,N_12368);
nor U18360 (N_18360,N_14470,N_15325);
and U18361 (N_18361,N_13627,N_17813);
nor U18362 (N_18362,N_14410,N_17586);
and U18363 (N_18363,N_14496,N_17049);
nand U18364 (N_18364,N_16988,N_16463);
nor U18365 (N_18365,N_17218,N_13203);
xnor U18366 (N_18366,N_15016,N_17653);
nor U18367 (N_18367,N_16804,N_17272);
and U18368 (N_18368,N_13224,N_16510);
or U18369 (N_18369,N_15757,N_14430);
nand U18370 (N_18370,N_17904,N_15981);
and U18371 (N_18371,N_16574,N_17565);
xor U18372 (N_18372,N_16993,N_14924);
xnor U18373 (N_18373,N_15132,N_14273);
and U18374 (N_18374,N_17573,N_14520);
and U18375 (N_18375,N_17012,N_15924);
nor U18376 (N_18376,N_12414,N_17616);
or U18377 (N_18377,N_16053,N_12647);
nand U18378 (N_18378,N_15014,N_12484);
or U18379 (N_18379,N_12528,N_13993);
and U18380 (N_18380,N_12298,N_17718);
xor U18381 (N_18381,N_13723,N_14100);
xor U18382 (N_18382,N_12945,N_13373);
nor U18383 (N_18383,N_17329,N_15322);
nor U18384 (N_18384,N_17580,N_15068);
nand U18385 (N_18385,N_15044,N_17890);
xnor U18386 (N_18386,N_16038,N_13509);
xnor U18387 (N_18387,N_15752,N_12100);
and U18388 (N_18388,N_13170,N_14773);
and U18389 (N_18389,N_13645,N_12013);
xnor U18390 (N_18390,N_12496,N_14963);
xnor U18391 (N_18391,N_12295,N_14633);
and U18392 (N_18392,N_13896,N_15247);
nor U18393 (N_18393,N_12071,N_17982);
or U18394 (N_18394,N_15224,N_13345);
and U18395 (N_18395,N_13813,N_12147);
nor U18396 (N_18396,N_17614,N_16352);
xor U18397 (N_18397,N_16734,N_17368);
or U18398 (N_18398,N_12963,N_13889);
xor U18399 (N_18399,N_17983,N_16369);
nand U18400 (N_18400,N_17832,N_16996);
nand U18401 (N_18401,N_12964,N_14805);
and U18402 (N_18402,N_12695,N_14461);
nand U18403 (N_18403,N_16497,N_16496);
nand U18404 (N_18404,N_17732,N_16356);
or U18405 (N_18405,N_16311,N_17765);
or U18406 (N_18406,N_15701,N_12569);
nand U18407 (N_18407,N_12284,N_16054);
and U18408 (N_18408,N_12476,N_13607);
nand U18409 (N_18409,N_16348,N_15805);
nor U18410 (N_18410,N_15253,N_13841);
and U18411 (N_18411,N_16620,N_15465);
or U18412 (N_18412,N_12248,N_12599);
nor U18413 (N_18413,N_16109,N_14223);
and U18414 (N_18414,N_12999,N_17140);
or U18415 (N_18415,N_14698,N_15369);
nor U18416 (N_18416,N_14179,N_15597);
and U18417 (N_18417,N_16770,N_15133);
nand U18418 (N_18418,N_14625,N_12207);
xor U18419 (N_18419,N_16404,N_14049);
and U18420 (N_18420,N_16614,N_13488);
nor U18421 (N_18421,N_13951,N_16378);
nor U18422 (N_18422,N_16316,N_17763);
or U18423 (N_18423,N_13704,N_17397);
nand U18424 (N_18424,N_15723,N_17981);
or U18425 (N_18425,N_13055,N_16631);
nand U18426 (N_18426,N_12680,N_12542);
nor U18427 (N_18427,N_15650,N_14488);
and U18428 (N_18428,N_15662,N_13568);
and U18429 (N_18429,N_14072,N_16270);
or U18430 (N_18430,N_14904,N_15908);
nor U18431 (N_18431,N_16658,N_17652);
nor U18432 (N_18432,N_16592,N_12213);
nand U18433 (N_18433,N_13486,N_16650);
and U18434 (N_18434,N_13554,N_15892);
nor U18435 (N_18435,N_15341,N_12835);
or U18436 (N_18436,N_15338,N_12707);
xnor U18437 (N_18437,N_12967,N_16513);
and U18438 (N_18438,N_17468,N_17343);
or U18439 (N_18439,N_13374,N_16465);
and U18440 (N_18440,N_16903,N_15847);
or U18441 (N_18441,N_14405,N_14936);
or U18442 (N_18442,N_12067,N_15603);
nor U18443 (N_18443,N_17255,N_16326);
nand U18444 (N_18444,N_12352,N_16632);
or U18445 (N_18445,N_13317,N_13732);
nor U18446 (N_18446,N_17903,N_14885);
xor U18447 (N_18447,N_14409,N_15314);
or U18448 (N_18448,N_16677,N_17437);
nor U18449 (N_18449,N_13228,N_15390);
nor U18450 (N_18450,N_17380,N_16231);
or U18451 (N_18451,N_13521,N_17773);
nor U18452 (N_18452,N_16966,N_15751);
nand U18453 (N_18453,N_12390,N_14703);
xnor U18454 (N_18454,N_13763,N_12296);
nor U18455 (N_18455,N_16363,N_14563);
nand U18456 (N_18456,N_13406,N_16980);
xnor U18457 (N_18457,N_16000,N_16933);
nor U18458 (N_18458,N_15273,N_15122);
and U18459 (N_18459,N_17143,N_16030);
and U18460 (N_18460,N_15295,N_13840);
nor U18461 (N_18461,N_17671,N_14415);
and U18462 (N_18462,N_15775,N_16782);
xor U18463 (N_18463,N_12458,N_12921);
and U18464 (N_18464,N_13761,N_13953);
nor U18465 (N_18465,N_13153,N_17407);
or U18466 (N_18466,N_16994,N_17146);
nor U18467 (N_18467,N_16078,N_17791);
nand U18468 (N_18468,N_12064,N_17584);
and U18469 (N_18469,N_15697,N_15164);
nand U18470 (N_18470,N_13937,N_15459);
nand U18471 (N_18471,N_15779,N_14829);
and U18472 (N_18472,N_13091,N_12021);
or U18473 (N_18473,N_15451,N_12822);
nand U18474 (N_18474,N_14471,N_14190);
nand U18475 (N_18475,N_15543,N_14513);
and U18476 (N_18476,N_16087,N_16283);
nand U18477 (N_18477,N_17830,N_14438);
or U18478 (N_18478,N_13728,N_12571);
or U18479 (N_18479,N_12417,N_17067);
nor U18480 (N_18480,N_12525,N_14097);
nand U18481 (N_18481,N_16692,N_17733);
nand U18482 (N_18482,N_12852,N_15142);
or U18483 (N_18483,N_14159,N_17454);
or U18484 (N_18484,N_17648,N_17638);
and U18485 (N_18485,N_16449,N_16433);
xor U18486 (N_18486,N_15942,N_15286);
nand U18487 (N_18487,N_14047,N_16144);
xor U18488 (N_18488,N_17589,N_17099);
and U18489 (N_18489,N_12395,N_16837);
nor U18490 (N_18490,N_15637,N_14998);
nor U18491 (N_18491,N_12703,N_12448);
xnor U18492 (N_18492,N_14884,N_12608);
nand U18493 (N_18493,N_16653,N_14794);
xnor U18494 (N_18494,N_14354,N_16550);
nor U18495 (N_18495,N_15726,N_12046);
nor U18496 (N_18496,N_15332,N_16253);
nand U18497 (N_18497,N_13018,N_13033);
xor U18498 (N_18498,N_12012,N_17123);
or U18499 (N_18499,N_15159,N_14719);
nor U18500 (N_18500,N_13267,N_12800);
xor U18501 (N_18501,N_17196,N_13535);
or U18502 (N_18502,N_15537,N_17942);
or U18503 (N_18503,N_12673,N_16705);
nand U18504 (N_18504,N_13340,N_17260);
nand U18505 (N_18505,N_12454,N_15143);
or U18506 (N_18506,N_13833,N_14342);
xor U18507 (N_18507,N_13327,N_14555);
or U18508 (N_18508,N_15781,N_12378);
and U18509 (N_18509,N_13026,N_16693);
xor U18510 (N_18510,N_14614,N_13092);
xnor U18511 (N_18511,N_13226,N_14081);
nand U18512 (N_18512,N_16153,N_17365);
nor U18513 (N_18513,N_17815,N_13351);
nand U18514 (N_18514,N_15079,N_17406);
nor U18515 (N_18515,N_16294,N_14307);
xor U18516 (N_18516,N_17333,N_17181);
xnor U18517 (N_18517,N_12211,N_16318);
nor U18518 (N_18518,N_12299,N_15255);
nor U18519 (N_18519,N_14138,N_15971);
nand U18520 (N_18520,N_14571,N_17185);
nor U18521 (N_18521,N_12910,N_13238);
and U18522 (N_18522,N_13490,N_12795);
nor U18523 (N_18523,N_12373,N_12239);
nor U18524 (N_18524,N_17361,N_17208);
xor U18525 (N_18525,N_17411,N_17840);
or U18526 (N_18526,N_17889,N_14859);
and U18527 (N_18527,N_17678,N_16654);
and U18528 (N_18528,N_15759,N_15423);
and U18529 (N_18529,N_17759,N_15048);
and U18530 (N_18530,N_12893,N_16493);
and U18531 (N_18531,N_17395,N_13615);
nand U18532 (N_18532,N_14212,N_13423);
nor U18533 (N_18533,N_16602,N_15954);
nand U18534 (N_18534,N_17604,N_17575);
nand U18535 (N_18535,N_16150,N_17785);
xnor U18536 (N_18536,N_14930,N_15549);
nand U18537 (N_18537,N_12166,N_13923);
nand U18538 (N_18538,N_15946,N_12238);
or U18539 (N_18539,N_17464,N_17318);
nor U18540 (N_18540,N_16851,N_13050);
or U18541 (N_18541,N_15739,N_12650);
xnor U18542 (N_18542,N_15047,N_15279);
xor U18543 (N_18543,N_15317,N_16520);
xor U18544 (N_18544,N_17920,N_15867);
or U18545 (N_18545,N_14407,N_13412);
or U18546 (N_18546,N_15740,N_15576);
nor U18547 (N_18547,N_17537,N_12049);
and U18548 (N_18548,N_12888,N_13987);
and U18549 (N_18549,N_15906,N_12324);
nand U18550 (N_18550,N_14497,N_14475);
or U18551 (N_18551,N_12728,N_12613);
and U18552 (N_18552,N_16134,N_15062);
nor U18553 (N_18553,N_16713,N_14926);
xnor U18554 (N_18554,N_16359,N_14600);
or U18555 (N_18555,N_13206,N_17430);
and U18556 (N_18556,N_13049,N_14076);
xor U18557 (N_18557,N_14736,N_17119);
and U18558 (N_18558,N_12977,N_15311);
and U18559 (N_18559,N_12360,N_12975);
or U18560 (N_18560,N_16887,N_17305);
and U18561 (N_18561,N_12620,N_13105);
nor U18562 (N_18562,N_13214,N_17923);
nor U18563 (N_18563,N_15380,N_17251);
and U18564 (N_18564,N_17121,N_14379);
or U18565 (N_18565,N_14780,N_17239);
nor U18566 (N_18566,N_14296,N_17378);
and U18567 (N_18567,N_14399,N_16357);
nor U18568 (N_18568,N_17866,N_16012);
or U18569 (N_18569,N_17173,N_17860);
or U18570 (N_18570,N_15764,N_13517);
nand U18571 (N_18571,N_16475,N_13027);
nor U18572 (N_18572,N_17076,N_12720);
xnor U18573 (N_18573,N_16504,N_13468);
or U18574 (N_18574,N_13957,N_14144);
xnor U18575 (N_18575,N_17080,N_13244);
and U18576 (N_18576,N_13711,N_14557);
or U18577 (N_18577,N_16936,N_13045);
and U18578 (N_18578,N_13137,N_17594);
nand U18579 (N_18579,N_16396,N_12078);
nor U18580 (N_18580,N_12831,N_14648);
nor U18581 (N_18581,N_13925,N_15282);
or U18582 (N_18582,N_16482,N_15026);
or U18583 (N_18583,N_15367,N_13817);
nor U18584 (N_18584,N_14498,N_15915);
nor U18585 (N_18585,N_17110,N_16551);
and U18586 (N_18586,N_13792,N_12223);
xor U18587 (N_18587,N_12494,N_15031);
nor U18588 (N_18588,N_16086,N_13725);
nor U18589 (N_18589,N_15432,N_16344);
nand U18590 (N_18590,N_14205,N_17472);
nand U18591 (N_18591,N_15793,N_13580);
xnor U18592 (N_18592,N_16004,N_16801);
xnor U18593 (N_18593,N_16061,N_15833);
and U18594 (N_18594,N_17392,N_13382);
nor U18595 (N_18595,N_14769,N_14566);
and U18596 (N_18596,N_14441,N_17267);
nand U18597 (N_18597,N_12915,N_17427);
or U18598 (N_18598,N_12381,N_17238);
xor U18599 (N_18599,N_16342,N_15574);
and U18600 (N_18600,N_15953,N_12407);
nor U18601 (N_18601,N_17058,N_16827);
xor U18602 (N_18602,N_15391,N_13463);
nand U18603 (N_18603,N_12559,N_15955);
nor U18604 (N_18604,N_13142,N_14745);
and U18605 (N_18605,N_16117,N_14502);
or U18606 (N_18606,N_15661,N_12596);
and U18607 (N_18607,N_13146,N_13000);
nor U18608 (N_18608,N_13269,N_12278);
nor U18609 (N_18609,N_15769,N_12828);
nor U18610 (N_18610,N_17888,N_15340);
xnor U18611 (N_18611,N_16293,N_14631);
or U18612 (N_18612,N_13865,N_16146);
and U18613 (N_18613,N_14982,N_16737);
xnor U18614 (N_18614,N_16274,N_16052);
and U18615 (N_18615,N_15951,N_17707);
or U18616 (N_18616,N_16891,N_16407);
and U18617 (N_18617,N_12734,N_14622);
and U18618 (N_18618,N_17317,N_14311);
nand U18619 (N_18619,N_13640,N_12083);
and U18620 (N_18620,N_13458,N_15534);
nor U18621 (N_18621,N_14185,N_16472);
or U18622 (N_18622,N_13592,N_15173);
nand U18623 (N_18623,N_12671,N_15123);
nor U18624 (N_18624,N_15658,N_15669);
xnor U18625 (N_18625,N_13846,N_17028);
and U18626 (N_18626,N_12136,N_16546);
and U18627 (N_18627,N_17848,N_15467);
nor U18628 (N_18628,N_15952,N_14634);
xor U18629 (N_18629,N_15824,N_16447);
nand U18630 (N_18630,N_12165,N_17516);
and U18631 (N_18631,N_12242,N_14725);
or U18632 (N_18632,N_17926,N_13671);
xor U18633 (N_18633,N_14526,N_13354);
xor U18634 (N_18634,N_13664,N_15555);
nor U18635 (N_18635,N_14588,N_13093);
and U18636 (N_18636,N_17935,N_17385);
nand U18637 (N_18637,N_15200,N_16228);
nand U18638 (N_18638,N_14721,N_16981);
nor U18639 (N_18639,N_14549,N_17354);
nor U18640 (N_18640,N_17592,N_12003);
xnor U18641 (N_18641,N_15036,N_15846);
or U18642 (N_18642,N_13736,N_14468);
or U18643 (N_18643,N_16266,N_13256);
or U18644 (N_18644,N_12402,N_13047);
nand U18645 (N_18645,N_17226,N_16216);
or U18646 (N_18646,N_13186,N_12833);
nand U18647 (N_18647,N_13898,N_17728);
or U18648 (N_18648,N_14678,N_14991);
or U18649 (N_18649,N_12654,N_13560);
xnor U18650 (N_18650,N_15709,N_14458);
nand U18651 (N_18651,N_14783,N_17896);
xnor U18652 (N_18652,N_14596,N_16760);
or U18653 (N_18653,N_15202,N_16978);
xnor U18654 (N_18654,N_15141,N_17842);
nor U18655 (N_18655,N_16554,N_16812);
xnor U18656 (N_18656,N_14320,N_15483);
nor U18657 (N_18657,N_17977,N_14877);
xnor U18658 (N_18658,N_15707,N_13920);
or U18659 (N_18659,N_17165,N_15645);
nor U18660 (N_18660,N_17349,N_15866);
or U18661 (N_18661,N_17770,N_16033);
nor U18662 (N_18662,N_13621,N_13122);
nand U18663 (N_18663,N_14084,N_14312);
nor U18664 (N_18664,N_14053,N_16880);
or U18665 (N_18665,N_12764,N_14760);
or U18666 (N_18666,N_13979,N_17327);
nand U18667 (N_18667,N_13318,N_13111);
nand U18668 (N_18668,N_15006,N_13653);
nand U18669 (N_18669,N_17127,N_12098);
and U18670 (N_18670,N_15001,N_12772);
xor U18671 (N_18671,N_16322,N_17649);
and U18672 (N_18672,N_14249,N_16791);
xnor U18673 (N_18673,N_14180,N_12081);
nor U18674 (N_18674,N_13429,N_15321);
nor U18675 (N_18675,N_15407,N_15765);
nand U18676 (N_18676,N_15109,N_16126);
or U18677 (N_18677,N_17937,N_15023);
nand U18678 (N_18678,N_16665,N_12919);
nor U18679 (N_18679,N_12188,N_15269);
and U18680 (N_18680,N_14785,N_17571);
xnor U18681 (N_18681,N_15469,N_16626);
nor U18682 (N_18682,N_17374,N_15546);
xnor U18683 (N_18683,N_17917,N_16956);
or U18684 (N_18684,N_14031,N_16084);
nor U18685 (N_18685,N_15641,N_14194);
and U18686 (N_18686,N_15536,N_15274);
and U18687 (N_18687,N_15819,N_12843);
and U18688 (N_18688,N_15207,N_13464);
or U18689 (N_18689,N_14064,N_17669);
nor U18690 (N_18690,N_13934,N_13790);
xor U18691 (N_18691,N_16422,N_15214);
and U18692 (N_18692,N_14911,N_14876);
or U18693 (N_18693,N_15830,N_12595);
nand U18694 (N_18694,N_16929,N_12733);
or U18695 (N_18695,N_13106,N_13127);
and U18696 (N_18696,N_14003,N_14484);
xor U18697 (N_18697,N_16011,N_17429);
nor U18698 (N_18698,N_17331,N_12867);
nor U18699 (N_18699,N_14718,N_15408);
or U18700 (N_18700,N_15989,N_12105);
xor U18701 (N_18701,N_12436,N_13063);
nand U18702 (N_18702,N_15480,N_15984);
nor U18703 (N_18703,N_15577,N_13322);
nand U18704 (N_18704,N_15012,N_16655);
nor U18705 (N_18705,N_15593,N_15653);
nand U18706 (N_18706,N_17953,N_17220);
nand U18707 (N_18707,N_14849,N_16193);
or U18708 (N_18708,N_13201,N_13410);
nor U18709 (N_18709,N_15125,N_17847);
xor U18710 (N_18710,N_17035,N_16056);
xor U18711 (N_18711,N_16072,N_16678);
nor U18712 (N_18712,N_16222,N_12361);
nor U18713 (N_18713,N_17457,N_16570);
nor U18714 (N_18714,N_17783,N_16651);
xor U18715 (N_18715,N_17100,N_16606);
and U18716 (N_18716,N_12723,N_17416);
nor U18717 (N_18717,N_17991,N_14938);
nor U18718 (N_18718,N_14820,N_14574);
or U18719 (N_18719,N_13109,N_14183);
nor U18720 (N_18720,N_15756,N_12158);
and U18721 (N_18721,N_16795,N_17914);
xor U18722 (N_18722,N_17984,N_17566);
nor U18723 (N_18723,N_17277,N_17326);
nor U18724 (N_18724,N_16198,N_13242);
nand U18725 (N_18725,N_16562,N_14629);
or U18726 (N_18726,N_15943,N_14242);
nand U18727 (N_18727,N_15682,N_13916);
nand U18728 (N_18728,N_14909,N_14516);
or U18729 (N_18729,N_14971,N_16110);
or U18730 (N_18730,N_14905,N_14929);
and U18731 (N_18731,N_17412,N_17781);
nand U18732 (N_18732,N_15018,N_17723);
xor U18733 (N_18733,N_16445,N_14983);
xnor U18734 (N_18734,N_13144,N_12110);
nor U18735 (N_18735,N_13416,N_12171);
and U18736 (N_18736,N_15983,N_12854);
xnor U18737 (N_18737,N_12874,N_17353);
nor U18738 (N_18738,N_14188,N_14440);
nor U18739 (N_18739,N_16467,N_15916);
nor U18740 (N_18740,N_13487,N_13507);
and U18741 (N_18741,N_15672,N_17453);
nor U18742 (N_18742,N_16296,N_12959);
xor U18743 (N_18743,N_15774,N_13895);
xnor U18744 (N_18744,N_13588,N_17351);
and U18745 (N_18745,N_16002,N_13997);
xor U18746 (N_18746,N_14061,N_13836);
or U18747 (N_18747,N_12788,N_12562);
and U18748 (N_18748,N_16944,N_12388);
xnor U18749 (N_18749,N_16001,N_13523);
nand U18750 (N_18750,N_12056,N_13013);
xor U18751 (N_18751,N_17495,N_12692);
nand U18752 (N_18752,N_15787,N_13990);
xnor U18753 (N_18753,N_16354,N_13320);
and U18754 (N_18754,N_13873,N_15518);
or U18755 (N_18755,N_12456,N_14740);
or U18756 (N_18756,N_13634,N_13022);
and U18757 (N_18757,N_12547,N_17319);
xor U18758 (N_18758,N_15070,N_15974);
nand U18759 (N_18759,N_17870,N_15330);
and U18760 (N_18760,N_15590,N_16398);
and U18761 (N_18761,N_12648,N_15581);
and U18762 (N_18762,N_15190,N_17149);
nand U18763 (N_18763,N_13905,N_14997);
nor U18764 (N_18764,N_15949,N_13518);
and U18765 (N_18765,N_14987,N_15716);
nor U18766 (N_18766,N_15431,N_17814);
and U18767 (N_18767,N_17061,N_17371);
and U18768 (N_18768,N_15310,N_16405);
or U18769 (N_18769,N_17974,N_15385);
and U18770 (N_18770,N_15278,N_14295);
or U18771 (N_18771,N_15342,N_13179);
or U18772 (N_18772,N_12209,N_16585);
or U18773 (N_18773,N_16802,N_13781);
nor U18774 (N_18774,N_13777,N_13003);
or U18775 (N_18775,N_14272,N_15710);
xnor U18776 (N_18776,N_14837,N_12652);
nor U18777 (N_18777,N_12568,N_15624);
nor U18778 (N_18778,N_12683,N_15982);
and U18779 (N_18779,N_14669,N_14697);
xor U18780 (N_18780,N_15492,N_14533);
and U18781 (N_18781,N_17686,N_17342);
nand U18782 (N_18782,N_13316,N_12235);
or U18783 (N_18783,N_15976,N_13368);
nand U18784 (N_18784,N_13823,N_15257);
nand U18785 (N_18785,N_16985,N_17038);
xor U18786 (N_18786,N_16267,N_16154);
nor U18787 (N_18787,N_12520,N_17120);
nor U18788 (N_18788,N_14028,N_15013);
and U18789 (N_18789,N_15615,N_12291);
nor U18790 (N_18790,N_14042,N_14107);
or U18791 (N_18791,N_13413,N_15557);
nor U18792 (N_18792,N_16310,N_14449);
nor U18793 (N_18793,N_16968,N_16533);
nor U18794 (N_18794,N_17724,N_16576);
or U18795 (N_18795,N_14433,N_14534);
nand U18796 (N_18796,N_17297,N_16014);
nand U18797 (N_18797,N_13489,N_15947);
nand U18798 (N_18798,N_15333,N_12289);
nand U18799 (N_18799,N_13064,N_16740);
nor U18800 (N_18800,N_17309,N_17363);
xor U18801 (N_18801,N_12108,N_12440);
nor U18802 (N_18802,N_13508,N_13829);
nor U18803 (N_18803,N_15858,N_13014);
and U18804 (N_18804,N_14013,N_15633);
nand U18805 (N_18805,N_16940,N_14811);
nor U18806 (N_18806,N_15761,N_17489);
or U18807 (N_18807,N_12186,N_15453);
nand U18808 (N_18808,N_16926,N_14290);
or U18809 (N_18809,N_16064,N_13212);
and U18810 (N_18810,N_17971,N_13085);
or U18811 (N_18811,N_13911,N_12506);
or U18812 (N_18812,N_17504,N_12659);
xnor U18813 (N_18813,N_14947,N_13851);
and U18814 (N_18814,N_15101,N_12371);
or U18815 (N_18815,N_16451,N_16531);
or U18816 (N_18816,N_13740,N_12111);
nand U18817 (N_18817,N_14646,N_12731);
or U18818 (N_18818,N_16305,N_13794);
and U18819 (N_18819,N_12839,N_14527);
xnor U18820 (N_18820,N_14124,N_14452);
nor U18821 (N_18821,N_15420,N_12618);
xor U18822 (N_18822,N_12574,N_17892);
and U18823 (N_18823,N_12129,N_14639);
nand U18824 (N_18824,N_14330,N_12990);
or U18825 (N_18825,N_14335,N_12459);
or U18826 (N_18826,N_17703,N_12894);
xor U18827 (N_18827,N_16859,N_13232);
xnor U18828 (N_18828,N_12546,N_12425);
or U18829 (N_18829,N_12500,N_12010);
xor U18830 (N_18830,N_13261,N_17524);
and U18831 (N_18831,N_16703,N_16285);
nand U18832 (N_18832,N_15102,N_15414);
and U18833 (N_18833,N_14465,N_12993);
nor U18834 (N_18834,N_13741,N_15786);
nor U18835 (N_18835,N_12906,N_17623);
or U18836 (N_18836,N_17270,N_13471);
or U18837 (N_18837,N_16361,N_16942);
or U18838 (N_18838,N_17299,N_13262);
nand U18839 (N_18839,N_15733,N_12881);
or U18840 (N_18840,N_15666,N_13702);
nand U18841 (N_18841,N_14208,N_13123);
and U18842 (N_18842,N_17950,N_12890);
or U18843 (N_18843,N_16898,N_17179);
and U18844 (N_18844,N_14522,N_15415);
nor U18845 (N_18845,N_13744,N_12987);
nand U18846 (N_18846,N_16333,N_12679);
xnor U18847 (N_18847,N_13623,N_16320);
nor U18848 (N_18848,N_15097,N_14724);
or U18849 (N_18849,N_15450,N_14700);
and U18850 (N_18850,N_14235,N_15236);
nor U18851 (N_18851,N_12363,N_14826);
or U18852 (N_18852,N_15839,N_12495);
nand U18853 (N_18853,N_17135,N_13596);
or U18854 (N_18854,N_15042,N_13886);
nor U18855 (N_18855,N_15463,N_14207);
nor U18856 (N_18856,N_17451,N_13797);
xor U18857 (N_18857,N_12099,N_13371);
nand U18858 (N_18858,N_16719,N_15754);
xnor U18859 (N_18859,N_16020,N_14898);
nor U18860 (N_18860,N_17911,N_15586);
nor U18861 (N_18861,N_15890,N_17744);
nor U18862 (N_18862,N_15898,N_16732);
or U18863 (N_18863,N_15475,N_13210);
nor U18864 (N_18864,N_15747,N_16200);
nor U18865 (N_18865,N_12464,N_14858);
nand U18866 (N_18866,N_12114,N_16372);
and U18867 (N_18867,N_14202,N_13424);
and U18868 (N_18868,N_16062,N_16736);
nor U18869 (N_18869,N_15928,N_16257);
or U18870 (N_18870,N_15022,N_17315);
nand U18871 (N_18871,N_12510,N_13407);
xnor U18872 (N_18872,N_16043,N_13428);
and U18873 (N_18873,N_17601,N_15046);
and U18874 (N_18874,N_17449,N_13658);
xnor U18875 (N_18875,N_13700,N_13447);
or U18876 (N_18876,N_17050,N_12042);
xor U18877 (N_18877,N_17657,N_14380);
nor U18878 (N_18878,N_16992,N_16829);
xnor U18879 (N_18879,N_12473,N_15933);
xnor U18880 (N_18880,N_16715,N_16649);
nand U18881 (N_18881,N_12404,N_14882);
or U18882 (N_18882,N_16685,N_17172);
and U18883 (N_18883,N_12797,N_16067);
xor U18884 (N_18884,N_14083,N_14933);
xnor U18885 (N_18885,N_12693,N_14638);
or U18886 (N_18886,N_17114,N_14755);
and U18887 (N_18887,N_13986,N_13930);
nand U18888 (N_18888,N_12643,N_17129);
nor U18889 (N_18889,N_13177,N_16068);
nand U18890 (N_18890,N_12377,N_15580);
xnor U18891 (N_18891,N_15860,N_12742);
xor U18892 (N_18892,N_15512,N_12043);
nand U18893 (N_18893,N_12865,N_16166);
xor U18894 (N_18894,N_12479,N_12641);
nand U18895 (N_18895,N_17178,N_13077);
nand U18896 (N_18896,N_16131,N_12047);
or U18897 (N_18897,N_15872,N_13579);
nand U18898 (N_18898,N_12621,N_12308);
xor U18899 (N_18899,N_13470,N_17877);
xnor U18900 (N_18900,N_12265,N_14123);
nor U18901 (N_18901,N_17730,N_12259);
nand U18902 (N_18902,N_17418,N_16175);
nor U18903 (N_18903,N_15508,N_15179);
nand U18904 (N_18904,N_16330,N_12980);
or U18905 (N_18905,N_13812,N_12383);
nor U18906 (N_18906,N_15235,N_16648);
nor U18907 (N_18907,N_16092,N_16938);
or U18908 (N_18908,N_12860,N_12801);
xnor U18909 (N_18909,N_13967,N_12809);
nand U18910 (N_18910,N_14897,N_14577);
xor U18911 (N_18911,N_14231,N_14601);
or U18912 (N_18912,N_13400,N_15392);
nand U18913 (N_18913,N_12985,N_17134);
or U18914 (N_18914,N_14044,N_12452);
xnor U18915 (N_18915,N_16104,N_16179);
and U18916 (N_18916,N_15681,N_16662);
and U18917 (N_18917,N_16613,N_15250);
nand U18918 (N_18918,N_13863,N_13882);
and U18919 (N_18919,N_14835,N_13644);
nand U18920 (N_18920,N_17019,N_17320);
and U18921 (N_18921,N_13180,N_14481);
or U18922 (N_18922,N_17868,N_16885);
nor U18923 (N_18923,N_12372,N_12790);
nand U18924 (N_18924,N_16246,N_14323);
xnor U18925 (N_18925,N_15854,N_12727);
xnor U18926 (N_18926,N_12721,N_16007);
xnor U18927 (N_18927,N_15060,N_12170);
or U18928 (N_18928,N_17000,N_12518);
and U18929 (N_18929,N_16339,N_12405);
or U18930 (N_18930,N_15698,N_12513);
xnor U18931 (N_18931,N_14328,N_15007);
or U18932 (N_18932,N_12517,N_14749);
or U18933 (N_18933,N_12018,N_12751);
and U18934 (N_18934,N_12148,N_13280);
nand U18935 (N_18935,N_15359,N_14543);
nor U18936 (N_18936,N_14705,N_12994);
or U18937 (N_18937,N_16501,N_16610);
nand U18938 (N_18938,N_14798,N_16790);
nand U18939 (N_18939,N_16024,N_13254);
nand U18940 (N_18940,N_14551,N_13978);
nand U18941 (N_18941,N_17428,N_17167);
nor U18942 (N_18942,N_12636,N_15218);
xnor U18943 (N_18943,N_12507,N_14535);
xnor U18944 (N_18944,N_12519,N_12694);
nand U18945 (N_18945,N_13196,N_13587);
and U18946 (N_18946,N_15029,N_15182);
or U18947 (N_18947,N_17227,N_13617);
nor U18948 (N_18948,N_13759,N_16441);
xnor U18949 (N_18949,N_16122,N_13246);
nor U18950 (N_18950,N_16256,N_15228);
and U18951 (N_18951,N_13768,N_17517);
and U18952 (N_18952,N_13343,N_14887);
or U18953 (N_18953,N_16233,N_14747);
nor U18954 (N_18954,N_14297,N_13825);
xor U18955 (N_18955,N_14658,N_14243);
and U18956 (N_18956,N_13009,N_17037);
nor U18957 (N_18957,N_13015,N_12610);
nor U18958 (N_18958,N_14608,N_15129);
or U18959 (N_18959,N_17221,N_12573);
nor U18960 (N_18960,N_17443,N_13870);
nand U18961 (N_18961,N_12848,N_12415);
and U18962 (N_18962,N_14960,N_12931);
nand U18963 (N_18963,N_17954,N_15679);
nor U18964 (N_18964,N_12208,N_16928);
xnor U18965 (N_18965,N_16918,N_13604);
or U18966 (N_18966,N_12437,N_12718);
or U18967 (N_18967,N_17280,N_16464);
or U18968 (N_18968,N_17263,N_15997);
and U18969 (N_18969,N_13281,N_15398);
nand U18970 (N_18970,N_15703,N_17341);
nand U18971 (N_18971,N_12077,N_13169);
nor U18972 (N_18972,N_14684,N_14797);
or U18973 (N_18973,N_15994,N_14151);
xor U18974 (N_18974,N_16221,N_12349);
nand U18975 (N_18975,N_13660,N_17112);
nor U18976 (N_18976,N_15706,N_14196);
or U18977 (N_18977,N_14919,N_16987);
and U18978 (N_18978,N_13052,N_15276);
and U18979 (N_18979,N_14052,N_12470);
xnor U18980 (N_18980,N_12970,N_13843);
xnor U18981 (N_18981,N_12323,N_15443);
and U18982 (N_18982,N_16268,N_15511);
and U18983 (N_18983,N_16275,N_12492);
or U18984 (N_18984,N_17751,N_14968);
or U18985 (N_18985,N_16991,N_15020);
and U18986 (N_18986,N_15874,N_15962);
or U18987 (N_18987,N_12499,N_13969);
nand U18988 (N_18988,N_14403,N_16998);
nor U18989 (N_18989,N_17828,N_13222);
nor U18990 (N_18990,N_13814,N_16192);
nor U18991 (N_18991,N_15242,N_16298);
xor U18992 (N_18992,N_12269,N_12498);
xor U18993 (N_18993,N_16088,N_16114);
and U18994 (N_18994,N_15080,N_12217);
or U18995 (N_18995,N_13323,N_16560);
nand U18996 (N_18996,N_14792,N_12957);
xor U18997 (N_18997,N_14224,N_14000);
nor U18998 (N_18998,N_17414,N_17283);
and U18999 (N_18999,N_17180,N_12367);
xnor U19000 (N_19000,N_16587,N_17662);
nand U19001 (N_19001,N_15357,N_16485);
xor U19002 (N_19002,N_15755,N_16629);
nor U19003 (N_19003,N_14432,N_15572);
and U19004 (N_19004,N_13787,N_15468);
xnor U19005 (N_19005,N_16567,N_17483);
or U19006 (N_19006,N_12998,N_13576);
or U19007 (N_19007,N_12973,N_14352);
nor U19008 (N_19008,N_12139,N_14881);
nor U19009 (N_19009,N_16409,N_16047);
nor U19010 (N_19010,N_17895,N_16798);
and U19011 (N_19011,N_12389,N_12583);
or U19012 (N_19012,N_17515,N_14071);
nand U19013 (N_19013,N_13563,N_17964);
nor U19014 (N_19014,N_17444,N_13753);
nor U19015 (N_19015,N_13031,N_16937);
xor U19016 (N_19016,N_13445,N_15794);
xor U19017 (N_19017,N_15552,N_16819);
and U19018 (N_19018,N_12882,N_17021);
nand U19019 (N_19019,N_14065,N_15320);
or U19020 (N_19020,N_13202,N_17447);
or U19021 (N_19021,N_16403,N_14506);
nor U19022 (N_19022,N_14784,N_13067);
or U19023 (N_19023,N_12199,N_12151);
and U19024 (N_19024,N_12825,N_17125);
xnor U19025 (N_19025,N_16120,N_14402);
nor U19026 (N_19026,N_17041,N_15623);
or U19027 (N_19027,N_12941,N_13376);
nand U19028 (N_19028,N_14787,N_16215);
xor U19029 (N_19029,N_13364,N_15039);
and U19030 (N_19030,N_15040,N_17933);
or U19031 (N_19031,N_14879,N_15584);
or U19032 (N_19032,N_16118,N_17383);
or U19033 (N_19033,N_15560,N_15965);
xor U19034 (N_19034,N_14447,N_16049);
xor U19035 (N_19035,N_16309,N_15021);
or U19036 (N_19036,N_14988,N_16578);
nor U19037 (N_19037,N_17204,N_14256);
nand U19038 (N_19038,N_13574,N_12684);
nor U19039 (N_19039,N_17989,N_17332);
and U19040 (N_19040,N_16597,N_15630);
xnor U19041 (N_19041,N_13586,N_14341);
nand U19042 (N_19042,N_17369,N_14404);
nand U19043 (N_19043,N_15156,N_14722);
nor U19044 (N_19044,N_13748,N_15472);
or U19045 (N_19045,N_15501,N_16579);
and U19046 (N_19046,N_13450,N_17235);
xor U19047 (N_19047,N_13217,N_13831);
xnor U19048 (N_19048,N_12340,N_16889);
nand U19049 (N_19049,N_16659,N_15315);
nand U19050 (N_19050,N_17284,N_15405);
nor U19051 (N_19051,N_16009,N_16406);
nor U19052 (N_19052,N_16394,N_12401);
or U19053 (N_19053,N_16375,N_17644);
or U19054 (N_19054,N_13684,N_15724);
xor U19055 (N_19055,N_14827,N_12034);
or U19056 (N_19056,N_14259,N_16123);
xnor U19057 (N_19057,N_16586,N_17645);
or U19058 (N_19058,N_14075,N_12488);
or U19059 (N_19059,N_15960,N_14309);
xor U19060 (N_19060,N_13370,N_16833);
nand U19061 (N_19061,N_13800,N_16129);
nor U19062 (N_19062,N_14743,N_17698);
or U19063 (N_19063,N_14187,N_13054);
or U19064 (N_19064,N_17060,N_17249);
nor U19065 (N_19065,N_12181,N_16866);
xnor U19066 (N_19066,N_17826,N_12020);
or U19067 (N_19067,N_16214,N_12740);
xnor U19068 (N_19068,N_17056,N_17308);
or U19069 (N_19069,N_15099,N_13453);
and U19070 (N_19070,N_15193,N_12302);
or U19071 (N_19071,N_13688,N_13799);
nor U19072 (N_19072,N_13821,N_14155);
nand U19073 (N_19073,N_15516,N_16100);
nor U19074 (N_19074,N_13665,N_14510);
and U19075 (N_19075,N_16679,N_12237);
nor U19076 (N_19076,N_17970,N_17008);
xor U19077 (N_19077,N_15302,N_17878);
or U19078 (N_19078,N_14951,N_17388);
xnor U19079 (N_19079,N_12124,N_13089);
or U19080 (N_19080,N_15073,N_17628);
and U19081 (N_19081,N_15806,N_12101);
or U19082 (N_19082,N_14270,N_17107);
or U19083 (N_19083,N_15715,N_17052);
nand U19084 (N_19084,N_17908,N_14935);
nand U19085 (N_19085,N_14812,N_15158);
or U19086 (N_19086,N_12455,N_12668);
and U19087 (N_19087,N_13710,N_13703);
nor U19088 (N_19088,N_12240,N_17939);
and U19089 (N_19089,N_14277,N_12862);
nor U19090 (N_19090,N_15183,N_12131);
xor U19091 (N_19091,N_12802,N_14240);
xnor U19092 (N_19092,N_12294,N_17716);
nor U19093 (N_19093,N_17295,N_14995);
nand U19094 (N_19094,N_13274,N_17615);
nor U19095 (N_19095,N_16428,N_15622);
and U19096 (N_19096,N_15476,N_14010);
or U19097 (N_19097,N_15523,N_16949);
and U19098 (N_19098,N_15541,N_17286);
nand U19099 (N_19099,N_15106,N_17560);
and U19100 (N_19100,N_13589,N_17549);
or U19101 (N_19101,N_15919,N_17477);
and U19102 (N_19102,N_16698,N_14863);
nand U19103 (N_19103,N_15568,N_12178);
nor U19104 (N_19104,N_16706,N_17627);
and U19105 (N_19105,N_16948,N_14972);
nor U19106 (N_19106,N_17803,N_17681);
nand U19107 (N_19107,N_15221,N_16483);
or U19108 (N_19108,N_16289,N_15538);
nand U19109 (N_19109,N_14332,N_15196);
nand U19110 (N_19110,N_13980,N_13198);
nor U19111 (N_19111,N_16552,N_13504);
xor U19112 (N_19112,N_17062,N_17636);
nor U19113 (N_19113,N_17992,N_14041);
and U19114 (N_19114,N_12944,N_17242);
nand U19115 (N_19115,N_12443,N_16337);
or U19116 (N_19116,N_12982,N_14038);
xor U19117 (N_19117,N_14788,N_13467);
xnor U19118 (N_19118,N_17697,N_15396);
and U19119 (N_19119,N_13084,N_16537);
or U19120 (N_19120,N_12930,N_16830);
nor U19121 (N_19121,N_16702,N_17508);
nor U19122 (N_19122,N_15280,N_13229);
or U19123 (N_19123,N_15673,N_15553);
nor U19124 (N_19124,N_12272,N_14206);
nor U19125 (N_19125,N_13435,N_14122);
nand U19126 (N_19126,N_17261,N_14772);
and U19127 (N_19127,N_17482,N_15944);
nand U19128 (N_19128,N_17667,N_13301);
nor U19129 (N_19129,N_17459,N_13926);
nor U19130 (N_19130,N_17175,N_15948);
nor U19131 (N_19131,N_16331,N_13183);
nand U19132 (N_19132,N_16460,N_13430);
xnor U19133 (N_19133,N_14893,N_17287);
and U19134 (N_19134,N_13940,N_16042);
nand U19135 (N_19135,N_12748,N_17543);
nor U19136 (N_19136,N_12133,N_15667);
xor U19137 (N_19137,N_16477,N_12107);
nand U19138 (N_19138,N_13867,N_17026);
or U19139 (N_19139,N_12091,N_16784);
xnor U19140 (N_19140,N_12397,N_14850);
xnor U19141 (N_19141,N_17339,N_12048);
nor U19142 (N_19142,N_14948,N_13506);
or U19143 (N_19143,N_17650,N_17156);
nand U19144 (N_19144,N_16498,N_14729);
nor U19145 (N_19145,N_17445,N_14198);
nand U19146 (N_19146,N_16090,N_12711);
xor U19147 (N_19147,N_16895,N_17205);
and U19148 (N_19148,N_13419,N_13965);
and U19149 (N_19149,N_17766,N_14570);
nor U19150 (N_19150,N_12630,N_16542);
or U19151 (N_19151,N_17460,N_15056);
xnor U19152 (N_19152,N_13473,N_13696);
xnor U19153 (N_19153,N_13290,N_17252);
or U19154 (N_19154,N_13330,N_15587);
xnor U19155 (N_19155,N_17709,N_13958);
nand U19156 (N_19156,N_15514,N_15882);
nor U19157 (N_19157,N_12029,N_13762);
nand U19158 (N_19158,N_17831,N_14766);
or U19159 (N_19159,N_12864,N_13171);
nand U19160 (N_19160,N_14716,N_12811);
nand U19161 (N_19161,N_12180,N_13906);
and U19162 (N_19162,N_15910,N_12887);
nor U19163 (N_19163,N_16295,N_13097);
nand U19164 (N_19164,N_15339,N_12135);
or U19165 (N_19165,N_14651,N_14655);
and U19166 (N_19166,N_15262,N_15437);
nand U19167 (N_19167,N_15059,N_16093);
xor U19168 (N_19168,N_12410,N_16417);
xnor U19169 (N_19169,N_17588,N_17556);
xor U19170 (N_19170,N_16227,N_15290);
nand U19171 (N_19171,N_13233,N_14390);
nand U19172 (N_19172,N_15801,N_16905);
nor U19173 (N_19173,N_12531,N_13695);
xnor U19174 (N_19174,N_17330,N_13939);
and U19175 (N_19175,N_16584,N_17301);
nor U19176 (N_19176,N_14524,N_13088);
nor U19177 (N_19177,N_14825,N_15896);
nor U19178 (N_19178,N_17382,N_17862);
or U19179 (N_19179,N_13789,N_13315);
nand U19180 (N_19180,N_13907,N_16984);
and U19181 (N_19181,N_12335,N_12717);
nor U19182 (N_19182,N_17213,N_13184);
and U19183 (N_19183,N_12714,N_15204);
nand U19184 (N_19184,N_12812,N_15900);
and U19185 (N_19185,N_13011,N_16575);
xor U19186 (N_19186,N_13279,N_15588);
nor U19187 (N_19187,N_17082,N_16724);
and U19188 (N_19188,N_17476,N_13838);
nand U19189 (N_19189,N_12953,N_17057);
and U19190 (N_19190,N_13824,N_15186);
nand U19191 (N_19191,N_16204,N_12080);
nor U19192 (N_19192,N_16742,N_16292);
and U19193 (N_19193,N_14426,N_13631);
nor U19194 (N_19194,N_17782,N_13505);
nor U19195 (N_19195,N_12543,N_14813);
or U19196 (N_19196,N_16174,N_17025);
xnor U19197 (N_19197,N_17618,N_13692);
nand U19198 (N_19198,N_16822,N_16045);
xor U19199 (N_19199,N_15421,N_17855);
nand U19200 (N_19200,N_12761,N_14848);
xnor U19201 (N_19201,N_16857,N_13165);
nand U19202 (N_19202,N_12468,N_15985);
nand U19203 (N_19203,N_12662,N_13178);
and U19204 (N_19204,N_17364,N_16608);
and U19205 (N_19205,N_13076,N_12369);
nand U19206 (N_19206,N_14586,N_12145);
nand U19207 (N_19207,N_12037,N_15137);
nand U19208 (N_19208,N_17811,N_13035);
or U19209 (N_19209,N_12206,N_13115);
or U19210 (N_19210,N_14679,N_14861);
xnor U19211 (N_19211,N_13963,N_16202);
nor U19212 (N_19212,N_15619,N_15072);
nor U19213 (N_19213,N_14153,N_12428);
nor U19214 (N_19214,N_12341,N_15995);
or U19215 (N_19215,N_14096,N_15719);
nor U19216 (N_19216,N_15124,N_17346);
nand U19217 (N_19217,N_14667,N_16448);
xnor U19218 (N_19218,N_14439,N_17492);
or U19219 (N_19219,N_12260,N_12121);
or U19220 (N_19220,N_14215,N_16003);
nor U19221 (N_19221,N_16571,N_17192);
and U19222 (N_19222,N_13185,N_16708);
xor U19223 (N_19223,N_12281,N_16941);
and U19224 (N_19224,N_17471,N_15203);
nand U19225 (N_19225,N_17626,N_13216);
nand U19226 (N_19226,N_17539,N_16910);
nand U19227 (N_19227,N_13192,N_15436);
or U19228 (N_19228,N_17596,N_14293);
and U19229 (N_19229,N_17921,N_14565);
and U19230 (N_19230,N_13380,N_15146);
and U19231 (N_19231,N_17470,N_13098);
nor U19232 (N_19232,N_13815,N_16674);
xnor U19233 (N_19233,N_15138,N_12039);
xor U19234 (N_19234,N_15239,N_17200);
xnor U19235 (N_19235,N_17217,N_14210);
xnor U19236 (N_19236,N_16901,N_12194);
nand U19237 (N_19237,N_13156,N_16877);
nand U19238 (N_19238,N_13599,N_14068);
xnor U19239 (N_19239,N_13131,N_12084);
or U19240 (N_19240,N_13575,N_17164);
or U19241 (N_19241,N_12481,N_17762);
and U19242 (N_19242,N_15119,N_16470);
nand U19243 (N_19243,N_12655,N_17234);
and U19244 (N_19244,N_17685,N_15522);
nor U19245 (N_19245,N_15449,N_16783);
and U19246 (N_19246,N_16103,N_12936);
nand U19247 (N_19247,N_17957,N_15005);
nand U19248 (N_19248,N_17948,N_14189);
xor U19249 (N_19249,N_16149,N_17073);
or U19250 (N_19250,N_17048,N_13947);
and U19251 (N_19251,N_12676,N_13892);
xnor U19252 (N_19252,N_15542,N_14291);
xor U19253 (N_19253,N_12577,N_16180);
or U19254 (N_19254,N_15730,N_15937);
nand U19255 (N_19255,N_12858,N_16112);
xnor U19256 (N_19256,N_14664,N_14347);
nor U19257 (N_19257,N_16031,N_13785);
or U19258 (N_19258,N_17421,N_13743);
or U19259 (N_19259,N_16852,N_16273);
or U19260 (N_19260,N_15135,N_17532);
or U19261 (N_19261,N_13713,N_14338);
and U19262 (N_19262,N_16663,N_12965);
xnor U19263 (N_19263,N_14102,N_13834);
and U19264 (N_19264,N_14868,N_15837);
or U19265 (N_19265,N_17613,N_14327);
xnor U19266 (N_19266,N_17345,N_13534);
and U19267 (N_19267,N_12935,N_14915);
and U19268 (N_19268,N_15201,N_12738);
nand U19269 (N_19269,N_13633,N_16313);
xnor U19270 (N_19270,N_15901,N_15504);
nor U19271 (N_19271,N_15305,N_13211);
or U19272 (N_19272,N_15304,N_14872);
and U19273 (N_19273,N_15799,N_15675);
xor U19274 (N_19274,N_13952,N_16397);
nor U19275 (N_19275,N_12137,N_16855);
and U19276 (N_19276,N_14182,N_17219);
and U19277 (N_19277,N_14579,N_16039);
or U19278 (N_19278,N_16474,N_17940);
and U19279 (N_19279,N_14211,N_17432);
and U19280 (N_19280,N_17656,N_13652);
nand U19281 (N_19281,N_16541,N_17032);
or U19282 (N_19282,N_14007,N_13600);
and U19283 (N_19283,N_12850,N_13415);
xnor U19284 (N_19284,N_15294,N_15090);
nand U19285 (N_19285,N_16490,N_13630);
xnor U19286 (N_19286,N_15879,N_14022);
or U19287 (N_19287,N_14545,N_17720);
nor U19288 (N_19288,N_14026,N_13529);
xor U19289 (N_19289,N_15911,N_13159);
or U19290 (N_19290,N_13474,N_17011);
and U19291 (N_19291,N_17337,N_14758);
xor U19292 (N_19292,N_16437,N_17336);
and U19293 (N_19293,N_15071,N_15484);
nor U19294 (N_19294,N_17861,N_12041);
nor U19295 (N_19295,N_14015,N_17088);
nand U19296 (N_19296,N_14824,N_16945);
nor U19297 (N_19297,N_14696,N_13369);
nand U19298 (N_19298,N_15825,N_16726);
nor U19299 (N_19299,N_15852,N_12537);
and U19300 (N_19300,N_13347,N_12215);
or U19301 (N_19301,N_14472,N_16411);
and U19302 (N_19302,N_14662,N_15084);
or U19303 (N_19303,N_16287,N_13459);
nand U19304 (N_19304,N_14874,N_15863);
and U19305 (N_19305,N_12750,N_13581);
nor U19306 (N_19306,N_16240,N_15654);
and U19307 (N_19307,N_12515,N_16913);
and U19308 (N_19308,N_14732,N_15027);
or U19309 (N_19309,N_14133,N_17413);
xnor U19310 (N_19310,N_15939,N_16171);
and U19311 (N_19311,N_16026,N_14781);
xnor U19312 (N_19312,N_14518,N_12570);
xnor U19313 (N_19313,N_14558,N_14529);
xor U19314 (N_19314,N_16057,N_13883);
or U19315 (N_19315,N_15789,N_15316);
and U19316 (N_19316,N_14125,N_17415);
and U19317 (N_19317,N_13285,N_12252);
nor U19318 (N_19318,N_17500,N_15992);
nor U19319 (N_19319,N_14305,N_13104);
nand U19320 (N_19320,N_16494,N_13769);
xor U19321 (N_19321,N_16779,N_16522);
nand U19322 (N_19322,N_12651,N_12258);
and U19323 (N_19323,N_12736,N_13855);
nor U19324 (N_19324,N_14702,N_15753);
xor U19325 (N_19325,N_13048,N_13037);
or U19326 (N_19326,N_17098,N_15371);
xor U19327 (N_19327,N_13782,N_16943);
xnor U19328 (N_19328,N_14306,N_16646);
or U19329 (N_19329,N_15440,N_12503);
xor U19330 (N_19330,N_17479,N_16495);
nor U19331 (N_19331,N_14852,N_12204);
nand U19332 (N_19332,N_13341,N_15791);
or U19333 (N_19333,N_15411,N_12580);
nand U19334 (N_19334,N_12735,N_16923);
and U19335 (N_19335,N_14217,N_17109);
nor U19336 (N_19336,N_12028,N_13864);
xnor U19337 (N_19337,N_14393,N_17731);
and U19338 (N_19338,N_17606,N_15728);
nor U19339 (N_19339,N_14103,N_14663);
and U19340 (N_19340,N_16279,N_12504);
and U19341 (N_19341,N_12184,N_14435);
nor U19342 (N_19342,N_14949,N_12853);
nor U19343 (N_19343,N_14314,N_17176);
nand U19344 (N_19344,N_12257,N_13182);
xnor U19345 (N_19345,N_13539,N_13977);
xnor U19346 (N_19346,N_12763,N_14121);
nor U19347 (N_19347,N_13454,N_12477);
nand U19348 (N_19348,N_16119,N_14649);
or U19349 (N_19349,N_14666,N_15884);
nor U19350 (N_19350,N_16601,N_16457);
nor U19351 (N_19351,N_12314,N_17182);
nor U19352 (N_19352,N_15249,N_13608);
xnor U19353 (N_19353,N_16489,N_14581);
and U19354 (N_19354,N_17400,N_13973);
nor U19355 (N_19355,N_17757,N_14319);
xor U19356 (N_19356,N_15762,N_17452);
and U19357 (N_19357,N_12997,N_14019);
and U19358 (N_19358,N_14017,N_16603);
nor U19359 (N_19359,N_12526,N_12918);
and U19360 (N_19360,N_17784,N_13324);
nand U19361 (N_19361,N_17375,N_16547);
nor U19362 (N_19362,N_17422,N_15627);
nand U19363 (N_19363,N_17540,N_12490);
xnor U19364 (N_19364,N_14778,N_17882);
or U19365 (N_19365,N_17480,N_13786);
and U19366 (N_19366,N_12466,N_12545);
xnor U19367 (N_19367,N_13657,N_16728);
nor U19368 (N_19368,N_14770,N_16258);
xor U19369 (N_19369,N_16291,N_14279);
nor U19370 (N_19370,N_13005,N_17367);
xor U19371 (N_19371,N_17721,N_14006);
nor U19372 (N_19372,N_15929,N_12635);
nor U19373 (N_19373,N_17228,N_17247);
nand U19374 (N_19374,N_15378,N_12779);
and U19375 (N_19375,N_15990,N_13312);
nor U19376 (N_19376,N_15112,N_14027);
and U19377 (N_19377,N_16573,N_17608);
xor U19378 (N_19378,N_15885,N_13227);
nor U19379 (N_19379,N_16604,N_13399);
nor U19380 (N_19380,N_13306,N_17115);
xor U19381 (N_19381,N_13403,N_15256);
nand U19382 (N_19382,N_13733,N_17250);
xor U19383 (N_19383,N_15629,N_13601);
nand U19384 (N_19384,N_16675,N_13972);
xnor U19385 (N_19385,N_17126,N_12304);
nand U19386 (N_19386,N_15091,N_17670);
or U19387 (N_19387,N_13803,N_13530);
nand U19388 (N_19388,N_12247,N_16453);
nor U19389 (N_19389,N_12737,N_12331);
nor U19390 (N_19390,N_16553,N_17253);
nand U19391 (N_19391,N_13956,N_17257);
or U19392 (N_19392,N_12913,N_12087);
and U19393 (N_19393,N_12085,N_16681);
nand U19394 (N_19394,N_15065,N_13443);
or U19395 (N_19395,N_13778,N_14612);
xor U19396 (N_19396,N_13175,N_16886);
nor U19397 (N_19397,N_17290,N_15384);
or U19398 (N_19398,N_12273,N_15605);
and U19399 (N_19399,N_14712,N_16660);
and U19400 (N_19400,N_14636,N_14412);
or U19401 (N_19401,N_16892,N_15474);
or U19402 (N_19402,N_16815,N_15487);
and U19403 (N_19403,N_17024,N_16906);
nand U19404 (N_19404,N_17611,N_16116);
or U19405 (N_19405,N_15416,N_14264);
and U19406 (N_19406,N_15430,N_14564);
nor U19407 (N_19407,N_13398,N_15711);
nand U19408 (N_19408,N_13335,N_14764);
nor U19409 (N_19409,N_16170,N_15979);
and U19410 (N_19410,N_17776,N_14087);
nand U19411 (N_19411,N_13258,N_17946);
xnor U19412 (N_19412,N_14425,N_13983);
nor U19413 (N_19413,N_14262,N_13847);
nand U19414 (N_19414,N_17348,N_14002);
and U19415 (N_19415,N_17599,N_12337);
or U19416 (N_19416,N_15243,N_16376);
xnor U19417 (N_19417,N_17741,N_14966);
nor U19418 (N_19418,N_14841,N_14495);
and U19419 (N_19419,N_15074,N_15987);
xor U19420 (N_19420,N_14967,N_13992);
nand U19421 (N_19421,N_14191,N_13342);
xor U19422 (N_19422,N_16101,N_14092);
xor U19423 (N_19423,N_15604,N_12926);
xnor U19424 (N_19424,N_14269,N_15778);
xor U19425 (N_19425,N_15932,N_14040);
nor U19426 (N_19426,N_16499,N_16128);
xnor U19427 (N_19427,N_15035,N_16187);
nor U19428 (N_19428,N_12146,N_17344);
and U19429 (N_19429,N_17637,N_14170);
xor U19430 (N_19430,N_15509,N_15695);
nand U19431 (N_19431,N_16544,N_13701);
nor U19432 (N_19432,N_15085,N_12609);
and U19433 (N_19433,N_13527,N_17796);
nand U19434 (N_19434,N_13602,N_17066);
nand U19435 (N_19435,N_15705,N_16556);
xor U19436 (N_19436,N_17159,N_17490);
and U19437 (N_19437,N_13948,N_12567);
nor U19438 (N_19438,N_16927,N_15258);
nand U19439 (N_19439,N_12321,N_15834);
nor U19440 (N_19440,N_15958,N_14392);
nand U19441 (N_19441,N_12590,N_14688);
nor U19442 (N_19442,N_17488,N_14228);
or U19443 (N_19443,N_14505,N_12290);
and U19444 (N_19444,N_12976,N_17423);
xnor U19445 (N_19445,N_15532,N_14261);
nor U19446 (N_19446,N_17124,N_15721);
and U19447 (N_19447,N_14448,N_14632);
and U19448 (N_19448,N_13385,N_13072);
nand U19449 (N_19449,N_13935,N_14350);
nand U19450 (N_19450,N_16368,N_16439);
nand U19451 (N_19451,N_13377,N_15840);
xnor U19452 (N_19452,N_14587,N_13780);
nor U19453 (N_19453,N_12878,N_13808);
nand U19454 (N_19454,N_17582,N_15404);
and U19455 (N_19455,N_16691,N_13605);
xnor U19456 (N_19456,N_14956,N_13205);
and U19457 (N_19457,N_13573,N_15206);
nor U19458 (N_19458,N_17725,N_12293);
or U19459 (N_19459,N_16500,N_14298);
nand U19460 (N_19460,N_17455,N_16076);
nand U19461 (N_19461,N_15130,N_16095);
nor U19462 (N_19462,N_13826,N_16444);
or U19463 (N_19463,N_16532,N_14954);
xor U19464 (N_19464,N_12154,N_17289);
xnor U19465 (N_19465,N_16459,N_13356);
or U19466 (N_19466,N_16251,N_15550);
and U19467 (N_19467,N_13672,N_14386);
or U19468 (N_19468,N_12666,N_16785);
or U19469 (N_19469,N_15240,N_12353);
nand U19470 (N_19470,N_16037,N_13402);
nor U19471 (N_19471,N_16343,N_16218);
or U19472 (N_19472,N_16588,N_17023);
or U19473 (N_19473,N_16514,N_12118);
nand U19474 (N_19474,N_14363,N_12868);
nor U19475 (N_19475,N_14746,N_12051);
and U19476 (N_19476,N_16894,N_12173);
and U19477 (N_19477,N_15301,N_13909);
and U19478 (N_19478,N_12924,N_16754);
nand U19479 (N_19479,N_16506,N_17141);
or U19480 (N_19480,N_17754,N_17568);
nor U19481 (N_19481,N_15521,N_14763);
nand U19482 (N_19482,N_15530,N_13805);
nor U19483 (N_19483,N_15482,N_17302);
and U19484 (N_19484,N_14660,N_16561);
or U19485 (N_19485,N_15212,N_13166);
or U19486 (N_19486,N_14200,N_13172);
xor U19487 (N_19487,N_14361,N_14143);
or U19488 (N_19488,N_12132,N_16976);
xnor U19489 (N_19489,N_14056,N_13541);
and U19490 (N_19490,N_16799,N_12327);
or U19491 (N_19491,N_13510,N_15094);
and U19492 (N_19492,N_13339,N_17655);
nor U19493 (N_19493,N_17823,N_17999);
xor U19494 (N_19494,N_12708,N_14466);
nand U19495 (N_19495,N_14486,N_16605);
and U19496 (N_19496,N_16596,N_12394);
nor U19497 (N_19497,N_15820,N_12951);
nor U19498 (N_19498,N_12193,N_15208);
nor U19499 (N_19499,N_17717,N_16879);
or U19500 (N_19500,N_16184,N_14349);
xnor U19501 (N_19501,N_17116,N_15277);
or U19502 (N_19502,N_15950,N_17366);
xor U19503 (N_19503,N_17666,N_16450);
nand U19504 (N_19504,N_14831,N_12557);
and U19505 (N_19505,N_13525,N_14193);
xnor U19506 (N_19506,N_17742,N_14048);
nand U19507 (N_19507,N_12851,N_13158);
nand U19508 (N_19508,N_16687,N_13511);
and U19509 (N_19509,N_15025,N_16236);
nand U19510 (N_19510,N_17046,N_12267);
nand U19511 (N_19511,N_13682,N_15354);
xor U19512 (N_19512,N_14227,N_13902);
and U19513 (N_19513,N_15089,N_15565);
xnor U19514 (N_19514,N_15386,N_14801);
nor U19515 (N_19515,N_14686,N_14681);
nor U19516 (N_19516,N_13524,N_16636);
and U19517 (N_19517,N_13497,N_17947);
nand U19518 (N_19518,N_16794,N_17045);
and U19519 (N_19519,N_17328,N_12625);
or U19520 (N_19520,N_14368,N_17527);
or U19521 (N_19521,N_14782,N_17230);
xor U19522 (N_19522,N_15967,N_16806);
xnor U19523 (N_19523,N_13313,N_16040);
and U19524 (N_19524,N_15893,N_13118);
nor U19525 (N_19525,N_12803,N_17865);
nor U19526 (N_19526,N_16102,N_13160);
xnor U19527 (N_19527,N_12122,N_17987);
and U19528 (N_19528,N_15676,N_16108);
or U19529 (N_19529,N_14822,N_14507);
nand U19530 (N_19530,N_14768,N_14902);
or U19531 (N_19531,N_14585,N_12552);
and U19532 (N_19532,N_14173,N_16868);
xnor U19533 (N_19533,N_16755,N_12730);
xnor U19534 (N_19534,N_15351,N_15010);
nor U19535 (N_19535,N_17834,N_15999);
or U19536 (N_19536,N_16558,N_13272);
or U19537 (N_19537,N_17680,N_15307);
and U19538 (N_19538,N_17665,N_15171);
nand U19539 (N_19539,N_15303,N_15748);
or U19540 (N_19540,N_17872,N_15864);
or U19541 (N_19541,N_14162,N_12222);
and U19542 (N_19542,N_13455,N_16505);
nor U19543 (N_19543,N_12849,N_16245);
nand U19544 (N_19544,N_14490,N_14894);
and U19545 (N_19545,N_15161,N_16364);
xor U19546 (N_19546,N_14865,N_14165);
xnor U19547 (N_19547,N_17672,N_14583);
xnor U19548 (N_19548,N_17695,N_17822);
xnor U19549 (N_19549,N_15388,N_12033);
or U19550 (N_19550,N_17064,N_17647);
nor U19551 (N_19551,N_12725,N_13500);
nand U19552 (N_19552,N_17154,N_12724);
and U19553 (N_19553,N_13625,N_17979);
or U19554 (N_19554,N_15489,N_16750);
or U19555 (N_19555,N_17473,N_15107);
nor U19556 (N_19556,N_15111,N_17998);
nor U19557 (N_19557,N_12014,N_12050);
nand U19558 (N_19558,N_17874,N_14444);
or U19559 (N_19559,N_13208,N_12061);
nand U19560 (N_19560,N_12191,N_15656);
nand U19561 (N_19561,N_15760,N_16209);
nor U19562 (N_19562,N_16212,N_14708);
or U19563 (N_19563,N_12691,N_14077);
nor U19564 (N_19564,N_12846,N_16974);
nand U19565 (N_19565,N_14959,N_17838);
and U19566 (N_19566,N_13571,N_12808);
xor U19567 (N_19567,N_15562,N_15168);
nand U19568 (N_19568,N_17222,N_15175);
and U19569 (N_19569,N_13409,N_17275);
nand U19570 (N_19570,N_17969,N_13135);
nor U19571 (N_19571,N_12904,N_13300);
nor U19572 (N_19572,N_13355,N_16317);
or U19573 (N_19573,N_16725,N_16803);
xor U19574 (N_19574,N_13042,N_12952);
nor U19575 (N_19575,N_14619,N_16735);
xor U19576 (N_19576,N_12231,N_17519);
xor U19577 (N_19577,N_13044,N_15938);
xor U19578 (N_19578,N_14617,N_16842);
xnor U19579 (N_19579,N_16232,N_12866);
or U19580 (N_19580,N_14213,N_13036);
nand U19581 (N_19581,N_14115,N_15318);
or U19582 (N_19582,N_15053,N_17956);
nor U19583 (N_19583,N_17393,N_14158);
and U19584 (N_19584,N_14442,N_12478);
or U19585 (N_19585,N_16527,N_16958);
xnor U19586 (N_19586,N_15904,N_12960);
nand U19587 (N_19587,N_17362,N_16934);
nand U19588 (N_19588,N_12859,N_16535);
nand U19589 (N_19589,N_17379,N_13820);
and U19590 (N_19590,N_14568,N_12805);
nor U19591 (N_19591,N_16113,N_13749);
or U19592 (N_19592,N_15796,N_12115);
xor U19593 (N_19593,N_13080,N_17474);
nor U19594 (N_19594,N_12075,N_13577);
nor U19595 (N_19595,N_15069,N_16066);
nor U19596 (N_19596,N_12760,N_17529);
nand U19597 (N_19597,N_14642,N_12243);
or U19598 (N_19598,N_14362,N_15595);
nand U19599 (N_19599,N_16288,N_13971);
or U19600 (N_19600,N_13982,N_12631);
nand U19601 (N_19601,N_13928,N_14671);
and U19602 (N_19602,N_14691,N_15803);
and U19603 (N_19603,N_14376,N_12221);
and U19604 (N_19604,N_16286,N_15481);
and U19605 (N_19605,N_16932,N_17852);
nor U19606 (N_19606,N_16058,N_16607);
nor U19607 (N_19607,N_17858,N_13477);
and U19608 (N_19608,N_16530,N_15868);
nor U19609 (N_19609,N_12292,N_14857);
nor U19610 (N_19610,N_14965,N_14373);
nand U19611 (N_19611,N_16438,N_14316);
nor U19612 (N_19612,N_14720,N_16652);
or U19613 (N_19613,N_14939,N_14624);
or U19614 (N_19614,N_17458,N_17387);
nor U19615 (N_19615,N_14233,N_15024);
xnor U19616 (N_19616,N_17799,N_14900);
or U19617 (N_19617,N_14676,N_14443);
xnor U19618 (N_19618,N_16048,N_12089);
nor U19619 (N_19619,N_17240,N_17635);
and U19620 (N_19620,N_16390,N_16346);
nor U19621 (N_19621,N_12461,N_13078);
xor U19622 (N_19622,N_15544,N_16381);
nor U19623 (N_19623,N_17469,N_17802);
xor U19624 (N_19624,N_15051,N_16924);
nand U19625 (N_19625,N_14241,N_14383);
nor U19626 (N_19626,N_14508,N_17997);
nand U19627 (N_19627,N_17096,N_15625);
nand U19628 (N_19628,N_13276,N_15772);
and U19629 (N_19629,N_13639,N_17001);
nor U19630 (N_19630,N_14735,N_14408);
xor U19631 (N_19631,N_15513,N_17886);
or U19632 (N_19632,N_15638,N_16639);
xnor U19633 (N_19633,N_17764,N_16022);
and U19634 (N_19634,N_17944,N_17002);
or U19635 (N_19635,N_12719,N_12008);
nor U19636 (N_19636,N_17918,N_16772);
or U19637 (N_19637,N_15188,N_13277);
or U19638 (N_19638,N_14974,N_16902);
nor U19639 (N_19639,N_12210,N_15582);
nor U19640 (N_19640,N_16410,N_14105);
xor U19641 (N_19641,N_12416,N_14301);
and U19642 (N_19642,N_13068,N_16878);
and U19643 (N_19643,N_13204,N_17664);
or U19644 (N_19644,N_12497,N_12364);
and U19645 (N_19645,N_13809,N_17506);
nand U19646 (N_19646,N_16349,N_12038);
nor U19647 (N_19647,N_17864,N_13017);
or U19648 (N_19648,N_14016,N_12587);
nor U19649 (N_19649,N_12109,N_14800);
or U19650 (N_19650,N_16201,N_14828);
xor U19651 (N_19651,N_16515,N_12305);
nor U19652 (N_19652,N_13138,N_17844);
nand U19653 (N_19653,N_14989,N_15446);
nand U19654 (N_19654,N_13673,N_15745);
xnor U19655 (N_19655,N_15464,N_12408);
nor U19656 (N_19656,N_16484,N_13656);
xnor U19657 (N_19657,N_13875,N_15827);
xnor U19658 (N_19658,N_16238,N_15043);
and U19659 (N_19659,N_13294,N_16182);
and U19660 (N_19660,N_16315,N_15776);
nor U19661 (N_19661,N_13961,N_17738);
nor U19662 (N_19662,N_16524,N_17980);
and U19663 (N_19663,N_17771,N_16255);
and U19664 (N_19664,N_13503,N_15180);
and U19665 (N_19665,N_14503,N_15545);
and U19666 (N_19666,N_16430,N_15356);
or U19667 (N_19667,N_12607,N_14992);
nor U19668 (N_19668,N_15926,N_17898);
nand U19669 (N_19669,N_14136,N_13936);
xor U19670 (N_19670,N_16731,N_12241);
and U19671 (N_19671,N_15750,N_15768);
nor U19672 (N_19672,N_17462,N_16680);
and U19673 (N_19673,N_16395,N_16329);
xnor U19674 (N_19674,N_14523,N_12411);
and U19675 (N_19675,N_13492,N_14009);
xnor U19676 (N_19676,N_17321,N_13984);
nor U19677 (N_19677,N_17694,N_14060);
or U19678 (N_19678,N_15413,N_15050);
nand U19679 (N_19679,N_15784,N_16063);
and U19680 (N_19680,N_14870,N_15353);
nor U19681 (N_19681,N_15011,N_13016);
nor U19682 (N_19682,N_12076,N_16971);
nor U19683 (N_19683,N_12626,N_17789);
and U19684 (N_19684,N_16436,N_16845);
xor U19685 (N_19685,N_17376,N_17128);
nor U19686 (N_19686,N_16758,N_13942);
nor U19687 (N_19687,N_12646,N_17094);
nand U19688 (N_19688,N_14613,N_16686);
nor U19689 (N_19689,N_13207,N_13101);
and U19690 (N_19690,N_16223,N_15189);
nor U19691 (N_19691,N_13666,N_14209);
and U19692 (N_19692,N_15912,N_15556);
nand U19693 (N_19693,N_17534,N_13991);
nand U19694 (N_19694,N_17910,N_16793);
nor U19695 (N_19695,N_17901,N_16338);
and U19696 (N_19696,N_16374,N_17509);
nand U19697 (N_19697,N_15033,N_16307);
nand U19698 (N_19698,N_13731,N_15515);
nor U19699 (N_19699,N_12979,N_13669);
nand U19700 (N_19700,N_12593,N_17885);
nor U19701 (N_19701,N_12117,N_17233);
and U19702 (N_19702,N_13619,N_13542);
xnor U19703 (N_19703,N_13637,N_13305);
nand U19704 (N_19704,N_14920,N_15598);
xnor U19705 (N_19705,N_17403,N_13110);
nand U19706 (N_19706,N_15444,N_14289);
xnor U19707 (N_19707,N_13451,N_12444);
nor U19708 (N_19708,N_14020,N_17873);
and U19709 (N_19709,N_16953,N_17936);
nand U19710 (N_19710,N_15349,N_17029);
xor U19711 (N_19711,N_16367,N_14359);
nor U19712 (N_19712,N_14375,N_13090);
xnor U19713 (N_19713,N_16854,N_15153);
and U19714 (N_19714,N_16580,N_16950);
xor U19715 (N_19715,N_12612,N_14690);
or U19716 (N_19716,N_16462,N_14512);
or U19717 (N_19717,N_13618,N_13572);
or U19718 (N_19718,N_13513,N_13564);
xor U19719 (N_19719,N_14494,N_14777);
nand U19720 (N_19720,N_15300,N_14222);
or U19721 (N_19721,N_13852,N_12538);
nor U19722 (N_19722,N_14744,N_15652);
nor U19723 (N_19723,N_15004,N_14203);
and U19724 (N_19724,N_13616,N_13282);
or U19725 (N_19725,N_12344,N_13885);
and U19726 (N_19726,N_17642,N_16008);
nor U19727 (N_19727,N_17083,N_16669);
and U19728 (N_19728,N_12054,N_12690);
xnor U19729 (N_19729,N_13603,N_14814);
nor U19730 (N_19730,N_12030,N_14025);
or U19731 (N_19731,N_14714,N_14908);
nor U19732 (N_19732,N_12006,N_16473);
and U19733 (N_19733,N_13057,N_15237);
or U19734 (N_19734,N_12306,N_14146);
nor U19735 (N_19735,N_13528,N_16224);
nand U19736 (N_19736,N_16172,N_15895);
and U19737 (N_19737,N_13887,N_17995);
and U19738 (N_19738,N_17334,N_12024);
nor U19739 (N_19739,N_14761,N_12889);
nor U19740 (N_19740,N_14336,N_17769);
nand U19741 (N_19741,N_13163,N_16502);
nand U19742 (N_19742,N_13597,N_14491);
nor U19743 (N_19743,N_14955,N_16186);
or U19744 (N_19744,N_17745,N_16751);
nand U19745 (N_19745,N_13903,N_17985);
or U19746 (N_19746,N_17007,N_12342);
or U19747 (N_19747,N_14292,N_12869);
xnor U19748 (N_19748,N_17215,N_14927);
nand U19749 (N_19749,N_15034,N_15381);
or U19750 (N_19750,N_16763,N_13460);
or U19751 (N_19751,N_16427,N_15602);
nand U19752 (N_19752,N_12196,N_17704);
xor U19753 (N_19753,N_16248,N_15909);
or U19754 (N_19754,N_12356,N_17632);
or U19755 (N_19755,N_14294,N_14572);
nor U19756 (N_19756,N_13372,N_17818);
or U19757 (N_19757,N_13296,N_13194);
and U19758 (N_19758,N_16899,N_16747);
xor U19759 (N_19759,N_16717,N_14901);
xor U19760 (N_19760,N_16765,N_16065);
nor U19761 (N_19761,N_13329,N_13551);
nor U19762 (N_19762,N_12055,N_12316);
and U19763 (N_19763,N_16759,N_17774);
or U19764 (N_19764,N_16930,N_17118);
xor U19765 (N_19765,N_13346,N_12053);
and U19766 (N_19766,N_13520,N_17792);
nor U19767 (N_19767,N_17928,N_14225);
and U19768 (N_19768,N_13879,N_14990);
or U19769 (N_19769,N_13155,N_15859);
xnor U19770 (N_19770,N_12423,N_13515);
or U19771 (N_19771,N_16107,N_15596);
and U19772 (N_19772,N_12834,N_14650);
or U19773 (N_19773,N_13558,N_15363);
and U19774 (N_19774,N_16324,N_16818);
and U19775 (N_19775,N_17578,N_12815);
nor U19776 (N_19776,N_16853,N_13622);
nor U19777 (N_19777,N_17402,N_14476);
nand U19778 (N_19778,N_17749,N_16939);
nor U19779 (N_19779,N_13818,N_14866);
xor U19780 (N_19780,N_13278,N_14492);
or U19781 (N_19781,N_16612,N_13779);
xnor U19782 (N_19782,N_12841,N_15360);
and U19783 (N_19783,N_14216,N_16085);
nand U19784 (N_19784,N_17485,N_16621);
nor U19785 (N_19785,N_12541,N_16365);
and U19786 (N_19786,N_13716,N_17761);
or U19787 (N_19787,N_13147,N_12907);
nor U19788 (N_19788,N_12409,N_16811);
and U19789 (N_19789,N_13717,N_16729);
nor U19790 (N_19790,N_16858,N_13537);
nand U19791 (N_19791,N_12886,N_16247);
xnor U19792 (N_19792,N_13452,N_16435);
nand U19793 (N_19793,N_15993,N_15966);
or U19794 (N_19794,N_15738,N_13121);
nor U19795 (N_19795,N_13167,N_14001);
or U19796 (N_19796,N_17693,N_13136);
and U19797 (N_19797,N_17794,N_13038);
nand U19798 (N_19798,N_15855,N_15015);
and U19799 (N_19799,N_12855,N_14499);
and U19800 (N_19800,N_15486,N_13613);
xnor U19801 (N_19801,N_13298,N_15327);
nand U19802 (N_19802,N_17102,N_16139);
or U19803 (N_19803,N_14741,N_17531);
nor U19804 (N_19804,N_17177,N_17229);
nand U19805 (N_19805,N_16051,N_15291);
and U19806 (N_19806,N_13307,N_17668);
and U19807 (N_19807,N_17973,N_17634);
and U19808 (N_19808,N_13099,N_14808);
xor U19809 (N_19809,N_17372,N_12287);
nor U19810 (N_19810,N_12922,N_13655);
and U19811 (N_19811,N_16010,N_16808);
or U19812 (N_19812,N_15299,N_17188);
nor U19813 (N_19813,N_14806,N_14428);
and U19814 (N_19814,N_16284,N_15222);
nand U19815 (N_19815,N_12667,N_12074);
nor U19816 (N_19816,N_13328,N_15655);
nand U19817 (N_19817,N_13816,N_16965);
nor U19818 (N_19818,N_16281,N_16377);
and U19819 (N_19819,N_12312,N_17131);
xnor U19820 (N_19820,N_16625,N_17546);
nor U19821 (N_19821,N_13215,N_13334);
nand U19822 (N_19822,N_13760,N_12262);
nand U19823 (N_19823,N_13632,N_12073);
xor U19824 (N_19824,N_12575,N_15292);
or U19825 (N_19825,N_16624,N_17478);
xor U19826 (N_19826,N_15812,N_15488);
nor U19827 (N_19827,N_14753,N_12983);
nor U19828 (N_19828,N_17142,N_14346);
xor U19829 (N_19829,N_16205,N_17837);
or U19830 (N_19830,N_17292,N_17518);
and U19831 (N_19831,N_12094,N_15616);
and U19832 (N_19832,N_14675,N_17237);
xnor U19833 (N_19833,N_14275,N_15578);
and U19834 (N_19834,N_13259,N_13832);
xor U19835 (N_19835,N_13807,N_13032);
or U19836 (N_19836,N_17360,N_15116);
nand U19837 (N_19837,N_13012,N_15265);
nand U19838 (N_19838,N_12026,N_12040);
or U19839 (N_19839,N_15742,N_16136);
or U19840 (N_19840,N_13056,N_16335);
and U19841 (N_19841,N_16138,N_17281);
and U19842 (N_19842,N_13966,N_13546);
or U19843 (N_19843,N_14742,N_16824);
nand U19844 (N_19844,N_15727,N_16780);
xor U19845 (N_19845,N_15284,N_15217);
nand U19846 (N_19846,N_12297,N_14431);
nand U19847 (N_19847,N_17163,N_17696);
nand U19848 (N_19848,N_14589,N_13556);
xnor U19849 (N_19849,N_12840,N_17835);
and U19850 (N_19850,N_13116,N_14385);
or U19851 (N_19851,N_14519,N_17017);
nand U19852 (N_19852,N_17498,N_14477);
nand U19853 (N_19853,N_13773,N_14252);
nand U19854 (N_19854,N_13791,N_15075);
nand U19855 (N_19855,N_14166,N_17202);
and U19856 (N_19856,N_12938,N_16543);
nand U19857 (N_19857,N_15551,N_17377);
nand U19858 (N_19858,N_12022,N_16383);
or U19859 (N_19859,N_13830,N_13670);
nand U19860 (N_19860,N_15996,N_12161);
nand U19861 (N_19861,N_15816,N_16700);
and U19862 (N_19862,N_16825,N_13336);
and U19863 (N_19863,N_17113,N_12787);
xnor U19864 (N_19864,N_13668,N_15176);
xor U19865 (N_19865,N_17081,N_16970);
and U19866 (N_19866,N_14059,N_14377);
nor U19867 (N_19867,N_17579,N_13614);
nor U19868 (N_19868,N_15923,N_12603);
xor U19869 (N_19869,N_12375,N_13366);
and U19870 (N_19870,N_16591,N_12796);
xnor U19871 (N_19871,N_15671,N_16640);
nand U19872 (N_19872,N_15461,N_16385);
nor U19873 (N_19873,N_12873,N_15589);
and U19874 (N_19874,N_16787,N_13842);
and U19875 (N_19875,N_13043,N_15927);
or U19876 (N_19876,N_17569,N_16919);
and U19877 (N_19877,N_12268,N_14855);
xor U19878 (N_19878,N_12615,N_16873);
nand U19879 (N_19879,N_16835,N_15163);
xnor U19880 (N_19880,N_13878,N_14647);
nor U19881 (N_19881,N_13197,N_12565);
nand U19882 (N_19882,N_13129,N_13811);
nand U19883 (N_19883,N_17259,N_14422);
and U19884 (N_19884,N_17994,N_16975);
nor U19885 (N_19885,N_17961,N_17133);
or U19886 (N_19886,N_14952,N_16979);
nand U19887 (N_19887,N_16016,N_16282);
xnor U19888 (N_19888,N_13584,N_12539);
and U19889 (N_19889,N_13874,N_12765);
and U19890 (N_19890,N_15592,N_13234);
and U19891 (N_19891,N_15000,N_16094);
and U19892 (N_19892,N_12313,N_14553);
nor U19893 (N_19893,N_14630,N_17679);
xor U19894 (N_19894,N_12232,N_14604);
or U19895 (N_19895,N_14981,N_12438);
nor U19896 (N_19896,N_16568,N_17619);
nor U19897 (N_19897,N_13718,N_15373);
xor U19898 (N_19898,N_13439,N_16156);
xor U19899 (N_19899,N_16730,N_17993);
nand U19900 (N_19900,N_14029,N_15162);
and U19901 (N_19901,N_14871,N_15849);
nor U19902 (N_19902,N_14606,N_13526);
nand U19903 (N_19903,N_13553,N_16809);
nand U19904 (N_19904,N_17016,N_17609);
or U19905 (N_19905,N_15425,N_14906);
nand U19906 (N_19906,N_16738,N_16617);
or U19907 (N_19907,N_12070,N_15098);
nor U19908 (N_19908,N_15964,N_12489);
or U19909 (N_19909,N_16897,N_12288);
xor U19910 (N_19910,N_13626,N_12824);
and U19911 (N_19911,N_15499,N_17298);
or U19912 (N_19912,N_15569,N_14322);
xnor U19913 (N_19913,N_12793,N_12336);
nor U19914 (N_19914,N_17748,N_12516);
nand U19915 (N_19915,N_15500,N_14267);
and U19916 (N_19916,N_15434,N_12283);
xor U19917 (N_19917,N_17790,N_12066);
or U19918 (N_19918,N_13598,N_16487);
and U19919 (N_19919,N_14360,N_15678);
or U19920 (N_19920,N_17340,N_13638);
nor U19921 (N_19921,N_17013,N_16657);
or U19922 (N_19922,N_16921,N_12271);
or U19923 (N_19923,N_17572,N_17700);
nand U19924 (N_19924,N_12560,N_17105);
nor U19925 (N_19925,N_15663,N_14088);
xnor U19926 (N_19926,N_14802,N_16177);
nor U19927 (N_19927,N_14659,N_13819);
and U19928 (N_19928,N_14715,N_17805);
nor U19929 (N_19929,N_13694,N_13845);
nor U19930 (N_19930,N_14201,N_15591);
xnor U19931 (N_19931,N_16140,N_12069);
or U19932 (N_19932,N_14559,N_15642);
or U19933 (N_19933,N_16856,N_16615);
and U19934 (N_19934,N_16132,N_15049);
and U19935 (N_19935,N_13877,N_13498);
or U19936 (N_19936,N_17879,N_15573);
and U19937 (N_19937,N_15873,N_12097);
nand U19938 (N_19938,N_14086,N_15248);
nor U19939 (N_19939,N_15389,N_15297);
nor U19940 (N_19940,N_12392,N_16373);
xnor U19941 (N_19941,N_16911,N_16616);
xor U19942 (N_19942,N_12601,N_17934);
nand U19943 (N_19943,N_12946,N_14560);
nand U19944 (N_19944,N_14853,N_16525);
nor U19945 (N_19945,N_15479,N_15268);
and U19946 (N_19946,N_13444,N_17779);
nand U19947 (N_19947,N_14912,N_13411);
nor U19948 (N_19948,N_12806,N_12387);
xor U19949 (N_19949,N_12203,N_12804);
nor U19950 (N_19950,N_17390,N_12674);
nand U19951 (N_19951,N_14054,N_16442);
nor U19952 (N_19952,N_17231,N_14840);
nor U19953 (N_19953,N_12236,N_14578);
or U19954 (N_19954,N_13040,N_17689);
and U19955 (N_19955,N_16071,N_17900);
nand U19956 (N_19956,N_17557,N_14343);
xnor U19957 (N_19957,N_13582,N_15871);
xor U19958 (N_19958,N_13549,N_13350);
nor U19959 (N_19959,N_15632,N_17491);
nor U19960 (N_19960,N_12445,N_16446);
or U19961 (N_19961,N_16142,N_16670);
or U19962 (N_19962,N_14023,N_17786);
or U19963 (N_19963,N_16589,N_14809);
nor U19964 (N_19964,N_12536,N_15225);
xnor U19965 (N_19965,N_14843,N_13029);
or U19966 (N_19966,N_13931,N_14635);
xor U19967 (N_19967,N_12365,N_13654);
nor U19968 (N_19968,N_17651,N_14163);
and U19969 (N_19969,N_14548,N_15842);
nand U19970 (N_19970,N_13924,N_13583);
xor U19971 (N_19971,N_15160,N_15972);
and U19972 (N_19972,N_17646,N_15150);
nand U19973 (N_19973,N_12582,N_12617);
xor U19974 (N_19974,N_16178,N_14530);
nor U19975 (N_19975,N_15808,N_16668);
xnor U19976 (N_19976,N_12431,N_14467);
and U19977 (N_19977,N_17225,N_16870);
or U19978 (N_19978,N_12420,N_15113);
xor U19979 (N_19979,N_15289,N_15185);
or U19980 (N_19980,N_17806,N_14547);
or U19981 (N_19981,N_17722,N_13675);
or U19982 (N_19982,N_17787,N_12623);
nand U19983 (N_19983,N_14644,N_12600);
xnor U19984 (N_19984,N_13408,N_17015);
xor U19985 (N_19985,N_15660,N_14101);
nand U19986 (N_19986,N_13065,N_12325);
xnor U19987 (N_19987,N_13764,N_13514);
nand U19988 (N_19988,N_13051,N_15177);
or U19989 (N_19989,N_15460,N_16124);
xor U19990 (N_19990,N_13436,N_13383);
nand U19991 (N_19991,N_17767,N_13449);
and U19992 (N_19992,N_16252,N_16353);
nand U19993 (N_19993,N_15766,N_17654);
xor U19994 (N_19994,N_13025,N_13481);
nand U19995 (N_19995,N_15337,N_13663);
xor U19996 (N_19996,N_12346,N_12187);
nand U19997 (N_19997,N_14880,N_12678);
nand U19998 (N_19998,N_12138,N_16269);
nand U19999 (N_19999,N_12453,N_13894);
nand U20000 (N_20000,N_14832,N_14333);
and U20001 (N_20001,N_15260,N_12715);
and U20002 (N_20002,N_12581,N_12696);
nand U20003 (N_20003,N_17945,N_13287);
nand U20004 (N_20004,N_13974,N_14552);
nor U20005 (N_20005,N_14739,N_12712);
or U20006 (N_20006,N_14643,N_14331);
nand U20007 (N_20007,N_14786,N_15174);
or U20008 (N_20008,N_12928,N_12558);
nor U20009 (N_20009,N_16345,N_15844);
nor U20010 (N_20010,N_13522,N_16714);
nand U20011 (N_20011,N_15287,N_12462);
or U20012 (N_20012,N_16121,N_12914);
xnor U20013 (N_20013,N_12351,N_14034);
or U20014 (N_20014,N_15554,N_14842);
nand U20015 (N_20015,N_16161,N_12991);
xnor U20016 (N_20016,N_12385,N_12996);
and U20017 (N_20017,N_12933,N_12891);
or U20018 (N_20018,N_14737,N_16748);
and U20019 (N_20019,N_13624,N_15973);
and U20020 (N_20020,N_15770,N_12384);
nor U20021 (N_20021,N_16035,N_15702);
or U20022 (N_20022,N_14677,N_12879);
or U20023 (N_20023,N_12449,N_16321);
or U20024 (N_20024,N_15393,N_15002);
nor U20025 (N_20025,N_14014,N_13796);
nand U20026 (N_20026,N_15197,N_16386);
nand U20027 (N_20027,N_16508,N_13108);
and U20028 (N_20028,N_12988,N_15061);
xor U20029 (N_20029,N_14339,N_14021);
and U20030 (N_20030,N_15166,N_12639);
xor U20031 (N_20031,N_17605,N_15442);
xor U20032 (N_20032,N_13021,N_14239);
xor U20033 (N_20033,N_13221,N_15288);
or U20034 (N_20034,N_12974,N_16013);
and U20035 (N_20035,N_14411,N_13927);
xor U20036 (N_20036,N_14066,N_17003);
nor U20037 (N_20037,N_13388,N_14286);
xor U20038 (N_20038,N_12689,N_15618);
and U20039 (N_20039,N_14310,N_17465);
and U20040 (N_20040,N_13395,N_12442);
and U20041 (N_20041,N_13344,N_14839);
nand U20042 (N_20042,N_17986,N_17966);
and U20043 (N_20043,N_12771,N_14620);
nor U20044 (N_20044,N_17788,N_16069);
nor U20045 (N_20045,N_17503,N_14457);
nand U20046 (N_20046,N_16402,N_14018);
xor U20047 (N_20047,N_14542,N_12954);
and U20048 (N_20048,N_13096,N_15853);
nand U20049 (N_20049,N_14710,N_16850);
xnor U20050 (N_20050,N_15395,N_17631);
xnor U20051 (N_20051,N_12482,N_14012);
xnor U20052 (N_20052,N_13606,N_17070);
or U20053 (N_20053,N_13712,N_12106);
nand U20054 (N_20054,N_17467,N_13628);
nand U20055 (N_20055,N_15968,N_14197);
or U20056 (N_20056,N_14276,N_16199);
xnor U20057 (N_20057,N_17448,N_15567);
nor U20058 (N_20058,N_12713,N_12432);
nand U20059 (N_20059,N_12640,N_14799);
xnor U20060 (N_20060,N_14401,N_12682);
and U20061 (N_20061,N_15525,N_17502);
nand U20062 (N_20062,N_14113,N_12152);
or U20063 (N_20063,N_17673,N_16821);
nand U20064 (N_20064,N_17699,N_17525);
xor U20065 (N_20065,N_16559,N_15379);
or U20066 (N_20066,N_16922,N_14394);
nor U20067 (N_20067,N_15621,N_16523);
nor U20068 (N_20068,N_16303,N_12642);
nor U20069 (N_20069,N_14157,N_16557);
nor U20070 (N_20070,N_17150,N_15783);
nand U20071 (N_20071,N_17241,N_16739);
and U20072 (N_20072,N_13932,N_13770);
xor U20073 (N_20073,N_12832,N_15902);
nand U20074 (N_20074,N_12301,N_14313);
nand U20075 (N_20075,N_13610,N_14540);
or U20076 (N_20076,N_14838,N_13899);
or U20077 (N_20077,N_14538,N_15306);
or U20078 (N_20078,N_15184,N_16021);
or U20079 (N_20079,N_17705,N_15329);
xor U20080 (N_20080,N_12142,N_17446);
or U20081 (N_20081,N_14039,N_14569);
nand U20082 (N_20082,N_13533,N_14531);
nor U20083 (N_20083,N_12063,N_13125);
xnor U20084 (N_20084,N_14856,N_15495);
and U20085 (N_20085,N_14883,N_16828);
or U20086 (N_20086,N_17808,N_14713);
and U20087 (N_20087,N_14419,N_13707);
and U20088 (N_20088,N_16957,N_13858);
or U20089 (N_20089,N_16044,N_15118);
nand U20090 (N_20090,N_14033,N_14554);
nor U20091 (N_20091,N_13241,N_15635);
xor U20092 (N_20092,N_12168,N_15350);
xor U20093 (N_20093,N_15213,N_17278);
nand U20094 (N_20094,N_13143,N_12116);
xor U20095 (N_20095,N_17304,N_16581);
nand U20096 (N_20096,N_12103,N_13126);
or U20097 (N_20097,N_17170,N_14126);
or U20098 (N_20098,N_15861,N_14489);
or U20099 (N_20099,N_16741,N_14726);
nand U20100 (N_20100,N_12120,N_13941);
and U20101 (N_20101,N_17273,N_15931);
nor U20102 (N_20102,N_14973,N_14970);
nor U20103 (N_20103,N_15233,N_12677);
nand U20104 (N_20104,N_13802,N_14098);
nor U20105 (N_20105,N_13674,N_13839);
xor U20106 (N_20106,N_15452,N_17551);
nand U20107 (N_20107,N_15961,N_13483);
xnor U20108 (N_20108,N_12493,N_17528);
and U20109 (N_20109,N_13922,N_14913);
nand U20110 (N_20110,N_14873,N_14748);
nand U20111 (N_20111,N_14420,N_13938);
xor U20112 (N_20112,N_14348,N_17191);
xnor U20113 (N_20113,N_14055,N_16864);
and U20114 (N_20114,N_15100,N_12422);
and U20115 (N_20115,N_15105,N_13028);
or U20116 (N_20116,N_15533,N_16169);
or U20117 (N_20117,N_15810,N_13871);
nand U20118 (N_20118,N_12088,N_16183);
nor U20119 (N_20119,N_14985,N_17505);
nor U20120 (N_20120,N_15918,N_12487);
or U20121 (N_20121,N_16229,N_17629);
nand U20122 (N_20122,N_16644,N_14129);
nand U20123 (N_20123,N_13752,N_14673);
nand U20124 (N_20124,N_17729,N_16871);
xnor U20125 (N_20125,N_16838,N_17497);
and U20126 (N_20126,N_16797,N_12157);
nand U20127 (N_20127,N_12523,N_16832);
nand U20128 (N_20128,N_16764,N_12175);
or U20129 (N_20129,N_17438,N_13173);
nand U20130 (N_20130,N_17775,N_13286);
and U20131 (N_20131,N_14274,N_12358);
xnor U20132 (N_20132,N_15427,N_12345);
nand U20133 (N_20133,N_16781,N_12159);
and U20134 (N_20134,N_13140,N_13856);
xor U20135 (N_20135,N_14977,N_15117);
or U20136 (N_20136,N_15664,N_12521);
or U20137 (N_20137,N_14116,N_17530);
xnor U20138 (N_20138,N_13218,N_15199);
nand U20139 (N_20139,N_12045,N_16380);
nor U20140 (N_20140,N_17203,N_12629);
nor U20141 (N_20141,N_12355,N_17027);
nand U20142 (N_20142,N_14111,N_16925);
or U20143 (N_20143,N_16454,N_15003);
or U20144 (N_20144,N_17296,N_17884);
xnor U20145 (N_20145,N_16917,N_13921);
nand U20146 (N_20146,N_17780,N_13866);
nor U20147 (N_20147,N_16244,N_14517);
and U20148 (N_20148,N_12446,N_13680);
or U20149 (N_20149,N_12637,N_12163);
and U20150 (N_20150,N_15077,N_16661);
xnor U20151 (N_20151,N_15507,N_15092);
or U20152 (N_20152,N_15506,N_16633);
xnor U20153 (N_20153,N_14218,N_16097);
nor U20154 (N_20154,N_14961,N_16159);
and U20155 (N_20155,N_12947,N_17258);
or U20156 (N_20156,N_16028,N_14357);
xnor U20157 (N_20157,N_15734,N_16989);
nand U20158 (N_20158,N_13426,N_15058);
and U20159 (N_20159,N_14953,N_15078);
or U20160 (N_20160,N_13235,N_16572);
nand U20161 (N_20161,N_14626,N_15151);
and U20162 (N_20162,N_16990,N_15017);
nor U20163 (N_20163,N_13248,N_15526);
or U20164 (N_20164,N_14063,N_16690);
nand U20165 (N_20165,N_14623,N_12244);
nor U20166 (N_20166,N_14964,N_12092);
xnor U20167 (N_20167,N_17396,N_13397);
nand U20168 (N_20168,N_17820,N_15096);
xor U20169 (N_20169,N_16341,N_12418);
and U20170 (N_20170,N_12611,N_17440);
nor U20171 (N_20171,N_13359,N_15448);
and U20172 (N_20172,N_14860,N_13659);
or U20173 (N_20173,N_16456,N_17827);
nand U20174 (N_20174,N_14247,N_16869);
nor U20175 (N_20175,N_14024,N_12749);
nand U20176 (N_20176,N_14073,N_13806);
and U20177 (N_20177,N_17661,N_13008);
nand U20178 (N_20178,N_16577,N_12280);
or U20179 (N_20179,N_16627,N_14258);
xnor U20180 (N_20180,N_12745,N_17514);
nor U20181 (N_20181,N_15988,N_16788);
or U20182 (N_20182,N_13950,N_14803);
and U20183 (N_20183,N_16962,N_14131);
or U20184 (N_20184,N_12966,N_12747);
xnor U20185 (N_20185,N_15331,N_13900);
nor U20186 (N_20186,N_13251,N_14810);
xor U20187 (N_20187,N_17639,N_13649);
and U20188 (N_20188,N_16302,N_13391);
or U20189 (N_20189,N_17547,N_12362);
or U20190 (N_20190,N_17988,N_13188);
or U20191 (N_20191,N_12366,N_12572);
nor U20192 (N_20192,N_17201,N_12883);
and U20193 (N_20193,N_15502,N_16276);
or U20194 (N_20194,N_15343,N_12958);
or U20195 (N_20195,N_12016,N_12564);
or U20196 (N_20196,N_17809,N_17335);
nand U20197 (N_20197,N_16419,N_15527);
and U20198 (N_20198,N_17659,N_15878);
nor U20199 (N_20199,N_15767,N_17311);
or U20200 (N_20200,N_13326,N_12884);
and U20201 (N_20201,N_13735,N_17189);
or U20202 (N_20202,N_15264,N_17034);
nor U20203 (N_20203,N_16032,N_17610);
nor U20204 (N_20204,N_15191,N_12319);
nor U20205 (N_20205,N_13687,N_15689);
xor U20206 (N_20206,N_17958,N_14795);
and U20207 (N_20207,N_16666,N_13193);
nand U20208 (N_20208,N_12755,N_14178);
or U20209 (N_20209,N_12475,N_12434);
or U20210 (N_20210,N_13996,N_17867);
nor U20211 (N_20211,N_12781,N_16826);
nor U20212 (N_20212,N_16805,N_17212);
nand U20213 (N_20213,N_16689,N_13552);
or U20214 (N_20214,N_17405,N_14287);
or U20215 (N_20215,N_14062,N_12644);
and U20216 (N_20216,N_14674,N_13512);
and U20217 (N_20217,N_17641,N_12604);
xnor U20218 (N_20218,N_12981,N_12653);
nor U20219 (N_20219,N_14030,N_13561);
or U20220 (N_20220,N_13438,N_12007);
nor U20221 (N_20221,N_14539,N_13679);
or U20222 (N_20222,N_12818,N_15140);
or U20223 (N_20223,N_17466,N_14640);
xor U20224 (N_20224,N_12729,N_13023);
and U20225 (N_20225,N_16836,N_15579);
nand U20226 (N_20226,N_17737,N_15599);
xnor U20227 (N_20227,N_15888,N_12672);
xnor U20228 (N_20228,N_12015,N_15529);
and U20229 (N_20229,N_15374,N_12079);
nand U20230 (N_20230,N_17323,N_13862);
or U20231 (N_20231,N_16350,N_15172);
xnor U20232 (N_20232,N_14370,N_13348);
nor U20233 (N_20233,N_14480,N_14986);
nor U20234 (N_20234,N_17536,N_17943);
and U20235 (N_20235,N_13250,N_17055);
nand U20236 (N_20236,N_14417,N_12929);
nor U20237 (N_20237,N_16167,N_15401);
and U20238 (N_20238,N_12467,N_15104);
xnor U20239 (N_20239,N_17513,N_13738);
or U20240 (N_20240,N_12934,N_12277);
and U20241 (N_20241,N_17545,N_14090);
xor U20242 (N_20242,N_14976,N_17859);
and U20243 (N_20243,N_12702,N_13034);
nand U20244 (N_20244,N_16190,N_16959);
xor U20245 (N_20245,N_13476,N_12143);
nor U20246 (N_20246,N_12134,N_17010);
nor U20247 (N_20247,N_17018,N_12766);
nand U20248 (N_20248,N_13053,N_17893);
xor U20249 (N_20249,N_15920,N_12563);
nor U20250 (N_20250,N_17254,N_15601);
and U20251 (N_20251,N_12903,N_16583);
and U20252 (N_20252,N_12201,N_17960);
nor U20253 (N_20253,N_12185,N_15692);
or U20254 (N_20254,N_15921,N_16145);
nand U20255 (N_20255,N_15963,N_12687);
and U20256 (N_20256,N_14487,N_16312);
or U20257 (N_20257,N_17743,N_14110);
xor U20258 (N_20258,N_16297,N_17194);
nor U20259 (N_20259,N_12616,N_16511);
xor U20260 (N_20260,N_17521,N_13566);
nor U20261 (N_20261,N_15308,N_15110);
nand U20262 (N_20262,N_15575,N_15227);
or U20263 (N_20263,N_12429,N_13437);
nand U20264 (N_20264,N_17931,N_17174);
xor U20265 (N_20265,N_17171,N_16718);
nor U20266 (N_20266,N_12778,N_15797);
xnor U20267 (N_20267,N_15843,N_14925);
nor U20268 (N_20268,N_15831,N_12249);
and U20269 (N_20269,N_14369,N_13239);
xnor U20270 (N_20270,N_16848,N_16429);
and U20271 (N_20271,N_14160,N_13876);
nor U20272 (N_20272,N_15870,N_16519);
or U20273 (N_20273,N_12807,N_12535);
or U20274 (N_20274,N_17849,N_13758);
nor U20275 (N_20275,N_12759,N_17684);
or U20276 (N_20276,N_12826,N_15313);
or U20277 (N_20277,N_16628,N_17541);
nor U20278 (N_20278,N_12942,N_15626);
and U20279 (N_20279,N_13139,N_14896);
and U20280 (N_20280,N_16034,N_13479);
and U20281 (N_20281,N_13472,N_12986);
xnor U20282 (N_20282,N_13708,N_14043);
xor U20283 (N_20283,N_16425,N_12968);
and U20284 (N_20284,N_16840,N_12579);
nand U20285 (N_20285,N_13240,N_12638);
nor U20286 (N_20286,N_16155,N_12334);
or U20287 (N_20287,N_15704,N_13117);
nand U20288 (N_20288,N_15410,N_13073);
and U20289 (N_20289,N_12009,N_17753);
or U20290 (N_20290,N_13393,N_17630);
xnor U20291 (N_20291,N_12005,N_12872);
nor U20292 (N_20292,N_14355,N_13358);
xor U20293 (N_20293,N_16384,N_17798);
nor U20294 (N_20294,N_17268,N_14134);
and U20295 (N_20295,N_15232,N_14653);
nand U20296 (N_20296,N_13676,N_16964);
or U20297 (N_20297,N_12357,N_14325);
or U20298 (N_20298,N_15030,N_12501);
and U20299 (N_20299,N_16813,N_14945);
nand U20300 (N_20300,N_12789,N_13697);
and U20301 (N_20301,N_13635,N_16516);
and U20302 (N_20302,N_15851,N_17633);
or U20303 (N_20303,N_14734,N_16127);
or U20304 (N_20304,N_15886,N_13798);
or U20305 (N_20305,N_17136,N_14236);
or U20306 (N_20306,N_12875,N_15850);
nand U20307 (N_20307,N_13319,N_12413);
nor U20308 (N_20308,N_17871,N_14562);
xor U20309 (N_20309,N_12035,N_13230);
xnor U20310 (N_20310,N_15223,N_15271);
nand U20311 (N_20311,N_17042,N_12253);
and U20312 (N_20312,N_17144,N_16865);
and U20313 (N_20313,N_17752,N_15462);
nand U20314 (N_20314,N_17020,N_14888);
nand U20315 (N_20315,N_13113,N_12794);
and U20316 (N_20316,N_17967,N_16471);
and U20317 (N_20317,N_17074,N_15647);
nor U20318 (N_20318,N_16466,N_15628);
xnor U20319 (N_20319,N_12202,N_15731);
nand U20320 (N_20320,N_13756,N_17736);
and U20321 (N_20321,N_13705,N_13019);
nand U20322 (N_20322,N_13392,N_13164);
xnor U20323 (N_20323,N_13754,N_16249);
nand U20324 (N_20324,N_16440,N_16388);
xor U20325 (N_20325,N_17711,N_17902);
nand U20326 (N_20326,N_12250,N_17279);
nor U20327 (N_20327,N_17719,N_13284);
xnor U20328 (N_20328,N_17824,N_13124);
and U20329 (N_20329,N_13357,N_17800);
nand U20330 (N_20330,N_13331,N_17168);
xnor U20331 (N_20331,N_17031,N_14940);
and U20332 (N_20332,N_12762,N_13457);
nand U20333 (N_20333,N_12898,N_15194);
nand U20334 (N_20334,N_12624,N_16997);
nor U20335 (N_20335,N_12777,N_15281);
xor U20336 (N_20336,N_17347,N_14993);
or U20337 (N_20337,N_13709,N_16909);
or U20338 (N_20338,N_17520,N_16151);
nor U20339 (N_20339,N_15540,N_15148);
xnor U20340 (N_20340,N_16225,N_14687);
or U20341 (N_20341,N_16912,N_13646);
nor U20342 (N_20342,N_17410,N_17755);
nand U20343 (N_20343,N_16671,N_14731);
xnor U20344 (N_20344,N_14266,N_13715);
nor U20345 (N_20345,N_16160,N_16701);
xor U20346 (N_20346,N_17408,N_15399);
and U20347 (N_20347,N_14791,N_17625);
xnor U20348 (N_20348,N_15471,N_12393);
or U20349 (N_20349,N_12658,N_12544);
nand U20350 (N_20350,N_13087,N_14095);
and U20351 (N_20351,N_14288,N_13570);
nand U20352 (N_20352,N_13706,N_16148);
nor U20353 (N_20353,N_16512,N_13314);
nor U20354 (N_20354,N_16347,N_15743);
nand U20355 (N_20355,N_17526,N_16478);
or U20356 (N_20356,N_17307,N_13349);
xor U20357 (N_20357,N_17499,N_12645);
nor U20358 (N_20358,N_16914,N_16888);
nand U20359 (N_20359,N_14616,N_15729);
and U20360 (N_20360,N_16480,N_14045);
xor U20361 (N_20361,N_15103,N_13594);
or U20362 (N_20362,N_14593,N_13061);
nor U20363 (N_20363,N_14899,N_16334);
and U20364 (N_20364,N_12972,N_14079);
nor U20365 (N_20365,N_16325,N_13859);
xor U20366 (N_20366,N_12286,N_17293);
xor U20367 (N_20367,N_16881,N_16299);
xnor U20368 (N_20368,N_12275,N_15956);
xor U20369 (N_20369,N_16977,N_12330);
nor U20370 (N_20370,N_16235,N_13569);
nor U20371 (N_20371,N_17915,N_14823);
or U20372 (N_20372,N_12072,N_12550);
xor U20373 (N_20373,N_13145,N_16413);
nand U20374 (N_20374,N_16135,N_17559);
or U20375 (N_20375,N_13360,N_14767);
nand U20376 (N_20376,N_16969,N_13225);
nor U20377 (N_20377,N_14561,N_17324);
nand U20378 (N_20378,N_17965,N_14251);
and U20379 (N_20379,N_12722,N_16814);
and U20380 (N_20380,N_12150,N_17424);
and U20381 (N_20381,N_12216,N_14423);
nor U20382 (N_20382,N_14693,N_17846);
nand U20383 (N_20383,N_15610,N_12791);
nand U20384 (N_20384,N_12899,N_16362);
xnor U20385 (N_20385,N_14661,N_17282);
xnor U20386 (N_20386,N_17598,N_12756);
nor U20387 (N_20387,N_17555,N_15245);
and U20388 (N_20388,N_12752,N_15665);
or U20389 (N_20389,N_14315,N_15167);
nor U20390 (N_20390,N_12019,N_17398);
xnor U20391 (N_20391,N_13094,N_15456);
or U20392 (N_20392,N_17603,N_13321);
xnor U20393 (N_20393,N_13494,N_15821);
or U20394 (N_20394,N_15780,N_15478);
xnor U20395 (N_20395,N_16676,N_17688);
or U20396 (N_20396,N_13074,N_16694);
or U20397 (N_20397,N_13134,N_12522);
xnor U20398 (N_20398,N_13431,N_15822);
xnor U20399 (N_20399,N_12227,N_16300);
nor U20400 (N_20400,N_17158,N_12059);
or U20401 (N_20401,N_14594,N_15998);
xnor U20402 (N_20402,N_15798,N_12255);
and U20403 (N_20403,N_16079,N_16672);
nor U20404 (N_20404,N_15441,N_14536);
and U20405 (N_20405,N_16323,N_13543);
or U20406 (N_20406,N_14248,N_12927);
nand U20407 (N_20407,N_12350,N_14229);
or U20408 (N_20408,N_15561,N_12190);
nor U20409 (N_20409,N_15700,N_15063);
xnor U20410 (N_20410,N_15771,N_14895);
and U20411 (N_20411,N_12002,N_15403);
nor U20412 (N_20412,N_16935,N_14400);
nor U20413 (N_20413,N_15346,N_15412);
xnor U20414 (N_20414,N_15336,N_17839);
nor U20415 (N_20415,N_17358,N_16673);
or U20416 (N_20416,N_14051,N_14996);
nand U20417 (N_20417,N_15713,N_15120);
and U20418 (N_20418,N_17833,N_16195);
xor U20419 (N_20419,N_17338,N_12400);
nor U20420 (N_20420,N_16314,N_14918);
nor U20421 (N_20421,N_13086,N_13338);
or U20422 (N_20422,N_12310,N_13112);
or U20423 (N_20423,N_14303,N_17941);
nand U20424 (N_20424,N_16189,N_14463);
nand U20425 (N_20425,N_16699,N_15037);
and U20426 (N_20426,N_17104,N_14907);
xor U20427 (N_20427,N_14397,N_17033);
or U20428 (N_20428,N_12398,N_14928);
and U20429 (N_20429,N_17389,N_16234);
and U20430 (N_20430,N_14395,N_13070);
or U20431 (N_20431,N_12329,N_15606);
nand U20432 (N_20432,N_12746,N_14365);
nand U20433 (N_20433,N_12814,N_12909);
xnor U20434 (N_20434,N_17758,N_15790);
nand U20435 (N_20435,N_15439,N_14421);
or U20436 (N_20436,N_13200,N_14682);
or U20437 (N_20437,N_17085,N_17005);
xnor U20438 (N_20438,N_12923,N_17899);
xnor U20439 (N_20439,N_15263,N_12533);
or U20440 (N_20440,N_12004,N_15402);
nand U20441 (N_20441,N_13401,N_16023);
or U20442 (N_20442,N_16260,N_12403);
or U20443 (N_20443,N_14371,N_13150);
nor U20444 (N_20444,N_15178,N_17715);
nor U20445 (N_20445,N_17044,N_13482);
xor U20446 (N_20446,N_17553,N_12149);
and U20447 (N_20447,N_15917,N_14921);
nor U20448 (N_20448,N_14532,N_15394);
nand U20449 (N_20449,N_15804,N_14127);
nor U20450 (N_20450,N_15082,N_14501);
nand U20451 (N_20451,N_12219,N_15744);
nand U20452 (N_20452,N_14344,N_13901);
or U20453 (N_20453,N_14821,N_14300);
xnor U20454 (N_20454,N_14941,N_16720);
and U20455 (N_20455,N_17676,N_13683);
and U20456 (N_20456,N_16564,N_16074);
and U20457 (N_20457,N_16036,N_14602);
xnor U20458 (N_20458,N_14573,N_16907);
xnor U20459 (N_20459,N_16277,N_14479);
nand U20460 (N_20460,N_14609,N_15424);
and U20461 (N_20461,N_15814,N_13390);
and U20462 (N_20462,N_17952,N_15894);
nand U20463 (N_20463,N_13265,N_16618);
nand U20464 (N_20464,N_12598,N_15922);
nand U20465 (N_20465,N_17030,N_12226);
and U20466 (N_20466,N_16391,N_13822);
nor U20467 (N_20467,N_16565,N_17356);
xnor U20468 (N_20468,N_13291,N_16635);
nor U20469 (N_20469,N_14923,N_14285);
xnor U20470 (N_20470,N_15041,N_15934);
and U20471 (N_20471,N_17274,N_14011);
xor U20472 (N_20472,N_16203,N_17687);
or U20473 (N_20473,N_15426,N_14137);
nand U20474 (N_20474,N_16768,N_15154);
nand U20475 (N_20475,N_12776,N_13448);
and U20476 (N_20476,N_12937,N_17184);
nor U20477 (N_20477,N_12011,N_12156);
nand U20478 (N_20478,N_15875,N_17600);
and U20479 (N_20479,N_16757,N_12532);
and U20480 (N_20480,N_13024,N_16158);
or U20481 (N_20481,N_15725,N_16414);
nor U20482 (N_20482,N_14117,N_16777);
nor U20483 (N_20483,N_16872,N_14304);
nor U20484 (N_20484,N_14707,N_17929);
and U20485 (N_20485,N_16834,N_12836);
xor U20486 (N_20486,N_17075,N_16528);
nor U20487 (N_20487,N_15634,N_15064);
or U20488 (N_20488,N_13362,N_17310);
nor U20489 (N_20489,N_17658,N_12780);
and U20490 (N_20490,N_14340,N_15535);
nor U20491 (N_20491,N_12017,N_17401);
nor U20492 (N_20492,N_17183,N_16082);
nand U20493 (N_20493,N_14482,N_16995);
or U20494 (N_20494,N_12589,N_16360);
xor U20495 (N_20495,N_15496,N_15454);
nor U20496 (N_20496,N_16340,N_16704);
nor U20497 (N_20497,N_15869,N_17352);
or U20498 (N_20498,N_12524,N_13417);
and U20499 (N_20499,N_13308,N_15856);
nor U20500 (N_20500,N_15737,N_17236);
and U20501 (N_20501,N_12307,N_12870);
xor U20502 (N_20502,N_15670,N_12514);
or U20503 (N_20503,N_14132,N_14078);
xor U20504 (N_20504,N_13788,N_17166);
nand U20505 (N_20505,N_12483,N_14265);
nor U20506 (N_20506,N_12701,N_12447);
nand U20507 (N_20507,N_13030,N_15358);
or U20508 (N_20508,N_17417,N_13249);
xnor U20509 (N_20509,N_13538,N_14164);
nor U20510 (N_20510,N_13130,N_16916);
or U20511 (N_20511,N_16503,N_14184);
nor U20512 (N_20512,N_13295,N_14250);
nand U20513 (N_20513,N_13828,N_15815);
or U20514 (N_20514,N_14130,N_16963);
and U20515 (N_20515,N_16308,N_13132);
nor U20516 (N_20516,N_14733,N_16846);
nor U20517 (N_20517,N_14109,N_12359);
nor U20518 (N_20518,N_15773,N_14567);
nand U20519 (N_20519,N_16075,N_17583);
or U20520 (N_20520,N_15558,N_12279);
or U20521 (N_20521,N_16563,N_14637);
and U20522 (N_20522,N_13075,N_16973);
and U20523 (N_20523,N_15229,N_15811);
nand U20524 (N_20524,N_12192,N_12670);
nand U20525 (N_20525,N_17441,N_15370);
nor U20526 (N_20526,N_14453,N_15782);
or U20527 (N_20527,N_12584,N_13404);
nand U20528 (N_20528,N_14937,N_17621);
and U20529 (N_20529,N_16265,N_12827);
nand U20530 (N_20530,N_16055,N_13502);
and U20531 (N_20531,N_12382,N_12328);
or U20532 (N_20532,N_17207,N_12234);
and U20533 (N_20533,N_16847,N_13578);
and U20534 (N_20534,N_15095,N_13946);
nand U20535 (N_20535,N_13719,N_17747);
nor U20536 (N_20536,N_17139,N_15045);
xnor U20537 (N_20537,N_17816,N_12774);
or U20538 (N_20538,N_16954,N_17913);
nor U20539 (N_20539,N_17246,N_12214);
and U20540 (N_20540,N_14381,N_16080);
xnor U20541 (N_20541,N_15032,N_14353);
nor U20542 (N_20542,N_12104,N_14751);
nor U20543 (N_20543,N_12950,N_17735);
xor U20544 (N_20544,N_15231,N_12767);
nor U20545 (N_20545,N_12885,N_15736);
nor U20546 (N_20546,N_12160,N_17190);
nand U20547 (N_20547,N_16619,N_16243);
xnor U20548 (N_20548,N_15445,N_12183);
and U20549 (N_20549,N_14628,N_13387);
and U20550 (N_20550,N_12311,N_16767);
nand U20551 (N_20551,N_12224,N_15991);
nand U20552 (N_20552,N_15251,N_12322);
xor U20553 (N_20553,N_15181,N_13154);
nor U20554 (N_20554,N_17068,N_14816);
xor U20555 (N_20555,N_13737,N_12739);
nor U20556 (N_20556,N_15283,N_13795);
xnor U20557 (N_20557,N_16147,N_15563);
and U20558 (N_20558,N_12511,N_12125);
or U20559 (N_20559,N_12726,N_13414);
nand U20560 (N_20560,N_17065,N_13531);
and U20561 (N_20561,N_12810,N_15696);
or U20562 (N_20562,N_17856,N_12757);
xnor U20563 (N_20563,N_13441,N_12813);
or U20564 (N_20564,N_17963,N_14576);
nor U20565 (N_20565,N_14329,N_13303);
or U20566 (N_20566,N_14268,N_17905);
nand U20567 (N_20567,N_13734,N_13648);
xnor U20568 (N_20568,N_13689,N_12978);
or U20569 (N_20569,N_17265,N_15564);
nor U20570 (N_20570,N_17894,N_15800);
nand U20571 (N_20571,N_12686,N_15785);
nor U20572 (N_20572,N_17674,N_16807);
nand U20573 (N_20573,N_13544,N_14112);
and U20574 (N_20574,N_12113,N_13854);
nor U20575 (N_20575,N_16327,N_17677);
and U20576 (N_20576,N_15809,N_14709);
nand U20577 (N_20577,N_17590,N_16967);
and U20578 (N_20578,N_13661,N_13333);
and U20579 (N_20579,N_16162,N_16432);
or U20580 (N_20580,N_17043,N_13219);
xor U20581 (N_20581,N_14796,N_12220);
nor U20582 (N_20582,N_15986,N_17256);
nor U20583 (N_20583,N_14074,N_14089);
nor U20584 (N_20584,N_16883,N_16181);
xnor U20585 (N_20585,N_16452,N_13547);
nor U20586 (N_20586,N_16946,N_17854);
nor U20587 (N_20587,N_12424,N_14478);
or U20588 (N_20588,N_12406,N_12876);
or U20589 (N_20589,N_12649,N_17810);
and U20590 (N_20590,N_16458,N_12661);
nor U20591 (N_20591,N_15646,N_17232);
and U20592 (N_20592,N_14485,N_17511);
xnor U20593 (N_20593,N_14119,N_17777);
xor U20594 (N_20594,N_15699,N_12095);
xor U20595 (N_20595,N_16306,N_12086);
nor U20596 (N_20596,N_14521,N_13881);
nand U20597 (N_20597,N_15978,N_17968);
and U20598 (N_20598,N_12940,N_14727);
nor U20599 (N_20599,N_17713,N_12555);
and U20600 (N_20600,N_15935,N_13910);
or U20601 (N_20601,N_15458,N_15334);
xor U20602 (N_20602,N_12182,N_15503);
nor U20603 (N_20603,N_17501,N_13381);
and U20604 (N_20604,N_12140,N_17089);
xor U20605 (N_20605,N_14008,N_16387);
nor U20606 (N_20606,N_14957,N_15155);
nor U20607 (N_20607,N_16401,N_15108);
nand U20608 (N_20608,N_13288,N_13908);
and U20609 (N_20609,N_15614,N_13283);
nor U20610 (N_20610,N_13861,N_16776);
or U20611 (N_20611,N_15493,N_12939);
or U20612 (N_20612,N_12228,N_15903);
xnor U20613 (N_20613,N_13849,N_13550);
nand U20614 (N_20614,N_12844,N_16271);
nor U20615 (N_20615,N_17683,N_12474);
nand U20616 (N_20616,N_15980,N_12126);
or U20617 (N_20617,N_13970,N_14984);
nand U20618 (N_20618,N_16099,N_17161);
xnor U20619 (N_20619,N_15905,N_17663);
and U20620 (N_20620,N_15838,N_16208);
or U20621 (N_20621,N_15498,N_12602);
nand U20622 (N_20622,N_14689,N_13650);
nor U20623 (N_20623,N_12000,N_13729);
xnor U20624 (N_20624,N_14283,N_12176);
xnor U20625 (N_20625,N_14980,N_14580);
nand U20626 (N_20626,N_16630,N_14765);
and U20627 (N_20627,N_16332,N_16096);
xor U20628 (N_20628,N_12036,N_13041);
or U20629 (N_20629,N_16336,N_13499);
and U20630 (N_20630,N_16707,N_13745);
and U20631 (N_20631,N_13069,N_17244);
xnor U20632 (N_20632,N_14818,N_13888);
nor U20633 (N_20633,N_15657,N_14424);
nand U20634 (N_20634,N_15144,N_14599);
or U20635 (N_20635,N_14704,N_12412);
nand U20636 (N_20636,N_16393,N_12969);
nor U20637 (N_20637,N_12457,N_15693);
and U20638 (N_20638,N_12838,N_16961);
and U20639 (N_20639,N_17804,N_12900);
and U20640 (N_20640,N_17829,N_13020);
nor U20641 (N_20641,N_16539,N_12326);
nor U20642 (N_20642,N_17595,N_13484);
nor U20643 (N_20643,N_12396,N_16538);
or U20644 (N_20644,N_15539,N_12665);
nand U20645 (N_20645,N_12025,N_15344);
xnor U20646 (N_20646,N_17493,N_15126);
xnor U20647 (N_20647,N_15763,N_14525);
or U20648 (N_20648,N_14050,N_14652);
or U20649 (N_20649,N_16304,N_17875);
xor U20650 (N_20650,N_13311,N_12093);
nor U20651 (N_20651,N_17071,N_16226);
or U20652 (N_20652,N_14752,N_12141);
or U20653 (N_20653,N_15835,N_15293);
or U20654 (N_20654,N_12338,N_16382);
and U20655 (N_20655,N_13999,N_13611);
xor U20656 (N_20656,N_13495,N_13975);
xor U20657 (N_20657,N_14582,N_17262);
and U20658 (N_20658,N_13810,N_14418);
and U20659 (N_20659,N_14833,N_12847);
xnor U20660 (N_20660,N_15466,N_14771);
or U20661 (N_20661,N_14192,N_14384);
or U20662 (N_20662,N_16716,N_16817);
and U20663 (N_20663,N_17210,N_14199);
and U20664 (N_20664,N_17660,N_14994);
or U20665 (N_20665,N_15818,N_13440);
nand U20666 (N_20666,N_12768,N_13289);
nor U20667 (N_20667,N_13960,N_13405);
or U20668 (N_20668,N_16641,N_15714);
or U20669 (N_20669,N_14147,N_16695);
and U20670 (N_20670,N_16549,N_14514);
xnor U20671 (N_20671,N_17072,N_13860);
nor U20672 (N_20672,N_14789,N_13904);
or U20673 (N_20673,N_16841,N_16623);
nor U20674 (N_20674,N_15008,N_13010);
xnor U20675 (N_20675,N_17243,N_16366);
or U20676 (N_20676,N_15355,N_15145);
nor U20677 (N_20677,N_13562,N_15957);
or U20678 (N_20678,N_16415,N_14597);
or U20679 (N_20679,N_17916,N_15326);
and U20680 (N_20680,N_14080,N_13714);
nor U20681 (N_20681,N_13189,N_16667);
and U20682 (N_20682,N_12430,N_15285);
nand U20683 (N_20683,N_15674,N_15136);
nor U20684 (N_20684,N_16545,N_15115);
nand U20685 (N_20685,N_17155,N_16540);
and U20686 (N_20686,N_12829,N_17624);
nand U20687 (N_20687,N_12451,N_16566);
or U20688 (N_20688,N_16185,N_13002);
nor U20689 (N_20689,N_13209,N_12585);
and U20690 (N_20690,N_14509,N_13446);
nand U20691 (N_20691,N_15945,N_13157);
or U20692 (N_20692,N_17132,N_12282);
xor U20693 (N_20693,N_17949,N_13119);
xnor U20694 (N_20694,N_12433,N_13433);
or U20695 (N_20695,N_13620,N_13396);
nand U20696 (N_20696,N_16721,N_12578);
or U20697 (N_20697,N_12130,N_12197);
xor U20698 (N_20698,N_16727,N_16831);
or U20699 (N_20699,N_12685,N_14436);
and U20700 (N_20700,N_12333,N_14324);
nor U20701 (N_20701,N_12380,N_14603);
or U20702 (N_20702,N_16070,N_16697);
xor U20703 (N_20703,N_17303,N_15361);
or U20704 (N_20704,N_17359,N_13190);
xnor U20705 (N_20705,N_17990,N_16399);
nand U20706 (N_20706,N_16642,N_16262);
and U20707 (N_20707,N_14817,N_14627);
xor U20708 (N_20708,N_12664,N_13775);
and U20709 (N_20709,N_15817,N_14120);
nand U20710 (N_20710,N_13420,N_14685);
xor U20711 (N_20711,N_12732,N_15127);
or U20712 (N_20712,N_13245,N_14851);
xnor U20713 (N_20713,N_17746,N_13857);
nand U20714 (N_20714,N_17675,N_13191);
and U20715 (N_20715,N_14793,N_12551);
and U20716 (N_20716,N_13432,N_12961);
xnor U20717 (N_20717,N_12309,N_14610);
and U20718 (N_20718,N_14450,N_14281);
and U20719 (N_20719,N_13100,N_12622);
nor U20720 (N_20720,N_15209,N_17090);
nand U20721 (N_20721,N_12276,N_15114);
and U20722 (N_20722,N_15758,N_14114);
nor U20723 (N_20723,N_14654,N_17439);
xnor U20724 (N_20724,N_16081,N_17122);
xnor U20725 (N_20725,N_13421,N_13174);
nand U20726 (N_20726,N_16073,N_12505);
nor U20727 (N_20727,N_16194,N_13302);
xnor U20728 (N_20728,N_15720,N_14282);
xnor U20729 (N_20729,N_17248,N_12261);
xnor U20730 (N_20730,N_13724,N_17951);
nand U20731 (N_20731,N_16844,N_14398);
nor U20732 (N_20732,N_17103,N_13962);
xor U20733 (N_20733,N_16745,N_15038);
and U20734 (N_20734,N_12663,N_16712);
nor U20735 (N_20735,N_16089,N_15220);
and U20736 (N_20736,N_15400,N_12469);
nor U20737 (N_20737,N_17938,N_13853);
nor U20738 (N_20738,N_14104,N_13456);
xor U20739 (N_20739,N_16595,N_13651);
nor U20740 (N_20740,N_16800,N_12675);
or U20741 (N_20741,N_17538,N_15319);
or U20742 (N_20742,N_14036,N_15433);
nand U20743 (N_20743,N_13469,N_12031);
nor U20744 (N_20744,N_15375,N_17682);
or U20745 (N_20745,N_13827,N_13880);
or U20746 (N_20746,N_14172,N_15717);
xnor U20747 (N_20747,N_14094,N_13004);
xor U20748 (N_20748,N_12992,N_17077);
nand U20749 (N_20749,N_17643,N_15246);
nor U20750 (N_20750,N_12450,N_12632);
nand U20751 (N_20751,N_14175,N_12823);
nor U20752 (N_20752,N_14366,N_17461);
xnor U20753 (N_20753,N_15857,N_14263);
nand U20754 (N_20754,N_13365,N_14728);
nand U20755 (N_20755,N_13893,N_12529);
nand U20756 (N_20756,N_14093,N_15531);
and U20757 (N_20757,N_15128,N_12627);
nand U20758 (N_20758,N_12955,N_14999);
nor U20759 (N_20759,N_16197,N_17151);
nand U20760 (N_20760,N_15749,N_12741);
or U20761 (N_20761,N_17442,N_14004);
and U20762 (N_20762,N_17550,N_13141);
nor U20763 (N_20763,N_15897,N_13913);
xnor U20764 (N_20764,N_15788,N_12177);
nor U20765 (N_20765,N_16141,N_17425);
xor U20766 (N_20766,N_16370,N_15195);
nor U20767 (N_20767,N_15087,N_16041);
and U20768 (N_20768,N_13083,N_13102);
or U20769 (N_20769,N_16867,N_13422);
and U20770 (N_20770,N_15234,N_12892);
xnor U20771 (N_20771,N_14145,N_16006);
xnor U20772 (N_20772,N_13945,N_14391);
and U20773 (N_20773,N_16491,N_16643);
xnor U20774 (N_20774,N_14656,N_14046);
xor U20775 (N_20775,N_13897,N_13771);
nand U20776 (N_20776,N_12586,N_14584);
nor U20777 (N_20777,N_13915,N_17314);
nor U20778 (N_20778,N_13079,N_16468);
nor U20779 (N_20779,N_16860,N_14169);
and U20780 (N_20780,N_17009,N_17111);
and U20781 (N_20781,N_17294,N_14260);
or U20782 (N_20782,N_12920,N_17206);
xnor U20783 (N_20783,N_15891,N_15631);
nor U20784 (N_20784,N_16876,N_16529);
nor U20785 (N_20785,N_15936,N_13478);
nor U20786 (N_20786,N_12633,N_17567);
nand U20787 (N_20787,N_14511,N_14204);
or U20788 (N_20788,N_14161,N_17264);
and U20789 (N_20789,N_16920,N_17819);
nand U20790 (N_20790,N_15639,N_15335);
xor U20791 (N_20791,N_13641,N_17426);
and U20792 (N_20792,N_13389,N_16683);
nand U20793 (N_20793,N_14762,N_13595);
nand U20794 (N_20794,N_17370,N_12370);
or U20795 (N_20795,N_13989,N_14611);
xnor U20796 (N_20796,N_16239,N_12871);
or U20797 (N_20797,N_14171,N_14378);
and U20798 (N_20798,N_17036,N_14683);
nor U20799 (N_20799,N_14118,N_16598);
or U20800 (N_20800,N_15057,N_13231);
and U20801 (N_20801,N_13352,N_15438);
nand U20802 (N_20802,N_17216,N_13266);
and U20803 (N_20803,N_13636,N_15028);
nand U20804 (N_20804,N_15205,N_12246);
and U20805 (N_20805,N_13783,N_12657);
or U20806 (N_20806,N_15152,N_17047);
xor U20807 (N_20807,N_16773,N_16469);
and U20808 (N_20808,N_15192,N_12391);
nor U20809 (N_20809,N_14672,N_16083);
and U20810 (N_20810,N_14358,N_13681);
and U20811 (N_20811,N_16952,N_17533);
or U20812 (N_20812,N_12534,N_15930);
nor U20813 (N_20813,N_15215,N_16947);
or U20814 (N_20814,N_16358,N_16137);
nor U20815 (N_20815,N_16762,N_15792);
and U20816 (N_20816,N_14148,N_17463);
nor U20817 (N_20817,N_14844,N_17863);
xor U20818 (N_20818,N_16999,N_13062);
nor U20819 (N_20819,N_13720,N_16983);
and U20820 (N_20820,N_17585,N_14754);
nor U20821 (N_20821,N_14469,N_14504);
nor U20822 (N_20822,N_17086,N_13685);
and U20823 (N_20823,N_15362,N_12949);
nor U20824 (N_20824,N_13293,N_12200);
nand U20825 (N_20825,N_16696,N_13848);
nor U20826 (N_20826,N_15473,N_14717);
nand U20827 (N_20827,N_15419,N_12857);
and U20828 (N_20828,N_15368,N_14645);
and U20829 (N_20829,N_16476,N_14220);
and U20830 (N_20830,N_15636,N_13133);
or U20831 (N_20831,N_14975,N_13367);
nor U20832 (N_20832,N_13066,N_12619);
nand U20833 (N_20833,N_17494,N_13891);
nor U20834 (N_20834,N_14830,N_12421);
xnor U20835 (N_20835,N_16688,N_17300);
xnor U20836 (N_20836,N_12508,N_17807);
or U20837 (N_20837,N_15270,N_12205);
xnor U20838 (N_20838,N_16481,N_13767);
or U20839 (N_20839,N_14318,N_17930);
nor U20840 (N_20840,N_13742,N_15170);
or U20841 (N_20841,N_13917,N_14670);
or U20842 (N_20842,N_13297,N_13766);
xnor U20843 (N_20843,N_14326,N_16756);
nor U20844 (N_20844,N_17325,N_12032);
nand U20845 (N_20845,N_12753,N_16412);
and U20846 (N_20846,N_12439,N_16792);
nand U20847 (N_20847,N_16915,N_16863);
nand U20848 (N_20848,N_14230,N_15659);
xor U20849 (N_20849,N_13059,N_12669);
xnor U20850 (N_20850,N_16152,N_12897);
or U20851 (N_20851,N_14834,N_12463);
xor U20852 (N_20852,N_13722,N_15406);
and U20853 (N_20853,N_12709,N_17355);
nand U20854 (N_20854,N_17574,N_12699);
nor U20855 (N_20855,N_17853,N_15211);
xor U20856 (N_20856,N_15668,N_14621);
or U20857 (N_20857,N_16029,N_15608);
xor U20858 (N_20858,N_12251,N_17857);
nand U20859 (N_20859,N_17160,N_15266);
and U20860 (N_20860,N_17431,N_16771);
xnor U20861 (N_20861,N_15685,N_17778);
nand U20862 (N_20862,N_16280,N_12861);
or U20863 (N_20863,N_14142,N_17912);
or U20864 (N_20864,N_13271,N_12153);
nand U20865 (N_20865,N_13243,N_12549);
and U20866 (N_20866,N_14226,N_17108);
or U20867 (N_20867,N_16862,N_17481);
xnor U20868 (N_20868,N_12485,N_13933);
or U20869 (N_20869,N_15267,N_15845);
and U20870 (N_20870,N_17271,N_14665);
nand U20871 (N_20871,N_17768,N_15418);
nand U20872 (N_20872,N_14271,N_14889);
nor U20873 (N_20873,N_14944,N_13475);
xnor U20874 (N_20874,N_15899,N_17577);
or U20875 (N_20875,N_16774,N_13727);
or U20876 (N_20876,N_17436,N_13058);
nor U20877 (N_20877,N_15735,N_12995);
nand U20878 (N_20878,N_12256,N_14979);
nand U20879 (N_20879,N_17510,N_17932);
and U20880 (N_20880,N_16752,N_17909);
nor U20881 (N_20881,N_12743,N_14546);
xnor U20882 (N_20882,N_16749,N_12027);
nor U20883 (N_20883,N_17486,N_13442);
xor U20884 (N_20884,N_13995,N_12989);
and U20885 (N_20885,N_14067,N_13532);
xor U20886 (N_20886,N_13491,N_13943);
or U20887 (N_20887,N_13006,N_12119);
and U20888 (N_20888,N_16278,N_15347);
or U20889 (N_20889,N_14776,N_14232);
or U20890 (N_20890,N_14962,N_16890);
xnor U20891 (N_20891,N_13260,N_14413);
and U20892 (N_20892,N_16882,N_15298);
nand U20893 (N_20893,N_12842,N_14694);
or U20894 (N_20894,N_13678,N_15226);
nor U20895 (N_20895,N_17825,N_13255);
xor U20896 (N_20896,N_16091,N_14607);
xor U20897 (N_20897,N_17193,N_15959);
or U20898 (N_20898,N_17475,N_16896);
or U20899 (N_20899,N_14299,N_12798);
xor U20900 (N_20900,N_13959,N_15841);
nor U20901 (N_20901,N_16157,N_14085);
and U20902 (N_20902,N_12971,N_17152);
nor U20903 (N_20903,N_15490,N_12597);
nand U20904 (N_20904,N_14950,N_14455);
and U20905 (N_20905,N_13168,N_16242);
xor U20906 (N_20906,N_12548,N_13998);
nor U20907 (N_20907,N_16355,N_16133);
or U20908 (N_20908,N_12001,N_16423);
xor U20909 (N_20909,N_15823,N_14544);
xor U20910 (N_20910,N_12591,N_16060);
nor U20911 (N_20911,N_14451,N_14847);
nand U20912 (N_20912,N_12318,N_12962);
nor U20913 (N_20913,N_17841,N_16019);
or U20914 (N_20914,N_14917,N_12614);
or U20915 (N_20915,N_15275,N_12896);
nor U20916 (N_20916,N_14483,N_14445);
or U20917 (N_20917,N_12263,N_12052);
or U20918 (N_20918,N_14701,N_16611);
nor U20919 (N_20919,N_12189,N_12332);
and U20920 (N_20920,N_14174,N_13545);
and U20921 (N_20921,N_14396,N_12948);
or U20922 (N_20922,N_17211,N_15067);
or U20923 (N_20923,N_16143,N_12233);
or U20924 (N_20924,N_12285,N_15643);
nand U20925 (N_20925,N_17793,N_12512);
nand U20926 (N_20926,N_14891,N_17419);
nor U20927 (N_20927,N_15570,N_12553);
nand U20928 (N_20928,N_13793,N_17450);
nand U20929 (N_20929,N_16418,N_15309);
nor U20930 (N_20930,N_16015,N_17399);
nor U20931 (N_20931,N_13555,N_12471);
nand U20932 (N_20932,N_13567,N_14167);
nor U20933 (N_20933,N_17739,N_14932);
and U20934 (N_20934,N_17850,N_13955);
xnor U20935 (N_20935,N_14775,N_12023);
nand U20936 (N_20936,N_13304,N_17456);
xnor U20937 (N_20937,N_17063,N_13516);
nor U20938 (N_20938,N_12819,N_15690);
nor U20939 (N_20939,N_16488,N_13890);
or U20940 (N_20940,N_12266,N_16492);
nand U20941 (N_20941,N_17386,N_12916);
xnor U20942 (N_20942,N_14389,N_15198);
or U20943 (N_20943,N_12588,N_14657);
xnor U20944 (N_20944,N_13667,N_16518);
xnor U20945 (N_20945,N_16908,N_12144);
or U20946 (N_20946,N_15364,N_15548);
xor U20947 (N_20947,N_17195,N_15081);
xor U20948 (N_20948,N_13263,N_13730);
xnor U20949 (N_20949,N_17727,N_17507);
nand U20950 (N_20950,N_12905,N_13114);
xnor U20951 (N_20951,N_16017,N_13361);
nand U20952 (N_20952,N_14317,N_12943);
or U20953 (N_20953,N_12374,N_13593);
nor U20954 (N_20954,N_16272,N_17756);
nor U20955 (N_20955,N_12491,N_14618);
nand U20956 (N_20956,N_12062,N_17797);
nor U20957 (N_20957,N_12799,N_12465);
or U20958 (N_20958,N_12705,N_15491);
nand U20959 (N_20959,N_16168,N_16647);
or U20960 (N_20960,N_16115,N_15149);
nand U20961 (N_20961,N_15387,N_17602);
xnor U20962 (N_20962,N_13434,N_12932);
or U20963 (N_20963,N_15694,N_17576);
nor U20964 (N_20964,N_12877,N_15612);
xnor U20965 (N_20965,N_14869,N_17801);
or U20966 (N_20966,N_17269,N_14804);
xnor U20967 (N_20967,N_17869,N_16371);
and U20968 (N_20968,N_15644,N_14168);
nand U20969 (N_20969,N_12486,N_14245);
xor U20970 (N_20970,N_16241,N_17022);
xor U20971 (N_20971,N_15913,N_14846);
or U20972 (N_20972,N_17101,N_14302);
xnor U20973 (N_20973,N_16637,N_17955);
xor U20974 (N_20974,N_16217,N_14254);
nand U20975 (N_20975,N_17209,N_13107);
or U20976 (N_20976,N_17006,N_16188);
or U20977 (N_20977,N_16165,N_16849);
or U20978 (N_20978,N_12198,N_14862);
and U20979 (N_20979,N_14886,N_15121);
or U20980 (N_20980,N_16548,N_13590);
xnor U20981 (N_20981,N_16609,N_14903);
xor U20982 (N_20982,N_14680,N_15829);
or U20983 (N_20983,N_14575,N_14692);
nor U20984 (N_20984,N_13060,N_15457);
nand U20985 (N_20985,N_12912,N_17845);
and U20986 (N_20986,N_17701,N_12561);
and U20987 (N_20987,N_15887,N_16746);
and U20988 (N_20988,N_13292,N_15348);
or U20989 (N_20989,N_13353,N_16416);
nand U20990 (N_20990,N_17876,N_14454);
or U20991 (N_20991,N_14057,N_17561);
or U20992 (N_20992,N_15566,N_16392);
xor U20993 (N_20993,N_12245,N_17051);
and U20994 (N_20994,N_17812,N_14181);
or U20995 (N_20995,N_15683,N_17137);
nand U20996 (N_20996,N_15940,N_13765);
xor U20997 (N_20997,N_14738,N_12264);
and U20998 (N_20998,N_14246,N_14615);
nor U20999 (N_20999,N_15795,N_12128);
or U21000 (N_21000,N_16974,N_14204);
nor U21001 (N_21001,N_12250,N_12050);
nor U21002 (N_21002,N_16414,N_12753);
nor U21003 (N_21003,N_14059,N_14746);
and U21004 (N_21004,N_17398,N_17435);
nand U21005 (N_21005,N_12491,N_14513);
nor U21006 (N_21006,N_15269,N_16380);
or U21007 (N_21007,N_13691,N_14731);
xor U21008 (N_21008,N_15583,N_16679);
and U21009 (N_21009,N_16531,N_17418);
xnor U21010 (N_21010,N_16560,N_15424);
and U21011 (N_21011,N_13713,N_17838);
and U21012 (N_21012,N_16042,N_17537);
or U21013 (N_21013,N_14624,N_15141);
nor U21014 (N_21014,N_12231,N_16565);
or U21015 (N_21015,N_17750,N_13506);
xnor U21016 (N_21016,N_13706,N_14217);
and U21017 (N_21017,N_14993,N_16099);
or U21018 (N_21018,N_13768,N_15899);
or U21019 (N_21019,N_17081,N_17947);
xor U21020 (N_21020,N_17908,N_13795);
or U21021 (N_21021,N_15957,N_12273);
xor U21022 (N_21022,N_16477,N_15434);
or U21023 (N_21023,N_15461,N_12937);
xor U21024 (N_21024,N_17823,N_12887);
or U21025 (N_21025,N_15268,N_14065);
nor U21026 (N_21026,N_16802,N_16645);
nand U21027 (N_21027,N_12440,N_14266);
xnor U21028 (N_21028,N_17487,N_12335);
nand U21029 (N_21029,N_17987,N_17732);
nand U21030 (N_21030,N_15650,N_14375);
xnor U21031 (N_21031,N_12352,N_12219);
xor U21032 (N_21032,N_13778,N_13891);
nand U21033 (N_21033,N_14200,N_13024);
or U21034 (N_21034,N_15214,N_16179);
xor U21035 (N_21035,N_15642,N_13651);
xnor U21036 (N_21036,N_15808,N_15495);
or U21037 (N_21037,N_13102,N_15143);
and U21038 (N_21038,N_17806,N_16610);
xor U21039 (N_21039,N_15893,N_17672);
xnor U21040 (N_21040,N_16176,N_15554);
nor U21041 (N_21041,N_13270,N_14318);
and U21042 (N_21042,N_13411,N_14306);
xor U21043 (N_21043,N_15209,N_13193);
and U21044 (N_21044,N_13142,N_12670);
nand U21045 (N_21045,N_15231,N_16809);
nor U21046 (N_21046,N_16055,N_14532);
nor U21047 (N_21047,N_16255,N_15525);
xor U21048 (N_21048,N_13374,N_13015);
and U21049 (N_21049,N_17019,N_17565);
nor U21050 (N_21050,N_16928,N_14306);
or U21051 (N_21051,N_13513,N_13699);
nand U21052 (N_21052,N_14554,N_16028);
nand U21053 (N_21053,N_12985,N_16721);
or U21054 (N_21054,N_14983,N_13820);
or U21055 (N_21055,N_16670,N_14999);
and U21056 (N_21056,N_15092,N_12587);
or U21057 (N_21057,N_13420,N_15624);
xnor U21058 (N_21058,N_13929,N_16108);
nor U21059 (N_21059,N_15933,N_14285);
and U21060 (N_21060,N_14830,N_12564);
and U21061 (N_21061,N_16440,N_14620);
and U21062 (N_21062,N_12119,N_14602);
nor U21063 (N_21063,N_16394,N_12619);
nor U21064 (N_21064,N_15759,N_12288);
and U21065 (N_21065,N_12258,N_14578);
nand U21066 (N_21066,N_12210,N_14769);
or U21067 (N_21067,N_12639,N_17573);
nand U21068 (N_21068,N_12042,N_16740);
nand U21069 (N_21069,N_13189,N_16003);
xnor U21070 (N_21070,N_15102,N_13149);
xor U21071 (N_21071,N_13698,N_13768);
or U21072 (N_21072,N_16638,N_12626);
nor U21073 (N_21073,N_17622,N_14215);
or U21074 (N_21074,N_13846,N_14458);
xor U21075 (N_21075,N_12014,N_17783);
and U21076 (N_21076,N_13509,N_15341);
or U21077 (N_21077,N_15640,N_12449);
nor U21078 (N_21078,N_17511,N_16012);
xor U21079 (N_21079,N_17653,N_15673);
nand U21080 (N_21080,N_14835,N_16391);
nand U21081 (N_21081,N_17586,N_14804);
xnor U21082 (N_21082,N_15263,N_17046);
xnor U21083 (N_21083,N_15685,N_15727);
nand U21084 (N_21084,N_12499,N_16064);
nand U21085 (N_21085,N_17302,N_15809);
xnor U21086 (N_21086,N_15841,N_17457);
xor U21087 (N_21087,N_13006,N_16083);
xnor U21088 (N_21088,N_14644,N_15431);
nand U21089 (N_21089,N_13051,N_15602);
or U21090 (N_21090,N_15132,N_17011);
xnor U21091 (N_21091,N_13292,N_13244);
and U21092 (N_21092,N_16446,N_12530);
and U21093 (N_21093,N_15675,N_13866);
and U21094 (N_21094,N_14666,N_17754);
and U21095 (N_21095,N_15208,N_15491);
nor U21096 (N_21096,N_12948,N_14464);
xor U21097 (N_21097,N_15003,N_15086);
xnor U21098 (N_21098,N_12097,N_16222);
or U21099 (N_21099,N_16206,N_15892);
xnor U21100 (N_21100,N_14847,N_16079);
or U21101 (N_21101,N_13155,N_13089);
nor U21102 (N_21102,N_14457,N_17689);
nor U21103 (N_21103,N_15868,N_17492);
nand U21104 (N_21104,N_14774,N_16114);
and U21105 (N_21105,N_15430,N_15526);
nor U21106 (N_21106,N_17028,N_13242);
xnor U21107 (N_21107,N_17925,N_17227);
xnor U21108 (N_21108,N_16079,N_12671);
xnor U21109 (N_21109,N_15830,N_16029);
nand U21110 (N_21110,N_15301,N_14304);
nand U21111 (N_21111,N_13027,N_15425);
or U21112 (N_21112,N_16939,N_15850);
and U21113 (N_21113,N_13370,N_14840);
and U21114 (N_21114,N_16187,N_12497);
xor U21115 (N_21115,N_14724,N_15475);
and U21116 (N_21116,N_13355,N_12884);
and U21117 (N_21117,N_13306,N_15109);
xor U21118 (N_21118,N_13480,N_16585);
nand U21119 (N_21119,N_13109,N_14322);
or U21120 (N_21120,N_14147,N_13927);
or U21121 (N_21121,N_13164,N_13165);
or U21122 (N_21122,N_16783,N_14083);
nor U21123 (N_21123,N_15216,N_12468);
xor U21124 (N_21124,N_15179,N_14874);
xnor U21125 (N_21125,N_16787,N_12230);
xor U21126 (N_21126,N_17739,N_15704);
and U21127 (N_21127,N_16838,N_14031);
nor U21128 (N_21128,N_17234,N_14121);
nor U21129 (N_21129,N_14653,N_13073);
nand U21130 (N_21130,N_12470,N_17852);
xnor U21131 (N_21131,N_13853,N_16621);
or U21132 (N_21132,N_13396,N_13102);
nor U21133 (N_21133,N_14352,N_17779);
xor U21134 (N_21134,N_17920,N_17983);
nor U21135 (N_21135,N_14401,N_15924);
or U21136 (N_21136,N_12765,N_13281);
xor U21137 (N_21137,N_12294,N_12148);
or U21138 (N_21138,N_14035,N_16556);
nand U21139 (N_21139,N_12538,N_16661);
nor U21140 (N_21140,N_15640,N_13874);
or U21141 (N_21141,N_12446,N_16327);
xor U21142 (N_21142,N_14099,N_17358);
nand U21143 (N_21143,N_16635,N_15424);
and U21144 (N_21144,N_12923,N_16026);
xor U21145 (N_21145,N_16189,N_13803);
nand U21146 (N_21146,N_15653,N_16014);
xnor U21147 (N_21147,N_14761,N_14140);
and U21148 (N_21148,N_12592,N_14559);
or U21149 (N_21149,N_13497,N_14543);
xnor U21150 (N_21150,N_13765,N_13413);
nand U21151 (N_21151,N_14650,N_14553);
nand U21152 (N_21152,N_16446,N_17511);
and U21153 (N_21153,N_12060,N_14428);
xor U21154 (N_21154,N_16930,N_17038);
nor U21155 (N_21155,N_15453,N_17252);
and U21156 (N_21156,N_14019,N_14864);
nand U21157 (N_21157,N_16240,N_14648);
or U21158 (N_21158,N_12925,N_14172);
xnor U21159 (N_21159,N_14028,N_14709);
and U21160 (N_21160,N_16390,N_12459);
or U21161 (N_21161,N_15278,N_12500);
or U21162 (N_21162,N_15079,N_14205);
nand U21163 (N_21163,N_13973,N_16364);
or U21164 (N_21164,N_12967,N_17812);
xnor U21165 (N_21165,N_15630,N_16315);
or U21166 (N_21166,N_13349,N_12640);
xnor U21167 (N_21167,N_16272,N_14775);
or U21168 (N_21168,N_12546,N_16538);
and U21169 (N_21169,N_13076,N_15870);
nand U21170 (N_21170,N_12838,N_12830);
and U21171 (N_21171,N_17469,N_13082);
nor U21172 (N_21172,N_12365,N_14369);
nand U21173 (N_21173,N_15216,N_12639);
and U21174 (N_21174,N_16799,N_15509);
xnor U21175 (N_21175,N_15698,N_14497);
or U21176 (N_21176,N_15191,N_12606);
or U21177 (N_21177,N_17095,N_12350);
or U21178 (N_21178,N_12698,N_16574);
xnor U21179 (N_21179,N_16478,N_17301);
nand U21180 (N_21180,N_12587,N_13767);
nand U21181 (N_21181,N_15395,N_14687);
xnor U21182 (N_21182,N_15552,N_15478);
nor U21183 (N_21183,N_15076,N_14126);
nor U21184 (N_21184,N_14724,N_14197);
or U21185 (N_21185,N_17933,N_14487);
xnor U21186 (N_21186,N_15780,N_14251);
xnor U21187 (N_21187,N_15588,N_15959);
xor U21188 (N_21188,N_12382,N_12477);
and U21189 (N_21189,N_13806,N_13260);
and U21190 (N_21190,N_17633,N_12004);
xnor U21191 (N_21191,N_17217,N_13370);
and U21192 (N_21192,N_13566,N_12786);
or U21193 (N_21193,N_15605,N_17081);
nand U21194 (N_21194,N_15901,N_12274);
xnor U21195 (N_21195,N_13846,N_15238);
and U21196 (N_21196,N_14947,N_16323);
and U21197 (N_21197,N_12693,N_14757);
or U21198 (N_21198,N_12822,N_13100);
xnor U21199 (N_21199,N_15753,N_13856);
or U21200 (N_21200,N_17381,N_16630);
nor U21201 (N_21201,N_13561,N_13087);
and U21202 (N_21202,N_16803,N_14100);
and U21203 (N_21203,N_12533,N_15225);
or U21204 (N_21204,N_17561,N_14141);
nor U21205 (N_21205,N_12592,N_16182);
or U21206 (N_21206,N_15395,N_14256);
and U21207 (N_21207,N_17704,N_12791);
xnor U21208 (N_21208,N_13536,N_12081);
and U21209 (N_21209,N_17629,N_17042);
xor U21210 (N_21210,N_17609,N_15992);
nand U21211 (N_21211,N_12215,N_14855);
nor U21212 (N_21212,N_13420,N_15316);
nand U21213 (N_21213,N_14874,N_17037);
xnor U21214 (N_21214,N_12715,N_14967);
nor U21215 (N_21215,N_15266,N_13136);
xnor U21216 (N_21216,N_14527,N_16758);
or U21217 (N_21217,N_16805,N_13431);
nor U21218 (N_21218,N_12118,N_16962);
nand U21219 (N_21219,N_15616,N_17360);
xor U21220 (N_21220,N_13719,N_15802);
nor U21221 (N_21221,N_13337,N_17784);
xor U21222 (N_21222,N_15030,N_16786);
nand U21223 (N_21223,N_14753,N_15775);
nor U21224 (N_21224,N_12472,N_14365);
or U21225 (N_21225,N_13243,N_14574);
nor U21226 (N_21226,N_15891,N_17533);
or U21227 (N_21227,N_16731,N_16498);
xnor U21228 (N_21228,N_16213,N_14040);
and U21229 (N_21229,N_15560,N_16711);
xor U21230 (N_21230,N_15365,N_17148);
nand U21231 (N_21231,N_13499,N_14121);
or U21232 (N_21232,N_15375,N_12111);
xor U21233 (N_21233,N_13846,N_14809);
or U21234 (N_21234,N_13348,N_13607);
xor U21235 (N_21235,N_17050,N_15694);
and U21236 (N_21236,N_15393,N_13138);
and U21237 (N_21237,N_16395,N_14458);
and U21238 (N_21238,N_14758,N_13024);
or U21239 (N_21239,N_16280,N_13500);
or U21240 (N_21240,N_16666,N_17855);
nor U21241 (N_21241,N_15073,N_13674);
and U21242 (N_21242,N_15478,N_12847);
nand U21243 (N_21243,N_13896,N_12124);
and U21244 (N_21244,N_17126,N_17409);
and U21245 (N_21245,N_17698,N_13570);
xor U21246 (N_21246,N_14920,N_14838);
or U21247 (N_21247,N_16471,N_14649);
xor U21248 (N_21248,N_16533,N_14237);
nand U21249 (N_21249,N_12223,N_16111);
and U21250 (N_21250,N_14256,N_15985);
nor U21251 (N_21251,N_15528,N_13471);
or U21252 (N_21252,N_17973,N_15209);
and U21253 (N_21253,N_13218,N_14326);
nand U21254 (N_21254,N_12107,N_17443);
and U21255 (N_21255,N_14724,N_13732);
and U21256 (N_21256,N_13687,N_16352);
nand U21257 (N_21257,N_16620,N_15402);
or U21258 (N_21258,N_17325,N_12080);
or U21259 (N_21259,N_15050,N_17032);
or U21260 (N_21260,N_14606,N_17493);
and U21261 (N_21261,N_15606,N_13330);
xnor U21262 (N_21262,N_12879,N_14196);
or U21263 (N_21263,N_13979,N_17000);
or U21264 (N_21264,N_12109,N_12400);
nand U21265 (N_21265,N_17082,N_15013);
and U21266 (N_21266,N_17515,N_14954);
nor U21267 (N_21267,N_15083,N_14202);
nor U21268 (N_21268,N_14163,N_16074);
nor U21269 (N_21269,N_12933,N_14440);
nand U21270 (N_21270,N_15360,N_15023);
and U21271 (N_21271,N_12156,N_17430);
nor U21272 (N_21272,N_17723,N_17410);
and U21273 (N_21273,N_15465,N_17443);
nand U21274 (N_21274,N_13061,N_15197);
xor U21275 (N_21275,N_15564,N_17681);
or U21276 (N_21276,N_16989,N_13541);
nor U21277 (N_21277,N_17403,N_17814);
or U21278 (N_21278,N_15640,N_13764);
nor U21279 (N_21279,N_15925,N_12054);
nand U21280 (N_21280,N_14818,N_14844);
and U21281 (N_21281,N_16463,N_14633);
nand U21282 (N_21282,N_12821,N_16348);
nand U21283 (N_21283,N_12667,N_17539);
or U21284 (N_21284,N_14733,N_15195);
xnor U21285 (N_21285,N_15386,N_12264);
and U21286 (N_21286,N_16282,N_17432);
and U21287 (N_21287,N_17404,N_14388);
nand U21288 (N_21288,N_16079,N_14354);
nor U21289 (N_21289,N_17306,N_14186);
nand U21290 (N_21290,N_17958,N_12042);
xnor U21291 (N_21291,N_13897,N_14422);
and U21292 (N_21292,N_12360,N_14630);
nand U21293 (N_21293,N_17888,N_12134);
or U21294 (N_21294,N_12005,N_13726);
and U21295 (N_21295,N_14219,N_15020);
nand U21296 (N_21296,N_12344,N_16621);
nor U21297 (N_21297,N_15047,N_13713);
and U21298 (N_21298,N_14280,N_16697);
and U21299 (N_21299,N_12721,N_15329);
nand U21300 (N_21300,N_12551,N_16863);
nor U21301 (N_21301,N_13192,N_13240);
and U21302 (N_21302,N_15747,N_12306);
or U21303 (N_21303,N_16734,N_14136);
xor U21304 (N_21304,N_15025,N_14022);
nor U21305 (N_21305,N_13994,N_15044);
and U21306 (N_21306,N_16793,N_12874);
or U21307 (N_21307,N_17200,N_15910);
or U21308 (N_21308,N_16862,N_14197);
and U21309 (N_21309,N_15674,N_15756);
nand U21310 (N_21310,N_16626,N_14070);
and U21311 (N_21311,N_15280,N_14419);
or U21312 (N_21312,N_15956,N_14681);
and U21313 (N_21313,N_17617,N_14512);
nor U21314 (N_21314,N_15672,N_14026);
and U21315 (N_21315,N_15753,N_13116);
xnor U21316 (N_21316,N_13995,N_13499);
and U21317 (N_21317,N_15338,N_17761);
nand U21318 (N_21318,N_13667,N_12031);
xnor U21319 (N_21319,N_14459,N_15443);
nand U21320 (N_21320,N_16496,N_13960);
xor U21321 (N_21321,N_15950,N_17719);
xor U21322 (N_21322,N_13572,N_17894);
nand U21323 (N_21323,N_17307,N_12953);
nand U21324 (N_21324,N_15947,N_13653);
or U21325 (N_21325,N_14693,N_14486);
nor U21326 (N_21326,N_12258,N_13899);
and U21327 (N_21327,N_16491,N_14865);
xor U21328 (N_21328,N_12095,N_15507);
xnor U21329 (N_21329,N_16919,N_15233);
or U21330 (N_21330,N_12533,N_12191);
nor U21331 (N_21331,N_13947,N_16524);
nand U21332 (N_21332,N_14917,N_12714);
nand U21333 (N_21333,N_16037,N_17254);
xor U21334 (N_21334,N_12686,N_14380);
and U21335 (N_21335,N_16895,N_13757);
nand U21336 (N_21336,N_17555,N_12843);
nand U21337 (N_21337,N_12755,N_14120);
xor U21338 (N_21338,N_13277,N_17206);
xnor U21339 (N_21339,N_16828,N_15335);
or U21340 (N_21340,N_12939,N_14456);
nand U21341 (N_21341,N_12541,N_14527);
nand U21342 (N_21342,N_14304,N_15551);
nand U21343 (N_21343,N_12761,N_15974);
or U21344 (N_21344,N_15636,N_14070);
xor U21345 (N_21345,N_15817,N_13510);
and U21346 (N_21346,N_15032,N_13864);
and U21347 (N_21347,N_13038,N_12167);
nand U21348 (N_21348,N_15656,N_13599);
and U21349 (N_21349,N_16625,N_15682);
nor U21350 (N_21350,N_14793,N_17783);
nor U21351 (N_21351,N_12932,N_12705);
nor U21352 (N_21352,N_13184,N_17969);
and U21353 (N_21353,N_15541,N_15309);
nor U21354 (N_21354,N_15160,N_12600);
or U21355 (N_21355,N_16718,N_15402);
xor U21356 (N_21356,N_17214,N_12945);
nor U21357 (N_21357,N_17461,N_12423);
xor U21358 (N_21358,N_13281,N_16942);
or U21359 (N_21359,N_17952,N_17408);
nor U21360 (N_21360,N_13921,N_15663);
and U21361 (N_21361,N_16563,N_17382);
xor U21362 (N_21362,N_12357,N_17889);
xnor U21363 (N_21363,N_16791,N_16749);
xor U21364 (N_21364,N_12025,N_14837);
and U21365 (N_21365,N_14561,N_16451);
or U21366 (N_21366,N_12977,N_17699);
or U21367 (N_21367,N_16950,N_14227);
xor U21368 (N_21368,N_16545,N_17438);
nand U21369 (N_21369,N_17526,N_13607);
or U21370 (N_21370,N_12689,N_15828);
or U21371 (N_21371,N_13593,N_15597);
and U21372 (N_21372,N_16522,N_12949);
nor U21373 (N_21373,N_14674,N_13088);
nand U21374 (N_21374,N_12346,N_14515);
nand U21375 (N_21375,N_16203,N_16273);
and U21376 (N_21376,N_17742,N_13700);
or U21377 (N_21377,N_14373,N_17346);
or U21378 (N_21378,N_13444,N_16951);
and U21379 (N_21379,N_17057,N_15620);
nor U21380 (N_21380,N_13956,N_13664);
xnor U21381 (N_21381,N_17983,N_16489);
and U21382 (N_21382,N_17242,N_13607);
and U21383 (N_21383,N_14717,N_12878);
or U21384 (N_21384,N_16775,N_14619);
nand U21385 (N_21385,N_16761,N_16476);
or U21386 (N_21386,N_15659,N_15577);
xor U21387 (N_21387,N_16347,N_13183);
and U21388 (N_21388,N_16638,N_16065);
and U21389 (N_21389,N_12909,N_16468);
nand U21390 (N_21390,N_16088,N_13649);
nand U21391 (N_21391,N_12251,N_16142);
nor U21392 (N_21392,N_17347,N_13465);
nor U21393 (N_21393,N_16774,N_16356);
nor U21394 (N_21394,N_14881,N_17951);
nor U21395 (N_21395,N_16686,N_15817);
or U21396 (N_21396,N_17864,N_13779);
nand U21397 (N_21397,N_12226,N_15322);
nor U21398 (N_21398,N_15397,N_12404);
xnor U21399 (N_21399,N_13431,N_17905);
and U21400 (N_21400,N_14323,N_13280);
and U21401 (N_21401,N_14013,N_13567);
and U21402 (N_21402,N_13306,N_17128);
and U21403 (N_21403,N_17344,N_14464);
or U21404 (N_21404,N_12857,N_14729);
nor U21405 (N_21405,N_15404,N_16719);
xnor U21406 (N_21406,N_17628,N_15114);
or U21407 (N_21407,N_17668,N_12686);
or U21408 (N_21408,N_16414,N_15855);
or U21409 (N_21409,N_13185,N_13860);
xor U21410 (N_21410,N_14258,N_15095);
nand U21411 (N_21411,N_13312,N_16185);
and U21412 (N_21412,N_12115,N_16972);
and U21413 (N_21413,N_12508,N_13363);
xnor U21414 (N_21414,N_16639,N_16733);
and U21415 (N_21415,N_17102,N_16662);
nand U21416 (N_21416,N_17491,N_14261);
xor U21417 (N_21417,N_12001,N_14014);
nand U21418 (N_21418,N_17360,N_14347);
or U21419 (N_21419,N_12091,N_14181);
xnor U21420 (N_21420,N_13650,N_13663);
nor U21421 (N_21421,N_16813,N_13535);
xnor U21422 (N_21422,N_16824,N_17838);
nor U21423 (N_21423,N_13517,N_17911);
or U21424 (N_21424,N_14491,N_17092);
and U21425 (N_21425,N_12228,N_13448);
xnor U21426 (N_21426,N_14885,N_13105);
and U21427 (N_21427,N_14417,N_12692);
or U21428 (N_21428,N_12870,N_17419);
nand U21429 (N_21429,N_13064,N_15050);
nand U21430 (N_21430,N_17810,N_16395);
or U21431 (N_21431,N_17214,N_16644);
nand U21432 (N_21432,N_16634,N_16918);
or U21433 (N_21433,N_17547,N_14763);
or U21434 (N_21434,N_17194,N_13064);
and U21435 (N_21435,N_14184,N_12188);
nor U21436 (N_21436,N_16458,N_12990);
or U21437 (N_21437,N_12675,N_16205);
nand U21438 (N_21438,N_15373,N_13405);
nor U21439 (N_21439,N_13536,N_16502);
nand U21440 (N_21440,N_17698,N_15918);
xnor U21441 (N_21441,N_13355,N_14978);
and U21442 (N_21442,N_12211,N_13715);
nor U21443 (N_21443,N_13326,N_17927);
xnor U21444 (N_21444,N_14439,N_14306);
and U21445 (N_21445,N_12662,N_12818);
or U21446 (N_21446,N_14186,N_15643);
xnor U21447 (N_21447,N_15094,N_12939);
nand U21448 (N_21448,N_14628,N_13941);
nand U21449 (N_21449,N_14111,N_14587);
or U21450 (N_21450,N_12558,N_12915);
nand U21451 (N_21451,N_15129,N_16443);
or U21452 (N_21452,N_17002,N_16731);
xor U21453 (N_21453,N_15808,N_12948);
nor U21454 (N_21454,N_14742,N_13497);
xor U21455 (N_21455,N_15396,N_13551);
nor U21456 (N_21456,N_15955,N_13664);
or U21457 (N_21457,N_15295,N_13339);
nor U21458 (N_21458,N_14032,N_17983);
xor U21459 (N_21459,N_12702,N_13854);
and U21460 (N_21460,N_16103,N_15916);
and U21461 (N_21461,N_17375,N_15925);
xnor U21462 (N_21462,N_16933,N_16963);
nand U21463 (N_21463,N_12368,N_14553);
xor U21464 (N_21464,N_16764,N_13318);
nand U21465 (N_21465,N_15166,N_16239);
or U21466 (N_21466,N_15987,N_17601);
xor U21467 (N_21467,N_14989,N_16965);
and U21468 (N_21468,N_16399,N_14148);
and U21469 (N_21469,N_16899,N_12142);
nand U21470 (N_21470,N_15289,N_16221);
and U21471 (N_21471,N_13098,N_16470);
nor U21472 (N_21472,N_17112,N_12507);
or U21473 (N_21473,N_15301,N_16159);
xnor U21474 (N_21474,N_13784,N_12399);
nor U21475 (N_21475,N_17767,N_15354);
nand U21476 (N_21476,N_13131,N_15486);
nand U21477 (N_21477,N_12000,N_15147);
xor U21478 (N_21478,N_16735,N_14672);
nor U21479 (N_21479,N_15190,N_12989);
xor U21480 (N_21480,N_14243,N_14850);
nand U21481 (N_21481,N_14200,N_12444);
nand U21482 (N_21482,N_15194,N_12980);
nand U21483 (N_21483,N_14818,N_16659);
and U21484 (N_21484,N_17205,N_12972);
nor U21485 (N_21485,N_15276,N_14944);
nor U21486 (N_21486,N_14145,N_17909);
nor U21487 (N_21487,N_16194,N_17654);
xnor U21488 (N_21488,N_17167,N_12933);
or U21489 (N_21489,N_15278,N_16402);
or U21490 (N_21490,N_14162,N_13444);
nor U21491 (N_21491,N_13270,N_15573);
nand U21492 (N_21492,N_16955,N_14007);
nor U21493 (N_21493,N_12632,N_13767);
or U21494 (N_21494,N_12446,N_12069);
xnor U21495 (N_21495,N_16333,N_16408);
nand U21496 (N_21496,N_15680,N_17634);
xnor U21497 (N_21497,N_12725,N_17515);
xnor U21498 (N_21498,N_13363,N_15546);
or U21499 (N_21499,N_16561,N_12746);
nand U21500 (N_21500,N_16666,N_13756);
xor U21501 (N_21501,N_13655,N_13691);
and U21502 (N_21502,N_14285,N_16535);
xor U21503 (N_21503,N_12573,N_15367);
or U21504 (N_21504,N_16719,N_14138);
nand U21505 (N_21505,N_12517,N_17269);
nand U21506 (N_21506,N_13150,N_17949);
xor U21507 (N_21507,N_16280,N_17166);
nor U21508 (N_21508,N_13181,N_13306);
nor U21509 (N_21509,N_14224,N_16504);
or U21510 (N_21510,N_13268,N_15626);
or U21511 (N_21511,N_12583,N_13954);
and U21512 (N_21512,N_13777,N_14193);
or U21513 (N_21513,N_13158,N_12039);
nand U21514 (N_21514,N_13193,N_16676);
or U21515 (N_21515,N_14318,N_15533);
or U21516 (N_21516,N_17848,N_15632);
nand U21517 (N_21517,N_13360,N_15276);
and U21518 (N_21518,N_16601,N_14798);
and U21519 (N_21519,N_14896,N_16975);
nor U21520 (N_21520,N_17766,N_17152);
nand U21521 (N_21521,N_14112,N_12019);
nor U21522 (N_21522,N_17969,N_12936);
xnor U21523 (N_21523,N_13811,N_16091);
nor U21524 (N_21524,N_16294,N_16530);
or U21525 (N_21525,N_16941,N_14052);
or U21526 (N_21526,N_17794,N_13434);
nand U21527 (N_21527,N_16940,N_13251);
and U21528 (N_21528,N_12278,N_12852);
and U21529 (N_21529,N_16285,N_13822);
or U21530 (N_21530,N_15011,N_15936);
nor U21531 (N_21531,N_16945,N_16294);
xor U21532 (N_21532,N_17506,N_15016);
nor U21533 (N_21533,N_12415,N_14117);
and U21534 (N_21534,N_14061,N_17422);
xnor U21535 (N_21535,N_13581,N_15146);
xor U21536 (N_21536,N_13377,N_16395);
and U21537 (N_21537,N_17311,N_15951);
nor U21538 (N_21538,N_16925,N_12528);
xor U21539 (N_21539,N_16393,N_12907);
and U21540 (N_21540,N_12163,N_12934);
or U21541 (N_21541,N_15461,N_16039);
xnor U21542 (N_21542,N_17729,N_12431);
xor U21543 (N_21543,N_14312,N_16673);
xor U21544 (N_21544,N_15624,N_12716);
or U21545 (N_21545,N_15319,N_15684);
nand U21546 (N_21546,N_16372,N_12412);
and U21547 (N_21547,N_13633,N_17861);
or U21548 (N_21548,N_16472,N_16212);
or U21549 (N_21549,N_13013,N_17044);
nand U21550 (N_21550,N_12026,N_13875);
nor U21551 (N_21551,N_15957,N_15833);
or U21552 (N_21552,N_14927,N_13015);
and U21553 (N_21553,N_13671,N_15384);
xnor U21554 (N_21554,N_13546,N_17887);
or U21555 (N_21555,N_17091,N_17311);
xor U21556 (N_21556,N_15925,N_15578);
xnor U21557 (N_21557,N_13360,N_12205);
and U21558 (N_21558,N_14446,N_15076);
and U21559 (N_21559,N_14031,N_14470);
xor U21560 (N_21560,N_12742,N_12911);
xor U21561 (N_21561,N_15199,N_15163);
nand U21562 (N_21562,N_14867,N_16509);
or U21563 (N_21563,N_13948,N_12769);
and U21564 (N_21564,N_12574,N_17508);
nand U21565 (N_21565,N_17970,N_14941);
nand U21566 (N_21566,N_13485,N_12119);
or U21567 (N_21567,N_13128,N_12678);
nand U21568 (N_21568,N_16100,N_15027);
or U21569 (N_21569,N_14271,N_12117);
xnor U21570 (N_21570,N_12510,N_14352);
xnor U21571 (N_21571,N_17504,N_15440);
or U21572 (N_21572,N_13358,N_17595);
nor U21573 (N_21573,N_14457,N_17290);
and U21574 (N_21574,N_17171,N_14782);
xor U21575 (N_21575,N_14633,N_13423);
nor U21576 (N_21576,N_17007,N_13112);
xor U21577 (N_21577,N_14338,N_15876);
or U21578 (N_21578,N_14623,N_13038);
or U21579 (N_21579,N_17807,N_15443);
or U21580 (N_21580,N_13166,N_13121);
or U21581 (N_21581,N_14870,N_14085);
and U21582 (N_21582,N_17233,N_16133);
and U21583 (N_21583,N_16266,N_14125);
xnor U21584 (N_21584,N_13092,N_15286);
and U21585 (N_21585,N_16238,N_12950);
and U21586 (N_21586,N_12143,N_16683);
xnor U21587 (N_21587,N_13612,N_14836);
nand U21588 (N_21588,N_15485,N_15824);
or U21589 (N_21589,N_14560,N_16536);
nand U21590 (N_21590,N_16504,N_15764);
nand U21591 (N_21591,N_13807,N_14527);
or U21592 (N_21592,N_12305,N_16888);
xnor U21593 (N_21593,N_14599,N_12782);
nor U21594 (N_21594,N_13194,N_17850);
or U21595 (N_21595,N_16527,N_14236);
and U21596 (N_21596,N_13807,N_13006);
and U21597 (N_21597,N_16224,N_15913);
and U21598 (N_21598,N_17373,N_14558);
or U21599 (N_21599,N_12753,N_16874);
and U21600 (N_21600,N_16714,N_13103);
xnor U21601 (N_21601,N_16604,N_15276);
and U21602 (N_21602,N_13145,N_12848);
nand U21603 (N_21603,N_14892,N_15898);
nand U21604 (N_21604,N_12862,N_13239);
or U21605 (N_21605,N_15681,N_15495);
or U21606 (N_21606,N_12327,N_12552);
nand U21607 (N_21607,N_17746,N_14752);
and U21608 (N_21608,N_15534,N_17974);
xnor U21609 (N_21609,N_12210,N_12486);
or U21610 (N_21610,N_16571,N_13533);
xnor U21611 (N_21611,N_16636,N_13030);
and U21612 (N_21612,N_17140,N_15631);
nand U21613 (N_21613,N_13014,N_16087);
or U21614 (N_21614,N_15065,N_14515);
nand U21615 (N_21615,N_13325,N_15102);
nor U21616 (N_21616,N_14524,N_13984);
nand U21617 (N_21617,N_13581,N_13911);
xor U21618 (N_21618,N_14116,N_15424);
or U21619 (N_21619,N_15152,N_17649);
xor U21620 (N_21620,N_14406,N_12531);
and U21621 (N_21621,N_15876,N_16969);
nor U21622 (N_21622,N_14797,N_16649);
and U21623 (N_21623,N_17185,N_15863);
nand U21624 (N_21624,N_15922,N_15318);
nor U21625 (N_21625,N_15423,N_12564);
nand U21626 (N_21626,N_14011,N_13777);
or U21627 (N_21627,N_14406,N_12454);
nand U21628 (N_21628,N_13489,N_15169);
nor U21629 (N_21629,N_17546,N_12028);
nand U21630 (N_21630,N_12902,N_15784);
nor U21631 (N_21631,N_16312,N_12648);
nand U21632 (N_21632,N_15089,N_14740);
or U21633 (N_21633,N_15698,N_12743);
or U21634 (N_21634,N_15733,N_16104);
and U21635 (N_21635,N_17131,N_12938);
xor U21636 (N_21636,N_14744,N_17707);
xor U21637 (N_21637,N_14261,N_14252);
nand U21638 (N_21638,N_15836,N_13461);
and U21639 (N_21639,N_17377,N_13826);
nand U21640 (N_21640,N_14363,N_16632);
nand U21641 (N_21641,N_17501,N_15306);
nor U21642 (N_21642,N_15383,N_13456);
xor U21643 (N_21643,N_15415,N_12455);
or U21644 (N_21644,N_15391,N_15131);
nand U21645 (N_21645,N_13810,N_13076);
nand U21646 (N_21646,N_16390,N_15137);
nand U21647 (N_21647,N_12402,N_13591);
nor U21648 (N_21648,N_16591,N_16661);
and U21649 (N_21649,N_13490,N_17960);
nand U21650 (N_21650,N_13593,N_13866);
and U21651 (N_21651,N_15245,N_15524);
xor U21652 (N_21652,N_14714,N_14485);
xnor U21653 (N_21653,N_16672,N_12283);
xor U21654 (N_21654,N_15315,N_16695);
nor U21655 (N_21655,N_14936,N_17794);
nor U21656 (N_21656,N_13458,N_17803);
nand U21657 (N_21657,N_14874,N_14502);
nor U21658 (N_21658,N_16861,N_13228);
and U21659 (N_21659,N_17207,N_14898);
xnor U21660 (N_21660,N_13394,N_17388);
and U21661 (N_21661,N_12326,N_12636);
or U21662 (N_21662,N_13042,N_12223);
xor U21663 (N_21663,N_15317,N_13050);
nand U21664 (N_21664,N_12140,N_13038);
or U21665 (N_21665,N_15814,N_15816);
nor U21666 (N_21666,N_16653,N_17971);
nand U21667 (N_21667,N_14132,N_12730);
xor U21668 (N_21668,N_14732,N_16096);
and U21669 (N_21669,N_12034,N_12591);
nor U21670 (N_21670,N_12147,N_13836);
or U21671 (N_21671,N_13198,N_14834);
and U21672 (N_21672,N_12655,N_14813);
and U21673 (N_21673,N_13174,N_16792);
nor U21674 (N_21674,N_12604,N_16425);
xor U21675 (N_21675,N_16011,N_16083);
nor U21676 (N_21676,N_14150,N_17295);
or U21677 (N_21677,N_14925,N_14126);
and U21678 (N_21678,N_16072,N_16947);
nand U21679 (N_21679,N_14659,N_12123);
nor U21680 (N_21680,N_14820,N_13999);
xnor U21681 (N_21681,N_15263,N_16057);
or U21682 (N_21682,N_13221,N_13839);
nor U21683 (N_21683,N_16725,N_16833);
xor U21684 (N_21684,N_12550,N_14906);
nor U21685 (N_21685,N_16850,N_15704);
nand U21686 (N_21686,N_16398,N_15580);
xor U21687 (N_21687,N_14259,N_16673);
xnor U21688 (N_21688,N_14915,N_14291);
or U21689 (N_21689,N_16624,N_14395);
xnor U21690 (N_21690,N_12763,N_13059);
xor U21691 (N_21691,N_13107,N_12970);
or U21692 (N_21692,N_12385,N_13261);
xnor U21693 (N_21693,N_13762,N_17190);
xnor U21694 (N_21694,N_13307,N_13584);
nor U21695 (N_21695,N_16357,N_13873);
and U21696 (N_21696,N_16628,N_14176);
and U21697 (N_21697,N_14920,N_16452);
and U21698 (N_21698,N_12374,N_13376);
nand U21699 (N_21699,N_14673,N_15216);
nor U21700 (N_21700,N_17259,N_17422);
nand U21701 (N_21701,N_12221,N_16925);
and U21702 (N_21702,N_15832,N_15825);
and U21703 (N_21703,N_17886,N_15946);
and U21704 (N_21704,N_12573,N_13911);
nor U21705 (N_21705,N_16188,N_15993);
nand U21706 (N_21706,N_13520,N_12701);
nand U21707 (N_21707,N_13500,N_13343);
nand U21708 (N_21708,N_14312,N_15306);
xor U21709 (N_21709,N_12949,N_14051);
nand U21710 (N_21710,N_14795,N_12335);
xor U21711 (N_21711,N_13326,N_12736);
or U21712 (N_21712,N_13125,N_16304);
nand U21713 (N_21713,N_14036,N_16966);
nor U21714 (N_21714,N_16097,N_12483);
nand U21715 (N_21715,N_14603,N_13487);
xor U21716 (N_21716,N_16529,N_13959);
and U21717 (N_21717,N_16687,N_17180);
nor U21718 (N_21718,N_15574,N_13191);
xor U21719 (N_21719,N_16501,N_14296);
nor U21720 (N_21720,N_14786,N_16643);
and U21721 (N_21721,N_17826,N_13012);
and U21722 (N_21722,N_17851,N_12302);
xnor U21723 (N_21723,N_17354,N_16588);
nor U21724 (N_21724,N_15664,N_12499);
nor U21725 (N_21725,N_17761,N_14685);
and U21726 (N_21726,N_16679,N_16519);
nand U21727 (N_21727,N_13232,N_16628);
or U21728 (N_21728,N_14405,N_13179);
nand U21729 (N_21729,N_14914,N_12644);
or U21730 (N_21730,N_16647,N_15677);
or U21731 (N_21731,N_14298,N_12688);
nand U21732 (N_21732,N_15793,N_17311);
or U21733 (N_21733,N_14269,N_15725);
and U21734 (N_21734,N_17913,N_15399);
nand U21735 (N_21735,N_16903,N_16990);
nand U21736 (N_21736,N_13258,N_17030);
and U21737 (N_21737,N_17635,N_14036);
or U21738 (N_21738,N_15406,N_14167);
nand U21739 (N_21739,N_16876,N_12494);
and U21740 (N_21740,N_17209,N_17972);
xor U21741 (N_21741,N_12009,N_14483);
nand U21742 (N_21742,N_12776,N_15188);
nand U21743 (N_21743,N_14862,N_13081);
and U21744 (N_21744,N_17026,N_17311);
nand U21745 (N_21745,N_15313,N_13074);
xnor U21746 (N_21746,N_16617,N_13122);
nor U21747 (N_21747,N_12988,N_14884);
nand U21748 (N_21748,N_16423,N_14443);
nor U21749 (N_21749,N_15272,N_16688);
nor U21750 (N_21750,N_16444,N_15802);
xnor U21751 (N_21751,N_15426,N_15307);
xnor U21752 (N_21752,N_13652,N_12352);
nor U21753 (N_21753,N_15044,N_15884);
nor U21754 (N_21754,N_16884,N_13970);
or U21755 (N_21755,N_13962,N_13240);
xor U21756 (N_21756,N_16269,N_15349);
nor U21757 (N_21757,N_15258,N_16319);
nor U21758 (N_21758,N_15038,N_14937);
or U21759 (N_21759,N_12776,N_12391);
or U21760 (N_21760,N_17611,N_16748);
or U21761 (N_21761,N_17819,N_12803);
or U21762 (N_21762,N_17239,N_12490);
nor U21763 (N_21763,N_16912,N_15223);
nor U21764 (N_21764,N_12764,N_15212);
xor U21765 (N_21765,N_14932,N_14872);
or U21766 (N_21766,N_13755,N_12222);
or U21767 (N_21767,N_16600,N_17812);
and U21768 (N_21768,N_17315,N_16988);
or U21769 (N_21769,N_14903,N_14361);
nor U21770 (N_21770,N_14867,N_16833);
and U21771 (N_21771,N_16510,N_15604);
and U21772 (N_21772,N_14354,N_16416);
nor U21773 (N_21773,N_17870,N_12979);
or U21774 (N_21774,N_17157,N_14123);
xnor U21775 (N_21775,N_12571,N_12064);
xor U21776 (N_21776,N_12533,N_17490);
xor U21777 (N_21777,N_16023,N_17902);
or U21778 (N_21778,N_13633,N_17487);
nand U21779 (N_21779,N_12116,N_13680);
xnor U21780 (N_21780,N_16477,N_13326);
nand U21781 (N_21781,N_12979,N_14695);
xnor U21782 (N_21782,N_16830,N_17857);
xnor U21783 (N_21783,N_14360,N_16413);
nor U21784 (N_21784,N_12387,N_17792);
and U21785 (N_21785,N_15722,N_14867);
nand U21786 (N_21786,N_17119,N_15761);
nand U21787 (N_21787,N_14582,N_13730);
nand U21788 (N_21788,N_12326,N_17221);
and U21789 (N_21789,N_13659,N_14183);
xnor U21790 (N_21790,N_17034,N_17525);
or U21791 (N_21791,N_15571,N_17067);
xor U21792 (N_21792,N_13821,N_17581);
and U21793 (N_21793,N_17963,N_13863);
or U21794 (N_21794,N_12239,N_14404);
xnor U21795 (N_21795,N_13524,N_12950);
nor U21796 (N_21796,N_16315,N_17566);
or U21797 (N_21797,N_17283,N_17069);
nor U21798 (N_21798,N_16185,N_16449);
xor U21799 (N_21799,N_17343,N_15958);
xnor U21800 (N_21800,N_17119,N_14855);
nor U21801 (N_21801,N_14800,N_17337);
or U21802 (N_21802,N_13180,N_13335);
or U21803 (N_21803,N_15349,N_17248);
or U21804 (N_21804,N_12981,N_16599);
and U21805 (N_21805,N_15258,N_12822);
nor U21806 (N_21806,N_14056,N_17972);
nand U21807 (N_21807,N_15002,N_17736);
or U21808 (N_21808,N_14937,N_13054);
or U21809 (N_21809,N_14163,N_14545);
xnor U21810 (N_21810,N_17844,N_13190);
nor U21811 (N_21811,N_17673,N_17754);
nand U21812 (N_21812,N_16504,N_15433);
nand U21813 (N_21813,N_12593,N_16282);
and U21814 (N_21814,N_14730,N_14519);
nand U21815 (N_21815,N_17541,N_17594);
or U21816 (N_21816,N_12669,N_14794);
xnor U21817 (N_21817,N_17493,N_15410);
nand U21818 (N_21818,N_17924,N_15330);
xor U21819 (N_21819,N_16544,N_13589);
xnor U21820 (N_21820,N_17138,N_12228);
xor U21821 (N_21821,N_17484,N_13870);
and U21822 (N_21822,N_12688,N_12148);
nand U21823 (N_21823,N_15519,N_16725);
or U21824 (N_21824,N_13910,N_17366);
nand U21825 (N_21825,N_17868,N_16218);
and U21826 (N_21826,N_16751,N_16621);
nor U21827 (N_21827,N_12265,N_13450);
nor U21828 (N_21828,N_12103,N_15345);
nand U21829 (N_21829,N_14291,N_12908);
and U21830 (N_21830,N_16201,N_14521);
or U21831 (N_21831,N_16977,N_12627);
and U21832 (N_21832,N_15903,N_16902);
xnor U21833 (N_21833,N_16029,N_16375);
nor U21834 (N_21834,N_16674,N_14486);
or U21835 (N_21835,N_15184,N_13077);
or U21836 (N_21836,N_14255,N_15019);
nand U21837 (N_21837,N_16925,N_15314);
nand U21838 (N_21838,N_13844,N_13182);
and U21839 (N_21839,N_12053,N_17143);
nand U21840 (N_21840,N_13957,N_14553);
and U21841 (N_21841,N_12007,N_15874);
xor U21842 (N_21842,N_15955,N_14472);
and U21843 (N_21843,N_13160,N_13213);
nor U21844 (N_21844,N_13357,N_14822);
and U21845 (N_21845,N_14977,N_13333);
xor U21846 (N_21846,N_17148,N_13302);
nand U21847 (N_21847,N_17775,N_17291);
nand U21848 (N_21848,N_13195,N_15638);
nor U21849 (N_21849,N_15970,N_14239);
xnor U21850 (N_21850,N_17594,N_15836);
nor U21851 (N_21851,N_15441,N_17090);
or U21852 (N_21852,N_15913,N_15646);
or U21853 (N_21853,N_13489,N_13091);
or U21854 (N_21854,N_15105,N_16441);
nand U21855 (N_21855,N_15373,N_12416);
nand U21856 (N_21856,N_12433,N_12145);
or U21857 (N_21857,N_13228,N_17222);
xnor U21858 (N_21858,N_14769,N_16211);
or U21859 (N_21859,N_12092,N_15497);
nor U21860 (N_21860,N_16713,N_16351);
nor U21861 (N_21861,N_16603,N_13040);
and U21862 (N_21862,N_16257,N_15520);
and U21863 (N_21863,N_16873,N_14663);
nand U21864 (N_21864,N_15339,N_16985);
and U21865 (N_21865,N_15246,N_13525);
nor U21866 (N_21866,N_17478,N_17757);
and U21867 (N_21867,N_14625,N_17431);
or U21868 (N_21868,N_17538,N_17194);
nor U21869 (N_21869,N_13884,N_17279);
xor U21870 (N_21870,N_12007,N_15544);
and U21871 (N_21871,N_13202,N_17431);
nor U21872 (N_21872,N_14053,N_12097);
and U21873 (N_21873,N_13932,N_16485);
nand U21874 (N_21874,N_12161,N_17239);
nand U21875 (N_21875,N_15825,N_16480);
or U21876 (N_21876,N_15250,N_14742);
and U21877 (N_21877,N_12534,N_15408);
nor U21878 (N_21878,N_17528,N_17753);
and U21879 (N_21879,N_16512,N_13602);
and U21880 (N_21880,N_12487,N_12464);
nor U21881 (N_21881,N_17900,N_17795);
nor U21882 (N_21882,N_17577,N_15427);
nand U21883 (N_21883,N_14249,N_15757);
and U21884 (N_21884,N_16581,N_14045);
and U21885 (N_21885,N_15221,N_16708);
nand U21886 (N_21886,N_15393,N_14591);
nand U21887 (N_21887,N_12321,N_15266);
xor U21888 (N_21888,N_16646,N_13005);
xor U21889 (N_21889,N_14308,N_12302);
and U21890 (N_21890,N_17758,N_12663);
or U21891 (N_21891,N_13246,N_13859);
or U21892 (N_21892,N_17094,N_13098);
and U21893 (N_21893,N_12997,N_16962);
nor U21894 (N_21894,N_15346,N_16033);
and U21895 (N_21895,N_14310,N_12633);
nand U21896 (N_21896,N_14870,N_12774);
and U21897 (N_21897,N_14417,N_16665);
nor U21898 (N_21898,N_14486,N_16936);
xor U21899 (N_21899,N_14148,N_15491);
and U21900 (N_21900,N_15862,N_17200);
nand U21901 (N_21901,N_16632,N_15223);
xor U21902 (N_21902,N_16024,N_12527);
and U21903 (N_21903,N_14367,N_17618);
and U21904 (N_21904,N_17685,N_14669);
nand U21905 (N_21905,N_12235,N_13814);
or U21906 (N_21906,N_17082,N_15047);
nor U21907 (N_21907,N_12038,N_16158);
xnor U21908 (N_21908,N_12200,N_14950);
xor U21909 (N_21909,N_16000,N_12044);
nand U21910 (N_21910,N_15240,N_14778);
nor U21911 (N_21911,N_16891,N_17505);
or U21912 (N_21912,N_14352,N_14392);
nor U21913 (N_21913,N_17464,N_16177);
or U21914 (N_21914,N_14555,N_17483);
nand U21915 (N_21915,N_12599,N_15425);
nand U21916 (N_21916,N_17762,N_17496);
nand U21917 (N_21917,N_14370,N_17990);
xor U21918 (N_21918,N_17571,N_14619);
nand U21919 (N_21919,N_17417,N_12169);
and U21920 (N_21920,N_12982,N_14289);
nor U21921 (N_21921,N_17524,N_14465);
xor U21922 (N_21922,N_15150,N_16644);
and U21923 (N_21923,N_12372,N_12629);
nand U21924 (N_21924,N_14734,N_15715);
nand U21925 (N_21925,N_13270,N_14996);
nand U21926 (N_21926,N_13701,N_13138);
nand U21927 (N_21927,N_12543,N_14828);
and U21928 (N_21928,N_12939,N_14655);
xnor U21929 (N_21929,N_14208,N_12919);
and U21930 (N_21930,N_17227,N_12287);
nand U21931 (N_21931,N_16609,N_16385);
nor U21932 (N_21932,N_13053,N_13557);
xor U21933 (N_21933,N_14686,N_16474);
and U21934 (N_21934,N_15963,N_14515);
and U21935 (N_21935,N_13934,N_17511);
and U21936 (N_21936,N_17898,N_16553);
nand U21937 (N_21937,N_17618,N_17947);
xnor U21938 (N_21938,N_15340,N_17728);
and U21939 (N_21939,N_14003,N_16368);
or U21940 (N_21940,N_17381,N_13476);
and U21941 (N_21941,N_15718,N_12095);
and U21942 (N_21942,N_16552,N_14601);
and U21943 (N_21943,N_13931,N_12763);
xnor U21944 (N_21944,N_16176,N_15090);
and U21945 (N_21945,N_15084,N_17619);
and U21946 (N_21946,N_17534,N_12130);
xnor U21947 (N_21947,N_12690,N_16545);
xor U21948 (N_21948,N_16747,N_16169);
or U21949 (N_21949,N_14106,N_15667);
and U21950 (N_21950,N_12283,N_15712);
or U21951 (N_21951,N_17871,N_17647);
and U21952 (N_21952,N_17658,N_15947);
nand U21953 (N_21953,N_13245,N_15339);
or U21954 (N_21954,N_16507,N_13979);
or U21955 (N_21955,N_14831,N_13476);
and U21956 (N_21956,N_16478,N_16443);
xor U21957 (N_21957,N_17685,N_13957);
nand U21958 (N_21958,N_12285,N_14584);
nor U21959 (N_21959,N_16267,N_12307);
xor U21960 (N_21960,N_16677,N_17619);
and U21961 (N_21961,N_14071,N_13403);
nand U21962 (N_21962,N_16939,N_14461);
nand U21963 (N_21963,N_16979,N_17361);
nand U21964 (N_21964,N_13112,N_16273);
xor U21965 (N_21965,N_14276,N_15148);
nand U21966 (N_21966,N_16257,N_15119);
nor U21967 (N_21967,N_13241,N_12583);
xor U21968 (N_21968,N_14164,N_16206);
nand U21969 (N_21969,N_15397,N_15937);
xor U21970 (N_21970,N_12771,N_14547);
nor U21971 (N_21971,N_17759,N_13023);
nor U21972 (N_21972,N_16239,N_13794);
or U21973 (N_21973,N_17813,N_16485);
and U21974 (N_21974,N_14796,N_12268);
nor U21975 (N_21975,N_12835,N_17362);
xor U21976 (N_21976,N_17037,N_15511);
or U21977 (N_21977,N_13412,N_15782);
or U21978 (N_21978,N_12318,N_17336);
xor U21979 (N_21979,N_17813,N_12636);
or U21980 (N_21980,N_17794,N_13562);
and U21981 (N_21981,N_13081,N_17635);
and U21982 (N_21982,N_12234,N_12177);
and U21983 (N_21983,N_17016,N_12741);
or U21984 (N_21984,N_17829,N_15866);
nand U21985 (N_21985,N_12316,N_16554);
or U21986 (N_21986,N_16599,N_15167);
nor U21987 (N_21987,N_13034,N_16100);
nand U21988 (N_21988,N_12483,N_16032);
nor U21989 (N_21989,N_17077,N_14364);
nor U21990 (N_21990,N_16062,N_17738);
xor U21991 (N_21991,N_15539,N_17655);
or U21992 (N_21992,N_13936,N_12371);
xor U21993 (N_21993,N_15721,N_15987);
nor U21994 (N_21994,N_12081,N_14560);
nand U21995 (N_21995,N_14251,N_15480);
nand U21996 (N_21996,N_15691,N_16047);
nand U21997 (N_21997,N_16767,N_14529);
or U21998 (N_21998,N_14498,N_16413);
xor U21999 (N_21999,N_12087,N_16983);
or U22000 (N_22000,N_12812,N_13260);
nand U22001 (N_22001,N_12370,N_13682);
nand U22002 (N_22002,N_16423,N_17483);
or U22003 (N_22003,N_12899,N_15306);
nand U22004 (N_22004,N_17330,N_15076);
or U22005 (N_22005,N_17671,N_15735);
nor U22006 (N_22006,N_17600,N_14920);
nand U22007 (N_22007,N_16117,N_15172);
xor U22008 (N_22008,N_13538,N_15417);
xor U22009 (N_22009,N_16980,N_12856);
xnor U22010 (N_22010,N_15887,N_12583);
nand U22011 (N_22011,N_17043,N_12133);
xnor U22012 (N_22012,N_15544,N_12343);
or U22013 (N_22013,N_15938,N_15322);
xor U22014 (N_22014,N_16635,N_16439);
nor U22015 (N_22015,N_14326,N_16225);
or U22016 (N_22016,N_15417,N_17830);
and U22017 (N_22017,N_16028,N_17750);
nand U22018 (N_22018,N_15006,N_17313);
or U22019 (N_22019,N_12696,N_12369);
nand U22020 (N_22020,N_13964,N_14252);
nand U22021 (N_22021,N_15344,N_12760);
nand U22022 (N_22022,N_14496,N_16903);
and U22023 (N_22023,N_15449,N_13739);
xnor U22024 (N_22024,N_12955,N_12128);
and U22025 (N_22025,N_16104,N_17847);
xnor U22026 (N_22026,N_13356,N_14631);
or U22027 (N_22027,N_13839,N_17776);
xor U22028 (N_22028,N_14064,N_17793);
nor U22029 (N_22029,N_13676,N_13863);
or U22030 (N_22030,N_13538,N_17640);
or U22031 (N_22031,N_17044,N_17994);
xor U22032 (N_22032,N_12908,N_13758);
xnor U22033 (N_22033,N_12571,N_17896);
nand U22034 (N_22034,N_12016,N_15912);
or U22035 (N_22035,N_15335,N_17623);
and U22036 (N_22036,N_17704,N_14459);
or U22037 (N_22037,N_13988,N_14707);
and U22038 (N_22038,N_15529,N_14294);
nor U22039 (N_22039,N_14188,N_13442);
nand U22040 (N_22040,N_14240,N_12670);
or U22041 (N_22041,N_13715,N_14435);
xor U22042 (N_22042,N_13937,N_17554);
nand U22043 (N_22043,N_16211,N_15587);
nor U22044 (N_22044,N_12797,N_15889);
and U22045 (N_22045,N_15738,N_13651);
or U22046 (N_22046,N_12565,N_12435);
nor U22047 (N_22047,N_15604,N_12081);
xnor U22048 (N_22048,N_17640,N_17587);
xor U22049 (N_22049,N_17599,N_12139);
or U22050 (N_22050,N_16606,N_15795);
xnor U22051 (N_22051,N_14013,N_12250);
or U22052 (N_22052,N_15317,N_15139);
xnor U22053 (N_22053,N_14496,N_12170);
nand U22054 (N_22054,N_12187,N_14042);
xor U22055 (N_22055,N_15135,N_14492);
nand U22056 (N_22056,N_13789,N_16568);
nand U22057 (N_22057,N_13551,N_14206);
or U22058 (N_22058,N_17042,N_16447);
nor U22059 (N_22059,N_12324,N_14838);
nand U22060 (N_22060,N_16149,N_15521);
or U22061 (N_22061,N_12638,N_15144);
or U22062 (N_22062,N_15808,N_17613);
nor U22063 (N_22063,N_13586,N_15800);
or U22064 (N_22064,N_17366,N_13311);
nor U22065 (N_22065,N_15564,N_13864);
xor U22066 (N_22066,N_15550,N_17867);
and U22067 (N_22067,N_15825,N_16338);
nand U22068 (N_22068,N_14032,N_14511);
nor U22069 (N_22069,N_12720,N_15693);
nor U22070 (N_22070,N_16342,N_14375);
or U22071 (N_22071,N_17873,N_16407);
nor U22072 (N_22072,N_16973,N_12582);
nor U22073 (N_22073,N_13429,N_15565);
or U22074 (N_22074,N_15046,N_16459);
and U22075 (N_22075,N_15511,N_17369);
and U22076 (N_22076,N_16680,N_13018);
nor U22077 (N_22077,N_14137,N_15159);
and U22078 (N_22078,N_13787,N_12845);
nand U22079 (N_22079,N_12691,N_13587);
or U22080 (N_22080,N_17805,N_15288);
nand U22081 (N_22081,N_15663,N_12503);
and U22082 (N_22082,N_16180,N_14012);
and U22083 (N_22083,N_14939,N_15439);
xnor U22084 (N_22084,N_17212,N_15321);
or U22085 (N_22085,N_13181,N_15656);
nor U22086 (N_22086,N_17726,N_15089);
nand U22087 (N_22087,N_16093,N_13844);
xnor U22088 (N_22088,N_12296,N_15397);
nand U22089 (N_22089,N_17075,N_16624);
nand U22090 (N_22090,N_13562,N_13513);
or U22091 (N_22091,N_12612,N_17802);
or U22092 (N_22092,N_15431,N_16536);
and U22093 (N_22093,N_16559,N_13735);
nand U22094 (N_22094,N_16718,N_13382);
nor U22095 (N_22095,N_14111,N_15620);
xor U22096 (N_22096,N_13603,N_17173);
and U22097 (N_22097,N_13489,N_13591);
and U22098 (N_22098,N_14483,N_15247);
and U22099 (N_22099,N_12799,N_15950);
nor U22100 (N_22100,N_14087,N_13596);
or U22101 (N_22101,N_13423,N_15359);
nor U22102 (N_22102,N_16126,N_12363);
nor U22103 (N_22103,N_14181,N_16227);
or U22104 (N_22104,N_17475,N_14871);
and U22105 (N_22105,N_14786,N_14506);
nor U22106 (N_22106,N_16082,N_15137);
xor U22107 (N_22107,N_14984,N_13922);
and U22108 (N_22108,N_15519,N_13259);
nand U22109 (N_22109,N_16969,N_17791);
and U22110 (N_22110,N_16897,N_16332);
xnor U22111 (N_22111,N_14107,N_13792);
xor U22112 (N_22112,N_13731,N_12170);
nand U22113 (N_22113,N_17250,N_12590);
nor U22114 (N_22114,N_17980,N_14331);
or U22115 (N_22115,N_17210,N_15837);
or U22116 (N_22116,N_14875,N_16487);
xnor U22117 (N_22117,N_14659,N_12584);
and U22118 (N_22118,N_16129,N_16518);
nor U22119 (N_22119,N_17951,N_12907);
or U22120 (N_22120,N_15444,N_17535);
and U22121 (N_22121,N_14469,N_15105);
and U22122 (N_22122,N_16581,N_17511);
nor U22123 (N_22123,N_13076,N_15517);
xnor U22124 (N_22124,N_15404,N_15635);
nand U22125 (N_22125,N_17905,N_15950);
nand U22126 (N_22126,N_17060,N_17166);
or U22127 (N_22127,N_16484,N_13800);
xor U22128 (N_22128,N_14094,N_12037);
and U22129 (N_22129,N_17987,N_17633);
xnor U22130 (N_22130,N_12406,N_12194);
nand U22131 (N_22131,N_14584,N_12626);
or U22132 (N_22132,N_15107,N_15032);
and U22133 (N_22133,N_17443,N_15404);
or U22134 (N_22134,N_17641,N_13404);
or U22135 (N_22135,N_16810,N_17815);
nand U22136 (N_22136,N_15925,N_14154);
nand U22137 (N_22137,N_15075,N_15955);
xor U22138 (N_22138,N_13860,N_14632);
xor U22139 (N_22139,N_14416,N_17650);
nand U22140 (N_22140,N_13862,N_14472);
nor U22141 (N_22141,N_12716,N_17700);
and U22142 (N_22142,N_17321,N_15215);
nor U22143 (N_22143,N_13831,N_15415);
nor U22144 (N_22144,N_15094,N_15638);
xor U22145 (N_22145,N_17066,N_14503);
or U22146 (N_22146,N_16747,N_14105);
nand U22147 (N_22147,N_14470,N_13724);
or U22148 (N_22148,N_12781,N_14300);
nand U22149 (N_22149,N_13357,N_14766);
xnor U22150 (N_22150,N_16311,N_12521);
nand U22151 (N_22151,N_12557,N_13389);
or U22152 (N_22152,N_13666,N_13553);
nor U22153 (N_22153,N_13143,N_13377);
nor U22154 (N_22154,N_15760,N_15621);
nand U22155 (N_22155,N_12031,N_15240);
xor U22156 (N_22156,N_14187,N_14099);
nand U22157 (N_22157,N_12921,N_12155);
nor U22158 (N_22158,N_12167,N_15839);
or U22159 (N_22159,N_17556,N_12602);
xor U22160 (N_22160,N_15337,N_14510);
nor U22161 (N_22161,N_14286,N_15168);
nor U22162 (N_22162,N_12966,N_15769);
nand U22163 (N_22163,N_15960,N_17478);
or U22164 (N_22164,N_15634,N_16678);
and U22165 (N_22165,N_15696,N_15249);
and U22166 (N_22166,N_12405,N_14649);
nand U22167 (N_22167,N_14849,N_13342);
nand U22168 (N_22168,N_17403,N_15763);
nor U22169 (N_22169,N_16858,N_15186);
xnor U22170 (N_22170,N_16825,N_16026);
nor U22171 (N_22171,N_13199,N_14240);
and U22172 (N_22172,N_14635,N_13576);
or U22173 (N_22173,N_13162,N_14913);
nand U22174 (N_22174,N_12324,N_14586);
nand U22175 (N_22175,N_17389,N_14407);
and U22176 (N_22176,N_12432,N_12608);
and U22177 (N_22177,N_12749,N_12150);
and U22178 (N_22178,N_13603,N_15813);
xnor U22179 (N_22179,N_12195,N_14214);
or U22180 (N_22180,N_13705,N_16153);
nand U22181 (N_22181,N_16466,N_13546);
nor U22182 (N_22182,N_14290,N_16744);
nor U22183 (N_22183,N_14830,N_17727);
nand U22184 (N_22184,N_17343,N_15137);
nor U22185 (N_22185,N_13626,N_14136);
nor U22186 (N_22186,N_15401,N_12441);
and U22187 (N_22187,N_15714,N_13398);
nand U22188 (N_22188,N_17140,N_16590);
and U22189 (N_22189,N_16507,N_17152);
nor U22190 (N_22190,N_15610,N_16757);
and U22191 (N_22191,N_14762,N_17103);
nand U22192 (N_22192,N_15949,N_16336);
nor U22193 (N_22193,N_16928,N_15764);
nand U22194 (N_22194,N_14952,N_17885);
and U22195 (N_22195,N_17076,N_17613);
nor U22196 (N_22196,N_17833,N_15124);
xnor U22197 (N_22197,N_15205,N_14431);
xor U22198 (N_22198,N_13849,N_14772);
nor U22199 (N_22199,N_14811,N_14017);
nand U22200 (N_22200,N_17238,N_17096);
nor U22201 (N_22201,N_16067,N_12224);
and U22202 (N_22202,N_13956,N_13943);
xor U22203 (N_22203,N_17286,N_17772);
or U22204 (N_22204,N_15704,N_15453);
xor U22205 (N_22205,N_16557,N_14395);
and U22206 (N_22206,N_17255,N_16700);
nand U22207 (N_22207,N_17939,N_14182);
and U22208 (N_22208,N_13622,N_14980);
nor U22209 (N_22209,N_16533,N_16430);
or U22210 (N_22210,N_12129,N_12420);
nor U22211 (N_22211,N_14332,N_17670);
and U22212 (N_22212,N_16815,N_17252);
xor U22213 (N_22213,N_17085,N_13947);
xor U22214 (N_22214,N_14862,N_13105);
and U22215 (N_22215,N_17374,N_14754);
xor U22216 (N_22216,N_15811,N_12393);
and U22217 (N_22217,N_17175,N_14051);
xor U22218 (N_22218,N_17506,N_17890);
xnor U22219 (N_22219,N_12870,N_14305);
nor U22220 (N_22220,N_17109,N_13197);
or U22221 (N_22221,N_17240,N_17844);
and U22222 (N_22222,N_12452,N_17620);
nor U22223 (N_22223,N_17033,N_13602);
and U22224 (N_22224,N_15922,N_16698);
xor U22225 (N_22225,N_13324,N_12241);
nor U22226 (N_22226,N_12175,N_16890);
xnor U22227 (N_22227,N_16153,N_13538);
nand U22228 (N_22228,N_17156,N_16480);
xnor U22229 (N_22229,N_15849,N_12128);
xor U22230 (N_22230,N_17473,N_16573);
or U22231 (N_22231,N_15570,N_12804);
nor U22232 (N_22232,N_13880,N_13439);
and U22233 (N_22233,N_13385,N_13876);
or U22234 (N_22234,N_13139,N_12015);
and U22235 (N_22235,N_12671,N_17805);
nor U22236 (N_22236,N_17567,N_15378);
or U22237 (N_22237,N_16602,N_13008);
nor U22238 (N_22238,N_17207,N_16481);
xnor U22239 (N_22239,N_17334,N_14165);
nor U22240 (N_22240,N_14383,N_12622);
or U22241 (N_22241,N_16223,N_16700);
or U22242 (N_22242,N_12279,N_12926);
and U22243 (N_22243,N_14185,N_13800);
xor U22244 (N_22244,N_16642,N_14149);
xor U22245 (N_22245,N_15395,N_16260);
and U22246 (N_22246,N_17678,N_15355);
and U22247 (N_22247,N_17691,N_12461);
nand U22248 (N_22248,N_13960,N_14100);
nand U22249 (N_22249,N_16715,N_14162);
or U22250 (N_22250,N_15553,N_13330);
or U22251 (N_22251,N_15911,N_13875);
nor U22252 (N_22252,N_15972,N_17511);
or U22253 (N_22253,N_14543,N_17423);
nor U22254 (N_22254,N_17728,N_12620);
xnor U22255 (N_22255,N_16056,N_15649);
and U22256 (N_22256,N_14887,N_15228);
xnor U22257 (N_22257,N_13508,N_13900);
and U22258 (N_22258,N_14944,N_16862);
nand U22259 (N_22259,N_15080,N_15902);
xnor U22260 (N_22260,N_17132,N_17177);
and U22261 (N_22261,N_12213,N_16804);
nor U22262 (N_22262,N_14660,N_14015);
nand U22263 (N_22263,N_16170,N_14960);
and U22264 (N_22264,N_12672,N_13994);
xor U22265 (N_22265,N_14343,N_12990);
or U22266 (N_22266,N_14990,N_15634);
or U22267 (N_22267,N_13490,N_16786);
nor U22268 (N_22268,N_14329,N_13362);
nand U22269 (N_22269,N_17576,N_13007);
nand U22270 (N_22270,N_16569,N_14019);
nand U22271 (N_22271,N_14448,N_13500);
xor U22272 (N_22272,N_14681,N_13704);
and U22273 (N_22273,N_16546,N_17002);
nand U22274 (N_22274,N_13206,N_16051);
nand U22275 (N_22275,N_17849,N_12363);
and U22276 (N_22276,N_17874,N_15585);
nor U22277 (N_22277,N_12718,N_14573);
nand U22278 (N_22278,N_17314,N_15125);
nand U22279 (N_22279,N_13116,N_15385);
and U22280 (N_22280,N_14029,N_16966);
nand U22281 (N_22281,N_14606,N_14101);
nand U22282 (N_22282,N_12644,N_12704);
xor U22283 (N_22283,N_17391,N_14260);
or U22284 (N_22284,N_13136,N_16032);
nand U22285 (N_22285,N_15372,N_12396);
nand U22286 (N_22286,N_12440,N_17981);
and U22287 (N_22287,N_16658,N_12399);
or U22288 (N_22288,N_12153,N_14967);
nor U22289 (N_22289,N_17495,N_17932);
xor U22290 (N_22290,N_17003,N_12238);
nor U22291 (N_22291,N_17652,N_16625);
xor U22292 (N_22292,N_17636,N_14983);
nor U22293 (N_22293,N_13268,N_17111);
xnor U22294 (N_22294,N_17622,N_14101);
nor U22295 (N_22295,N_16324,N_14658);
nand U22296 (N_22296,N_12535,N_12887);
nor U22297 (N_22297,N_14647,N_12077);
or U22298 (N_22298,N_12823,N_12859);
or U22299 (N_22299,N_12380,N_17790);
and U22300 (N_22300,N_13668,N_15080);
or U22301 (N_22301,N_14542,N_17403);
or U22302 (N_22302,N_17379,N_17207);
xnor U22303 (N_22303,N_13020,N_13423);
xnor U22304 (N_22304,N_15123,N_12774);
and U22305 (N_22305,N_15974,N_12913);
or U22306 (N_22306,N_17105,N_13190);
and U22307 (N_22307,N_15826,N_13169);
nor U22308 (N_22308,N_17106,N_13599);
or U22309 (N_22309,N_14216,N_13426);
nand U22310 (N_22310,N_17208,N_12764);
nand U22311 (N_22311,N_13918,N_14592);
nor U22312 (N_22312,N_14127,N_13784);
nor U22313 (N_22313,N_13264,N_16520);
and U22314 (N_22314,N_12747,N_14327);
or U22315 (N_22315,N_17161,N_13437);
or U22316 (N_22316,N_12576,N_13715);
nor U22317 (N_22317,N_16724,N_13870);
xnor U22318 (N_22318,N_15315,N_13446);
and U22319 (N_22319,N_16842,N_17825);
or U22320 (N_22320,N_12755,N_13203);
nor U22321 (N_22321,N_16554,N_15426);
nand U22322 (N_22322,N_17641,N_13289);
nand U22323 (N_22323,N_16459,N_13848);
nand U22324 (N_22324,N_16518,N_17248);
xor U22325 (N_22325,N_14491,N_14167);
nor U22326 (N_22326,N_15966,N_12862);
or U22327 (N_22327,N_16815,N_13989);
or U22328 (N_22328,N_14728,N_15796);
and U22329 (N_22329,N_14884,N_16272);
or U22330 (N_22330,N_12004,N_16257);
nand U22331 (N_22331,N_15100,N_12385);
or U22332 (N_22332,N_14328,N_13140);
or U22333 (N_22333,N_15100,N_16642);
and U22334 (N_22334,N_16374,N_14213);
nand U22335 (N_22335,N_15132,N_14092);
nand U22336 (N_22336,N_16851,N_13268);
or U22337 (N_22337,N_13311,N_17149);
nor U22338 (N_22338,N_12140,N_14100);
or U22339 (N_22339,N_16050,N_16277);
nor U22340 (N_22340,N_12944,N_16891);
xnor U22341 (N_22341,N_13712,N_12165);
xor U22342 (N_22342,N_15612,N_13039);
nor U22343 (N_22343,N_14199,N_17228);
or U22344 (N_22344,N_13620,N_15960);
nand U22345 (N_22345,N_12686,N_12013);
or U22346 (N_22346,N_17187,N_16864);
and U22347 (N_22347,N_15576,N_13594);
or U22348 (N_22348,N_17180,N_13621);
xor U22349 (N_22349,N_13968,N_12014);
or U22350 (N_22350,N_16642,N_14295);
xnor U22351 (N_22351,N_12873,N_12255);
or U22352 (N_22352,N_15292,N_16014);
or U22353 (N_22353,N_13490,N_13150);
xor U22354 (N_22354,N_14936,N_12594);
nor U22355 (N_22355,N_12536,N_12711);
nand U22356 (N_22356,N_14564,N_16499);
xor U22357 (N_22357,N_13033,N_16457);
xnor U22358 (N_22358,N_15641,N_16656);
and U22359 (N_22359,N_14306,N_15226);
xor U22360 (N_22360,N_13730,N_15115);
and U22361 (N_22361,N_17955,N_17621);
nor U22362 (N_22362,N_13117,N_13801);
or U22363 (N_22363,N_15203,N_14314);
and U22364 (N_22364,N_16793,N_15681);
xnor U22365 (N_22365,N_16467,N_17150);
and U22366 (N_22366,N_14668,N_15364);
or U22367 (N_22367,N_14872,N_12809);
and U22368 (N_22368,N_14931,N_12705);
xnor U22369 (N_22369,N_13484,N_12289);
or U22370 (N_22370,N_16016,N_12815);
xnor U22371 (N_22371,N_16588,N_13669);
nand U22372 (N_22372,N_13889,N_12295);
and U22373 (N_22373,N_16278,N_13832);
nor U22374 (N_22374,N_15954,N_15564);
nand U22375 (N_22375,N_16707,N_16669);
xnor U22376 (N_22376,N_15136,N_15955);
and U22377 (N_22377,N_12365,N_15126);
xnor U22378 (N_22378,N_16786,N_13420);
and U22379 (N_22379,N_15218,N_14364);
xor U22380 (N_22380,N_15782,N_17279);
or U22381 (N_22381,N_14905,N_16706);
nand U22382 (N_22382,N_14910,N_14031);
nor U22383 (N_22383,N_14880,N_15928);
and U22384 (N_22384,N_16865,N_17168);
or U22385 (N_22385,N_13676,N_13428);
or U22386 (N_22386,N_17236,N_16726);
and U22387 (N_22387,N_17320,N_13145);
xor U22388 (N_22388,N_14563,N_12582);
nand U22389 (N_22389,N_16970,N_14323);
nor U22390 (N_22390,N_17691,N_13903);
xnor U22391 (N_22391,N_14926,N_15371);
or U22392 (N_22392,N_17430,N_13508);
nor U22393 (N_22393,N_12431,N_14417);
xor U22394 (N_22394,N_16553,N_13011);
or U22395 (N_22395,N_17988,N_14888);
nor U22396 (N_22396,N_17136,N_14434);
and U22397 (N_22397,N_17702,N_13122);
and U22398 (N_22398,N_17742,N_13940);
and U22399 (N_22399,N_15050,N_12017);
nor U22400 (N_22400,N_12862,N_15375);
xor U22401 (N_22401,N_14973,N_17006);
nor U22402 (N_22402,N_13405,N_12093);
nor U22403 (N_22403,N_17861,N_12220);
or U22404 (N_22404,N_15531,N_14442);
or U22405 (N_22405,N_15512,N_13982);
nand U22406 (N_22406,N_15939,N_14322);
and U22407 (N_22407,N_16856,N_17101);
or U22408 (N_22408,N_17811,N_15779);
or U22409 (N_22409,N_15806,N_15625);
xor U22410 (N_22410,N_14090,N_12039);
nor U22411 (N_22411,N_16613,N_16323);
xor U22412 (N_22412,N_17381,N_14691);
or U22413 (N_22413,N_12573,N_16954);
or U22414 (N_22414,N_17070,N_14049);
or U22415 (N_22415,N_12280,N_17813);
nand U22416 (N_22416,N_17638,N_13048);
and U22417 (N_22417,N_14160,N_12927);
nor U22418 (N_22418,N_16934,N_16956);
or U22419 (N_22419,N_15002,N_17078);
nor U22420 (N_22420,N_13768,N_17734);
xnor U22421 (N_22421,N_14141,N_12187);
xor U22422 (N_22422,N_16064,N_13917);
nand U22423 (N_22423,N_14704,N_16083);
nor U22424 (N_22424,N_14897,N_15219);
or U22425 (N_22425,N_13490,N_16160);
or U22426 (N_22426,N_17387,N_13879);
or U22427 (N_22427,N_17088,N_14028);
nor U22428 (N_22428,N_15793,N_13882);
nand U22429 (N_22429,N_13557,N_13297);
nor U22430 (N_22430,N_13825,N_13618);
xnor U22431 (N_22431,N_13887,N_12493);
or U22432 (N_22432,N_14979,N_15240);
xor U22433 (N_22433,N_17011,N_15199);
or U22434 (N_22434,N_12241,N_16596);
nand U22435 (N_22435,N_15216,N_16642);
nor U22436 (N_22436,N_15353,N_17875);
xnor U22437 (N_22437,N_16715,N_12879);
and U22438 (N_22438,N_17671,N_16243);
and U22439 (N_22439,N_12734,N_13434);
and U22440 (N_22440,N_15242,N_13592);
nand U22441 (N_22441,N_16472,N_14158);
and U22442 (N_22442,N_13337,N_14826);
or U22443 (N_22443,N_15362,N_13520);
nor U22444 (N_22444,N_16230,N_12994);
and U22445 (N_22445,N_12367,N_12260);
or U22446 (N_22446,N_12370,N_16704);
or U22447 (N_22447,N_15251,N_16571);
or U22448 (N_22448,N_15690,N_15570);
xnor U22449 (N_22449,N_17448,N_14585);
xnor U22450 (N_22450,N_15992,N_13324);
nand U22451 (N_22451,N_14871,N_16025);
xnor U22452 (N_22452,N_13216,N_17344);
xnor U22453 (N_22453,N_13059,N_14843);
nor U22454 (N_22454,N_17150,N_12812);
nand U22455 (N_22455,N_17015,N_17463);
and U22456 (N_22456,N_13342,N_13030);
or U22457 (N_22457,N_13034,N_14232);
nand U22458 (N_22458,N_16215,N_17210);
and U22459 (N_22459,N_12943,N_17857);
xor U22460 (N_22460,N_15729,N_14789);
nand U22461 (N_22461,N_14299,N_14012);
nor U22462 (N_22462,N_13367,N_16073);
and U22463 (N_22463,N_16521,N_13886);
and U22464 (N_22464,N_17763,N_17579);
and U22465 (N_22465,N_15482,N_14725);
or U22466 (N_22466,N_16729,N_13930);
or U22467 (N_22467,N_12591,N_17227);
and U22468 (N_22468,N_16512,N_12535);
nand U22469 (N_22469,N_17837,N_13293);
nand U22470 (N_22470,N_14904,N_14692);
xor U22471 (N_22471,N_16117,N_15922);
xor U22472 (N_22472,N_12154,N_12597);
or U22473 (N_22473,N_15397,N_13048);
nand U22474 (N_22474,N_12689,N_17000);
xnor U22475 (N_22475,N_13661,N_15960);
xor U22476 (N_22476,N_14615,N_12837);
xnor U22477 (N_22477,N_17760,N_16752);
xor U22478 (N_22478,N_17868,N_12533);
nand U22479 (N_22479,N_17237,N_14386);
xnor U22480 (N_22480,N_16577,N_15265);
xnor U22481 (N_22481,N_15441,N_13438);
and U22482 (N_22482,N_15000,N_17380);
nor U22483 (N_22483,N_15356,N_12993);
and U22484 (N_22484,N_14073,N_16328);
xnor U22485 (N_22485,N_14545,N_12795);
nor U22486 (N_22486,N_13772,N_16827);
nand U22487 (N_22487,N_14166,N_16033);
and U22488 (N_22488,N_12367,N_13519);
nor U22489 (N_22489,N_16742,N_14314);
xnor U22490 (N_22490,N_16167,N_14155);
nand U22491 (N_22491,N_14709,N_16688);
nor U22492 (N_22492,N_17621,N_17389);
or U22493 (N_22493,N_14131,N_14691);
or U22494 (N_22494,N_17076,N_13422);
xnor U22495 (N_22495,N_16908,N_13202);
nand U22496 (N_22496,N_15517,N_16440);
nor U22497 (N_22497,N_15199,N_13611);
nor U22498 (N_22498,N_16299,N_15392);
nor U22499 (N_22499,N_14744,N_17864);
and U22500 (N_22500,N_14794,N_16573);
and U22501 (N_22501,N_15687,N_15983);
or U22502 (N_22502,N_17111,N_16170);
and U22503 (N_22503,N_15167,N_13855);
xnor U22504 (N_22504,N_16921,N_16633);
and U22505 (N_22505,N_15195,N_15719);
nand U22506 (N_22506,N_14729,N_13778);
and U22507 (N_22507,N_13526,N_13229);
xor U22508 (N_22508,N_12634,N_14688);
or U22509 (N_22509,N_16063,N_14464);
nand U22510 (N_22510,N_13916,N_15434);
and U22511 (N_22511,N_13513,N_14464);
or U22512 (N_22512,N_12285,N_15162);
nand U22513 (N_22513,N_14386,N_16336);
and U22514 (N_22514,N_16717,N_15972);
and U22515 (N_22515,N_12150,N_16048);
and U22516 (N_22516,N_14670,N_15006);
xnor U22517 (N_22517,N_12811,N_13440);
xor U22518 (N_22518,N_13976,N_17923);
xnor U22519 (N_22519,N_16818,N_16301);
or U22520 (N_22520,N_15519,N_17505);
or U22521 (N_22521,N_13786,N_17856);
nand U22522 (N_22522,N_17665,N_14026);
and U22523 (N_22523,N_15860,N_13084);
and U22524 (N_22524,N_15138,N_16091);
and U22525 (N_22525,N_15852,N_15577);
or U22526 (N_22526,N_16082,N_12046);
or U22527 (N_22527,N_16818,N_17926);
nand U22528 (N_22528,N_14729,N_15031);
nor U22529 (N_22529,N_16822,N_13305);
and U22530 (N_22530,N_16716,N_13220);
or U22531 (N_22531,N_13000,N_15730);
nor U22532 (N_22532,N_12807,N_14332);
or U22533 (N_22533,N_15571,N_14930);
or U22534 (N_22534,N_17359,N_17645);
xnor U22535 (N_22535,N_15725,N_13991);
nand U22536 (N_22536,N_12951,N_16723);
xor U22537 (N_22537,N_13018,N_16256);
and U22538 (N_22538,N_15942,N_17999);
xnor U22539 (N_22539,N_12165,N_14656);
nand U22540 (N_22540,N_14624,N_13536);
nand U22541 (N_22541,N_16421,N_13524);
nor U22542 (N_22542,N_13612,N_13684);
nand U22543 (N_22543,N_15083,N_16291);
or U22544 (N_22544,N_17323,N_17862);
nand U22545 (N_22545,N_16648,N_15952);
nand U22546 (N_22546,N_16871,N_15739);
or U22547 (N_22547,N_12342,N_17542);
nand U22548 (N_22548,N_14153,N_16431);
or U22549 (N_22549,N_15521,N_16051);
xnor U22550 (N_22550,N_14652,N_17412);
nor U22551 (N_22551,N_12126,N_12314);
or U22552 (N_22552,N_15992,N_12868);
nand U22553 (N_22553,N_12153,N_15449);
nand U22554 (N_22554,N_14324,N_15012);
xor U22555 (N_22555,N_15195,N_12675);
nand U22556 (N_22556,N_13541,N_15963);
nor U22557 (N_22557,N_13156,N_12617);
nor U22558 (N_22558,N_14903,N_13244);
nor U22559 (N_22559,N_17031,N_12146);
nand U22560 (N_22560,N_17964,N_12007);
xor U22561 (N_22561,N_14399,N_15171);
xor U22562 (N_22562,N_13031,N_14065);
xor U22563 (N_22563,N_16988,N_13990);
nand U22564 (N_22564,N_14937,N_16327);
and U22565 (N_22565,N_15906,N_15733);
or U22566 (N_22566,N_14807,N_16548);
or U22567 (N_22567,N_15620,N_13460);
and U22568 (N_22568,N_12132,N_14591);
xor U22569 (N_22569,N_15900,N_16141);
and U22570 (N_22570,N_15436,N_17128);
or U22571 (N_22571,N_16751,N_17950);
and U22572 (N_22572,N_15005,N_14364);
or U22573 (N_22573,N_17520,N_12050);
nand U22574 (N_22574,N_12615,N_12659);
or U22575 (N_22575,N_16495,N_14087);
nor U22576 (N_22576,N_15952,N_17599);
xor U22577 (N_22577,N_13749,N_13406);
or U22578 (N_22578,N_17691,N_12524);
xor U22579 (N_22579,N_16374,N_12783);
and U22580 (N_22580,N_13538,N_15324);
nor U22581 (N_22581,N_12406,N_16593);
or U22582 (N_22582,N_14366,N_15779);
nand U22583 (N_22583,N_12944,N_15606);
nor U22584 (N_22584,N_17007,N_15804);
nor U22585 (N_22585,N_15986,N_12454);
xor U22586 (N_22586,N_16306,N_12206);
or U22587 (N_22587,N_15037,N_13866);
and U22588 (N_22588,N_16484,N_16415);
or U22589 (N_22589,N_17734,N_15400);
xor U22590 (N_22590,N_15175,N_14783);
nand U22591 (N_22591,N_13997,N_12399);
nor U22592 (N_22592,N_16091,N_14169);
or U22593 (N_22593,N_16808,N_14752);
nand U22594 (N_22594,N_14948,N_14113);
or U22595 (N_22595,N_17111,N_13916);
xor U22596 (N_22596,N_14437,N_15945);
and U22597 (N_22597,N_13177,N_12156);
xor U22598 (N_22598,N_17220,N_15657);
nand U22599 (N_22599,N_15126,N_12233);
and U22600 (N_22600,N_13107,N_15786);
xor U22601 (N_22601,N_14190,N_15615);
nand U22602 (N_22602,N_15719,N_13552);
nand U22603 (N_22603,N_15836,N_12063);
and U22604 (N_22604,N_16692,N_17852);
or U22605 (N_22605,N_12363,N_17665);
nor U22606 (N_22606,N_12393,N_12536);
and U22607 (N_22607,N_12853,N_14026);
or U22608 (N_22608,N_14634,N_15685);
or U22609 (N_22609,N_15056,N_16383);
nor U22610 (N_22610,N_14218,N_16189);
or U22611 (N_22611,N_14913,N_17217);
or U22612 (N_22612,N_15899,N_16635);
nor U22613 (N_22613,N_13417,N_12856);
or U22614 (N_22614,N_13142,N_16593);
or U22615 (N_22615,N_13432,N_16869);
or U22616 (N_22616,N_15735,N_17309);
or U22617 (N_22617,N_14905,N_16948);
xnor U22618 (N_22618,N_16191,N_16284);
nand U22619 (N_22619,N_17031,N_17278);
and U22620 (N_22620,N_12573,N_17296);
and U22621 (N_22621,N_14146,N_12386);
or U22622 (N_22622,N_14388,N_14382);
and U22623 (N_22623,N_14412,N_14209);
or U22624 (N_22624,N_16574,N_12195);
xnor U22625 (N_22625,N_15448,N_15481);
or U22626 (N_22626,N_12488,N_12754);
or U22627 (N_22627,N_16991,N_17305);
xor U22628 (N_22628,N_14751,N_14690);
or U22629 (N_22629,N_16633,N_14396);
nand U22630 (N_22630,N_15311,N_16831);
xnor U22631 (N_22631,N_14311,N_13003);
and U22632 (N_22632,N_12085,N_14607);
and U22633 (N_22633,N_17991,N_17738);
or U22634 (N_22634,N_12869,N_14568);
nor U22635 (N_22635,N_13422,N_17033);
nand U22636 (N_22636,N_15528,N_15838);
nor U22637 (N_22637,N_12212,N_17614);
xor U22638 (N_22638,N_13460,N_12860);
or U22639 (N_22639,N_13524,N_13483);
or U22640 (N_22640,N_12181,N_17923);
nand U22641 (N_22641,N_12769,N_17482);
nor U22642 (N_22642,N_15372,N_14048);
or U22643 (N_22643,N_13301,N_14603);
or U22644 (N_22644,N_16257,N_12865);
nor U22645 (N_22645,N_12252,N_15308);
or U22646 (N_22646,N_12286,N_15087);
and U22647 (N_22647,N_14495,N_15006);
or U22648 (N_22648,N_14769,N_16949);
nor U22649 (N_22649,N_14948,N_16583);
nand U22650 (N_22650,N_12859,N_14863);
nor U22651 (N_22651,N_13686,N_12682);
or U22652 (N_22652,N_12876,N_12215);
nand U22653 (N_22653,N_12410,N_15649);
or U22654 (N_22654,N_15319,N_12700);
xor U22655 (N_22655,N_13617,N_14583);
nand U22656 (N_22656,N_12527,N_15827);
and U22657 (N_22657,N_17785,N_12679);
xor U22658 (N_22658,N_13068,N_14633);
or U22659 (N_22659,N_16604,N_16499);
or U22660 (N_22660,N_12540,N_13447);
nand U22661 (N_22661,N_12349,N_12657);
nand U22662 (N_22662,N_14613,N_15022);
nor U22663 (N_22663,N_13799,N_17198);
nand U22664 (N_22664,N_14910,N_17906);
nand U22665 (N_22665,N_15485,N_14271);
xor U22666 (N_22666,N_16927,N_17709);
nand U22667 (N_22667,N_17639,N_12563);
nor U22668 (N_22668,N_14044,N_13258);
or U22669 (N_22669,N_14341,N_13309);
nor U22670 (N_22670,N_13495,N_16371);
or U22671 (N_22671,N_12962,N_13273);
or U22672 (N_22672,N_17654,N_12456);
xnor U22673 (N_22673,N_12567,N_15989);
and U22674 (N_22674,N_15638,N_13543);
or U22675 (N_22675,N_17974,N_17865);
nor U22676 (N_22676,N_16019,N_14742);
and U22677 (N_22677,N_14888,N_14310);
xor U22678 (N_22678,N_17999,N_13479);
nor U22679 (N_22679,N_12160,N_14706);
or U22680 (N_22680,N_16464,N_14522);
nor U22681 (N_22681,N_15938,N_12088);
or U22682 (N_22682,N_12830,N_15788);
nand U22683 (N_22683,N_13531,N_16907);
nor U22684 (N_22684,N_12635,N_15340);
nor U22685 (N_22685,N_15921,N_14630);
nand U22686 (N_22686,N_13506,N_14679);
or U22687 (N_22687,N_15651,N_13165);
and U22688 (N_22688,N_12898,N_14252);
and U22689 (N_22689,N_14571,N_14286);
and U22690 (N_22690,N_16631,N_13403);
and U22691 (N_22691,N_12238,N_16158);
or U22692 (N_22692,N_14001,N_16624);
xnor U22693 (N_22693,N_17577,N_13081);
xor U22694 (N_22694,N_12403,N_13785);
xor U22695 (N_22695,N_13903,N_14185);
nand U22696 (N_22696,N_12659,N_17773);
and U22697 (N_22697,N_13779,N_15881);
or U22698 (N_22698,N_14938,N_13448);
nand U22699 (N_22699,N_16045,N_12733);
and U22700 (N_22700,N_17629,N_14643);
nor U22701 (N_22701,N_13442,N_15172);
xor U22702 (N_22702,N_13087,N_13711);
and U22703 (N_22703,N_17107,N_12418);
xor U22704 (N_22704,N_14258,N_16855);
nand U22705 (N_22705,N_12683,N_17056);
nand U22706 (N_22706,N_12639,N_16540);
xnor U22707 (N_22707,N_13641,N_13163);
xor U22708 (N_22708,N_14396,N_13258);
xnor U22709 (N_22709,N_12338,N_15101);
nor U22710 (N_22710,N_16736,N_17186);
nand U22711 (N_22711,N_15847,N_14216);
and U22712 (N_22712,N_15208,N_15619);
nand U22713 (N_22713,N_13541,N_12650);
nor U22714 (N_22714,N_14122,N_17772);
nor U22715 (N_22715,N_15941,N_14354);
xnor U22716 (N_22716,N_17281,N_16420);
and U22717 (N_22717,N_17184,N_15815);
and U22718 (N_22718,N_16417,N_12006);
nand U22719 (N_22719,N_15419,N_17598);
and U22720 (N_22720,N_14571,N_14701);
nor U22721 (N_22721,N_16241,N_16945);
or U22722 (N_22722,N_16326,N_12622);
or U22723 (N_22723,N_16547,N_14026);
nor U22724 (N_22724,N_17699,N_17483);
nor U22725 (N_22725,N_13801,N_12906);
nand U22726 (N_22726,N_15302,N_15860);
nand U22727 (N_22727,N_15214,N_14133);
nand U22728 (N_22728,N_12700,N_17950);
xor U22729 (N_22729,N_15022,N_17122);
nor U22730 (N_22730,N_15839,N_15318);
xnor U22731 (N_22731,N_17201,N_12688);
or U22732 (N_22732,N_13759,N_15240);
nor U22733 (N_22733,N_14440,N_16130);
nand U22734 (N_22734,N_17235,N_14490);
nor U22735 (N_22735,N_15632,N_14573);
or U22736 (N_22736,N_14169,N_12537);
xnor U22737 (N_22737,N_13362,N_16623);
and U22738 (N_22738,N_12573,N_15831);
nor U22739 (N_22739,N_13484,N_17959);
nor U22740 (N_22740,N_17230,N_12715);
or U22741 (N_22741,N_13615,N_12741);
nor U22742 (N_22742,N_17501,N_14034);
xnor U22743 (N_22743,N_16671,N_15610);
or U22744 (N_22744,N_17721,N_13277);
nand U22745 (N_22745,N_15721,N_14051);
and U22746 (N_22746,N_15360,N_16176);
xor U22747 (N_22747,N_12309,N_15249);
and U22748 (N_22748,N_13930,N_17390);
or U22749 (N_22749,N_13912,N_16246);
or U22750 (N_22750,N_14647,N_17182);
nor U22751 (N_22751,N_12242,N_17945);
nor U22752 (N_22752,N_12355,N_15154);
or U22753 (N_22753,N_15041,N_16230);
or U22754 (N_22754,N_14859,N_14362);
nor U22755 (N_22755,N_13772,N_15497);
nand U22756 (N_22756,N_13586,N_16192);
or U22757 (N_22757,N_13343,N_16037);
or U22758 (N_22758,N_13302,N_12854);
and U22759 (N_22759,N_13265,N_16486);
and U22760 (N_22760,N_15672,N_13197);
nor U22761 (N_22761,N_16072,N_16046);
nor U22762 (N_22762,N_16019,N_16260);
xnor U22763 (N_22763,N_17509,N_15253);
nor U22764 (N_22764,N_13423,N_13425);
nor U22765 (N_22765,N_16330,N_14245);
nor U22766 (N_22766,N_16113,N_16841);
nor U22767 (N_22767,N_12648,N_16238);
and U22768 (N_22768,N_12594,N_16370);
nand U22769 (N_22769,N_13109,N_13983);
xor U22770 (N_22770,N_13833,N_16062);
nor U22771 (N_22771,N_14717,N_16025);
nand U22772 (N_22772,N_13881,N_13320);
nand U22773 (N_22773,N_16346,N_13016);
nor U22774 (N_22774,N_13397,N_14337);
nand U22775 (N_22775,N_13793,N_13082);
nand U22776 (N_22776,N_16030,N_16359);
nand U22777 (N_22777,N_12032,N_16375);
xnor U22778 (N_22778,N_15811,N_12627);
nand U22779 (N_22779,N_13946,N_16079);
nor U22780 (N_22780,N_16052,N_17373);
or U22781 (N_22781,N_16754,N_15791);
nor U22782 (N_22782,N_12424,N_12014);
or U22783 (N_22783,N_15097,N_13999);
and U22784 (N_22784,N_14500,N_12458);
nand U22785 (N_22785,N_15392,N_13500);
nand U22786 (N_22786,N_15240,N_17257);
nand U22787 (N_22787,N_14168,N_14457);
and U22788 (N_22788,N_15248,N_16564);
and U22789 (N_22789,N_17427,N_15701);
nor U22790 (N_22790,N_16222,N_15998);
and U22791 (N_22791,N_16901,N_16131);
xnor U22792 (N_22792,N_16336,N_12624);
nand U22793 (N_22793,N_15242,N_14908);
or U22794 (N_22794,N_12413,N_12730);
and U22795 (N_22795,N_15654,N_17239);
nand U22796 (N_22796,N_13456,N_17935);
or U22797 (N_22797,N_13869,N_13469);
xnor U22798 (N_22798,N_12290,N_15727);
xor U22799 (N_22799,N_14583,N_15053);
xnor U22800 (N_22800,N_12763,N_14787);
nand U22801 (N_22801,N_15545,N_17007);
and U22802 (N_22802,N_14011,N_14656);
xnor U22803 (N_22803,N_14240,N_15482);
nor U22804 (N_22804,N_12866,N_15564);
or U22805 (N_22805,N_16183,N_14910);
nor U22806 (N_22806,N_15955,N_15977);
nand U22807 (N_22807,N_14667,N_14106);
xor U22808 (N_22808,N_17940,N_13726);
nor U22809 (N_22809,N_17372,N_16412);
xor U22810 (N_22810,N_13651,N_12844);
xor U22811 (N_22811,N_13766,N_15802);
and U22812 (N_22812,N_13693,N_15534);
nand U22813 (N_22813,N_17801,N_13888);
and U22814 (N_22814,N_15096,N_15048);
nand U22815 (N_22815,N_12532,N_17046);
nor U22816 (N_22816,N_16604,N_16151);
nand U22817 (N_22817,N_17875,N_12298);
or U22818 (N_22818,N_17747,N_14503);
or U22819 (N_22819,N_16748,N_14209);
and U22820 (N_22820,N_15617,N_13903);
xor U22821 (N_22821,N_14156,N_14404);
nor U22822 (N_22822,N_16064,N_13077);
or U22823 (N_22823,N_16482,N_16514);
nor U22824 (N_22824,N_16182,N_12017);
and U22825 (N_22825,N_12015,N_15282);
nor U22826 (N_22826,N_15670,N_17579);
and U22827 (N_22827,N_15964,N_16578);
or U22828 (N_22828,N_12091,N_15994);
or U22829 (N_22829,N_16143,N_17168);
xor U22830 (N_22830,N_16203,N_16556);
nand U22831 (N_22831,N_16660,N_15017);
nand U22832 (N_22832,N_12352,N_13895);
nand U22833 (N_22833,N_14274,N_16714);
nor U22834 (N_22834,N_13707,N_15141);
and U22835 (N_22835,N_12738,N_13010);
or U22836 (N_22836,N_17175,N_14496);
nor U22837 (N_22837,N_17393,N_16689);
nand U22838 (N_22838,N_13813,N_15788);
nand U22839 (N_22839,N_15949,N_16384);
nor U22840 (N_22840,N_12154,N_12648);
or U22841 (N_22841,N_17615,N_17742);
or U22842 (N_22842,N_15771,N_13393);
or U22843 (N_22843,N_17063,N_17127);
nand U22844 (N_22844,N_13529,N_17508);
nand U22845 (N_22845,N_16193,N_12947);
nand U22846 (N_22846,N_13219,N_17298);
or U22847 (N_22847,N_12639,N_14238);
nor U22848 (N_22848,N_14697,N_13403);
or U22849 (N_22849,N_17324,N_16089);
or U22850 (N_22850,N_14552,N_16620);
xnor U22851 (N_22851,N_12871,N_13575);
xnor U22852 (N_22852,N_13054,N_15133);
nand U22853 (N_22853,N_12814,N_16595);
and U22854 (N_22854,N_17808,N_16020);
nand U22855 (N_22855,N_17263,N_17977);
nand U22856 (N_22856,N_14434,N_12929);
and U22857 (N_22857,N_17683,N_15590);
or U22858 (N_22858,N_14729,N_13645);
xnor U22859 (N_22859,N_14782,N_16814);
or U22860 (N_22860,N_16487,N_12371);
or U22861 (N_22861,N_17143,N_14576);
and U22862 (N_22862,N_16725,N_13651);
nand U22863 (N_22863,N_12937,N_14646);
or U22864 (N_22864,N_13595,N_17885);
and U22865 (N_22865,N_16634,N_12954);
nand U22866 (N_22866,N_12805,N_16809);
nand U22867 (N_22867,N_14435,N_15540);
nand U22868 (N_22868,N_14091,N_12269);
nor U22869 (N_22869,N_16860,N_17058);
and U22870 (N_22870,N_13700,N_17439);
nand U22871 (N_22871,N_13920,N_17167);
and U22872 (N_22872,N_14942,N_13975);
nor U22873 (N_22873,N_16947,N_15671);
or U22874 (N_22874,N_15235,N_14596);
xnor U22875 (N_22875,N_13102,N_14259);
nor U22876 (N_22876,N_16993,N_16812);
and U22877 (N_22877,N_14827,N_16398);
and U22878 (N_22878,N_17713,N_14238);
nor U22879 (N_22879,N_15671,N_13476);
or U22880 (N_22880,N_17437,N_14120);
xnor U22881 (N_22881,N_16741,N_12716);
nor U22882 (N_22882,N_14135,N_13585);
or U22883 (N_22883,N_17290,N_13520);
nor U22884 (N_22884,N_13825,N_14967);
or U22885 (N_22885,N_14285,N_16962);
nand U22886 (N_22886,N_13984,N_16093);
nand U22887 (N_22887,N_12516,N_14395);
and U22888 (N_22888,N_13131,N_17113);
nor U22889 (N_22889,N_13503,N_12160);
or U22890 (N_22890,N_17075,N_14860);
xnor U22891 (N_22891,N_15877,N_15854);
and U22892 (N_22892,N_16897,N_12553);
nand U22893 (N_22893,N_15224,N_13251);
nand U22894 (N_22894,N_15417,N_16277);
nand U22895 (N_22895,N_14135,N_13900);
nand U22896 (N_22896,N_16455,N_15256);
xnor U22897 (N_22897,N_13383,N_17486);
or U22898 (N_22898,N_16472,N_15852);
nor U22899 (N_22899,N_17409,N_12216);
nor U22900 (N_22900,N_12591,N_17119);
nor U22901 (N_22901,N_14362,N_15932);
nor U22902 (N_22902,N_17124,N_15583);
nor U22903 (N_22903,N_16422,N_15010);
nand U22904 (N_22904,N_16742,N_12557);
nand U22905 (N_22905,N_14255,N_16974);
nand U22906 (N_22906,N_17977,N_14246);
nor U22907 (N_22907,N_13123,N_14694);
nor U22908 (N_22908,N_13652,N_17940);
xor U22909 (N_22909,N_15332,N_17647);
nand U22910 (N_22910,N_13798,N_16285);
and U22911 (N_22911,N_13930,N_15475);
nor U22912 (N_22912,N_17197,N_12221);
or U22913 (N_22913,N_12150,N_15839);
or U22914 (N_22914,N_15776,N_12639);
and U22915 (N_22915,N_16210,N_16775);
or U22916 (N_22916,N_15437,N_15102);
nor U22917 (N_22917,N_17999,N_17438);
or U22918 (N_22918,N_12909,N_14911);
nand U22919 (N_22919,N_17149,N_14002);
or U22920 (N_22920,N_17004,N_17332);
or U22921 (N_22921,N_17113,N_12829);
nand U22922 (N_22922,N_17806,N_15366);
or U22923 (N_22923,N_16331,N_17113);
or U22924 (N_22924,N_16382,N_17513);
xnor U22925 (N_22925,N_12256,N_16234);
and U22926 (N_22926,N_13600,N_12500);
nor U22927 (N_22927,N_17302,N_12424);
xor U22928 (N_22928,N_14667,N_12764);
and U22929 (N_22929,N_17889,N_12654);
nand U22930 (N_22930,N_17825,N_12386);
or U22931 (N_22931,N_12107,N_16802);
nand U22932 (N_22932,N_15548,N_15222);
nor U22933 (N_22933,N_14566,N_14227);
or U22934 (N_22934,N_15554,N_17024);
and U22935 (N_22935,N_17369,N_12314);
xnor U22936 (N_22936,N_12906,N_12722);
or U22937 (N_22937,N_17397,N_16968);
xor U22938 (N_22938,N_15375,N_16951);
xnor U22939 (N_22939,N_16701,N_16869);
and U22940 (N_22940,N_16703,N_16945);
xnor U22941 (N_22941,N_17947,N_14832);
xor U22942 (N_22942,N_17240,N_17909);
or U22943 (N_22943,N_17579,N_14284);
and U22944 (N_22944,N_14781,N_12661);
and U22945 (N_22945,N_13505,N_13128);
or U22946 (N_22946,N_12606,N_13485);
and U22947 (N_22947,N_16122,N_17690);
nor U22948 (N_22948,N_15748,N_17386);
or U22949 (N_22949,N_15237,N_14144);
or U22950 (N_22950,N_15216,N_17859);
nor U22951 (N_22951,N_17275,N_17916);
and U22952 (N_22952,N_13654,N_16707);
or U22953 (N_22953,N_14998,N_12709);
xnor U22954 (N_22954,N_13375,N_14535);
and U22955 (N_22955,N_13369,N_13441);
nor U22956 (N_22956,N_12382,N_16386);
nor U22957 (N_22957,N_13880,N_14638);
nor U22958 (N_22958,N_13182,N_12043);
and U22959 (N_22959,N_12735,N_16136);
nand U22960 (N_22960,N_17465,N_13590);
or U22961 (N_22961,N_14878,N_12835);
nor U22962 (N_22962,N_15609,N_17068);
nand U22963 (N_22963,N_13207,N_17229);
and U22964 (N_22964,N_15518,N_13628);
nor U22965 (N_22965,N_12447,N_12471);
and U22966 (N_22966,N_15889,N_14298);
nor U22967 (N_22967,N_13609,N_14743);
or U22968 (N_22968,N_17291,N_13222);
nand U22969 (N_22969,N_17092,N_14908);
xor U22970 (N_22970,N_13764,N_12378);
or U22971 (N_22971,N_17406,N_16005);
nand U22972 (N_22972,N_16751,N_15424);
and U22973 (N_22973,N_15121,N_15250);
and U22974 (N_22974,N_14065,N_14070);
and U22975 (N_22975,N_13671,N_12917);
and U22976 (N_22976,N_16916,N_14865);
nor U22977 (N_22977,N_12575,N_13950);
nor U22978 (N_22978,N_12430,N_12739);
xnor U22979 (N_22979,N_16086,N_12565);
and U22980 (N_22980,N_12086,N_15898);
nor U22981 (N_22981,N_16983,N_12929);
and U22982 (N_22982,N_14751,N_12312);
nand U22983 (N_22983,N_12641,N_12307);
nor U22984 (N_22984,N_14556,N_17637);
or U22985 (N_22985,N_17942,N_13153);
or U22986 (N_22986,N_16368,N_13975);
xnor U22987 (N_22987,N_12507,N_16460);
or U22988 (N_22988,N_13722,N_15442);
nand U22989 (N_22989,N_15616,N_17896);
nor U22990 (N_22990,N_13320,N_17901);
and U22991 (N_22991,N_16995,N_13350);
nor U22992 (N_22992,N_17795,N_17870);
and U22993 (N_22993,N_12586,N_15995);
xnor U22994 (N_22994,N_15925,N_15207);
nor U22995 (N_22995,N_14087,N_16001);
or U22996 (N_22996,N_12336,N_12345);
or U22997 (N_22997,N_13570,N_12601);
nand U22998 (N_22998,N_13891,N_17394);
and U22999 (N_22999,N_12630,N_16006);
nand U23000 (N_23000,N_13498,N_12468);
and U23001 (N_23001,N_17897,N_13198);
or U23002 (N_23002,N_13431,N_15071);
xor U23003 (N_23003,N_14288,N_17043);
nand U23004 (N_23004,N_16457,N_16994);
nor U23005 (N_23005,N_12638,N_12270);
xnor U23006 (N_23006,N_16101,N_14073);
nor U23007 (N_23007,N_13399,N_14302);
nor U23008 (N_23008,N_13730,N_14051);
xor U23009 (N_23009,N_15545,N_15619);
nand U23010 (N_23010,N_12698,N_14060);
nand U23011 (N_23011,N_15929,N_16691);
nand U23012 (N_23012,N_13523,N_13436);
and U23013 (N_23013,N_16304,N_12701);
nor U23014 (N_23014,N_16500,N_12926);
nand U23015 (N_23015,N_13387,N_16266);
xnor U23016 (N_23016,N_14721,N_14054);
nand U23017 (N_23017,N_12155,N_16937);
nor U23018 (N_23018,N_13434,N_14301);
nand U23019 (N_23019,N_13133,N_15779);
xor U23020 (N_23020,N_17980,N_17362);
nand U23021 (N_23021,N_13144,N_17722);
and U23022 (N_23022,N_13881,N_12525);
or U23023 (N_23023,N_14328,N_12321);
or U23024 (N_23024,N_15034,N_17223);
or U23025 (N_23025,N_12681,N_16067);
or U23026 (N_23026,N_13288,N_14803);
and U23027 (N_23027,N_16211,N_16428);
nand U23028 (N_23028,N_15304,N_12027);
nand U23029 (N_23029,N_15634,N_14110);
nor U23030 (N_23030,N_12329,N_13949);
or U23031 (N_23031,N_12794,N_15745);
nand U23032 (N_23032,N_14735,N_16832);
nor U23033 (N_23033,N_12335,N_16691);
or U23034 (N_23034,N_13665,N_16913);
nor U23035 (N_23035,N_13125,N_17809);
and U23036 (N_23036,N_12949,N_13562);
or U23037 (N_23037,N_17816,N_13827);
nor U23038 (N_23038,N_12336,N_16753);
nor U23039 (N_23039,N_15271,N_14896);
nand U23040 (N_23040,N_15820,N_15486);
xor U23041 (N_23041,N_14139,N_14956);
or U23042 (N_23042,N_12794,N_13880);
and U23043 (N_23043,N_13382,N_15173);
nor U23044 (N_23044,N_14668,N_14046);
xnor U23045 (N_23045,N_15835,N_16304);
or U23046 (N_23046,N_14540,N_13397);
nand U23047 (N_23047,N_17483,N_17846);
xor U23048 (N_23048,N_17931,N_16881);
and U23049 (N_23049,N_12662,N_13246);
nor U23050 (N_23050,N_14630,N_17833);
or U23051 (N_23051,N_15351,N_16503);
or U23052 (N_23052,N_17271,N_12033);
nand U23053 (N_23053,N_17002,N_13949);
nor U23054 (N_23054,N_14813,N_14306);
or U23055 (N_23055,N_17431,N_14717);
and U23056 (N_23056,N_13370,N_15734);
xnor U23057 (N_23057,N_17200,N_15328);
nor U23058 (N_23058,N_16915,N_16930);
or U23059 (N_23059,N_17390,N_17035);
and U23060 (N_23060,N_14201,N_13781);
nor U23061 (N_23061,N_14903,N_14899);
nor U23062 (N_23062,N_14682,N_16814);
xor U23063 (N_23063,N_17835,N_13695);
or U23064 (N_23064,N_16501,N_16138);
nand U23065 (N_23065,N_12712,N_13667);
and U23066 (N_23066,N_14127,N_14375);
nand U23067 (N_23067,N_13755,N_12973);
nand U23068 (N_23068,N_15596,N_12322);
and U23069 (N_23069,N_13886,N_12774);
nor U23070 (N_23070,N_12257,N_13792);
nand U23071 (N_23071,N_16211,N_12626);
xnor U23072 (N_23072,N_17194,N_17308);
nor U23073 (N_23073,N_15864,N_17045);
xnor U23074 (N_23074,N_14257,N_15531);
xor U23075 (N_23075,N_14269,N_14694);
or U23076 (N_23076,N_15585,N_13713);
and U23077 (N_23077,N_12745,N_12063);
and U23078 (N_23078,N_12673,N_14854);
or U23079 (N_23079,N_13425,N_17425);
or U23080 (N_23080,N_17522,N_13682);
and U23081 (N_23081,N_14558,N_14941);
xnor U23082 (N_23082,N_12082,N_14989);
xor U23083 (N_23083,N_16448,N_13056);
and U23084 (N_23084,N_14884,N_17974);
or U23085 (N_23085,N_15257,N_17307);
nor U23086 (N_23086,N_12112,N_14112);
nor U23087 (N_23087,N_12689,N_17373);
or U23088 (N_23088,N_17034,N_14874);
nor U23089 (N_23089,N_12243,N_17520);
nand U23090 (N_23090,N_13451,N_14423);
and U23091 (N_23091,N_15250,N_13012);
nor U23092 (N_23092,N_16771,N_14883);
xor U23093 (N_23093,N_17941,N_14318);
xor U23094 (N_23094,N_14339,N_17458);
or U23095 (N_23095,N_13830,N_13307);
nand U23096 (N_23096,N_12935,N_16757);
xnor U23097 (N_23097,N_15081,N_12299);
or U23098 (N_23098,N_15900,N_12050);
xor U23099 (N_23099,N_15353,N_14485);
or U23100 (N_23100,N_17804,N_17446);
nor U23101 (N_23101,N_14988,N_17831);
nor U23102 (N_23102,N_12269,N_12650);
xnor U23103 (N_23103,N_13198,N_16896);
nor U23104 (N_23104,N_16470,N_17131);
xor U23105 (N_23105,N_16234,N_14209);
nor U23106 (N_23106,N_15867,N_14716);
nor U23107 (N_23107,N_14084,N_14078);
xnor U23108 (N_23108,N_16537,N_17837);
nor U23109 (N_23109,N_17858,N_17394);
xnor U23110 (N_23110,N_17087,N_13364);
nand U23111 (N_23111,N_15822,N_13058);
nor U23112 (N_23112,N_17485,N_16397);
nand U23113 (N_23113,N_17205,N_16235);
or U23114 (N_23114,N_17923,N_13162);
nor U23115 (N_23115,N_17826,N_12757);
nor U23116 (N_23116,N_15767,N_14646);
and U23117 (N_23117,N_16662,N_17458);
nand U23118 (N_23118,N_16229,N_14883);
or U23119 (N_23119,N_14108,N_15110);
nand U23120 (N_23120,N_17507,N_12244);
and U23121 (N_23121,N_16997,N_14236);
or U23122 (N_23122,N_13724,N_14601);
nand U23123 (N_23123,N_14817,N_13491);
nand U23124 (N_23124,N_16237,N_12562);
nand U23125 (N_23125,N_16075,N_13071);
nand U23126 (N_23126,N_16850,N_12501);
nor U23127 (N_23127,N_17688,N_15232);
nand U23128 (N_23128,N_16913,N_14678);
xnor U23129 (N_23129,N_17910,N_15997);
nand U23130 (N_23130,N_13478,N_16902);
nor U23131 (N_23131,N_13763,N_16431);
nand U23132 (N_23132,N_16782,N_12124);
or U23133 (N_23133,N_14927,N_14772);
nor U23134 (N_23134,N_17621,N_14274);
and U23135 (N_23135,N_17503,N_15319);
nand U23136 (N_23136,N_13407,N_14799);
nor U23137 (N_23137,N_12521,N_16879);
and U23138 (N_23138,N_12139,N_12916);
nor U23139 (N_23139,N_16001,N_16837);
and U23140 (N_23140,N_17894,N_16995);
nor U23141 (N_23141,N_16536,N_15862);
xor U23142 (N_23142,N_14892,N_17106);
nor U23143 (N_23143,N_17170,N_15072);
and U23144 (N_23144,N_15255,N_12246);
and U23145 (N_23145,N_17836,N_13810);
nand U23146 (N_23146,N_15490,N_13588);
xor U23147 (N_23147,N_13947,N_12086);
and U23148 (N_23148,N_17443,N_14608);
nand U23149 (N_23149,N_14440,N_13565);
nand U23150 (N_23150,N_15400,N_14625);
nor U23151 (N_23151,N_17625,N_12969);
or U23152 (N_23152,N_14522,N_16096);
nor U23153 (N_23153,N_13131,N_15323);
nor U23154 (N_23154,N_15689,N_15708);
or U23155 (N_23155,N_15366,N_13849);
and U23156 (N_23156,N_13038,N_16676);
and U23157 (N_23157,N_12943,N_12193);
nand U23158 (N_23158,N_14528,N_17982);
nand U23159 (N_23159,N_17937,N_15866);
or U23160 (N_23160,N_14342,N_12255);
or U23161 (N_23161,N_12917,N_14202);
and U23162 (N_23162,N_13955,N_16679);
xnor U23163 (N_23163,N_12566,N_17207);
or U23164 (N_23164,N_17117,N_14688);
nand U23165 (N_23165,N_13799,N_14498);
nand U23166 (N_23166,N_13407,N_13904);
nand U23167 (N_23167,N_17334,N_16643);
or U23168 (N_23168,N_13107,N_13867);
or U23169 (N_23169,N_16331,N_17963);
nand U23170 (N_23170,N_16545,N_12682);
nor U23171 (N_23171,N_12042,N_17477);
or U23172 (N_23172,N_14226,N_15945);
xnor U23173 (N_23173,N_17188,N_13100);
xor U23174 (N_23174,N_12952,N_12019);
or U23175 (N_23175,N_15590,N_17533);
xnor U23176 (N_23176,N_15925,N_13108);
or U23177 (N_23177,N_17773,N_15920);
nor U23178 (N_23178,N_15690,N_17531);
and U23179 (N_23179,N_14212,N_16268);
nand U23180 (N_23180,N_14517,N_16742);
and U23181 (N_23181,N_16403,N_14264);
nand U23182 (N_23182,N_17765,N_17561);
and U23183 (N_23183,N_17028,N_13349);
nor U23184 (N_23184,N_13826,N_17949);
nand U23185 (N_23185,N_14367,N_14776);
nor U23186 (N_23186,N_13846,N_15305);
and U23187 (N_23187,N_16152,N_15134);
xor U23188 (N_23188,N_17066,N_13329);
nand U23189 (N_23189,N_16531,N_15342);
nand U23190 (N_23190,N_13265,N_15042);
and U23191 (N_23191,N_16081,N_13867);
or U23192 (N_23192,N_16988,N_17815);
and U23193 (N_23193,N_17000,N_14790);
and U23194 (N_23194,N_16252,N_17626);
nand U23195 (N_23195,N_13525,N_13810);
or U23196 (N_23196,N_14576,N_16392);
nand U23197 (N_23197,N_12820,N_14471);
or U23198 (N_23198,N_13667,N_12310);
or U23199 (N_23199,N_12976,N_13649);
nor U23200 (N_23200,N_14497,N_15766);
and U23201 (N_23201,N_17261,N_15053);
or U23202 (N_23202,N_14875,N_16342);
and U23203 (N_23203,N_13179,N_16682);
nand U23204 (N_23204,N_13781,N_14688);
and U23205 (N_23205,N_17194,N_15030);
or U23206 (N_23206,N_14939,N_17722);
nand U23207 (N_23207,N_12639,N_14298);
nor U23208 (N_23208,N_17289,N_16206);
xnor U23209 (N_23209,N_12863,N_17437);
nand U23210 (N_23210,N_12210,N_13014);
nor U23211 (N_23211,N_14665,N_14232);
or U23212 (N_23212,N_17773,N_12121);
nor U23213 (N_23213,N_13784,N_14313);
or U23214 (N_23214,N_15936,N_12043);
and U23215 (N_23215,N_16737,N_13038);
xor U23216 (N_23216,N_17363,N_15969);
nor U23217 (N_23217,N_13438,N_12087);
nor U23218 (N_23218,N_17378,N_12147);
and U23219 (N_23219,N_17991,N_14846);
xnor U23220 (N_23220,N_15961,N_17721);
nor U23221 (N_23221,N_14395,N_16322);
and U23222 (N_23222,N_12701,N_14531);
nand U23223 (N_23223,N_12082,N_13353);
nor U23224 (N_23224,N_16270,N_14016);
xnor U23225 (N_23225,N_12394,N_15118);
and U23226 (N_23226,N_14548,N_13974);
nand U23227 (N_23227,N_12411,N_16191);
nand U23228 (N_23228,N_15902,N_12845);
and U23229 (N_23229,N_12490,N_14896);
nand U23230 (N_23230,N_12384,N_12469);
or U23231 (N_23231,N_13730,N_12532);
or U23232 (N_23232,N_13567,N_15621);
and U23233 (N_23233,N_17537,N_16220);
nor U23234 (N_23234,N_13310,N_13091);
xor U23235 (N_23235,N_16294,N_16718);
nor U23236 (N_23236,N_15058,N_15224);
nand U23237 (N_23237,N_15979,N_15998);
or U23238 (N_23238,N_12712,N_15646);
xnor U23239 (N_23239,N_17089,N_12907);
and U23240 (N_23240,N_16082,N_14332);
and U23241 (N_23241,N_17171,N_14537);
and U23242 (N_23242,N_12740,N_17418);
nand U23243 (N_23243,N_13920,N_16926);
or U23244 (N_23244,N_14899,N_17053);
or U23245 (N_23245,N_13903,N_16936);
xnor U23246 (N_23246,N_12838,N_15294);
or U23247 (N_23247,N_14876,N_15757);
or U23248 (N_23248,N_14238,N_13301);
or U23249 (N_23249,N_16564,N_14173);
or U23250 (N_23250,N_13176,N_16197);
xor U23251 (N_23251,N_15673,N_12770);
nor U23252 (N_23252,N_12219,N_17486);
xor U23253 (N_23253,N_17309,N_12541);
or U23254 (N_23254,N_12137,N_12293);
xnor U23255 (N_23255,N_12536,N_16976);
and U23256 (N_23256,N_14555,N_13833);
and U23257 (N_23257,N_16369,N_12675);
xnor U23258 (N_23258,N_15213,N_17206);
nand U23259 (N_23259,N_15503,N_12207);
nand U23260 (N_23260,N_15351,N_17437);
nor U23261 (N_23261,N_16381,N_12074);
xnor U23262 (N_23262,N_12120,N_17006);
or U23263 (N_23263,N_15708,N_12062);
or U23264 (N_23264,N_12591,N_13988);
nor U23265 (N_23265,N_17704,N_13304);
and U23266 (N_23266,N_13443,N_16378);
and U23267 (N_23267,N_15050,N_16305);
and U23268 (N_23268,N_13903,N_17026);
xnor U23269 (N_23269,N_17476,N_16191);
nor U23270 (N_23270,N_17244,N_17748);
and U23271 (N_23271,N_16724,N_16206);
and U23272 (N_23272,N_12037,N_12102);
xnor U23273 (N_23273,N_15030,N_14876);
and U23274 (N_23274,N_12078,N_16844);
nand U23275 (N_23275,N_16461,N_13370);
xnor U23276 (N_23276,N_13565,N_12800);
nand U23277 (N_23277,N_17315,N_16219);
xnor U23278 (N_23278,N_15756,N_12788);
xnor U23279 (N_23279,N_13470,N_16191);
and U23280 (N_23280,N_17227,N_15821);
nor U23281 (N_23281,N_12852,N_16673);
and U23282 (N_23282,N_17435,N_12934);
and U23283 (N_23283,N_17973,N_14296);
xor U23284 (N_23284,N_17588,N_17239);
nand U23285 (N_23285,N_17693,N_15697);
or U23286 (N_23286,N_12305,N_17030);
nand U23287 (N_23287,N_13195,N_13176);
or U23288 (N_23288,N_17393,N_16009);
nor U23289 (N_23289,N_12944,N_15312);
nand U23290 (N_23290,N_16119,N_17889);
and U23291 (N_23291,N_15755,N_16710);
nand U23292 (N_23292,N_13435,N_13739);
or U23293 (N_23293,N_17743,N_17626);
and U23294 (N_23294,N_13748,N_16485);
and U23295 (N_23295,N_17889,N_14218);
nor U23296 (N_23296,N_17420,N_15927);
nor U23297 (N_23297,N_16914,N_12724);
nor U23298 (N_23298,N_15819,N_15261);
nand U23299 (N_23299,N_15033,N_17095);
xnor U23300 (N_23300,N_14699,N_16385);
nand U23301 (N_23301,N_17651,N_14293);
or U23302 (N_23302,N_15158,N_17695);
nand U23303 (N_23303,N_14584,N_14794);
or U23304 (N_23304,N_14653,N_12215);
and U23305 (N_23305,N_15015,N_17576);
nor U23306 (N_23306,N_16732,N_16305);
nor U23307 (N_23307,N_12844,N_17423);
and U23308 (N_23308,N_14874,N_12724);
xnor U23309 (N_23309,N_16694,N_17659);
nor U23310 (N_23310,N_16492,N_13549);
and U23311 (N_23311,N_14099,N_17464);
nor U23312 (N_23312,N_14769,N_12430);
or U23313 (N_23313,N_14185,N_12207);
nor U23314 (N_23314,N_14799,N_12404);
or U23315 (N_23315,N_12954,N_17093);
nand U23316 (N_23316,N_13442,N_15248);
nand U23317 (N_23317,N_15850,N_17949);
nor U23318 (N_23318,N_15437,N_17506);
xor U23319 (N_23319,N_15774,N_16996);
xor U23320 (N_23320,N_16874,N_16545);
nor U23321 (N_23321,N_15912,N_14947);
and U23322 (N_23322,N_17627,N_16299);
nor U23323 (N_23323,N_12218,N_12357);
nor U23324 (N_23324,N_15804,N_12921);
nor U23325 (N_23325,N_12437,N_12585);
or U23326 (N_23326,N_16841,N_17961);
xnor U23327 (N_23327,N_13860,N_17541);
or U23328 (N_23328,N_17703,N_15487);
and U23329 (N_23329,N_17345,N_14595);
nor U23330 (N_23330,N_14107,N_15149);
nor U23331 (N_23331,N_14541,N_17669);
xor U23332 (N_23332,N_14020,N_15365);
and U23333 (N_23333,N_15788,N_15912);
xnor U23334 (N_23334,N_14967,N_17691);
or U23335 (N_23335,N_15500,N_16565);
nor U23336 (N_23336,N_17121,N_16342);
nand U23337 (N_23337,N_17442,N_15600);
and U23338 (N_23338,N_12453,N_16212);
xor U23339 (N_23339,N_12322,N_14673);
xor U23340 (N_23340,N_15448,N_15678);
or U23341 (N_23341,N_15735,N_13645);
and U23342 (N_23342,N_15293,N_16858);
nand U23343 (N_23343,N_12971,N_14795);
or U23344 (N_23344,N_17340,N_16062);
or U23345 (N_23345,N_13023,N_16278);
xor U23346 (N_23346,N_13370,N_15719);
or U23347 (N_23347,N_14258,N_15609);
or U23348 (N_23348,N_16301,N_14525);
nand U23349 (N_23349,N_12362,N_16534);
nand U23350 (N_23350,N_13630,N_15582);
nand U23351 (N_23351,N_15448,N_15941);
nor U23352 (N_23352,N_13905,N_14318);
nand U23353 (N_23353,N_14700,N_17581);
and U23354 (N_23354,N_16892,N_13057);
xor U23355 (N_23355,N_17783,N_16621);
nand U23356 (N_23356,N_17323,N_12911);
nor U23357 (N_23357,N_16216,N_16589);
nand U23358 (N_23358,N_17016,N_12053);
nor U23359 (N_23359,N_12268,N_17548);
nor U23360 (N_23360,N_14319,N_17785);
xnor U23361 (N_23361,N_14271,N_17266);
nor U23362 (N_23362,N_16594,N_17804);
nor U23363 (N_23363,N_12158,N_15532);
nand U23364 (N_23364,N_13696,N_14902);
or U23365 (N_23365,N_16098,N_13188);
nor U23366 (N_23366,N_14915,N_16005);
nand U23367 (N_23367,N_13743,N_15838);
nor U23368 (N_23368,N_12861,N_14478);
and U23369 (N_23369,N_15512,N_15396);
xor U23370 (N_23370,N_17882,N_14743);
and U23371 (N_23371,N_16332,N_13522);
nand U23372 (N_23372,N_12306,N_13047);
nor U23373 (N_23373,N_14408,N_14214);
xnor U23374 (N_23374,N_15426,N_14929);
and U23375 (N_23375,N_17066,N_16491);
nand U23376 (N_23376,N_16507,N_13635);
nor U23377 (N_23377,N_15555,N_17621);
or U23378 (N_23378,N_13332,N_14837);
nor U23379 (N_23379,N_12065,N_16487);
xor U23380 (N_23380,N_16714,N_12210);
nand U23381 (N_23381,N_12553,N_13792);
nand U23382 (N_23382,N_16729,N_12652);
nor U23383 (N_23383,N_12116,N_14547);
nand U23384 (N_23384,N_13468,N_15400);
nand U23385 (N_23385,N_16152,N_15666);
and U23386 (N_23386,N_12664,N_16589);
or U23387 (N_23387,N_15508,N_12827);
nand U23388 (N_23388,N_12885,N_13478);
xor U23389 (N_23389,N_12513,N_17823);
xnor U23390 (N_23390,N_12636,N_16767);
or U23391 (N_23391,N_12057,N_16422);
nand U23392 (N_23392,N_12074,N_14126);
nor U23393 (N_23393,N_14358,N_15338);
or U23394 (N_23394,N_12472,N_14626);
nand U23395 (N_23395,N_17003,N_17241);
nor U23396 (N_23396,N_15727,N_16547);
or U23397 (N_23397,N_16615,N_13571);
and U23398 (N_23398,N_13005,N_15390);
nand U23399 (N_23399,N_13179,N_12214);
or U23400 (N_23400,N_15486,N_16293);
xnor U23401 (N_23401,N_13130,N_14051);
or U23402 (N_23402,N_16104,N_12527);
and U23403 (N_23403,N_15320,N_13910);
or U23404 (N_23404,N_14914,N_14379);
nor U23405 (N_23405,N_12938,N_16567);
or U23406 (N_23406,N_12953,N_14969);
and U23407 (N_23407,N_16169,N_14656);
xor U23408 (N_23408,N_16032,N_14877);
xor U23409 (N_23409,N_15865,N_12282);
nand U23410 (N_23410,N_16586,N_16951);
nor U23411 (N_23411,N_14454,N_14335);
or U23412 (N_23412,N_14253,N_14503);
or U23413 (N_23413,N_13021,N_17960);
or U23414 (N_23414,N_13910,N_14701);
xnor U23415 (N_23415,N_16105,N_15437);
nor U23416 (N_23416,N_12847,N_15503);
or U23417 (N_23417,N_17924,N_13695);
nor U23418 (N_23418,N_14453,N_16051);
nand U23419 (N_23419,N_13319,N_15787);
or U23420 (N_23420,N_13550,N_16680);
nor U23421 (N_23421,N_12760,N_16920);
or U23422 (N_23422,N_15551,N_12554);
or U23423 (N_23423,N_12873,N_17403);
and U23424 (N_23424,N_16830,N_15815);
xnor U23425 (N_23425,N_16457,N_14691);
or U23426 (N_23426,N_16217,N_12758);
nor U23427 (N_23427,N_14599,N_16574);
or U23428 (N_23428,N_14976,N_12771);
nor U23429 (N_23429,N_16363,N_13242);
nand U23430 (N_23430,N_12450,N_15728);
or U23431 (N_23431,N_14200,N_17872);
xor U23432 (N_23432,N_16261,N_14559);
and U23433 (N_23433,N_12961,N_16131);
nor U23434 (N_23434,N_13484,N_17725);
xor U23435 (N_23435,N_17382,N_17800);
nand U23436 (N_23436,N_17499,N_17236);
and U23437 (N_23437,N_12263,N_16903);
nand U23438 (N_23438,N_16459,N_13133);
xor U23439 (N_23439,N_17306,N_16714);
and U23440 (N_23440,N_13551,N_14109);
and U23441 (N_23441,N_15023,N_17964);
nor U23442 (N_23442,N_13841,N_14037);
xnor U23443 (N_23443,N_15363,N_16336);
xnor U23444 (N_23444,N_12610,N_13319);
and U23445 (N_23445,N_13737,N_17950);
and U23446 (N_23446,N_12886,N_12636);
and U23447 (N_23447,N_12516,N_16544);
nand U23448 (N_23448,N_13957,N_13153);
nand U23449 (N_23449,N_14359,N_13577);
nor U23450 (N_23450,N_12207,N_16409);
and U23451 (N_23451,N_12419,N_16517);
xnor U23452 (N_23452,N_14581,N_15096);
or U23453 (N_23453,N_17936,N_13327);
nand U23454 (N_23454,N_14044,N_17214);
xor U23455 (N_23455,N_14072,N_12180);
nand U23456 (N_23456,N_12394,N_15290);
and U23457 (N_23457,N_12714,N_16158);
or U23458 (N_23458,N_17050,N_13471);
nor U23459 (N_23459,N_12732,N_12975);
nand U23460 (N_23460,N_16467,N_17019);
nand U23461 (N_23461,N_13014,N_16327);
xnor U23462 (N_23462,N_12295,N_13746);
nor U23463 (N_23463,N_16149,N_16216);
nand U23464 (N_23464,N_17263,N_15149);
and U23465 (N_23465,N_16614,N_16147);
and U23466 (N_23466,N_13768,N_13688);
xnor U23467 (N_23467,N_12754,N_17272);
nor U23468 (N_23468,N_17030,N_13046);
xnor U23469 (N_23469,N_15937,N_16404);
nor U23470 (N_23470,N_14032,N_16020);
nor U23471 (N_23471,N_14160,N_12364);
nor U23472 (N_23472,N_16777,N_12346);
nor U23473 (N_23473,N_17163,N_13168);
xor U23474 (N_23474,N_17427,N_17055);
or U23475 (N_23475,N_13640,N_16518);
nand U23476 (N_23476,N_16885,N_13533);
xor U23477 (N_23477,N_13337,N_15656);
nand U23478 (N_23478,N_12765,N_14127);
nor U23479 (N_23479,N_12210,N_12524);
and U23480 (N_23480,N_12190,N_12891);
xnor U23481 (N_23481,N_14275,N_15761);
or U23482 (N_23482,N_15603,N_14662);
nand U23483 (N_23483,N_13096,N_13004);
nor U23484 (N_23484,N_16917,N_14769);
xnor U23485 (N_23485,N_15641,N_15534);
nor U23486 (N_23486,N_15295,N_13408);
nand U23487 (N_23487,N_13302,N_13042);
and U23488 (N_23488,N_12220,N_17181);
nand U23489 (N_23489,N_17653,N_16425);
or U23490 (N_23490,N_13284,N_16729);
and U23491 (N_23491,N_12535,N_12107);
xor U23492 (N_23492,N_13830,N_14224);
xor U23493 (N_23493,N_16883,N_13213);
or U23494 (N_23494,N_12506,N_15243);
nor U23495 (N_23495,N_17686,N_14809);
nor U23496 (N_23496,N_13215,N_17214);
xnor U23497 (N_23497,N_15931,N_13465);
xnor U23498 (N_23498,N_13737,N_12533);
xnor U23499 (N_23499,N_12954,N_12631);
and U23500 (N_23500,N_13706,N_13850);
xor U23501 (N_23501,N_15993,N_16117);
or U23502 (N_23502,N_17530,N_13968);
nor U23503 (N_23503,N_14559,N_17244);
and U23504 (N_23504,N_13373,N_13179);
or U23505 (N_23505,N_17432,N_13571);
xor U23506 (N_23506,N_17901,N_16307);
and U23507 (N_23507,N_17785,N_14942);
nor U23508 (N_23508,N_12862,N_15321);
or U23509 (N_23509,N_17289,N_17828);
xnor U23510 (N_23510,N_17979,N_16331);
nor U23511 (N_23511,N_13911,N_14669);
xnor U23512 (N_23512,N_15580,N_17046);
nor U23513 (N_23513,N_15586,N_17334);
and U23514 (N_23514,N_15469,N_16901);
nand U23515 (N_23515,N_17707,N_14061);
nor U23516 (N_23516,N_17579,N_15799);
and U23517 (N_23517,N_15201,N_14248);
or U23518 (N_23518,N_17077,N_15840);
xnor U23519 (N_23519,N_14309,N_12945);
and U23520 (N_23520,N_15010,N_16867);
nand U23521 (N_23521,N_15059,N_17455);
and U23522 (N_23522,N_12908,N_14579);
nand U23523 (N_23523,N_14148,N_17285);
xnor U23524 (N_23524,N_17655,N_14966);
and U23525 (N_23525,N_17579,N_12328);
nand U23526 (N_23526,N_12980,N_14607);
nor U23527 (N_23527,N_13447,N_13062);
and U23528 (N_23528,N_13506,N_16980);
and U23529 (N_23529,N_15914,N_15267);
nand U23530 (N_23530,N_12074,N_12478);
or U23531 (N_23531,N_12427,N_12748);
and U23532 (N_23532,N_12950,N_13966);
and U23533 (N_23533,N_13856,N_17146);
and U23534 (N_23534,N_12047,N_17736);
xor U23535 (N_23535,N_13426,N_15098);
or U23536 (N_23536,N_16661,N_17873);
nor U23537 (N_23537,N_16113,N_14933);
or U23538 (N_23538,N_14469,N_15943);
nand U23539 (N_23539,N_14213,N_17896);
or U23540 (N_23540,N_12493,N_17872);
nor U23541 (N_23541,N_12151,N_14508);
xor U23542 (N_23542,N_17613,N_17104);
nand U23543 (N_23543,N_13080,N_14484);
nand U23544 (N_23544,N_14397,N_17696);
nor U23545 (N_23545,N_15635,N_12821);
nor U23546 (N_23546,N_17328,N_16320);
and U23547 (N_23547,N_13700,N_15167);
xnor U23548 (N_23548,N_13541,N_13944);
nor U23549 (N_23549,N_14935,N_13671);
nor U23550 (N_23550,N_17997,N_17237);
or U23551 (N_23551,N_16317,N_16571);
xnor U23552 (N_23552,N_14193,N_15140);
nor U23553 (N_23553,N_12156,N_15686);
nand U23554 (N_23554,N_15869,N_17778);
nor U23555 (N_23555,N_14961,N_15482);
xor U23556 (N_23556,N_14739,N_17328);
nand U23557 (N_23557,N_16445,N_16821);
nor U23558 (N_23558,N_16138,N_14240);
and U23559 (N_23559,N_16840,N_16318);
xor U23560 (N_23560,N_17178,N_12009);
nor U23561 (N_23561,N_16828,N_14856);
nor U23562 (N_23562,N_12628,N_17388);
nor U23563 (N_23563,N_17855,N_17550);
and U23564 (N_23564,N_12241,N_17339);
nand U23565 (N_23565,N_14923,N_17547);
xor U23566 (N_23566,N_12731,N_14688);
and U23567 (N_23567,N_14488,N_16865);
nor U23568 (N_23568,N_16111,N_13896);
or U23569 (N_23569,N_13253,N_13920);
and U23570 (N_23570,N_15642,N_17079);
or U23571 (N_23571,N_17079,N_16343);
xnor U23572 (N_23572,N_13243,N_13329);
or U23573 (N_23573,N_17195,N_13366);
and U23574 (N_23574,N_17955,N_14476);
and U23575 (N_23575,N_13795,N_16815);
and U23576 (N_23576,N_16215,N_12361);
nor U23577 (N_23577,N_16772,N_17981);
or U23578 (N_23578,N_14117,N_13465);
nor U23579 (N_23579,N_17777,N_14004);
or U23580 (N_23580,N_12988,N_13845);
and U23581 (N_23581,N_16931,N_16984);
and U23582 (N_23582,N_12923,N_15651);
xor U23583 (N_23583,N_15021,N_16715);
xnor U23584 (N_23584,N_14490,N_13854);
or U23585 (N_23585,N_13992,N_12375);
xor U23586 (N_23586,N_14886,N_15598);
nand U23587 (N_23587,N_12239,N_15775);
nand U23588 (N_23588,N_13946,N_13574);
xnor U23589 (N_23589,N_14116,N_14371);
xnor U23590 (N_23590,N_17375,N_14289);
nand U23591 (N_23591,N_12459,N_16121);
and U23592 (N_23592,N_12811,N_12376);
nand U23593 (N_23593,N_15640,N_17861);
and U23594 (N_23594,N_12866,N_13437);
xor U23595 (N_23595,N_17305,N_13601);
and U23596 (N_23596,N_15909,N_14054);
and U23597 (N_23597,N_17048,N_12854);
nor U23598 (N_23598,N_12026,N_15616);
or U23599 (N_23599,N_15177,N_14154);
nor U23600 (N_23600,N_16436,N_13470);
and U23601 (N_23601,N_12983,N_14654);
nor U23602 (N_23602,N_17644,N_15847);
xor U23603 (N_23603,N_12502,N_13750);
nor U23604 (N_23604,N_13513,N_14913);
or U23605 (N_23605,N_16556,N_17070);
and U23606 (N_23606,N_13797,N_17210);
or U23607 (N_23607,N_12614,N_14806);
nor U23608 (N_23608,N_14237,N_15592);
and U23609 (N_23609,N_16082,N_14766);
xor U23610 (N_23610,N_14370,N_16593);
nand U23611 (N_23611,N_12169,N_17380);
and U23612 (N_23612,N_13305,N_14247);
and U23613 (N_23613,N_12073,N_16823);
nand U23614 (N_23614,N_13036,N_12644);
xnor U23615 (N_23615,N_12989,N_14065);
xnor U23616 (N_23616,N_12816,N_16417);
xor U23617 (N_23617,N_13769,N_12218);
and U23618 (N_23618,N_13962,N_12581);
or U23619 (N_23619,N_16107,N_14093);
and U23620 (N_23620,N_13797,N_14278);
xnor U23621 (N_23621,N_15017,N_13175);
nand U23622 (N_23622,N_16451,N_16733);
or U23623 (N_23623,N_13850,N_13177);
or U23624 (N_23624,N_14674,N_13830);
or U23625 (N_23625,N_13878,N_13431);
or U23626 (N_23626,N_13691,N_12690);
and U23627 (N_23627,N_15420,N_13067);
nand U23628 (N_23628,N_13043,N_16197);
nor U23629 (N_23629,N_16031,N_12538);
nor U23630 (N_23630,N_13928,N_14888);
or U23631 (N_23631,N_17546,N_16448);
nand U23632 (N_23632,N_15581,N_12423);
or U23633 (N_23633,N_12953,N_15529);
and U23634 (N_23634,N_14456,N_13062);
or U23635 (N_23635,N_15727,N_17428);
or U23636 (N_23636,N_17336,N_12586);
xnor U23637 (N_23637,N_16659,N_15516);
nand U23638 (N_23638,N_13672,N_12525);
xnor U23639 (N_23639,N_15862,N_14037);
and U23640 (N_23640,N_13942,N_17279);
nor U23641 (N_23641,N_17223,N_13033);
xor U23642 (N_23642,N_17211,N_15152);
nand U23643 (N_23643,N_16184,N_13458);
and U23644 (N_23644,N_13469,N_12821);
nand U23645 (N_23645,N_12616,N_12167);
nor U23646 (N_23646,N_13566,N_17181);
and U23647 (N_23647,N_15317,N_12664);
nor U23648 (N_23648,N_12585,N_13802);
or U23649 (N_23649,N_17174,N_12887);
nor U23650 (N_23650,N_15659,N_13235);
xor U23651 (N_23651,N_17489,N_15945);
nor U23652 (N_23652,N_17529,N_12437);
nor U23653 (N_23653,N_16871,N_14548);
nor U23654 (N_23654,N_15485,N_17344);
or U23655 (N_23655,N_16623,N_17354);
and U23656 (N_23656,N_15635,N_13610);
nor U23657 (N_23657,N_15731,N_15946);
nand U23658 (N_23658,N_16766,N_17026);
nand U23659 (N_23659,N_14731,N_14391);
nor U23660 (N_23660,N_16168,N_13789);
nand U23661 (N_23661,N_14146,N_15528);
or U23662 (N_23662,N_15710,N_13648);
nor U23663 (N_23663,N_13202,N_13988);
or U23664 (N_23664,N_17041,N_13522);
and U23665 (N_23665,N_13380,N_12303);
and U23666 (N_23666,N_13737,N_16654);
xnor U23667 (N_23667,N_13429,N_17882);
xor U23668 (N_23668,N_17745,N_17761);
or U23669 (N_23669,N_12665,N_17200);
and U23670 (N_23670,N_17375,N_17130);
xor U23671 (N_23671,N_12898,N_15213);
nor U23672 (N_23672,N_15098,N_13042);
and U23673 (N_23673,N_17904,N_13056);
xor U23674 (N_23674,N_16935,N_14567);
or U23675 (N_23675,N_15072,N_14759);
nor U23676 (N_23676,N_12597,N_17935);
and U23677 (N_23677,N_17764,N_16917);
xor U23678 (N_23678,N_12978,N_14987);
nor U23679 (N_23679,N_15952,N_12925);
xnor U23680 (N_23680,N_14123,N_17705);
or U23681 (N_23681,N_14064,N_13969);
and U23682 (N_23682,N_17903,N_12554);
nor U23683 (N_23683,N_13395,N_16537);
nor U23684 (N_23684,N_12783,N_14098);
nor U23685 (N_23685,N_17320,N_17164);
nand U23686 (N_23686,N_12355,N_15157);
or U23687 (N_23687,N_16948,N_14312);
xor U23688 (N_23688,N_15950,N_17298);
nor U23689 (N_23689,N_12027,N_17184);
nand U23690 (N_23690,N_15215,N_17939);
or U23691 (N_23691,N_12574,N_16481);
nand U23692 (N_23692,N_12659,N_13884);
nand U23693 (N_23693,N_12230,N_17381);
or U23694 (N_23694,N_14204,N_16887);
nor U23695 (N_23695,N_17558,N_15037);
nor U23696 (N_23696,N_16366,N_15843);
nand U23697 (N_23697,N_12630,N_13968);
nor U23698 (N_23698,N_13557,N_13757);
xnor U23699 (N_23699,N_17475,N_13018);
xnor U23700 (N_23700,N_16387,N_12806);
nor U23701 (N_23701,N_13733,N_17049);
or U23702 (N_23702,N_17412,N_13209);
nor U23703 (N_23703,N_16409,N_17334);
and U23704 (N_23704,N_16064,N_14082);
and U23705 (N_23705,N_12416,N_14349);
or U23706 (N_23706,N_15633,N_17033);
nor U23707 (N_23707,N_12254,N_12142);
nor U23708 (N_23708,N_13496,N_12734);
nand U23709 (N_23709,N_13669,N_12812);
and U23710 (N_23710,N_16798,N_13894);
nand U23711 (N_23711,N_15781,N_15826);
xor U23712 (N_23712,N_15658,N_16648);
and U23713 (N_23713,N_15314,N_15474);
nor U23714 (N_23714,N_15398,N_17460);
nand U23715 (N_23715,N_15243,N_17631);
xnor U23716 (N_23716,N_16061,N_17969);
or U23717 (N_23717,N_12381,N_13832);
nand U23718 (N_23718,N_13601,N_17389);
xnor U23719 (N_23719,N_14077,N_14255);
nand U23720 (N_23720,N_13852,N_17251);
nor U23721 (N_23721,N_16495,N_12236);
nor U23722 (N_23722,N_12618,N_17469);
nor U23723 (N_23723,N_15884,N_15916);
and U23724 (N_23724,N_13566,N_12350);
and U23725 (N_23725,N_14676,N_15523);
nor U23726 (N_23726,N_12348,N_14804);
nand U23727 (N_23727,N_16099,N_14551);
or U23728 (N_23728,N_17601,N_15786);
nor U23729 (N_23729,N_12054,N_16263);
nor U23730 (N_23730,N_12598,N_12177);
xor U23731 (N_23731,N_13374,N_16874);
or U23732 (N_23732,N_14977,N_16988);
nand U23733 (N_23733,N_16009,N_15632);
or U23734 (N_23734,N_13276,N_15046);
or U23735 (N_23735,N_13246,N_12765);
and U23736 (N_23736,N_15946,N_12842);
or U23737 (N_23737,N_15141,N_15826);
and U23738 (N_23738,N_14074,N_17443);
and U23739 (N_23739,N_15507,N_15301);
or U23740 (N_23740,N_16388,N_14611);
nand U23741 (N_23741,N_15108,N_17130);
nor U23742 (N_23742,N_13462,N_16251);
or U23743 (N_23743,N_14890,N_14144);
xnor U23744 (N_23744,N_14169,N_15687);
and U23745 (N_23745,N_16237,N_13100);
and U23746 (N_23746,N_17905,N_16183);
and U23747 (N_23747,N_15502,N_15848);
or U23748 (N_23748,N_17265,N_15848);
xnor U23749 (N_23749,N_16631,N_15082);
nand U23750 (N_23750,N_15641,N_12849);
nand U23751 (N_23751,N_12375,N_12001);
and U23752 (N_23752,N_16505,N_12487);
nor U23753 (N_23753,N_12805,N_16756);
nand U23754 (N_23754,N_16960,N_17115);
and U23755 (N_23755,N_13927,N_16562);
or U23756 (N_23756,N_16520,N_14637);
and U23757 (N_23757,N_14227,N_16477);
nor U23758 (N_23758,N_17725,N_12527);
or U23759 (N_23759,N_12714,N_17770);
or U23760 (N_23760,N_13843,N_15033);
and U23761 (N_23761,N_14386,N_14841);
or U23762 (N_23762,N_13765,N_15831);
or U23763 (N_23763,N_13873,N_13208);
nor U23764 (N_23764,N_15785,N_17558);
or U23765 (N_23765,N_14576,N_14541);
or U23766 (N_23766,N_12015,N_12760);
nor U23767 (N_23767,N_17684,N_15864);
or U23768 (N_23768,N_12853,N_16928);
nor U23769 (N_23769,N_17242,N_14634);
xnor U23770 (N_23770,N_12350,N_15935);
or U23771 (N_23771,N_16544,N_15049);
or U23772 (N_23772,N_17893,N_16415);
or U23773 (N_23773,N_14982,N_12278);
nand U23774 (N_23774,N_14161,N_15718);
xnor U23775 (N_23775,N_16020,N_16707);
xor U23776 (N_23776,N_14183,N_12138);
nor U23777 (N_23777,N_17057,N_12013);
or U23778 (N_23778,N_13755,N_14117);
and U23779 (N_23779,N_15373,N_14746);
nor U23780 (N_23780,N_16039,N_15472);
and U23781 (N_23781,N_12627,N_13380);
xnor U23782 (N_23782,N_14569,N_12445);
or U23783 (N_23783,N_17175,N_15644);
xnor U23784 (N_23784,N_14241,N_13462);
nor U23785 (N_23785,N_16391,N_13458);
nand U23786 (N_23786,N_12546,N_17383);
nor U23787 (N_23787,N_15117,N_13779);
and U23788 (N_23788,N_13511,N_15281);
nand U23789 (N_23789,N_16989,N_16612);
nor U23790 (N_23790,N_17868,N_17791);
nand U23791 (N_23791,N_12726,N_16661);
nand U23792 (N_23792,N_13639,N_13523);
nor U23793 (N_23793,N_13707,N_15794);
and U23794 (N_23794,N_15711,N_15391);
xor U23795 (N_23795,N_15497,N_12869);
xor U23796 (N_23796,N_15200,N_16807);
and U23797 (N_23797,N_15405,N_14127);
nand U23798 (N_23798,N_16286,N_17378);
nor U23799 (N_23799,N_13958,N_12822);
nand U23800 (N_23800,N_13170,N_12907);
and U23801 (N_23801,N_14464,N_12289);
or U23802 (N_23802,N_15280,N_15586);
and U23803 (N_23803,N_12033,N_13617);
and U23804 (N_23804,N_17825,N_14653);
or U23805 (N_23805,N_14065,N_17139);
nand U23806 (N_23806,N_16558,N_16794);
nor U23807 (N_23807,N_13668,N_12072);
nor U23808 (N_23808,N_17904,N_16193);
and U23809 (N_23809,N_13704,N_13019);
xnor U23810 (N_23810,N_12965,N_12282);
and U23811 (N_23811,N_14853,N_16292);
nor U23812 (N_23812,N_15495,N_16789);
xnor U23813 (N_23813,N_15987,N_16330);
or U23814 (N_23814,N_15743,N_12476);
or U23815 (N_23815,N_16964,N_17543);
and U23816 (N_23816,N_12588,N_15966);
xor U23817 (N_23817,N_15134,N_12939);
nor U23818 (N_23818,N_14374,N_12970);
and U23819 (N_23819,N_13802,N_16230);
nand U23820 (N_23820,N_13506,N_15249);
and U23821 (N_23821,N_17771,N_12032);
and U23822 (N_23822,N_15961,N_12250);
xnor U23823 (N_23823,N_12586,N_15478);
and U23824 (N_23824,N_14323,N_16686);
nor U23825 (N_23825,N_13315,N_14190);
nand U23826 (N_23826,N_17673,N_13682);
or U23827 (N_23827,N_13269,N_13553);
or U23828 (N_23828,N_12973,N_17580);
or U23829 (N_23829,N_17403,N_15742);
nand U23830 (N_23830,N_17195,N_17785);
and U23831 (N_23831,N_17407,N_13811);
xnor U23832 (N_23832,N_17464,N_15881);
nor U23833 (N_23833,N_16780,N_13491);
nor U23834 (N_23834,N_17568,N_12593);
and U23835 (N_23835,N_12116,N_16478);
xnor U23836 (N_23836,N_14132,N_12499);
xnor U23837 (N_23837,N_17982,N_14981);
xnor U23838 (N_23838,N_12535,N_14598);
nand U23839 (N_23839,N_17474,N_12759);
nor U23840 (N_23840,N_17769,N_14625);
and U23841 (N_23841,N_15184,N_15062);
or U23842 (N_23842,N_12764,N_14000);
nand U23843 (N_23843,N_14798,N_13772);
xnor U23844 (N_23844,N_17436,N_15290);
xor U23845 (N_23845,N_13481,N_13630);
or U23846 (N_23846,N_17765,N_15927);
nand U23847 (N_23847,N_12324,N_14806);
xor U23848 (N_23848,N_13621,N_12587);
and U23849 (N_23849,N_13507,N_16878);
nand U23850 (N_23850,N_14004,N_13226);
nor U23851 (N_23851,N_13415,N_12689);
nand U23852 (N_23852,N_12951,N_17208);
xor U23853 (N_23853,N_15568,N_12696);
xor U23854 (N_23854,N_15567,N_15739);
nand U23855 (N_23855,N_17966,N_16653);
xor U23856 (N_23856,N_17767,N_16347);
or U23857 (N_23857,N_17280,N_13479);
nor U23858 (N_23858,N_15019,N_15554);
nand U23859 (N_23859,N_16112,N_15746);
nor U23860 (N_23860,N_15614,N_16974);
or U23861 (N_23861,N_14410,N_13674);
nand U23862 (N_23862,N_13703,N_13308);
xnor U23863 (N_23863,N_15387,N_15552);
and U23864 (N_23864,N_17218,N_17005);
nor U23865 (N_23865,N_12438,N_12396);
or U23866 (N_23866,N_17163,N_13917);
xor U23867 (N_23867,N_16242,N_13508);
or U23868 (N_23868,N_15375,N_15903);
nand U23869 (N_23869,N_14559,N_13256);
nand U23870 (N_23870,N_13727,N_15581);
xor U23871 (N_23871,N_12442,N_17185);
xor U23872 (N_23872,N_13058,N_17176);
nand U23873 (N_23873,N_14181,N_16162);
and U23874 (N_23874,N_12126,N_17552);
nand U23875 (N_23875,N_16994,N_17305);
or U23876 (N_23876,N_16263,N_16578);
nand U23877 (N_23877,N_17078,N_13991);
or U23878 (N_23878,N_14494,N_15162);
or U23879 (N_23879,N_15588,N_14749);
nand U23880 (N_23880,N_17840,N_15054);
and U23881 (N_23881,N_12438,N_16928);
or U23882 (N_23882,N_17318,N_17362);
nand U23883 (N_23883,N_12154,N_17307);
xor U23884 (N_23884,N_17041,N_16355);
or U23885 (N_23885,N_17708,N_17996);
nand U23886 (N_23886,N_15440,N_14095);
nand U23887 (N_23887,N_13590,N_13179);
xnor U23888 (N_23888,N_13514,N_12642);
nand U23889 (N_23889,N_16255,N_15520);
or U23890 (N_23890,N_12119,N_16029);
nor U23891 (N_23891,N_17895,N_17583);
nor U23892 (N_23892,N_17117,N_16799);
xnor U23893 (N_23893,N_12952,N_13182);
or U23894 (N_23894,N_16954,N_12462);
xor U23895 (N_23895,N_12074,N_13891);
nand U23896 (N_23896,N_15663,N_14283);
or U23897 (N_23897,N_15045,N_12280);
xnor U23898 (N_23898,N_13772,N_17959);
or U23899 (N_23899,N_12766,N_17199);
nand U23900 (N_23900,N_15853,N_15193);
nand U23901 (N_23901,N_12684,N_15660);
xnor U23902 (N_23902,N_14467,N_17827);
or U23903 (N_23903,N_15638,N_14524);
and U23904 (N_23904,N_15225,N_14200);
xor U23905 (N_23905,N_16436,N_14409);
nand U23906 (N_23906,N_15387,N_16912);
or U23907 (N_23907,N_17079,N_13540);
nor U23908 (N_23908,N_12048,N_13938);
nand U23909 (N_23909,N_15118,N_16051);
nor U23910 (N_23910,N_15450,N_13489);
or U23911 (N_23911,N_17481,N_15698);
or U23912 (N_23912,N_14332,N_14645);
and U23913 (N_23913,N_14259,N_13541);
and U23914 (N_23914,N_17705,N_13078);
or U23915 (N_23915,N_15839,N_14705);
nor U23916 (N_23916,N_17420,N_16364);
nor U23917 (N_23917,N_14489,N_15813);
and U23918 (N_23918,N_16052,N_15140);
xnor U23919 (N_23919,N_12090,N_17861);
nor U23920 (N_23920,N_17485,N_16469);
nand U23921 (N_23921,N_16818,N_16962);
nand U23922 (N_23922,N_15359,N_16559);
or U23923 (N_23923,N_12419,N_13682);
and U23924 (N_23924,N_15897,N_16852);
xnor U23925 (N_23925,N_15887,N_15790);
or U23926 (N_23926,N_17680,N_13335);
nor U23927 (N_23927,N_14266,N_17775);
xnor U23928 (N_23928,N_16674,N_17348);
nor U23929 (N_23929,N_12420,N_12251);
or U23930 (N_23930,N_15635,N_15971);
or U23931 (N_23931,N_16850,N_13706);
xor U23932 (N_23932,N_16518,N_12586);
and U23933 (N_23933,N_16256,N_13947);
xor U23934 (N_23934,N_14183,N_12076);
and U23935 (N_23935,N_17787,N_17117);
nand U23936 (N_23936,N_13005,N_17831);
xnor U23937 (N_23937,N_13432,N_17372);
nor U23938 (N_23938,N_16811,N_14413);
xnor U23939 (N_23939,N_15496,N_15381);
xor U23940 (N_23940,N_13854,N_17210);
or U23941 (N_23941,N_14484,N_13694);
and U23942 (N_23942,N_16381,N_17863);
nand U23943 (N_23943,N_17734,N_17097);
xor U23944 (N_23944,N_16909,N_16614);
or U23945 (N_23945,N_12369,N_12932);
or U23946 (N_23946,N_12990,N_17388);
and U23947 (N_23947,N_14177,N_15909);
or U23948 (N_23948,N_16251,N_17790);
or U23949 (N_23949,N_17929,N_16650);
nand U23950 (N_23950,N_14060,N_13734);
xnor U23951 (N_23951,N_17690,N_17308);
or U23952 (N_23952,N_13867,N_12549);
or U23953 (N_23953,N_17461,N_13684);
xnor U23954 (N_23954,N_13478,N_15522);
nor U23955 (N_23955,N_16855,N_12182);
or U23956 (N_23956,N_16370,N_16899);
xor U23957 (N_23957,N_12474,N_14384);
or U23958 (N_23958,N_14040,N_17841);
nor U23959 (N_23959,N_16302,N_16149);
nand U23960 (N_23960,N_13312,N_17155);
nor U23961 (N_23961,N_13586,N_12204);
nand U23962 (N_23962,N_16168,N_12159);
nand U23963 (N_23963,N_15395,N_16790);
nor U23964 (N_23964,N_17583,N_12913);
xor U23965 (N_23965,N_13435,N_17867);
xnor U23966 (N_23966,N_17043,N_14451);
and U23967 (N_23967,N_15332,N_12173);
nand U23968 (N_23968,N_15566,N_16286);
nand U23969 (N_23969,N_13135,N_15881);
xor U23970 (N_23970,N_17105,N_12083);
xor U23971 (N_23971,N_14639,N_16775);
nand U23972 (N_23972,N_14861,N_12330);
or U23973 (N_23973,N_17760,N_12018);
xnor U23974 (N_23974,N_12139,N_12737);
xnor U23975 (N_23975,N_15701,N_13901);
nand U23976 (N_23976,N_14176,N_17075);
nor U23977 (N_23977,N_13210,N_17531);
and U23978 (N_23978,N_12384,N_17477);
nand U23979 (N_23979,N_15953,N_13753);
xor U23980 (N_23980,N_12824,N_16426);
nand U23981 (N_23981,N_16477,N_15488);
nor U23982 (N_23982,N_13192,N_14071);
or U23983 (N_23983,N_15087,N_17704);
nor U23984 (N_23984,N_12891,N_16466);
xor U23985 (N_23985,N_17939,N_12476);
xor U23986 (N_23986,N_13279,N_12286);
nor U23987 (N_23987,N_17707,N_13172);
and U23988 (N_23988,N_17457,N_14609);
nand U23989 (N_23989,N_13425,N_13063);
nand U23990 (N_23990,N_14202,N_17125);
or U23991 (N_23991,N_15367,N_15239);
nand U23992 (N_23992,N_14195,N_16512);
nor U23993 (N_23993,N_15893,N_17549);
and U23994 (N_23994,N_15674,N_12791);
nor U23995 (N_23995,N_14852,N_14290);
xnor U23996 (N_23996,N_16878,N_14624);
nand U23997 (N_23997,N_16267,N_17633);
xor U23998 (N_23998,N_12118,N_17226);
nand U23999 (N_23999,N_15317,N_17011);
xnor U24000 (N_24000,N_19806,N_23423);
nand U24001 (N_24001,N_21536,N_22309);
and U24002 (N_24002,N_19810,N_21880);
nand U24003 (N_24003,N_21455,N_20755);
and U24004 (N_24004,N_21177,N_22680);
xnor U24005 (N_24005,N_23112,N_20730);
or U24006 (N_24006,N_22209,N_20861);
nor U24007 (N_24007,N_19306,N_23122);
or U24008 (N_24008,N_23509,N_21261);
xor U24009 (N_24009,N_19857,N_19072);
or U24010 (N_24010,N_22946,N_22546);
nor U24011 (N_24011,N_23125,N_23272);
nand U24012 (N_24012,N_19916,N_22390);
nand U24013 (N_24013,N_19530,N_22374);
and U24014 (N_24014,N_19025,N_21319);
xnor U24015 (N_24015,N_21675,N_20920);
nand U24016 (N_24016,N_22221,N_18972);
or U24017 (N_24017,N_23073,N_22692);
nor U24018 (N_24018,N_23088,N_20814);
or U24019 (N_24019,N_22564,N_21890);
and U24020 (N_24020,N_18005,N_19574);
or U24021 (N_24021,N_22170,N_23761);
nor U24022 (N_24022,N_19187,N_19179);
nand U24023 (N_24023,N_22869,N_19561);
nand U24024 (N_24024,N_20988,N_20830);
nor U24025 (N_24025,N_19040,N_21271);
xnor U24026 (N_24026,N_22046,N_20364);
or U24027 (N_24027,N_20515,N_23180);
and U24028 (N_24028,N_22882,N_20202);
xor U24029 (N_24029,N_18224,N_23139);
nor U24030 (N_24030,N_18455,N_21649);
or U24031 (N_24031,N_20622,N_20062);
or U24032 (N_24032,N_19017,N_23947);
or U24033 (N_24033,N_21673,N_23358);
nand U24034 (N_24034,N_19816,N_21564);
or U24035 (N_24035,N_19153,N_19499);
nand U24036 (N_24036,N_19336,N_23254);
nor U24037 (N_24037,N_19411,N_21907);
or U24038 (N_24038,N_21061,N_22833);
and U24039 (N_24039,N_21566,N_22240);
nand U24040 (N_24040,N_21069,N_20793);
xnor U24041 (N_24041,N_21705,N_20575);
xnor U24042 (N_24042,N_19898,N_21137);
nand U24043 (N_24043,N_19844,N_18017);
or U24044 (N_24044,N_19679,N_19964);
xnor U24045 (N_24045,N_20758,N_21243);
and U24046 (N_24046,N_19947,N_18195);
or U24047 (N_24047,N_23937,N_20632);
nand U24048 (N_24048,N_18174,N_23347);
and U24049 (N_24049,N_18469,N_22455);
or U24050 (N_24050,N_20293,N_19963);
nor U24051 (N_24051,N_22536,N_21016);
xor U24052 (N_24052,N_19569,N_23703);
and U24053 (N_24053,N_19211,N_20578);
nand U24054 (N_24054,N_20907,N_21959);
nand U24055 (N_24055,N_19297,N_23051);
nor U24056 (N_24056,N_21173,N_23827);
xnor U24057 (N_24057,N_22395,N_19827);
xnor U24058 (N_24058,N_23202,N_21635);
xor U24059 (N_24059,N_22207,N_19647);
and U24060 (N_24060,N_23666,N_23571);
nor U24061 (N_24061,N_22949,N_23265);
nand U24062 (N_24062,N_19912,N_21923);
and U24063 (N_24063,N_18205,N_21614);
nand U24064 (N_24064,N_21236,N_18103);
or U24065 (N_24065,N_23374,N_23094);
nor U24066 (N_24066,N_19973,N_21870);
or U24067 (N_24067,N_20156,N_18733);
nand U24068 (N_24068,N_18593,N_19609);
nor U24069 (N_24069,N_21134,N_20876);
nand U24070 (N_24070,N_22615,N_22573);
xor U24071 (N_24071,N_22785,N_18487);
nand U24072 (N_24072,N_18098,N_18441);
nor U24073 (N_24073,N_19730,N_19502);
and U24074 (N_24074,N_19444,N_22172);
or U24075 (N_24075,N_19497,N_20948);
nand U24076 (N_24076,N_22270,N_18875);
or U24077 (N_24077,N_18340,N_22657);
nand U24078 (N_24078,N_19261,N_20238);
nand U24079 (N_24079,N_21706,N_23917);
nor U24080 (N_24080,N_21035,N_23205);
or U24081 (N_24081,N_23054,N_21715);
or U24082 (N_24082,N_23880,N_19624);
or U24083 (N_24083,N_18400,N_22154);
and U24084 (N_24084,N_21252,N_23999);
xor U24085 (N_24085,N_21485,N_22348);
and U24086 (N_24086,N_21508,N_19450);
nor U24087 (N_24087,N_23941,N_20648);
and U24088 (N_24088,N_21884,N_20250);
or U24089 (N_24089,N_23206,N_21553);
nor U24090 (N_24090,N_19314,N_18414);
nor U24091 (N_24091,N_19426,N_21579);
nand U24092 (N_24092,N_21938,N_20174);
and U24093 (N_24093,N_22089,N_23842);
nor U24094 (N_24094,N_19889,N_21151);
nand U24095 (N_24095,N_20408,N_22444);
and U24096 (N_24096,N_21644,N_22503);
nand U24097 (N_24097,N_19563,N_20034);
and U24098 (N_24098,N_21217,N_18659);
xnor U24099 (N_24099,N_19068,N_21431);
nor U24100 (N_24100,N_20474,N_18442);
nand U24101 (N_24101,N_21707,N_23150);
xor U24102 (N_24102,N_18906,N_22721);
nand U24103 (N_24103,N_23533,N_23126);
nand U24104 (N_24104,N_19553,N_18988);
or U24105 (N_24105,N_18268,N_22386);
and U24106 (N_24106,N_19071,N_21053);
or U24107 (N_24107,N_23969,N_21269);
or U24108 (N_24108,N_18001,N_18927);
or U24109 (N_24109,N_21459,N_22838);
or U24110 (N_24110,N_20136,N_18585);
and U24111 (N_24111,N_23096,N_20239);
xor U24112 (N_24112,N_18996,N_20232);
xor U24113 (N_24113,N_21500,N_23497);
and U24114 (N_24114,N_19505,N_18355);
nor U24115 (N_24115,N_19724,N_22187);
nand U24116 (N_24116,N_18373,N_21648);
nand U24117 (N_24117,N_20801,N_18130);
or U24118 (N_24118,N_18405,N_19155);
nand U24119 (N_24119,N_23047,N_20946);
and U24120 (N_24120,N_22191,N_22350);
xnor U24121 (N_24121,N_23040,N_18738);
and U24122 (N_24122,N_23671,N_18903);
and U24123 (N_24123,N_21031,N_21462);
and U24124 (N_24124,N_20764,N_20373);
nor U24125 (N_24125,N_19169,N_20874);
nand U24126 (N_24126,N_18257,N_21495);
xnor U24127 (N_24127,N_19494,N_22610);
xnor U24128 (N_24128,N_20199,N_18770);
xnor U24129 (N_24129,N_21121,N_23199);
xnor U24130 (N_24130,N_23894,N_22658);
nand U24131 (N_24131,N_22550,N_21781);
nand U24132 (N_24132,N_23219,N_20012);
and U24133 (N_24133,N_23567,N_23460);
xnor U24134 (N_24134,N_18795,N_20669);
xnor U24135 (N_24135,N_23481,N_23344);
and U24136 (N_24136,N_20840,N_21468);
xnor U24137 (N_24137,N_21384,N_21279);
or U24138 (N_24138,N_22320,N_23997);
nand U24139 (N_24139,N_18311,N_20165);
xor U24140 (N_24140,N_23470,N_18870);
nor U24141 (N_24141,N_21244,N_18682);
nor U24142 (N_24142,N_23617,N_21539);
xnor U24143 (N_24143,N_18681,N_21913);
and U24144 (N_24144,N_22488,N_19231);
nor U24145 (N_24145,N_19214,N_22160);
nand U24146 (N_24146,N_20898,N_21807);
xnor U24147 (N_24147,N_22813,N_23298);
and U24148 (N_24148,N_23149,N_20391);
and U24149 (N_24149,N_18486,N_19202);
nor U24150 (N_24150,N_23644,N_21258);
and U24151 (N_24151,N_22644,N_23992);
or U24152 (N_24152,N_22566,N_22719);
or U24153 (N_24153,N_20548,N_19802);
and U24154 (N_24154,N_18356,N_19055);
nand U24155 (N_24155,N_19037,N_19051);
and U24156 (N_24156,N_18489,N_23756);
nand U24157 (N_24157,N_22186,N_20301);
or U24158 (N_24158,N_19510,N_21247);
nor U24159 (N_24159,N_23142,N_21795);
xor U24160 (N_24160,N_20828,N_20997);
xor U24161 (N_24161,N_23170,N_21803);
nor U24162 (N_24162,N_19937,N_22865);
and U24163 (N_24163,N_18668,N_19390);
nor U24164 (N_24164,N_23609,N_23258);
nor U24165 (N_24165,N_19078,N_21792);
xnor U24166 (N_24166,N_18891,N_22297);
nor U24167 (N_24167,N_19999,N_21902);
nand U24168 (N_24168,N_18346,N_20978);
and U24169 (N_24169,N_22327,N_21710);
and U24170 (N_24170,N_20502,N_20075);
nand U24171 (N_24171,N_23608,N_19812);
and U24172 (N_24172,N_18705,N_23758);
xnor U24173 (N_24173,N_20722,N_21680);
nor U24174 (N_24174,N_21263,N_23817);
nand U24175 (N_24175,N_23314,N_18791);
nand U24176 (N_24176,N_21514,N_21526);
nor U24177 (N_24177,N_18690,N_21272);
and U24178 (N_24178,N_21313,N_20172);
nand U24179 (N_24179,N_22183,N_22913);
nor U24180 (N_24180,N_23920,N_22323);
nand U24181 (N_24181,N_23572,N_20141);
nor U24182 (N_24182,N_19992,N_20124);
xor U24183 (N_24183,N_18408,N_21481);
xnor U24184 (N_24184,N_21740,N_21989);
xnor U24185 (N_24185,N_22013,N_22747);
xnor U24186 (N_24186,N_21749,N_18986);
nand U24187 (N_24187,N_22391,N_22963);
or U24188 (N_24188,N_18748,N_22756);
nand U24189 (N_24189,N_21647,N_22370);
nand U24190 (N_24190,N_23841,N_18097);
and U24191 (N_24191,N_18712,N_20573);
nand U24192 (N_24192,N_21062,N_19642);
nor U24193 (N_24193,N_18104,N_22019);
nand U24194 (N_24194,N_19566,N_22858);
nand U24195 (N_24195,N_21360,N_19330);
or U24196 (N_24196,N_18815,N_23673);
xnor U24197 (N_24197,N_19950,N_21419);
nor U24198 (N_24198,N_18888,N_20719);
xor U24199 (N_24199,N_20393,N_22804);
nor U24200 (N_24200,N_18350,N_19601);
nor U24201 (N_24201,N_23591,N_19462);
xor U24202 (N_24202,N_23006,N_19075);
nor U24203 (N_24203,N_21797,N_21717);
and U24204 (N_24204,N_21947,N_18561);
and U24205 (N_24205,N_18573,N_21399);
nor U24206 (N_24206,N_22956,N_22164);
and U24207 (N_24207,N_19678,N_23251);
xor U24208 (N_24208,N_22333,N_21697);
or U24209 (N_24209,N_19392,N_22402);
nand U24210 (N_24210,N_20045,N_19033);
nor U24211 (N_24211,N_18380,N_22159);
and U24212 (N_24212,N_19855,N_20128);
nand U24213 (N_24213,N_22773,N_20712);
xnor U24214 (N_24214,N_21070,N_20101);
nor U24215 (N_24215,N_20973,N_19456);
nand U24216 (N_24216,N_22577,N_18566);
nand U24217 (N_24217,N_18364,N_18994);
nor U24218 (N_24218,N_20409,N_18899);
or U24219 (N_24219,N_22096,N_19757);
or U24220 (N_24220,N_19098,N_22472);
and U24221 (N_24221,N_18691,N_18204);
and U24222 (N_24222,N_18417,N_23773);
nand U24223 (N_24223,N_18190,N_20964);
nor U24224 (N_24224,N_22372,N_19317);
xor U24225 (N_24225,N_21837,N_22733);
and U24226 (N_24226,N_19848,N_18043);
nand U24227 (N_24227,N_23027,N_22881);
xor U24228 (N_24228,N_21701,N_18855);
and U24229 (N_24229,N_23410,N_21420);
and U24230 (N_24230,N_23132,N_19175);
xor U24231 (N_24231,N_19209,N_23988);
and U24232 (N_24232,N_20646,N_18175);
xor U24233 (N_24233,N_21354,N_20475);
or U24234 (N_24234,N_23975,N_19759);
nand U24235 (N_24235,N_21527,N_20899);
nor U24236 (N_24236,N_22912,N_22421);
nor U24237 (N_24237,N_20201,N_22490);
or U24238 (N_24238,N_22245,N_23475);
and U24239 (N_24239,N_23085,N_23267);
nand U24240 (N_24240,N_21371,N_22722);
nand U24241 (N_24241,N_18032,N_18019);
nand U24242 (N_24242,N_23377,N_18166);
xnor U24243 (N_24243,N_18030,N_18153);
or U24244 (N_24244,N_18020,N_19644);
nor U24245 (N_24245,N_20659,N_20883);
or U24246 (N_24246,N_19993,N_19027);
nor U24247 (N_24247,N_21733,N_18950);
and U24248 (N_24248,N_19005,N_20927);
nor U24249 (N_24249,N_18272,N_19259);
or U24250 (N_24250,N_20950,N_23906);
xnor U24251 (N_24251,N_18128,N_21366);
or U24252 (N_24252,N_22924,N_21568);
xnor U24253 (N_24253,N_19804,N_19268);
nor U24254 (N_24254,N_19448,N_21873);
or U24255 (N_24255,N_18299,N_21201);
or U24256 (N_24256,N_21197,N_20461);
and U24257 (N_24257,N_18660,N_19092);
and U24258 (N_24258,N_19953,N_21861);
xor U24259 (N_24259,N_19171,N_20564);
nand U24260 (N_24260,N_18079,N_18471);
xnor U24261 (N_24261,N_19064,N_20778);
and U24262 (N_24262,N_19221,N_23456);
and U24263 (N_24263,N_23484,N_23425);
and U24264 (N_24264,N_21406,N_19754);
nand U24265 (N_24265,N_20647,N_23434);
nand U24266 (N_24266,N_19349,N_18133);
and U24267 (N_24267,N_18995,N_23165);
or U24268 (N_24268,N_18510,N_22492);
or U24269 (N_24269,N_19486,N_22015);
and U24270 (N_24270,N_23158,N_18752);
and U24271 (N_24271,N_21392,N_23315);
nand U24272 (N_24272,N_19913,N_20425);
or U24273 (N_24273,N_19861,N_21007);
nor U24274 (N_24274,N_23637,N_19696);
nand U24275 (N_24275,N_23127,N_21698);
nor U24276 (N_24276,N_18285,N_18431);
xor U24277 (N_24277,N_22887,N_18597);
nor U24278 (N_24278,N_23858,N_21628);
nor U24279 (N_24279,N_21932,N_21933);
and U24280 (N_24280,N_18035,N_21941);
xnor U24281 (N_24281,N_23035,N_21897);
and U24282 (N_24282,N_20923,N_21067);
and U24283 (N_24283,N_18794,N_19047);
and U24284 (N_24284,N_23411,N_20015);
xor U24285 (N_24285,N_21556,N_20493);
and U24286 (N_24286,N_20765,N_18689);
or U24287 (N_24287,N_22636,N_18251);
nand U24288 (N_24288,N_20077,N_18416);
nor U24289 (N_24289,N_21223,N_20057);
and U24290 (N_24290,N_22802,N_20256);
and U24291 (N_24291,N_18067,N_21856);
xor U24292 (N_24292,N_23722,N_20476);
or U24293 (N_24293,N_20346,N_20565);
nand U24294 (N_24294,N_23683,N_21091);
xnor U24295 (N_24295,N_19032,N_18173);
nor U24296 (N_24296,N_20970,N_20139);
and U24297 (N_24297,N_18762,N_22378);
nor U24298 (N_24298,N_21616,N_20686);
xnor U24299 (N_24299,N_21100,N_19252);
and U24300 (N_24300,N_23734,N_20234);
or U24301 (N_24301,N_22620,N_18812);
or U24302 (N_24302,N_23688,N_20951);
xnor U24303 (N_24303,N_23657,N_20741);
nor U24304 (N_24304,N_19764,N_22583);
or U24305 (N_24305,N_21809,N_20772);
or U24306 (N_24306,N_22548,N_23083);
nand U24307 (N_24307,N_19255,N_18858);
xnor U24308 (N_24308,N_18223,N_21828);
nor U24309 (N_24309,N_23565,N_19034);
nor U24310 (N_24310,N_22587,N_19132);
or U24311 (N_24311,N_23919,N_23925);
nor U24312 (N_24312,N_23828,N_18367);
nor U24313 (N_24313,N_18277,N_21674);
nor U24314 (N_24314,N_20246,N_23432);
and U24315 (N_24315,N_20248,N_22398);
nor U24316 (N_24316,N_22124,N_22764);
or U24317 (N_24317,N_21569,N_23412);
nand U24318 (N_24318,N_22000,N_21445);
nor U24319 (N_24319,N_18436,N_19215);
nor U24320 (N_24320,N_22695,N_19024);
nand U24321 (N_24321,N_22334,N_19781);
and U24322 (N_24322,N_23524,N_20300);
nand U24323 (N_24323,N_18298,N_18160);
nand U24324 (N_24324,N_20842,N_22415);
or U24325 (N_24325,N_20760,N_20415);
nor U24326 (N_24326,N_23469,N_23763);
or U24327 (N_24327,N_18341,N_20630);
nor U24328 (N_24328,N_19290,N_23217);
or U24329 (N_24329,N_22414,N_19083);
and U24330 (N_24330,N_22338,N_21024);
and U24331 (N_24331,N_23620,N_18241);
nand U24332 (N_24332,N_20167,N_22222);
nand U24333 (N_24333,N_23564,N_18640);
nand U24334 (N_24334,N_23901,N_20553);
xnor U24335 (N_24335,N_21582,N_20266);
xor U24336 (N_24336,N_22387,N_20386);
xnor U24337 (N_24337,N_18558,N_21713);
nand U24338 (N_24338,N_20452,N_21138);
and U24339 (N_24339,N_23596,N_23653);
and U24340 (N_24340,N_20921,N_21704);
nor U24341 (N_24341,N_22770,N_20517);
nor U24342 (N_24342,N_18283,N_18799);
xnor U24343 (N_24343,N_23812,N_19395);
or U24344 (N_24344,N_20429,N_18465);
nor U24345 (N_24345,N_23339,N_20473);
nand U24346 (N_24346,N_22941,N_20990);
or U24347 (N_24347,N_22317,N_20032);
xor U24348 (N_24348,N_21280,N_22246);
and U24349 (N_24349,N_18866,N_21490);
nand U24350 (N_24350,N_21023,N_22382);
or U24351 (N_24351,N_20982,N_22758);
and U24352 (N_24352,N_21824,N_18650);
and U24353 (N_24353,N_18523,N_23686);
nand U24354 (N_24354,N_23197,N_20091);
xor U24355 (N_24355,N_22273,N_21022);
nor U24356 (N_24356,N_20699,N_20694);
or U24357 (N_24357,N_19639,N_19906);
nor U24358 (N_24358,N_19608,N_20210);
xor U24359 (N_24359,N_21469,N_22759);
and U24360 (N_24360,N_22847,N_18096);
and U24361 (N_24361,N_20785,N_18915);
and U24362 (N_24362,N_19895,N_19551);
or U24363 (N_24363,N_21990,N_19659);
and U24364 (N_24364,N_19596,N_18813);
nor U24365 (N_24365,N_22094,N_23635);
nor U24366 (N_24366,N_19968,N_20086);
nand U24367 (N_24367,N_18049,N_23874);
or U24368 (N_24368,N_21779,N_20866);
and U24369 (N_24369,N_19399,N_21182);
nor U24370 (N_24370,N_19925,N_19449);
xnor U24371 (N_24371,N_19847,N_20198);
or U24372 (N_24372,N_22741,N_20370);
nor U24373 (N_24373,N_23077,N_22675);
xor U24374 (N_24374,N_22039,N_20454);
and U24375 (N_24375,N_20017,N_22040);
and U24376 (N_24376,N_23513,N_21098);
nor U24377 (N_24377,N_18165,N_23859);
nor U24378 (N_24378,N_18804,N_23923);
or U24379 (N_24379,N_21551,N_22713);
nor U24380 (N_24380,N_20311,N_23805);
xor U24381 (N_24381,N_19875,N_22362);
nor U24382 (N_24382,N_21814,N_18765);
and U24383 (N_24383,N_19790,N_18628);
nand U24384 (N_24384,N_22903,N_20912);
nor U24385 (N_24385,N_19996,N_19763);
or U24386 (N_24386,N_18232,N_18075);
nand U24387 (N_24387,N_19287,N_18832);
nand U24388 (N_24388,N_22514,N_18699);
xnor U24389 (N_24389,N_22939,N_21865);
or U24390 (N_24390,N_23560,N_18540);
xnor U24391 (N_24391,N_23806,N_18222);
and U24392 (N_24392,N_18100,N_18594);
xnor U24393 (N_24393,N_19514,N_20120);
or U24394 (N_24394,N_21337,N_20931);
and U24395 (N_24395,N_22210,N_23733);
xor U24396 (N_24396,N_20689,N_18099);
and U24397 (N_24397,N_22617,N_19272);
xor U24398 (N_24398,N_21358,N_18530);
nand U24399 (N_24399,N_18537,N_21850);
nor U24400 (N_24400,N_20316,N_23575);
nor U24401 (N_24401,N_21175,N_19203);
xor U24402 (N_24402,N_20222,N_23863);
nor U24403 (N_24403,N_19195,N_20320);
or U24404 (N_24404,N_23636,N_20860);
nor U24405 (N_24405,N_20835,N_20598);
nand U24406 (N_24406,N_20439,N_20225);
and U24407 (N_24407,N_18239,N_23607);
nand U24408 (N_24408,N_22163,N_20549);
nor U24409 (N_24409,N_18315,N_22064);
or U24410 (N_24410,N_19674,N_23129);
nor U24411 (N_24411,N_19910,N_18830);
nor U24412 (N_24412,N_19531,N_22888);
nand U24413 (N_24413,N_22753,N_22959);
and U24414 (N_24414,N_22034,N_23599);
or U24415 (N_24415,N_19304,N_22641);
and U24416 (N_24416,N_20154,N_19970);
nor U24417 (N_24417,N_22237,N_23514);
xnor U24418 (N_24418,N_21216,N_21922);
xnor U24419 (N_24419,N_21590,N_22581);
xnor U24420 (N_24420,N_18621,N_19637);
nor U24421 (N_24421,N_18039,N_19533);
nor U24422 (N_24422,N_19124,N_22408);
nor U24423 (N_24423,N_20112,N_23273);
xnor U24424 (N_24424,N_22346,N_20420);
nor U24425 (N_24425,N_19247,N_23566);
nand U24426 (N_24426,N_21557,N_20371);
xor U24427 (N_24427,N_18737,N_22679);
nor U24428 (N_24428,N_20902,N_21924);
or U24429 (N_24429,N_19156,N_19664);
xor U24430 (N_24430,N_20639,N_18494);
nor U24431 (N_24431,N_18665,N_22475);
nand U24432 (N_24432,N_19059,N_22556);
xor U24433 (N_24433,N_19382,N_18088);
nand U24434 (N_24434,N_22467,N_22557);
or U24435 (N_24435,N_22003,N_18159);
nand U24436 (N_24436,N_20466,N_18884);
and U24437 (N_24437,N_22216,N_20875);
or U24438 (N_24438,N_19159,N_23612);
or U24439 (N_24439,N_19424,N_22481);
or U24440 (N_24440,N_18894,N_19779);
or U24441 (N_24441,N_19481,N_21535);
nand U24442 (N_24442,N_23355,N_21344);
xor U24443 (N_24443,N_23264,N_19492);
or U24444 (N_24444,N_23690,N_20271);
nand U24445 (N_24445,N_19962,N_23252);
nor U24446 (N_24446,N_22302,N_19309);
xor U24447 (N_24447,N_20286,N_20710);
nand U24448 (N_24448,N_21544,N_22194);
nor U24449 (N_24449,N_23046,N_21726);
xnor U24450 (N_24450,N_23134,N_23577);
and U24451 (N_24451,N_19325,N_23697);
nand U24452 (N_24452,N_23606,N_19630);
and U24453 (N_24453,N_22079,N_21802);
and U24454 (N_24454,N_20367,N_22950);
and U24455 (N_24455,N_18507,N_21405);
or U24456 (N_24456,N_19008,N_22528);
or U24457 (N_24457,N_22706,N_18521);
xnor U24458 (N_24458,N_22545,N_18238);
xor U24459 (N_24459,N_18536,N_20688);
or U24460 (N_24460,N_22182,N_20538);
or U24461 (N_24461,N_21058,N_20093);
nor U24462 (N_24462,N_19969,N_21593);
xnor U24463 (N_24463,N_20497,N_19625);
nand U24464 (N_24464,N_18983,N_20609);
xnor U24465 (N_24465,N_21039,N_21096);
xnor U24466 (N_24466,N_22099,N_22397);
and U24467 (N_24467,N_20095,N_21855);
and U24468 (N_24468,N_23101,N_20520);
nand U24469 (N_24469,N_20240,N_21187);
and U24470 (N_24470,N_18267,N_22884);
and U24471 (N_24471,N_21686,N_23752);
or U24472 (N_24472,N_18955,N_21532);
or U24473 (N_24473,N_18513,N_23154);
xnor U24474 (N_24474,N_20580,N_18393);
or U24475 (N_24475,N_20733,N_19073);
xor U24476 (N_24476,N_19603,N_23965);
or U24477 (N_24477,N_23926,N_18047);
or U24478 (N_24478,N_21831,N_18289);
or U24479 (N_24479,N_22144,N_22697);
nor U24480 (N_24480,N_22591,N_20941);
nand U24481 (N_24481,N_19599,N_19157);
and U24482 (N_24482,N_22749,N_22523);
nand U24483 (N_24483,N_19076,N_20011);
nand U24484 (N_24484,N_20711,N_19543);
nor U24485 (N_24485,N_21677,N_19415);
or U24486 (N_24486,N_19717,N_22872);
nor U24487 (N_24487,N_21885,N_19578);
nor U24488 (N_24488,N_21631,N_21194);
or U24489 (N_24489,N_18898,N_21832);
and U24490 (N_24490,N_21038,N_20255);
nand U24491 (N_24491,N_18822,N_22890);
or U24492 (N_24492,N_18674,N_22150);
and U24493 (N_24493,N_20662,N_19355);
or U24494 (N_24494,N_19108,N_19589);
nand U24495 (N_24495,N_19504,N_21232);
xor U24496 (N_24496,N_23024,N_19134);
or U24497 (N_24497,N_20306,N_18270);
xnor U24498 (N_24498,N_18951,N_20972);
xor U24499 (N_24499,N_18136,N_21460);
nor U24500 (N_24500,N_19170,N_20030);
nand U24501 (N_24501,N_23285,N_22988);
nor U24502 (N_24502,N_21492,N_21926);
and U24503 (N_24503,N_23266,N_20910);
and U24504 (N_24504,N_19769,N_18422);
nand U24505 (N_24505,N_22707,N_18716);
and U24506 (N_24506,N_22930,N_21574);
xnor U24507 (N_24507,N_18004,N_23098);
nor U24508 (N_24508,N_21268,N_21391);
or U24509 (N_24509,N_18549,N_19516);
nor U24510 (N_24510,N_19918,N_20361);
and U24511 (N_24511,N_21013,N_20228);
and U24512 (N_24512,N_23297,N_21109);
or U24513 (N_24513,N_21872,N_18745);
xor U24514 (N_24514,N_20696,N_22471);
and U24515 (N_24515,N_19522,N_22968);
and U24516 (N_24516,N_18488,N_21424);
nand U24517 (N_24517,N_19727,N_19740);
nor U24518 (N_24518,N_19508,N_18933);
and U24519 (N_24519,N_18724,N_20004);
or U24520 (N_24520,N_23507,N_18491);
and U24521 (N_24521,N_18252,N_19461);
nand U24522 (N_24522,N_20365,N_18811);
nand U24523 (N_24523,N_19267,N_19663);
nand U24524 (N_24524,N_18755,N_19229);
nand U24525 (N_24525,N_20612,N_22354);
nand U24526 (N_24526,N_21484,N_19432);
nand U24527 (N_24527,N_23232,N_20060);
nand U24528 (N_24528,N_22752,N_18118);
nor U24529 (N_24529,N_21606,N_20080);
or U24530 (N_24530,N_23472,N_22037);
nor U24531 (N_24531,N_21470,N_22321);
xnor U24532 (N_24532,N_22105,N_21168);
or U24533 (N_24533,N_18661,N_19666);
nor U24534 (N_24534,N_19319,N_21835);
nor U24535 (N_24535,N_18102,N_22050);
nand U24536 (N_24536,N_22519,N_21008);
or U24537 (N_24537,N_18575,N_21754);
and U24538 (N_24538,N_21122,N_19859);
or U24539 (N_24539,N_23595,N_22628);
nand U24540 (N_24540,N_19271,N_22477);
and U24541 (N_24541,N_18146,N_20945);
nor U24542 (N_24542,N_19286,N_22824);
nor U24543 (N_24543,N_23240,N_19417);
nand U24544 (N_24544,N_19782,N_22148);
or U24545 (N_24545,N_22329,N_23921);
nand U24546 (N_24546,N_19243,N_19837);
nand U24547 (N_24547,N_22727,N_20302);
or U24548 (N_24548,N_20241,N_21956);
xnor U24549 (N_24549,N_23585,N_20868);
and U24550 (N_24550,N_19021,N_22268);
or U24551 (N_24551,N_19590,N_18135);
and U24552 (N_24552,N_18619,N_19586);
xnor U24553 (N_24553,N_18259,N_18715);
and U24554 (N_24554,N_18332,N_18505);
nand U24555 (N_24555,N_18610,N_20818);
and U24556 (N_24556,N_23646,N_23530);
and U24557 (N_24557,N_19423,N_22718);
nor U24558 (N_24558,N_19090,N_19705);
or U24559 (N_24559,N_18750,N_20108);
or U24560 (N_24560,N_22894,N_22554);
or U24561 (N_24561,N_18763,N_20752);
xor U24562 (N_24562,N_22817,N_19154);
nor U24563 (N_24563,N_18424,N_22025);
or U24564 (N_24564,N_19052,N_20288);
xor U24565 (N_24565,N_20066,N_22112);
xor U24566 (N_24566,N_18514,N_23891);
xor U24567 (N_24567,N_21295,N_18688);
nor U24568 (N_24568,N_19206,N_20656);
or U24569 (N_24569,N_23754,N_22982);
xor U24570 (N_24570,N_20267,N_23043);
xnor U24571 (N_24571,N_23225,N_21050);
nand U24572 (N_24572,N_23723,N_22134);
nand U24573 (N_24573,N_23028,N_22388);
and U24574 (N_24574,N_18700,N_23457);
or U24575 (N_24575,N_22765,N_21165);
and U24576 (N_24576,N_19016,N_22137);
nand U24577 (N_24577,N_18461,N_20747);
or U24578 (N_24578,N_22337,N_18717);
nand U24579 (N_24579,N_20102,N_22505);
nor U24580 (N_24580,N_20703,N_21571);
and U24581 (N_24581,N_23562,N_18145);
nand U24582 (N_24582,N_19568,N_20928);
xnor U24583 (N_24583,N_22960,N_20099);
nor U24584 (N_24584,N_21374,N_23584);
nand U24585 (N_24585,N_19095,N_18913);
and U24586 (N_24586,N_23537,N_22673);
xnor U24587 (N_24587,N_23319,N_23067);
nand U24588 (N_24588,N_19184,N_20725);
or U24589 (N_24589,N_21825,N_23550);
xnor U24590 (N_24590,N_22742,N_21901);
nor U24591 (N_24591,N_20519,N_22189);
or U24592 (N_24592,N_22531,N_20322);
nand U24593 (N_24593,N_22811,N_22107);
nor U24594 (N_24594,N_22132,N_23654);
and U24595 (N_24595,N_23549,N_18565);
and U24596 (N_24596,N_18654,N_19610);
xnor U24597 (N_24597,N_21104,N_22592);
nand U24598 (N_24598,N_18821,N_23415);
xnor U24599 (N_24599,N_22147,N_21477);
nand U24600 (N_24600,N_21962,N_23304);
or U24601 (N_24601,N_22355,N_21979);
xor U24602 (N_24602,N_18864,N_18111);
xnor U24603 (N_24603,N_21141,N_21401);
xor U24604 (N_24604,N_18977,N_19189);
xnor U24605 (N_24605,N_19220,N_23176);
or U24606 (N_24606,N_21145,N_21410);
and U24607 (N_24607,N_19793,N_18378);
or U24608 (N_24608,N_23201,N_18900);
and U24609 (N_24609,N_21306,N_23075);
nor U24610 (N_24610,N_19941,N_19629);
nor U24611 (N_24611,N_20446,N_20433);
or U24612 (N_24612,N_21845,N_22702);
nor U24613 (N_24613,N_21474,N_18788);
nand U24614 (N_24614,N_21597,N_20394);
and U24615 (N_24615,N_23007,N_18759);
and U24616 (N_24616,N_18194,N_23463);
nand U24617 (N_24617,N_20372,N_23797);
nand U24618 (N_24618,N_19117,N_18493);
xnor U24619 (N_24619,N_20533,N_18313);
nand U24620 (N_24620,N_23869,N_19796);
xor U24621 (N_24621,N_20588,N_22624);
xnor U24622 (N_24622,N_19275,N_18630);
nor U24623 (N_24623,N_23243,N_22938);
xnor U24624 (N_24624,N_23402,N_19658);
and U24625 (N_24625,N_21382,N_19560);
or U24626 (N_24626,N_18182,N_19633);
nand U24627 (N_24627,N_23709,N_21842);
nand U24628 (N_24628,N_18632,N_19147);
xnor U24629 (N_24629,N_19833,N_22358);
nor U24630 (N_24630,N_18749,N_21620);
xnor U24631 (N_24631,N_20697,N_23451);
nand U24632 (N_24632,N_20449,N_18844);
nand U24633 (N_24633,N_20282,N_19832);
nand U24634 (N_24634,N_23229,N_23640);
nor U24635 (N_24635,N_21504,N_22940);
nand U24636 (N_24636,N_22463,N_21523);
nor U24637 (N_24637,N_19413,N_21278);
nor U24638 (N_24638,N_19246,N_18389);
nand U24639 (N_24639,N_20081,N_20059);
nor U24640 (N_24640,N_22409,N_18263);
and U24641 (N_24641,N_23548,N_21747);
nor U24642 (N_24642,N_20559,N_21622);
or U24643 (N_24643,N_22818,N_18848);
and U24644 (N_24644,N_23799,N_19123);
nor U24645 (N_24645,N_21284,N_19784);
xor U24646 (N_24646,N_19028,N_21136);
nor U24647 (N_24647,N_19538,N_18533);
xor U24648 (N_24648,N_22954,N_20016);
and U24649 (N_24649,N_19116,N_22986);
nand U24650 (N_24650,N_21032,N_20008);
nand U24651 (N_24651,N_20904,N_23017);
nor U24652 (N_24652,N_18365,N_21226);
nand U24653 (N_24653,N_21903,N_19544);
nand U24654 (N_24654,N_20324,N_19577);
or U24655 (N_24655,N_19069,N_20528);
and U24656 (N_24656,N_23311,N_23450);
nand U24657 (N_24657,N_20581,N_21642);
nor U24658 (N_24658,N_21995,N_19780);
xnor U24659 (N_24659,N_20005,N_20960);
nand U24660 (N_24660,N_20637,N_22510);
nor U24661 (N_24661,N_23708,N_21951);
and U24662 (N_24662,N_23053,N_19228);
nand U24663 (N_24663,N_19737,N_21975);
or U24664 (N_24664,N_23439,N_18670);
and U24665 (N_24665,N_19346,N_19988);
xor U24666 (N_24666,N_18055,N_21563);
nor U24667 (N_24667,N_20723,N_18390);
or U24668 (N_24668,N_23843,N_18109);
xor U24669 (N_24669,N_19929,N_19618);
nor U24670 (N_24670,N_18964,N_23915);
and U24671 (N_24671,N_19687,N_22322);
and U24672 (N_24672,N_21664,N_20122);
and U24673 (N_24673,N_23393,N_18633);
xor U24674 (N_24674,N_19934,N_23956);
nand U24675 (N_24675,N_18948,N_21356);
nor U24676 (N_24676,N_20481,N_22606);
xnor U24677 (N_24677,N_22406,N_22608);
xnor U24678 (N_24678,N_22217,N_18545);
xnor U24679 (N_24679,N_18403,N_22361);
nand U24680 (N_24680,N_20315,N_22682);
nor U24681 (N_24681,N_23036,N_23517);
nor U24682 (N_24682,N_21510,N_21056);
nand U24683 (N_24683,N_22683,N_22901);
xor U24684 (N_24684,N_21587,N_21330);
nor U24685 (N_24685,N_22158,N_23333);
and U24686 (N_24686,N_21952,N_20547);
nor U24687 (N_24687,N_23940,N_23767);
or U24688 (N_24688,N_20512,N_22899);
and U24689 (N_24689,N_20362,N_22684);
nor U24690 (N_24690,N_21403,N_20438);
nor U24691 (N_24691,N_19614,N_22330);
xor U24692 (N_24692,N_22999,N_23072);
nand U24693 (N_24693,N_22836,N_22995);
nor U24694 (N_24694,N_22128,N_23802);
or U24695 (N_24695,N_19320,N_21696);
and U24696 (N_24696,N_21129,N_20052);
nand U24697 (N_24697,N_19891,N_20839);
and U24698 (N_24698,N_20652,N_23551);
or U24699 (N_24699,N_18784,N_23212);
xor U24700 (N_24700,N_18671,N_23226);
and U24701 (N_24701,N_22994,N_20781);
and U24702 (N_24702,N_21874,N_18433);
or U24703 (N_24703,N_22795,N_23780);
or U24704 (N_24704,N_19241,N_18392);
nor U24705 (N_24705,N_22312,N_22532);
nand U24706 (N_24706,N_20038,N_21154);
and U24707 (N_24707,N_22202,N_22613);
nor U24708 (N_24708,N_19410,N_18059);
xnor U24709 (N_24709,N_20591,N_21155);
xor U24710 (N_24710,N_20563,N_20961);
nor U24711 (N_24711,N_23724,N_23334);
nor U24712 (N_24712,N_23519,N_18407);
xor U24713 (N_24713,N_19770,N_22060);
or U24714 (N_24714,N_22768,N_21921);
nand U24715 (N_24715,N_21997,N_23521);
nor U24716 (N_24716,N_23331,N_19692);
or U24717 (N_24717,N_18429,N_21537);
nand U24718 (N_24718,N_23787,N_20775);
nor U24719 (N_24719,N_23574,N_23579);
and U24720 (N_24720,N_21117,N_22278);
nand U24721 (N_24721,N_20774,N_23210);
nand U24722 (N_24722,N_21115,N_22874);
and U24723 (N_24723,N_21240,N_20044);
xor U24724 (N_24724,N_20157,N_19407);
nor U24725 (N_24725,N_20673,N_22909);
or U24726 (N_24726,N_19899,N_18072);
nor U24727 (N_24727,N_22454,N_22996);
or U24728 (N_24728,N_23633,N_19734);
nand U24729 (N_24729,N_19901,N_21819);
nand U24730 (N_24730,N_19631,N_20943);
xor U24731 (N_24731,N_19299,N_18728);
nand U24732 (N_24732,N_23638,N_22165);
xor U24733 (N_24733,N_23911,N_23866);
and U24734 (N_24734,N_18583,N_23598);
or U24735 (N_24735,N_18334,N_18760);
and U24736 (N_24736,N_18217,N_19645);
and U24737 (N_24737,N_19460,N_21844);
or U24738 (N_24738,N_23650,N_23818);
or U24739 (N_24739,N_22456,N_23114);
nand U24740 (N_24740,N_23953,N_18835);
xnor U24741 (N_24741,N_23401,N_23123);
nor U24742 (N_24742,N_21270,N_18457);
nor U24743 (N_24743,N_22493,N_19829);
xnor U24744 (N_24744,N_20209,N_19534);
and U24745 (N_24745,N_22286,N_23622);
or U24746 (N_24746,N_20097,N_19760);
nand U24747 (N_24747,N_19182,N_18552);
nor U24748 (N_24748,N_22737,N_19846);
nand U24749 (N_24749,N_20327,N_18384);
and U24750 (N_24750,N_19101,N_21063);
or U24751 (N_24751,N_19783,N_23628);
or U24752 (N_24752,N_21172,N_18647);
or U24753 (N_24753,N_22319,N_19628);
and U24754 (N_24754,N_18612,N_21560);
nand U24755 (N_24755,N_23223,N_22405);
and U24756 (N_24756,N_22254,N_22558);
nand U24757 (N_24757,N_20761,N_20576);
and U24758 (N_24758,N_20313,N_18284);
or U24759 (N_24759,N_22637,N_21638);
nand U24760 (N_24760,N_18329,N_19127);
nor U24761 (N_24761,N_19579,N_19292);
nor U24762 (N_24762,N_18309,N_23336);
nand U24763 (N_24763,N_23409,N_23368);
nor U24764 (N_24764,N_18580,N_23163);
xor U24765 (N_24765,N_23803,N_19080);
or U24766 (N_24766,N_18810,N_21395);
nor U24767 (N_24767,N_18401,N_20989);
xnor U24768 (N_24768,N_20430,N_19924);
xnor U24769 (N_24769,N_21660,N_23173);
xor U24770 (N_24770,N_21829,N_19015);
nor U24771 (N_24771,N_18879,N_19805);
nand U24772 (N_24772,N_20718,N_21670);
and U24773 (N_24773,N_19959,N_19113);
nor U24774 (N_24774,N_22543,N_19345);
nand U24775 (N_24775,N_21370,N_20221);
and U24776 (N_24776,N_22211,N_19870);
nor U24777 (N_24777,N_22023,N_23536);
or U24778 (N_24778,N_21326,N_22951);
or U24779 (N_24779,N_19892,N_19056);
or U24780 (N_24780,N_19669,N_18872);
nand U24781 (N_24781,N_22303,N_23976);
and U24782 (N_24782,N_19775,N_21033);
and U24783 (N_24783,N_23967,N_20850);
xnor U24784 (N_24784,N_23305,N_21082);
nor U24785 (N_24785,N_21531,N_20242);
xor U24786 (N_24786,N_21159,N_21503);
and U24787 (N_24787,N_23903,N_19443);
and U24788 (N_24788,N_21336,N_18198);
and U24789 (N_24789,N_20333,N_18893);
nor U24790 (N_24790,N_20145,N_22265);
nand U24791 (N_24791,N_20993,N_21059);
nor U24792 (N_24792,N_21090,N_19239);
or U24793 (N_24793,N_23867,N_20882);
or U24794 (N_24794,N_18244,N_20073);
and U24795 (N_24795,N_19006,N_20887);
and U24796 (N_24796,N_21937,N_20680);
nand U24797 (N_24797,N_18188,N_19381);
and U24798 (N_24798,N_21254,N_22595);
and U24799 (N_24799,N_20903,N_18023);
nor U24800 (N_24800,N_23449,N_21776);
and U24801 (N_24801,N_22274,N_19150);
and U24802 (N_24802,N_22970,N_19405);
nand U24803 (N_24803,N_18761,N_23056);
and U24804 (N_24804,N_20090,N_18658);
nand U24805 (N_24805,N_18557,N_19366);
xor U24806 (N_24806,N_21157,N_18579);
and U24807 (N_24807,N_18087,N_18000);
nand U24808 (N_24808,N_22486,N_23277);
xnor U24809 (N_24809,N_20954,N_20511);
or U24810 (N_24810,N_23345,N_18074);
xor U24811 (N_24811,N_18141,N_20061);
or U24812 (N_24812,N_23532,N_18082);
and U24813 (N_24813,N_22602,N_20427);
nor U24814 (N_24814,N_22307,N_22448);
nand U24815 (N_24815,N_20670,N_18326);
nor U24816 (N_24816,N_23826,N_23274);
nand U24817 (N_24817,N_21625,N_23932);
or U24818 (N_24818,N_20942,N_22757);
nand U24819 (N_24819,N_21572,N_21516);
or U24820 (N_24820,N_20164,N_19376);
and U24821 (N_24821,N_18496,N_20490);
nor U24822 (N_24822,N_20654,N_20480);
nor U24823 (N_24823,N_22755,N_22723);
and U24824 (N_24824,N_21255,N_18219);
nand U24825 (N_24825,N_18834,N_23068);
nand U24826 (N_24826,N_19888,N_22572);
nor U24827 (N_24827,N_19112,N_18282);
and U24828 (N_24828,N_19691,N_18162);
nand U24829 (N_24829,N_20836,N_19884);
or U24830 (N_24830,N_23616,N_21262);
nand U24831 (N_24831,N_18154,N_18980);
nor U24832 (N_24832,N_22009,N_20215);
nor U24833 (N_24833,N_21609,N_20253);
or U24834 (N_24834,N_23592,N_23601);
and U24835 (N_24835,N_20486,N_21246);
or U24836 (N_24836,N_23854,N_23692);
xor U24837 (N_24837,N_21257,N_22975);
and U24838 (N_24838,N_18925,N_20541);
xnor U24839 (N_24839,N_23255,N_21207);
nand U24840 (N_24840,N_22915,N_18312);
xnor U24841 (N_24841,N_23458,N_20806);
and U24842 (N_24842,N_21549,N_22509);
or U24843 (N_24843,N_21559,N_21777);
and U24844 (N_24844,N_20187,N_19334);
nor U24845 (N_24845,N_18910,N_22442);
or U24846 (N_24846,N_23021,N_21515);
and U24847 (N_24847,N_20488,N_22041);
and U24848 (N_24848,N_21799,N_19199);
or U24849 (N_24849,N_22977,N_20949);
nor U24850 (N_24850,N_20103,N_22082);
nand U24851 (N_24851,N_21911,N_23400);
nand U24852 (N_24852,N_19347,N_23505);
and U24853 (N_24853,N_19894,N_21520);
xor U24854 (N_24854,N_22937,N_23665);
and U24855 (N_24855,N_22712,N_22502);
or U24856 (N_24856,N_20063,N_20304);
and U24857 (N_24857,N_20031,N_19341);
xor U24858 (N_24858,N_21908,N_18740);
and U24859 (N_24859,N_19430,N_20838);
nand U24860 (N_24860,N_22815,N_22068);
xnor U24861 (N_24861,N_21123,N_21276);
nand U24862 (N_24862,N_18957,N_23383);
xnor U24863 (N_24863,N_21291,N_18027);
nand U24864 (N_24864,N_23699,N_20147);
nand U24865 (N_24865,N_20069,N_20808);
and U24866 (N_24866,N_19398,N_18199);
and U24867 (N_24867,N_19791,N_19305);
nand U24868 (N_24868,N_23299,N_22087);
and U24869 (N_24869,N_23216,N_19311);
nor U24870 (N_24870,N_18281,N_23448);
nand U24871 (N_24871,N_18985,N_20281);
nand U24872 (N_24872,N_21533,N_20888);
and U24873 (N_24873,N_20397,N_23506);
and U24874 (N_24874,N_22866,N_22306);
nand U24875 (N_24875,N_21005,N_21413);
and U24876 (N_24876,N_22038,N_19718);
xor U24877 (N_24877,N_21040,N_21221);
or U24878 (N_24878,N_20738,N_18008);
or U24879 (N_24879,N_20000,N_18954);
nor U24880 (N_24880,N_22958,N_19863);
nand U24881 (N_24881,N_23885,N_19269);
and U24882 (N_24882,N_19867,N_19488);
nand U24883 (N_24883,N_18789,N_20597);
and U24884 (N_24884,N_18614,N_21542);
xnor U24885 (N_24885,N_18534,N_19457);
xor U24886 (N_24886,N_20233,N_21265);
nand U24887 (N_24887,N_23846,N_20894);
or U24888 (N_24888,N_23008,N_19886);
nand U24889 (N_24889,N_18168,N_18060);
and U24890 (N_24890,N_19029,N_22511);
and U24891 (N_24891,N_23253,N_20153);
nor U24892 (N_24892,N_22072,N_18140);
nand U24893 (N_24893,N_21287,N_18235);
xor U24894 (N_24894,N_19111,N_19329);
or U24895 (N_24895,N_19979,N_23030);
or U24896 (N_24896,N_20896,N_19665);
and U24897 (N_24897,N_23515,N_23185);
and U24898 (N_24898,N_22745,N_22594);
nand U24899 (N_24899,N_21044,N_19657);
nand U24900 (N_24900,N_21188,N_20249);
nand U24901 (N_24901,N_23726,N_19088);
or U24902 (N_24902,N_20618,N_23485);
nor U24903 (N_24903,N_19483,N_20556);
nor U24904 (N_24904,N_19598,N_23162);
nand U24905 (N_24905,N_23394,N_23032);
xor U24906 (N_24906,N_21234,N_22762);
or U24907 (N_24907,N_21667,N_23348);
xnor U24908 (N_24908,N_21426,N_21086);
nand U24909 (N_24909,N_18840,N_22856);
nor U24910 (N_24910,N_19852,N_21655);
nor U24911 (N_24911,N_20812,N_20478);
xor U24912 (N_24912,N_18820,N_22195);
and U24913 (N_24913,N_19940,N_22139);
or U24914 (N_24914,N_19732,N_19026);
xnor U24915 (N_24915,N_20054,N_19851);
xnor U24916 (N_24916,N_20185,N_22863);
nor U24917 (N_24917,N_23325,N_20414);
xnor U24918 (N_24918,N_22917,N_21105);
nand U24919 (N_24919,N_20307,N_21205);
and U24920 (N_24920,N_22296,N_23949);
or U24921 (N_24921,N_19547,N_19619);
and U24922 (N_24922,N_20610,N_18800);
xnor U24923 (N_24923,N_18406,N_20220);
nor U24924 (N_24924,N_23222,N_19915);
or U24925 (N_24925,N_23586,N_21839);
and U24926 (N_24926,N_18622,N_19803);
nand U24927 (N_24927,N_21624,N_21928);
nand U24928 (N_24928,N_19391,N_23016);
nor U24929 (N_24929,N_19830,N_18316);
nor U24930 (N_24930,N_21589,N_22184);
and U24931 (N_24931,N_18729,N_19315);
nand U24932 (N_24932,N_20375,N_19493);
xnor U24933 (N_24933,N_21378,N_20713);
nor U24934 (N_24934,N_20837,N_21721);
xnor U24935 (N_24935,N_20273,N_22396);
xor U24936 (N_24936,N_22131,N_21339);
xor U24937 (N_24937,N_19340,N_19470);
or U24938 (N_24938,N_22460,N_18377);
nor U24939 (N_24939,N_22005,N_23813);
xnor U24940 (N_24940,N_19792,N_20460);
or U24941 (N_24941,N_22630,N_21325);
xnor U24942 (N_24942,N_18989,N_21800);
xor U24943 (N_24943,N_20767,N_18307);
and U24944 (N_24944,N_19012,N_18825);
xnor U24945 (N_24945,N_21830,N_19896);
nor U24946 (N_24946,N_21851,N_18412);
nand U24947 (N_24947,N_22114,N_23037);
or U24948 (N_24948,N_23510,N_23615);
nand U24949 (N_24949,N_19823,N_23498);
or U24950 (N_24950,N_20640,N_18197);
or U24951 (N_24951,N_20649,N_18944);
xnor U24952 (N_24952,N_21641,N_22784);
xor U24953 (N_24953,N_23459,N_21309);
and U24954 (N_24954,N_19125,N_22133);
nand U24955 (N_24955,N_20791,N_22479);
xor U24956 (N_24956,N_22055,N_22280);
or U24957 (N_24957,N_19923,N_20503);
xnor U24958 (N_24958,N_18817,N_22054);
nor U24959 (N_24959,N_21896,N_23010);
nand U24960 (N_24960,N_22411,N_23091);
nand U24961 (N_24961,N_23676,N_20557);
or U24962 (N_24962,N_22948,N_21428);
nand U24963 (N_24963,N_21077,N_18895);
xnor U24964 (N_24964,N_20514,N_19731);
xor U24965 (N_24965,N_22582,N_20918);
xor U24966 (N_24966,N_23675,N_19270);
nor U24967 (N_24967,N_20116,N_19739);
xor U24968 (N_24968,N_20783,N_19860);
nor U24969 (N_24969,N_21690,N_18002);
nor U24970 (N_24970,N_21708,N_18456);
nand U24971 (N_24971,N_20002,N_19049);
and U24972 (N_24972,N_23308,N_22552);
nor U24973 (N_24973,N_23014,N_19594);
nor U24974 (N_24974,N_20594,N_19911);
nand U24975 (N_24975,N_21001,N_18711);
and U24976 (N_24976,N_23012,N_19365);
or U24977 (N_24977,N_20957,N_22925);
or U24978 (N_24978,N_23049,N_23316);
or U24979 (N_24979,N_19749,N_19926);
nor U24980 (N_24980,N_22365,N_20962);
xor U24981 (N_24981,N_23203,N_20084);
and U24982 (N_24982,N_22969,N_23271);
and U24983 (N_24983,N_20352,N_22792);
nor U24984 (N_24984,N_22110,N_22394);
xnor U24985 (N_24985,N_23766,N_20963);
nor U24986 (N_24986,N_20111,N_22944);
nand U24987 (N_24987,N_19070,N_19181);
or U24988 (N_24988,N_21438,N_23164);
nand U24989 (N_24989,N_19713,N_18701);
nand U24990 (N_24990,N_19212,N_19868);
nand U24991 (N_24991,N_19582,N_19084);
nor U24992 (N_24992,N_20170,N_20087);
xnor U24993 (N_24993,N_20690,N_22449);
nand U24994 (N_24994,N_18777,N_19853);
xnor U24995 (N_24995,N_19667,N_18502);
and U24996 (N_24996,N_21744,N_20832);
or U24997 (N_24997,N_19377,N_23907);
nor U24998 (N_24998,N_19126,N_18180);
and U24999 (N_24999,N_21718,N_18914);
nand U25000 (N_25000,N_21450,N_22103);
and U25001 (N_25001,N_20441,N_21286);
xor U25002 (N_25002,N_22373,N_21183);
and U25003 (N_25003,N_19995,N_21632);
or U25004 (N_25004,N_18710,N_19054);
or U25005 (N_25005,N_21689,N_21160);
nor U25006 (N_25006,N_23087,N_21353);
nor U25007 (N_25007,N_19869,N_19276);
nor U25008 (N_25008,N_22618,N_18126);
and U25009 (N_25009,N_22936,N_20826);
and U25010 (N_25010,N_18751,N_21264);
nor U25011 (N_25011,N_22920,N_22705);
nand U25012 (N_25012,N_20418,N_22616);
xnor U25013 (N_25013,N_22313,N_21910);
or U25014 (N_25014,N_20260,N_20390);
and U25015 (N_25015,N_20025,N_21994);
or U25016 (N_25016,N_23712,N_18591);
or U25017 (N_25017,N_23528,N_22200);
nor U25018 (N_25018,N_22480,N_22748);
and U25019 (N_25019,N_21021,N_22867);
nor U25020 (N_25020,N_21592,N_21600);
xnor U25021 (N_25021,N_23375,N_23076);
nand U25022 (N_25022,N_22750,N_22316);
nor U25023 (N_25023,N_21653,N_19429);
or U25024 (N_25024,N_20022,N_18076);
nor U25025 (N_25025,N_23833,N_23369);
nor U25026 (N_25026,N_18073,N_20844);
and U25027 (N_25027,N_23759,N_21895);
nor U25028 (N_25028,N_22645,N_20330);
nor U25029 (N_25029,N_19344,N_18388);
nor U25030 (N_25030,N_21054,N_18054);
nand U25031 (N_25031,N_18498,N_19436);
or U25032 (N_25032,N_21588,N_20489);
or U25033 (N_25033,N_22831,N_20299);
nand U25034 (N_25034,N_18029,N_18993);
and U25035 (N_25035,N_20368,N_21722);
or U25036 (N_25036,N_23639,N_19293);
nor U25037 (N_25037,N_22366,N_19158);
nand U25038 (N_25038,N_20334,N_19524);
nor U25039 (N_25039,N_21102,N_20421);
nand U25040 (N_25040,N_22854,N_22436);
and U25041 (N_25041,N_23488,N_19536);
and U25042 (N_25042,N_23140,N_23130);
or U25043 (N_25043,N_19653,N_21818);
and U25044 (N_25044,N_21199,N_18323);
and U25045 (N_25045,N_19980,N_20224);
and U25046 (N_25046,N_19693,N_20258);
and U25047 (N_25047,N_21882,N_19373);
or U25048 (N_25048,N_23390,N_20522);
and U25049 (N_25049,N_22279,N_20168);
or U25050 (N_25050,N_21307,N_21525);
or U25051 (N_25051,N_18783,N_19372);
xnor U25052 (N_25052,N_19230,N_21416);
xnor U25053 (N_25053,N_20636,N_18946);
or U25054 (N_25054,N_20020,N_22671);
or U25055 (N_25055,N_21218,N_21241);
nor U25056 (N_25056,N_22599,N_22410);
and U25057 (N_25057,N_23246,N_21581);
nor U25058 (N_25058,N_20872,N_23667);
nand U25059 (N_25059,N_23106,N_22026);
or U25060 (N_25060,N_20678,N_20230);
and U25061 (N_25061,N_20374,N_19482);
or U25062 (N_25062,N_22914,N_23800);
xor U25063 (N_25063,N_23486,N_23193);
nor U25064 (N_25064,N_20700,N_19162);
xnor U25065 (N_25065,N_19471,N_21037);
and U25066 (N_25066,N_19756,N_19591);
or U25067 (N_25067,N_23504,N_22206);
or U25068 (N_25068,N_18497,N_21213);
and U25069 (N_25069,N_23233,N_18038);
nor U25070 (N_25070,N_22423,N_21321);
xor U25071 (N_25071,N_22633,N_18953);
xor U25072 (N_25072,N_19253,N_23740);
xnor U25073 (N_25073,N_21208,N_18697);
or U25074 (N_25074,N_22860,N_19177);
nor U25075 (N_25075,N_20750,N_22326);
or U25076 (N_25076,N_21364,N_23909);
or U25077 (N_25077,N_22539,N_19933);
or U25078 (N_25078,N_23104,N_19041);
nor U25079 (N_25079,N_20264,N_22031);
nor U25080 (N_25080,N_23384,N_19490);
and U25081 (N_25081,N_19441,N_21078);
or U25082 (N_25082,N_22585,N_20484);
or U25083 (N_25083,N_22676,N_22997);
or U25084 (N_25084,N_22052,N_23025);
nor U25085 (N_25085,N_19668,N_18769);
nor U25086 (N_25086,N_18935,N_23379);
nor U25087 (N_25087,N_20593,N_20847);
nand U25088 (N_25088,N_23159,N_21699);
nor U25089 (N_25089,N_23850,N_21550);
nand U25090 (N_25090,N_22868,N_19632);
xor U25091 (N_25091,N_22929,N_20027);
and U25092 (N_25092,N_22291,N_23270);
nor U25093 (N_25093,N_19592,N_21193);
nand U25094 (N_25094,N_21275,N_19303);
nor U25095 (N_25095,N_19338,N_18846);
or U25096 (N_25096,N_18882,N_23178);
nor U25097 (N_25097,N_20259,N_23670);
nor U25098 (N_25098,N_23655,N_21788);
and U25099 (N_25099,N_18924,N_23141);
xnor U25100 (N_25100,N_20905,N_22674);
or U25101 (N_25101,N_18058,N_20261);
xnor U25102 (N_25102,N_19302,N_23627);
nor U25103 (N_25103,N_21665,N_22484);
nand U25104 (N_25104,N_21057,N_21277);
xor U25105 (N_25105,N_22893,N_21629);
and U25106 (N_25106,N_19567,N_22100);
xnor U25107 (N_25107,N_19479,N_18181);
or U25108 (N_25108,N_22570,N_19396);
nor U25109 (N_25109,N_22962,N_23578);
nand U25110 (N_25110,N_19110,N_21534);
and U25111 (N_25111,N_19065,N_18527);
or U25112 (N_25112,N_18264,N_20705);
or U25113 (N_25113,N_20492,N_21909);
or U25114 (N_25114,N_21530,N_22115);
nor U25115 (N_25115,N_20026,N_23778);
and U25116 (N_25116,N_22001,N_23427);
and U25117 (N_25117,N_19809,N_19512);
nor U25118 (N_25118,N_19323,N_18036);
or U25119 (N_25119,N_23771,N_21774);
xnor U25120 (N_25120,N_19035,N_18351);
xnor U25121 (N_25121,N_23876,N_22652);
xor U25122 (N_25122,N_21784,N_21162);
and U25123 (N_25123,N_23183,N_20585);
or U25124 (N_25124,N_18451,N_18031);
and U25125 (N_25125,N_21623,N_23309);
xor U25126 (N_25126,N_19971,N_19326);
xor U25127 (N_25127,N_23174,N_21083);
nor U25128 (N_25128,N_23587,N_18050);
nor U25129 (N_25129,N_21206,N_22369);
nand U25130 (N_25130,N_23593,N_20213);
or U25131 (N_25131,N_20584,N_20569);
nand U25132 (N_25132,N_21087,N_19023);
nand U25133 (N_25133,N_19009,N_21458);
xor U25134 (N_25134,N_18248,N_23980);
or U25135 (N_25135,N_18548,N_18928);
or U25136 (N_25136,N_18186,N_18007);
nand U25137 (N_25137,N_22006,N_19105);
and U25138 (N_25138,N_18448,N_22698);
xnor U25139 (N_25139,N_19956,N_22522);
and U25140 (N_25140,N_19698,N_23137);
nor U25141 (N_25141,N_20714,N_22953);
nand U25142 (N_25142,N_18034,N_23011);
xor U25143 (N_25143,N_21834,N_23944);
nor U25144 (N_25144,N_23191,N_19542);
nor U25145 (N_25145,N_23784,N_18803);
nor U25146 (N_25146,N_18437,N_20265);
xor U25147 (N_25147,N_18926,N_23120);
or U25148 (N_25148,N_22923,N_22081);
nand U25149 (N_25149,N_18278,N_18131);
nand U25150 (N_25150,N_21712,N_22111);
nor U25151 (N_25151,N_23181,N_22255);
nand U25152 (N_25152,N_19602,N_18958);
and U25153 (N_25153,N_22453,N_23895);
xor U25154 (N_25154,N_20815,N_18420);
nand U25155 (N_25155,N_21596,N_19617);
and U25156 (N_25156,N_22981,N_20929);
and U25157 (N_25157,N_23822,N_22812);
nand U25158 (N_25158,N_22113,N_19938);
nand U25159 (N_25159,N_19333,N_22135);
nand U25160 (N_25160,N_21186,N_22934);
xor U25161 (N_25161,N_19104,N_23658);
or U25162 (N_25162,N_22021,N_22127);
or U25163 (N_25163,N_21385,N_23704);
and U25164 (N_25164,N_19897,N_20217);
nand U25165 (N_25165,N_20204,N_18161);
nor U25166 (N_25166,N_20423,N_20395);
nand U25167 (N_25167,N_19103,N_21290);
and U25168 (N_25168,N_19356,N_20715);
nor U25169 (N_25169,N_19706,N_21003);
nand U25170 (N_25170,N_21041,N_20191);
or U25171 (N_25171,N_23649,N_20245);
nor U25172 (N_25172,N_20341,N_19670);
and U25173 (N_25173,N_20189,N_21219);
nor U25174 (N_25174,N_21266,N_23256);
or U25175 (N_25175,N_19222,N_19018);
or U25176 (N_25176,N_18562,N_19079);
nor U25177 (N_25177,N_23651,N_21759);
nor U25178 (N_25178,N_22029,N_18997);
nor U25179 (N_25179,N_19513,N_22910);
xor U25180 (N_25180,N_18397,N_23263);
nor U25181 (N_25181,N_21380,N_20192);
or U25182 (N_25182,N_23987,N_20456);
and U25183 (N_25183,N_21394,N_21869);
or U25184 (N_25184,N_22343,N_20566);
or U25185 (N_25185,N_18107,N_19057);
and U25186 (N_25186,N_22897,N_19676);
nand U25187 (N_25187,N_18736,N_20629);
xor U25188 (N_25188,N_22734,N_23107);
xor U25189 (N_25189,N_21700,N_23853);
nor U25190 (N_25190,N_21577,N_21993);
nor U25191 (N_25191,N_21456,N_20780);
nor U25192 (N_25192,N_22138,N_19500);
or U25193 (N_25193,N_18236,N_23777);
or U25194 (N_25194,N_23195,N_21434);
and U25195 (N_25195,N_22198,N_18904);
nand U25196 (N_25196,N_23050,N_18509);
and U25197 (N_25197,N_21256,N_21734);
nand U25198 (N_25198,N_20074,N_19967);
nor U25199 (N_25199,N_19121,N_18675);
and U25200 (N_25200,N_22156,N_23604);
nor U25201 (N_25201,N_23063,N_19359);
and U25202 (N_25202,N_22282,N_18354);
or U25203 (N_25203,N_23590,N_23839);
xnor U25204 (N_25204,N_18646,N_21594);
xor U25205 (N_25205,N_19186,N_23064);
nand U25206 (N_25206,N_20958,N_19661);
or U25207 (N_25207,N_18201,N_19942);
xor U25208 (N_25208,N_19527,N_19096);
or U25209 (N_25209,N_23701,N_20039);
or U25210 (N_25210,N_18564,N_22422);
and U25211 (N_25211,N_22196,N_20231);
or U25212 (N_25212,N_21961,N_19420);
or U25213 (N_25213,N_22010,N_23198);
or U25214 (N_25214,N_22655,N_18555);
xor U25215 (N_25215,N_23234,N_22754);
and U25216 (N_25216,N_20638,N_19541);
nor U25217 (N_25217,N_19178,N_22822);
or U25218 (N_25218,N_22524,N_18631);
nor U25219 (N_25219,N_23553,N_23729);
xnor U25220 (N_25220,N_18157,N_23570);
nor U25221 (N_25221,N_20955,N_18292);
or U25222 (N_25222,N_23660,N_21757);
or U25223 (N_25223,N_23428,N_21954);
nand U25224 (N_25224,N_21887,N_23904);
xor U25225 (N_25225,N_19745,N_19031);
nor U25226 (N_25226,N_18805,N_19097);
xnor U25227 (N_25227,N_20679,N_19735);
and U25228 (N_25228,N_20605,N_19273);
nor U25229 (N_25229,N_23115,N_21002);
nor U25230 (N_25230,N_18987,N_20650);
and U25231 (N_25231,N_20590,N_23436);
or U25232 (N_25232,N_22984,N_19141);
xor U25233 (N_25233,N_20822,N_21362);
nor U25234 (N_25234,N_23111,N_19371);
nand U25235 (N_25235,N_21111,N_23003);
and U25236 (N_25236,N_22224,N_22714);
and U25237 (N_25237,N_22814,N_21604);
nand U25238 (N_25238,N_22739,N_23597);
or U25239 (N_25239,N_23093,N_21765);
nor U25240 (N_25240,N_20321,N_19480);
nor U25241 (N_25241,N_19207,N_21745);
and U25242 (N_25242,N_19890,N_22793);
and U25243 (N_25243,N_19742,N_22384);
nor U25244 (N_25244,N_21915,N_18860);
nor U25245 (N_25245,N_23019,N_21064);
and U25246 (N_25246,N_23062,N_18409);
xnor U25247 (N_25247,N_20769,N_18077);
nor U25248 (N_25248,N_20959,N_22363);
and U25249 (N_25249,N_19714,N_21732);
nor U25250 (N_25250,N_22578,N_19086);
nand U25251 (N_25251,N_21501,N_21073);
nor U25252 (N_25252,N_18666,N_22169);
nor U25253 (N_25253,N_20825,N_20759);
or U25254 (N_25254,N_18184,N_21402);
or U25255 (N_25255,N_21652,N_23287);
and U25256 (N_25256,N_19130,N_18742);
and U25257 (N_25257,N_20600,N_19725);
nor U25258 (N_25258,N_18163,N_18395);
nor U25259 (N_25259,N_23493,N_23531);
nand U25260 (N_25260,N_18942,N_22843);
and U25261 (N_25261,N_18303,N_21347);
or U25262 (N_25262,N_22871,N_20257);
nand U25263 (N_25263,N_18679,N_18818);
xnor U25264 (N_25264,N_21512,N_22310);
nand U25265 (N_25265,N_22426,N_18503);
nand U25266 (N_25266,N_18518,N_18669);
nor U25267 (N_25267,N_19165,N_22635);
or U25268 (N_25268,N_21094,N_18726);
nor U25269 (N_25269,N_21489,N_21099);
nand U25270 (N_25270,N_21446,N_23259);
nor U25271 (N_25271,N_23060,N_21918);
xor U25272 (N_25272,N_18727,N_23291);
nor U25273 (N_25273,N_18359,N_22538);
xor U25274 (N_25274,N_18063,N_20996);
or U25275 (N_25275,N_19468,N_22276);
and U25276 (N_25276,N_19849,N_22961);
or U25277 (N_25277,N_22036,N_22826);
or U25278 (N_25278,N_19951,N_21785);
and U25279 (N_25279,N_22336,N_20089);
nand U25280 (N_25280,N_21342,N_21787);
nand U25281 (N_25281,N_21253,N_22403);
and U25282 (N_25282,N_21143,N_20841);
or U25283 (N_25283,N_18234,N_22731);
or U25284 (N_25284,N_21293,N_23238);
nor U25285 (N_25285,N_18015,N_20865);
nor U25286 (N_25286,N_22253,N_22841);
xor U25287 (N_25287,N_22786,N_23861);
xor U25288 (N_25288,N_22880,N_19003);
or U25289 (N_25289,N_20118,N_22235);
nand U25290 (N_25290,N_22568,N_22829);
and U25291 (N_25291,N_21981,N_22458);
nand U25292 (N_25292,N_23042,N_20348);
nand U25293 (N_25293,N_20657,N_23857);
nor U25294 (N_25294,N_23931,N_20789);
nand U25295 (N_25295,N_22638,N_23103);
and U25296 (N_25296,N_20163,N_23760);
nor U25297 (N_25297,N_20190,N_20197);
nand U25298 (N_25298,N_21108,N_21755);
or U25299 (N_25299,N_23554,N_23407);
or U25300 (N_25300,N_19404,N_21482);
xor U25301 (N_25301,N_21610,N_18438);
xor U25302 (N_25302,N_22284,N_23922);
nor U25303 (N_25303,N_19282,N_20937);
and U25304 (N_25304,N_22588,N_23710);
or U25305 (N_25305,N_21498,N_23698);
xor U25306 (N_25306,N_23026,N_23138);
nand U25307 (N_25307,N_19787,N_19484);
nor U25308 (N_25308,N_18604,N_19744);
and U25309 (N_25309,N_21408,N_21317);
nor U25310 (N_25310,N_21860,N_23769);
xor U25311 (N_25311,N_19266,N_18132);
xor U25312 (N_25312,N_22688,N_18381);
or U25313 (N_25313,N_18837,N_22989);
nor U25314 (N_25314,N_22744,N_21080);
nand U25315 (N_25315,N_18129,N_20509);
and U25316 (N_25316,N_20796,N_19765);
nor U25317 (N_25317,N_23605,N_20110);
xnor U25318 (N_25318,N_19082,N_23626);
or U25319 (N_25319,N_19350,N_21867);
xnor U25320 (N_25320,N_20183,N_18645);
and U25321 (N_25321,N_21425,N_20617);
xnor U25322 (N_25322,N_18823,N_21815);
nor U25323 (N_25323,N_22565,N_20574);
xnor U25324 (N_25324,N_22457,N_20353);
and U25325 (N_25325,N_19650,N_20126);
and U25326 (N_25326,N_20417,N_18192);
xor U25327 (N_25327,N_23039,N_23069);
nor U25328 (N_25328,N_22151,N_21429);
nor U25329 (N_25329,N_21976,N_22895);
xnor U25330 (N_25330,N_20645,N_20194);
nand U25331 (N_25331,N_19452,N_21238);
xor U25332 (N_25332,N_21131,N_18947);
xnor U25333 (N_25333,N_22120,N_18125);
xor U25334 (N_25334,N_20754,N_20055);
or U25335 (N_25335,N_22495,N_21178);
or U25336 (N_25336,N_19300,N_23954);
nor U25337 (N_25337,N_18218,N_22432);
or U25338 (N_25338,N_19571,N_18841);
xor U25339 (N_25339,N_23057,N_21404);
and U25340 (N_25340,N_19331,N_21473);
nand U25341 (N_25341,N_20660,N_20053);
nor U25342 (N_25342,N_19585,N_23283);
nand U25343 (N_25343,N_20855,N_21068);
or U25344 (N_25344,N_22513,N_23852);
nand U25345 (N_25345,N_23981,N_21135);
nand U25346 (N_25346,N_21735,N_19839);
or U25347 (N_25347,N_22190,N_20909);
nand U25348 (N_25348,N_21081,N_18070);
xnor U25349 (N_25349,N_19828,N_23542);
nor U25350 (N_25350,N_20366,N_19240);
and U25351 (N_25351,N_21528,N_23020);
nor U25352 (N_25352,N_21454,N_23303);
or U25353 (N_25353,N_18220,N_21934);
nand U25354 (N_25354,N_21565,N_21169);
xnor U25355 (N_25355,N_18142,N_23735);
nor U25356 (N_25356,N_19007,N_22033);
nand U25357 (N_25357,N_19662,N_21840);
xor U25358 (N_25358,N_19379,N_21640);
nor U25359 (N_25359,N_23961,N_23952);
and U25360 (N_25360,N_20021,N_18143);
or U25361 (N_25361,N_22850,N_21076);
and U25362 (N_25362,N_23478,N_21852);
or U25363 (N_25363,N_18753,N_22879);
or U25364 (N_25364,N_23929,N_22098);
nand U25365 (N_25365,N_20803,N_20155);
or U25366 (N_25366,N_18200,N_20802);
or U25367 (N_25367,N_21703,N_23973);
or U25368 (N_25368,N_23559,N_18637);
and U25369 (N_25369,N_22439,N_20381);
and U25370 (N_25370,N_20331,N_20106);
nand U25371 (N_25371,N_18816,N_23357);
nand U25372 (N_25372,N_23883,N_18693);
or U25373 (N_25373,N_23742,N_19274);
nand U25374 (N_25374,N_18170,N_23023);
nor U25375 (N_25375,N_22266,N_21060);
and U25376 (N_25376,N_20407,N_19546);
nand U25377 (N_25377,N_19532,N_20207);
and U25378 (N_25378,N_18706,N_18807);
nand U25379 (N_25379,N_19900,N_23061);
and U25380 (N_25380,N_21750,N_20529);
and U25381 (N_25381,N_18237,N_20358);
or U25382 (N_25382,N_18275,N_21478);
nand U25383 (N_25383,N_23196,N_19053);
or U25384 (N_25384,N_18570,N_22071);
and U25385 (N_25385,N_23097,N_22080);
nand U25386 (N_25386,N_18797,N_23836);
nand U25387 (N_25387,N_23089,N_20577);
nor U25388 (N_25388,N_20615,N_23496);
xnor U25389 (N_25389,N_18037,N_21042);
and U25390 (N_25390,N_21036,N_23005);
or U25391 (N_25391,N_20867,N_20624);
nor U25392 (N_25392,N_21189,N_21101);
nand U25393 (N_25393,N_20067,N_23643);
or U25394 (N_25394,N_23433,N_19367);
nor U25395 (N_25395,N_18648,N_19419);
xor U25396 (N_25396,N_19958,N_18969);
and U25397 (N_25397,N_19776,N_18624);
nor U25398 (N_25398,N_18454,N_19093);
and U25399 (N_25399,N_20227,N_23522);
and U25400 (N_25400,N_23313,N_20843);
nand U25401 (N_25401,N_21437,N_21463);
or U25402 (N_25402,N_20272,N_20773);
xor U25403 (N_25403,N_18061,N_19495);
nor U25404 (N_25404,N_23135,N_19038);
and U25405 (N_25405,N_18048,N_20524);
nor U25406 (N_25406,N_19312,N_18550);
nor U25407 (N_25407,N_18766,N_23441);
or U25408 (N_25408,N_23386,N_22781);
xnor U25409 (N_25409,N_18152,N_23200);
nor U25410 (N_25410,N_20208,N_22285);
nor U25411 (N_25411,N_21004,N_21158);
xor U25412 (N_25412,N_22527,N_22299);
nor U25413 (N_25413,N_22516,N_19862);
xor U25414 (N_25414,N_21299,N_23362);
nand U25415 (N_25415,N_21107,N_21308);
or U25416 (N_25416,N_18101,N_22476);
nand U25417 (N_25417,N_18026,N_20987);
and U25418 (N_25418,N_21010,N_22123);
or U25419 (N_25419,N_21939,N_19152);
xor U25420 (N_25420,N_19921,N_22032);
xnor U25421 (N_25421,N_19386,N_21071);
or U25422 (N_25422,N_20276,N_23018);
nor U25423 (N_25423,N_18453,N_18480);
or U25424 (N_25424,N_18685,N_18719);
nand U25425 (N_25425,N_20337,N_23985);
and U25426 (N_25426,N_21751,N_21302);
nor U25427 (N_25427,N_18206,N_23899);
xor U25428 (N_25428,N_20287,N_18897);
or U25429 (N_25429,N_20885,N_22663);
nand U25430 (N_25430,N_21051,N_20602);
and U25431 (N_25431,N_21381,N_19509);
or U25432 (N_25432,N_18652,N_21554);
nand U25433 (N_25433,N_20971,N_21711);
xnor U25434 (N_25434,N_19388,N_19673);
nor U25435 (N_25435,N_22435,N_21964);
nor U25436 (N_25436,N_23220,N_19808);
nand U25437 (N_25437,N_20325,N_21584);
nand U25438 (N_25438,N_23442,N_22101);
nor U25439 (N_25439,N_20739,N_21447);
and U25440 (N_25440,N_22555,N_23936);
and U25441 (N_25441,N_23465,N_19160);
xnor U25442 (N_25442,N_21627,N_19952);
or U25443 (N_25443,N_22857,N_20130);
and U25444 (N_25444,N_18476,N_19232);
nor U25445 (N_25445,N_22434,N_18569);
or U25446 (N_25446,N_22228,N_23613);
or U25447 (N_25447,N_21267,N_21719);
nand U25448 (N_25448,N_20518,N_20879);
nor U25449 (N_25449,N_23972,N_22640);
or U25450 (N_25450,N_23480,N_23768);
or U25451 (N_25451,N_19248,N_20510);
or U25452 (N_25452,N_20864,N_23161);
nor U25453 (N_25453,N_21297,N_23438);
nand U25454 (N_25454,N_18490,N_20471);
nor U25455 (N_25455,N_18629,N_21771);
or U25456 (N_25456,N_21519,N_23398);
nand U25457 (N_25457,N_22482,N_18572);
nor U25458 (N_25458,N_18782,N_18998);
xnor U25459 (N_25459,N_23491,N_19795);
or U25460 (N_25460,N_21181,N_19920);
or U25461 (N_25461,N_21611,N_18231);
nor U25462 (N_25462,N_18547,N_19451);
nor U25463 (N_25463,N_18771,N_23634);
or U25464 (N_25464,N_18767,N_19148);
nand U25465 (N_25465,N_21331,N_22807);
nor U25466 (N_25466,N_23145,N_20323);
or U25467 (N_25467,N_22335,N_19877);
and U25468 (N_25468,N_21868,N_22244);
or U25469 (N_25469,N_18187,N_23361);
nand U25470 (N_25470,N_23884,N_19129);
nand U25471 (N_25471,N_23730,N_18402);
or U25472 (N_25472,N_19646,N_18641);
or U25473 (N_25473,N_18470,N_18121);
nand U25474 (N_25474,N_22916,N_20314);
nor U25475 (N_25475,N_22474,N_22263);
nor U25476 (N_25476,N_22998,N_19288);
or U25477 (N_25477,N_18778,N_22992);
xor U25478 (N_25478,N_23563,N_23462);
or U25479 (N_25479,N_21499,N_20521);
xor U25480 (N_25480,N_21917,N_22385);
nand U25481 (N_25481,N_23166,N_18687);
nand U25482 (N_25482,N_23231,N_23795);
nand U25483 (N_25483,N_23719,N_21770);
xnor U25484 (N_25484,N_23968,N_23765);
nor U25485 (N_25485,N_23978,N_23804);
and U25486 (N_25486,N_19190,N_22301);
nor U25487 (N_25487,N_21948,N_21220);
xnor U25488 (N_25488,N_22586,N_18554);
nor U25489 (N_25489,N_19142,N_22450);
xnor U25490 (N_25490,N_18428,N_19686);
nand U25491 (N_25491,N_21639,N_23824);
nand U25492 (N_25492,N_21576,N_22035);
nand U25493 (N_25493,N_20254,N_18539);
nand U25494 (N_25494,N_20162,N_23467);
and U25495 (N_25495,N_19876,N_19383);
xnor U25496 (N_25496,N_19375,N_18601);
and U25497 (N_25497,N_22964,N_21643);
and U25498 (N_25498,N_20344,N_21858);
or U25499 (N_25499,N_21982,N_22294);
nand U25500 (N_25500,N_23289,N_21876);
nor U25501 (N_25501,N_20953,N_20829);
or U25502 (N_25502,N_23739,N_20040);
and U25503 (N_25503,N_19385,N_22425);
nor U25504 (N_25504,N_22227,N_22048);
and U25505 (N_25505,N_20681,N_19507);
or U25506 (N_25506,N_18068,N_23373);
xnor U25507 (N_25507,N_20435,N_18308);
nand U25508 (N_25508,N_19612,N_19236);
and U25509 (N_25509,N_18909,N_18961);
nand U25510 (N_25510,N_18636,N_22441);
nor U25511 (N_25511,N_18524,N_20196);
and U25512 (N_25512,N_18419,N_19545);
nor U25513 (N_25513,N_20572,N_22258);
nand U25514 (N_25514,N_21666,N_20779);
xor U25515 (N_25515,N_22687,N_22562);
nor U25516 (N_25516,N_19576,N_22469);
xnor U25517 (N_25517,N_19729,N_23479);
nand U25518 (N_25518,N_21782,N_23645);
or U25519 (N_25519,N_23144,N_22331);
or U25520 (N_25520,N_20805,N_23794);
nor U25521 (N_25521,N_21084,N_22689);
or U25522 (N_25522,N_18345,N_21185);
or U25523 (N_25523,N_21603,N_20926);
and U25524 (N_25524,N_20083,N_21914);
or U25525 (N_25525,N_22349,N_22603);
xor U25526 (N_25526,N_20702,N_20309);
and U25527 (N_25527,N_21506,N_23886);
and U25528 (N_25528,N_18322,N_20655);
or U25529 (N_25529,N_18255,N_19871);
nand U25530 (N_25530,N_20788,N_23155);
or U25531 (N_25531,N_20925,N_20595);
nor U25532 (N_25532,N_18541,N_18683);
xor U25533 (N_25533,N_18626,N_23420);
xnor U25534 (N_25534,N_19296,N_19984);
nand U25535 (N_25535,N_22979,N_18016);
nor U25536 (N_25536,N_23128,N_20068);
and U25537 (N_25537,N_22102,N_23647);
or U25538 (N_25538,N_18347,N_22508);
or U25539 (N_25539,N_20862,N_23749);
and U25540 (N_25540,N_23190,N_21400);
or U25541 (N_25541,N_18773,N_23329);
nand U25542 (N_25542,N_20751,N_18065);
nor U25543 (N_25543,N_23933,N_23791);
nor U25544 (N_25544,N_23902,N_22715);
nand U25545 (N_25545,N_19301,N_19944);
nor U25546 (N_25546,N_19526,N_18169);
nand U25547 (N_25547,N_18723,N_19066);
xor U25548 (N_25548,N_23581,N_20863);
nor U25549 (N_25549,N_18703,N_21762);
xnor U25550 (N_25550,N_19520,N_22097);
xor U25551 (N_25551,N_22823,N_22806);
and U25552 (N_25552,N_18430,N_20975);
and U25553 (N_25553,N_20668,N_19251);
xor U25554 (N_25554,N_20665,N_21957);
xnor U25555 (N_25555,N_20029,N_22371);
xnor U25556 (N_25556,N_21848,N_20305);
or U25557 (N_25557,N_23950,N_19743);
nor U25558 (N_25558,N_20911,N_19651);
or U25559 (N_25559,N_20043,N_22878);
and U25560 (N_25560,N_23065,N_21191);
nor U25561 (N_25561,N_21124,N_19414);
nor U25562 (N_25562,N_22844,N_21929);
nor U25563 (N_25563,N_23312,N_21464);
and U25564 (N_25564,N_23545,N_18515);
and U25565 (N_25565,N_19826,N_21112);
and U25566 (N_25566,N_21048,N_19289);
or U25567 (N_25567,N_18202,N_21359);
nor U25568 (N_25568,N_18542,N_21305);
nand U25569 (N_25569,N_23582,N_23476);
and U25570 (N_25570,N_18010,N_19176);
nor U25571 (N_25571,N_23482,N_18337);
and U25572 (N_25572,N_23055,N_19245);
nand U25573 (N_25573,N_22821,N_20177);
xnor U25574 (N_25574,N_20729,N_18333);
or U25575 (N_25575,N_19708,N_18137);
xor U25576 (N_25576,N_23546,N_23156);
xnor U25577 (N_25577,N_18327,N_21968);
nor U25578 (N_25578,N_22553,N_19397);
or U25579 (N_25579,N_22497,N_19208);
and U25580 (N_25580,N_18033,N_20088);
nand U25581 (N_25581,N_23445,N_23600);
or U25582 (N_25582,N_20734,N_19932);
nand U25583 (N_25583,N_20448,N_21756);
nand U25584 (N_25584,N_22030,N_21014);
xnor U25585 (N_25585,N_18940,N_18372);
and U25586 (N_25586,N_18598,N_23244);
xor U25587 (N_25587,N_18304,N_22701);
nand U25588 (N_25588,N_23179,N_19478);
and U25589 (N_25589,N_20658,N_19575);
xnor U25590 (N_25590,N_21940,N_19265);
nor U25591 (N_25591,N_22241,N_21332);
and U25592 (N_25592,N_21467,N_20740);
or U25593 (N_25593,N_22597,N_21916);
and U25594 (N_25594,N_18758,N_19881);
or U25595 (N_25595,N_21942,N_19416);
xor U25596 (N_25596,N_20457,N_21407);
nand U25597 (N_25597,N_18483,N_22117);
or U25598 (N_25598,N_20744,N_19408);
xor U25599 (N_25599,N_19464,N_22250);
nand U25600 (N_25600,N_20685,N_22877);
nor U25601 (N_25601,N_18071,N_23748);
nor U25602 (N_25602,N_22870,N_18922);
or U25603 (N_25603,N_22167,N_18707);
or U25604 (N_25604,N_19879,N_20431);
and U25605 (N_25605,N_22743,N_22085);
nand U25606 (N_25606,N_19278,N_22561);
nor U25607 (N_25607,N_18734,N_23927);
nand U25608 (N_25608,N_23074,N_19106);
nand U25609 (N_25609,N_21092,N_22392);
and U25610 (N_25610,N_21618,N_19002);
xnor U25611 (N_25611,N_21541,N_22324);
and U25612 (N_25612,N_18741,N_23224);
nand U25613 (N_25613,N_18361,N_23576);
and U25614 (N_25614,N_19728,N_19726);
nand U25615 (N_25615,N_20536,N_23678);
nand U25616 (N_25616,N_22277,N_21509);
nor U25617 (N_25617,N_19565,N_22907);
and U25618 (N_25618,N_19352,N_19785);
nor U25619 (N_25619,N_18892,N_21026);
xnor U25620 (N_25620,N_22972,N_19283);
and U25621 (N_25621,N_19721,N_22693);
nand U25622 (N_25622,N_22574,N_22703);
nand U25623 (N_25623,N_23770,N_23732);
xnor U25624 (N_25624,N_22118,N_22898);
and U25625 (N_25625,N_22700,N_21816);
or U25626 (N_25626,N_22943,N_18615);
or U25627 (N_25627,N_21066,N_18567);
xnor U25628 (N_25628,N_18444,N_21443);
nand U25629 (N_25629,N_23403,N_20792);
or U25630 (N_25630,N_21355,N_22662);
nand U25631 (N_25631,N_19681,N_19022);
nor U25632 (N_25632,N_19324,N_21152);
xor U25633 (N_25633,N_20856,N_23395);
nor U25634 (N_25634,N_23589,N_18321);
nand U25635 (N_25635,N_20171,N_21820);
nor U25636 (N_25636,N_22708,N_22056);
xor U25637 (N_25637,N_20877,N_18302);
or U25638 (N_25638,N_18295,N_23148);
xnor U25639 (N_25639,N_20582,N_23728);
or U25640 (N_25640,N_21889,N_18644);
xnor U25641 (N_25641,N_23785,N_22647);
and U25642 (N_25642,N_23152,N_20820);
or U25643 (N_25643,N_23963,N_21996);
nor U25644 (N_25644,N_23951,N_22672);
or U25645 (N_25645,N_22904,N_19813);
or U25646 (N_25646,N_19322,N_23694);
nor U25647 (N_25647,N_23619,N_23443);
nand U25648 (N_25648,N_21679,N_22728);
and U25649 (N_25649,N_23490,N_19475);
and U25650 (N_25650,N_23674,N_19866);
or U25651 (N_25651,N_23796,N_23058);
nor U25652 (N_25652,N_19167,N_20787);
nor U25653 (N_25653,N_21476,N_23376);
nor U25654 (N_25654,N_20516,N_18287);
nand U25655 (N_25655,N_19814,N_23535);
nand U25656 (N_25656,N_19487,N_21180);
nor U25657 (N_25657,N_23966,N_22489);
nand U25658 (N_25658,N_18120,N_18651);
nor U25659 (N_25659,N_18446,N_20146);
xor U25660 (N_25660,N_21020,N_19821);
nand U25661 (N_25661,N_21209,N_18827);
or U25662 (N_25662,N_20203,N_20037);
or U25663 (N_25663,N_21846,N_21190);
and U25664 (N_25664,N_23871,N_18376);
and U25665 (N_25665,N_20291,N_23641);
and U25666 (N_25666,N_18115,N_21204);
and U25667 (N_25667,N_20200,N_19198);
xor U25668 (N_25668,N_18516,N_23873);
nand U25669 (N_25669,N_22656,N_19085);
xor U25670 (N_25670,N_23534,N_23623);
nor U25671 (N_25671,N_23707,N_22226);
nand U25672 (N_25672,N_18318,N_23741);
or U25673 (N_25673,N_21179,N_18247);
nor U25674 (N_25674,N_21906,N_21025);
nor U25675 (N_25675,N_22906,N_22549);
nand U25676 (N_25676,N_23809,N_22259);
or U25677 (N_25677,N_23300,N_21318);
nor U25678 (N_25678,N_19225,N_20440);
xor U25679 (N_25679,N_20552,N_21612);
or U25680 (N_25680,N_21148,N_23831);
or U25681 (N_25681,N_23512,N_22983);
nand U25682 (N_25682,N_20663,N_20443);
and U25683 (N_25683,N_19766,N_19335);
nor U25684 (N_25684,N_21681,N_20205);
nand U25685 (N_25685,N_19751,N_19496);
and U25686 (N_25686,N_22153,N_22506);
nand U25687 (N_25687,N_18478,N_18328);
or U25688 (N_25688,N_23568,N_20447);
nand U25689 (N_25689,N_19515,N_22945);
xor U25690 (N_25690,N_20901,N_23776);
or U25691 (N_25691,N_21808,N_22840);
nor U25692 (N_25692,N_23182,N_21095);
and U25693 (N_25693,N_18463,N_21074);
xor U25694 (N_25694,N_21315,N_22289);
xor U25695 (N_25695,N_23359,N_20119);
or U25696 (N_25696,N_21683,N_23382);
nand U25697 (N_25697,N_18466,N_20508);
xnor U25698 (N_25698,N_21743,N_20554);
xnor U25699 (N_25699,N_23747,N_22443);
xnor U25700 (N_25700,N_20396,N_20064);
and U25701 (N_25701,N_21772,N_20406);
nand U25702 (N_25702,N_21224,N_22236);
and U25703 (N_25703,N_21875,N_23100);
nor U25704 (N_25704,N_22157,N_19797);
and U25705 (N_25705,N_19824,N_21274);
or U25706 (N_25706,N_22197,N_22547);
or U25707 (N_25707,N_22799,N_23119);
nor U25708 (N_25708,N_20285,N_23189);
or U25709 (N_25709,N_19446,N_22600);
nor U25710 (N_25710,N_18046,N_21348);
or U25711 (N_25711,N_23668,N_19873);
nand U25712 (N_25712,N_18057,N_22763);
xor U25713 (N_25713,N_18582,N_21006);
xnor U25714 (N_25714,N_20994,N_22942);
or U25715 (N_25715,N_21383,N_21300);
nand U25716 (N_25716,N_23716,N_19994);
nand U25717 (N_25717,N_22283,N_19985);
nand U25718 (N_25718,N_20458,N_20072);
nor U25719 (N_25719,N_19463,N_20625);
and U25720 (N_25720,N_20939,N_22077);
nor U25721 (N_25721,N_21617,N_23547);
and U25722 (N_25722,N_18833,N_22428);
nand U25723 (N_25723,N_20223,N_23365);
nand U25724 (N_25724,N_18216,N_18721);
or U25725 (N_25725,N_22896,N_18185);
and U25726 (N_25726,N_22014,N_19946);
nor U25727 (N_25727,N_23717,N_21586);
xnor U25728 (N_25728,N_21769,N_18012);
or U25729 (N_25729,N_18876,N_21289);
nor U25730 (N_25730,N_23540,N_18730);
nor U25731 (N_25731,N_18106,N_23461);
nand U25732 (N_25732,N_20506,N_22579);
and U25733 (N_25733,N_20596,N_21304);
xor U25734 (N_25734,N_22751,N_22654);
nand U25735 (N_25735,N_23121,N_21018);
xnor U25736 (N_25736,N_19466,N_18847);
and U25737 (N_25737,N_23737,N_21963);
and U25738 (N_25738,N_19237,N_19694);
and U25739 (N_25739,N_21497,N_23079);
nor U25740 (N_25740,N_22356,N_21871);
and U25741 (N_25741,N_21513,N_20766);
or U25742 (N_25742,N_22076,N_19872);
xnor U25743 (N_25743,N_21214,N_18911);
or U25744 (N_25744,N_23029,N_18546);
nor U25745 (N_25745,N_21303,N_20411);
nand U25746 (N_25746,N_22192,N_20977);
nand U25747 (N_25747,N_20218,N_23474);
and U25748 (N_25748,N_20583,N_20701);
nor U25749 (N_25749,N_21731,N_22012);
and U25750 (N_25750,N_21052,N_22201);
nand U25751 (N_25751,N_21229,N_19611);
nor U25752 (N_25752,N_21849,N_22590);
nand U25753 (N_25753,N_18867,N_18663);
and U25754 (N_25754,N_22494,N_18095);
nand U25755 (N_25755,N_19472,N_21298);
and U25756 (N_25756,N_20356,N_22709);
nor U25757 (N_25757,N_18240,N_20704);
or U25758 (N_25758,N_23834,N_22776);
nor U25759 (N_25759,N_21943,N_18108);
and U25760 (N_25760,N_19620,N_22544);
xor U25761 (N_25761,N_23955,N_23893);
nand U25762 (N_25762,N_20092,N_21475);
nand U25763 (N_25763,N_18852,N_19904);
or U25764 (N_25764,N_20426,N_19369);
nand U25765 (N_25765,N_22413,N_19427);
xor U25766 (N_25766,N_23847,N_21575);
and U25767 (N_25767,N_19753,N_23898);
xor U25768 (N_25768,N_19778,N_21493);
nand U25769 (N_25769,N_20504,N_19907);
xor U25770 (N_25770,N_22116,N_22142);
nand U25771 (N_25771,N_21511,N_21441);
nor U25772 (N_25772,N_23632,N_18139);
and U25773 (N_25773,N_23405,N_22704);
or U25774 (N_25774,N_19425,N_20672);
and U25775 (N_25775,N_18044,N_18838);
xor U25776 (N_25776,N_19403,N_21433);
xor U25777 (N_25777,N_23351,N_22861);
or U25778 (N_25778,N_18209,N_19528);
nand U25779 (N_25779,N_21488,N_23731);
nand U25780 (N_25780,N_18862,N_18398);
nor U25781 (N_25781,N_23110,N_21607);
or U25782 (N_25782,N_18616,N_18280);
xor U25783 (N_25783,N_21595,N_20180);
nand U25784 (N_25784,N_18349,N_18831);
nor U25785 (N_25785,N_18709,N_18526);
xor U25786 (N_25786,N_20892,N_22625);
nand U25787 (N_25787,N_21621,N_19264);
nand U25788 (N_25788,N_21423,N_23870);
xnor U25789 (N_25789,N_23414,N_22845);
and U25790 (N_25790,N_20913,N_23629);
nor U25791 (N_25791,N_18568,N_22816);
nor U25792 (N_25792,N_20109,N_21768);
and U25793 (N_25793,N_22670,N_22551);
nand U25794 (N_25794,N_23529,N_23807);
or U25795 (N_25795,N_19939,N_23143);
nand U25796 (N_25796,N_19820,N_22404);
nor U25797 (N_25797,N_22769,N_20523);
nor U25798 (N_25798,N_18305,N_20469);
or U25799 (N_25799,N_23652,N_21390);
or U25800 (N_25800,N_22271,N_23257);
xnor U25801 (N_25801,N_20413,N_22855);
or U25802 (N_25802,N_20094,N_22049);
xnor U25803 (N_25803,N_20014,N_22433);
nand U25804 (N_25804,N_19122,N_22332);
nand U25805 (N_25805,N_19310,N_20310);
or U25806 (N_25806,N_19972,N_22659);
nor U25807 (N_25807,N_21397,N_21125);
nand U25808 (N_25808,N_20379,N_18021);
and U25809 (N_25809,N_20494,N_21920);
and U25810 (N_25810,N_23751,N_20895);
or U25811 (N_25811,N_19989,N_18936);
or U25812 (N_25812,N_21110,N_19627);
nor U25813 (N_25813,N_18342,N_22069);
nand U25814 (N_25814,N_21130,N_21415);
nor U25815 (N_25815,N_20969,N_23328);
and U25816 (N_25816,N_20794,N_21365);
or U25817 (N_25817,N_22267,N_20604);
nor U25818 (N_25818,N_18279,N_20007);
or U25819 (N_25819,N_20303,N_21034);
nor U25820 (N_25820,N_20419,N_23782);
and U25821 (N_25821,N_18343,N_23092);
and U25822 (N_25822,N_18962,N_23860);
nor U25823 (N_25823,N_22011,N_21442);
or U25824 (N_25824,N_20551,N_20827);
xnor U25825 (N_25825,N_21368,N_20871);
nand U25826 (N_25826,N_19205,N_20144);
nand U25827 (N_25827,N_23837,N_18260);
xnor U25828 (N_25828,N_21055,N_19045);
xor U25829 (N_25829,N_20403,N_20530);
and U25830 (N_25830,N_19258,N_18731);
xnor U25831 (N_25831,N_21613,N_18643);
or U25832 (N_25832,N_21324,N_21043);
xor U25833 (N_25833,N_22846,N_18865);
nor U25834 (N_25834,N_18443,N_23280);
nand U25835 (N_25835,N_19649,N_18504);
xor U25836 (N_25836,N_21389,N_19930);
nand U25837 (N_25837,N_18138,N_22215);
or U25838 (N_25838,N_18191,N_21791);
xnor U25839 (N_25839,N_21888,N_21491);
nand U25840 (N_25840,N_23989,N_20667);
nand U25841 (N_25841,N_18127,N_18854);
xnor U25842 (N_25842,N_20915,N_23343);
xnor U25843 (N_25843,N_21233,N_21457);
and U25844 (N_25844,N_20579,N_21088);
and U25845 (N_25845,N_23109,N_18743);
xor U25846 (N_25846,N_23889,N_23844);
nor U25847 (N_25847,N_21694,N_22643);
nand U25848 (N_25848,N_22067,N_21723);
and U25849 (N_25849,N_22446,N_22711);
nor U25850 (N_25850,N_21411,N_19168);
and U25851 (N_25851,N_20345,N_19058);
and U25852 (N_25852,N_21285,N_21283);
nand U25853 (N_25853,N_18664,N_22020);
or U25854 (N_25854,N_19295,N_23663);
nor U25855 (N_25855,N_22375,N_22314);
and U25856 (N_25856,N_19244,N_23399);
nor U25857 (N_25857,N_23516,N_19660);
xnor U25858 (N_25858,N_22084,N_20889);
nand U25859 (N_25859,N_23942,N_20692);
nor U25860 (N_25860,N_19798,N_21630);
or U25861 (N_25861,N_20070,N_21085);
nand U25862 (N_25862,N_18819,N_20727);
nor U25863 (N_25863,N_22499,N_21688);
or U25864 (N_25864,N_22368,N_19210);
nand U25865 (N_25865,N_22125,N_20501);
and U25866 (N_25866,N_18949,N_18117);
nand U25867 (N_25867,N_20499,N_19955);
xnor U25868 (N_25868,N_19767,N_19535);
or U25869 (N_25869,N_19945,N_19332);
or U25870 (N_25870,N_21656,N_20857);
and U25871 (N_25871,N_20114,N_23669);
nor U25872 (N_25872,N_21806,N_22061);
nand U25873 (N_25873,N_20682,N_21421);
xnor U25874 (N_25874,N_18212,N_22178);
and U25875 (N_25875,N_22229,N_19831);
and U25876 (N_25876,N_19801,N_22257);
or U25877 (N_25877,N_23426,N_21742);
nor U25878 (N_25878,N_19961,N_23241);
and U25879 (N_25879,N_21813,N_18901);
xnor U25880 (N_25880,N_19192,N_21925);
nor U25881 (N_25881,N_20277,N_19965);
and U25882 (N_25882,N_20799,N_21969);
nand U25883 (N_25883,N_20380,N_20601);
and U25884 (N_25884,N_19284,N_20412);
nor U25885 (N_25885,N_22777,N_19874);
nor U25886 (N_25886,N_23762,N_23279);
xor U25887 (N_25887,N_18806,N_22205);
and U25888 (N_25888,N_23071,N_22955);
xnor U25889 (N_25889,N_20104,N_19525);
nand U25890 (N_25890,N_18779,N_20746);
nand U25891 (N_25891,N_23691,N_21598);
nor U25892 (N_25892,N_21132,N_22571);
nor U25893 (N_25893,N_19260,N_19172);
nand U25894 (N_25894,N_22921,N_21015);
or U25895 (N_25895,N_22176,N_23664);
xor U25896 (N_25896,N_21585,N_23038);
nor U25897 (N_25897,N_19552,N_23538);
and U25898 (N_25898,N_23454,N_23715);
nand U25899 (N_25899,N_23453,N_21282);
and U25900 (N_25900,N_19161,N_20500);
nor U25901 (N_25901,N_19433,N_23569);
nand U25902 (N_25902,N_20698,N_20160);
and U25903 (N_25903,N_23275,N_18396);
and U25904 (N_25904,N_18856,N_21881);
and U25905 (N_25905,N_20295,N_21650);
nand U25906 (N_25906,N_20076,N_18253);
and U25907 (N_25907,N_19328,N_21449);
and U25908 (N_25908,N_21166,N_21794);
nand U25909 (N_25909,N_19982,N_21387);
nor U25910 (N_25910,N_22842,N_23872);
nand U25911 (N_25911,N_22051,N_22152);
xnor U25912 (N_25912,N_20404,N_19133);
xor U25913 (N_25913,N_22293,N_21955);
nand U25914 (N_25914,N_18931,N_19641);
and U25915 (N_25915,N_22598,N_18809);
nor U25916 (N_25916,N_20984,N_19491);
xor U25917 (N_25917,N_22242,N_22666);
or U25918 (N_25918,N_20422,N_22935);
nand U25919 (N_25919,N_22710,N_23924);
xor U25920 (N_25920,N_22065,N_22485);
nand U25921 (N_25921,N_22567,N_23695);
nor U25922 (N_25922,N_18114,N_23555);
or U25923 (N_25923,N_18383,N_22420);
nand U25924 (N_25924,N_22605,N_20800);
nor U25925 (N_25925,N_20193,N_20614);
nand U25926 (N_25926,N_18434,N_21668);
or U25927 (N_25927,N_23108,N_20768);
or U25928 (N_25928,N_22238,N_21149);
nand U25929 (N_25929,N_22584,N_22430);
or U25930 (N_25930,N_21692,N_23526);
xnor U25931 (N_25931,N_21195,N_22646);
and U25932 (N_25932,N_20743,N_20736);
and U25933 (N_25933,N_21736,N_23672);
nand U25934 (N_25934,N_22119,N_18836);
or U25935 (N_25935,N_19856,N_19249);
xor U25936 (N_25936,N_20813,N_18702);
nor U25937 (N_25937,N_20558,N_22290);
xnor U25938 (N_25938,N_18873,N_18147);
xor U25939 (N_25939,N_23682,N_20065);
nand U25940 (N_25940,N_21761,N_19020);
nand U25941 (N_25941,N_19640,N_23774);
xor U25942 (N_25942,N_20777,N_21046);
nor U25943 (N_25943,N_23207,N_23378);
nand U25944 (N_25944,N_19588,N_19353);
nand U25945 (N_25945,N_21615,N_21011);
nand U25946 (N_25946,N_18415,N_19606);
or U25947 (N_25947,N_22788,N_19409);
nor U25948 (N_25948,N_19788,N_23324);
nor U25949 (N_25949,N_20611,N_22919);
or U25950 (N_25950,N_19557,N_18028);
xor U25951 (N_25951,N_19204,N_23523);
nor U25952 (N_25952,N_23048,N_19043);
nand U25953 (N_25953,N_22859,N_23370);
and U25954 (N_25954,N_21758,N_22161);
xnor U25955 (N_25955,N_22213,N_20846);
xnor U25956 (N_25956,N_19523,N_18696);
and U25957 (N_25957,N_20432,N_23242);
nand U25958 (N_25958,N_23918,N_23133);
nor U25959 (N_25959,N_22918,N_19354);
or U25960 (N_25960,N_19655,N_19558);
nand U25961 (N_25961,N_20019,N_19777);
nor U25962 (N_25962,N_21144,N_18531);
and U25963 (N_25963,N_19914,N_21974);
or U25964 (N_25964,N_22720,N_18853);
or U25965 (N_25965,N_23301,N_18618);
nand U25966 (N_25966,N_22298,N_22782);
or U25967 (N_25967,N_20568,N_20900);
xnor U25968 (N_25968,N_21658,N_23520);
nand U25969 (N_25969,N_19238,N_19864);
nand U25970 (N_25970,N_19011,N_21215);
and U25971 (N_25971,N_19583,N_19418);
or U25972 (N_25972,N_18952,N_20735);
xor U25973 (N_25973,N_18756,N_21373);
xor U25974 (N_25974,N_22452,N_23851);
xnor U25975 (N_25975,N_22028,N_22623);
nor U25976 (N_25976,N_20916,N_21608);
and U25977 (N_25977,N_18085,N_20687);
nor U25978 (N_25978,N_18620,N_18739);
xnor U25979 (N_25979,N_19039,N_20182);
and U25980 (N_25980,N_22272,N_20853);
and U25981 (N_25981,N_22611,N_22464);
nand U25982 (N_25982,N_23998,N_21780);
and U25983 (N_25983,N_23558,N_22540);
xor U25984 (N_25984,N_18824,N_20858);
nand U25985 (N_25985,N_18506,N_19094);
nand U25986 (N_25986,N_19164,N_21260);
nor U25987 (N_25987,N_19936,N_18520);
xor U25988 (N_25988,N_20616,N_19902);
and U25989 (N_25989,N_22440,N_18609);
nor U25990 (N_25990,N_20462,N_20980);
xnor U25991 (N_25991,N_18871,N_20526);
nor U25992 (N_25992,N_21567,N_19438);
nand U25993 (N_25993,N_23815,N_19307);
xnor U25994 (N_25994,N_18423,N_20003);
or U25995 (N_25995,N_18432,N_21323);
or U25996 (N_25996,N_18588,N_23679);
xnor U25997 (N_25997,N_18720,N_21691);
and U25998 (N_25998,N_23346,N_19387);
and U25999 (N_25999,N_21605,N_18780);
nor U26000 (N_26000,N_19838,N_18112);
xnor U26001 (N_26001,N_20935,N_20216);
nand U26002 (N_26002,N_18522,N_20643);
xor U26003 (N_26003,N_19752,N_20823);
xnor U26004 (N_26004,N_19091,N_20296);
or U26005 (N_26005,N_21783,N_21156);
and U26006 (N_26006,N_18938,N_20724);
nand U26007 (N_26007,N_19680,N_23781);
or U26008 (N_26008,N_19643,N_20924);
xor U26009 (N_26009,N_22609,N_18581);
xor U26010 (N_26010,N_19327,N_21106);
and U26011 (N_26011,N_18678,N_19044);
or U26012 (N_26012,N_19363,N_22093);
nor U26013 (N_26013,N_21310,N_19511);
nand U26014 (N_26014,N_22143,N_18584);
nor U26015 (N_26015,N_20999,N_21507);
nand U26016 (N_26016,N_21854,N_20453);
nand U26017 (N_26017,N_20401,N_23102);
xnor U26018 (N_26018,N_20851,N_23835);
or U26019 (N_26019,N_19046,N_22849);
nand U26020 (N_26020,N_18254,N_21414);
xor U26021 (N_26021,N_20355,N_19949);
xnor U26022 (N_26022,N_22155,N_21439);
xnor U26023 (N_26023,N_23820,N_18692);
or U26024 (N_26024,N_18290,N_23167);
or U26025 (N_26025,N_20006,N_21790);
or U26026 (N_26026,N_18801,N_22487);
xnor U26027 (N_26027,N_21789,N_18868);
nor U26028 (N_26028,N_21097,N_22876);
or U26029 (N_26029,N_19099,N_20416);
xnor U26030 (N_26030,N_18440,N_20041);
and U26031 (N_26031,N_20455,N_18394);
nand U26032 (N_26032,N_18966,N_21453);
or U26033 (N_26033,N_21836,N_23419);
xnor U26034 (N_26034,N_18324,N_22171);
nand U26035 (N_26035,N_18519,N_23830);
xor U26036 (N_26036,N_20881,N_18786);
nor U26037 (N_26037,N_20028,N_23086);
or U26038 (N_26038,N_18425,N_21838);
and U26039 (N_26039,N_23845,N_22664);
nand U26040 (N_26040,N_23984,N_21654);
and U26041 (N_26041,N_22341,N_19191);
xor U26042 (N_26042,N_20166,N_18634);
or U26043 (N_26043,N_18164,N_23990);
or U26044 (N_26044,N_22886,N_19922);
xor U26045 (N_26045,N_20354,N_23116);
xor U26046 (N_26046,N_23986,N_23117);
nor U26047 (N_26047,N_19131,N_21992);
and U26048 (N_26048,N_20890,N_18839);
or U26049 (N_26049,N_19358,N_18623);
xnor U26050 (N_26050,N_21984,N_18492);
or U26051 (N_26051,N_22491,N_19138);
nor U26052 (N_26052,N_20143,N_23268);
nand U26053 (N_26053,N_23235,N_19854);
xor U26054 (N_26054,N_18695,N_22418);
and U26055 (N_26055,N_23296,N_19685);
or U26056 (N_26056,N_19539,N_18686);
and U26057 (N_26057,N_20385,N_21720);
or U26058 (N_26058,N_20550,N_22589);
and U26059 (N_26059,N_20376,N_20749);
nand U26060 (N_26060,N_20934,N_18981);
or U26061 (N_26061,N_21496,N_19233);
nand U26062 (N_26062,N_22766,N_20544);
or U26063 (N_26063,N_20159,N_20378);
and U26064 (N_26064,N_22095,N_20445);
nand U26065 (N_26065,N_20891,N_20383);
and U26066 (N_26066,N_21346,N_22808);
or U26067 (N_26067,N_19216,N_20135);
nand U26068 (N_26068,N_23685,N_23779);
and U26069 (N_26069,N_21192,N_21971);
nand U26070 (N_26070,N_21351,N_19747);
and U26071 (N_26071,N_23580,N_23939);
and U26072 (N_26072,N_19200,N_21936);
nand U26073 (N_26073,N_18714,N_22730);
xnor U26074 (N_26074,N_18611,N_18189);
nand U26075 (N_26075,N_23693,N_18246);
or U26076 (N_26076,N_21019,N_20804);
and U26077 (N_26077,N_21878,N_23213);
xnor U26078 (N_26078,N_18144,N_19771);
and U26079 (N_26079,N_20477,N_18081);
nor U26080 (N_26080,N_18774,N_20708);
xnor U26081 (N_26081,N_18258,N_20235);
xor U26082 (N_26082,N_20627,N_19800);
and U26083 (N_26083,N_22140,N_22520);
nor U26084 (N_26084,N_18878,N_20810);
or U26085 (N_26085,N_23887,N_22974);
or U26086 (N_26086,N_20487,N_19746);
nor U26087 (N_26087,N_19469,N_23878);
nor U26088 (N_26088,N_21601,N_21687);
nand U26089 (N_26089,N_23900,N_23727);
and U26090 (N_26090,N_21927,N_19887);
and U26091 (N_26091,N_23186,N_22825);
xnor U26092 (N_26092,N_22180,N_18657);
and U26093 (N_26093,N_23417,N_18449);
or U26094 (N_26094,N_22008,N_20195);
nand U26095 (N_26095,N_22364,N_21977);
xor U26096 (N_26096,N_23725,N_19835);
nor U26097 (N_26097,N_22496,N_23447);
nand U26098 (N_26098,N_21311,N_21440);
nor U26099 (N_26099,N_20219,N_21702);
xor U26100 (N_26100,N_22232,N_18458);
or U26101 (N_26101,N_20651,N_20795);
nor U26102 (N_26102,N_20212,N_18276);
xnor U26103 (N_26103,N_21760,N_20562);
and U26104 (N_26104,N_20013,N_23455);
nand U26105 (N_26105,N_19501,N_23295);
xnor U26106 (N_26106,N_23250,N_20974);
nand U26107 (N_26107,N_23353,N_22791);
or U26108 (N_26108,N_23877,N_20748);
nand U26109 (N_26109,N_20956,N_22642);
and U26110 (N_26110,N_23821,N_21335);
xnor U26111 (N_26111,N_20525,N_20908);
or U26112 (N_26112,N_23556,N_19281);
or U26113 (N_26113,N_18776,N_23473);
xor U26114 (N_26114,N_19789,N_22066);
nor U26115 (N_26115,N_22092,N_20326);
xor U26116 (N_26116,N_18473,N_21338);
or U26117 (N_26117,N_18317,N_21322);
nor U26118 (N_26118,N_21634,N_21714);
and U26119 (N_26119,N_20542,N_23052);
nor U26120 (N_26120,N_23192,N_19977);
nor U26121 (N_26121,N_23188,N_22275);
nand U26122 (N_26122,N_22340,N_21716);
xnor U26123 (N_26123,N_22614,N_18435);
nor U26124 (N_26124,N_20247,N_19437);
nor U26125 (N_26125,N_23364,N_22717);
xnor U26126 (N_26126,N_21651,N_21119);
nand U26127 (N_26127,N_19613,N_23838);
xnor U26128 (N_26128,N_22800,N_22318);
and U26129 (N_26129,N_21422,N_22517);
xnor U26130 (N_26130,N_22515,N_20485);
nor U26131 (N_26131,N_21357,N_18802);
xor U26132 (N_26132,N_19521,N_21847);
nor U26133 (N_26133,N_20079,N_23001);
xor U26134 (N_26134,N_19850,N_19166);
xnor U26135 (N_26135,N_23962,N_18485);
nand U26136 (N_26136,N_21367,N_18959);
and U26137 (N_26137,N_19339,N_23388);
xnor U26138 (N_26138,N_19519,N_22057);
nor U26139 (N_26139,N_22108,N_18445);
and U26140 (N_26140,N_19562,N_19671);
nand U26141 (N_26141,N_20363,N_20465);
nor U26142 (N_26142,N_23000,N_20807);
nor U26143 (N_26143,N_20382,N_20312);
nand U26144 (N_26144,N_21142,N_21793);
nor U26145 (N_26145,N_18177,N_23611);
nor U26146 (N_26146,N_23702,N_18291);
nor U26147 (N_26147,N_20770,N_22648);
nand U26148 (N_26148,N_21637,N_18920);
xnor U26149 (N_26149,N_20621,N_22820);
xnor U26150 (N_26150,N_22819,N_21966);
and U26151 (N_26151,N_22694,N_22047);
and U26152 (N_26152,N_20757,N_22223);
or U26153 (N_26153,N_22927,N_21949);
nand U26154 (N_26154,N_18460,N_19506);
or U26155 (N_26155,N_19118,N_23397);
nand U26156 (N_26156,N_20852,N_20771);
or U26157 (N_26157,N_23518,N_18501);
nand U26158 (N_26158,N_23066,N_19722);
nor U26159 (N_26159,N_23811,N_20459);
or U26160 (N_26160,N_22243,N_21983);
and U26161 (N_26161,N_20051,N_19978);
nor U26162 (N_26162,N_21545,N_20726);
xor U26163 (N_26163,N_19256,N_20507);
or U26164 (N_26164,N_19815,N_20009);
nor U26165 (N_26165,N_18052,N_18908);
and U26166 (N_26166,N_18877,N_20906);
nor U26167 (N_26167,N_19218,N_23175);
or U26168 (N_26168,N_22973,N_22468);
or U26169 (N_26169,N_20319,N_20134);
or U26170 (N_26170,N_22188,N_22780);
and U26171 (N_26171,N_18123,N_18418);
nand U26172 (N_26172,N_19684,N_18559);
xor U26173 (N_26173,N_20870,N_18479);
and U26174 (N_26174,N_20173,N_21417);
nand U26175 (N_26175,N_20979,N_23330);
or U26176 (N_26176,N_18211,N_20532);
or U26177 (N_26177,N_18379,N_18676);
and U26178 (N_26178,N_21027,N_21746);
nand U26179 (N_26179,N_18735,N_21363);
xor U26180 (N_26180,N_22902,N_20117);
and U26181 (N_26181,N_21695,N_19761);
and U26182 (N_26182,N_23276,N_21905);
nor U26183 (N_26183,N_22853,N_22214);
or U26184 (N_26184,N_21945,N_19623);
or U26185 (N_26185,N_20571,N_23755);
and U26186 (N_26186,N_19503,N_22256);
xnor U26187 (N_26187,N_18294,N_23237);
or U26188 (N_26188,N_23689,N_18025);
xnor U26189 (N_26189,N_21879,N_23471);
or U26190 (N_26190,N_18193,N_20033);
and U26191 (N_26191,N_22779,N_18213);
nor U26192 (N_26192,N_21029,N_19146);
and U26193 (N_26193,N_19704,N_18167);
nor U26194 (N_26194,N_19010,N_19981);
and U26195 (N_26195,N_22419,N_22075);
or U26196 (N_26196,N_23823,N_22281);
xnor U26197 (N_26197,N_19459,N_18596);
nor U26198 (N_26198,N_23750,N_18042);
nand U26199 (N_26199,N_20211,N_23840);
nor U26200 (N_26200,N_19843,N_20024);
xnor U26201 (N_26201,N_21965,N_18599);
nand U26202 (N_26202,N_23789,N_21766);
xor U26203 (N_26203,N_20716,N_23059);
nor U26204 (N_26204,N_19120,N_22193);
nor U26205 (N_26205,N_21524,N_23793);
and U26206 (N_26206,N_18973,N_23979);
xor U26207 (N_26207,N_18916,N_22512);
and U26208 (N_26208,N_21237,N_18851);
xnor U26209 (N_26209,N_21671,N_22353);
or U26210 (N_26210,N_18009,N_20620);
or U26211 (N_26211,N_20644,N_21804);
or U26212 (N_26212,N_20880,N_23890);
or U26213 (N_26213,N_21451,N_18551);
nor U26214 (N_26214,N_21633,N_23943);
xor U26215 (N_26215,N_19400,N_22634);
nand U26216 (N_26216,N_19149,N_23408);
nor U26217 (N_26217,N_18375,N_18314);
nor U26218 (N_26218,N_21883,N_19197);
and U26219 (N_26219,N_22908,N_19712);
nor U26220 (N_26220,N_18426,N_20631);
xnor U26221 (N_26221,N_22262,N_21919);
or U26222 (N_26222,N_22220,N_18574);
nor U26223 (N_26223,N_22058,N_20150);
xnor U26224 (N_26224,N_21432,N_22621);
or U26225 (N_26225,N_23440,N_18357);
nor U26226 (N_26226,N_18210,N_21210);
and U26227 (N_26227,N_20121,N_21773);
and U26228 (N_26228,N_20402,N_22122);
nor U26229 (N_26229,N_18775,N_22130);
nor U26230 (N_26230,N_22760,N_18481);
nor U26231 (N_26231,N_20991,N_22401);
xnor U26232 (N_26232,N_19768,N_23810);
or U26233 (N_26233,N_23705,N_19885);
nand U26234 (N_26234,N_22007,N_18941);
xor U26235 (N_26235,N_21950,N_20967);
nor U26236 (N_26236,N_23677,N_20707);
and U26237 (N_26237,N_20127,N_19139);
or U26238 (N_26238,N_23539,N_22177);
nand U26239 (N_26239,N_23045,N_18982);
or U26240 (N_26240,N_19738,N_23541);
and U26241 (N_26241,N_21352,N_23249);
and U26242 (N_26242,N_18656,N_19402);
or U26243 (N_26243,N_22109,N_23230);
xor U26244 (N_26244,N_20428,N_21823);
or U26245 (N_26245,N_20834,N_21436);
nand U26246 (N_26246,N_21361,N_19136);
and U26247 (N_26247,N_20854,N_21396);
or U26248 (N_26248,N_19719,N_22798);
nand U26249 (N_26249,N_18603,N_22622);
nand U26250 (N_26250,N_23208,N_22794);
nand U26251 (N_26251,N_19605,N_21388);
and U26252 (N_26252,N_22261,N_18084);
nor U26253 (N_26253,N_21393,N_18606);
nor U26254 (N_26254,N_22325,N_20653);
nand U26255 (N_26255,N_21709,N_21301);
and U26256 (N_26256,N_21676,N_23775);
nor U26257 (N_26257,N_18677,N_19107);
nor U26258 (N_26258,N_23464,N_21864);
and U26259 (N_26259,N_21047,N_19517);
nor U26260 (N_26260,N_20387,N_23323);
nor U26261 (N_26261,N_21398,N_19715);
or U26262 (N_26262,N_23090,N_18078);
or U26263 (N_26263,N_18262,N_23897);
xnor U26264 (N_26264,N_20100,N_18905);
xnor U26265 (N_26265,N_18178,N_22168);
xnor U26266 (N_26266,N_19570,N_23335);
xnor U26267 (N_26267,N_18439,N_23856);
nor U26268 (N_26268,N_21970,N_19702);
nor U26269 (N_26269,N_20641,N_20359);
nand U26270 (N_26270,N_22991,N_23033);
and U26271 (N_26271,N_19622,N_21972);
nand U26272 (N_26272,N_23993,N_23718);
nand U26273 (N_26273,N_22740,N_22725);
nand U26274 (N_26274,N_18885,N_20050);
nor U26275 (N_26275,N_18306,N_23009);
nand U26276 (N_26276,N_20270,N_19672);
and U26277 (N_26277,N_20444,N_19348);
and U26278 (N_26278,N_22461,N_23209);
and U26279 (N_26279,N_21343,N_20175);
or U26280 (N_26280,N_19581,N_22852);
xnor U26281 (N_26281,N_23959,N_18850);
or U26282 (N_26282,N_18148,N_19227);
nand U26283 (N_26283,N_22971,N_20046);
or U26284 (N_26284,N_18274,N_18529);
nand U26285 (N_26285,N_19014,N_22315);
xnor U26286 (N_26286,N_18225,N_19998);
or U26287 (N_26287,N_21222,N_21900);
xor U26288 (N_26288,N_19277,N_22834);
and U26289 (N_26289,N_21841,N_19819);
xor U26290 (N_26290,N_23194,N_22789);
xnor U26291 (N_26291,N_21775,N_20914);
xor U26292 (N_26292,N_21801,N_22104);
nand U26293 (N_26293,N_22525,N_22518);
xnor U26294 (N_26294,N_19580,N_21645);
nand U26295 (N_26295,N_20410,N_18869);
nand U26296 (N_26296,N_22146,N_19183);
nand U26297 (N_26297,N_18149,N_23819);
nand U26298 (N_26298,N_18635,N_19067);
nor U26299 (N_26299,N_21127,N_22767);
nor U26300 (N_26300,N_23004,N_19151);
nand U26301 (N_26301,N_20332,N_22952);
xnor U26302 (N_26302,N_20263,N_19723);
or U26303 (N_26303,N_21748,N_23808);
and U26304 (N_26304,N_20555,N_22185);
nor U26305 (N_26305,N_19393,N_19173);
nand U26306 (N_26306,N_22966,N_23625);
and U26307 (N_26307,N_23317,N_20599);
xor U26308 (N_26308,N_19145,N_23868);
xor U26309 (N_26309,N_18467,N_20534);
nand U26310 (N_26310,N_21891,N_19143);
xnor U26311 (N_26311,N_18156,N_20798);
nand U26312 (N_26312,N_18586,N_21494);
xor U26313 (N_26313,N_20384,N_22407);
xor U26314 (N_26314,N_23648,N_23713);
xnor U26315 (N_26315,N_19697,N_23746);
nand U26316 (N_26316,N_19550,N_19587);
nand U26317 (N_26317,N_23483,N_21430);
nor U26318 (N_26318,N_23721,N_19836);
or U26319 (N_26319,N_20176,N_23437);
nand U26320 (N_26320,N_23875,N_19262);
or U26321 (N_26321,N_22560,N_23825);
or U26322 (N_26322,N_21862,N_20762);
xor U26323 (N_26323,N_20570,N_18793);
and U26324 (N_26324,N_19498,N_18512);
and U26325 (N_26325,N_22070,N_23239);
and U26326 (N_26326,N_19842,N_21502);
nand U26327 (N_26327,N_18918,N_21684);
and U26328 (N_26328,N_21811,N_19957);
xnor U26329 (N_26329,N_23738,N_18069);
nand U26330 (N_26330,N_20181,N_22126);
and U26331 (N_26331,N_18094,N_22810);
or U26332 (N_26332,N_23389,N_19597);
nor U26333 (N_26333,N_19652,N_19600);
xor U26334 (N_26334,N_18018,N_22726);
xnor U26335 (N_26335,N_21540,N_19928);
or U26336 (N_26336,N_20845,N_22529);
and U26337 (N_26337,N_20283,N_19954);
xor U26338 (N_26338,N_18080,N_18592);
and U26339 (N_26339,N_18617,N_23916);
nand U26340 (N_26340,N_22063,N_19465);
nand U26341 (N_26341,N_20952,N_19656);
or U26342 (N_26342,N_19374,N_19695);
and U26343 (N_26343,N_18203,N_18970);
nor U26344 (N_26344,N_20968,N_22247);
nand U26345 (N_26345,N_19263,N_20824);
nor U26346 (N_26346,N_22074,N_21646);
nand U26347 (N_26347,N_23583,N_23544);
or U26348 (N_26348,N_23468,N_23882);
xor U26349 (N_26349,N_22931,N_20535);
nand U26350 (N_26350,N_18553,N_18608);
nor U26351 (N_26351,N_18917,N_22086);
and U26352 (N_26352,N_23489,N_22377);
nand U26353 (N_26353,N_19677,N_23772);
xnor U26354 (N_26354,N_21316,N_20442);
nand U26355 (N_26355,N_20878,N_20776);
and U26356 (N_26356,N_18544,N_18842);
nand U26357 (N_26357,N_20998,N_23552);
and U26358 (N_26358,N_20405,N_19975);
xor U26359 (N_26359,N_21812,N_20786);
xnor U26360 (N_26360,N_20279,N_22797);
xnor U26361 (N_26361,N_21250,N_20297);
xnor U26362 (N_26362,N_20317,N_18360);
or U26363 (N_26363,N_20753,N_22933);
xor U26364 (N_26364,N_18764,N_19703);
nand U26365 (N_26365,N_21412,N_22412);
nand U26366 (N_26366,N_22889,N_18242);
xor U26367 (N_26367,N_19445,N_22832);
or U26368 (N_26368,N_19128,N_20113);
nor U26369 (N_26369,N_19489,N_19291);
xnor U26370 (N_26370,N_18912,N_19100);
xor U26371 (N_26371,N_18366,N_20336);
or U26372 (N_26372,N_23948,N_20129);
or U26373 (N_26373,N_20932,N_22249);
nand U26374 (N_26374,N_22650,N_19135);
nor U26375 (N_26375,N_21273,N_18358);
nor U26376 (N_26376,N_23151,N_20308);
nand U26377 (N_26377,N_22535,N_23327);
nand U26378 (N_26378,N_19474,N_18013);
nand U26379 (N_26379,N_21312,N_21843);
or U26380 (N_26380,N_18083,N_20936);
xnor U26381 (N_26381,N_21153,N_18427);
nand U26382 (N_26382,N_20613,N_23662);
nand U26383 (N_26383,N_18768,N_23908);
nor U26384 (N_26384,N_23466,N_19428);
or U26385 (N_26385,N_22885,N_23354);
nor U26386 (N_26386,N_23084,N_23034);
xnor U26387 (N_26387,N_22612,N_18369);
or U26388 (N_26388,N_21225,N_20274);
or U26389 (N_26389,N_21231,N_22078);
nand U26390 (N_26390,N_18828,N_23172);
and U26391 (N_26391,N_20137,N_22199);
and U26392 (N_26392,N_20985,N_20695);
nor U26393 (N_26393,N_18221,N_18886);
and U26394 (N_26394,N_23435,N_23146);
and U26395 (N_26395,N_22736,N_19548);
xnor U26396 (N_26396,N_20133,N_19987);
and U26397 (N_26397,N_23391,N_19318);
nor U26398 (N_26398,N_20350,N_19974);
or U26399 (N_26399,N_22862,N_21072);
nand U26400 (N_26400,N_20468,N_20947);
and U26401 (N_26401,N_19087,N_23501);
xor U26402 (N_26402,N_21466,N_22175);
nand U26403 (N_26403,N_19000,N_19089);
and U26404 (N_26404,N_18370,N_19865);
xnor U26405 (N_26405,N_22292,N_18968);
xnor U26406 (N_26406,N_22835,N_22787);
or U26407 (N_26407,N_23404,N_18881);
xor U26408 (N_26408,N_21886,N_21935);
nand U26409 (N_26409,N_19174,N_21251);
or U26410 (N_26410,N_18421,N_21333);
and U26411 (N_26411,N_19001,N_22166);
nand U26412 (N_26412,N_23736,N_22661);
nand U26413 (N_26413,N_21636,N_21126);
xnor U26414 (N_26414,N_22219,N_23356);
or U26415 (N_26415,N_22891,N_20731);
or U26416 (N_26416,N_23502,N_23082);
nand U26417 (N_26417,N_19422,N_21375);
xor U26418 (N_26418,N_23015,N_22839);
nand U26419 (N_26419,N_21376,N_23184);
or U26420 (N_26420,N_21529,N_23700);
nor U26421 (N_26421,N_20184,N_18482);
nor U26422 (N_26422,N_18344,N_19654);
or U26423 (N_26423,N_18859,N_21386);
xor U26424 (N_26424,N_20292,N_23124);
xnor U26425 (N_26425,N_22447,N_20619);
nor U26426 (N_26426,N_23881,N_21591);
xor U26427 (N_26427,N_19774,N_23687);
or U26428 (N_26428,N_20226,N_22381);
xnor U26429 (N_26429,N_22004,N_19298);
nand U26430 (N_26430,N_21377,N_22451);
and U26431 (N_26431,N_21678,N_20078);
nor U26432 (N_26432,N_22295,N_19909);
or U26433 (N_26433,N_18413,N_22399);
or U26434 (N_26434,N_19364,N_20628);
xnor U26435 (N_26435,N_23418,N_19223);
xnor U26436 (N_26436,N_22500,N_18991);
or U26437 (N_26437,N_19250,N_22696);
nor U26438 (N_26438,N_20188,N_23928);
or U26439 (N_26439,N_23494,N_18293);
xor U26440 (N_26440,N_19564,N_18158);
nor U26441 (N_26441,N_20933,N_22771);
xnor U26442 (N_26442,N_20138,N_21727);
nor U26443 (N_26443,N_23292,N_18122);
nand U26444 (N_26444,N_23352,N_21294);
xnor U26445 (N_26445,N_22129,N_18976);
nand U26446 (N_26446,N_20244,N_18348);
and U26447 (N_26447,N_21427,N_20606);
nand U26448 (N_26448,N_23610,N_22225);
or U26449 (N_26449,N_20873,N_19394);
xor U26450 (N_26450,N_20347,N_18447);
nand U26451 (N_26451,N_19615,N_21017);
and U26452 (N_26452,N_18649,N_20349);
nor U26453 (N_26453,N_20339,N_18124);
or U26454 (N_26454,N_20098,N_19337);
nor U26455 (N_26455,N_18963,N_19799);
nand U26456 (N_26456,N_20944,N_19254);
or U26457 (N_26457,N_20464,N_18229);
xor U26458 (N_26458,N_20360,N_19370);
and U26459 (N_26459,N_18919,N_21796);
or U26460 (N_26460,N_18890,N_19690);
xor U26461 (N_26461,N_19549,N_20229);
xor U26462 (N_26462,N_23013,N_18543);
nand U26463 (N_26463,N_22900,N_20035);
xor U26464 (N_26464,N_20608,N_22775);
nor U26465 (N_26465,N_18116,N_22304);
nand U26466 (N_26466,N_23446,N_21174);
nand U26467 (N_26467,N_18757,N_23684);
nor U26468 (N_26468,N_21259,N_18243);
and U26469 (N_26469,N_22090,N_23078);
nor U26470 (N_26470,N_19013,N_18233);
and U26471 (N_26471,N_21170,N_18450);
or U26472 (N_26472,N_19368,N_21877);
or U26473 (N_26473,N_18330,N_23081);
or U26474 (N_26474,N_23381,N_22796);
nand U26475 (N_26475,N_22498,N_19042);
nand U26476 (N_26476,N_18014,N_18452);
xnor U26477 (N_26477,N_18352,N_18960);
and U26478 (N_26478,N_21242,N_20056);
xnor U26479 (N_26479,N_23211,N_18746);
or U26480 (N_26480,N_23788,N_22173);
and U26481 (N_26481,N_21113,N_19960);
nand U26482 (N_26482,N_22465,N_21778);
or U26483 (N_26483,N_18979,N_21065);
or U26484 (N_26484,N_18732,N_23996);
and U26485 (N_26485,N_18410,N_18863);
nand U26486 (N_26486,N_18214,N_23970);
nand U26487 (N_26487,N_20782,N_22424);
and U26488 (N_26488,N_20342,N_18091);
and U26489 (N_26489,N_23326,N_18698);
nand U26490 (N_26490,N_20294,N_22990);
and U26491 (N_26491,N_21486,N_20546);
nand U26492 (N_26492,N_21580,N_19109);
or U26493 (N_26493,N_20531,N_20107);
nor U26494 (N_26494,N_22686,N_19638);
and U26495 (N_26495,N_22987,N_18672);
nor U26496 (N_26496,N_23912,N_22649);
nand U26497 (N_26497,N_20152,N_21767);
xnor U26498 (N_26498,N_20819,N_23310);
xor U26499 (N_26499,N_20472,N_19431);
nor U26500 (N_26500,N_21573,N_21752);
nand U26501 (N_26501,N_22145,N_19280);
and U26502 (N_26502,N_19226,N_23958);
nor U26503 (N_26503,N_21863,N_20869);
nor U26504 (N_26504,N_19219,N_19061);
or U26505 (N_26505,N_20706,N_18226);
or U26506 (N_26506,N_23372,N_22305);
nand U26507 (N_26507,N_23322,N_21517);
nor U26508 (N_26508,N_18404,N_20893);
nand U26509 (N_26509,N_21249,N_22083);
or U26510 (N_26510,N_18975,N_21146);
nor U26511 (N_26511,N_20105,N_22478);
and U26512 (N_26512,N_22174,N_18387);
xor U26513 (N_26513,N_22016,N_20797);
nor U26514 (N_26514,N_20149,N_22864);
nor U26515 (N_26515,N_18196,N_22922);
nor U26516 (N_26516,N_20042,N_18325);
or U26517 (N_26517,N_23366,N_20467);
nor U26518 (N_26518,N_23290,N_20289);
or U26519 (N_26519,N_18230,N_22665);
nor U26520 (N_26520,N_21973,N_18538);
nand U26521 (N_26521,N_18310,N_23814);
nand U26522 (N_26522,N_22601,N_18297);
and U26523 (N_26523,N_23177,N_21893);
nand U26524 (N_26524,N_21826,N_18744);
xor U26525 (N_26525,N_20940,N_18468);
nor U26526 (N_26526,N_23262,N_20340);
or U26527 (N_26527,N_19476,N_19762);
xor U26528 (N_26528,N_23974,N_22024);
and U26529 (N_26529,N_22300,N_23413);
or U26530 (N_26530,N_23508,N_18713);
or U26531 (N_26531,N_21946,N_20683);
xor U26532 (N_26532,N_23350,N_23743);
and U26533 (N_26533,N_18965,N_22563);
xnor U26534 (N_26534,N_19794,N_20626);
or U26535 (N_26535,N_18787,N_22043);
nor U26536 (N_26536,N_20742,N_18051);
or U26537 (N_26537,N_20922,N_23261);
and U26538 (N_26538,N_23892,N_22732);
nor U26539 (N_26539,N_22892,N_19442);
and U26540 (N_26540,N_23169,N_18477);
xor U26541 (N_26541,N_23349,N_19362);
xnor U26542 (N_26542,N_19750,N_19903);
and U26543 (N_26543,N_21558,N_22389);
and U26544 (N_26544,N_18857,N_23588);
and U26545 (N_26545,N_18887,N_18411);
nor U26546 (N_26546,N_20983,N_21522);
and U26547 (N_26547,N_19019,N_18066);
or U26548 (N_26548,N_21548,N_18943);
nor U26549 (N_26549,N_23168,N_23215);
xor U26550 (N_26550,N_21230,N_23661);
nand U26551 (N_26551,N_19626,N_22462);
or U26552 (N_26552,N_18150,N_21988);
nand U26553 (N_26553,N_23406,N_20018);
and U26554 (N_26554,N_20495,N_20399);
nand U26555 (N_26555,N_23286,N_21626);
nand U26556 (N_26556,N_20463,N_21372);
and U26557 (N_26557,N_22042,N_19201);
nor U26558 (N_26558,N_21049,N_18600);
and U26559 (N_26559,N_22957,N_22724);
or U26560 (N_26560,N_20290,N_23248);
and U26561 (N_26561,N_23452,N_23801);
nor U26562 (N_26562,N_19185,N_23070);
nand U26563 (N_26563,N_20115,N_21521);
nand U26564 (N_26564,N_19004,N_19905);
and U26565 (N_26565,N_20545,N_19188);
nand U26566 (N_26566,N_20817,N_22027);
nand U26567 (N_26567,N_23430,N_19434);
nor U26568 (N_26568,N_20140,N_22809);
or U26569 (N_26569,N_21985,N_23913);
xor U26570 (N_26570,N_21958,N_22053);
nand U26571 (N_26571,N_19224,N_19455);
nor U26572 (N_26572,N_18286,N_21730);
or U26573 (N_26573,N_22575,N_18151);
nor U26574 (N_26574,N_23282,N_21685);
or U26575 (N_26575,N_23905,N_19786);
nand U26576 (N_26576,N_18589,N_22783);
and U26577 (N_26577,N_19036,N_22218);
nand U26578 (N_26578,N_22431,N_20816);
or U26579 (N_26579,N_20721,N_18861);
and U26580 (N_26580,N_21140,N_18320);
or U26581 (N_26581,N_18602,N_22619);
nor U26582 (N_26582,N_19559,N_21235);
nand U26583 (N_26583,N_21045,N_21786);
nor U26584 (N_26584,N_21171,N_18269);
nand U26585 (N_26585,N_19242,N_22526);
xnor U26586 (N_26586,N_21899,N_19048);
nor U26587 (N_26587,N_23696,N_23786);
xor U26588 (N_26588,N_20298,N_22993);
nor U26589 (N_26589,N_18625,N_21461);
or U26590 (N_26590,N_19467,N_18273);
xor U26591 (N_26591,N_22928,N_20505);
nand U26592 (N_26592,N_21741,N_21379);
nor U26593 (N_26593,N_22632,N_22851);
or U26594 (N_26594,N_22360,N_22716);
or U26595 (N_26595,N_20161,N_20278);
xor U26596 (N_26596,N_20269,N_21998);
and U26597 (N_26597,N_19556,N_22288);
xor U26598 (N_26598,N_20252,N_22260);
or U26599 (N_26599,N_23603,N_18937);
nand U26600 (N_26600,N_20831,N_22967);
nand U26601 (N_26601,N_20451,N_22521);
nor U26602 (N_26602,N_19380,N_22533);
or U26603 (N_26603,N_20338,N_18391);
nor U26604 (N_26604,N_22264,N_19077);
nand U26605 (N_26605,N_18627,N_19701);
nor U26606 (N_26606,N_20388,N_23934);
and U26607 (N_26607,N_23879,N_22668);
nor U26608 (N_26608,N_22604,N_23946);
or U26609 (N_26609,N_23630,N_20677);
nand U26610 (N_26610,N_22541,N_19818);
nor U26611 (N_26611,N_21739,N_22978);
or U26612 (N_26612,N_19593,N_18386);
nor U26613 (N_26613,N_23862,N_19700);
xor U26614 (N_26614,N_18974,N_18368);
xnor U26615 (N_26615,N_19144,N_21328);
nand U26616 (N_26616,N_23332,N_23099);
or U26617 (N_26617,N_18249,N_23360);
nand U26618 (N_26618,N_21827,N_21184);
and U26619 (N_26619,N_23044,N_20676);
nand U26620 (N_26620,N_20543,N_19213);
and U26621 (N_26621,N_21725,N_21281);
or U26622 (N_26622,N_22429,N_18508);
nand U26623 (N_26623,N_19194,N_18796);
nand U26624 (N_26624,N_20450,N_21853);
nand U26625 (N_26625,N_18930,N_19882);
nor U26626 (N_26626,N_18849,N_18517);
nor U26627 (N_26627,N_20592,N_18335);
and U26628 (N_26628,N_20369,N_23848);
and U26629 (N_26629,N_21619,N_23424);
nor U26630 (N_26630,N_23227,N_20010);
nand U26631 (N_26631,N_22678,N_23422);
or U26632 (N_26632,N_18725,N_22501);
nand U26633 (N_26633,N_18399,N_20132);
and U26634 (N_26634,N_20001,N_23187);
or U26635 (N_26635,N_21682,N_23342);
or U26636 (N_26636,N_18722,N_21663);
nor U26637 (N_26637,N_18113,N_20048);
xnor U26638 (N_26638,N_19733,N_21000);
nor U26639 (N_26639,N_22774,N_19689);
xor U26640 (N_26640,N_19976,N_23656);
or U26641 (N_26641,N_18605,N_18371);
nor U26642 (N_26642,N_20329,N_21999);
and U26643 (N_26643,N_22136,N_18607);
or U26644 (N_26644,N_20357,N_18183);
or U26645 (N_26645,N_18843,N_18300);
or U26646 (N_26646,N_19115,N_18499);
nor U26647 (N_26647,N_22699,N_23221);
nand U26648 (N_26648,N_18829,N_19931);
and U26649 (N_26649,N_23832,N_23764);
or U26650 (N_26650,N_18781,N_18684);
nor U26651 (N_26651,N_20058,N_20343);
and U26652 (N_26652,N_21167,N_22651);
nand U26653 (N_26653,N_22677,N_23680);
nor U26654 (N_26654,N_18062,N_18642);
xnor U26655 (N_26655,N_23153,N_20642);
nand U26656 (N_26656,N_22204,N_18896);
nand U26657 (N_26657,N_19755,N_20635);
nand U26658 (N_26658,N_22438,N_21931);
nor U26659 (N_26659,N_20284,N_22504);
nor U26660 (N_26660,N_18653,N_23790);
nor U26661 (N_26661,N_19983,N_22530);
or U26662 (N_26662,N_21930,N_18747);
or U26663 (N_26663,N_22252,N_22179);
and U26664 (N_26664,N_22883,N_20809);
nand U26665 (N_26665,N_18845,N_18578);
xor U26666 (N_26666,N_23659,N_21314);
nor U26667 (N_26667,N_22542,N_22607);
nand U26668 (N_26668,N_23499,N_22311);
nand U26669 (N_26669,N_22181,N_18155);
xnor U26670 (N_26670,N_20986,N_21120);
and U26671 (N_26671,N_21079,N_18003);
nand U26672 (N_26672,N_22287,N_21737);
xnor U26673 (N_26673,N_20540,N_18923);
xor U26674 (N_26674,N_22483,N_19807);
xor U26675 (N_26675,N_23113,N_21543);
nor U26676 (N_26676,N_22875,N_22352);
nor U26677 (N_26677,N_21212,N_19114);
nor U26678 (N_26678,N_20023,N_22580);
nand U26679 (N_26679,N_22328,N_22121);
nor U26680 (N_26680,N_20917,N_21075);
nor U26681 (N_26681,N_22251,N_21471);
nor U26682 (N_26682,N_20400,N_21409);
or U26683 (N_26683,N_19308,N_21472);
nand U26684 (N_26684,N_20237,N_18382);
xor U26685 (N_26685,N_22416,N_22427);
xnor U26686 (N_26686,N_19773,N_19682);
xnor U26687 (N_26687,N_23573,N_18556);
or U26688 (N_26688,N_18883,N_20720);
nor U26689 (N_26689,N_18921,N_23171);
nand U26690 (N_26690,N_22790,N_21986);
or U26691 (N_26691,N_18929,N_23757);
and U26692 (N_26692,N_23792,N_18176);
nand U26693 (N_26693,N_21583,N_19707);
or U26694 (N_26694,N_21518,N_18301);
xnor U26695 (N_26695,N_23957,N_21479);
or U26696 (N_26696,N_18992,N_20483);
nor U26697 (N_26697,N_19817,N_21196);
nand U26698 (N_26698,N_18792,N_21729);
xor U26699 (N_26699,N_21103,N_23711);
nor U26700 (N_26700,N_22681,N_22746);
or U26701 (N_26701,N_20280,N_20496);
nor U26702 (N_26702,N_19180,N_20859);
nand U26703 (N_26703,N_19573,N_18119);
nor U26704 (N_26704,N_18971,N_22507);
nand U26705 (N_26705,N_22576,N_18011);
xnor U26706 (N_26706,N_23855,N_18808);
nor U26707 (N_26707,N_18978,N_23642);
xnor U26708 (N_26708,N_22437,N_20560);
nand U26709 (N_26709,N_19908,N_19342);
xor U26710 (N_26710,N_21487,N_19748);
and U26711 (N_26711,N_20849,N_21465);
xnor U26712 (N_26712,N_20434,N_21570);
and U26713 (N_26713,N_18532,N_19063);
nor U26714 (N_26714,N_18939,N_22669);
and U26715 (N_26715,N_20071,N_18475);
nor U26716 (N_26716,N_20833,N_22248);
xor U26717 (N_26717,N_23621,N_23492);
nor U26718 (N_26718,N_21248,N_21662);
or U26719 (N_26719,N_19572,N_23204);
xnor U26720 (N_26720,N_23218,N_18956);
nand U26721 (N_26721,N_21892,N_19257);
and U26722 (N_26722,N_21176,N_19406);
nor U26723 (N_26723,N_22059,N_18772);
nor U26724 (N_26724,N_20178,N_22830);
and U26725 (N_26725,N_19234,N_22269);
nand U26726 (N_26726,N_23527,N_21894);
and U26727 (N_26727,N_21239,N_18694);
nand U26728 (N_26728,N_21320,N_22803);
nand U26729 (N_26729,N_23783,N_18265);
nand U26730 (N_26730,N_21798,N_21435);
nand U26731 (N_26731,N_23888,N_21245);
and U26732 (N_26732,N_22537,N_23503);
and U26733 (N_26733,N_18798,N_22828);
or U26734 (N_26734,N_18459,N_21547);
xor U26735 (N_26735,N_20848,N_18250);
xor U26736 (N_26736,N_20981,N_19102);
nor U26737 (N_26737,N_18967,N_22639);
and U26738 (N_26738,N_19688,N_21578);
nand U26739 (N_26739,N_19384,N_23385);
nand U26740 (N_26740,N_18089,N_21028);
and U26741 (N_26741,N_18472,N_22559);
and U26742 (N_26742,N_19294,N_19811);
nand U26743 (N_26743,N_19878,N_23983);
nand U26744 (N_26744,N_18179,N_21448);
and U26745 (N_26745,N_19485,N_22357);
and U26746 (N_26746,N_22735,N_18680);
xnor U26747 (N_26747,N_23706,N_20131);
xnor U26748 (N_26748,N_18093,N_23829);
and U26749 (N_26749,N_23371,N_23031);
or U26750 (N_26750,N_21128,N_19584);
and U26751 (N_26751,N_21552,N_18363);
xnor U26752 (N_26752,N_20096,N_20717);
nand U26753 (N_26753,N_23095,N_23745);
xor U26754 (N_26754,N_18595,N_21859);
or U26755 (N_26755,N_19193,N_19473);
or U26756 (N_26756,N_21953,N_21538);
nand U26757 (N_26757,N_18814,N_22827);
xnor U26758 (N_26758,N_18511,N_18261);
nor U26759 (N_26759,N_22459,N_21753);
nand U26760 (N_26760,N_19990,N_23798);
and U26761 (N_26761,N_20236,N_22044);
and U26762 (N_26762,N_20561,N_23288);
nand U26763 (N_26763,N_19858,N_18525);
xor U26764 (N_26764,N_18271,N_20607);
and U26765 (N_26765,N_20243,N_19060);
xor U26766 (N_26766,N_19453,N_21693);
nor U26767 (N_26767,N_21203,N_22367);
nand U26768 (N_26768,N_23896,N_23849);
and U26769 (N_26769,N_20603,N_20537);
or U26770 (N_26770,N_21960,N_23321);
nor U26771 (N_26771,N_21728,N_21349);
nor U26772 (N_26772,N_20318,N_20790);
nor U26773 (N_26773,N_19119,N_19279);
xnor U26774 (N_26774,N_19943,N_19840);
xnor U26775 (N_26775,N_22376,N_20745);
and U26776 (N_26776,N_20424,N_21350);
nor U26777 (N_26777,N_21150,N_19421);
and U26778 (N_26778,N_20123,N_20634);
or U26779 (N_26779,N_18056,N_22593);
and U26780 (N_26780,N_18474,N_18560);
and U26781 (N_26781,N_22685,N_20142);
and U26782 (N_26782,N_19440,N_22400);
nor U26783 (N_26783,N_20966,N_20527);
nand U26784 (N_26784,N_22738,N_19595);
xor U26785 (N_26785,N_23294,N_22141);
or U26786 (N_26786,N_18353,N_22772);
and U26787 (N_26787,N_20328,N_18655);
nor U26788 (N_26788,N_23714,N_18639);
or U26789 (N_26789,N_22691,N_22629);
xnor U26790 (N_26790,N_19361,N_18022);
xor U26791 (N_26791,N_23500,N_18528);
nor U26792 (N_26792,N_23157,N_23511);
and U26793 (N_26793,N_23293,N_22801);
or U26794 (N_26794,N_19883,N_21967);
or U26795 (N_26795,N_23367,N_18064);
or U26796 (N_26796,N_22805,N_23614);
xor U26797 (N_26797,N_19321,N_19683);
xnor U26798 (N_26798,N_20884,N_20732);
nor U26799 (N_26799,N_18673,N_21912);
nor U26800 (N_26800,N_23487,N_19081);
xnor U26801 (N_26801,N_23994,N_21763);
xor U26802 (N_26802,N_21340,N_22091);
or U26803 (N_26803,N_21116,N_19062);
xnor U26804 (N_26804,N_21898,N_19343);
nand U26805 (N_26805,N_23431,N_22212);
and U26806 (N_26806,N_21369,N_22470);
and U26807 (N_26807,N_23557,N_22345);
or U26808 (N_26808,N_18587,N_18880);
or U26809 (N_26809,N_21657,N_23982);
or U26810 (N_26810,N_23938,N_20513);
nor U26811 (N_26811,N_19447,N_21118);
nor U26812 (N_26812,N_21659,N_22848);
and U26813 (N_26813,N_18228,N_21139);
nand U26814 (N_26814,N_19285,N_22351);
or U26815 (N_26815,N_19518,N_19834);
or U26816 (N_26816,N_18339,N_20587);
nor U26817 (N_26817,N_21089,N_21555);
nand U26818 (N_26818,N_23594,N_21483);
and U26819 (N_26819,N_22980,N_21980);
nor U26820 (N_26820,N_21810,N_18638);
and U26821 (N_26821,N_23214,N_22342);
nand U26822 (N_26822,N_22653,N_22837);
or U26823 (N_26823,N_22761,N_21228);
xor U26824 (N_26824,N_19880,N_19140);
or U26825 (N_26825,N_20186,N_23340);
xnor U26826 (N_26826,N_21672,N_21561);
nor U26827 (N_26827,N_21944,N_23960);
nand U26828 (N_26828,N_22690,N_19529);
or U26829 (N_26829,N_18245,N_23429);
and U26830 (N_26830,N_18662,N_20684);
xor U26831 (N_26831,N_18288,N_22062);
or U26832 (N_26832,N_19555,N_21341);
nand U26833 (N_26833,N_19927,N_23080);
and U26834 (N_26834,N_18331,N_23444);
nor U26835 (N_26835,N_23306,N_20693);
or U26836 (N_26836,N_22017,N_18790);
nand U26837 (N_26837,N_23561,N_21602);
nand U26838 (N_26838,N_23753,N_21738);
nand U26839 (N_26839,N_18464,N_19822);
xnor U26840 (N_26840,N_18577,N_18207);
or U26841 (N_26841,N_18754,N_19163);
or U26842 (N_26842,N_23245,N_23914);
and U26843 (N_26843,N_18785,N_20251);
nor U26844 (N_26844,N_22380,N_23387);
and U26845 (N_26845,N_22239,N_22985);
nor U26846 (N_26846,N_22667,N_21546);
or U26847 (N_26847,N_23160,N_19986);
xnor U26848 (N_26848,N_18105,N_23864);
xnor U26849 (N_26849,N_18990,N_22932);
xnor U26850 (N_26850,N_20206,N_20158);
nand U26851 (N_26851,N_21822,N_20763);
xnor U26852 (N_26852,N_23284,N_20047);
or U26853 (N_26853,N_20036,N_20479);
or U26854 (N_26854,N_19439,N_20633);
nor U26855 (N_26855,N_22347,N_20965);
xor U26856 (N_26856,N_22162,N_23477);
and U26857 (N_26857,N_21292,N_18090);
nor U26858 (N_26858,N_18590,N_22926);
xor U26859 (N_26859,N_19607,N_19050);
nand U26860 (N_26860,N_20709,N_20737);
and U26861 (N_26861,N_19997,N_20335);
xnor U26862 (N_26862,N_20691,N_18704);
and U26863 (N_26863,N_22947,N_20589);
and U26864 (N_26864,N_21147,N_20784);
and U26865 (N_26865,N_22344,N_20674);
nor U26866 (N_26866,N_19636,N_20567);
and U26867 (N_26867,N_21661,N_22445);
nand U26868 (N_26868,N_20214,N_18006);
or U26869 (N_26869,N_19709,N_19710);
nand U26870 (N_26870,N_21163,N_23910);
xor U26871 (N_26871,N_21599,N_23543);
nand U26872 (N_26872,N_18215,N_20125);
nand U26873 (N_26873,N_19841,N_18500);
and U26874 (N_26874,N_23421,N_22339);
nor U26875 (N_26875,N_21093,N_20671);
nand U26876 (N_26876,N_19401,N_21114);
xnor U26877 (N_26877,N_18092,N_21200);
nor U26878 (N_26878,N_21133,N_22022);
or U26879 (N_26879,N_18945,N_23495);
nor U26880 (N_26880,N_23935,N_21202);
and U26881 (N_26881,N_18462,N_18667);
nor U26882 (N_26882,N_21452,N_18999);
xor U26883 (N_26883,N_22230,N_18907);
or U26884 (N_26884,N_21505,N_20623);
xnor U26885 (N_26885,N_20661,N_19711);
or U26886 (N_26886,N_20377,N_19966);
xnor U26887 (N_26887,N_23318,N_21805);
or U26888 (N_26888,N_21161,N_23228);
nand U26889 (N_26889,N_22873,N_19758);
xor U26890 (N_26890,N_18826,N_21562);
or U26891 (N_26891,N_22018,N_19313);
nor U26892 (N_26892,N_22729,N_20262);
nor U26893 (N_26893,N_23320,N_22203);
nand U26894 (N_26894,N_19616,N_23337);
nand U26895 (N_26895,N_22231,N_21345);
or U26896 (N_26896,N_23236,N_23865);
and U26897 (N_26897,N_18319,N_21009);
or U26898 (N_26898,N_19360,N_19736);
and U26899 (N_26899,N_22393,N_21817);
nand U26900 (N_26900,N_18053,N_19699);
xor U26901 (N_26901,N_18874,N_22233);
xor U26902 (N_26902,N_18535,N_20082);
nand U26903 (N_26903,N_20389,N_20436);
and U26904 (N_26904,N_18889,N_23118);
xor U26905 (N_26905,N_20811,N_22106);
and U26906 (N_26906,N_20437,N_23022);
or U26907 (N_26907,N_18362,N_20351);
nand U26908 (N_26908,N_20992,N_19074);
or U26909 (N_26909,N_18045,N_23602);
xnor U26910 (N_26910,N_22976,N_23136);
xor U26911 (N_26911,N_20498,N_23525);
or U26912 (N_26912,N_23307,N_23281);
and U26913 (N_26913,N_23278,N_21288);
or U26914 (N_26914,N_23247,N_21334);
nand U26915 (N_26915,N_21724,N_21764);
or U26916 (N_26916,N_22965,N_18338);
nor U26917 (N_26917,N_22905,N_18266);
nand U26918 (N_26918,N_18934,N_19635);
xor U26919 (N_26919,N_23105,N_22208);
xnor U26920 (N_26920,N_21327,N_20938);
nand U26921 (N_26921,N_21978,N_18484);
or U26922 (N_26922,N_23991,N_22627);
nor U26923 (N_26923,N_18336,N_21012);
and U26924 (N_26924,N_19477,N_19621);
and U26925 (N_26925,N_22073,N_23341);
nand U26926 (N_26926,N_22002,N_20268);
nand U26927 (N_26927,N_19893,N_19351);
xor U26928 (N_26928,N_19634,N_22149);
nand U26929 (N_26929,N_18296,N_19537);
nand U26930 (N_26930,N_20664,N_20169);
nor U26931 (N_26931,N_21480,N_18227);
and U26932 (N_26932,N_21418,N_18563);
nor U26933 (N_26933,N_23720,N_19554);
xor U26934 (N_26934,N_18172,N_20049);
xnor U26935 (N_26935,N_21904,N_23995);
and U26936 (N_26936,N_21833,N_22379);
or U26937 (N_26937,N_22631,N_19741);
nand U26938 (N_26938,N_23147,N_19357);
xor U26939 (N_26939,N_21987,N_19772);
and U26940 (N_26940,N_18041,N_19675);
nand U26941 (N_26941,N_18576,N_20491);
and U26942 (N_26942,N_20151,N_21296);
nand U26943 (N_26943,N_21030,N_19825);
or U26944 (N_26944,N_23631,N_18613);
or U26945 (N_26945,N_18374,N_22569);
or U26946 (N_26946,N_22596,N_20821);
and U26947 (N_26947,N_20976,N_21227);
xnor U26948 (N_26948,N_23260,N_23380);
nor U26949 (N_26949,N_20586,N_20897);
nor U26950 (N_26950,N_22088,N_23041);
xnor U26951 (N_26951,N_23930,N_22534);
nand U26952 (N_26952,N_19316,N_23338);
nand U26953 (N_26953,N_19196,N_22466);
and U26954 (N_26954,N_20666,N_19217);
nor U26955 (N_26955,N_20085,N_23945);
or U26956 (N_26956,N_19991,N_18110);
nor U26957 (N_26957,N_21198,N_19389);
nor U26958 (N_26958,N_23971,N_23269);
or U26959 (N_26959,N_22383,N_20886);
nand U26960 (N_26960,N_23416,N_22359);
or U26961 (N_26961,N_19435,N_18902);
nand U26962 (N_26962,N_20930,N_23816);
and U26963 (N_26963,N_20539,N_20482);
xnor U26964 (N_26964,N_22234,N_19648);
or U26965 (N_26965,N_23302,N_23363);
nand U26966 (N_26966,N_23681,N_21211);
or U26967 (N_26967,N_18208,N_19412);
xnor U26968 (N_26968,N_19604,N_22778);
nand U26969 (N_26969,N_18718,N_20275);
nand U26970 (N_26970,N_20398,N_20470);
or U26971 (N_26971,N_18495,N_23977);
and U26972 (N_26972,N_22911,N_19235);
or U26973 (N_26973,N_21164,N_20179);
or U26974 (N_26974,N_20392,N_19935);
nor U26975 (N_26975,N_18040,N_19540);
xor U26976 (N_26976,N_23744,N_23002);
nor U26977 (N_26977,N_20728,N_19919);
xor U26978 (N_26978,N_19030,N_20995);
nor U26979 (N_26979,N_19378,N_18086);
nor U26980 (N_26980,N_18932,N_21866);
and U26981 (N_26981,N_22473,N_19720);
nor U26982 (N_26982,N_22308,N_23131);
xnor U26983 (N_26983,N_20919,N_19458);
nor U26984 (N_26984,N_21821,N_23396);
or U26985 (N_26985,N_19917,N_19454);
nand U26986 (N_26986,N_19137,N_18256);
and U26987 (N_26987,N_22417,N_21329);
nor U26988 (N_26988,N_23618,N_18134);
xor U26989 (N_26989,N_18708,N_20756);
or U26990 (N_26990,N_19845,N_23964);
xor U26991 (N_26991,N_22626,N_21669);
nor U26992 (N_26992,N_18571,N_20148);
or U26993 (N_26993,N_20675,N_18984);
nand U26994 (N_26994,N_18024,N_22660);
and U26995 (N_26995,N_19716,N_22045);
nor U26996 (N_26996,N_18385,N_19948);
nand U26997 (N_26997,N_21444,N_23392);
or U26998 (N_26998,N_21857,N_23624);
nand U26999 (N_26999,N_21991,N_18171);
nor U27000 (N_27000,N_23949,N_22763);
and U27001 (N_27001,N_22766,N_18132);
xor U27002 (N_27002,N_21307,N_21950);
or U27003 (N_27003,N_23647,N_22950);
nand U27004 (N_27004,N_22232,N_18536);
nor U27005 (N_27005,N_20615,N_19375);
nor U27006 (N_27006,N_23305,N_20070);
xnor U27007 (N_27007,N_18126,N_18337);
nand U27008 (N_27008,N_19742,N_22967);
and U27009 (N_27009,N_23723,N_22737);
nor U27010 (N_27010,N_19483,N_19592);
nor U27011 (N_27011,N_23638,N_19843);
xnor U27012 (N_27012,N_23275,N_23592);
or U27013 (N_27013,N_21972,N_22694);
and U27014 (N_27014,N_18977,N_18127);
and U27015 (N_27015,N_18856,N_19820);
nand U27016 (N_27016,N_18219,N_21815);
or U27017 (N_27017,N_21382,N_20621);
nand U27018 (N_27018,N_18771,N_20100);
or U27019 (N_27019,N_21726,N_21914);
nand U27020 (N_27020,N_23150,N_18319);
nand U27021 (N_27021,N_20179,N_19584);
or U27022 (N_27022,N_22412,N_23599);
and U27023 (N_27023,N_18511,N_19250);
xor U27024 (N_27024,N_21187,N_18850);
nor U27025 (N_27025,N_21334,N_20316);
and U27026 (N_27026,N_21981,N_20972);
xnor U27027 (N_27027,N_19088,N_18376);
nor U27028 (N_27028,N_21916,N_20202);
nor U27029 (N_27029,N_19426,N_22100);
or U27030 (N_27030,N_18953,N_23865);
xor U27031 (N_27031,N_20436,N_19700);
xor U27032 (N_27032,N_23512,N_19359);
nor U27033 (N_27033,N_19408,N_23703);
xor U27034 (N_27034,N_19242,N_21354);
nand U27035 (N_27035,N_19430,N_21188);
and U27036 (N_27036,N_22242,N_23787);
nand U27037 (N_27037,N_22028,N_19964);
xnor U27038 (N_27038,N_23152,N_22249);
or U27039 (N_27039,N_18013,N_19064);
nand U27040 (N_27040,N_23915,N_23627);
nand U27041 (N_27041,N_21319,N_18286);
xor U27042 (N_27042,N_20241,N_21041);
nand U27043 (N_27043,N_21257,N_21122);
xnor U27044 (N_27044,N_23389,N_21403);
and U27045 (N_27045,N_21558,N_19563);
or U27046 (N_27046,N_23700,N_18592);
nand U27047 (N_27047,N_19601,N_21871);
xor U27048 (N_27048,N_21176,N_20377);
nor U27049 (N_27049,N_18339,N_22991);
nor U27050 (N_27050,N_22574,N_20390);
and U27051 (N_27051,N_18367,N_19377);
xor U27052 (N_27052,N_22710,N_22940);
nor U27053 (N_27053,N_20908,N_21633);
and U27054 (N_27054,N_23139,N_21373);
nor U27055 (N_27055,N_19603,N_19255);
xnor U27056 (N_27056,N_20220,N_21048);
nor U27057 (N_27057,N_20508,N_20712);
nor U27058 (N_27058,N_20951,N_22012);
or U27059 (N_27059,N_18658,N_18203);
nand U27060 (N_27060,N_18636,N_22501);
nor U27061 (N_27061,N_18239,N_23221);
nand U27062 (N_27062,N_19707,N_22327);
nor U27063 (N_27063,N_22205,N_22779);
or U27064 (N_27064,N_18086,N_22406);
and U27065 (N_27065,N_19423,N_23598);
or U27066 (N_27066,N_23015,N_18665);
nor U27067 (N_27067,N_23381,N_19264);
nand U27068 (N_27068,N_18655,N_22422);
xnor U27069 (N_27069,N_18394,N_19581);
xor U27070 (N_27070,N_19668,N_19506);
and U27071 (N_27071,N_23907,N_21418);
nor U27072 (N_27072,N_22651,N_20525);
xor U27073 (N_27073,N_22160,N_19500);
and U27074 (N_27074,N_20428,N_22561);
nor U27075 (N_27075,N_22070,N_23537);
nor U27076 (N_27076,N_18519,N_21019);
xor U27077 (N_27077,N_18737,N_23151);
xor U27078 (N_27078,N_23807,N_22378);
xnor U27079 (N_27079,N_18458,N_20055);
nor U27080 (N_27080,N_23149,N_21279);
nand U27081 (N_27081,N_21479,N_18072);
nand U27082 (N_27082,N_20641,N_19101);
nor U27083 (N_27083,N_19668,N_23806);
and U27084 (N_27084,N_19113,N_21609);
nand U27085 (N_27085,N_22896,N_22807);
xnor U27086 (N_27086,N_20933,N_22727);
and U27087 (N_27087,N_22810,N_23182);
nand U27088 (N_27088,N_23889,N_18875);
nor U27089 (N_27089,N_18289,N_19237);
nor U27090 (N_27090,N_21554,N_18677);
xnor U27091 (N_27091,N_23835,N_22136);
or U27092 (N_27092,N_23572,N_21805);
and U27093 (N_27093,N_18075,N_21259);
and U27094 (N_27094,N_19075,N_23066);
nand U27095 (N_27095,N_22224,N_21282);
or U27096 (N_27096,N_23731,N_22647);
nor U27097 (N_27097,N_20715,N_20820);
nand U27098 (N_27098,N_22828,N_18440);
and U27099 (N_27099,N_18851,N_20264);
nand U27100 (N_27100,N_21250,N_18658);
nand U27101 (N_27101,N_22640,N_21481);
and U27102 (N_27102,N_22247,N_18739);
nor U27103 (N_27103,N_22882,N_18671);
and U27104 (N_27104,N_23541,N_22598);
or U27105 (N_27105,N_23881,N_21941);
or U27106 (N_27106,N_19327,N_21210);
xnor U27107 (N_27107,N_18633,N_18352);
nand U27108 (N_27108,N_19088,N_18761);
and U27109 (N_27109,N_21772,N_19107);
nor U27110 (N_27110,N_20043,N_21758);
and U27111 (N_27111,N_22909,N_20362);
nor U27112 (N_27112,N_19182,N_20957);
and U27113 (N_27113,N_22834,N_23078);
nand U27114 (N_27114,N_21864,N_19421);
nor U27115 (N_27115,N_21982,N_22750);
and U27116 (N_27116,N_23669,N_19537);
or U27117 (N_27117,N_21918,N_20756);
and U27118 (N_27118,N_22809,N_22075);
nor U27119 (N_27119,N_20401,N_20580);
and U27120 (N_27120,N_18437,N_22298);
nand U27121 (N_27121,N_18103,N_18186);
xor U27122 (N_27122,N_23467,N_18377);
xnor U27123 (N_27123,N_18181,N_21090);
or U27124 (N_27124,N_23175,N_21224);
xnor U27125 (N_27125,N_20495,N_20624);
and U27126 (N_27126,N_22497,N_22024);
nand U27127 (N_27127,N_19278,N_21387);
xor U27128 (N_27128,N_23521,N_23048);
xnor U27129 (N_27129,N_23694,N_21180);
xor U27130 (N_27130,N_21853,N_23665);
nor U27131 (N_27131,N_22490,N_21606);
or U27132 (N_27132,N_18601,N_21969);
nand U27133 (N_27133,N_23470,N_21571);
nand U27134 (N_27134,N_18264,N_22512);
or U27135 (N_27135,N_18630,N_19560);
nor U27136 (N_27136,N_18820,N_23949);
or U27137 (N_27137,N_20960,N_23576);
nand U27138 (N_27138,N_21405,N_22059);
xnor U27139 (N_27139,N_21221,N_21668);
nor U27140 (N_27140,N_18401,N_19545);
or U27141 (N_27141,N_18032,N_23407);
xor U27142 (N_27142,N_19007,N_18284);
and U27143 (N_27143,N_18330,N_19714);
xor U27144 (N_27144,N_21333,N_22766);
nand U27145 (N_27145,N_21236,N_23432);
nand U27146 (N_27146,N_19699,N_18181);
nand U27147 (N_27147,N_21707,N_18777);
nor U27148 (N_27148,N_21042,N_21344);
or U27149 (N_27149,N_20399,N_19235);
and U27150 (N_27150,N_21136,N_22131);
and U27151 (N_27151,N_20275,N_22824);
nand U27152 (N_27152,N_19895,N_18598);
and U27153 (N_27153,N_23807,N_21424);
xnor U27154 (N_27154,N_23811,N_18733);
nor U27155 (N_27155,N_20961,N_21598);
nand U27156 (N_27156,N_18753,N_19638);
nor U27157 (N_27157,N_21641,N_20282);
nand U27158 (N_27158,N_22016,N_23964);
nor U27159 (N_27159,N_19811,N_23715);
and U27160 (N_27160,N_19355,N_23302);
xnor U27161 (N_27161,N_20712,N_21822);
xnor U27162 (N_27162,N_19917,N_19708);
nor U27163 (N_27163,N_22582,N_18043);
and U27164 (N_27164,N_21581,N_19270);
xnor U27165 (N_27165,N_20096,N_20850);
nor U27166 (N_27166,N_19878,N_19670);
nor U27167 (N_27167,N_18565,N_22347);
nand U27168 (N_27168,N_23869,N_21836);
and U27169 (N_27169,N_18227,N_21084);
xor U27170 (N_27170,N_23342,N_20194);
nand U27171 (N_27171,N_18010,N_22245);
nor U27172 (N_27172,N_19974,N_23637);
or U27173 (N_27173,N_21729,N_23442);
and U27174 (N_27174,N_18664,N_19930);
nor U27175 (N_27175,N_21651,N_18048);
nor U27176 (N_27176,N_21634,N_18081);
and U27177 (N_27177,N_19777,N_22160);
and U27178 (N_27178,N_18736,N_23083);
xnor U27179 (N_27179,N_20232,N_23228);
xor U27180 (N_27180,N_22790,N_20572);
or U27181 (N_27181,N_18065,N_19803);
xor U27182 (N_27182,N_21661,N_20383);
xor U27183 (N_27183,N_23729,N_21749);
xnor U27184 (N_27184,N_22341,N_22466);
and U27185 (N_27185,N_20636,N_21297);
nand U27186 (N_27186,N_22080,N_21749);
or U27187 (N_27187,N_21092,N_21005);
nor U27188 (N_27188,N_19861,N_18389);
and U27189 (N_27189,N_22438,N_23655);
or U27190 (N_27190,N_22099,N_22034);
xor U27191 (N_27191,N_19542,N_22074);
nor U27192 (N_27192,N_23518,N_21602);
and U27193 (N_27193,N_20632,N_20239);
or U27194 (N_27194,N_18576,N_19557);
nor U27195 (N_27195,N_21027,N_22757);
nand U27196 (N_27196,N_18748,N_22771);
or U27197 (N_27197,N_19359,N_22109);
nor U27198 (N_27198,N_18100,N_19645);
nand U27199 (N_27199,N_21870,N_22088);
nand U27200 (N_27200,N_20999,N_18550);
or U27201 (N_27201,N_21849,N_21416);
and U27202 (N_27202,N_22942,N_23087);
xor U27203 (N_27203,N_20102,N_20912);
nand U27204 (N_27204,N_22322,N_22044);
or U27205 (N_27205,N_19293,N_21746);
and U27206 (N_27206,N_19074,N_22695);
nor U27207 (N_27207,N_21339,N_18991);
and U27208 (N_27208,N_21945,N_21167);
and U27209 (N_27209,N_18931,N_20034);
or U27210 (N_27210,N_22442,N_22163);
xnor U27211 (N_27211,N_21298,N_22360);
nand U27212 (N_27212,N_21875,N_18317);
or U27213 (N_27213,N_19227,N_19807);
and U27214 (N_27214,N_21239,N_23910);
nand U27215 (N_27215,N_20513,N_18686);
and U27216 (N_27216,N_21496,N_21774);
or U27217 (N_27217,N_19615,N_20201);
nor U27218 (N_27218,N_21759,N_23221);
or U27219 (N_27219,N_21004,N_21978);
xor U27220 (N_27220,N_21109,N_21941);
or U27221 (N_27221,N_18919,N_23568);
xor U27222 (N_27222,N_22117,N_23449);
and U27223 (N_27223,N_20154,N_18443);
nor U27224 (N_27224,N_19376,N_18524);
nor U27225 (N_27225,N_22658,N_20049);
or U27226 (N_27226,N_19280,N_23516);
nor U27227 (N_27227,N_23678,N_22677);
xnor U27228 (N_27228,N_23623,N_20316);
xor U27229 (N_27229,N_20421,N_23980);
or U27230 (N_27230,N_23468,N_21624);
or U27231 (N_27231,N_19085,N_21053);
nor U27232 (N_27232,N_18131,N_20388);
nand U27233 (N_27233,N_19448,N_19848);
or U27234 (N_27234,N_18349,N_20963);
and U27235 (N_27235,N_21799,N_19045);
nand U27236 (N_27236,N_21399,N_20316);
xor U27237 (N_27237,N_23800,N_21340);
xnor U27238 (N_27238,N_23165,N_23953);
nand U27239 (N_27239,N_20834,N_23285);
nand U27240 (N_27240,N_22005,N_19232);
and U27241 (N_27241,N_23479,N_23973);
nor U27242 (N_27242,N_22669,N_18035);
nand U27243 (N_27243,N_19127,N_19326);
nand U27244 (N_27244,N_18310,N_21018);
xnor U27245 (N_27245,N_21152,N_21890);
and U27246 (N_27246,N_18012,N_22387);
xor U27247 (N_27247,N_20572,N_21363);
or U27248 (N_27248,N_18427,N_21563);
and U27249 (N_27249,N_18744,N_18266);
nand U27250 (N_27250,N_23149,N_21778);
nand U27251 (N_27251,N_22268,N_19178);
and U27252 (N_27252,N_23067,N_23009);
nand U27253 (N_27253,N_23810,N_19212);
or U27254 (N_27254,N_20162,N_20435);
xnor U27255 (N_27255,N_20885,N_21504);
and U27256 (N_27256,N_19621,N_22201);
or U27257 (N_27257,N_22218,N_21667);
nor U27258 (N_27258,N_20711,N_20443);
nor U27259 (N_27259,N_19316,N_19150);
nand U27260 (N_27260,N_21918,N_19175);
nand U27261 (N_27261,N_20946,N_22600);
and U27262 (N_27262,N_21287,N_19052);
nand U27263 (N_27263,N_19244,N_18477);
xnor U27264 (N_27264,N_21350,N_20915);
nor U27265 (N_27265,N_18025,N_18768);
or U27266 (N_27266,N_23946,N_22430);
or U27267 (N_27267,N_23910,N_20782);
nand U27268 (N_27268,N_23537,N_23136);
nor U27269 (N_27269,N_19325,N_18076);
xnor U27270 (N_27270,N_22718,N_19118);
and U27271 (N_27271,N_18936,N_20343);
or U27272 (N_27272,N_18872,N_18041);
xor U27273 (N_27273,N_21971,N_20902);
xor U27274 (N_27274,N_22928,N_19349);
nand U27275 (N_27275,N_20819,N_21460);
nand U27276 (N_27276,N_22577,N_19310);
or U27277 (N_27277,N_21753,N_19703);
nand U27278 (N_27278,N_23263,N_19829);
and U27279 (N_27279,N_18371,N_23537);
and U27280 (N_27280,N_21298,N_22752);
and U27281 (N_27281,N_18522,N_20797);
nand U27282 (N_27282,N_18514,N_20140);
nand U27283 (N_27283,N_23635,N_22784);
nor U27284 (N_27284,N_23113,N_23959);
nand U27285 (N_27285,N_23014,N_19885);
nor U27286 (N_27286,N_19449,N_23084);
or U27287 (N_27287,N_18613,N_21379);
or U27288 (N_27288,N_22614,N_18672);
nand U27289 (N_27289,N_22569,N_22554);
or U27290 (N_27290,N_21355,N_23374);
nor U27291 (N_27291,N_21618,N_22692);
nor U27292 (N_27292,N_20774,N_19081);
and U27293 (N_27293,N_18154,N_22602);
xor U27294 (N_27294,N_20866,N_23829);
or U27295 (N_27295,N_23291,N_18254);
and U27296 (N_27296,N_18993,N_21711);
xnor U27297 (N_27297,N_18386,N_21951);
xor U27298 (N_27298,N_23484,N_23413);
nor U27299 (N_27299,N_19548,N_23917);
or U27300 (N_27300,N_19879,N_20001);
and U27301 (N_27301,N_23560,N_21561);
xor U27302 (N_27302,N_20092,N_20992);
nor U27303 (N_27303,N_23181,N_19863);
nand U27304 (N_27304,N_18873,N_21873);
or U27305 (N_27305,N_19105,N_22653);
xor U27306 (N_27306,N_22725,N_19305);
and U27307 (N_27307,N_23438,N_21521);
or U27308 (N_27308,N_23469,N_20519);
nor U27309 (N_27309,N_23373,N_23747);
or U27310 (N_27310,N_21407,N_22065);
xor U27311 (N_27311,N_23381,N_19678);
or U27312 (N_27312,N_21604,N_21923);
xor U27313 (N_27313,N_18873,N_21198);
xor U27314 (N_27314,N_21587,N_23538);
or U27315 (N_27315,N_19737,N_19333);
nor U27316 (N_27316,N_23725,N_23644);
nor U27317 (N_27317,N_23498,N_22080);
nand U27318 (N_27318,N_20812,N_23032);
xor U27319 (N_27319,N_20814,N_20949);
nor U27320 (N_27320,N_18327,N_20433);
nor U27321 (N_27321,N_21595,N_21351);
nand U27322 (N_27322,N_23829,N_21158);
or U27323 (N_27323,N_20454,N_21390);
or U27324 (N_27324,N_18810,N_20093);
nor U27325 (N_27325,N_21761,N_20645);
xor U27326 (N_27326,N_20119,N_22631);
or U27327 (N_27327,N_20399,N_18590);
nand U27328 (N_27328,N_21122,N_22241);
and U27329 (N_27329,N_19661,N_18428);
nor U27330 (N_27330,N_18876,N_21695);
or U27331 (N_27331,N_23355,N_19083);
or U27332 (N_27332,N_22439,N_22708);
or U27333 (N_27333,N_22627,N_23868);
or U27334 (N_27334,N_23556,N_23402);
or U27335 (N_27335,N_23803,N_23323);
nand U27336 (N_27336,N_23458,N_18573);
nor U27337 (N_27337,N_19649,N_19259);
and U27338 (N_27338,N_21489,N_20244);
nor U27339 (N_27339,N_23888,N_18817);
and U27340 (N_27340,N_23827,N_21615);
nand U27341 (N_27341,N_22423,N_22008);
nor U27342 (N_27342,N_20798,N_19955);
or U27343 (N_27343,N_22622,N_21775);
and U27344 (N_27344,N_23917,N_20859);
nand U27345 (N_27345,N_21769,N_22914);
nand U27346 (N_27346,N_22030,N_21333);
or U27347 (N_27347,N_23325,N_18722);
xor U27348 (N_27348,N_22309,N_18076);
xor U27349 (N_27349,N_18807,N_23735);
or U27350 (N_27350,N_22050,N_18952);
nand U27351 (N_27351,N_18992,N_20810);
nor U27352 (N_27352,N_20491,N_22073);
xor U27353 (N_27353,N_18957,N_22297);
nor U27354 (N_27354,N_22144,N_21214);
and U27355 (N_27355,N_18185,N_22964);
nand U27356 (N_27356,N_22798,N_18667);
xnor U27357 (N_27357,N_18814,N_20049);
xor U27358 (N_27358,N_22535,N_22836);
and U27359 (N_27359,N_20631,N_20225);
and U27360 (N_27360,N_22683,N_19932);
or U27361 (N_27361,N_18927,N_19740);
or U27362 (N_27362,N_19786,N_19436);
nand U27363 (N_27363,N_21252,N_20881);
nor U27364 (N_27364,N_19648,N_23891);
and U27365 (N_27365,N_23243,N_18731);
nor U27366 (N_27366,N_23182,N_19641);
nand U27367 (N_27367,N_21577,N_22614);
nand U27368 (N_27368,N_19785,N_22800);
and U27369 (N_27369,N_22474,N_20951);
nor U27370 (N_27370,N_22255,N_22523);
and U27371 (N_27371,N_22048,N_19176);
or U27372 (N_27372,N_23474,N_20862);
and U27373 (N_27373,N_19053,N_23587);
and U27374 (N_27374,N_18303,N_21467);
xnor U27375 (N_27375,N_18247,N_23933);
or U27376 (N_27376,N_23007,N_18224);
or U27377 (N_27377,N_18469,N_23064);
nor U27378 (N_27378,N_20295,N_18533);
nand U27379 (N_27379,N_23381,N_22771);
and U27380 (N_27380,N_19210,N_19455);
and U27381 (N_27381,N_20886,N_18836);
nand U27382 (N_27382,N_22946,N_22745);
or U27383 (N_27383,N_21350,N_22304);
nand U27384 (N_27384,N_23089,N_21673);
nand U27385 (N_27385,N_20584,N_20766);
or U27386 (N_27386,N_22358,N_19145);
nand U27387 (N_27387,N_22014,N_21475);
nor U27388 (N_27388,N_18295,N_21651);
or U27389 (N_27389,N_21241,N_18671);
xor U27390 (N_27390,N_21575,N_21858);
nand U27391 (N_27391,N_20169,N_21840);
or U27392 (N_27392,N_22835,N_19161);
nor U27393 (N_27393,N_22608,N_19569);
or U27394 (N_27394,N_21161,N_19329);
or U27395 (N_27395,N_23586,N_22264);
and U27396 (N_27396,N_22078,N_19984);
nor U27397 (N_27397,N_23188,N_21408);
nor U27398 (N_27398,N_21820,N_20132);
or U27399 (N_27399,N_18651,N_23959);
xor U27400 (N_27400,N_19454,N_20825);
or U27401 (N_27401,N_18446,N_22301);
nor U27402 (N_27402,N_23934,N_19712);
or U27403 (N_27403,N_23474,N_20231);
and U27404 (N_27404,N_23128,N_23431);
nand U27405 (N_27405,N_18233,N_20860);
nand U27406 (N_27406,N_19566,N_20985);
and U27407 (N_27407,N_21009,N_18009);
or U27408 (N_27408,N_21297,N_20195);
xor U27409 (N_27409,N_22726,N_19584);
and U27410 (N_27410,N_22184,N_23850);
xor U27411 (N_27411,N_19273,N_20631);
or U27412 (N_27412,N_20602,N_21702);
xor U27413 (N_27413,N_19558,N_20948);
and U27414 (N_27414,N_18271,N_18633);
or U27415 (N_27415,N_19153,N_20382);
and U27416 (N_27416,N_20543,N_19220);
and U27417 (N_27417,N_19155,N_20023);
nand U27418 (N_27418,N_20391,N_18364);
xor U27419 (N_27419,N_23981,N_21374);
nand U27420 (N_27420,N_19785,N_23577);
and U27421 (N_27421,N_20820,N_21743);
nor U27422 (N_27422,N_19879,N_23742);
and U27423 (N_27423,N_23400,N_22725);
xnor U27424 (N_27424,N_19985,N_19366);
or U27425 (N_27425,N_18049,N_21097);
nor U27426 (N_27426,N_23839,N_21591);
nor U27427 (N_27427,N_21234,N_20255);
nor U27428 (N_27428,N_21500,N_20255);
xor U27429 (N_27429,N_22844,N_21071);
and U27430 (N_27430,N_23852,N_21063);
or U27431 (N_27431,N_19232,N_20095);
xnor U27432 (N_27432,N_21089,N_20356);
nand U27433 (N_27433,N_18890,N_19840);
xnor U27434 (N_27434,N_23647,N_20819);
and U27435 (N_27435,N_19513,N_20640);
xor U27436 (N_27436,N_21766,N_22188);
nor U27437 (N_27437,N_22412,N_19173);
xnor U27438 (N_27438,N_21883,N_19350);
or U27439 (N_27439,N_23088,N_22707);
nand U27440 (N_27440,N_19203,N_23636);
or U27441 (N_27441,N_22789,N_19617);
nor U27442 (N_27442,N_19785,N_23551);
nand U27443 (N_27443,N_18222,N_20059);
xor U27444 (N_27444,N_18335,N_23197);
or U27445 (N_27445,N_18971,N_18360);
nand U27446 (N_27446,N_23011,N_23143);
nand U27447 (N_27447,N_20331,N_18828);
nand U27448 (N_27448,N_23136,N_20439);
xnor U27449 (N_27449,N_20880,N_21118);
nand U27450 (N_27450,N_19624,N_21538);
xor U27451 (N_27451,N_22391,N_19389);
or U27452 (N_27452,N_18787,N_21608);
and U27453 (N_27453,N_19269,N_20792);
or U27454 (N_27454,N_22235,N_22079);
nor U27455 (N_27455,N_22720,N_19564);
nand U27456 (N_27456,N_18649,N_21016);
nand U27457 (N_27457,N_19426,N_21057);
xor U27458 (N_27458,N_22113,N_22892);
or U27459 (N_27459,N_23284,N_23480);
nand U27460 (N_27460,N_21055,N_22518);
nor U27461 (N_27461,N_19051,N_20936);
nor U27462 (N_27462,N_23641,N_19543);
nor U27463 (N_27463,N_19217,N_19022);
nand U27464 (N_27464,N_22915,N_18982);
or U27465 (N_27465,N_21879,N_21689);
and U27466 (N_27466,N_19629,N_22483);
and U27467 (N_27467,N_21471,N_18502);
or U27468 (N_27468,N_18222,N_22104);
nor U27469 (N_27469,N_22319,N_18691);
nand U27470 (N_27470,N_22578,N_19727);
xnor U27471 (N_27471,N_21105,N_23066);
or U27472 (N_27472,N_18360,N_22855);
nor U27473 (N_27473,N_19945,N_23133);
nor U27474 (N_27474,N_21258,N_19152);
or U27475 (N_27475,N_18232,N_19454);
xor U27476 (N_27476,N_20001,N_18840);
nand U27477 (N_27477,N_23836,N_21648);
or U27478 (N_27478,N_23769,N_19393);
nor U27479 (N_27479,N_19256,N_19700);
xor U27480 (N_27480,N_21854,N_21348);
nor U27481 (N_27481,N_21127,N_21589);
and U27482 (N_27482,N_23570,N_20982);
and U27483 (N_27483,N_19786,N_19409);
and U27484 (N_27484,N_23283,N_23863);
nand U27485 (N_27485,N_23390,N_19050);
xnor U27486 (N_27486,N_23138,N_21081);
and U27487 (N_27487,N_22229,N_18727);
nor U27488 (N_27488,N_20731,N_18619);
xnor U27489 (N_27489,N_23385,N_20181);
or U27490 (N_27490,N_21059,N_20808);
and U27491 (N_27491,N_22871,N_18034);
nor U27492 (N_27492,N_21273,N_19377);
nor U27493 (N_27493,N_22996,N_23631);
nand U27494 (N_27494,N_20467,N_20129);
and U27495 (N_27495,N_18966,N_23524);
or U27496 (N_27496,N_18701,N_22711);
nor U27497 (N_27497,N_21077,N_22818);
xor U27498 (N_27498,N_19155,N_23788);
or U27499 (N_27499,N_19612,N_20728);
nor U27500 (N_27500,N_20138,N_20631);
xnor U27501 (N_27501,N_23305,N_20398);
nand U27502 (N_27502,N_19917,N_22659);
xnor U27503 (N_27503,N_23911,N_20420);
or U27504 (N_27504,N_18230,N_23767);
and U27505 (N_27505,N_18709,N_21738);
or U27506 (N_27506,N_19280,N_20430);
xor U27507 (N_27507,N_18340,N_20254);
and U27508 (N_27508,N_19527,N_20662);
and U27509 (N_27509,N_21968,N_22701);
xnor U27510 (N_27510,N_23677,N_18342);
xor U27511 (N_27511,N_20569,N_23544);
and U27512 (N_27512,N_20111,N_20554);
xor U27513 (N_27513,N_23035,N_19266);
nor U27514 (N_27514,N_22096,N_21108);
and U27515 (N_27515,N_23198,N_23697);
nand U27516 (N_27516,N_22200,N_21243);
nand U27517 (N_27517,N_23156,N_23786);
and U27518 (N_27518,N_20857,N_20391);
nor U27519 (N_27519,N_21319,N_22836);
nor U27520 (N_27520,N_18753,N_20816);
and U27521 (N_27521,N_20056,N_18683);
or U27522 (N_27522,N_19750,N_19214);
nor U27523 (N_27523,N_23017,N_21603);
and U27524 (N_27524,N_21913,N_19682);
or U27525 (N_27525,N_18545,N_23157);
xor U27526 (N_27526,N_18953,N_22279);
nor U27527 (N_27527,N_18843,N_18929);
or U27528 (N_27528,N_21006,N_23671);
xnor U27529 (N_27529,N_23179,N_23306);
or U27530 (N_27530,N_22855,N_21136);
nor U27531 (N_27531,N_18997,N_18003);
nand U27532 (N_27532,N_18695,N_20551);
nand U27533 (N_27533,N_19688,N_18055);
or U27534 (N_27534,N_20144,N_23568);
nand U27535 (N_27535,N_19875,N_23521);
or U27536 (N_27536,N_20683,N_23947);
or U27537 (N_27537,N_20371,N_18623);
nand U27538 (N_27538,N_18373,N_23867);
xor U27539 (N_27539,N_20713,N_21588);
xor U27540 (N_27540,N_23219,N_18671);
xor U27541 (N_27541,N_21399,N_18945);
or U27542 (N_27542,N_20598,N_21075);
nand U27543 (N_27543,N_23769,N_19751);
nor U27544 (N_27544,N_23378,N_21321);
or U27545 (N_27545,N_23255,N_18705);
nor U27546 (N_27546,N_19049,N_21057);
or U27547 (N_27547,N_18688,N_21409);
or U27548 (N_27548,N_20365,N_19647);
and U27549 (N_27549,N_18859,N_20414);
nand U27550 (N_27550,N_18387,N_21012);
nor U27551 (N_27551,N_23148,N_22366);
xor U27552 (N_27552,N_21259,N_19779);
and U27553 (N_27553,N_21843,N_20658);
nor U27554 (N_27554,N_23103,N_21424);
or U27555 (N_27555,N_19563,N_21018);
xor U27556 (N_27556,N_22159,N_19789);
and U27557 (N_27557,N_23572,N_21243);
xor U27558 (N_27558,N_20795,N_21453);
xor U27559 (N_27559,N_20017,N_21732);
or U27560 (N_27560,N_20323,N_22250);
nand U27561 (N_27561,N_19973,N_21684);
nor U27562 (N_27562,N_20124,N_22030);
nand U27563 (N_27563,N_19222,N_18805);
and U27564 (N_27564,N_23702,N_21800);
and U27565 (N_27565,N_20934,N_23921);
and U27566 (N_27566,N_20244,N_22737);
nor U27567 (N_27567,N_20011,N_18157);
xor U27568 (N_27568,N_18314,N_22766);
and U27569 (N_27569,N_21195,N_22651);
nand U27570 (N_27570,N_22440,N_21485);
xnor U27571 (N_27571,N_20311,N_23262);
xnor U27572 (N_27572,N_18734,N_23249);
nor U27573 (N_27573,N_18050,N_20844);
and U27574 (N_27574,N_20020,N_21591);
and U27575 (N_27575,N_18096,N_23262);
nor U27576 (N_27576,N_20420,N_22956);
nand U27577 (N_27577,N_23848,N_23790);
nor U27578 (N_27578,N_22278,N_19932);
and U27579 (N_27579,N_19561,N_19982);
and U27580 (N_27580,N_20221,N_20739);
and U27581 (N_27581,N_18871,N_22729);
nand U27582 (N_27582,N_23006,N_18923);
nor U27583 (N_27583,N_20588,N_23940);
or U27584 (N_27584,N_23442,N_20478);
nand U27585 (N_27585,N_19927,N_18146);
or U27586 (N_27586,N_22933,N_18766);
nand U27587 (N_27587,N_23945,N_22009);
or U27588 (N_27588,N_23394,N_20761);
nand U27589 (N_27589,N_20249,N_21363);
or U27590 (N_27590,N_23576,N_18072);
xnor U27591 (N_27591,N_19545,N_23612);
and U27592 (N_27592,N_18959,N_20304);
and U27593 (N_27593,N_20895,N_22991);
or U27594 (N_27594,N_21765,N_22124);
nand U27595 (N_27595,N_23732,N_19752);
or U27596 (N_27596,N_20762,N_21452);
and U27597 (N_27597,N_23552,N_19205);
and U27598 (N_27598,N_23795,N_23405);
or U27599 (N_27599,N_19553,N_19276);
nand U27600 (N_27600,N_20824,N_19256);
xnor U27601 (N_27601,N_18005,N_22761);
nor U27602 (N_27602,N_20811,N_20766);
and U27603 (N_27603,N_21531,N_20118);
or U27604 (N_27604,N_21871,N_18632);
nor U27605 (N_27605,N_19139,N_20332);
or U27606 (N_27606,N_20999,N_21899);
nand U27607 (N_27607,N_21948,N_20870);
or U27608 (N_27608,N_22316,N_23342);
nor U27609 (N_27609,N_18730,N_22875);
and U27610 (N_27610,N_23243,N_18392);
or U27611 (N_27611,N_23833,N_20944);
or U27612 (N_27612,N_18231,N_19666);
xnor U27613 (N_27613,N_23666,N_18524);
and U27614 (N_27614,N_21252,N_22944);
and U27615 (N_27615,N_19791,N_22892);
and U27616 (N_27616,N_18674,N_22300);
nand U27617 (N_27617,N_21905,N_18754);
or U27618 (N_27618,N_20335,N_20294);
nor U27619 (N_27619,N_18808,N_23753);
nor U27620 (N_27620,N_22177,N_18878);
xnor U27621 (N_27621,N_23641,N_20899);
and U27622 (N_27622,N_22326,N_18152);
and U27623 (N_27623,N_19493,N_19309);
nor U27624 (N_27624,N_18907,N_19411);
nor U27625 (N_27625,N_22695,N_20996);
and U27626 (N_27626,N_23886,N_21127);
nor U27627 (N_27627,N_21174,N_18123);
and U27628 (N_27628,N_18520,N_23056);
and U27629 (N_27629,N_21071,N_19786);
nor U27630 (N_27630,N_19061,N_20333);
and U27631 (N_27631,N_19179,N_18219);
and U27632 (N_27632,N_22590,N_23277);
or U27633 (N_27633,N_19995,N_21074);
or U27634 (N_27634,N_20434,N_18497);
xor U27635 (N_27635,N_21869,N_18580);
nor U27636 (N_27636,N_21252,N_23271);
nand U27637 (N_27637,N_19388,N_20883);
nor U27638 (N_27638,N_22126,N_19611);
or U27639 (N_27639,N_18709,N_21326);
xnor U27640 (N_27640,N_18882,N_20779);
nor U27641 (N_27641,N_21422,N_22558);
or U27642 (N_27642,N_23293,N_21433);
nand U27643 (N_27643,N_19348,N_22844);
nor U27644 (N_27644,N_19611,N_18421);
xor U27645 (N_27645,N_18537,N_23836);
and U27646 (N_27646,N_18191,N_22181);
xor U27647 (N_27647,N_22950,N_21510);
and U27648 (N_27648,N_18995,N_18588);
xor U27649 (N_27649,N_19800,N_22469);
nand U27650 (N_27650,N_19249,N_22881);
nand U27651 (N_27651,N_20543,N_20744);
nand U27652 (N_27652,N_21464,N_21028);
or U27653 (N_27653,N_21726,N_23926);
xor U27654 (N_27654,N_18095,N_19556);
nand U27655 (N_27655,N_21581,N_22229);
or U27656 (N_27656,N_21988,N_21184);
or U27657 (N_27657,N_22300,N_18334);
nand U27658 (N_27658,N_21192,N_18620);
nor U27659 (N_27659,N_18424,N_19712);
and U27660 (N_27660,N_20961,N_22761);
or U27661 (N_27661,N_22266,N_21695);
or U27662 (N_27662,N_22312,N_22681);
nand U27663 (N_27663,N_20125,N_23549);
nand U27664 (N_27664,N_21019,N_18832);
and U27665 (N_27665,N_22901,N_21804);
or U27666 (N_27666,N_20622,N_19264);
nor U27667 (N_27667,N_22825,N_20511);
nand U27668 (N_27668,N_22804,N_23621);
nand U27669 (N_27669,N_23981,N_21946);
xor U27670 (N_27670,N_21761,N_21272);
xor U27671 (N_27671,N_19724,N_21086);
nor U27672 (N_27672,N_18910,N_21297);
nand U27673 (N_27673,N_20616,N_22975);
nor U27674 (N_27674,N_18524,N_20883);
xnor U27675 (N_27675,N_21153,N_21468);
xor U27676 (N_27676,N_18454,N_19952);
and U27677 (N_27677,N_19619,N_22303);
xnor U27678 (N_27678,N_20831,N_19734);
or U27679 (N_27679,N_21616,N_21883);
xnor U27680 (N_27680,N_18461,N_18093);
nor U27681 (N_27681,N_18091,N_23414);
xor U27682 (N_27682,N_23432,N_18320);
or U27683 (N_27683,N_23326,N_19046);
or U27684 (N_27684,N_22321,N_23754);
xnor U27685 (N_27685,N_21744,N_20427);
nor U27686 (N_27686,N_22901,N_22795);
nand U27687 (N_27687,N_18052,N_19722);
xnor U27688 (N_27688,N_23932,N_21187);
and U27689 (N_27689,N_21968,N_18793);
nor U27690 (N_27690,N_23950,N_18460);
or U27691 (N_27691,N_20039,N_19991);
and U27692 (N_27692,N_20076,N_23189);
nor U27693 (N_27693,N_19243,N_23520);
nand U27694 (N_27694,N_19794,N_23042);
xor U27695 (N_27695,N_19930,N_21160);
or U27696 (N_27696,N_23853,N_23700);
and U27697 (N_27697,N_22174,N_23387);
nor U27698 (N_27698,N_22017,N_22802);
and U27699 (N_27699,N_18503,N_22115);
or U27700 (N_27700,N_21632,N_19734);
xnor U27701 (N_27701,N_19570,N_23719);
or U27702 (N_27702,N_22604,N_19414);
and U27703 (N_27703,N_19533,N_19029);
nor U27704 (N_27704,N_18911,N_21524);
or U27705 (N_27705,N_19071,N_18989);
nor U27706 (N_27706,N_22385,N_18085);
nand U27707 (N_27707,N_23775,N_20532);
nor U27708 (N_27708,N_20399,N_20608);
nand U27709 (N_27709,N_18308,N_19025);
xor U27710 (N_27710,N_23843,N_22970);
nor U27711 (N_27711,N_23115,N_18190);
nand U27712 (N_27712,N_21187,N_22733);
nor U27713 (N_27713,N_21956,N_18525);
or U27714 (N_27714,N_23098,N_23935);
and U27715 (N_27715,N_22374,N_18648);
and U27716 (N_27716,N_22273,N_23060);
xor U27717 (N_27717,N_18945,N_18487);
xor U27718 (N_27718,N_21520,N_22315);
xnor U27719 (N_27719,N_22693,N_23048);
xnor U27720 (N_27720,N_18650,N_21156);
and U27721 (N_27721,N_21120,N_20346);
and U27722 (N_27722,N_20631,N_19987);
nor U27723 (N_27723,N_23055,N_22241);
xor U27724 (N_27724,N_19644,N_20002);
nor U27725 (N_27725,N_19002,N_18166);
nand U27726 (N_27726,N_19997,N_18621);
nor U27727 (N_27727,N_23804,N_20955);
nand U27728 (N_27728,N_22080,N_22134);
nand U27729 (N_27729,N_19419,N_21433);
nor U27730 (N_27730,N_19224,N_21465);
and U27731 (N_27731,N_20888,N_19509);
nor U27732 (N_27732,N_23071,N_19353);
xnor U27733 (N_27733,N_21952,N_20034);
and U27734 (N_27734,N_19424,N_19707);
and U27735 (N_27735,N_19114,N_22297);
nor U27736 (N_27736,N_21417,N_23548);
nand U27737 (N_27737,N_18190,N_20563);
or U27738 (N_27738,N_22893,N_20448);
xnor U27739 (N_27739,N_21984,N_22388);
nand U27740 (N_27740,N_22605,N_22165);
or U27741 (N_27741,N_23483,N_23628);
xnor U27742 (N_27742,N_23737,N_22921);
or U27743 (N_27743,N_22407,N_19697);
and U27744 (N_27744,N_20814,N_21594);
and U27745 (N_27745,N_20496,N_23826);
nand U27746 (N_27746,N_23534,N_23920);
xnor U27747 (N_27747,N_22340,N_21791);
nor U27748 (N_27748,N_22692,N_23884);
nor U27749 (N_27749,N_20760,N_19848);
or U27750 (N_27750,N_19221,N_22850);
and U27751 (N_27751,N_19489,N_23239);
nor U27752 (N_27752,N_20521,N_21447);
xnor U27753 (N_27753,N_22159,N_19301);
nor U27754 (N_27754,N_23683,N_20374);
xor U27755 (N_27755,N_21811,N_19052);
xnor U27756 (N_27756,N_23505,N_21673);
xor U27757 (N_27757,N_18457,N_20042);
nand U27758 (N_27758,N_18980,N_19089);
and U27759 (N_27759,N_20707,N_21806);
or U27760 (N_27760,N_23856,N_20228);
and U27761 (N_27761,N_21141,N_20949);
xor U27762 (N_27762,N_23172,N_23498);
and U27763 (N_27763,N_19111,N_22079);
nand U27764 (N_27764,N_21530,N_20067);
or U27765 (N_27765,N_18268,N_21093);
nor U27766 (N_27766,N_19356,N_21025);
nand U27767 (N_27767,N_23683,N_21316);
or U27768 (N_27768,N_20049,N_18720);
nor U27769 (N_27769,N_19223,N_23831);
and U27770 (N_27770,N_20871,N_22719);
and U27771 (N_27771,N_18725,N_23492);
xor U27772 (N_27772,N_23126,N_19085);
xnor U27773 (N_27773,N_21366,N_21602);
nand U27774 (N_27774,N_19267,N_21590);
or U27775 (N_27775,N_23557,N_23165);
xor U27776 (N_27776,N_19109,N_18342);
xor U27777 (N_27777,N_23209,N_23991);
or U27778 (N_27778,N_23552,N_20246);
nand U27779 (N_27779,N_19885,N_22564);
nand U27780 (N_27780,N_23231,N_23330);
nand U27781 (N_27781,N_22900,N_22790);
nand U27782 (N_27782,N_20745,N_20835);
xnor U27783 (N_27783,N_19735,N_19379);
and U27784 (N_27784,N_23783,N_23075);
or U27785 (N_27785,N_22095,N_23440);
and U27786 (N_27786,N_23392,N_22246);
xor U27787 (N_27787,N_18244,N_22237);
or U27788 (N_27788,N_23899,N_23642);
nor U27789 (N_27789,N_21610,N_23146);
or U27790 (N_27790,N_19265,N_20445);
nand U27791 (N_27791,N_22761,N_21630);
nand U27792 (N_27792,N_18788,N_21372);
and U27793 (N_27793,N_20554,N_18285);
and U27794 (N_27794,N_19343,N_18475);
xor U27795 (N_27795,N_22145,N_23883);
nor U27796 (N_27796,N_23808,N_22129);
nor U27797 (N_27797,N_21442,N_18362);
and U27798 (N_27798,N_19541,N_20288);
and U27799 (N_27799,N_18178,N_19023);
and U27800 (N_27800,N_18546,N_18099);
or U27801 (N_27801,N_23630,N_19137);
nand U27802 (N_27802,N_18720,N_20005);
xor U27803 (N_27803,N_20286,N_20302);
xor U27804 (N_27804,N_20485,N_22216);
xor U27805 (N_27805,N_18682,N_20464);
nand U27806 (N_27806,N_19022,N_22852);
nand U27807 (N_27807,N_23066,N_21184);
and U27808 (N_27808,N_21256,N_22754);
xor U27809 (N_27809,N_18500,N_20041);
and U27810 (N_27810,N_18201,N_23160);
or U27811 (N_27811,N_20214,N_20557);
nor U27812 (N_27812,N_19794,N_22370);
and U27813 (N_27813,N_20750,N_18894);
and U27814 (N_27814,N_19375,N_20711);
xnor U27815 (N_27815,N_18758,N_19621);
xnor U27816 (N_27816,N_20393,N_18192);
and U27817 (N_27817,N_20765,N_20488);
or U27818 (N_27818,N_18055,N_21463);
xnor U27819 (N_27819,N_23236,N_21531);
or U27820 (N_27820,N_19491,N_22722);
or U27821 (N_27821,N_23718,N_23788);
and U27822 (N_27822,N_19946,N_20678);
and U27823 (N_27823,N_18100,N_19429);
or U27824 (N_27824,N_21806,N_18885);
xnor U27825 (N_27825,N_21230,N_18222);
and U27826 (N_27826,N_22661,N_19394);
and U27827 (N_27827,N_23304,N_20472);
xor U27828 (N_27828,N_19286,N_22141);
nor U27829 (N_27829,N_23900,N_20217);
nor U27830 (N_27830,N_23404,N_20745);
xnor U27831 (N_27831,N_21498,N_21247);
xnor U27832 (N_27832,N_20259,N_23152);
nor U27833 (N_27833,N_23270,N_23482);
or U27834 (N_27834,N_20647,N_19685);
nand U27835 (N_27835,N_23724,N_21807);
nor U27836 (N_27836,N_23235,N_22247);
or U27837 (N_27837,N_21014,N_23534);
and U27838 (N_27838,N_23102,N_18929);
xor U27839 (N_27839,N_20820,N_19825);
or U27840 (N_27840,N_22919,N_19104);
xor U27841 (N_27841,N_19586,N_21498);
xnor U27842 (N_27842,N_19243,N_20031);
xnor U27843 (N_27843,N_19107,N_18415);
nor U27844 (N_27844,N_23840,N_23049);
and U27845 (N_27845,N_18719,N_22046);
xor U27846 (N_27846,N_18100,N_23301);
nor U27847 (N_27847,N_19711,N_19984);
nor U27848 (N_27848,N_18807,N_23544);
or U27849 (N_27849,N_22328,N_21256);
xor U27850 (N_27850,N_20936,N_20229);
or U27851 (N_27851,N_20457,N_20733);
and U27852 (N_27852,N_22936,N_22885);
nor U27853 (N_27853,N_22245,N_21760);
xnor U27854 (N_27854,N_21036,N_19363);
and U27855 (N_27855,N_19042,N_20805);
and U27856 (N_27856,N_19203,N_23853);
nor U27857 (N_27857,N_22723,N_18476);
or U27858 (N_27858,N_19458,N_23383);
xor U27859 (N_27859,N_23245,N_23827);
and U27860 (N_27860,N_23409,N_22709);
nor U27861 (N_27861,N_22850,N_18248);
xnor U27862 (N_27862,N_18676,N_22221);
xor U27863 (N_27863,N_20712,N_21924);
nor U27864 (N_27864,N_20471,N_22812);
or U27865 (N_27865,N_19121,N_20690);
and U27866 (N_27866,N_19977,N_18287);
or U27867 (N_27867,N_21963,N_19997);
nor U27868 (N_27868,N_18510,N_19996);
nor U27869 (N_27869,N_22930,N_22256);
xnor U27870 (N_27870,N_18298,N_19290);
nand U27871 (N_27871,N_18076,N_19392);
nor U27872 (N_27872,N_18673,N_19999);
xnor U27873 (N_27873,N_22895,N_20696);
nor U27874 (N_27874,N_22400,N_18231);
or U27875 (N_27875,N_21561,N_18031);
nand U27876 (N_27876,N_23018,N_22908);
and U27877 (N_27877,N_23548,N_20658);
and U27878 (N_27878,N_22172,N_18909);
xnor U27879 (N_27879,N_18632,N_23603);
nand U27880 (N_27880,N_22883,N_23983);
and U27881 (N_27881,N_18556,N_20936);
nand U27882 (N_27882,N_21239,N_21472);
and U27883 (N_27883,N_21190,N_22575);
nor U27884 (N_27884,N_19755,N_23382);
nor U27885 (N_27885,N_18515,N_22600);
xnor U27886 (N_27886,N_18500,N_19705);
xnor U27887 (N_27887,N_23953,N_18531);
xor U27888 (N_27888,N_18735,N_22034);
or U27889 (N_27889,N_18234,N_21098);
nor U27890 (N_27890,N_23609,N_19489);
nand U27891 (N_27891,N_20278,N_18016);
or U27892 (N_27892,N_18927,N_19721);
nand U27893 (N_27893,N_23290,N_22893);
nand U27894 (N_27894,N_18831,N_23666);
or U27895 (N_27895,N_21742,N_21933);
nor U27896 (N_27896,N_19336,N_19108);
xnor U27897 (N_27897,N_23772,N_19248);
xnor U27898 (N_27898,N_19045,N_23056);
xor U27899 (N_27899,N_23699,N_21749);
xor U27900 (N_27900,N_18413,N_20985);
and U27901 (N_27901,N_18487,N_20100);
nor U27902 (N_27902,N_20750,N_23415);
nor U27903 (N_27903,N_19311,N_22597);
or U27904 (N_27904,N_21709,N_21992);
or U27905 (N_27905,N_19958,N_18293);
xor U27906 (N_27906,N_23495,N_18468);
nand U27907 (N_27907,N_20085,N_21603);
nand U27908 (N_27908,N_20370,N_20034);
or U27909 (N_27909,N_21368,N_18996);
nand U27910 (N_27910,N_20861,N_21156);
nor U27911 (N_27911,N_19799,N_19747);
or U27912 (N_27912,N_19395,N_21983);
nor U27913 (N_27913,N_21279,N_21534);
nand U27914 (N_27914,N_21180,N_18048);
and U27915 (N_27915,N_20826,N_23244);
or U27916 (N_27916,N_21618,N_18576);
or U27917 (N_27917,N_19112,N_22521);
and U27918 (N_27918,N_18486,N_19171);
xnor U27919 (N_27919,N_20424,N_22702);
or U27920 (N_27920,N_19181,N_23841);
nor U27921 (N_27921,N_19352,N_18877);
xnor U27922 (N_27922,N_20332,N_20746);
or U27923 (N_27923,N_21108,N_22917);
nand U27924 (N_27924,N_23668,N_23712);
xor U27925 (N_27925,N_18653,N_20926);
and U27926 (N_27926,N_20941,N_21563);
or U27927 (N_27927,N_21991,N_18609);
xnor U27928 (N_27928,N_22988,N_18085);
or U27929 (N_27929,N_20463,N_18452);
nand U27930 (N_27930,N_23052,N_22500);
nand U27931 (N_27931,N_18170,N_20396);
nand U27932 (N_27932,N_19782,N_23978);
and U27933 (N_27933,N_20052,N_23934);
and U27934 (N_27934,N_19921,N_18688);
nor U27935 (N_27935,N_21714,N_23990);
and U27936 (N_27936,N_23953,N_23067);
or U27937 (N_27937,N_19067,N_20145);
and U27938 (N_27938,N_22538,N_21954);
xnor U27939 (N_27939,N_20544,N_20869);
nor U27940 (N_27940,N_19349,N_22189);
nand U27941 (N_27941,N_20925,N_22365);
nor U27942 (N_27942,N_21282,N_18901);
and U27943 (N_27943,N_18889,N_20654);
and U27944 (N_27944,N_21072,N_20339);
xor U27945 (N_27945,N_21865,N_21087);
xor U27946 (N_27946,N_19104,N_20540);
xor U27947 (N_27947,N_19034,N_18237);
nand U27948 (N_27948,N_22877,N_23693);
nor U27949 (N_27949,N_18519,N_19287);
nor U27950 (N_27950,N_23827,N_20821);
nand U27951 (N_27951,N_18087,N_23619);
xor U27952 (N_27952,N_19838,N_20820);
nor U27953 (N_27953,N_19740,N_23071);
xor U27954 (N_27954,N_21504,N_19419);
or U27955 (N_27955,N_18224,N_19062);
nand U27956 (N_27956,N_18770,N_20376);
xnor U27957 (N_27957,N_21617,N_21638);
or U27958 (N_27958,N_21351,N_23312);
and U27959 (N_27959,N_18563,N_21863);
xor U27960 (N_27960,N_23688,N_18834);
nand U27961 (N_27961,N_20089,N_18690);
or U27962 (N_27962,N_22338,N_18311);
nor U27963 (N_27963,N_19253,N_20322);
nand U27964 (N_27964,N_22307,N_22302);
nand U27965 (N_27965,N_18026,N_18777);
or U27966 (N_27966,N_19026,N_19444);
and U27967 (N_27967,N_18356,N_22379);
nand U27968 (N_27968,N_21727,N_19637);
nor U27969 (N_27969,N_21843,N_20759);
and U27970 (N_27970,N_18863,N_22162);
and U27971 (N_27971,N_22852,N_21680);
nor U27972 (N_27972,N_22575,N_19758);
and U27973 (N_27973,N_18192,N_21474);
or U27974 (N_27974,N_23185,N_23724);
nor U27975 (N_27975,N_23223,N_18238);
xor U27976 (N_27976,N_18446,N_22123);
xor U27977 (N_27977,N_21596,N_18616);
or U27978 (N_27978,N_21781,N_19086);
and U27979 (N_27979,N_21081,N_21781);
nand U27980 (N_27980,N_22556,N_21543);
nor U27981 (N_27981,N_21567,N_22669);
and U27982 (N_27982,N_19854,N_22794);
nor U27983 (N_27983,N_21573,N_22428);
xnor U27984 (N_27984,N_19434,N_18352);
nor U27985 (N_27985,N_18828,N_19851);
nor U27986 (N_27986,N_22861,N_20459);
and U27987 (N_27987,N_23407,N_19785);
and U27988 (N_27988,N_21852,N_19999);
or U27989 (N_27989,N_19311,N_18100);
nor U27990 (N_27990,N_20019,N_22027);
nand U27991 (N_27991,N_23075,N_18934);
and U27992 (N_27992,N_18676,N_20630);
and U27993 (N_27993,N_18077,N_21185);
or U27994 (N_27994,N_19869,N_22857);
nor U27995 (N_27995,N_19662,N_23608);
and U27996 (N_27996,N_21270,N_20821);
nor U27997 (N_27997,N_23420,N_20343);
or U27998 (N_27998,N_22898,N_23476);
xor U27999 (N_27999,N_22129,N_21301);
xor U28000 (N_28000,N_19431,N_22503);
xor U28001 (N_28001,N_18813,N_22859);
or U28002 (N_28002,N_19179,N_21649);
and U28003 (N_28003,N_18972,N_21469);
nand U28004 (N_28004,N_21328,N_18792);
or U28005 (N_28005,N_21173,N_23765);
nor U28006 (N_28006,N_20320,N_23907);
nand U28007 (N_28007,N_20844,N_19199);
or U28008 (N_28008,N_22681,N_23740);
or U28009 (N_28009,N_19237,N_19190);
nand U28010 (N_28010,N_23668,N_18035);
or U28011 (N_28011,N_23206,N_20640);
or U28012 (N_28012,N_18949,N_21174);
and U28013 (N_28013,N_21526,N_21245);
or U28014 (N_28014,N_23658,N_22240);
nand U28015 (N_28015,N_19556,N_23835);
or U28016 (N_28016,N_22218,N_23214);
and U28017 (N_28017,N_18790,N_21434);
and U28018 (N_28018,N_18478,N_21039);
nand U28019 (N_28019,N_18883,N_18927);
and U28020 (N_28020,N_23340,N_19367);
nand U28021 (N_28021,N_22304,N_21709);
nand U28022 (N_28022,N_22248,N_19757);
xor U28023 (N_28023,N_23299,N_23265);
nand U28024 (N_28024,N_23613,N_19736);
and U28025 (N_28025,N_23593,N_20491);
nand U28026 (N_28026,N_23145,N_20539);
nor U28027 (N_28027,N_23165,N_19786);
nand U28028 (N_28028,N_23808,N_23427);
or U28029 (N_28029,N_18526,N_23595);
and U28030 (N_28030,N_22271,N_19647);
xor U28031 (N_28031,N_21411,N_23627);
or U28032 (N_28032,N_20380,N_18551);
or U28033 (N_28033,N_18299,N_20685);
nand U28034 (N_28034,N_19269,N_19597);
xor U28035 (N_28035,N_23933,N_20801);
nand U28036 (N_28036,N_22243,N_20334);
nor U28037 (N_28037,N_21859,N_20982);
or U28038 (N_28038,N_19436,N_23610);
and U28039 (N_28039,N_20020,N_19211);
or U28040 (N_28040,N_20007,N_19200);
nor U28041 (N_28041,N_21415,N_22013);
or U28042 (N_28042,N_19329,N_19141);
nor U28043 (N_28043,N_18750,N_20384);
xor U28044 (N_28044,N_23528,N_21178);
nand U28045 (N_28045,N_19143,N_21646);
nor U28046 (N_28046,N_19346,N_19214);
xnor U28047 (N_28047,N_23239,N_23592);
and U28048 (N_28048,N_20746,N_19707);
or U28049 (N_28049,N_21257,N_21719);
nor U28050 (N_28050,N_22846,N_18079);
and U28051 (N_28051,N_18797,N_18225);
nor U28052 (N_28052,N_23377,N_21111);
nor U28053 (N_28053,N_20461,N_21988);
and U28054 (N_28054,N_23895,N_18480);
nor U28055 (N_28055,N_18305,N_22619);
nand U28056 (N_28056,N_21609,N_23307);
nand U28057 (N_28057,N_23686,N_18534);
xnor U28058 (N_28058,N_19658,N_21793);
and U28059 (N_28059,N_22937,N_22538);
nor U28060 (N_28060,N_23483,N_18603);
xor U28061 (N_28061,N_20125,N_20465);
xnor U28062 (N_28062,N_23588,N_20360);
and U28063 (N_28063,N_21973,N_20025);
or U28064 (N_28064,N_23295,N_22656);
and U28065 (N_28065,N_18231,N_20475);
xor U28066 (N_28066,N_19883,N_20105);
nand U28067 (N_28067,N_19059,N_19415);
and U28068 (N_28068,N_18767,N_20474);
or U28069 (N_28069,N_22681,N_20474);
xor U28070 (N_28070,N_22573,N_19675);
or U28071 (N_28071,N_20355,N_18402);
or U28072 (N_28072,N_22103,N_20410);
nor U28073 (N_28073,N_21093,N_22548);
and U28074 (N_28074,N_19867,N_21632);
nor U28075 (N_28075,N_22985,N_22950);
or U28076 (N_28076,N_20833,N_22877);
or U28077 (N_28077,N_23464,N_21592);
or U28078 (N_28078,N_21369,N_22476);
nand U28079 (N_28079,N_22665,N_23323);
or U28080 (N_28080,N_20519,N_19767);
nand U28081 (N_28081,N_21842,N_22210);
nand U28082 (N_28082,N_23936,N_18304);
nand U28083 (N_28083,N_21373,N_22054);
or U28084 (N_28084,N_18873,N_20107);
or U28085 (N_28085,N_20470,N_19140);
xnor U28086 (N_28086,N_20613,N_22896);
xnor U28087 (N_28087,N_22259,N_18849);
nand U28088 (N_28088,N_22985,N_19046);
and U28089 (N_28089,N_21002,N_23135);
nand U28090 (N_28090,N_23310,N_20704);
and U28091 (N_28091,N_22621,N_19096);
nand U28092 (N_28092,N_19572,N_23180);
or U28093 (N_28093,N_20647,N_22502);
or U28094 (N_28094,N_19609,N_21989);
nand U28095 (N_28095,N_20007,N_21200);
and U28096 (N_28096,N_23074,N_22022);
and U28097 (N_28097,N_18100,N_21871);
or U28098 (N_28098,N_20332,N_18261);
nor U28099 (N_28099,N_18161,N_19507);
nor U28100 (N_28100,N_19127,N_22851);
or U28101 (N_28101,N_20992,N_20205);
xor U28102 (N_28102,N_18838,N_20914);
nor U28103 (N_28103,N_19597,N_23768);
nand U28104 (N_28104,N_18762,N_20519);
and U28105 (N_28105,N_20314,N_22119);
nor U28106 (N_28106,N_20889,N_21056);
or U28107 (N_28107,N_23089,N_21461);
xnor U28108 (N_28108,N_19876,N_21333);
or U28109 (N_28109,N_19280,N_23095);
nand U28110 (N_28110,N_19778,N_22341);
xor U28111 (N_28111,N_18585,N_19030);
nand U28112 (N_28112,N_18949,N_19763);
or U28113 (N_28113,N_20812,N_18332);
nand U28114 (N_28114,N_18638,N_19455);
nor U28115 (N_28115,N_23244,N_22068);
or U28116 (N_28116,N_21485,N_21813);
or U28117 (N_28117,N_20372,N_20719);
and U28118 (N_28118,N_23489,N_19161);
nand U28119 (N_28119,N_21511,N_18504);
or U28120 (N_28120,N_21724,N_19307);
nand U28121 (N_28121,N_21263,N_23378);
xnor U28122 (N_28122,N_21243,N_20265);
nor U28123 (N_28123,N_21843,N_22494);
nand U28124 (N_28124,N_20352,N_18431);
xnor U28125 (N_28125,N_20738,N_20858);
nor U28126 (N_28126,N_22108,N_22478);
nand U28127 (N_28127,N_19131,N_18855);
nor U28128 (N_28128,N_18065,N_22192);
and U28129 (N_28129,N_21320,N_22842);
xor U28130 (N_28130,N_18678,N_19857);
and U28131 (N_28131,N_20903,N_19991);
xnor U28132 (N_28132,N_18175,N_21343);
or U28133 (N_28133,N_20672,N_22282);
and U28134 (N_28134,N_18823,N_23583);
nand U28135 (N_28135,N_22905,N_23620);
and U28136 (N_28136,N_19090,N_22171);
and U28137 (N_28137,N_20932,N_19060);
or U28138 (N_28138,N_23991,N_19928);
or U28139 (N_28139,N_18499,N_20039);
xnor U28140 (N_28140,N_19486,N_22021);
xor U28141 (N_28141,N_18463,N_18829);
nor U28142 (N_28142,N_21378,N_20652);
nor U28143 (N_28143,N_21005,N_21185);
nor U28144 (N_28144,N_20345,N_20797);
or U28145 (N_28145,N_21942,N_20740);
and U28146 (N_28146,N_23810,N_23203);
nand U28147 (N_28147,N_19704,N_22060);
or U28148 (N_28148,N_20676,N_21287);
xnor U28149 (N_28149,N_19671,N_20669);
nand U28150 (N_28150,N_19594,N_22259);
xnor U28151 (N_28151,N_21151,N_18364);
or U28152 (N_28152,N_22235,N_23270);
nor U28153 (N_28153,N_19877,N_19339);
nor U28154 (N_28154,N_23116,N_20998);
nor U28155 (N_28155,N_23391,N_19165);
or U28156 (N_28156,N_23833,N_22284);
xor U28157 (N_28157,N_20146,N_20368);
nand U28158 (N_28158,N_18462,N_22149);
or U28159 (N_28159,N_18051,N_20509);
or U28160 (N_28160,N_19976,N_18874);
nand U28161 (N_28161,N_20610,N_22166);
and U28162 (N_28162,N_18342,N_19361);
nor U28163 (N_28163,N_23143,N_21751);
xor U28164 (N_28164,N_23598,N_22066);
or U28165 (N_28165,N_22229,N_23446);
nor U28166 (N_28166,N_20429,N_22259);
or U28167 (N_28167,N_23225,N_19487);
xor U28168 (N_28168,N_20521,N_18214);
or U28169 (N_28169,N_22325,N_20820);
and U28170 (N_28170,N_19314,N_19355);
nand U28171 (N_28171,N_23765,N_21621);
nand U28172 (N_28172,N_18110,N_20367);
and U28173 (N_28173,N_19707,N_19171);
nand U28174 (N_28174,N_19744,N_21000);
or U28175 (N_28175,N_23602,N_21322);
nor U28176 (N_28176,N_22495,N_21567);
and U28177 (N_28177,N_20537,N_19520);
nand U28178 (N_28178,N_23731,N_22694);
or U28179 (N_28179,N_19806,N_18730);
or U28180 (N_28180,N_20216,N_21818);
or U28181 (N_28181,N_19887,N_22597);
or U28182 (N_28182,N_20918,N_21519);
and U28183 (N_28183,N_18685,N_21052);
or U28184 (N_28184,N_19191,N_20224);
nand U28185 (N_28185,N_22579,N_22474);
nand U28186 (N_28186,N_22133,N_19284);
xor U28187 (N_28187,N_22436,N_21649);
and U28188 (N_28188,N_22523,N_20931);
nand U28189 (N_28189,N_20890,N_20271);
or U28190 (N_28190,N_18692,N_21108);
xor U28191 (N_28191,N_21923,N_18900);
nand U28192 (N_28192,N_22952,N_19065);
and U28193 (N_28193,N_19301,N_19190);
and U28194 (N_28194,N_21892,N_20399);
and U28195 (N_28195,N_21856,N_23106);
nand U28196 (N_28196,N_22293,N_23774);
xor U28197 (N_28197,N_21671,N_21830);
nand U28198 (N_28198,N_21307,N_22605);
or U28199 (N_28199,N_22836,N_20872);
and U28200 (N_28200,N_23341,N_20496);
xnor U28201 (N_28201,N_21513,N_21794);
and U28202 (N_28202,N_20103,N_20595);
xor U28203 (N_28203,N_22861,N_19561);
xor U28204 (N_28204,N_18326,N_21657);
nor U28205 (N_28205,N_18340,N_19864);
and U28206 (N_28206,N_23843,N_22577);
nand U28207 (N_28207,N_23923,N_23121);
and U28208 (N_28208,N_19719,N_23127);
or U28209 (N_28209,N_20630,N_23432);
or U28210 (N_28210,N_18441,N_23695);
nor U28211 (N_28211,N_21229,N_19463);
or U28212 (N_28212,N_20843,N_22431);
nor U28213 (N_28213,N_19305,N_22832);
nand U28214 (N_28214,N_23541,N_20141);
or U28215 (N_28215,N_21045,N_18576);
nor U28216 (N_28216,N_22801,N_23116);
and U28217 (N_28217,N_23822,N_22277);
nand U28218 (N_28218,N_18026,N_19609);
or U28219 (N_28219,N_22799,N_21399);
and U28220 (N_28220,N_19350,N_18828);
nor U28221 (N_28221,N_18726,N_19612);
nand U28222 (N_28222,N_18044,N_20476);
xnor U28223 (N_28223,N_19924,N_20043);
nand U28224 (N_28224,N_23029,N_21495);
nand U28225 (N_28225,N_23054,N_21580);
or U28226 (N_28226,N_20121,N_23223);
nand U28227 (N_28227,N_22599,N_19896);
or U28228 (N_28228,N_20964,N_23158);
and U28229 (N_28229,N_22925,N_22993);
or U28230 (N_28230,N_22855,N_18779);
xnor U28231 (N_28231,N_22400,N_18119);
or U28232 (N_28232,N_18193,N_18809);
xor U28233 (N_28233,N_23461,N_19742);
or U28234 (N_28234,N_18671,N_20358);
nand U28235 (N_28235,N_19979,N_18023);
nand U28236 (N_28236,N_20694,N_23434);
nand U28237 (N_28237,N_18777,N_22393);
nor U28238 (N_28238,N_21204,N_23669);
xnor U28239 (N_28239,N_20513,N_22494);
and U28240 (N_28240,N_19097,N_22348);
xnor U28241 (N_28241,N_20776,N_20919);
nand U28242 (N_28242,N_23948,N_20407);
and U28243 (N_28243,N_20173,N_18650);
and U28244 (N_28244,N_20637,N_21722);
nand U28245 (N_28245,N_18600,N_19449);
or U28246 (N_28246,N_19944,N_21224);
and U28247 (N_28247,N_20533,N_18350);
nor U28248 (N_28248,N_19659,N_22354);
and U28249 (N_28249,N_21238,N_19075);
nor U28250 (N_28250,N_19307,N_22241);
and U28251 (N_28251,N_21907,N_18661);
nor U28252 (N_28252,N_22935,N_21796);
nand U28253 (N_28253,N_22256,N_23081);
nand U28254 (N_28254,N_23053,N_19194);
or U28255 (N_28255,N_18509,N_18158);
xnor U28256 (N_28256,N_20028,N_19311);
nand U28257 (N_28257,N_23810,N_23115);
and U28258 (N_28258,N_19242,N_18284);
nor U28259 (N_28259,N_21963,N_20234);
nand U28260 (N_28260,N_22457,N_22408);
nand U28261 (N_28261,N_19605,N_20005);
xor U28262 (N_28262,N_19562,N_23953);
nor U28263 (N_28263,N_21389,N_21569);
nand U28264 (N_28264,N_21873,N_23520);
nor U28265 (N_28265,N_19179,N_22840);
or U28266 (N_28266,N_18505,N_18946);
nand U28267 (N_28267,N_23223,N_19355);
and U28268 (N_28268,N_22740,N_20692);
nor U28269 (N_28269,N_18895,N_21778);
and U28270 (N_28270,N_21092,N_19461);
and U28271 (N_28271,N_22913,N_20680);
nor U28272 (N_28272,N_18937,N_22942);
and U28273 (N_28273,N_20299,N_21883);
or U28274 (N_28274,N_21381,N_19951);
and U28275 (N_28275,N_20626,N_19977);
and U28276 (N_28276,N_21004,N_19555);
and U28277 (N_28277,N_21734,N_18064);
nand U28278 (N_28278,N_19341,N_22407);
or U28279 (N_28279,N_21661,N_19768);
and U28280 (N_28280,N_23370,N_23632);
nor U28281 (N_28281,N_22232,N_18978);
or U28282 (N_28282,N_23143,N_20965);
and U28283 (N_28283,N_21449,N_23752);
nor U28284 (N_28284,N_22314,N_22680);
and U28285 (N_28285,N_23732,N_23522);
nand U28286 (N_28286,N_22037,N_19963);
or U28287 (N_28287,N_23149,N_20816);
nor U28288 (N_28288,N_22141,N_18796);
nor U28289 (N_28289,N_19917,N_20217);
nand U28290 (N_28290,N_18433,N_19762);
xor U28291 (N_28291,N_22509,N_21815);
nor U28292 (N_28292,N_20665,N_23629);
xnor U28293 (N_28293,N_19681,N_19500);
nor U28294 (N_28294,N_19196,N_20231);
xnor U28295 (N_28295,N_20709,N_19506);
and U28296 (N_28296,N_23949,N_18305);
nand U28297 (N_28297,N_21500,N_19968);
nand U28298 (N_28298,N_21381,N_23916);
nand U28299 (N_28299,N_20201,N_19080);
or U28300 (N_28300,N_21445,N_20955);
nor U28301 (N_28301,N_19207,N_18240);
nand U28302 (N_28302,N_22968,N_18076);
or U28303 (N_28303,N_20971,N_22981);
nor U28304 (N_28304,N_20535,N_20143);
nor U28305 (N_28305,N_19106,N_22888);
nor U28306 (N_28306,N_21234,N_23385);
xor U28307 (N_28307,N_18586,N_20092);
or U28308 (N_28308,N_23981,N_22253);
and U28309 (N_28309,N_18939,N_18257);
nand U28310 (N_28310,N_20535,N_21852);
and U28311 (N_28311,N_21565,N_20132);
nor U28312 (N_28312,N_21599,N_23304);
and U28313 (N_28313,N_19126,N_18046);
and U28314 (N_28314,N_22802,N_19371);
nand U28315 (N_28315,N_23568,N_20457);
and U28316 (N_28316,N_18095,N_20073);
xnor U28317 (N_28317,N_20148,N_21246);
or U28318 (N_28318,N_23077,N_18746);
nand U28319 (N_28319,N_18403,N_21348);
and U28320 (N_28320,N_19893,N_19796);
nand U28321 (N_28321,N_22254,N_18971);
and U28322 (N_28322,N_20904,N_23291);
or U28323 (N_28323,N_23020,N_20411);
or U28324 (N_28324,N_21470,N_21924);
nor U28325 (N_28325,N_21786,N_22717);
or U28326 (N_28326,N_23973,N_18092);
nor U28327 (N_28327,N_20534,N_23954);
and U28328 (N_28328,N_22387,N_23656);
xor U28329 (N_28329,N_22239,N_19426);
or U28330 (N_28330,N_19242,N_19304);
xnor U28331 (N_28331,N_22797,N_21796);
or U28332 (N_28332,N_21323,N_23914);
or U28333 (N_28333,N_23720,N_21199);
nand U28334 (N_28334,N_21084,N_23568);
xor U28335 (N_28335,N_21046,N_22145);
and U28336 (N_28336,N_18863,N_18257);
nor U28337 (N_28337,N_19607,N_18093);
xnor U28338 (N_28338,N_23889,N_19562);
xor U28339 (N_28339,N_20654,N_18865);
and U28340 (N_28340,N_19212,N_19705);
xor U28341 (N_28341,N_18093,N_23933);
nor U28342 (N_28342,N_19231,N_19007);
and U28343 (N_28343,N_23402,N_21656);
nor U28344 (N_28344,N_23405,N_18853);
xnor U28345 (N_28345,N_18362,N_23858);
nand U28346 (N_28346,N_18443,N_19573);
or U28347 (N_28347,N_19345,N_19290);
or U28348 (N_28348,N_21695,N_21995);
nand U28349 (N_28349,N_22436,N_23655);
xor U28350 (N_28350,N_21321,N_21097);
xor U28351 (N_28351,N_20685,N_18909);
nand U28352 (N_28352,N_23711,N_18536);
and U28353 (N_28353,N_20253,N_21549);
or U28354 (N_28354,N_18762,N_19533);
or U28355 (N_28355,N_19684,N_20211);
and U28356 (N_28356,N_21064,N_23764);
or U28357 (N_28357,N_22847,N_19102);
nand U28358 (N_28358,N_20089,N_23031);
nand U28359 (N_28359,N_22459,N_20678);
nand U28360 (N_28360,N_22702,N_23094);
xnor U28361 (N_28361,N_23881,N_23237);
or U28362 (N_28362,N_19055,N_19376);
or U28363 (N_28363,N_19227,N_18933);
or U28364 (N_28364,N_23975,N_22881);
nor U28365 (N_28365,N_20168,N_23778);
and U28366 (N_28366,N_20511,N_23121);
nand U28367 (N_28367,N_23505,N_23014);
or U28368 (N_28368,N_18201,N_21585);
nor U28369 (N_28369,N_18623,N_21036);
or U28370 (N_28370,N_22068,N_22939);
or U28371 (N_28371,N_19726,N_19811);
xnor U28372 (N_28372,N_18982,N_19076);
nand U28373 (N_28373,N_22781,N_22335);
xnor U28374 (N_28374,N_19823,N_21396);
and U28375 (N_28375,N_23515,N_19232);
or U28376 (N_28376,N_18886,N_18971);
and U28377 (N_28377,N_18839,N_22503);
nand U28378 (N_28378,N_21130,N_18074);
nand U28379 (N_28379,N_21502,N_23596);
and U28380 (N_28380,N_23022,N_22591);
or U28381 (N_28381,N_18822,N_19180);
nor U28382 (N_28382,N_21375,N_21791);
and U28383 (N_28383,N_23912,N_20835);
xnor U28384 (N_28384,N_22880,N_20905);
nor U28385 (N_28385,N_22988,N_18328);
and U28386 (N_28386,N_20952,N_20008);
nand U28387 (N_28387,N_19963,N_23026);
nand U28388 (N_28388,N_22748,N_19274);
xnor U28389 (N_28389,N_23913,N_23646);
nand U28390 (N_28390,N_23602,N_19428);
xnor U28391 (N_28391,N_19602,N_21435);
xor U28392 (N_28392,N_19406,N_21160);
xor U28393 (N_28393,N_20794,N_22834);
nand U28394 (N_28394,N_21133,N_19480);
and U28395 (N_28395,N_20846,N_21681);
nand U28396 (N_28396,N_23658,N_23396);
nor U28397 (N_28397,N_23366,N_18191);
nor U28398 (N_28398,N_19642,N_23560);
or U28399 (N_28399,N_19024,N_21474);
nand U28400 (N_28400,N_23514,N_19658);
or U28401 (N_28401,N_18074,N_21172);
xor U28402 (N_28402,N_22293,N_20371);
or U28403 (N_28403,N_21403,N_21474);
nand U28404 (N_28404,N_19465,N_23863);
xnor U28405 (N_28405,N_18437,N_23092);
nand U28406 (N_28406,N_19702,N_23089);
and U28407 (N_28407,N_19025,N_23554);
xor U28408 (N_28408,N_20535,N_20703);
nand U28409 (N_28409,N_23622,N_22666);
nand U28410 (N_28410,N_18069,N_19162);
and U28411 (N_28411,N_22642,N_19729);
nand U28412 (N_28412,N_18294,N_21740);
xor U28413 (N_28413,N_22220,N_21095);
nor U28414 (N_28414,N_22429,N_21894);
nand U28415 (N_28415,N_22793,N_22340);
or U28416 (N_28416,N_21011,N_19634);
xor U28417 (N_28417,N_20295,N_19032);
nor U28418 (N_28418,N_18845,N_18345);
and U28419 (N_28419,N_22872,N_20228);
nor U28420 (N_28420,N_20111,N_18926);
xor U28421 (N_28421,N_23177,N_20982);
nand U28422 (N_28422,N_23990,N_22919);
and U28423 (N_28423,N_19837,N_18522);
nand U28424 (N_28424,N_23847,N_21008);
xnor U28425 (N_28425,N_23263,N_19728);
and U28426 (N_28426,N_18161,N_20676);
and U28427 (N_28427,N_19689,N_23727);
nor U28428 (N_28428,N_20953,N_22028);
nor U28429 (N_28429,N_20337,N_21088);
xor U28430 (N_28430,N_22855,N_23357);
nor U28431 (N_28431,N_21910,N_23561);
nand U28432 (N_28432,N_18116,N_19203);
xor U28433 (N_28433,N_19889,N_18310);
or U28434 (N_28434,N_22355,N_23520);
and U28435 (N_28435,N_18284,N_21132);
and U28436 (N_28436,N_22152,N_23623);
nand U28437 (N_28437,N_22447,N_21079);
and U28438 (N_28438,N_23530,N_22717);
or U28439 (N_28439,N_20187,N_19628);
nor U28440 (N_28440,N_19746,N_21937);
nand U28441 (N_28441,N_20647,N_18800);
nor U28442 (N_28442,N_20913,N_20255);
nor U28443 (N_28443,N_22857,N_22269);
or U28444 (N_28444,N_21088,N_23127);
and U28445 (N_28445,N_19077,N_18521);
nand U28446 (N_28446,N_22604,N_22724);
nand U28447 (N_28447,N_20166,N_22075);
nor U28448 (N_28448,N_18188,N_20733);
xnor U28449 (N_28449,N_23361,N_22750);
nand U28450 (N_28450,N_19143,N_19790);
and U28451 (N_28451,N_20290,N_20465);
xor U28452 (N_28452,N_19296,N_19829);
nor U28453 (N_28453,N_20487,N_20139);
and U28454 (N_28454,N_19588,N_22654);
or U28455 (N_28455,N_22765,N_22188);
nand U28456 (N_28456,N_19921,N_18154);
xor U28457 (N_28457,N_18966,N_19714);
and U28458 (N_28458,N_18579,N_20806);
and U28459 (N_28459,N_18187,N_22744);
nand U28460 (N_28460,N_20804,N_23947);
and U28461 (N_28461,N_20269,N_19120);
nor U28462 (N_28462,N_21183,N_21439);
nor U28463 (N_28463,N_22629,N_21633);
xnor U28464 (N_28464,N_18491,N_23272);
nor U28465 (N_28465,N_20988,N_19123);
xor U28466 (N_28466,N_19817,N_20912);
nand U28467 (N_28467,N_19368,N_21884);
and U28468 (N_28468,N_19589,N_20186);
or U28469 (N_28469,N_23035,N_20410);
nand U28470 (N_28470,N_19817,N_22919);
xnor U28471 (N_28471,N_22795,N_23221);
nand U28472 (N_28472,N_18314,N_20228);
or U28473 (N_28473,N_21415,N_22378);
nand U28474 (N_28474,N_23235,N_20704);
xor U28475 (N_28475,N_19297,N_20481);
nor U28476 (N_28476,N_19543,N_22175);
xnor U28477 (N_28477,N_23728,N_22400);
nor U28478 (N_28478,N_18163,N_22258);
nand U28479 (N_28479,N_22982,N_19198);
xnor U28480 (N_28480,N_23378,N_19611);
or U28481 (N_28481,N_18983,N_19473);
and U28482 (N_28482,N_21482,N_18955);
and U28483 (N_28483,N_22562,N_18369);
xor U28484 (N_28484,N_21046,N_21703);
xnor U28485 (N_28485,N_22698,N_19675);
or U28486 (N_28486,N_18765,N_20518);
nand U28487 (N_28487,N_18499,N_19179);
or U28488 (N_28488,N_18662,N_20643);
nor U28489 (N_28489,N_21757,N_18624);
xnor U28490 (N_28490,N_18584,N_21952);
and U28491 (N_28491,N_18669,N_19599);
nand U28492 (N_28492,N_18331,N_19288);
xor U28493 (N_28493,N_22452,N_18671);
nand U28494 (N_28494,N_18748,N_19116);
and U28495 (N_28495,N_21734,N_21515);
nor U28496 (N_28496,N_23084,N_18085);
nand U28497 (N_28497,N_18211,N_23778);
or U28498 (N_28498,N_18514,N_19375);
nand U28499 (N_28499,N_23905,N_19130);
and U28500 (N_28500,N_21756,N_22455);
xnor U28501 (N_28501,N_19157,N_21622);
xnor U28502 (N_28502,N_20085,N_22726);
or U28503 (N_28503,N_23978,N_19170);
or U28504 (N_28504,N_18197,N_21228);
and U28505 (N_28505,N_19402,N_18321);
and U28506 (N_28506,N_20953,N_18105);
and U28507 (N_28507,N_20439,N_22097);
nand U28508 (N_28508,N_18861,N_18592);
xnor U28509 (N_28509,N_20026,N_20346);
nand U28510 (N_28510,N_22493,N_20267);
xor U28511 (N_28511,N_22037,N_19718);
nand U28512 (N_28512,N_19859,N_22864);
xnor U28513 (N_28513,N_23427,N_23407);
or U28514 (N_28514,N_20117,N_21378);
xor U28515 (N_28515,N_22735,N_21540);
nand U28516 (N_28516,N_23833,N_23012);
xnor U28517 (N_28517,N_19546,N_18249);
nand U28518 (N_28518,N_22436,N_18209);
xor U28519 (N_28519,N_23785,N_19273);
nand U28520 (N_28520,N_18043,N_19564);
or U28521 (N_28521,N_23634,N_21131);
or U28522 (N_28522,N_23100,N_23728);
or U28523 (N_28523,N_21268,N_23311);
nand U28524 (N_28524,N_20787,N_18642);
nand U28525 (N_28525,N_21228,N_21782);
nand U28526 (N_28526,N_18379,N_18799);
and U28527 (N_28527,N_18312,N_23628);
and U28528 (N_28528,N_21839,N_21967);
and U28529 (N_28529,N_20651,N_22587);
or U28530 (N_28530,N_20464,N_23544);
nor U28531 (N_28531,N_18379,N_20247);
or U28532 (N_28532,N_20048,N_23365);
or U28533 (N_28533,N_22618,N_23630);
or U28534 (N_28534,N_19975,N_19698);
and U28535 (N_28535,N_22062,N_22504);
nor U28536 (N_28536,N_19491,N_23757);
and U28537 (N_28537,N_19863,N_18318);
nor U28538 (N_28538,N_20303,N_21110);
nor U28539 (N_28539,N_18235,N_19661);
and U28540 (N_28540,N_19918,N_22555);
nor U28541 (N_28541,N_18003,N_22923);
nor U28542 (N_28542,N_20763,N_21941);
or U28543 (N_28543,N_20993,N_20338);
xnor U28544 (N_28544,N_21033,N_23543);
and U28545 (N_28545,N_19816,N_21735);
xor U28546 (N_28546,N_22757,N_18671);
or U28547 (N_28547,N_23745,N_18222);
or U28548 (N_28548,N_19040,N_22759);
and U28549 (N_28549,N_20235,N_20955);
nor U28550 (N_28550,N_19091,N_18964);
or U28551 (N_28551,N_22591,N_18036);
nand U28552 (N_28552,N_21257,N_21038);
or U28553 (N_28553,N_19506,N_19265);
and U28554 (N_28554,N_20268,N_22009);
and U28555 (N_28555,N_22099,N_21912);
or U28556 (N_28556,N_20584,N_21292);
or U28557 (N_28557,N_23529,N_22203);
nand U28558 (N_28558,N_22210,N_22567);
or U28559 (N_28559,N_19153,N_23580);
and U28560 (N_28560,N_20549,N_20356);
or U28561 (N_28561,N_23065,N_20685);
nor U28562 (N_28562,N_22248,N_21003);
xnor U28563 (N_28563,N_22472,N_23766);
or U28564 (N_28564,N_23940,N_19665);
xnor U28565 (N_28565,N_19455,N_21107);
nor U28566 (N_28566,N_23444,N_19213);
nand U28567 (N_28567,N_18354,N_21536);
or U28568 (N_28568,N_23413,N_22463);
or U28569 (N_28569,N_22096,N_18105);
and U28570 (N_28570,N_22309,N_22340);
and U28571 (N_28571,N_19746,N_23956);
xnor U28572 (N_28572,N_20129,N_23402);
and U28573 (N_28573,N_18765,N_20593);
and U28574 (N_28574,N_20275,N_20362);
or U28575 (N_28575,N_22550,N_21319);
or U28576 (N_28576,N_20764,N_20461);
and U28577 (N_28577,N_22601,N_23901);
or U28578 (N_28578,N_20565,N_21673);
or U28579 (N_28579,N_23535,N_20742);
xor U28580 (N_28580,N_19051,N_20505);
or U28581 (N_28581,N_23164,N_19855);
and U28582 (N_28582,N_18761,N_19734);
or U28583 (N_28583,N_22164,N_22142);
xor U28584 (N_28584,N_18330,N_18133);
xor U28585 (N_28585,N_20077,N_23291);
or U28586 (N_28586,N_21537,N_23659);
nor U28587 (N_28587,N_22517,N_21874);
xnor U28588 (N_28588,N_22307,N_19218);
nand U28589 (N_28589,N_23630,N_23312);
or U28590 (N_28590,N_21702,N_18525);
nor U28591 (N_28591,N_23187,N_18935);
nor U28592 (N_28592,N_23482,N_23180);
or U28593 (N_28593,N_21700,N_22479);
and U28594 (N_28594,N_18722,N_19437);
and U28595 (N_28595,N_20496,N_19247);
or U28596 (N_28596,N_23602,N_20283);
and U28597 (N_28597,N_18383,N_21335);
xor U28598 (N_28598,N_20606,N_18831);
or U28599 (N_28599,N_22716,N_18827);
nand U28600 (N_28600,N_20114,N_18103);
xnor U28601 (N_28601,N_18729,N_23537);
nand U28602 (N_28602,N_23930,N_23838);
and U28603 (N_28603,N_21552,N_19097);
xnor U28604 (N_28604,N_23547,N_20601);
nand U28605 (N_28605,N_22589,N_23739);
nand U28606 (N_28606,N_20834,N_20812);
nand U28607 (N_28607,N_23918,N_23318);
nand U28608 (N_28608,N_18761,N_18641);
xnor U28609 (N_28609,N_19785,N_20635);
or U28610 (N_28610,N_23138,N_19795);
and U28611 (N_28611,N_21057,N_19001);
nand U28612 (N_28612,N_20178,N_19091);
or U28613 (N_28613,N_22469,N_23295);
nor U28614 (N_28614,N_21405,N_18453);
xnor U28615 (N_28615,N_23515,N_21609);
or U28616 (N_28616,N_19401,N_21306);
nor U28617 (N_28617,N_18623,N_18995);
and U28618 (N_28618,N_22134,N_20119);
nand U28619 (N_28619,N_20438,N_21161);
nor U28620 (N_28620,N_23600,N_23780);
xnor U28621 (N_28621,N_19825,N_20859);
xnor U28622 (N_28622,N_22017,N_22350);
nor U28623 (N_28623,N_19402,N_19389);
nand U28624 (N_28624,N_22815,N_20113);
nand U28625 (N_28625,N_22291,N_20529);
and U28626 (N_28626,N_22076,N_18487);
nor U28627 (N_28627,N_22794,N_18776);
xor U28628 (N_28628,N_23248,N_23223);
nand U28629 (N_28629,N_19212,N_22616);
and U28630 (N_28630,N_20707,N_21877);
nor U28631 (N_28631,N_23369,N_19934);
nand U28632 (N_28632,N_22298,N_18623);
nand U28633 (N_28633,N_19301,N_22296);
or U28634 (N_28634,N_23182,N_18099);
nor U28635 (N_28635,N_19710,N_22321);
nand U28636 (N_28636,N_18989,N_18316);
and U28637 (N_28637,N_20030,N_20115);
nor U28638 (N_28638,N_19940,N_23520);
or U28639 (N_28639,N_18766,N_18416);
xor U28640 (N_28640,N_23114,N_19288);
nand U28641 (N_28641,N_19233,N_18028);
and U28642 (N_28642,N_18893,N_21041);
xnor U28643 (N_28643,N_19562,N_22529);
nand U28644 (N_28644,N_18517,N_20349);
or U28645 (N_28645,N_21930,N_20652);
xor U28646 (N_28646,N_19619,N_22286);
or U28647 (N_28647,N_22173,N_19659);
nand U28648 (N_28648,N_18074,N_19572);
nand U28649 (N_28649,N_20465,N_19750);
nand U28650 (N_28650,N_20788,N_21150);
nor U28651 (N_28651,N_19446,N_22984);
xnor U28652 (N_28652,N_19745,N_23905);
and U28653 (N_28653,N_21183,N_18570);
xnor U28654 (N_28654,N_19458,N_23505);
nand U28655 (N_28655,N_22991,N_23975);
nor U28656 (N_28656,N_21742,N_20722);
and U28657 (N_28657,N_20885,N_19310);
or U28658 (N_28658,N_19325,N_23810);
and U28659 (N_28659,N_20624,N_20790);
xor U28660 (N_28660,N_19803,N_21705);
nor U28661 (N_28661,N_22343,N_21413);
or U28662 (N_28662,N_23272,N_23684);
nor U28663 (N_28663,N_20001,N_21980);
xor U28664 (N_28664,N_22368,N_22729);
and U28665 (N_28665,N_18988,N_18513);
nor U28666 (N_28666,N_20654,N_22716);
and U28667 (N_28667,N_18573,N_21345);
xnor U28668 (N_28668,N_21692,N_19356);
xnor U28669 (N_28669,N_19043,N_18556);
nand U28670 (N_28670,N_18574,N_19480);
or U28671 (N_28671,N_18511,N_18735);
or U28672 (N_28672,N_23616,N_22405);
nand U28673 (N_28673,N_23038,N_21986);
xnor U28674 (N_28674,N_23455,N_22327);
xor U28675 (N_28675,N_22814,N_21428);
or U28676 (N_28676,N_23880,N_22351);
xor U28677 (N_28677,N_20580,N_19971);
or U28678 (N_28678,N_19340,N_19908);
or U28679 (N_28679,N_21296,N_22970);
nand U28680 (N_28680,N_19868,N_19176);
or U28681 (N_28681,N_22408,N_19165);
and U28682 (N_28682,N_18117,N_20060);
xnor U28683 (N_28683,N_18393,N_20802);
nor U28684 (N_28684,N_21802,N_22040);
or U28685 (N_28685,N_20945,N_22211);
xor U28686 (N_28686,N_19463,N_19285);
or U28687 (N_28687,N_18023,N_23432);
or U28688 (N_28688,N_19562,N_18911);
xnor U28689 (N_28689,N_21919,N_18848);
or U28690 (N_28690,N_21443,N_20814);
nand U28691 (N_28691,N_21352,N_18075);
or U28692 (N_28692,N_23068,N_22541);
nor U28693 (N_28693,N_21829,N_23095);
or U28694 (N_28694,N_23333,N_18303);
or U28695 (N_28695,N_23088,N_20344);
nor U28696 (N_28696,N_23156,N_18692);
and U28697 (N_28697,N_18025,N_20783);
and U28698 (N_28698,N_20221,N_19237);
nor U28699 (N_28699,N_18874,N_22171);
nor U28700 (N_28700,N_21979,N_21677);
nand U28701 (N_28701,N_23001,N_21696);
nand U28702 (N_28702,N_18756,N_20111);
nor U28703 (N_28703,N_19957,N_23564);
nand U28704 (N_28704,N_22655,N_18536);
nor U28705 (N_28705,N_21249,N_20852);
and U28706 (N_28706,N_21331,N_21215);
or U28707 (N_28707,N_20006,N_18032);
and U28708 (N_28708,N_22428,N_19929);
xnor U28709 (N_28709,N_20663,N_19908);
nor U28710 (N_28710,N_23102,N_21759);
xor U28711 (N_28711,N_21669,N_18900);
nand U28712 (N_28712,N_20325,N_21809);
xor U28713 (N_28713,N_23971,N_19251);
nand U28714 (N_28714,N_19290,N_19933);
nand U28715 (N_28715,N_18362,N_19418);
and U28716 (N_28716,N_19895,N_18643);
xnor U28717 (N_28717,N_21368,N_18700);
and U28718 (N_28718,N_18471,N_20721);
nor U28719 (N_28719,N_22416,N_23471);
nand U28720 (N_28720,N_23765,N_18134);
nand U28721 (N_28721,N_20344,N_22477);
nor U28722 (N_28722,N_19509,N_21528);
and U28723 (N_28723,N_22761,N_19079);
nor U28724 (N_28724,N_21076,N_21696);
or U28725 (N_28725,N_20541,N_22186);
xor U28726 (N_28726,N_23765,N_20608);
nor U28727 (N_28727,N_18741,N_21798);
nand U28728 (N_28728,N_18809,N_21253);
and U28729 (N_28729,N_22020,N_22148);
or U28730 (N_28730,N_20180,N_22881);
and U28731 (N_28731,N_19608,N_19384);
nand U28732 (N_28732,N_21030,N_23099);
nor U28733 (N_28733,N_22709,N_21835);
and U28734 (N_28734,N_19188,N_20913);
and U28735 (N_28735,N_20597,N_19441);
or U28736 (N_28736,N_18369,N_18896);
or U28737 (N_28737,N_21176,N_20510);
and U28738 (N_28738,N_21923,N_19231);
nand U28739 (N_28739,N_21522,N_19363);
nand U28740 (N_28740,N_18996,N_22598);
and U28741 (N_28741,N_18532,N_22262);
or U28742 (N_28742,N_21082,N_18887);
nand U28743 (N_28743,N_22957,N_19594);
nor U28744 (N_28744,N_19947,N_20780);
nand U28745 (N_28745,N_23595,N_18576);
or U28746 (N_28746,N_18527,N_19368);
xnor U28747 (N_28747,N_21732,N_19312);
and U28748 (N_28748,N_20636,N_23293);
nand U28749 (N_28749,N_19144,N_18929);
or U28750 (N_28750,N_18561,N_20786);
and U28751 (N_28751,N_19840,N_18130);
xor U28752 (N_28752,N_22136,N_23456);
nor U28753 (N_28753,N_18314,N_22800);
nand U28754 (N_28754,N_21522,N_20572);
nor U28755 (N_28755,N_22008,N_20720);
xnor U28756 (N_28756,N_18581,N_23240);
nor U28757 (N_28757,N_22734,N_19530);
or U28758 (N_28758,N_20725,N_19428);
or U28759 (N_28759,N_22450,N_22233);
nand U28760 (N_28760,N_19886,N_23169);
or U28761 (N_28761,N_19592,N_19229);
nand U28762 (N_28762,N_20780,N_18615);
and U28763 (N_28763,N_20279,N_18661);
nor U28764 (N_28764,N_21714,N_18038);
nor U28765 (N_28765,N_20094,N_21737);
nor U28766 (N_28766,N_20856,N_22671);
nor U28767 (N_28767,N_18545,N_23854);
xnor U28768 (N_28768,N_23641,N_20773);
xnor U28769 (N_28769,N_19909,N_21780);
and U28770 (N_28770,N_18844,N_20906);
xor U28771 (N_28771,N_23593,N_18453);
or U28772 (N_28772,N_20481,N_21114);
nand U28773 (N_28773,N_20912,N_20181);
and U28774 (N_28774,N_21900,N_19358);
xor U28775 (N_28775,N_22723,N_22718);
or U28776 (N_28776,N_23061,N_20173);
nor U28777 (N_28777,N_19200,N_18882);
nor U28778 (N_28778,N_23454,N_22433);
nor U28779 (N_28779,N_23660,N_23268);
or U28780 (N_28780,N_20610,N_18015);
nor U28781 (N_28781,N_18814,N_18886);
nand U28782 (N_28782,N_22997,N_18668);
and U28783 (N_28783,N_18530,N_23375);
and U28784 (N_28784,N_23507,N_23560);
xor U28785 (N_28785,N_21268,N_20088);
or U28786 (N_28786,N_19933,N_21780);
and U28787 (N_28787,N_18792,N_22571);
nand U28788 (N_28788,N_19840,N_21901);
nand U28789 (N_28789,N_19348,N_19186);
nor U28790 (N_28790,N_21082,N_19436);
xor U28791 (N_28791,N_21451,N_22503);
nor U28792 (N_28792,N_21220,N_23927);
xor U28793 (N_28793,N_22071,N_19859);
xor U28794 (N_28794,N_22385,N_20844);
xnor U28795 (N_28795,N_20241,N_19639);
and U28796 (N_28796,N_21926,N_22163);
nor U28797 (N_28797,N_21883,N_20543);
xnor U28798 (N_28798,N_19658,N_18639);
and U28799 (N_28799,N_19072,N_19930);
or U28800 (N_28800,N_20577,N_20636);
nand U28801 (N_28801,N_19372,N_23250);
and U28802 (N_28802,N_21742,N_23452);
or U28803 (N_28803,N_19061,N_22290);
or U28804 (N_28804,N_19557,N_22597);
and U28805 (N_28805,N_19107,N_19287);
xnor U28806 (N_28806,N_21677,N_20713);
and U28807 (N_28807,N_21372,N_23859);
xor U28808 (N_28808,N_18117,N_20509);
and U28809 (N_28809,N_20378,N_19850);
and U28810 (N_28810,N_21522,N_19532);
and U28811 (N_28811,N_21405,N_23815);
or U28812 (N_28812,N_19174,N_20929);
nor U28813 (N_28813,N_23052,N_20748);
xor U28814 (N_28814,N_18165,N_21541);
nor U28815 (N_28815,N_19366,N_23480);
or U28816 (N_28816,N_21056,N_21237);
and U28817 (N_28817,N_19909,N_23375);
or U28818 (N_28818,N_19335,N_21432);
xnor U28819 (N_28819,N_23194,N_21333);
or U28820 (N_28820,N_19298,N_22182);
nor U28821 (N_28821,N_20001,N_21075);
or U28822 (N_28822,N_20663,N_21763);
and U28823 (N_28823,N_18410,N_20088);
nand U28824 (N_28824,N_23456,N_19283);
or U28825 (N_28825,N_18755,N_23145);
and U28826 (N_28826,N_19466,N_20602);
and U28827 (N_28827,N_21430,N_19715);
nor U28828 (N_28828,N_23906,N_23073);
and U28829 (N_28829,N_19758,N_21842);
xor U28830 (N_28830,N_20762,N_20732);
nand U28831 (N_28831,N_19081,N_23115);
nand U28832 (N_28832,N_19395,N_22913);
and U28833 (N_28833,N_22671,N_20395);
or U28834 (N_28834,N_20393,N_23708);
or U28835 (N_28835,N_20937,N_18938);
nor U28836 (N_28836,N_19718,N_22584);
or U28837 (N_28837,N_23534,N_19894);
nor U28838 (N_28838,N_22069,N_19677);
and U28839 (N_28839,N_23078,N_20751);
nand U28840 (N_28840,N_18950,N_23079);
nand U28841 (N_28841,N_21641,N_21922);
nor U28842 (N_28842,N_18321,N_23620);
or U28843 (N_28843,N_20520,N_21860);
or U28844 (N_28844,N_21438,N_23549);
and U28845 (N_28845,N_20773,N_19449);
or U28846 (N_28846,N_20486,N_23227);
nand U28847 (N_28847,N_20073,N_21746);
xor U28848 (N_28848,N_18538,N_21708);
nor U28849 (N_28849,N_18803,N_20710);
nand U28850 (N_28850,N_19225,N_18492);
and U28851 (N_28851,N_20768,N_21853);
xor U28852 (N_28852,N_21365,N_21764);
nand U28853 (N_28853,N_23880,N_22925);
xnor U28854 (N_28854,N_18794,N_20043);
or U28855 (N_28855,N_22071,N_19419);
nor U28856 (N_28856,N_23532,N_23911);
xor U28857 (N_28857,N_22570,N_21052);
xor U28858 (N_28858,N_18009,N_21849);
or U28859 (N_28859,N_21354,N_21084);
or U28860 (N_28860,N_21680,N_21980);
or U28861 (N_28861,N_21620,N_22935);
nor U28862 (N_28862,N_22231,N_20887);
xnor U28863 (N_28863,N_18774,N_19746);
and U28864 (N_28864,N_20563,N_18148);
xnor U28865 (N_28865,N_18935,N_19351);
and U28866 (N_28866,N_21317,N_20655);
or U28867 (N_28867,N_23673,N_23723);
xor U28868 (N_28868,N_22516,N_19859);
and U28869 (N_28869,N_22268,N_23368);
nand U28870 (N_28870,N_23493,N_18369);
or U28871 (N_28871,N_23831,N_21178);
or U28872 (N_28872,N_21633,N_23649);
and U28873 (N_28873,N_22407,N_21418);
nand U28874 (N_28874,N_22738,N_18418);
or U28875 (N_28875,N_23120,N_23544);
nand U28876 (N_28876,N_18173,N_22158);
nand U28877 (N_28877,N_23330,N_22012);
nor U28878 (N_28878,N_22811,N_22736);
nor U28879 (N_28879,N_20790,N_21533);
nor U28880 (N_28880,N_23460,N_18566);
nand U28881 (N_28881,N_22448,N_23893);
xor U28882 (N_28882,N_22859,N_18022);
or U28883 (N_28883,N_18893,N_18957);
and U28884 (N_28884,N_20013,N_22137);
nand U28885 (N_28885,N_21012,N_22911);
nor U28886 (N_28886,N_22831,N_18703);
and U28887 (N_28887,N_23335,N_19087);
nor U28888 (N_28888,N_23813,N_21625);
nor U28889 (N_28889,N_23119,N_21467);
xnor U28890 (N_28890,N_22576,N_23963);
nand U28891 (N_28891,N_22406,N_21634);
or U28892 (N_28892,N_18350,N_21714);
nand U28893 (N_28893,N_21643,N_23539);
and U28894 (N_28894,N_20636,N_19575);
nand U28895 (N_28895,N_20085,N_22631);
nor U28896 (N_28896,N_18311,N_23667);
nand U28897 (N_28897,N_22452,N_20542);
nor U28898 (N_28898,N_23314,N_20196);
or U28899 (N_28899,N_20476,N_21925);
xnor U28900 (N_28900,N_22847,N_23394);
nand U28901 (N_28901,N_20599,N_22980);
or U28902 (N_28902,N_19410,N_18098);
xnor U28903 (N_28903,N_18378,N_19102);
and U28904 (N_28904,N_21421,N_18269);
nor U28905 (N_28905,N_19723,N_19993);
nand U28906 (N_28906,N_19169,N_23447);
nand U28907 (N_28907,N_19825,N_18835);
nand U28908 (N_28908,N_20994,N_23674);
nand U28909 (N_28909,N_18006,N_20668);
or U28910 (N_28910,N_19442,N_23507);
xor U28911 (N_28911,N_19730,N_21106);
or U28912 (N_28912,N_20041,N_19958);
nand U28913 (N_28913,N_18929,N_21338);
and U28914 (N_28914,N_23804,N_20872);
nor U28915 (N_28915,N_22259,N_20286);
nand U28916 (N_28916,N_22271,N_19781);
xor U28917 (N_28917,N_19752,N_21701);
xor U28918 (N_28918,N_18279,N_22394);
nand U28919 (N_28919,N_22970,N_22736);
and U28920 (N_28920,N_21567,N_21409);
or U28921 (N_28921,N_23485,N_23718);
xnor U28922 (N_28922,N_21354,N_20221);
and U28923 (N_28923,N_23902,N_23749);
nor U28924 (N_28924,N_21828,N_22739);
nor U28925 (N_28925,N_19950,N_23550);
and U28926 (N_28926,N_22582,N_18530);
and U28927 (N_28927,N_20108,N_18303);
xor U28928 (N_28928,N_23561,N_19144);
or U28929 (N_28929,N_21654,N_22056);
nor U28930 (N_28930,N_22621,N_23088);
or U28931 (N_28931,N_20718,N_23037);
xnor U28932 (N_28932,N_19348,N_22223);
nand U28933 (N_28933,N_22311,N_23564);
and U28934 (N_28934,N_19777,N_20310);
nor U28935 (N_28935,N_22786,N_18791);
nor U28936 (N_28936,N_23642,N_18668);
and U28937 (N_28937,N_23787,N_19642);
xor U28938 (N_28938,N_20244,N_21180);
or U28939 (N_28939,N_23396,N_23719);
or U28940 (N_28940,N_19799,N_22867);
nand U28941 (N_28941,N_23366,N_22023);
nor U28942 (N_28942,N_18296,N_22100);
and U28943 (N_28943,N_22668,N_23233);
or U28944 (N_28944,N_20638,N_18652);
nand U28945 (N_28945,N_20088,N_18465);
and U28946 (N_28946,N_19703,N_20446);
nor U28947 (N_28947,N_21626,N_19568);
or U28948 (N_28948,N_23195,N_21218);
nand U28949 (N_28949,N_20506,N_19361);
nand U28950 (N_28950,N_19086,N_23007);
xor U28951 (N_28951,N_20209,N_22362);
xor U28952 (N_28952,N_20409,N_18474);
xnor U28953 (N_28953,N_19916,N_21180);
nand U28954 (N_28954,N_19059,N_18450);
or U28955 (N_28955,N_19738,N_18975);
or U28956 (N_28956,N_22853,N_20972);
or U28957 (N_28957,N_21877,N_23247);
and U28958 (N_28958,N_20277,N_20444);
or U28959 (N_28959,N_22446,N_21531);
nor U28960 (N_28960,N_23113,N_21615);
nor U28961 (N_28961,N_23259,N_18661);
nand U28962 (N_28962,N_18254,N_20732);
or U28963 (N_28963,N_23559,N_19722);
nor U28964 (N_28964,N_18786,N_20045);
and U28965 (N_28965,N_23698,N_22690);
or U28966 (N_28966,N_19717,N_19516);
nand U28967 (N_28967,N_19778,N_19396);
or U28968 (N_28968,N_21022,N_20639);
and U28969 (N_28969,N_23337,N_19281);
or U28970 (N_28970,N_20845,N_18859);
nand U28971 (N_28971,N_19762,N_23634);
nand U28972 (N_28972,N_20900,N_20691);
nor U28973 (N_28973,N_21591,N_19929);
or U28974 (N_28974,N_18373,N_19709);
nor U28975 (N_28975,N_19692,N_23235);
or U28976 (N_28976,N_18191,N_19634);
xnor U28977 (N_28977,N_20828,N_20245);
and U28978 (N_28978,N_20635,N_23757);
nor U28979 (N_28979,N_23302,N_22049);
xnor U28980 (N_28980,N_21477,N_20090);
nor U28981 (N_28981,N_21739,N_22835);
or U28982 (N_28982,N_22590,N_21425);
nand U28983 (N_28983,N_19776,N_21772);
or U28984 (N_28984,N_22482,N_18894);
or U28985 (N_28985,N_21434,N_21695);
nand U28986 (N_28986,N_18073,N_21521);
nand U28987 (N_28987,N_23736,N_20038);
xnor U28988 (N_28988,N_23002,N_23319);
nor U28989 (N_28989,N_18973,N_21851);
nor U28990 (N_28990,N_23545,N_19547);
or U28991 (N_28991,N_21175,N_22903);
nor U28992 (N_28992,N_21834,N_22150);
xnor U28993 (N_28993,N_21779,N_20417);
xnor U28994 (N_28994,N_22899,N_20986);
xnor U28995 (N_28995,N_22501,N_18985);
xnor U28996 (N_28996,N_19653,N_23999);
and U28997 (N_28997,N_22350,N_21775);
nand U28998 (N_28998,N_22675,N_20243);
xor U28999 (N_28999,N_20803,N_20853);
nor U29000 (N_29000,N_18806,N_19252);
nor U29001 (N_29001,N_22718,N_22636);
and U29002 (N_29002,N_22676,N_21163);
nor U29003 (N_29003,N_19092,N_20736);
or U29004 (N_29004,N_21649,N_19475);
nor U29005 (N_29005,N_20006,N_20994);
nor U29006 (N_29006,N_19340,N_23268);
xor U29007 (N_29007,N_18919,N_22286);
nor U29008 (N_29008,N_22494,N_21247);
xor U29009 (N_29009,N_22878,N_21515);
nand U29010 (N_29010,N_22108,N_19350);
and U29011 (N_29011,N_20623,N_20968);
or U29012 (N_29012,N_23637,N_23415);
or U29013 (N_29013,N_20321,N_23258);
nand U29014 (N_29014,N_23554,N_21468);
nand U29015 (N_29015,N_20822,N_21326);
nand U29016 (N_29016,N_23557,N_23637);
nor U29017 (N_29017,N_18053,N_20290);
and U29018 (N_29018,N_18892,N_21455);
nor U29019 (N_29019,N_21122,N_20077);
and U29020 (N_29020,N_22477,N_18012);
nand U29021 (N_29021,N_21845,N_19888);
nand U29022 (N_29022,N_22304,N_20766);
or U29023 (N_29023,N_20423,N_22018);
nor U29024 (N_29024,N_23804,N_22059);
nor U29025 (N_29025,N_19529,N_18222);
and U29026 (N_29026,N_18229,N_21374);
nor U29027 (N_29027,N_23353,N_19533);
nand U29028 (N_29028,N_19467,N_20939);
or U29029 (N_29029,N_18474,N_19390);
nand U29030 (N_29030,N_23984,N_18171);
or U29031 (N_29031,N_21226,N_23500);
xor U29032 (N_29032,N_18007,N_22591);
nor U29033 (N_29033,N_23711,N_19101);
nor U29034 (N_29034,N_18991,N_20976);
xnor U29035 (N_29035,N_20398,N_19715);
xnor U29036 (N_29036,N_23431,N_20850);
and U29037 (N_29037,N_19590,N_18443);
xnor U29038 (N_29038,N_21741,N_18148);
and U29039 (N_29039,N_21927,N_18017);
xnor U29040 (N_29040,N_18620,N_18752);
nor U29041 (N_29041,N_21724,N_18174);
and U29042 (N_29042,N_22348,N_23329);
xnor U29043 (N_29043,N_21865,N_21259);
nor U29044 (N_29044,N_18274,N_19690);
nand U29045 (N_29045,N_19476,N_19623);
xnor U29046 (N_29046,N_20827,N_23432);
xor U29047 (N_29047,N_19510,N_19783);
and U29048 (N_29048,N_23010,N_21614);
and U29049 (N_29049,N_21505,N_23966);
or U29050 (N_29050,N_18237,N_18497);
xor U29051 (N_29051,N_23265,N_19496);
or U29052 (N_29052,N_20635,N_19225);
or U29053 (N_29053,N_20502,N_21057);
and U29054 (N_29054,N_19821,N_19980);
nand U29055 (N_29055,N_23730,N_23055);
or U29056 (N_29056,N_18578,N_21315);
nand U29057 (N_29057,N_18092,N_21118);
xnor U29058 (N_29058,N_22672,N_22068);
or U29059 (N_29059,N_18423,N_20357);
nor U29060 (N_29060,N_19729,N_18509);
and U29061 (N_29061,N_21666,N_18153);
xor U29062 (N_29062,N_18963,N_21099);
or U29063 (N_29063,N_21021,N_21697);
nand U29064 (N_29064,N_21953,N_18848);
and U29065 (N_29065,N_21851,N_20242);
nand U29066 (N_29066,N_23596,N_20169);
nand U29067 (N_29067,N_20277,N_18554);
nand U29068 (N_29068,N_22805,N_22964);
and U29069 (N_29069,N_18580,N_18586);
xor U29070 (N_29070,N_22020,N_18843);
or U29071 (N_29071,N_23814,N_22396);
and U29072 (N_29072,N_21023,N_22919);
nand U29073 (N_29073,N_21205,N_19739);
xor U29074 (N_29074,N_21458,N_21795);
nand U29075 (N_29075,N_23745,N_21576);
or U29076 (N_29076,N_18755,N_20669);
or U29077 (N_29077,N_20575,N_18481);
xor U29078 (N_29078,N_23606,N_21527);
and U29079 (N_29079,N_22898,N_20727);
nor U29080 (N_29080,N_18097,N_20620);
and U29081 (N_29081,N_19779,N_20637);
or U29082 (N_29082,N_22978,N_19445);
or U29083 (N_29083,N_21203,N_23400);
and U29084 (N_29084,N_21984,N_18745);
and U29085 (N_29085,N_22827,N_23866);
and U29086 (N_29086,N_18723,N_19669);
xor U29087 (N_29087,N_22511,N_21878);
or U29088 (N_29088,N_23158,N_18202);
and U29089 (N_29089,N_22756,N_22271);
and U29090 (N_29090,N_21319,N_20634);
nor U29091 (N_29091,N_23605,N_22827);
or U29092 (N_29092,N_18704,N_19821);
nor U29093 (N_29093,N_23856,N_19381);
and U29094 (N_29094,N_23728,N_19834);
nand U29095 (N_29095,N_22143,N_22506);
nor U29096 (N_29096,N_21727,N_21046);
nor U29097 (N_29097,N_19507,N_19233);
nor U29098 (N_29098,N_18585,N_23856);
and U29099 (N_29099,N_23240,N_22580);
or U29100 (N_29100,N_21942,N_18798);
nand U29101 (N_29101,N_23608,N_18230);
and U29102 (N_29102,N_18283,N_18369);
nor U29103 (N_29103,N_21206,N_20007);
or U29104 (N_29104,N_18340,N_23191);
or U29105 (N_29105,N_18217,N_19009);
nor U29106 (N_29106,N_20013,N_19712);
and U29107 (N_29107,N_22685,N_20231);
or U29108 (N_29108,N_23393,N_18472);
xor U29109 (N_29109,N_23551,N_23220);
and U29110 (N_29110,N_19000,N_23146);
nor U29111 (N_29111,N_21211,N_21833);
nor U29112 (N_29112,N_20522,N_20663);
or U29113 (N_29113,N_20300,N_19934);
nand U29114 (N_29114,N_21132,N_19912);
and U29115 (N_29115,N_22712,N_21003);
xor U29116 (N_29116,N_23573,N_18316);
nor U29117 (N_29117,N_18104,N_23108);
nor U29118 (N_29118,N_20520,N_18985);
and U29119 (N_29119,N_20489,N_23059);
and U29120 (N_29120,N_23584,N_23714);
and U29121 (N_29121,N_21977,N_23316);
nand U29122 (N_29122,N_20996,N_23714);
nor U29123 (N_29123,N_23143,N_21499);
nand U29124 (N_29124,N_19278,N_21921);
or U29125 (N_29125,N_19724,N_23820);
nand U29126 (N_29126,N_21526,N_23529);
nand U29127 (N_29127,N_22228,N_22283);
and U29128 (N_29128,N_20723,N_23097);
nand U29129 (N_29129,N_20197,N_19774);
and U29130 (N_29130,N_22012,N_21353);
xnor U29131 (N_29131,N_19316,N_18287);
nor U29132 (N_29132,N_22106,N_18203);
or U29133 (N_29133,N_22593,N_18708);
nand U29134 (N_29134,N_21152,N_23524);
nand U29135 (N_29135,N_23346,N_19206);
or U29136 (N_29136,N_19967,N_19371);
nor U29137 (N_29137,N_22874,N_22776);
or U29138 (N_29138,N_19597,N_22006);
or U29139 (N_29139,N_20861,N_18141);
or U29140 (N_29140,N_20185,N_19044);
nor U29141 (N_29141,N_19921,N_18796);
or U29142 (N_29142,N_22690,N_21816);
or U29143 (N_29143,N_22449,N_19968);
xnor U29144 (N_29144,N_19518,N_23395);
and U29145 (N_29145,N_18349,N_21840);
xnor U29146 (N_29146,N_21409,N_23949);
xor U29147 (N_29147,N_22660,N_22013);
or U29148 (N_29148,N_19159,N_18126);
nand U29149 (N_29149,N_23530,N_23884);
or U29150 (N_29150,N_22750,N_21790);
and U29151 (N_29151,N_21991,N_22331);
or U29152 (N_29152,N_22747,N_18245);
nand U29153 (N_29153,N_18379,N_18156);
xnor U29154 (N_29154,N_21975,N_19506);
nand U29155 (N_29155,N_20571,N_22814);
nand U29156 (N_29156,N_23594,N_21101);
nor U29157 (N_29157,N_22710,N_19397);
nand U29158 (N_29158,N_23824,N_20957);
or U29159 (N_29159,N_21407,N_20911);
and U29160 (N_29160,N_19034,N_22800);
nor U29161 (N_29161,N_22055,N_22212);
and U29162 (N_29162,N_20280,N_19007);
nor U29163 (N_29163,N_22483,N_23151);
nand U29164 (N_29164,N_23675,N_20172);
xor U29165 (N_29165,N_22019,N_21950);
xor U29166 (N_29166,N_21182,N_18512);
nand U29167 (N_29167,N_23603,N_21494);
and U29168 (N_29168,N_20100,N_18784);
or U29169 (N_29169,N_22133,N_18323);
nand U29170 (N_29170,N_22869,N_23207);
or U29171 (N_29171,N_23142,N_22241);
nor U29172 (N_29172,N_18013,N_18882);
nor U29173 (N_29173,N_18199,N_20867);
nor U29174 (N_29174,N_20872,N_18845);
or U29175 (N_29175,N_18445,N_20112);
xor U29176 (N_29176,N_20953,N_23588);
or U29177 (N_29177,N_20126,N_19758);
xnor U29178 (N_29178,N_18100,N_23993);
nand U29179 (N_29179,N_19057,N_22330);
and U29180 (N_29180,N_22374,N_22208);
nand U29181 (N_29181,N_20821,N_23681);
or U29182 (N_29182,N_20997,N_19096);
xor U29183 (N_29183,N_18148,N_19645);
xnor U29184 (N_29184,N_22737,N_21034);
nor U29185 (N_29185,N_18179,N_21750);
nand U29186 (N_29186,N_23583,N_22241);
nand U29187 (N_29187,N_18055,N_19040);
xor U29188 (N_29188,N_20910,N_19532);
nand U29189 (N_29189,N_18790,N_20270);
or U29190 (N_29190,N_20417,N_18049);
or U29191 (N_29191,N_23972,N_20281);
nand U29192 (N_29192,N_21100,N_22359);
and U29193 (N_29193,N_21372,N_21180);
or U29194 (N_29194,N_21822,N_19681);
xnor U29195 (N_29195,N_19882,N_19875);
xor U29196 (N_29196,N_23635,N_22236);
nand U29197 (N_29197,N_21152,N_21010);
nor U29198 (N_29198,N_23901,N_19023);
xor U29199 (N_29199,N_19662,N_22141);
xor U29200 (N_29200,N_18309,N_23283);
nand U29201 (N_29201,N_22956,N_18896);
nand U29202 (N_29202,N_19157,N_23842);
nand U29203 (N_29203,N_21320,N_19812);
and U29204 (N_29204,N_20748,N_20117);
and U29205 (N_29205,N_23409,N_18822);
nand U29206 (N_29206,N_21265,N_20235);
xor U29207 (N_29207,N_18697,N_21117);
nor U29208 (N_29208,N_18158,N_18104);
and U29209 (N_29209,N_21140,N_20893);
nor U29210 (N_29210,N_21921,N_21530);
nand U29211 (N_29211,N_20003,N_23546);
and U29212 (N_29212,N_20199,N_22614);
or U29213 (N_29213,N_21182,N_18509);
nand U29214 (N_29214,N_19742,N_20545);
or U29215 (N_29215,N_21125,N_21079);
xnor U29216 (N_29216,N_20859,N_23752);
nor U29217 (N_29217,N_21239,N_19170);
xor U29218 (N_29218,N_23018,N_21285);
or U29219 (N_29219,N_20023,N_20939);
nand U29220 (N_29220,N_23365,N_23196);
nand U29221 (N_29221,N_20089,N_21584);
nor U29222 (N_29222,N_23418,N_22826);
or U29223 (N_29223,N_21312,N_22703);
nand U29224 (N_29224,N_22443,N_18405);
or U29225 (N_29225,N_19974,N_18969);
and U29226 (N_29226,N_19973,N_21191);
xnor U29227 (N_29227,N_19076,N_21433);
xnor U29228 (N_29228,N_21683,N_19001);
nor U29229 (N_29229,N_23207,N_23386);
or U29230 (N_29230,N_21748,N_18544);
and U29231 (N_29231,N_23705,N_20632);
and U29232 (N_29232,N_20610,N_18266);
nand U29233 (N_29233,N_22421,N_21148);
nand U29234 (N_29234,N_20031,N_22648);
xor U29235 (N_29235,N_20588,N_23567);
nand U29236 (N_29236,N_19830,N_19576);
or U29237 (N_29237,N_20074,N_19754);
or U29238 (N_29238,N_20133,N_21968);
and U29239 (N_29239,N_20711,N_21289);
and U29240 (N_29240,N_19954,N_20721);
and U29241 (N_29241,N_19009,N_23844);
nand U29242 (N_29242,N_18963,N_22424);
or U29243 (N_29243,N_18138,N_23334);
xor U29244 (N_29244,N_21571,N_21564);
and U29245 (N_29245,N_19904,N_22455);
or U29246 (N_29246,N_23149,N_19206);
xor U29247 (N_29247,N_19921,N_21365);
nand U29248 (N_29248,N_21185,N_21461);
or U29249 (N_29249,N_18111,N_22113);
or U29250 (N_29250,N_18306,N_18462);
nand U29251 (N_29251,N_21708,N_19051);
xor U29252 (N_29252,N_20886,N_22188);
nand U29253 (N_29253,N_18706,N_18149);
nor U29254 (N_29254,N_21619,N_21981);
or U29255 (N_29255,N_21229,N_20992);
nand U29256 (N_29256,N_20458,N_19896);
xnor U29257 (N_29257,N_19737,N_18124);
nor U29258 (N_29258,N_22667,N_22067);
or U29259 (N_29259,N_22678,N_21199);
xor U29260 (N_29260,N_23361,N_18381);
or U29261 (N_29261,N_22810,N_22728);
and U29262 (N_29262,N_23754,N_20861);
xor U29263 (N_29263,N_21369,N_18763);
nor U29264 (N_29264,N_23305,N_23496);
or U29265 (N_29265,N_23137,N_20256);
or U29266 (N_29266,N_23435,N_21486);
and U29267 (N_29267,N_18476,N_21313);
xnor U29268 (N_29268,N_21934,N_22855);
xnor U29269 (N_29269,N_20200,N_22055);
nand U29270 (N_29270,N_19533,N_22195);
or U29271 (N_29271,N_20139,N_19939);
xnor U29272 (N_29272,N_18319,N_18092);
nand U29273 (N_29273,N_20556,N_18995);
nand U29274 (N_29274,N_22541,N_18770);
and U29275 (N_29275,N_20333,N_22380);
xnor U29276 (N_29276,N_18599,N_23666);
xnor U29277 (N_29277,N_21852,N_21419);
nor U29278 (N_29278,N_23821,N_22848);
or U29279 (N_29279,N_21193,N_21130);
xnor U29280 (N_29280,N_22624,N_18394);
nor U29281 (N_29281,N_20547,N_20171);
nand U29282 (N_29282,N_20911,N_22265);
or U29283 (N_29283,N_22905,N_18009);
and U29284 (N_29284,N_21274,N_22291);
nand U29285 (N_29285,N_18754,N_20903);
and U29286 (N_29286,N_22879,N_21962);
nor U29287 (N_29287,N_21696,N_19484);
xor U29288 (N_29288,N_21769,N_19279);
xor U29289 (N_29289,N_19591,N_22621);
and U29290 (N_29290,N_21731,N_21621);
xor U29291 (N_29291,N_19051,N_19356);
xnor U29292 (N_29292,N_19125,N_18477);
nand U29293 (N_29293,N_23029,N_23839);
or U29294 (N_29294,N_22985,N_19505);
nand U29295 (N_29295,N_23183,N_20249);
xor U29296 (N_29296,N_20755,N_20336);
or U29297 (N_29297,N_18553,N_18204);
xor U29298 (N_29298,N_20962,N_21899);
xnor U29299 (N_29299,N_18111,N_23428);
or U29300 (N_29300,N_23967,N_23554);
and U29301 (N_29301,N_23253,N_22127);
or U29302 (N_29302,N_23318,N_23821);
and U29303 (N_29303,N_21020,N_22164);
nand U29304 (N_29304,N_20686,N_18584);
nor U29305 (N_29305,N_22850,N_20283);
or U29306 (N_29306,N_22704,N_22717);
xor U29307 (N_29307,N_22883,N_20050);
nor U29308 (N_29308,N_18111,N_18625);
nand U29309 (N_29309,N_20936,N_21145);
xor U29310 (N_29310,N_23948,N_20037);
and U29311 (N_29311,N_20205,N_19612);
and U29312 (N_29312,N_18995,N_20987);
nand U29313 (N_29313,N_21574,N_18441);
and U29314 (N_29314,N_21909,N_19577);
xor U29315 (N_29315,N_18866,N_23420);
xor U29316 (N_29316,N_18077,N_18797);
nand U29317 (N_29317,N_21627,N_20774);
nand U29318 (N_29318,N_19560,N_23201);
xnor U29319 (N_29319,N_18557,N_19505);
or U29320 (N_29320,N_21773,N_18226);
xnor U29321 (N_29321,N_19990,N_21718);
nand U29322 (N_29322,N_20740,N_19455);
nor U29323 (N_29323,N_19316,N_20798);
nand U29324 (N_29324,N_20122,N_21306);
nor U29325 (N_29325,N_22372,N_22921);
and U29326 (N_29326,N_21949,N_21627);
nor U29327 (N_29327,N_21692,N_19996);
nand U29328 (N_29328,N_21470,N_20176);
and U29329 (N_29329,N_23834,N_19171);
xor U29330 (N_29330,N_21435,N_19556);
nor U29331 (N_29331,N_21664,N_23733);
nand U29332 (N_29332,N_21134,N_19966);
nand U29333 (N_29333,N_23883,N_20514);
xor U29334 (N_29334,N_21352,N_23178);
or U29335 (N_29335,N_18728,N_21071);
xor U29336 (N_29336,N_23497,N_20724);
or U29337 (N_29337,N_18228,N_21064);
xor U29338 (N_29338,N_18117,N_19869);
or U29339 (N_29339,N_22914,N_21652);
nand U29340 (N_29340,N_21513,N_18473);
nand U29341 (N_29341,N_22577,N_18998);
nor U29342 (N_29342,N_22222,N_18307);
xnor U29343 (N_29343,N_19946,N_20456);
or U29344 (N_29344,N_18834,N_20957);
or U29345 (N_29345,N_19893,N_18357);
nand U29346 (N_29346,N_22541,N_23027);
xnor U29347 (N_29347,N_18792,N_18532);
nand U29348 (N_29348,N_23309,N_21560);
nand U29349 (N_29349,N_20171,N_20787);
nand U29350 (N_29350,N_22352,N_19925);
xnor U29351 (N_29351,N_19042,N_22880);
nor U29352 (N_29352,N_20526,N_21419);
and U29353 (N_29353,N_23382,N_23679);
xnor U29354 (N_29354,N_23378,N_18289);
and U29355 (N_29355,N_21290,N_18788);
xnor U29356 (N_29356,N_23289,N_23850);
nand U29357 (N_29357,N_20469,N_19639);
and U29358 (N_29358,N_19237,N_19362);
nor U29359 (N_29359,N_20090,N_19719);
and U29360 (N_29360,N_21084,N_21563);
or U29361 (N_29361,N_19645,N_22854);
xor U29362 (N_29362,N_18431,N_19431);
nor U29363 (N_29363,N_21817,N_19131);
and U29364 (N_29364,N_20964,N_18389);
or U29365 (N_29365,N_20810,N_20260);
xor U29366 (N_29366,N_22543,N_21754);
or U29367 (N_29367,N_22797,N_20924);
nor U29368 (N_29368,N_22211,N_23049);
or U29369 (N_29369,N_18991,N_22238);
xor U29370 (N_29370,N_22282,N_22858);
nand U29371 (N_29371,N_20285,N_22378);
or U29372 (N_29372,N_18645,N_19785);
nand U29373 (N_29373,N_18023,N_21925);
xor U29374 (N_29374,N_20376,N_21003);
nor U29375 (N_29375,N_23042,N_18520);
nor U29376 (N_29376,N_23348,N_22164);
nand U29377 (N_29377,N_19394,N_20740);
and U29378 (N_29378,N_21223,N_22482);
or U29379 (N_29379,N_23082,N_22728);
nor U29380 (N_29380,N_19719,N_23041);
and U29381 (N_29381,N_23565,N_23423);
nand U29382 (N_29382,N_22731,N_20719);
xnor U29383 (N_29383,N_19704,N_22344);
or U29384 (N_29384,N_23316,N_20056);
nand U29385 (N_29385,N_22642,N_22503);
and U29386 (N_29386,N_20151,N_20939);
xor U29387 (N_29387,N_22016,N_23154);
or U29388 (N_29388,N_19162,N_21921);
xor U29389 (N_29389,N_21358,N_20567);
or U29390 (N_29390,N_18570,N_22544);
nand U29391 (N_29391,N_20578,N_20839);
or U29392 (N_29392,N_20890,N_22897);
nor U29393 (N_29393,N_21603,N_20322);
xnor U29394 (N_29394,N_23527,N_20646);
nor U29395 (N_29395,N_20645,N_18124);
or U29396 (N_29396,N_18712,N_21573);
or U29397 (N_29397,N_18887,N_20992);
or U29398 (N_29398,N_18927,N_19880);
nand U29399 (N_29399,N_20239,N_19026);
or U29400 (N_29400,N_23779,N_18989);
and U29401 (N_29401,N_22567,N_19453);
xnor U29402 (N_29402,N_18378,N_19610);
nor U29403 (N_29403,N_20762,N_20748);
xnor U29404 (N_29404,N_18822,N_22070);
xnor U29405 (N_29405,N_20487,N_21821);
nand U29406 (N_29406,N_19208,N_20084);
nor U29407 (N_29407,N_22936,N_22470);
nand U29408 (N_29408,N_21872,N_23015);
nand U29409 (N_29409,N_23816,N_19199);
xnor U29410 (N_29410,N_23870,N_23619);
xor U29411 (N_29411,N_22615,N_18578);
and U29412 (N_29412,N_18719,N_21848);
nor U29413 (N_29413,N_19490,N_21626);
nand U29414 (N_29414,N_20176,N_22346);
nand U29415 (N_29415,N_20360,N_19938);
xnor U29416 (N_29416,N_21326,N_22398);
and U29417 (N_29417,N_21448,N_20263);
nand U29418 (N_29418,N_23279,N_20222);
nor U29419 (N_29419,N_19033,N_22494);
xor U29420 (N_29420,N_21565,N_20388);
nand U29421 (N_29421,N_21692,N_23249);
or U29422 (N_29422,N_23734,N_21177);
nor U29423 (N_29423,N_19791,N_20829);
nand U29424 (N_29424,N_19045,N_18016);
and U29425 (N_29425,N_20147,N_18649);
or U29426 (N_29426,N_19925,N_20130);
nor U29427 (N_29427,N_20171,N_20424);
nor U29428 (N_29428,N_19104,N_23236);
and U29429 (N_29429,N_21384,N_23806);
nand U29430 (N_29430,N_22274,N_19896);
or U29431 (N_29431,N_23764,N_21288);
and U29432 (N_29432,N_20516,N_22726);
or U29433 (N_29433,N_19946,N_18886);
xnor U29434 (N_29434,N_22416,N_20931);
and U29435 (N_29435,N_21113,N_19229);
xnor U29436 (N_29436,N_21602,N_22084);
and U29437 (N_29437,N_18095,N_23758);
xor U29438 (N_29438,N_20598,N_18296);
or U29439 (N_29439,N_18702,N_19346);
nand U29440 (N_29440,N_19281,N_20768);
and U29441 (N_29441,N_19337,N_21068);
or U29442 (N_29442,N_22211,N_18856);
nand U29443 (N_29443,N_18922,N_23510);
nor U29444 (N_29444,N_21091,N_23506);
nand U29445 (N_29445,N_20722,N_23689);
nor U29446 (N_29446,N_22055,N_23992);
nand U29447 (N_29447,N_20984,N_22268);
and U29448 (N_29448,N_23714,N_22493);
and U29449 (N_29449,N_21806,N_23543);
xnor U29450 (N_29450,N_23529,N_22595);
nor U29451 (N_29451,N_20350,N_19928);
or U29452 (N_29452,N_20506,N_19605);
nand U29453 (N_29453,N_21610,N_19774);
xor U29454 (N_29454,N_22137,N_23322);
xnor U29455 (N_29455,N_21646,N_23684);
xor U29456 (N_29456,N_18854,N_20752);
nand U29457 (N_29457,N_22168,N_20933);
nand U29458 (N_29458,N_21170,N_21664);
and U29459 (N_29459,N_20883,N_21057);
or U29460 (N_29460,N_23603,N_22612);
and U29461 (N_29461,N_22423,N_21129);
or U29462 (N_29462,N_18444,N_20571);
nor U29463 (N_29463,N_18826,N_23931);
nand U29464 (N_29464,N_19712,N_20391);
nand U29465 (N_29465,N_18922,N_23067);
or U29466 (N_29466,N_22756,N_22093);
or U29467 (N_29467,N_22828,N_22163);
nand U29468 (N_29468,N_22716,N_22116);
xnor U29469 (N_29469,N_19236,N_19762);
nor U29470 (N_29470,N_22671,N_23174);
nor U29471 (N_29471,N_23462,N_23408);
nand U29472 (N_29472,N_20797,N_22589);
nor U29473 (N_29473,N_20324,N_22009);
xor U29474 (N_29474,N_19844,N_19724);
nand U29475 (N_29475,N_23817,N_19660);
nand U29476 (N_29476,N_19736,N_19461);
nor U29477 (N_29477,N_20622,N_22275);
xnor U29478 (N_29478,N_19261,N_18497);
or U29479 (N_29479,N_21364,N_20464);
xnor U29480 (N_29480,N_23200,N_23816);
xnor U29481 (N_29481,N_19900,N_23520);
nand U29482 (N_29482,N_19229,N_19177);
nor U29483 (N_29483,N_20625,N_19876);
or U29484 (N_29484,N_20388,N_22851);
and U29485 (N_29485,N_20322,N_22306);
xnor U29486 (N_29486,N_22733,N_21279);
nor U29487 (N_29487,N_18223,N_23898);
nand U29488 (N_29488,N_22264,N_22432);
or U29489 (N_29489,N_18934,N_18220);
nor U29490 (N_29490,N_23263,N_23241);
nor U29491 (N_29491,N_23203,N_19376);
and U29492 (N_29492,N_21328,N_18846);
nor U29493 (N_29493,N_20566,N_22935);
and U29494 (N_29494,N_23445,N_19934);
nand U29495 (N_29495,N_19710,N_21759);
or U29496 (N_29496,N_21909,N_22532);
xnor U29497 (N_29497,N_19866,N_22051);
nand U29498 (N_29498,N_21980,N_21828);
nand U29499 (N_29499,N_22371,N_20180);
nand U29500 (N_29500,N_18149,N_18174);
xnor U29501 (N_29501,N_20070,N_23179);
or U29502 (N_29502,N_23012,N_21856);
xnor U29503 (N_29503,N_22800,N_21425);
and U29504 (N_29504,N_20127,N_19720);
xor U29505 (N_29505,N_21335,N_22080);
nand U29506 (N_29506,N_19699,N_18650);
nand U29507 (N_29507,N_20037,N_19678);
xor U29508 (N_29508,N_20118,N_21690);
and U29509 (N_29509,N_19903,N_22112);
and U29510 (N_29510,N_18598,N_20671);
or U29511 (N_29511,N_19686,N_23965);
nand U29512 (N_29512,N_18951,N_22338);
nand U29513 (N_29513,N_19299,N_21164);
or U29514 (N_29514,N_19495,N_20522);
and U29515 (N_29515,N_23901,N_20758);
nand U29516 (N_29516,N_18194,N_23263);
and U29517 (N_29517,N_21293,N_21104);
and U29518 (N_29518,N_19469,N_18517);
nor U29519 (N_29519,N_18388,N_19770);
nand U29520 (N_29520,N_21458,N_19691);
or U29521 (N_29521,N_20657,N_22969);
nand U29522 (N_29522,N_22610,N_18220);
xor U29523 (N_29523,N_21944,N_20350);
or U29524 (N_29524,N_20620,N_23601);
and U29525 (N_29525,N_18109,N_23733);
nand U29526 (N_29526,N_18312,N_19023);
xor U29527 (N_29527,N_18707,N_23848);
or U29528 (N_29528,N_22529,N_23438);
nor U29529 (N_29529,N_19781,N_21624);
and U29530 (N_29530,N_22696,N_22022);
xnor U29531 (N_29531,N_23517,N_22789);
or U29532 (N_29532,N_18728,N_20270);
nor U29533 (N_29533,N_21688,N_19161);
or U29534 (N_29534,N_23135,N_22255);
and U29535 (N_29535,N_21649,N_22681);
nor U29536 (N_29536,N_20052,N_22812);
or U29537 (N_29537,N_19837,N_22688);
or U29538 (N_29538,N_22846,N_20213);
and U29539 (N_29539,N_20494,N_22609);
or U29540 (N_29540,N_23734,N_20721);
and U29541 (N_29541,N_20350,N_21850);
xor U29542 (N_29542,N_19206,N_20718);
nor U29543 (N_29543,N_22074,N_20850);
and U29544 (N_29544,N_22187,N_18923);
xor U29545 (N_29545,N_20271,N_21864);
nor U29546 (N_29546,N_18877,N_21747);
nand U29547 (N_29547,N_19873,N_19564);
xor U29548 (N_29548,N_23548,N_22229);
nand U29549 (N_29549,N_21918,N_18010);
xnor U29550 (N_29550,N_21472,N_19725);
and U29551 (N_29551,N_23641,N_23839);
and U29552 (N_29552,N_19681,N_21113);
or U29553 (N_29553,N_18538,N_22237);
or U29554 (N_29554,N_19911,N_22773);
or U29555 (N_29555,N_23374,N_21987);
or U29556 (N_29556,N_19152,N_23094);
or U29557 (N_29557,N_19476,N_22570);
and U29558 (N_29558,N_20824,N_22425);
nor U29559 (N_29559,N_21630,N_18134);
xnor U29560 (N_29560,N_21180,N_18365);
nand U29561 (N_29561,N_18602,N_20479);
nand U29562 (N_29562,N_23893,N_23040);
or U29563 (N_29563,N_19517,N_21914);
nor U29564 (N_29564,N_20225,N_22467);
nand U29565 (N_29565,N_20544,N_18425);
nor U29566 (N_29566,N_23310,N_21110);
nor U29567 (N_29567,N_23811,N_21550);
or U29568 (N_29568,N_21807,N_22118);
xnor U29569 (N_29569,N_22995,N_21040);
nand U29570 (N_29570,N_22135,N_19220);
and U29571 (N_29571,N_23726,N_21735);
and U29572 (N_29572,N_18519,N_18810);
nor U29573 (N_29573,N_22855,N_20989);
nor U29574 (N_29574,N_23830,N_23312);
or U29575 (N_29575,N_19872,N_19169);
nand U29576 (N_29576,N_20773,N_19755);
xor U29577 (N_29577,N_23323,N_18426);
and U29578 (N_29578,N_19535,N_20112);
or U29579 (N_29579,N_18282,N_22351);
or U29580 (N_29580,N_20797,N_22279);
and U29581 (N_29581,N_23526,N_22786);
or U29582 (N_29582,N_19076,N_18022);
nand U29583 (N_29583,N_23949,N_23033);
or U29584 (N_29584,N_21322,N_18201);
or U29585 (N_29585,N_20011,N_22577);
nand U29586 (N_29586,N_22975,N_23111);
or U29587 (N_29587,N_20008,N_19889);
and U29588 (N_29588,N_20174,N_19678);
or U29589 (N_29589,N_23667,N_23453);
or U29590 (N_29590,N_18509,N_18931);
xnor U29591 (N_29591,N_18306,N_23174);
nand U29592 (N_29592,N_20197,N_20823);
nor U29593 (N_29593,N_21807,N_18339);
or U29594 (N_29594,N_20699,N_18162);
or U29595 (N_29595,N_22749,N_20242);
nand U29596 (N_29596,N_21720,N_23047);
and U29597 (N_29597,N_21638,N_21243);
nand U29598 (N_29598,N_20025,N_22327);
xnor U29599 (N_29599,N_19226,N_22348);
nand U29600 (N_29600,N_18693,N_23409);
xnor U29601 (N_29601,N_22359,N_22238);
or U29602 (N_29602,N_23051,N_23767);
or U29603 (N_29603,N_22196,N_19605);
and U29604 (N_29604,N_19176,N_20863);
or U29605 (N_29605,N_21855,N_20091);
and U29606 (N_29606,N_21944,N_21400);
and U29607 (N_29607,N_21485,N_18411);
or U29608 (N_29608,N_20496,N_22676);
and U29609 (N_29609,N_23672,N_19328);
nor U29610 (N_29610,N_21796,N_22555);
or U29611 (N_29611,N_22744,N_20889);
or U29612 (N_29612,N_18106,N_22762);
or U29613 (N_29613,N_22913,N_18330);
xor U29614 (N_29614,N_19364,N_22963);
nand U29615 (N_29615,N_19243,N_18154);
nand U29616 (N_29616,N_18663,N_19603);
nand U29617 (N_29617,N_21764,N_22133);
xor U29618 (N_29618,N_21221,N_18066);
xnor U29619 (N_29619,N_23583,N_20018);
nor U29620 (N_29620,N_18409,N_22783);
or U29621 (N_29621,N_19498,N_20271);
and U29622 (N_29622,N_20817,N_19985);
or U29623 (N_29623,N_18469,N_23568);
and U29624 (N_29624,N_18510,N_20531);
xnor U29625 (N_29625,N_18334,N_18518);
or U29626 (N_29626,N_18277,N_21362);
nand U29627 (N_29627,N_19200,N_20499);
nor U29628 (N_29628,N_18640,N_19457);
xnor U29629 (N_29629,N_23166,N_22327);
and U29630 (N_29630,N_19101,N_19404);
or U29631 (N_29631,N_20806,N_22057);
nor U29632 (N_29632,N_20177,N_19773);
nor U29633 (N_29633,N_22203,N_21966);
xor U29634 (N_29634,N_20010,N_22082);
or U29635 (N_29635,N_19099,N_19864);
xnor U29636 (N_29636,N_23407,N_22570);
xnor U29637 (N_29637,N_22198,N_18059);
nor U29638 (N_29638,N_22920,N_23236);
and U29639 (N_29639,N_20896,N_19499);
nand U29640 (N_29640,N_23542,N_23118);
nor U29641 (N_29641,N_19695,N_21370);
nor U29642 (N_29642,N_23136,N_21067);
nand U29643 (N_29643,N_21312,N_19834);
or U29644 (N_29644,N_22482,N_22789);
nor U29645 (N_29645,N_18869,N_22774);
xnor U29646 (N_29646,N_20250,N_23287);
or U29647 (N_29647,N_18533,N_23068);
or U29648 (N_29648,N_23617,N_20082);
nand U29649 (N_29649,N_22580,N_23977);
and U29650 (N_29650,N_20122,N_19111);
xnor U29651 (N_29651,N_18498,N_22421);
nand U29652 (N_29652,N_22454,N_20507);
or U29653 (N_29653,N_19846,N_22936);
xor U29654 (N_29654,N_19397,N_21962);
nand U29655 (N_29655,N_19365,N_18130);
or U29656 (N_29656,N_20377,N_19716);
nor U29657 (N_29657,N_22290,N_20070);
xor U29658 (N_29658,N_19788,N_19406);
nor U29659 (N_29659,N_21162,N_18341);
or U29660 (N_29660,N_21828,N_19777);
nand U29661 (N_29661,N_22102,N_21105);
nand U29662 (N_29662,N_22168,N_19337);
nand U29663 (N_29663,N_21647,N_18051);
xnor U29664 (N_29664,N_20579,N_19862);
and U29665 (N_29665,N_22066,N_23837);
or U29666 (N_29666,N_22513,N_21302);
xor U29667 (N_29667,N_20959,N_22683);
nand U29668 (N_29668,N_21306,N_18945);
nand U29669 (N_29669,N_23799,N_21893);
nand U29670 (N_29670,N_23270,N_18142);
xor U29671 (N_29671,N_18395,N_22636);
or U29672 (N_29672,N_22721,N_22825);
xor U29673 (N_29673,N_18080,N_21581);
xnor U29674 (N_29674,N_21223,N_20697);
or U29675 (N_29675,N_19756,N_23491);
xnor U29676 (N_29676,N_19728,N_18169);
and U29677 (N_29677,N_22218,N_23847);
nor U29678 (N_29678,N_22407,N_19589);
nand U29679 (N_29679,N_18997,N_19292);
nor U29680 (N_29680,N_22156,N_23318);
nor U29681 (N_29681,N_20350,N_22591);
xnor U29682 (N_29682,N_21061,N_22722);
xnor U29683 (N_29683,N_20318,N_20595);
and U29684 (N_29684,N_20221,N_18414);
and U29685 (N_29685,N_20205,N_23654);
or U29686 (N_29686,N_22259,N_20679);
or U29687 (N_29687,N_23965,N_19057);
and U29688 (N_29688,N_19147,N_20155);
or U29689 (N_29689,N_20812,N_23133);
or U29690 (N_29690,N_23507,N_20811);
nand U29691 (N_29691,N_23607,N_20876);
nand U29692 (N_29692,N_20703,N_22686);
nor U29693 (N_29693,N_20486,N_20787);
nor U29694 (N_29694,N_21404,N_21215);
or U29695 (N_29695,N_18075,N_21928);
nor U29696 (N_29696,N_23549,N_21475);
or U29697 (N_29697,N_20077,N_22760);
and U29698 (N_29698,N_21947,N_20783);
xnor U29699 (N_29699,N_20260,N_21982);
and U29700 (N_29700,N_19200,N_22447);
nor U29701 (N_29701,N_18483,N_23505);
nand U29702 (N_29702,N_18392,N_23341);
xnor U29703 (N_29703,N_18278,N_18018);
nor U29704 (N_29704,N_21439,N_22506);
and U29705 (N_29705,N_22664,N_23984);
or U29706 (N_29706,N_18828,N_23140);
nor U29707 (N_29707,N_18943,N_23742);
xnor U29708 (N_29708,N_23638,N_20068);
xnor U29709 (N_29709,N_18416,N_21166);
nor U29710 (N_29710,N_23938,N_20751);
or U29711 (N_29711,N_23635,N_18412);
nand U29712 (N_29712,N_18448,N_22746);
and U29713 (N_29713,N_18295,N_23958);
nor U29714 (N_29714,N_19180,N_20651);
and U29715 (N_29715,N_21672,N_19634);
xor U29716 (N_29716,N_23729,N_18323);
nor U29717 (N_29717,N_19328,N_18905);
nor U29718 (N_29718,N_23825,N_18217);
xnor U29719 (N_29719,N_23865,N_19184);
and U29720 (N_29720,N_20363,N_20486);
nor U29721 (N_29721,N_22356,N_21548);
nand U29722 (N_29722,N_18005,N_20346);
nand U29723 (N_29723,N_19336,N_18993);
and U29724 (N_29724,N_23207,N_20501);
or U29725 (N_29725,N_20066,N_19945);
nand U29726 (N_29726,N_22665,N_18172);
nor U29727 (N_29727,N_22958,N_23385);
nand U29728 (N_29728,N_19229,N_19999);
nand U29729 (N_29729,N_18942,N_21421);
xor U29730 (N_29730,N_23406,N_22432);
or U29731 (N_29731,N_22568,N_22746);
and U29732 (N_29732,N_23397,N_21952);
nand U29733 (N_29733,N_21155,N_21142);
nand U29734 (N_29734,N_20752,N_19782);
nor U29735 (N_29735,N_20133,N_21909);
nand U29736 (N_29736,N_23028,N_22568);
and U29737 (N_29737,N_21070,N_23561);
or U29738 (N_29738,N_19958,N_22823);
or U29739 (N_29739,N_23941,N_19614);
xor U29740 (N_29740,N_22850,N_20145);
xnor U29741 (N_29741,N_19153,N_21060);
nand U29742 (N_29742,N_19796,N_22033);
nor U29743 (N_29743,N_23802,N_21807);
nor U29744 (N_29744,N_19052,N_22063);
or U29745 (N_29745,N_19146,N_18837);
nand U29746 (N_29746,N_18395,N_20881);
or U29747 (N_29747,N_21021,N_18485);
nand U29748 (N_29748,N_21669,N_23822);
nand U29749 (N_29749,N_19728,N_20518);
nor U29750 (N_29750,N_21592,N_21335);
nor U29751 (N_29751,N_20103,N_18229);
xnor U29752 (N_29752,N_18809,N_19087);
or U29753 (N_29753,N_20934,N_22020);
or U29754 (N_29754,N_22201,N_22775);
nand U29755 (N_29755,N_19511,N_19488);
xor U29756 (N_29756,N_18719,N_19232);
nor U29757 (N_29757,N_20488,N_19652);
nor U29758 (N_29758,N_22386,N_20880);
and U29759 (N_29759,N_23161,N_19793);
nor U29760 (N_29760,N_19560,N_21287);
xor U29761 (N_29761,N_18132,N_19258);
nor U29762 (N_29762,N_18072,N_21657);
xnor U29763 (N_29763,N_23850,N_23288);
nand U29764 (N_29764,N_21243,N_23388);
xor U29765 (N_29765,N_19200,N_19606);
xnor U29766 (N_29766,N_21766,N_21254);
xor U29767 (N_29767,N_20729,N_18219);
nor U29768 (N_29768,N_19031,N_21038);
and U29769 (N_29769,N_22397,N_19596);
nor U29770 (N_29770,N_23829,N_22020);
or U29771 (N_29771,N_20172,N_19916);
and U29772 (N_29772,N_20719,N_22262);
xnor U29773 (N_29773,N_20746,N_21974);
xnor U29774 (N_29774,N_22012,N_20292);
xnor U29775 (N_29775,N_20066,N_19287);
nand U29776 (N_29776,N_18993,N_23763);
and U29777 (N_29777,N_21580,N_22175);
nand U29778 (N_29778,N_20834,N_23139);
or U29779 (N_29779,N_18033,N_22352);
or U29780 (N_29780,N_21790,N_19946);
xnor U29781 (N_29781,N_19039,N_21687);
or U29782 (N_29782,N_18972,N_20172);
nand U29783 (N_29783,N_21450,N_19308);
or U29784 (N_29784,N_22384,N_18849);
or U29785 (N_29785,N_21566,N_23612);
nand U29786 (N_29786,N_23760,N_20913);
xnor U29787 (N_29787,N_21932,N_18222);
or U29788 (N_29788,N_18375,N_23737);
xnor U29789 (N_29789,N_20857,N_22430);
and U29790 (N_29790,N_20103,N_23275);
and U29791 (N_29791,N_19933,N_20907);
xnor U29792 (N_29792,N_19259,N_23832);
nor U29793 (N_29793,N_19268,N_22202);
nor U29794 (N_29794,N_18332,N_18279);
xnor U29795 (N_29795,N_23538,N_18231);
and U29796 (N_29796,N_20763,N_23960);
xor U29797 (N_29797,N_21465,N_21298);
and U29798 (N_29798,N_19216,N_18055);
or U29799 (N_29799,N_20846,N_21036);
nand U29800 (N_29800,N_18623,N_23661);
nand U29801 (N_29801,N_22596,N_18037);
or U29802 (N_29802,N_21948,N_21899);
nor U29803 (N_29803,N_20894,N_22745);
nor U29804 (N_29804,N_20583,N_23617);
nand U29805 (N_29805,N_23947,N_23117);
or U29806 (N_29806,N_19582,N_19120);
xnor U29807 (N_29807,N_18624,N_21730);
nand U29808 (N_29808,N_22547,N_21939);
or U29809 (N_29809,N_23392,N_22313);
xnor U29810 (N_29810,N_19889,N_18342);
nor U29811 (N_29811,N_20867,N_22542);
xor U29812 (N_29812,N_21309,N_18301);
nand U29813 (N_29813,N_22859,N_19084);
nor U29814 (N_29814,N_18950,N_23510);
nor U29815 (N_29815,N_22208,N_22579);
and U29816 (N_29816,N_18636,N_19912);
and U29817 (N_29817,N_22233,N_19862);
and U29818 (N_29818,N_19098,N_20174);
or U29819 (N_29819,N_18404,N_22788);
nand U29820 (N_29820,N_22578,N_18769);
and U29821 (N_29821,N_23033,N_20315);
or U29822 (N_29822,N_23574,N_21466);
nand U29823 (N_29823,N_23092,N_23970);
and U29824 (N_29824,N_20517,N_22105);
nor U29825 (N_29825,N_20169,N_22313);
or U29826 (N_29826,N_23038,N_19787);
nor U29827 (N_29827,N_19897,N_23024);
nor U29828 (N_29828,N_19897,N_23996);
or U29829 (N_29829,N_23254,N_18613);
nand U29830 (N_29830,N_23494,N_19063);
xor U29831 (N_29831,N_20816,N_23771);
and U29832 (N_29832,N_21969,N_22552);
or U29833 (N_29833,N_20667,N_22279);
xor U29834 (N_29834,N_21279,N_22794);
nand U29835 (N_29835,N_20552,N_22697);
nand U29836 (N_29836,N_20048,N_20636);
nand U29837 (N_29837,N_20598,N_20005);
nand U29838 (N_29838,N_21412,N_19523);
xnor U29839 (N_29839,N_20211,N_23406);
or U29840 (N_29840,N_19263,N_21483);
nand U29841 (N_29841,N_18522,N_23647);
nand U29842 (N_29842,N_18181,N_21373);
and U29843 (N_29843,N_18397,N_22771);
nand U29844 (N_29844,N_22940,N_20527);
and U29845 (N_29845,N_21241,N_19389);
nor U29846 (N_29846,N_19394,N_22248);
or U29847 (N_29847,N_21979,N_19921);
xor U29848 (N_29848,N_19470,N_21424);
nor U29849 (N_29849,N_19368,N_19619);
nor U29850 (N_29850,N_22859,N_18051);
nor U29851 (N_29851,N_22027,N_18237);
nand U29852 (N_29852,N_20658,N_21909);
nor U29853 (N_29853,N_22088,N_21349);
nand U29854 (N_29854,N_22769,N_18608);
or U29855 (N_29855,N_18593,N_23847);
or U29856 (N_29856,N_22962,N_21637);
xnor U29857 (N_29857,N_18223,N_18211);
or U29858 (N_29858,N_18679,N_20776);
nand U29859 (N_29859,N_21215,N_22107);
nand U29860 (N_29860,N_19112,N_21862);
nor U29861 (N_29861,N_21953,N_23295);
and U29862 (N_29862,N_22456,N_18228);
nand U29863 (N_29863,N_20050,N_22763);
xnor U29864 (N_29864,N_18659,N_22602);
nand U29865 (N_29865,N_19052,N_22451);
or U29866 (N_29866,N_20332,N_23227);
or U29867 (N_29867,N_21566,N_22897);
nand U29868 (N_29868,N_19537,N_20996);
and U29869 (N_29869,N_18735,N_20070);
or U29870 (N_29870,N_23310,N_20812);
nor U29871 (N_29871,N_20660,N_21171);
nor U29872 (N_29872,N_22928,N_22110);
nor U29873 (N_29873,N_21834,N_23882);
or U29874 (N_29874,N_20831,N_19038);
nor U29875 (N_29875,N_18851,N_21035);
xnor U29876 (N_29876,N_18209,N_21664);
nor U29877 (N_29877,N_21262,N_22673);
or U29878 (N_29878,N_20769,N_22981);
nand U29879 (N_29879,N_22432,N_19940);
nor U29880 (N_29880,N_21065,N_18631);
xnor U29881 (N_29881,N_22837,N_19612);
nor U29882 (N_29882,N_22515,N_19405);
xnor U29883 (N_29883,N_23501,N_23560);
xnor U29884 (N_29884,N_23701,N_23786);
xor U29885 (N_29885,N_23871,N_22990);
xor U29886 (N_29886,N_20065,N_23125);
and U29887 (N_29887,N_20643,N_22554);
and U29888 (N_29888,N_22144,N_18672);
and U29889 (N_29889,N_19227,N_18815);
nor U29890 (N_29890,N_19684,N_18376);
nor U29891 (N_29891,N_23776,N_21348);
xor U29892 (N_29892,N_23538,N_22607);
xnor U29893 (N_29893,N_20541,N_18468);
or U29894 (N_29894,N_23670,N_23748);
or U29895 (N_29895,N_18909,N_23025);
or U29896 (N_29896,N_21029,N_20175);
nor U29897 (N_29897,N_21670,N_21908);
and U29898 (N_29898,N_20277,N_22880);
nand U29899 (N_29899,N_21310,N_20491);
and U29900 (N_29900,N_21754,N_22230);
nand U29901 (N_29901,N_21173,N_19759);
xor U29902 (N_29902,N_22845,N_23367);
and U29903 (N_29903,N_20373,N_22984);
nand U29904 (N_29904,N_22625,N_20775);
nor U29905 (N_29905,N_20776,N_22116);
xnor U29906 (N_29906,N_18542,N_20153);
xnor U29907 (N_29907,N_18477,N_23577);
nand U29908 (N_29908,N_21943,N_20494);
nand U29909 (N_29909,N_18277,N_21566);
and U29910 (N_29910,N_21301,N_23816);
or U29911 (N_29911,N_21581,N_18553);
xor U29912 (N_29912,N_22341,N_22280);
xnor U29913 (N_29913,N_20136,N_22781);
or U29914 (N_29914,N_18144,N_20741);
nor U29915 (N_29915,N_19712,N_21639);
xnor U29916 (N_29916,N_23838,N_22130);
and U29917 (N_29917,N_23510,N_20365);
nor U29918 (N_29918,N_22367,N_18995);
nor U29919 (N_29919,N_20305,N_18742);
xnor U29920 (N_29920,N_18324,N_19201);
xnor U29921 (N_29921,N_21406,N_21156);
nor U29922 (N_29922,N_21660,N_18974);
nor U29923 (N_29923,N_21991,N_21535);
and U29924 (N_29924,N_18884,N_18603);
nor U29925 (N_29925,N_19832,N_21522);
or U29926 (N_29926,N_19985,N_22112);
and U29927 (N_29927,N_19726,N_22021);
and U29928 (N_29928,N_19908,N_19007);
nor U29929 (N_29929,N_18815,N_20684);
nand U29930 (N_29930,N_20212,N_21070);
or U29931 (N_29931,N_23382,N_23425);
xor U29932 (N_29932,N_22420,N_23510);
xnor U29933 (N_29933,N_21068,N_21514);
xnor U29934 (N_29934,N_19504,N_23526);
nor U29935 (N_29935,N_23463,N_21033);
nor U29936 (N_29936,N_23067,N_22589);
and U29937 (N_29937,N_19260,N_23745);
nor U29938 (N_29938,N_18897,N_23504);
nand U29939 (N_29939,N_18050,N_20458);
and U29940 (N_29940,N_23388,N_19067);
and U29941 (N_29941,N_20848,N_22847);
nor U29942 (N_29942,N_22554,N_22573);
nor U29943 (N_29943,N_18019,N_23636);
nor U29944 (N_29944,N_18789,N_19279);
nor U29945 (N_29945,N_18237,N_22711);
nor U29946 (N_29946,N_23573,N_23089);
and U29947 (N_29947,N_23011,N_18318);
xnor U29948 (N_29948,N_18171,N_21811);
and U29949 (N_29949,N_18831,N_19462);
xnor U29950 (N_29950,N_23086,N_21812);
nand U29951 (N_29951,N_19973,N_21249);
nand U29952 (N_29952,N_18999,N_19048);
or U29953 (N_29953,N_23240,N_21932);
and U29954 (N_29954,N_19624,N_23416);
nand U29955 (N_29955,N_20991,N_23219);
and U29956 (N_29956,N_21461,N_22780);
nor U29957 (N_29957,N_18821,N_19234);
nor U29958 (N_29958,N_19001,N_21942);
or U29959 (N_29959,N_23531,N_18513);
or U29960 (N_29960,N_22852,N_19087);
nand U29961 (N_29961,N_21195,N_18055);
nor U29962 (N_29962,N_19170,N_19820);
nor U29963 (N_29963,N_19862,N_20417);
and U29964 (N_29964,N_22420,N_18026);
and U29965 (N_29965,N_18170,N_20374);
nor U29966 (N_29966,N_22282,N_20071);
xnor U29967 (N_29967,N_19961,N_18714);
and U29968 (N_29968,N_20652,N_21103);
nor U29969 (N_29969,N_22560,N_18299);
nand U29970 (N_29970,N_20852,N_23391);
nand U29971 (N_29971,N_18572,N_22138);
nor U29972 (N_29972,N_22397,N_23871);
xnor U29973 (N_29973,N_19320,N_18974);
xor U29974 (N_29974,N_22252,N_22399);
and U29975 (N_29975,N_19034,N_21711);
nor U29976 (N_29976,N_19690,N_21137);
xnor U29977 (N_29977,N_20927,N_23206);
nand U29978 (N_29978,N_18776,N_22808);
or U29979 (N_29979,N_23400,N_23865);
and U29980 (N_29980,N_20519,N_21939);
nand U29981 (N_29981,N_18630,N_18317);
xnor U29982 (N_29982,N_19337,N_23172);
xnor U29983 (N_29983,N_20027,N_18270);
or U29984 (N_29984,N_22203,N_22334);
and U29985 (N_29985,N_23719,N_19178);
and U29986 (N_29986,N_23120,N_19465);
nand U29987 (N_29987,N_21762,N_22718);
and U29988 (N_29988,N_18415,N_18062);
nor U29989 (N_29989,N_18764,N_23233);
nor U29990 (N_29990,N_21837,N_20077);
or U29991 (N_29991,N_22649,N_22046);
nand U29992 (N_29992,N_20795,N_20432);
xor U29993 (N_29993,N_20193,N_23015);
or U29994 (N_29994,N_18456,N_18243);
xor U29995 (N_29995,N_18275,N_19937);
or U29996 (N_29996,N_22728,N_22413);
xor U29997 (N_29997,N_23065,N_19891);
or U29998 (N_29998,N_20848,N_19160);
nand U29999 (N_29999,N_23097,N_20000);
or UO_0 (O_0,N_29212,N_25038);
nand UO_1 (O_1,N_28496,N_26521);
xor UO_2 (O_2,N_27537,N_24059);
nand UO_3 (O_3,N_28977,N_29826);
and UO_4 (O_4,N_28864,N_28655);
nand UO_5 (O_5,N_28383,N_28741);
nor UO_6 (O_6,N_26022,N_29442);
or UO_7 (O_7,N_27837,N_25120);
nor UO_8 (O_8,N_25986,N_24919);
or UO_9 (O_9,N_28503,N_26239);
nand UO_10 (O_10,N_25010,N_26444);
and UO_11 (O_11,N_26366,N_29043);
xor UO_12 (O_12,N_27791,N_27689);
or UO_13 (O_13,N_29423,N_26465);
nor UO_14 (O_14,N_29074,N_26960);
or UO_15 (O_15,N_25092,N_28315);
nand UO_16 (O_16,N_29628,N_28127);
nand UO_17 (O_17,N_29360,N_26194);
xnor UO_18 (O_18,N_29534,N_28836);
and UO_19 (O_19,N_28153,N_29509);
nor UO_20 (O_20,N_28087,N_24193);
nor UO_21 (O_21,N_26349,N_26724);
or UO_22 (O_22,N_25341,N_26193);
xor UO_23 (O_23,N_25366,N_25125);
xnor UO_24 (O_24,N_27684,N_29825);
xor UO_25 (O_25,N_25937,N_25242);
and UO_26 (O_26,N_26028,N_26075);
xnor UO_27 (O_27,N_28615,N_24970);
or UO_28 (O_28,N_27561,N_28043);
nand UO_29 (O_29,N_29807,N_24190);
or UO_30 (O_30,N_27571,N_29992);
xor UO_31 (O_31,N_29218,N_29105);
or UO_32 (O_32,N_28438,N_27275);
and UO_33 (O_33,N_29560,N_25916);
nor UO_34 (O_34,N_28228,N_25773);
xnor UO_35 (O_35,N_24213,N_29226);
xnor UO_36 (O_36,N_29741,N_24824);
and UO_37 (O_37,N_29202,N_26266);
nand UO_38 (O_38,N_24460,N_26766);
xnor UO_39 (O_39,N_27905,N_24790);
nand UO_40 (O_40,N_24172,N_26264);
nand UO_41 (O_41,N_27935,N_26810);
and UO_42 (O_42,N_26974,N_27906);
nor UO_43 (O_43,N_29932,N_24145);
xnor UO_44 (O_44,N_28282,N_24712);
nor UO_45 (O_45,N_27121,N_27546);
nand UO_46 (O_46,N_24323,N_26692);
xnor UO_47 (O_47,N_24903,N_29211);
xnor UO_48 (O_48,N_29362,N_28005);
nand UO_49 (O_49,N_27181,N_26614);
and UO_50 (O_50,N_28140,N_24705);
nand UO_51 (O_51,N_27487,N_29134);
xnor UO_52 (O_52,N_26233,N_24104);
nand UO_53 (O_53,N_29852,N_27196);
or UO_54 (O_54,N_28855,N_28587);
nand UO_55 (O_55,N_29849,N_29890);
xnor UO_56 (O_56,N_24252,N_29173);
or UO_57 (O_57,N_28968,N_27520);
xnor UO_58 (O_58,N_27719,N_25380);
nor UO_59 (O_59,N_26751,N_25741);
and UO_60 (O_60,N_27336,N_26676);
nor UO_61 (O_61,N_29735,N_25776);
nand UO_62 (O_62,N_26740,N_29650);
nand UO_63 (O_63,N_25255,N_28782);
and UO_64 (O_64,N_27038,N_27293);
and UO_65 (O_65,N_29129,N_28622);
nand UO_66 (O_66,N_24862,N_24174);
or UO_67 (O_67,N_28547,N_28419);
and UO_68 (O_68,N_25067,N_26402);
and UO_69 (O_69,N_24277,N_28812);
or UO_70 (O_70,N_24444,N_25737);
and UO_71 (O_71,N_29749,N_25110);
or UO_72 (O_72,N_27399,N_26454);
xor UO_73 (O_73,N_26338,N_24958);
nor UO_74 (O_74,N_26341,N_26330);
nor UO_75 (O_75,N_24209,N_24463);
or UO_76 (O_76,N_26917,N_24877);
nand UO_77 (O_77,N_26360,N_27156);
and UO_78 (O_78,N_25686,N_24118);
and UO_79 (O_79,N_25562,N_24366);
xnor UO_80 (O_80,N_25188,N_27084);
nand UO_81 (O_81,N_29032,N_27506);
nand UO_82 (O_82,N_26520,N_27144);
xor UO_83 (O_83,N_25166,N_27712);
xnor UO_84 (O_84,N_24244,N_26382);
or UO_85 (O_85,N_29305,N_28976);
nand UO_86 (O_86,N_24287,N_27030);
nand UO_87 (O_87,N_24803,N_27702);
and UO_88 (O_88,N_27957,N_28200);
xnor UO_89 (O_89,N_26284,N_26448);
and UO_90 (O_90,N_27620,N_29346);
xor UO_91 (O_91,N_28959,N_25088);
nand UO_92 (O_92,N_27381,N_28771);
xor UO_93 (O_93,N_27106,N_29791);
xnor UO_94 (O_94,N_29200,N_28159);
nor UO_95 (O_95,N_28355,N_28400);
and UO_96 (O_96,N_24815,N_28004);
nand UO_97 (O_97,N_29088,N_29175);
xnor UO_98 (O_98,N_27840,N_25457);
and UO_99 (O_99,N_24844,N_28360);
nand UO_100 (O_100,N_25684,N_29819);
nand UO_101 (O_101,N_26260,N_29958);
xnor UO_102 (O_102,N_27198,N_29050);
nand UO_103 (O_103,N_27243,N_25960);
or UO_104 (O_104,N_25841,N_26359);
nor UO_105 (O_105,N_29926,N_28962);
nor UO_106 (O_106,N_28709,N_24294);
or UO_107 (O_107,N_28000,N_26802);
xor UO_108 (O_108,N_24312,N_25585);
nor UO_109 (O_109,N_28745,N_26643);
nor UO_110 (O_110,N_27061,N_27298);
nand UO_111 (O_111,N_25448,N_26946);
nor UO_112 (O_112,N_28134,N_28204);
and UO_113 (O_113,N_27825,N_27942);
xnor UO_114 (O_114,N_29702,N_26579);
and UO_115 (O_115,N_25261,N_25049);
and UO_116 (O_116,N_27480,N_25523);
nand UO_117 (O_117,N_28729,N_29917);
nor UO_118 (O_118,N_28521,N_25648);
or UO_119 (O_119,N_26700,N_24881);
nand UO_120 (O_120,N_26673,N_26224);
xor UO_121 (O_121,N_26298,N_24084);
or UO_122 (O_122,N_24381,N_26098);
nor UO_123 (O_123,N_28452,N_27975);
nand UO_124 (O_124,N_26540,N_29995);
and UO_125 (O_125,N_24820,N_27968);
xnor UO_126 (O_126,N_27730,N_24330);
or UO_127 (O_127,N_27530,N_25520);
nand UO_128 (O_128,N_28230,N_25138);
nor UO_129 (O_129,N_28209,N_26154);
nor UO_130 (O_130,N_28088,N_26555);
and UO_131 (O_131,N_24101,N_29303);
nand UO_132 (O_132,N_25427,N_27971);
or UO_133 (O_133,N_26843,N_27227);
and UO_134 (O_134,N_26009,N_26404);
and UO_135 (O_135,N_26425,N_27019);
nand UO_136 (O_136,N_27751,N_27648);
xor UO_137 (O_137,N_26007,N_29607);
nor UO_138 (O_138,N_27956,N_26162);
nand UO_139 (O_139,N_28735,N_24432);
xor UO_140 (O_140,N_29492,N_29788);
and UO_141 (O_141,N_25671,N_26563);
nand UO_142 (O_142,N_26636,N_26267);
xnor UO_143 (O_143,N_27586,N_27257);
nor UO_144 (O_144,N_26778,N_26706);
xnor UO_145 (O_145,N_24069,N_29642);
or UO_146 (O_146,N_24063,N_26829);
nor UO_147 (O_147,N_29051,N_27829);
or UO_148 (O_148,N_27394,N_28131);
nand UO_149 (O_149,N_29014,N_24818);
nand UO_150 (O_150,N_24907,N_27043);
or UO_151 (O_151,N_24886,N_27570);
xor UO_152 (O_152,N_26570,N_28664);
or UO_153 (O_153,N_29945,N_29431);
or UO_154 (O_154,N_28386,N_27070);
or UO_155 (O_155,N_26453,N_27961);
and UO_156 (O_156,N_25325,N_29424);
and UO_157 (O_157,N_25678,N_27636);
nand UO_158 (O_158,N_29794,N_27550);
and UO_159 (O_159,N_27296,N_29367);
and UO_160 (O_160,N_25158,N_29946);
xnor UO_161 (O_161,N_29839,N_24028);
and UO_162 (O_162,N_29304,N_25269);
xor UO_163 (O_163,N_26245,N_25506);
xnor UO_164 (O_164,N_27461,N_27585);
and UO_165 (O_165,N_29462,N_24737);
nor UO_166 (O_166,N_28757,N_26683);
or UO_167 (O_167,N_27619,N_24834);
or UO_168 (O_168,N_26305,N_24533);
and UO_169 (O_169,N_28732,N_27912);
and UO_170 (O_170,N_27511,N_26400);
and UO_171 (O_171,N_25938,N_29656);
nor UO_172 (O_172,N_26696,N_27077);
nor UO_173 (O_173,N_29066,N_29520);
xor UO_174 (O_174,N_25935,N_27678);
nor UO_175 (O_175,N_25486,N_25783);
xnor UO_176 (O_176,N_26278,N_24730);
nand UO_177 (O_177,N_29372,N_25211);
and UO_178 (O_178,N_29883,N_27265);
or UO_179 (O_179,N_26455,N_27143);
nor UO_180 (O_180,N_29556,N_27765);
nor UO_181 (O_181,N_27414,N_27855);
or UO_182 (O_182,N_26628,N_26450);
and UO_183 (O_183,N_25328,N_29856);
nand UO_184 (O_184,N_29308,N_27380);
or UO_185 (O_185,N_29836,N_28966);
or UO_186 (O_186,N_27563,N_25665);
xor UO_187 (O_187,N_24991,N_27781);
nor UO_188 (O_188,N_26471,N_26482);
nor UO_189 (O_189,N_29001,N_29652);
nor UO_190 (O_190,N_28198,N_27788);
or UO_191 (O_191,N_28486,N_27523);
nor UO_192 (O_192,N_24857,N_27587);
nand UO_193 (O_193,N_25844,N_28338);
or UO_194 (O_194,N_27710,N_29624);
xnor UO_195 (O_195,N_26263,N_28356);
nand UO_196 (O_196,N_24466,N_28196);
and UO_197 (O_197,N_26408,N_26259);
nand UO_198 (O_198,N_27989,N_27090);
nand UO_199 (O_199,N_26847,N_29625);
and UO_200 (O_200,N_27708,N_28985);
xnor UO_201 (O_201,N_28094,N_25690);
or UO_202 (O_202,N_24679,N_28441);
or UO_203 (O_203,N_28916,N_29888);
xnor UO_204 (O_204,N_29815,N_25253);
or UO_205 (O_205,N_29457,N_26253);
and UO_206 (O_206,N_24643,N_24915);
or UO_207 (O_207,N_28256,N_28633);
nor UO_208 (O_208,N_28826,N_28493);
xor UO_209 (O_209,N_24331,N_28425);
nand UO_210 (O_210,N_25928,N_29497);
nand UO_211 (O_211,N_28744,N_25271);
nand UO_212 (O_212,N_24863,N_29910);
nand UO_213 (O_213,N_26530,N_24576);
nor UO_214 (O_214,N_24518,N_29990);
xor UO_215 (O_215,N_26241,N_28460);
and UO_216 (O_216,N_25335,N_27002);
and UO_217 (O_217,N_25393,N_25435);
or UO_218 (O_218,N_26844,N_26593);
and UO_219 (O_219,N_25742,N_28853);
xor UO_220 (O_220,N_29953,N_29366);
or UO_221 (O_221,N_27192,N_29260);
xnor UO_222 (O_222,N_27656,N_25514);
and UO_223 (O_223,N_25617,N_25066);
xnor UO_224 (O_224,N_28764,N_25022);
nor UO_225 (O_225,N_29964,N_24885);
xor UO_226 (O_226,N_26424,N_25672);
or UO_227 (O_227,N_28108,N_25870);
nand UO_228 (O_228,N_29673,N_29444);
or UO_229 (O_229,N_25172,N_24667);
nand UO_230 (O_230,N_25473,N_26783);
nor UO_231 (O_231,N_24508,N_29393);
xnor UO_232 (O_232,N_29750,N_26719);
xor UO_233 (O_233,N_27015,N_24562);
nand UO_234 (O_234,N_28669,N_24509);
xnor UO_235 (O_235,N_28007,N_26542);
xor UO_236 (O_236,N_25679,N_26927);
nand UO_237 (O_237,N_28728,N_29712);
and UO_238 (O_238,N_29023,N_25029);
nor UO_239 (O_239,N_29668,N_29510);
xor UO_240 (O_240,N_25812,N_26189);
xor UO_241 (O_241,N_26979,N_24399);
nor UO_242 (O_242,N_24453,N_29635);
nor UO_243 (O_243,N_26935,N_25397);
and UO_244 (O_244,N_27185,N_25804);
and UO_245 (O_245,N_27016,N_28803);
nor UO_246 (O_246,N_25477,N_29760);
or UO_247 (O_247,N_29236,N_24767);
and UO_248 (O_248,N_28848,N_28036);
and UO_249 (O_249,N_24128,N_29486);
nor UO_250 (O_250,N_29550,N_28746);
nand UO_251 (O_251,N_29344,N_26097);
xor UO_252 (O_252,N_28321,N_28789);
nor UO_253 (O_253,N_26665,N_29041);
xnor UO_254 (O_254,N_27013,N_27735);
nor UO_255 (O_255,N_24214,N_26617);
nor UO_256 (O_256,N_28023,N_25145);
nor UO_257 (O_257,N_28090,N_27037);
and UO_258 (O_258,N_25183,N_24723);
or UO_259 (O_259,N_25577,N_24935);
or UO_260 (O_260,N_25368,N_28594);
nor UO_261 (O_261,N_29940,N_28469);
nand UO_262 (O_262,N_28630,N_25755);
nor UO_263 (O_263,N_25511,N_26965);
and UO_264 (O_264,N_25717,N_28822);
and UO_265 (O_265,N_24969,N_24302);
and UO_266 (O_266,N_29232,N_29908);
or UO_267 (O_267,N_28278,N_29600);
nand UO_268 (O_268,N_24720,N_29925);
and UO_269 (O_269,N_29927,N_27771);
or UO_270 (O_270,N_29118,N_28894);
nor UO_271 (O_271,N_24695,N_27998);
nor UO_272 (O_272,N_25867,N_28257);
nand UO_273 (O_273,N_29508,N_26871);
xor UO_274 (O_274,N_27488,N_24414);
nor UO_275 (O_275,N_25354,N_26833);
nor UO_276 (O_276,N_25074,N_27929);
nor UO_277 (O_277,N_26793,N_25208);
xor UO_278 (O_278,N_24071,N_28676);
xor UO_279 (O_279,N_28212,N_25519);
xnor UO_280 (O_280,N_29104,N_25784);
and UO_281 (O_281,N_29403,N_25861);
nand UO_282 (O_282,N_29732,N_27035);
or UO_283 (O_283,N_28265,N_29469);
or UO_284 (O_284,N_24872,N_26878);
nand UO_285 (O_285,N_25787,N_25089);
or UO_286 (O_286,N_26609,N_26115);
nor UO_287 (O_287,N_25749,N_29265);
nand UO_288 (O_288,N_27369,N_29827);
nor UO_289 (O_289,N_24501,N_25611);
xor UO_290 (O_290,N_28473,N_27711);
or UO_291 (O_291,N_28941,N_27311);
nor UO_292 (O_292,N_27299,N_27897);
and UO_293 (O_293,N_29296,N_29706);
nor UO_294 (O_294,N_28681,N_29555);
nor UO_295 (O_295,N_24557,N_29857);
xor UO_296 (O_296,N_28385,N_27934);
nor UO_297 (O_297,N_25663,N_28592);
and UO_298 (O_298,N_24105,N_28289);
or UO_299 (O_299,N_27927,N_24457);
xnor UO_300 (O_300,N_27830,N_24814);
nor UO_301 (O_301,N_26205,N_27376);
or UO_302 (O_302,N_28387,N_26779);
xnor UO_303 (O_303,N_26608,N_28561);
or UO_304 (O_304,N_29401,N_25304);
nand UO_305 (O_305,N_26013,N_25996);
nor UO_306 (O_306,N_25370,N_24925);
or UO_307 (O_307,N_27747,N_27465);
and UO_308 (O_308,N_24655,N_25516);
nand UO_309 (O_309,N_26368,N_26414);
nor UO_310 (O_310,N_27101,N_26438);
nor UO_311 (O_311,N_24391,N_28297);
nor UO_312 (O_312,N_29752,N_27877);
nor UO_313 (O_313,N_29714,N_26145);
nor UO_314 (O_314,N_24204,N_26499);
and UO_315 (O_315,N_24228,N_25869);
xor UO_316 (O_316,N_29195,N_29592);
and UO_317 (O_317,N_24517,N_29021);
nor UO_318 (O_318,N_25973,N_28115);
or UO_319 (O_319,N_26822,N_28897);
nor UO_320 (O_320,N_25399,N_25987);
and UO_321 (O_321,N_29008,N_28427);
and UO_322 (O_322,N_26672,N_29152);
or UO_323 (O_323,N_28544,N_27372);
or UO_324 (O_324,N_28406,N_25326);
and UO_325 (O_325,N_29655,N_26983);
or UO_326 (O_326,N_28984,N_25279);
nand UO_327 (O_327,N_27976,N_29037);
nor UO_328 (O_328,N_26987,N_26350);
or UO_329 (O_329,N_26486,N_26926);
nand UO_330 (O_330,N_25568,N_29898);
xnor UO_331 (O_331,N_28605,N_29568);
or UO_332 (O_332,N_25860,N_25962);
nand UO_333 (O_333,N_28668,N_24591);
nand UO_334 (O_334,N_24434,N_29539);
and UO_335 (O_335,N_29280,N_24053);
nor UO_336 (O_336,N_26774,N_24550);
xnor UO_337 (O_337,N_29047,N_29433);
nand UO_338 (O_338,N_26911,N_24464);
nand UO_339 (O_339,N_28055,N_25006);
xnor UO_340 (O_340,N_29095,N_29817);
nand UO_341 (O_341,N_24574,N_24709);
nor UO_342 (O_342,N_28832,N_26762);
nand UO_343 (O_343,N_25754,N_28505);
and UO_344 (O_344,N_25410,N_28781);
nand UO_345 (O_345,N_26303,N_24589);
or UO_346 (O_346,N_24014,N_29078);
or UO_347 (O_347,N_24369,N_27021);
and UO_348 (O_348,N_28060,N_27431);
or UO_349 (O_349,N_29699,N_26637);
and UO_350 (O_350,N_24904,N_28589);
and UO_351 (O_351,N_24644,N_29334);
nor UO_352 (O_352,N_26120,N_28957);
nor UO_353 (O_353,N_28214,N_25768);
nand UO_354 (O_354,N_29079,N_25956);
xnor UO_355 (O_355,N_29025,N_25813);
nor UO_356 (O_356,N_29793,N_27325);
or UO_357 (O_357,N_28736,N_24560);
or UO_358 (O_358,N_25015,N_25636);
and UO_359 (O_359,N_26738,N_24532);
nand UO_360 (O_360,N_26393,N_28494);
and UO_361 (O_361,N_27749,N_27580);
and UO_362 (O_362,N_24371,N_24718);
xor UO_363 (O_363,N_29179,N_27445);
and UO_364 (O_364,N_27756,N_29676);
nand UO_365 (O_365,N_26122,N_27460);
or UO_366 (O_366,N_29385,N_28501);
nand UO_367 (O_367,N_24853,N_26769);
and UO_368 (O_368,N_24087,N_24119);
xor UO_369 (O_369,N_26331,N_27979);
or UO_370 (O_370,N_29956,N_24774);
and UO_371 (O_371,N_25296,N_27273);
nand UO_372 (O_372,N_24048,N_28234);
nor UO_373 (O_373,N_29601,N_27672);
nor UO_374 (O_374,N_25180,N_29693);
xnor UO_375 (O_375,N_29980,N_27657);
and UO_376 (O_376,N_28080,N_25213);
and UO_377 (O_377,N_28291,N_29086);
xor UO_378 (O_378,N_29689,N_28654);
and UO_379 (O_379,N_28111,N_25609);
or UO_380 (O_380,N_26051,N_25883);
or UO_381 (O_381,N_25699,N_26014);
or UO_382 (O_382,N_24531,N_24687);
nand UO_383 (O_383,N_24127,N_25373);
and UO_384 (O_384,N_24941,N_25441);
xor UO_385 (O_385,N_24047,N_24164);
or UO_386 (O_386,N_28275,N_28980);
nand UO_387 (O_387,N_28382,N_29778);
and UO_388 (O_388,N_25235,N_29802);
nor UO_389 (O_389,N_26685,N_24416);
nor UO_390 (O_390,N_24243,N_27110);
xor UO_391 (O_391,N_26849,N_26717);
or UO_392 (O_392,N_25982,N_28918);
nand UO_393 (O_393,N_25897,N_28133);
and UO_394 (O_394,N_25329,N_28084);
xor UO_395 (O_395,N_27500,N_27824);
nor UO_396 (O_396,N_24627,N_29833);
xor UO_397 (O_397,N_29414,N_28333);
or UO_398 (O_398,N_24765,N_29087);
nand UO_399 (O_399,N_24749,N_26436);
or UO_400 (O_400,N_29251,N_25542);
nor UO_401 (O_401,N_28990,N_27297);
xor UO_402 (O_402,N_29197,N_29746);
and UO_403 (O_403,N_29279,N_25412);
or UO_404 (O_404,N_27249,N_27304);
nor UO_405 (O_405,N_24044,N_29016);
xnor UO_406 (O_406,N_27800,N_28266);
nand UO_407 (O_407,N_25574,N_29868);
or UO_408 (O_408,N_27028,N_27007);
nand UO_409 (O_409,N_29068,N_27029);
nor UO_410 (O_410,N_24448,N_25774);
or UO_411 (O_411,N_25789,N_25534);
or UO_412 (O_412,N_24217,N_26040);
and UO_413 (O_413,N_27759,N_29426);
nand UO_414 (O_414,N_27239,N_29184);
or UO_415 (O_415,N_29850,N_25992);
nor UO_416 (O_416,N_26524,N_25706);
nor UO_417 (O_417,N_25418,N_29420);
nor UO_418 (O_418,N_25102,N_29022);
or UO_419 (O_419,N_27644,N_26526);
or UO_420 (O_420,N_24895,N_27051);
nand UO_421 (O_421,N_25829,N_29713);
nand UO_422 (O_422,N_24600,N_27456);
or UO_423 (O_423,N_29233,N_25311);
xor UO_424 (O_424,N_26615,N_25549);
xnor UO_425 (O_425,N_28331,N_27491);
or UO_426 (O_426,N_28193,N_26619);
nand UO_427 (O_427,N_29075,N_24019);
xnor UO_428 (O_428,N_29797,N_26651);
xnor UO_429 (O_429,N_26680,N_25785);
or UO_430 (O_430,N_28788,N_25876);
nand UO_431 (O_431,N_28490,N_29643);
nor UO_432 (O_432,N_26859,N_27387);
xnor UO_433 (O_433,N_29879,N_25673);
and UO_434 (O_434,N_28430,N_24514);
or UO_435 (O_435,N_27876,N_24425);
or UO_436 (O_436,N_25472,N_26140);
nor UO_437 (O_437,N_27923,N_29842);
nand UO_438 (O_438,N_28670,N_27229);
nor UO_439 (O_439,N_27789,N_28931);
nor UO_440 (O_440,N_24265,N_27050);
and UO_441 (O_441,N_29496,N_29342);
nor UO_442 (O_442,N_25414,N_27661);
nand UO_443 (O_443,N_27024,N_25443);
and UO_444 (O_444,N_26556,N_26012);
nor UO_445 (O_445,N_26679,N_29666);
nor UO_446 (O_446,N_25465,N_25406);
nand UO_447 (O_447,N_26046,N_28071);
or UO_448 (O_448,N_26959,N_25426);
xor UO_449 (O_449,N_25078,N_26909);
xor UO_450 (O_450,N_26668,N_26202);
and UO_451 (O_451,N_24304,N_29349);
xor UO_452 (O_452,N_25420,N_28028);
nand UO_453 (O_453,N_26693,N_27870);
nor UO_454 (O_454,N_24083,N_27111);
or UO_455 (O_455,N_24382,N_25163);
nand UO_456 (O_456,N_29163,N_26481);
or UO_457 (O_457,N_28927,N_25793);
or UO_458 (O_458,N_25605,N_27251);
nor UO_459 (O_459,N_24739,N_24337);
nand UO_460 (O_460,N_24171,N_27107);
and UO_461 (O_461,N_28763,N_24882);
or UO_462 (O_462,N_25278,N_29004);
or UO_463 (O_463,N_28439,N_27569);
and UO_464 (O_464,N_26033,N_24951);
xor UO_465 (O_465,N_26541,N_25763);
nor UO_466 (O_466,N_27610,N_28251);
nand UO_467 (O_467,N_27553,N_25898);
and UO_468 (O_468,N_28591,N_26925);
and UO_469 (O_469,N_26883,N_28138);
nor UO_470 (O_470,N_25434,N_27396);
and UO_471 (O_471,N_25280,N_25238);
nand UO_472 (O_472,N_26958,N_29514);
nand UO_473 (O_473,N_24937,N_29489);
nor UO_474 (O_474,N_26602,N_24947);
nand UO_475 (O_475,N_27300,N_25892);
nor UO_476 (O_476,N_29172,N_29532);
and UO_477 (O_477,N_24959,N_25135);
xnor UO_478 (O_478,N_25178,N_26509);
and UO_479 (O_479,N_28484,N_24811);
or UO_480 (O_480,N_25584,N_26067);
or UO_481 (O_481,N_29805,N_24153);
or UO_482 (O_482,N_26708,N_29804);
and UO_483 (O_483,N_26389,N_26613);
nor UO_484 (O_484,N_26403,N_29769);
nor UO_485 (O_485,N_24511,N_25769);
nand UO_486 (O_486,N_24394,N_25361);
or UO_487 (O_487,N_29939,N_28286);
xnor UO_488 (O_488,N_29217,N_28048);
and UO_489 (O_489,N_27400,N_25517);
nand UO_490 (O_490,N_27447,N_25217);
xnor UO_491 (O_491,N_26969,N_25203);
xor UO_492 (O_492,N_24408,N_25091);
or UO_493 (O_493,N_26136,N_28020);
nor UO_494 (O_494,N_25228,N_28773);
nor UO_495 (O_495,N_25714,N_28336);
or UO_496 (O_496,N_28524,N_26928);
nand UO_497 (O_497,N_25739,N_28653);
xnor UO_498 (O_498,N_25174,N_29895);
xnor UO_499 (O_499,N_28556,N_26568);
nor UO_500 (O_500,N_27108,N_27823);
and UO_501 (O_501,N_25411,N_24849);
nand UO_502 (O_502,N_27986,N_28872);
and UO_503 (O_503,N_26944,N_25118);
nor UO_504 (O_504,N_28079,N_28250);
xor UO_505 (O_505,N_26644,N_29764);
nor UO_506 (O_506,N_26899,N_27668);
nor UO_507 (O_507,N_26112,N_29731);
xor UO_508 (O_508,N_24165,N_24492);
or UO_509 (O_509,N_25433,N_24353);
and UO_510 (O_510,N_27462,N_25129);
xor UO_511 (O_511,N_26785,N_28528);
nor UO_512 (O_512,N_25849,N_24035);
nor UO_513 (O_513,N_25833,N_24218);
xnor UO_514 (O_514,N_26003,N_26798);
nor UO_515 (O_515,N_25291,N_28969);
nor UO_516 (O_516,N_24505,N_27764);
nand UO_517 (O_517,N_28687,N_29038);
and UO_518 (O_518,N_28139,N_27011);
or UO_519 (O_519,N_29222,N_26328);
nor UO_520 (O_520,N_26016,N_25744);
nor UO_521 (O_521,N_28562,N_27034);
and UO_522 (O_522,N_29314,N_27856);
nor UO_523 (O_523,N_26276,N_24481);
nor UO_524 (O_524,N_25028,N_25976);
and UO_525 (O_525,N_28703,N_24017);
nor UO_526 (O_526,N_24734,N_25186);
or UO_527 (O_527,N_28666,N_25264);
and UO_528 (O_528,N_27152,N_27471);
nor UO_529 (O_529,N_26200,N_24634);
nor UO_530 (O_530,N_25529,N_24772);
or UO_531 (O_531,N_24953,N_27092);
or UO_532 (O_532,N_25848,N_27053);
xnor UO_533 (O_533,N_24040,N_28190);
or UO_534 (O_534,N_26121,N_25512);
and UO_535 (O_535,N_27947,N_26777);
or UO_536 (O_536,N_25734,N_24356);
nand UO_537 (O_537,N_25207,N_24282);
xor UO_538 (O_538,N_29092,N_28628);
or UO_539 (O_539,N_24160,N_28619);
xor UO_540 (O_540,N_25277,N_28551);
xnor UO_541 (O_541,N_27256,N_29239);
nor UO_542 (O_542,N_29962,N_27333);
nand UO_543 (O_543,N_25111,N_25447);
and UO_544 (O_544,N_25500,N_28328);
xor UO_545 (O_545,N_27221,N_24604);
nand UO_546 (O_546,N_26083,N_26753);
nand UO_547 (O_547,N_26603,N_25199);
nand UO_548 (O_548,N_26410,N_25582);
nand UO_549 (O_549,N_24022,N_29459);
nand UO_550 (O_550,N_25194,N_28498);
and UO_551 (O_551,N_24890,N_26898);
and UO_552 (O_552,N_24583,N_28737);
nor UO_553 (O_553,N_28413,N_24944);
nand UO_554 (O_554,N_26734,N_27260);
nand UO_555 (O_555,N_27655,N_26826);
and UO_556 (O_556,N_29036,N_26870);
xor UO_557 (O_557,N_27810,N_25788);
or UO_558 (O_558,N_27210,N_29498);
or UO_559 (O_559,N_26144,N_29138);
and UO_560 (O_560,N_27266,N_24784);
nor UO_561 (O_561,N_27535,N_24155);
or UO_562 (O_562,N_25864,N_25002);
or UO_563 (O_563,N_29262,N_26257);
or UO_564 (O_564,N_27930,N_24923);
or UO_565 (O_565,N_29448,N_29575);
nor UO_566 (O_566,N_24307,N_28983);
nor UO_567 (O_567,N_25588,N_29863);
and UO_568 (O_568,N_27081,N_27258);
xnor UO_569 (O_569,N_28804,N_27131);
nand UO_570 (O_570,N_27475,N_27573);
nand UO_571 (O_571,N_28261,N_28049);
nand UO_572 (O_572,N_27150,N_27952);
or UO_573 (O_573,N_28565,N_29144);
nor UO_574 (O_574,N_28888,N_28724);
and UO_575 (O_575,N_29743,N_29331);
and UO_576 (O_576,N_26709,N_27801);
or UO_577 (O_577,N_27413,N_25001);
and UO_578 (O_578,N_25603,N_24728);
or UO_579 (O_579,N_29187,N_24738);
xnor UO_580 (O_580,N_24011,N_26495);
nand UO_581 (O_581,N_27130,N_28810);
nor UO_582 (O_582,N_28939,N_28530);
and UO_583 (O_583,N_27262,N_26886);
nor UO_584 (O_584,N_24336,N_29872);
or UO_585 (O_585,N_25231,N_27315);
xnor UO_586 (O_586,N_26431,N_26788);
nor UO_587 (O_587,N_25195,N_26446);
nand UO_588 (O_588,N_28099,N_26288);
nor UO_589 (O_589,N_29874,N_24582);
nand UO_590 (O_590,N_25879,N_29640);
nor UO_591 (O_591,N_27344,N_27207);
nor UO_592 (O_592,N_27845,N_29470);
xnor UO_593 (O_593,N_26817,N_29010);
nor UO_594 (O_594,N_24779,N_27835);
or UO_595 (O_595,N_26346,N_24202);
and UO_596 (O_596,N_29970,N_27232);
nor UO_597 (O_597,N_26392,N_24592);
xnor UO_598 (O_598,N_27858,N_28022);
or UO_599 (O_599,N_29353,N_25702);
nand UO_600 (O_600,N_29739,N_25371);
or UO_601 (O_601,N_27323,N_29546);
xnor UO_602 (O_602,N_26825,N_28816);
and UO_603 (O_603,N_24446,N_28695);
or UO_604 (O_604,N_24598,N_26168);
xor UO_605 (O_605,N_29573,N_29914);
nand UO_606 (O_606,N_27900,N_24392);
and UO_607 (O_607,N_24152,N_28847);
or UO_608 (O_608,N_28326,N_26739);
nand UO_609 (O_609,N_28052,N_29647);
or UO_610 (O_610,N_29090,N_24081);
xor UO_611 (O_611,N_24789,N_25175);
nor UO_612 (O_612,N_26084,N_29323);
nand UO_613 (O_613,N_24752,N_25378);
nand UO_614 (O_614,N_29950,N_26184);
xnor UO_615 (O_615,N_27426,N_24280);
nand UO_616 (O_616,N_25115,N_28861);
nor UO_617 (O_617,N_25683,N_27102);
or UO_618 (O_618,N_24185,N_29456);
nand UO_619 (O_619,N_28248,N_26261);
or UO_620 (O_620,N_28518,N_29324);
xnor UO_621 (O_621,N_26496,N_27993);
xor UO_622 (O_622,N_29255,N_24373);
xnor UO_623 (O_623,N_27008,N_24563);
nand UO_624 (O_624,N_24144,N_24838);
nand UO_625 (O_625,N_27969,N_28458);
nand UO_626 (O_626,N_24438,N_25456);
nor UO_627 (O_627,N_24299,N_29847);
xor UO_628 (O_628,N_26999,N_26271);
nand UO_629 (O_629,N_24112,N_24565);
nor UO_630 (O_630,N_24465,N_27161);
nand UO_631 (O_631,N_26721,N_27446);
and UO_632 (O_632,N_27324,N_26065);
or UO_633 (O_633,N_25917,N_27331);
xor UO_634 (O_634,N_28914,N_29810);
or UO_635 (O_635,N_26150,N_27485);
xnor UO_636 (O_636,N_26045,N_26884);
nor UO_637 (O_637,N_26277,N_29564);
nand UO_638 (O_638,N_25452,N_26091);
xor UO_639 (O_639,N_24626,N_24701);
nor UO_640 (O_640,N_28899,N_26674);
or UO_641 (O_641,N_28073,N_24039);
and UO_642 (O_642,N_27200,N_27409);
nand UO_643 (O_643,N_25141,N_24461);
nor UO_644 (O_644,N_26029,N_28322);
xnor UO_645 (O_645,N_26327,N_26544);
or UO_646 (O_646,N_29157,N_27201);
and UO_647 (O_647,N_24556,N_29521);
xnor UO_648 (O_648,N_26291,N_26720);
xor UO_649 (O_649,N_26323,N_27980);
nand UO_650 (O_650,N_25358,N_28814);
nand UO_651 (O_651,N_25794,N_27023);
xnor UO_652 (O_652,N_24227,N_25934);
xor UO_653 (O_653,N_24226,N_28921);
xor UO_654 (O_654,N_29558,N_24628);
nand UO_655 (O_655,N_28327,N_25623);
nor UO_656 (O_656,N_29434,N_24298);
xor UO_657 (O_657,N_24607,N_24281);
xor UO_658 (O_658,N_25113,N_27223);
or UO_659 (O_659,N_25945,N_28097);
xnor UO_660 (O_660,N_25797,N_28924);
or UO_661 (O_661,N_25190,N_24581);
and UO_662 (O_662,N_29224,N_24833);
and UO_663 (O_663,N_27147,N_26816);
and UO_664 (O_664,N_24996,N_27390);
xnor UO_665 (O_665,N_27354,N_25062);
nand UO_666 (O_666,N_26552,N_29604);
and UO_667 (O_667,N_28423,N_25518);
nor UO_668 (O_668,N_24891,N_24625);
and UO_669 (O_669,N_24177,N_28740);
or UO_670 (O_670,N_26841,N_24076);
or UO_671 (O_671,N_24681,N_28118);
nand UO_672 (O_672,N_29180,N_25347);
and UO_673 (O_673,N_28156,N_26605);
and UO_674 (O_674,N_27303,N_27466);
nand UO_675 (O_675,N_24293,N_28476);
and UO_676 (O_676,N_26659,N_24852);
and UO_677 (O_677,N_29028,N_25748);
xor UO_678 (O_678,N_27752,N_25273);
xor UO_679 (O_679,N_29130,N_24805);
and UO_680 (O_680,N_26854,N_24007);
nand UO_681 (O_681,N_28553,N_28369);
and UO_682 (O_682,N_27495,N_26686);
nand UO_683 (O_683,N_29419,N_26573);
and UO_684 (O_684,N_27448,N_24559);
xor UO_685 (O_685,N_29286,N_28273);
nor UO_686 (O_686,N_26066,N_25920);
nor UO_687 (O_687,N_27302,N_29478);
xor UO_688 (O_688,N_24763,N_24699);
or UO_689 (O_689,N_27691,N_26661);
xnor UO_690 (O_690,N_29516,N_25246);
nor UO_691 (O_691,N_28032,N_28402);
or UO_692 (O_692,N_28951,N_29891);
nand UO_693 (O_693,N_27317,N_27847);
nor UO_694 (O_694,N_24787,N_27499);
or UO_695 (O_695,N_29013,N_29924);
and UO_696 (O_696,N_24555,N_25726);
and UO_697 (O_697,N_27795,N_25640);
and UO_698 (O_698,N_28839,N_26996);
and UO_699 (O_699,N_28779,N_25583);
nor UO_700 (O_700,N_25669,N_28571);
nand UO_701 (O_701,N_29566,N_25889);
nand UO_702 (O_702,N_29114,N_24472);
nand UO_703 (O_703,N_24449,N_27866);
nand UO_704 (O_704,N_29168,N_28418);
or UO_705 (O_705,N_24956,N_25547);
nor UO_706 (O_706,N_27109,N_29873);
nand UO_707 (O_707,N_24736,N_24978);
xnor UO_708 (O_708,N_25119,N_24181);
nor UO_709 (O_709,N_29537,N_27745);
nor UO_710 (O_710,N_24260,N_27205);
and UO_711 (O_711,N_27528,N_28167);
nor UO_712 (O_712,N_29881,N_24691);
and UO_713 (O_713,N_24782,N_24497);
nor UO_714 (O_714,N_29757,N_28281);
xor UO_715 (O_715,N_25193,N_28199);
or UO_716 (O_716,N_28375,N_26319);
and UO_717 (O_717,N_26590,N_27006);
nand UO_718 (O_718,N_26176,N_29283);
or UO_719 (O_719,N_27532,N_26689);
nor UO_720 (O_720,N_26159,N_29972);
and UO_721 (O_721,N_25856,N_26477);
xor UO_722 (O_722,N_24865,N_24621);
or UO_723 (O_723,N_27355,N_29859);
xor UO_724 (O_724,N_26557,N_24315);
xnor UO_725 (O_725,N_29846,N_25628);
xnor UO_726 (O_726,N_27513,N_27531);
nor UO_727 (O_727,N_25137,N_24162);
nand UO_728 (O_728,N_26395,N_27424);
nand UO_729 (O_729,N_29775,N_25818);
xnor UO_730 (O_730,N_29292,N_26729);
and UO_731 (O_731,N_26160,N_29756);
xor UO_732 (O_732,N_29035,N_28599);
or UO_733 (O_733,N_25413,N_29267);
or UO_734 (O_734,N_26714,N_29428);
nand UO_735 (O_735,N_25564,N_24700);
xor UO_736 (O_736,N_28875,N_28301);
nor UO_737 (O_737,N_29397,N_26601);
nand UO_738 (O_738,N_29340,N_26550);
xor UO_739 (O_739,N_29453,N_26308);
or UO_740 (O_740,N_26836,N_24305);
xnor UO_741 (O_741,N_27617,N_29072);
and UO_742 (O_742,N_28169,N_25364);
xnor UO_743 (O_743,N_25011,N_28993);
or UO_744 (O_744,N_29409,N_29229);
xor UO_745 (O_745,N_26489,N_28259);
nor UO_746 (O_746,N_26094,N_28237);
nor UO_747 (O_747,N_27071,N_27099);
xnor UO_748 (O_748,N_24906,N_24950);
nor UO_749 (O_749,N_28459,N_24436);
nor UO_750 (O_750,N_28233,N_29322);
or UO_751 (O_751,N_24714,N_24066);
nand UO_752 (O_752,N_25777,N_26748);
xnor UO_753 (O_753,N_29975,N_27838);
xnor UO_754 (O_754,N_25643,N_24783);
and UO_755 (O_755,N_28919,N_27869);
nand UO_756 (O_756,N_25313,N_29185);
or UO_757 (O_757,N_29181,N_27479);
nor UO_758 (O_758,N_24785,N_25187);
or UO_759 (O_759,N_26867,N_26469);
nand UO_760 (O_760,N_24283,N_25340);
or UO_761 (O_761,N_26089,N_27504);
nor UO_762 (O_762,N_27680,N_25914);
or UO_763 (O_763,N_26510,N_29003);
nand UO_764 (O_764,N_26581,N_27278);
nor UO_765 (O_765,N_27326,N_25462);
and UO_766 (O_766,N_27478,N_27695);
and UO_767 (O_767,N_24418,N_26135);
nand UO_768 (O_768,N_28850,N_27902);
nor UO_769 (O_769,N_27182,N_28098);
nand UO_770 (O_770,N_25316,N_28933);
xor UO_771 (O_771,N_28462,N_25352);
nand UO_772 (O_772,N_25558,N_24055);
nor UO_773 (O_773,N_24178,N_26699);
xnor UO_774 (O_774,N_26441,N_26799);
and UO_775 (O_775,N_27225,N_29390);
or UO_776 (O_776,N_24222,N_24870);
xor UO_777 (O_777,N_25630,N_29111);
or UO_778 (O_778,N_25980,N_28009);
nand UO_779 (O_779,N_26732,N_29913);
or UO_780 (O_780,N_25214,N_26986);
and UO_781 (O_781,N_28357,N_24622);
nand UO_782 (O_782,N_29422,N_27705);
xor UO_783 (O_783,N_24522,N_27616);
xor UO_784 (O_784,N_29808,N_24403);
nor UO_785 (O_785,N_24571,N_25334);
nand UO_786 (O_786,N_25470,N_29410);
xnor UO_787 (O_787,N_26698,N_27212);
or UO_788 (O_788,N_24900,N_27089);
or UO_789 (O_789,N_24909,N_29616);
or UO_790 (O_790,N_26283,N_24491);
nor UO_791 (O_791,N_26247,N_24211);
nor UO_792 (O_792,N_29787,N_28359);
nor UO_793 (O_793,N_27415,N_25048);
xor UO_794 (O_794,N_27271,N_28244);
or UO_795 (O_795,N_28815,N_28157);
or UO_796 (O_796,N_28342,N_26805);
nand UO_797 (O_797,N_28407,N_26417);
nor UO_798 (O_798,N_27862,N_24668);
nand UO_799 (O_799,N_26405,N_27017);
and UO_800 (O_800,N_26853,N_28761);
nor UO_801 (O_801,N_28444,N_28880);
and UO_802 (O_802,N_26971,N_29495);
and UO_803 (O_803,N_26268,N_29330);
or UO_804 (O_804,N_27983,N_29482);
nor UO_805 (O_805,N_29317,N_27073);
or UO_806 (O_806,N_25725,N_27605);
xnor UO_807 (O_807,N_29717,N_26099);
nand UO_808 (O_808,N_26458,N_24715);
xor UO_809 (O_809,N_26981,N_26157);
nor UO_810 (O_810,N_26747,N_25866);
xor UO_811 (O_811,N_25543,N_28570);
nor UO_812 (O_812,N_25539,N_27158);
nor UO_813 (O_813,N_29518,N_26384);
or UO_814 (O_814,N_25747,N_29599);
nand UO_815 (O_815,N_26874,N_26004);
and UO_816 (O_816,N_24445,N_26462);
nor UO_817 (O_817,N_25027,N_25041);
or UO_818 (O_818,N_24359,N_24010);
xnor UO_819 (O_819,N_28231,N_28708);
or UO_820 (O_820,N_28363,N_25929);
or UO_821 (O_821,N_28258,N_25896);
nor UO_822 (O_822,N_25167,N_29110);
and UO_823 (O_823,N_24278,N_28271);
and UO_824 (O_824,N_25565,N_24639);
nor UO_825 (O_825,N_29745,N_25780);
and UO_826 (O_826,N_27386,N_27254);
nand UO_827 (O_827,N_28978,N_24846);
or UO_828 (O_828,N_24086,N_26130);
nor UO_829 (O_829,N_24809,N_27464);
nor UO_830 (O_830,N_27049,N_28994);
nor UO_831 (O_831,N_25333,N_27558);
or UO_832 (O_832,N_27673,N_24372);
nand UO_833 (O_833,N_27455,N_24708);
nor UO_834 (O_834,N_25627,N_27699);
nor UO_835 (O_835,N_29720,N_29194);
nand UO_836 (O_836,N_28559,N_26061);
nor UO_837 (O_837,N_29002,N_27883);
and UO_838 (O_838,N_26227,N_27757);
nor UO_839 (O_839,N_29554,N_24939);
xnor UO_840 (O_840,N_26881,N_24578);
xnor UO_841 (O_841,N_28027,N_25451);
nor UO_842 (O_842,N_24317,N_24021);
or UO_843 (O_843,N_28949,N_25647);
xor UO_844 (O_844,N_24036,N_27140);
xor UO_845 (O_845,N_29708,N_29824);
xor UO_846 (O_846,N_26188,N_26005);
nor UO_847 (O_847,N_29081,N_24725);
or UO_848 (O_848,N_27663,N_28038);
and UO_849 (O_849,N_26534,N_26713);
xor UO_850 (O_850,N_26662,N_27816);
or UO_851 (O_851,N_24759,N_27652);
xnor UO_852 (O_852,N_28799,N_26741);
nand UO_853 (O_853,N_28614,N_25407);
xor UO_854 (O_854,N_25939,N_26299);
and UO_855 (O_855,N_26181,N_27555);
xor UO_856 (O_856,N_28210,N_25745);
nand UO_857 (O_857,N_27893,N_24345);
nand UO_858 (O_858,N_28317,N_26694);
xnor UO_859 (O_859,N_29225,N_26626);
xor UO_860 (O_860,N_29252,N_24673);
or UO_861 (O_861,N_26914,N_26546);
xor UO_862 (O_862,N_29467,N_25507);
xnor UO_863 (O_863,N_27498,N_28785);
or UO_864 (O_864,N_25384,N_27638);
nand UO_865 (O_865,N_27601,N_26571);
nor UO_866 (O_866,N_29395,N_26113);
nand UO_867 (O_867,N_25438,N_25483);
and UO_868 (O_868,N_26073,N_28675);
nor UO_869 (O_869,N_26494,N_24268);
and UO_870 (O_870,N_25659,N_29528);
xor UO_871 (O_871,N_24088,N_27626);
xor UO_872 (O_872,N_28637,N_25030);
and UO_873 (O_873,N_24374,N_28961);
nor UO_874 (O_874,N_24623,N_27769);
nor UO_875 (O_875,N_27194,N_24058);
xnor UO_876 (O_876,N_29795,N_24801);
and UO_877 (O_877,N_27780,N_25127);
nor UO_878 (O_878,N_26664,N_24685);
xor UO_879 (O_879,N_26480,N_25877);
nor UO_880 (O_880,N_24724,N_28372);
nor UO_881 (O_881,N_26894,N_27173);
and UO_882 (O_882,N_24270,N_27240);
nor UO_883 (O_883,N_28811,N_26173);
xnor UO_884 (O_884,N_24540,N_29621);
or UO_885 (O_885,N_26924,N_28091);
nand UO_886 (O_886,N_26695,N_24631);
and UO_887 (O_887,N_29663,N_26048);
and UO_888 (O_888,N_24795,N_26006);
xor UO_889 (O_889,N_28416,N_29132);
xnor UO_890 (O_890,N_29477,N_25546);
nor UO_891 (O_891,N_27483,N_24358);
nand UO_892 (O_892,N_29978,N_24296);
xnor UO_893 (O_893,N_26789,N_28721);
nand UO_894 (O_894,N_26596,N_24879);
xor UO_895 (O_895,N_29595,N_25757);
and UO_896 (O_896,N_24004,N_26310);
or UO_897 (O_897,N_26677,N_25432);
or UO_898 (O_898,N_25339,N_25918);
and UO_899 (O_899,N_26682,N_29394);
nor UO_900 (O_900,N_24292,N_27482);
nor UO_901 (O_901,N_25626,N_29678);
nor UO_902 (O_902,N_29934,N_27463);
xnor UO_903 (O_903,N_24473,N_24239);
xor UO_904 (O_904,N_27832,N_28128);
nor UO_905 (O_905,N_24250,N_28064);
nand UO_906 (O_906,N_27775,N_26912);
and UO_907 (O_907,N_27629,N_29981);
xor UO_908 (O_908,N_25467,N_26956);
or UO_909 (O_909,N_25830,N_27421);
nor UO_910 (O_910,N_25191,N_27202);
xor UO_911 (O_911,N_28380,N_26710);
nand UO_912 (O_912,N_29965,N_28165);
or UO_913 (O_913,N_25153,N_26758);
nand UO_914 (O_914,N_26916,N_28120);
or UO_915 (O_915,N_25639,N_25687);
xor UO_916 (O_916,N_24750,N_25592);
xor UO_917 (O_917,N_25023,N_24856);
nand UO_918 (O_918,N_24777,N_28805);
nand UO_919 (O_919,N_26819,N_26857);
xor UO_920 (O_920,N_27951,N_29042);
nand UO_921 (O_921,N_26569,N_27078);
or UO_922 (O_922,N_28464,N_26500);
and UO_923 (O_923,N_29109,N_25336);
and UO_924 (O_924,N_29096,N_27020);
nor UO_925 (O_925,N_27590,N_26332);
nor UO_926 (O_926,N_27435,N_28175);
nand UO_927 (O_927,N_28426,N_24295);
xnor UO_928 (O_928,N_27700,N_27217);
nor UO_929 (O_929,N_29112,N_26050);
nor UO_930 (O_930,N_28513,N_27472);
or UO_931 (O_931,N_25032,N_29475);
nor UO_932 (O_932,N_29116,N_29961);
nand UO_933 (O_933,N_27032,N_26292);
nand UO_934 (O_934,N_27430,N_29671);
nand UO_935 (O_935,N_25820,N_29590);
nand UO_936 (O_936,N_26702,N_24134);
and UO_937 (O_937,N_24942,N_24974);
xnor UO_938 (O_938,N_25719,N_24395);
and UO_939 (O_939,N_25471,N_26634);
and UO_940 (O_940,N_26010,N_25112);
nor UO_941 (O_941,N_25791,N_24649);
and UO_942 (O_942,N_29502,N_28627);
nor UO_943 (O_943,N_29271,N_28609);
nor UO_944 (O_944,N_25008,N_26092);
or UO_945 (O_945,N_26231,N_25392);
nand UO_946 (O_946,N_25306,N_29227);
nor UO_947 (O_947,N_25993,N_26440);
or UO_948 (O_948,N_25349,N_25250);
and UO_949 (O_949,N_29687,N_28077);
and UO_950 (O_950,N_29645,N_24577);
and UO_951 (O_951,N_25530,N_25910);
nor UO_952 (O_952,N_27941,N_25974);
nor UO_953 (O_953,N_27510,N_25003);
nand UO_954 (O_954,N_25045,N_25670);
nand UO_955 (O_955,N_24831,N_27276);
nand UO_956 (O_956,N_24423,N_27401);
xor UO_957 (O_957,N_24624,N_29241);
xnor UO_958 (O_958,N_24860,N_28515);
and UO_959 (O_959,N_26980,N_29928);
or UO_960 (O_960,N_25144,N_28029);
xnor UO_961 (O_961,N_24349,N_24409);
nand UO_962 (O_962,N_26047,N_28854);
nor UO_963 (O_963,N_25589,N_27978);
nor UO_964 (O_964,N_27065,N_26767);
nand UO_965 (O_965,N_29033,N_28909);
or UO_966 (O_966,N_29052,N_25807);
nor UO_967 (O_967,N_24766,N_24892);
xnor UO_968 (O_968,N_24344,N_27190);
nand UO_969 (O_969,N_29125,N_24440);
xnor UO_970 (O_970,N_26839,N_24660);
xnor UO_971 (O_971,N_28218,N_29641);
xnor UO_972 (O_972,N_28747,N_26795);
nor UO_973 (O_973,N_26922,N_26511);
and UO_974 (O_974,N_29918,N_27402);
and UO_975 (O_975,N_26529,N_25886);
and UO_976 (O_976,N_29877,N_28595);
nor UO_977 (O_977,N_24754,N_27389);
xnor UO_978 (O_978,N_29973,N_29683);
nor UO_979 (O_979,N_29103,N_29894);
nand UO_980 (O_980,N_28833,N_26574);
nor UO_981 (O_981,N_26873,N_26430);
nor UO_982 (O_982,N_26087,N_28603);
or UO_983 (O_983,N_28903,N_28838);
xnor UO_984 (O_984,N_26756,N_28643);
nand UO_985 (O_985,N_25731,N_29091);
nor UO_986 (O_986,N_27085,N_24546);
nand UO_987 (O_987,N_28207,N_24318);
nand UO_988 (O_988,N_28249,N_27717);
nor UO_989 (O_989,N_24041,N_24771);
nand UO_990 (O_990,N_24286,N_28989);
nand UO_991 (O_991,N_25234,N_25184);
xor UO_992 (O_992,N_24910,N_25722);
or UO_993 (O_993,N_27721,N_29501);
xor UO_994 (O_994,N_25236,N_27516);
xor UO_995 (O_995,N_25300,N_29149);
or UO_996 (O_996,N_26800,N_29341);
nand UO_997 (O_997,N_26476,N_25318);
nor UO_998 (O_998,N_26564,N_27992);
and UO_999 (O_999,N_29463,N_25020);
and UO_1000 (O_1000,N_25948,N_28869);
and UO_1001 (O_1001,N_29586,N_24192);
xnor UO_1002 (O_1002,N_29685,N_29161);
or UO_1003 (O_1003,N_28621,N_24415);
or UO_1004 (O_1004,N_28543,N_29967);
or UO_1005 (O_1005,N_26761,N_28232);
xor UO_1006 (O_1006,N_24755,N_29614);
or UO_1007 (O_1007,N_29084,N_26931);
nor UO_1008 (O_1008,N_26964,N_29553);
or UO_1009 (O_1009,N_24586,N_24642);
and UO_1010 (O_1010,N_27872,N_27518);
nand UO_1011 (O_1011,N_24003,N_26102);
xnor UO_1012 (O_1012,N_27468,N_28431);
or UO_1013 (O_1013,N_25431,N_24327);
xor UO_1014 (O_1014,N_27815,N_27784);
and UO_1015 (O_1015,N_26208,N_25535);
nor UO_1016 (O_1016,N_27069,N_26681);
nand UO_1017 (O_1017,N_25243,N_27588);
and UO_1018 (O_1018,N_28136,N_28905);
or UO_1019 (O_1019,N_25657,N_25635);
xnor UO_1020 (O_1020,N_26370,N_28830);
xnor UO_1021 (O_1021,N_29633,N_24670);
xor UO_1022 (O_1022,N_26074,N_25622);
nor UO_1023 (O_1023,N_28146,N_27583);
or UO_1024 (O_1024,N_25838,N_24799);
and UO_1025 (O_1025,N_26642,N_25245);
nand UO_1026 (O_1026,N_27164,N_28965);
or UO_1027 (O_1027,N_25281,N_26901);
or UO_1028 (O_1028,N_24871,N_25390);
nand UO_1029 (O_1029,N_29893,N_27341);
xor UO_1030 (O_1030,N_26831,N_24821);
xor UO_1031 (O_1031,N_24424,N_24187);
nand UO_1032 (O_1032,N_26472,N_27665);
or UO_1033 (O_1033,N_27692,N_29803);
or UO_1034 (O_1034,N_29786,N_24341);
or UO_1035 (O_1035,N_28631,N_25156);
nor UO_1036 (O_1036,N_25136,N_25162);
nor UO_1037 (O_1037,N_24121,N_27643);
or UO_1038 (O_1038,N_26473,N_29759);
nor UO_1039 (O_1039,N_26137,N_24661);
xnor UO_1040 (O_1040,N_24406,N_29162);
or UO_1041 (O_1041,N_27142,N_24163);
xor UO_1042 (O_1042,N_26293,N_29899);
or UO_1043 (O_1043,N_27625,N_28012);
and UO_1044 (O_1044,N_28307,N_28780);
or UO_1045 (O_1045,N_25970,N_28045);
and UO_1046 (O_1046,N_25069,N_28723);
nor UO_1047 (O_1047,N_26727,N_25385);
xnor UO_1048 (O_1048,N_24316,N_27087);
or UO_1049 (O_1049,N_25283,N_25097);
xor UO_1050 (O_1050,N_24471,N_27197);
nand UO_1051 (O_1051,N_28856,N_28608);
and UO_1052 (O_1052,N_28715,N_28396);
nor UO_1053 (O_1053,N_26085,N_26246);
xor UO_1054 (O_1054,N_28150,N_25682);
nand UO_1055 (O_1055,N_24588,N_26835);
or UO_1056 (O_1056,N_28516,N_25107);
or UO_1057 (O_1057,N_25895,N_27072);
nand UO_1058 (O_1058,N_27357,N_29494);
or UO_1059 (O_1059,N_25039,N_28858);
and UO_1060 (O_1060,N_27097,N_26728);
xnor UO_1061 (O_1061,N_26275,N_27338);
xor UO_1062 (O_1062,N_26169,N_29045);
and UO_1063 (O_1063,N_25360,N_25650);
or UO_1064 (O_1064,N_26021,N_26621);
nand UO_1065 (O_1065,N_28335,N_24231);
and UO_1066 (O_1066,N_27859,N_29253);
and UO_1067 (O_1067,N_29329,N_26124);
nand UO_1068 (O_1068,N_25185,N_29017);
or UO_1069 (O_1069,N_29373,N_27666);
and UO_1070 (O_1070,N_28294,N_24769);
xor UO_1071 (O_1071,N_28454,N_29996);
nand UO_1072 (O_1072,N_27337,N_26174);
nand UO_1073 (O_1073,N_27247,N_26057);
or UO_1074 (O_1074,N_28229,N_25468);
nand UO_1075 (O_1075,N_26235,N_29911);
and UO_1076 (O_1076,N_27310,N_27289);
or UO_1077 (O_1077,N_24469,N_26314);
and UO_1078 (O_1078,N_28130,N_25845);
xor UO_1079 (O_1079,N_26892,N_28264);
or UO_1080 (O_1080,N_26562,N_29243);
nand UO_1081 (O_1081,N_29060,N_26380);
and UO_1082 (O_1082,N_26345,N_27067);
nor UO_1083 (O_1083,N_28844,N_27754);
and UO_1084 (O_1084,N_25556,N_28436);
or UO_1085 (O_1085,N_24340,N_27044);
or UO_1086 (O_1086,N_24617,N_24945);
xnor UO_1087 (O_1087,N_24241,N_28468);
and UO_1088 (O_1088,N_28572,N_28296);
or UO_1089 (O_1089,N_25024,N_27703);
xnor UO_1090 (O_1090,N_24965,N_25476);
and UO_1091 (O_1091,N_25337,N_25154);
or UO_1092 (O_1092,N_24806,N_26811);
nand UO_1093 (O_1093,N_29370,N_26442);
nand UO_1094 (O_1094,N_24646,N_27508);
nor UO_1095 (O_1095,N_25808,N_26207);
or UO_1096 (O_1096,N_25967,N_26025);
nor UO_1097 (O_1097,N_28738,N_29455);
nand UO_1098 (O_1098,N_27999,N_29565);
nand UO_1099 (O_1099,N_24710,N_28573);
and UO_1100 (O_1100,N_24220,N_28711);
and UO_1101 (O_1101,N_29941,N_27058);
nand UO_1102 (O_1102,N_28656,N_28255);
xnor UO_1103 (O_1103,N_25270,N_24037);
and UO_1104 (O_1104,N_25176,N_25498);
nand UO_1105 (O_1105,N_27676,N_27364);
xor UO_1106 (O_1106,N_25408,N_29858);
nand UO_1107 (O_1107,N_29027,N_29355);
or UO_1108 (O_1108,N_26104,N_29376);
and UO_1109 (O_1109,N_26842,N_24103);
or UO_1110 (O_1110,N_26279,N_24079);
or UO_1111 (O_1111,N_27871,N_27329);
and UO_1112 (O_1112,N_24308,N_25362);
nand UO_1113 (O_1113,N_26468,N_26059);
nor UO_1114 (O_1114,N_27291,N_24154);
xnor UO_1115 (O_1115,N_24490,N_27373);
xor UO_1116 (O_1116,N_27132,N_25157);
and UO_1117 (O_1117,N_29270,N_29480);
xnor UO_1118 (O_1118,N_28106,N_29659);
xnor UO_1119 (O_1119,N_25058,N_29291);
or UO_1120 (O_1120,N_26479,N_25553);
nor UO_1121 (O_1121,N_29193,N_25389);
nor UO_1122 (O_1122,N_28293,N_29471);
xnor UO_1123 (O_1123,N_26525,N_28579);
or UO_1124 (O_1124,N_28227,N_28793);
nand UO_1125 (O_1125,N_28174,N_25688);
nor UO_1126 (O_1126,N_29256,N_26251);
nor UO_1127 (O_1127,N_28834,N_25952);
or UO_1128 (O_1128,N_24276,N_25063);
nand UO_1129 (O_1129,N_29784,N_28975);
and UO_1130 (O_1130,N_26416,N_24198);
xnor UO_1131 (O_1131,N_24876,N_24499);
nor UO_1132 (O_1132,N_25801,N_29959);
xnor UO_1133 (O_1133,N_26219,N_27005);
nor UO_1134 (O_1134,N_25658,N_29302);
and UO_1135 (O_1135,N_27512,N_26938);
xor UO_1136 (O_1136,N_26492,N_28395);
nor UO_1137 (O_1137,N_25926,N_27036);
nand UO_1138 (O_1138,N_29191,N_27474);
and UO_1139 (O_1139,N_24201,N_26105);
xnor UO_1140 (O_1140,N_24864,N_27567);
xnor UO_1141 (O_1141,N_26375,N_24123);
xor UO_1142 (O_1142,N_26523,N_27544);
xor UO_1143 (O_1143,N_25202,N_27696);
xnor UO_1144 (O_1144,N_25555,N_26342);
and UO_1145 (O_1145,N_28308,N_24129);
nor UO_1146 (O_1146,N_27686,N_24599);
or UO_1147 (O_1147,N_27220,N_27850);
or UO_1148 (O_1148,N_28510,N_27904);
nand UO_1149 (O_1149,N_26226,N_27393);
nand UO_1150 (O_1150,N_26387,N_28247);
and UO_1151 (O_1151,N_25143,N_28696);
xnor UO_1152 (O_1152,N_24092,N_24608);
xor UO_1153 (O_1153,N_26443,N_26678);
nor UO_1154 (O_1154,N_24561,N_26383);
nand UO_1155 (O_1155,N_29040,N_27609);
and UO_1156 (O_1156,N_24770,N_28311);
nor UO_1157 (O_1157,N_25173,N_27403);
and UO_1158 (O_1158,N_27568,N_28325);
or UO_1159 (O_1159,N_29531,N_24311);
nand UO_1160 (O_1160,N_24898,N_24800);
and UO_1161 (O_1161,N_28825,N_27566);
xnor UO_1162 (O_1162,N_25105,N_29374);
xnor UO_1163 (O_1163,N_24375,N_29930);
xor UO_1164 (O_1164,N_25554,N_27670);
nand UO_1165 (O_1165,N_29147,N_29923);
nor UO_1166 (O_1166,N_27564,N_24704);
xnor UO_1167 (O_1167,N_28718,N_26858);
or UO_1168 (O_1168,N_25911,N_28378);
or UO_1169 (O_1169,N_27539,N_27094);
nor UO_1170 (O_1170,N_25538,N_25212);
nand UO_1171 (O_1171,N_27603,N_25422);
or UO_1172 (O_1172,N_26487,N_27494);
and UO_1173 (O_1173,N_25274,N_24232);
nor UO_1174 (O_1174,N_25198,N_24496);
nand UO_1175 (O_1175,N_29589,N_28546);
xnor UO_1176 (O_1176,N_24527,N_25417);
and UO_1177 (O_1177,N_26657,N_27536);
xor UO_1178 (O_1178,N_27294,N_25205);
and UO_1179 (O_1179,N_25515,N_25551);
nor UO_1180 (O_1180,N_24807,N_27153);
xnor UO_1181 (O_1181,N_29007,N_28137);
or UO_1182 (O_1182,N_28751,N_28222);
nand UO_1183 (O_1183,N_26081,N_26357);
nand UO_1184 (O_1184,N_29389,N_25863);
and UO_1185 (O_1185,N_27726,N_28755);
nor UO_1186 (O_1186,N_28896,N_27224);
or UO_1187 (O_1187,N_26604,N_25846);
or UO_1188 (O_1188,N_28596,N_27651);
and UO_1189 (O_1189,N_28245,N_24339);
xor UO_1190 (O_1190,N_25289,N_29878);
and UO_1191 (O_1191,N_26336,N_29257);
and UO_1192 (O_1192,N_29705,N_26533);
and UO_1193 (O_1193,N_25192,N_25946);
xnor UO_1194 (O_1194,N_24493,N_28692);
nor UO_1195 (O_1195,N_27187,N_24106);
and UO_1196 (O_1196,N_27907,N_24485);
xnor UO_1197 (O_1197,N_27822,N_24142);
or UO_1198 (O_1198,N_29630,N_27785);
or UO_1199 (O_1199,N_25160,N_24541);
xnor UO_1200 (O_1200,N_25695,N_29525);
or UO_1201 (O_1201,N_24149,N_25007);
or UO_1202 (O_1202,N_26420,N_27848);
and UO_1203 (O_1203,N_29864,N_24537);
and UO_1204 (O_1204,N_24413,N_29266);
nand UO_1205 (O_1205,N_27242,N_25703);
nand UO_1206 (O_1206,N_25475,N_25718);
nand UO_1207 (O_1207,N_25654,N_26199);
nor UO_1208 (O_1208,N_24050,N_26646);
or UO_1209 (O_1209,N_25668,N_25310);
xnor UO_1210 (O_1210,N_25197,N_25317);
or UO_1211 (O_1211,N_25735,N_27014);
and UO_1212 (O_1212,N_24360,N_26281);
nor UO_1213 (O_1213,N_24376,N_24828);
nor UO_1214 (O_1214,N_29289,N_25709);
nor UO_1215 (O_1215,N_25545,N_24109);
or UO_1216 (O_1216,N_25085,N_25258);
nand UO_1217 (O_1217,N_24837,N_28932);
and UO_1218 (O_1218,N_28828,N_27367);
nand UO_1219 (O_1219,N_26880,N_29377);
xor UO_1220 (O_1220,N_29882,N_26653);
and UO_1221 (O_1221,N_24343,N_27104);
nor UO_1222 (O_1222,N_29061,N_26882);
nand UO_1223 (O_1223,N_28283,N_28195);
nand UO_1224 (O_1224,N_26961,N_27737);
and UO_1225 (O_1225,N_26797,N_26660);
or UO_1226 (O_1226,N_24901,N_27836);
nor UO_1227 (O_1227,N_24633,N_28843);
and UO_1228 (O_1228,N_28435,N_26750);
and UO_1229 (O_1229,N_29148,N_25484);
nor UO_1230 (O_1230,N_27063,N_25239);
and UO_1231 (O_1231,N_29719,N_27761);
and UO_1232 (O_1232,N_25862,N_24025);
or UO_1233 (O_1233,N_26304,N_29880);
and UO_1234 (O_1234,N_25130,N_29005);
nor UO_1235 (O_1235,N_27593,N_24819);
and UO_1236 (O_1236,N_24753,N_24585);
or UO_1237 (O_1237,N_27443,N_28660);
nand UO_1238 (O_1238,N_24321,N_29513);
and UO_1239 (O_1239,N_27449,N_25795);
xnor UO_1240 (O_1240,N_26229,N_28474);
or UO_1241 (O_1241,N_27141,N_25730);
nor UO_1242 (O_1242,N_24435,N_26743);
and UO_1243 (O_1243,N_24285,N_26947);
xor UO_1244 (O_1244,N_24967,N_24810);
nand UO_1245 (O_1245,N_28182,N_25758);
xor UO_1246 (O_1246,N_26329,N_25131);
or UO_1247 (O_1247,N_26165,N_25821);
or UO_1248 (O_1248,N_25031,N_28731);
or UO_1249 (O_1249,N_26391,N_28263);
or UO_1250 (O_1250,N_27473,N_24322);
xnor UO_1251 (O_1251,N_28999,N_28219);
or UO_1252 (O_1252,N_26334,N_29915);
or UO_1253 (O_1253,N_27199,N_24552);
or UO_1254 (O_1254,N_27937,N_26063);
or UO_1255 (O_1255,N_26736,N_27096);
nor UO_1256 (O_1256,N_24057,N_26321);
nand UO_1257 (O_1257,N_28845,N_26248);
nor UO_1258 (O_1258,N_28792,N_29117);
nor UO_1259 (O_1259,N_25017,N_25095);
xor UO_1260 (O_1260,N_27122,N_28948);
or UO_1261 (O_1261,N_24398,N_27453);
and UO_1262 (O_1262,N_27738,N_24074);
nand UO_1263 (O_1263,N_25814,N_27576);
xnor UO_1264 (O_1264,N_29391,N_29164);
nand UO_1265 (O_1265,N_28534,N_24929);
nor UO_1266 (O_1266,N_25738,N_25522);
or UO_1267 (O_1267,N_25455,N_27234);
xor UO_1268 (O_1268,N_26155,N_29115);
and UO_1269 (O_1269,N_27425,N_27441);
nor UO_1270 (O_1270,N_27554,N_25423);
or UO_1271 (O_1271,N_26918,N_27615);
xnor UO_1272 (O_1272,N_27720,N_25054);
xor UO_1273 (O_1273,N_29639,N_26933);
or UO_1274 (O_1274,N_26988,N_29049);
nor UO_1275 (O_1275,N_26451,N_27334);
or UO_1276 (O_1276,N_24396,N_27176);
nand UO_1277 (O_1277,N_29695,N_29626);
nand UO_1278 (O_1278,N_27722,N_26069);
nor UO_1279 (O_1279,N_29998,N_28163);
or UO_1280 (O_1280,N_27578,N_26343);
nand UO_1281 (O_1281,N_29993,N_26554);
nand UO_1282 (O_1282,N_27408,N_28758);
nor UO_1283 (O_1283,N_29474,N_26921);
nor UO_1284 (O_1284,N_28787,N_26138);
and UO_1285 (O_1285,N_29481,N_24125);
or UO_1286 (O_1286,N_24183,N_24439);
xor UO_1287 (O_1287,N_28292,N_25499);
nand UO_1288 (O_1288,N_24570,N_26904);
and UO_1289 (O_1289,N_24858,N_24553);
nor UO_1290 (O_1290,N_28320,N_28749);
and UO_1291 (O_1291,N_28310,N_29994);
xnor UO_1292 (O_1292,N_27292,N_26538);
or UO_1293 (O_1293,N_27704,N_25215);
and UO_1294 (O_1294,N_27370,N_29336);
or UO_1295 (O_1295,N_28929,N_26250);
or UO_1296 (O_1296,N_27345,N_28824);
nor UO_1297 (O_1297,N_27033,N_29718);
xnor UO_1298 (O_1298,N_28103,N_25204);
and UO_1299 (O_1299,N_25247,N_24348);
or UO_1300 (O_1300,N_27660,N_29293);
nand UO_1301 (O_1301,N_29567,N_29722);
xor UO_1302 (O_1302,N_24635,N_25241);
xnor UO_1303 (O_1303,N_27556,N_27547);
and UO_1304 (O_1304,N_29418,N_29141);
and UO_1305 (O_1305,N_25633,N_27206);
nand UO_1306 (O_1306,N_25053,N_27879);
xor UO_1307 (O_1307,N_26178,N_24219);
xnor UO_1308 (O_1308,N_24648,N_24474);
xor UO_1309 (O_1309,N_25350,N_27343);
nor UO_1310 (O_1310,N_27339,N_25096);
xnor UO_1311 (O_1311,N_29158,N_29503);
xor UO_1312 (O_1312,N_28982,N_29077);
nand UO_1313 (O_1313,N_25071,N_28549);
xor UO_1314 (O_1314,N_28667,N_25893);
and UO_1315 (O_1315,N_24636,N_26466);
nand UO_1316 (O_1316,N_28754,N_29452);
nor UO_1317 (O_1317,N_28884,N_26017);
xnor UO_1318 (O_1318,N_29948,N_24271);
or UO_1319 (O_1319,N_25921,N_29094);
xnor UO_1320 (O_1320,N_27889,N_25170);
and UO_1321 (O_1321,N_27308,N_28560);
nor UO_1322 (O_1322,N_26704,N_29860);
and UO_1323 (O_1323,N_25224,N_24138);
nand UO_1324 (O_1324,N_26163,N_29951);
or UO_1325 (O_1325,N_24210,N_25405);
nand UO_1326 (O_1326,N_24912,N_28168);
or UO_1327 (O_1327,N_25999,N_26090);
nor UO_1328 (O_1328,N_27091,N_29327);
xnor UO_1329 (O_1329,N_29454,N_25147);
or UO_1330 (O_1330,N_25968,N_24238);
or UO_1331 (O_1331,N_25218,N_29167);
nor UO_1332 (O_1332,N_27079,N_26372);
nor UO_1333 (O_1333,N_24618,N_29783);
xnor UO_1334 (O_1334,N_29240,N_26776);
nor UO_1335 (O_1335,N_28522,N_27597);
nand UO_1336 (O_1336,N_26427,N_29617);
or UO_1337 (O_1337,N_28016,N_26703);
nor UO_1338 (O_1338,N_25047,N_25943);
nor UO_1339 (O_1339,N_27496,N_28057);
nor UO_1340 (O_1340,N_25649,N_28646);
xor UO_1341 (O_1341,N_25453,N_28116);
or UO_1342 (O_1342,N_27621,N_26828);
or UO_1343 (O_1343,N_28170,N_26997);
nand UO_1344 (O_1344,N_24836,N_24692);
nor UO_1345 (O_1345,N_27579,N_25450);
xor UO_1346 (O_1346,N_24868,N_24873);
or UO_1347 (O_1347,N_28937,N_29536);
nor UO_1348 (O_1348,N_27804,N_29729);
nor UO_1349 (O_1349,N_26108,N_25013);
or UO_1350 (O_1350,N_25834,N_24516);
nor UO_1351 (O_1351,N_29679,N_29404);
xnor UO_1352 (O_1352,N_28100,N_25677);
nand UO_1353 (O_1353,N_26650,N_28337);
nand UO_1354 (O_1354,N_28381,N_25084);
or UO_1355 (O_1355,N_27340,N_26252);
and UO_1356 (O_1356,N_29844,N_27250);
xor UO_1357 (O_1357,N_28350,N_27129);
xnor UO_1358 (O_1358,N_27290,N_24166);
or UO_1359 (O_1359,N_24158,N_25798);
nand UO_1360 (O_1360,N_24001,N_24273);
nand UO_1361 (O_1361,N_27863,N_28160);
xor UO_1362 (O_1362,N_29306,N_28700);
nor UO_1363 (O_1363,N_26690,N_29835);
xor UO_1364 (O_1364,N_29665,N_29661);
nand UO_1365 (O_1365,N_24997,N_28566);
and UO_1366 (O_1366,N_28767,N_28683);
nand UO_1367 (O_1367,N_28930,N_29955);
or UO_1368 (O_1368,N_28506,N_29242);
xor UO_1369 (O_1369,N_29220,N_25345);
and UO_1370 (O_1370,N_24512,N_29576);
nor UO_1371 (O_1371,N_27093,N_29288);
or UO_1372 (O_1372,N_25836,N_25675);
and UO_1373 (O_1373,N_25338,N_26437);
or UO_1374 (O_1374,N_26457,N_26396);
xnor UO_1375 (O_1375,N_24822,N_24256);
and UO_1376 (O_1376,N_24262,N_29215);
xnor UO_1377 (O_1377,N_29830,N_29210);
xnor UO_1378 (O_1378,N_28479,N_25348);
and UO_1379 (O_1379,N_24090,N_29439);
nor UO_1380 (O_1380,N_27115,N_24689);
nand UO_1381 (O_1381,N_28063,N_26192);
and UO_1382 (O_1382,N_28526,N_27163);
nor UO_1383 (O_1383,N_25513,N_26749);
and UO_1384 (O_1384,N_27458,N_24133);
nor UO_1385 (O_1385,N_25599,N_24717);
nand UO_1386 (O_1386,N_25817,N_24189);
nor UO_1387 (O_1387,N_29751,N_28447);
xor UO_1388 (O_1388,N_29772,N_29264);
nand UO_1389 (O_1389,N_26151,N_25404);
and UO_1390 (O_1390,N_24038,N_29504);
nand UO_1391 (O_1391,N_29449,N_26906);
nand UO_1392 (O_1392,N_25873,N_29335);
xnor UO_1393 (O_1393,N_28145,N_29700);
nor UO_1394 (O_1394,N_25014,N_25727);
xor UO_1395 (O_1395,N_26770,N_26256);
or UO_1396 (O_1396,N_24659,N_27740);
nor UO_1397 (O_1397,N_26611,N_27436);
xnor UO_1398 (O_1398,N_24664,N_27944);
or UO_1399 (O_1399,N_25827,N_24794);
nor UO_1400 (O_1400,N_25025,N_29127);
or UO_1401 (O_1401,N_26167,N_28096);
nor UO_1402 (O_1402,N_26512,N_29952);
nand UO_1403 (O_1403,N_24662,N_27382);
or UO_1404 (O_1404,N_28164,N_27632);
nor UO_1405 (O_1405,N_24146,N_27226);
or UO_1406 (O_1406,N_24475,N_24259);
xnor UO_1407 (O_1407,N_25891,N_29505);
and UO_1408 (O_1408,N_26865,N_27054);
nor UO_1409 (O_1409,N_25026,N_26952);
nor UO_1410 (O_1410,N_26326,N_25729);
and UO_1411 (O_1411,N_29627,N_26771);
nand UO_1412 (O_1412,N_27667,N_26982);
or UO_1413 (O_1413,N_25315,N_26972);
nor UO_1414 (O_1414,N_27042,N_24513);
nand UO_1415 (O_1415,N_25284,N_25200);
and UO_1416 (O_1416,N_29704,N_28783);
nor UO_1417 (O_1417,N_25667,N_29904);
nor UO_1418 (O_1418,N_25913,N_24253);
nor UO_1419 (O_1419,N_27000,N_24179);
xnor UO_1420 (O_1420,N_26945,N_27284);
nor UO_1421 (O_1421,N_24719,N_24176);
and UO_1422 (O_1422,N_24745,N_28370);
xnor UO_1423 (O_1423,N_28302,N_29488);
or UO_1424 (O_1424,N_28276,N_28707);
and UO_1425 (O_1425,N_27313,N_27817);
and UO_1426 (O_1426,N_28086,N_26422);
xor UO_1427 (O_1427,N_28470,N_28862);
nor UO_1428 (O_1428,N_24690,N_27385);
nor UO_1429 (O_1429,N_27486,N_28652);
nand UO_1430 (O_1430,N_26365,N_25925);
or UO_1431 (O_1431,N_26670,N_25882);
xnor UO_1432 (O_1432,N_29667,N_26934);
and UO_1433 (O_1433,N_25732,N_27286);
and UO_1434 (O_1434,N_25828,N_24911);
and UO_1435 (O_1435,N_26813,N_28502);
or UO_1436 (O_1436,N_24567,N_25298);
and UO_1437 (O_1437,N_24905,N_27162);
xnor UO_1438 (O_1438,N_28877,N_28109);
nand UO_1439 (O_1439,N_25263,N_28113);
nor UO_1440 (O_1440,N_26502,N_27255);
or UO_1441 (O_1441,N_29059,N_25051);
xnor UO_1442 (O_1442,N_24242,N_29867);
and UO_1443 (O_1443,N_26561,N_28456);
nor UO_1444 (O_1444,N_27890,N_27145);
and UO_1445 (O_1445,N_25822,N_27925);
xor UO_1446 (O_1446,N_24095,N_27327);
xor UO_1447 (O_1447,N_24606,N_26962);
and UO_1448 (O_1448,N_28176,N_29715);
xnor UO_1449 (O_1449,N_26306,N_25488);
or UO_1450 (O_1450,N_28072,N_26153);
and UO_1451 (O_1451,N_24350,N_24140);
nor UO_1452 (O_1452,N_29690,N_24973);
nor UO_1453 (O_1453,N_28093,N_24212);
nor UO_1454 (O_1454,N_26645,N_29189);
and UO_1455 (O_1455,N_28031,N_29561);
nor UO_1456 (O_1456,N_24016,N_25712);
or UO_1457 (O_1457,N_24234,N_28576);
nor UO_1458 (O_1458,N_25855,N_29527);
xnor UO_1459 (O_1459,N_28001,N_25485);
xnor UO_1460 (O_1460,N_25221,N_25761);
or UO_1461 (O_1461,N_28520,N_24869);
nand UO_1462 (O_1462,N_29174,N_26801);
or UO_1463 (O_1463,N_27910,N_29594);
xnor UO_1464 (O_1464,N_28389,N_24507);
nand UO_1465 (O_1465,N_26143,N_28226);
and UO_1466 (O_1466,N_29999,N_27193);
nand UO_1467 (O_1467,N_25480,N_27116);
xor UO_1468 (O_1468,N_28809,N_26464);
or UO_1469 (O_1469,N_28642,N_28495);
or UO_1470 (O_1470,N_29269,N_28907);
nor UO_1471 (O_1471,N_26588,N_29300);
or UO_1472 (O_1472,N_26639,N_26062);
or UO_1473 (O_1473,N_25076,N_26790);
xor UO_1474 (O_1474,N_24147,N_25531);
and UO_1475 (O_1475,N_29382,N_26625);
or UO_1476 (O_1476,N_25398,N_25000);
and UO_1477 (O_1477,N_25033,N_25984);
xnor UO_1478 (O_1478,N_29865,N_29724);
nor UO_1479 (O_1479,N_27790,N_29615);
and UO_1480 (O_1480,N_24184,N_26697);
nand UO_1481 (O_1481,N_27577,N_25134);
or UO_1482 (O_1482,N_26589,N_29192);
or UO_1483 (O_1483,N_26110,N_24538);
xnor UO_1484 (O_1484,N_27418,N_24422);
xnor UO_1485 (O_1485,N_29073,N_28684);
xnor UO_1486 (O_1486,N_26285,N_25953);
and UO_1487 (O_1487,N_26309,N_25990);
and UO_1488 (O_1488,N_27082,N_26294);
and UO_1489 (O_1489,N_28986,N_28569);
and UO_1490 (O_1490,N_25037,N_25109);
xnor UO_1491 (O_1491,N_27839,N_24102);
nor UO_1492 (O_1492,N_29447,N_24332);
nor UO_1493 (O_1493,N_25805,N_27248);
nor UO_1494 (O_1494,N_29831,N_28584);
nand UO_1495 (O_1495,N_29024,N_28577);
xor UO_1496 (O_1496,N_24137,N_29165);
and UO_1497 (O_1497,N_27047,N_27209);
and UO_1498 (O_1498,N_24680,N_29907);
nor UO_1499 (O_1499,N_28189,N_25685);
nor UO_1500 (O_1500,N_27716,N_25449);
nand UO_1501 (O_1501,N_25503,N_24150);
nor UO_1502 (O_1502,N_28860,N_25124);
and UO_1503 (O_1503,N_27314,N_24122);
and UO_1504 (O_1504,N_28191,N_25557);
xnor UO_1505 (O_1505,N_29737,N_24096);
and UO_1506 (O_1506,N_26648,N_24267);
xor UO_1507 (O_1507,N_27318,N_24707);
nand UO_1508 (O_1508,N_27527,N_27312);
or UO_1509 (O_1509,N_27988,N_26146);
nor UO_1510 (O_1510,N_24990,N_28039);
and UO_1511 (O_1511,N_25248,N_26211);
nand UO_1512 (O_1512,N_25949,N_26001);
and UO_1513 (O_1513,N_28772,N_24788);
and UO_1514 (O_1514,N_24180,N_29721);
nand UO_1515 (O_1515,N_26297,N_24933);
nand UO_1516 (O_1516,N_29800,N_29244);
and UO_1517 (O_1517,N_24430,N_25374);
and UO_1518 (O_1518,N_26488,N_25305);
nand UO_1519 (O_1519,N_27031,N_29762);
or UO_1520 (O_1520,N_25723,N_28645);
nand UO_1521 (O_1521,N_24006,N_29540);
and UO_1522 (O_1522,N_28717,N_28602);
xnor UO_1523 (O_1523,N_26311,N_26607);
nor UO_1524 (O_1524,N_25819,N_27598);
nor UO_1525 (O_1525,N_27896,N_28868);
nor UO_1526 (O_1526,N_28629,N_25837);
and UO_1527 (O_1527,N_27384,N_25615);
or UO_1528 (O_1528,N_24986,N_27701);
nor UO_1529 (O_1529,N_27330,N_26716);
xor UO_1530 (O_1530,N_24043,N_28272);
xor UO_1531 (O_1531,N_25099,N_24603);
or UO_1532 (O_1532,N_26223,N_25601);
and UO_1533 (O_1533,N_25052,N_28842);
or UO_1534 (O_1534,N_24402,N_27806);
or UO_1535 (O_1535,N_28678,N_26791);
nor UO_1536 (O_1536,N_28155,N_28466);
nor UO_1537 (O_1537,N_29369,N_28786);
nand UO_1538 (O_1538,N_24731,N_29949);
nand UO_1539 (O_1539,N_25254,N_28030);
and UO_1540 (O_1540,N_29407,N_28742);
and UO_1541 (O_1541,N_26386,N_28753);
nand UO_1542 (O_1542,N_28300,N_28525);
nor UO_1543 (O_1543,N_24762,N_24999);
nand UO_1544 (O_1544,N_29733,N_28482);
nor UO_1545 (O_1545,N_28874,N_26821);
xor UO_1546 (O_1546,N_29649,N_24619);
or UO_1547 (O_1547,N_29921,N_28035);
nand UO_1548 (O_1548,N_24523,N_28374);
or UO_1549 (O_1549,N_25132,N_25899);
or UO_1550 (O_1550,N_27269,N_26656);
nand UO_1551 (O_1551,N_27538,N_26034);
nor UO_1552 (O_1552,N_26497,N_24542);
xor UO_1553 (O_1553,N_27411,N_27347);
and UO_1554 (O_1554,N_27914,N_25954);
or UO_1555 (O_1555,N_28415,N_24255);
or UO_1556 (O_1556,N_28489,N_24568);
nor UO_1557 (O_1557,N_26994,N_28998);
or UO_1558 (O_1558,N_29684,N_29436);
xnor UO_1559 (O_1559,N_28034,N_24248);
nor UO_1560 (O_1560,N_26026,N_25344);
nor UO_1561 (O_1561,N_26037,N_26794);
nor UO_1562 (O_1562,N_27921,N_26616);
or UO_1563 (O_1563,N_25552,N_26966);
and UO_1564 (O_1564,N_24023,N_27846);
and UO_1565 (O_1565,N_24387,N_28610);
nor UO_1566 (O_1566,N_25121,N_27233);
and UO_1567 (O_1567,N_27529,N_28002);
nand UO_1568 (O_1568,N_27748,N_27342);
and UO_1569 (O_1569,N_25046,N_25600);
xor UO_1570 (O_1570,N_28756,N_29862);
nand UO_1571 (O_1571,N_29585,N_27671);
nand UO_1572 (O_1572,N_29048,N_29461);
nor UO_1573 (O_1573,N_25644,N_26039);
nor UO_1574 (O_1574,N_24672,N_29053);
nand UO_1575 (O_1575,N_29281,N_25544);
nand UO_1576 (O_1576,N_27574,N_28623);
nand UO_1577 (O_1577,N_28574,N_27782);
nand UO_1578 (O_1578,N_24437,N_26745);
nor UO_1579 (O_1579,N_28702,N_24595);
nand UO_1580 (O_1580,N_29609,N_24875);
nor UO_1581 (O_1581,N_29359,N_26459);
or UO_1582 (O_1582,N_24861,N_25985);
xor UO_1583 (O_1583,N_27607,N_27267);
xnor UO_1584 (O_1584,N_26490,N_25843);
and UO_1585 (O_1585,N_24510,N_26196);
and UO_1586 (O_1586,N_27208,N_27395);
or UO_1587 (O_1587,N_26214,N_28964);
nand UO_1588 (O_1588,N_25376,N_26082);
nand UO_1589 (O_1589,N_25056,N_25430);
and UO_1590 (O_1590,N_28024,N_25966);
xor UO_1591 (O_1591,N_24421,N_27614);
and UO_1592 (O_1592,N_25621,N_24936);
nand UO_1593 (O_1593,N_25998,N_29897);
xnor UO_1594 (O_1594,N_29137,N_26272);
or UO_1595 (O_1595,N_28491,N_26340);
xor UO_1596 (O_1596,N_24020,N_29357);
or UO_1597 (O_1597,N_27155,N_28344);
and UO_1598 (O_1598,N_25429,N_26376);
nor UO_1599 (O_1599,N_28778,N_26846);
nand UO_1600 (O_1600,N_29919,N_27562);
or UO_1601 (O_1601,N_26990,N_29499);
nor UO_1602 (O_1602,N_29055,N_28437);
or UO_1603 (O_1603,N_25681,N_29108);
nor UO_1604 (O_1604,N_25227,N_29790);
or UO_1605 (O_1605,N_25469,N_24756);
xnor UO_1606 (O_1606,N_28141,N_25707);
xor UO_1607 (O_1607,N_28776,N_29785);
or UO_1608 (O_1608,N_25537,N_29837);
nor UO_1609 (O_1609,N_24117,N_24385);
nor UO_1610 (O_1610,N_29246,N_26970);
nand UO_1611 (O_1611,N_29957,N_28112);
xor UO_1612 (O_1612,N_24988,N_28597);
xor UO_1613 (O_1613,N_25799,N_29620);
and UO_1614 (O_1614,N_28923,N_28243);
or UO_1615 (O_1615,N_29943,N_28578);
xor UO_1616 (O_1616,N_28947,N_24355);
nand UO_1617 (O_1617,N_29199,N_24167);
or UO_1618 (O_1618,N_24961,N_25612);
nor UO_1619 (O_1619,N_25122,N_24191);
nor UO_1620 (O_1620,N_28367,N_26803);
and UO_1621 (O_1621,N_27707,N_24611);
nand UO_1622 (O_1622,N_28186,N_28988);
or UO_1623 (O_1623,N_24170,N_26505);
nand UO_1624 (O_1624,N_28616,N_29960);
nand UO_1625 (O_1625,N_24955,N_27821);
nand UO_1626 (O_1626,N_24261,N_27095);
xnor UO_1627 (O_1627,N_29889,N_24169);
and UO_1628 (O_1628,N_24097,N_27909);
nor UO_1629 (O_1629,N_24908,N_27467);
nor UO_1630 (O_1630,N_26578,N_29657);
nor UO_1631 (O_1631,N_25720,N_24203);
or UO_1632 (O_1632,N_25566,N_28635);
nor UO_1633 (O_1633,N_28420,N_29171);
nor UO_1634 (O_1634,N_26107,N_24080);
or UO_1635 (O_1635,N_27798,N_29736);
nand UO_1636 (O_1636,N_28026,N_28991);
nand UO_1637 (O_1637,N_26195,N_27362);
nor UO_1638 (O_1638,N_25796,N_26255);
or UO_1639 (O_1639,N_28185,N_24310);
or UO_1640 (O_1640,N_27724,N_24686);
xor UO_1641 (O_1641,N_25930,N_24257);
xnor UO_1642 (O_1642,N_28428,N_24764);
and UO_1643 (O_1643,N_26565,N_29944);
nor UO_1644 (O_1644,N_24495,N_24602);
nand UO_1645 (O_1645,N_27157,N_27404);
nor UO_1646 (O_1646,N_25363,N_29747);
nor UO_1647 (O_1647,N_24506,N_29186);
or UO_1648 (O_1648,N_29067,N_28564);
nand UO_1649 (O_1649,N_26423,N_25375);
or UO_1650 (O_1650,N_28593,N_28076);
nand UO_1651 (O_1651,N_26222,N_26204);
or UO_1652 (O_1652,N_27148,N_28519);
nor UO_1653 (O_1653,N_24977,N_26493);
xnor UO_1654 (O_1654,N_29287,N_25691);
nor UO_1655 (O_1655,N_26041,N_27794);
or UO_1656 (O_1656,N_29533,N_26234);
or UO_1657 (O_1657,N_27359,N_28151);
and UO_1658 (O_1658,N_27739,N_24124);
nand UO_1659 (O_1659,N_28588,N_26812);
or UO_1660 (O_1660,N_29198,N_28917);
and UO_1661 (O_1661,N_25149,N_28117);
and UO_1662 (O_1662,N_26582,N_28523);
or UO_1663 (O_1663,N_28996,N_25093);
and UO_1664 (O_1664,N_26910,N_25494);
nand UO_1665 (O_1665,N_25700,N_27423);
nor UO_1666 (O_1666,N_28085,N_29169);
xnor UO_1667 (O_1667,N_24980,N_29012);
and UO_1668 (O_1668,N_28618,N_28791);
and UO_1669 (O_1669,N_25550,N_26198);
nand UO_1670 (O_1670,N_25307,N_24380);
xnor UO_1671 (O_1671,N_24476,N_25580);
or UO_1672 (O_1672,N_27420,N_27826);
and UO_1673 (O_1673,N_28481,N_25179);
nand UO_1674 (O_1674,N_29587,N_27932);
nor UO_1675 (O_1675,N_27948,N_27059);
or UO_1676 (O_1676,N_29982,N_27786);
xor UO_1677 (O_1677,N_29464,N_27805);
or UO_1678 (O_1678,N_26744,N_25823);
xor UO_1679 (O_1679,N_28279,N_25567);
and UO_1680 (O_1680,N_27773,N_25504);
nand UO_1681 (O_1681,N_29479,N_26475);
xor UO_1682 (O_1682,N_27117,N_24199);
xnor UO_1683 (O_1683,N_29339,N_24215);
and UO_1684 (O_1684,N_25806,N_25206);
and UO_1685 (O_1685,N_26456,N_28434);
and UO_1686 (O_1686,N_25701,N_29020);
and UO_1687 (O_1687,N_24029,N_25331);
xor UO_1688 (O_1688,N_25871,N_24652);
nand UO_1689 (O_1689,N_25210,N_24194);
nor UO_1690 (O_1690,N_27012,N_25816);
xnor UO_1691 (O_1691,N_29131,N_29686);
nor UO_1692 (O_1692,N_29298,N_28397);
or UO_1693 (O_1693,N_28673,N_24972);
nand UO_1694 (O_1694,N_26237,N_24535);
nand UO_1695 (O_1695,N_26127,N_25177);
nor UO_1696 (O_1696,N_26452,N_28636);
xor UO_1697 (O_1697,N_28166,N_27991);
xnor UO_1698 (O_1698,N_24984,N_29598);
or UO_1699 (O_1699,N_25265,N_28463);
nor UO_1700 (O_1700,N_29058,N_27407);
and UO_1701 (O_1701,N_28819,N_26862);
xnor UO_1702 (O_1702,N_29933,N_27427);
nor UO_1703 (O_1703,N_27349,N_24657);
nand UO_1704 (O_1704,N_24033,N_25908);
and UO_1705 (O_1705,N_25505,N_27611);
xnor UO_1706 (O_1706,N_24135,N_25466);
xnor UO_1707 (O_1707,N_29155,N_25576);
xor UO_1708 (O_1708,N_26712,N_27706);
and UO_1709 (O_1709,N_27868,N_28532);
and UO_1710 (O_1710,N_27894,N_29938);
nor UO_1711 (O_1711,N_26134,N_27940);
xor UO_1712 (O_1712,N_28647,N_24291);
nor UO_1713 (O_1713,N_25021,N_28913);
xor UO_1714 (O_1714,N_27041,N_28206);
xor UO_1715 (O_1715,N_25232,N_27787);
nand UO_1716 (O_1716,N_25680,N_28624);
nor UO_1717 (O_1717,N_28443,N_28352);
and UO_1718 (O_1718,N_27492,N_24830);
xnor UO_1719 (O_1719,N_25080,N_27915);
or UO_1720 (O_1720,N_29675,N_26072);
or UO_1721 (O_1721,N_24186,N_27928);
nand UO_1722 (O_1722,N_27584,N_26035);
xnor UO_1723 (O_1723,N_25790,N_28124);
nand UO_1724 (O_1724,N_29557,N_27365);
and UO_1725 (O_1725,N_27216,N_27174);
nand UO_1726 (O_1726,N_24963,N_25944);
nand UO_1727 (O_1727,N_25978,N_29254);
nand UO_1728 (O_1728,N_24456,N_25302);
nand UO_1729 (O_1729,N_24698,N_26572);
or UO_1730 (O_1730,N_24269,N_28648);
nor UO_1731 (O_1731,N_28239,N_25593);
or UO_1732 (O_1732,N_29295,N_24985);
xnor UO_1733 (O_1733,N_24426,N_27287);
xnor UO_1734 (O_1734,N_26353,N_28104);
and UO_1735 (O_1735,N_25614,N_24502);
or UO_1736 (O_1736,N_29205,N_29866);
nand UO_1737 (O_1737,N_26583,N_29399);
nand UO_1738 (O_1738,N_26576,N_24264);
or UO_1739 (O_1739,N_25591,N_27662);
nor UO_1740 (O_1740,N_28712,N_27172);
nand UO_1741 (O_1741,N_28598,N_29188);
nor UO_1742 (O_1742,N_29310,N_27592);
nor UO_1743 (O_1743,N_29563,N_26517);
xnor UO_1744 (O_1744,N_29580,N_26815);
xor UO_1745 (O_1745,N_29029,N_24031);
xnor UO_1746 (O_1746,N_26638,N_26932);
nand UO_1747 (O_1747,N_26182,N_27175);
and UO_1748 (O_1748,N_27864,N_27682);
and UO_1749 (O_1749,N_26445,N_25563);
nor UO_1750 (O_1750,N_24927,N_25040);
xnor UO_1751 (O_1751,N_28686,N_29754);
nor UO_1752 (O_1752,N_29107,N_26535);
and UO_1753 (O_1753,N_27631,N_29100);
nor UO_1754 (O_1754,N_24976,N_24665);
nor UO_1755 (O_1755,N_25981,N_26221);
or UO_1756 (O_1756,N_26027,N_28658);
nor UO_1757 (O_1757,N_29664,N_26183);
and UO_1758 (O_1758,N_29796,N_29771);
or UO_1759 (O_1759,N_29411,N_24727);
xnor UO_1760 (O_1760,N_29106,N_29400);
and UO_1761 (O_1761,N_29352,N_29082);
or UO_1762 (O_1762,N_29691,N_25268);
xor UO_1763 (O_1763,N_26814,N_26254);
and UO_1764 (O_1764,N_28110,N_27368);
and UO_1765 (O_1765,N_27945,N_24450);
nor UO_1766 (O_1766,N_29309,N_29988);
nand UO_1767 (O_1767,N_28693,N_25810);
xnor UO_1768 (O_1768,N_28211,N_28769);
nand UO_1769 (O_1769,N_27545,N_26606);
and UO_1770 (O_1770,N_27259,N_26118);
nand UO_1771 (O_1771,N_25226,N_26133);
xnor UO_1772 (O_1772,N_24151,N_24263);
xor UO_1773 (O_1773,N_28177,N_28934);
and UO_1774 (O_1774,N_25082,N_28640);
and UO_1775 (O_1775,N_25394,N_24251);
nand UO_1776 (O_1776,N_27742,N_29143);
nor UO_1777 (O_1777,N_26539,N_28324);
nand UO_1778 (O_1778,N_29726,N_29203);
or UO_1779 (O_1779,N_28017,N_27450);
nand UO_1780 (O_1780,N_25559,N_27543);
xnor UO_1781 (O_1781,N_26119,N_29519);
and UO_1782 (O_1782,N_25915,N_26318);
nor UO_1783 (O_1783,N_28863,N_29991);
and UO_1784 (O_1784,N_26044,N_28568);
nor UO_1785 (O_1785,N_24804,N_26411);
or UO_1786 (O_1786,N_24775,N_27575);
xnor UO_1787 (O_1787,N_27391,N_28171);
and UO_1788 (O_1788,N_27637,N_26851);
xor UO_1789 (O_1789,N_27955,N_29440);
nand UO_1790 (O_1790,N_28590,N_28743);
nand UO_1791 (O_1791,N_26612,N_29133);
or UO_1792 (O_1792,N_29406,N_24520);
nand UO_1793 (O_1793,N_27052,N_26879);
nor UO_1794 (O_1794,N_27972,N_26989);
nor UO_1795 (O_1795,N_25716,N_27167);
xnor UO_1796 (O_1796,N_28013,N_26984);
nor UO_1797 (O_1797,N_28943,N_27439);
or UO_1798 (O_1798,N_26513,N_28552);
nand UO_1799 (O_1799,N_24946,N_27882);
and UO_1800 (O_1800,N_24247,N_29581);
or UO_1801 (O_1801,N_25409,N_27186);
or UO_1802 (O_1802,N_25065,N_24741);
xor UO_1803 (O_1803,N_24854,N_29491);
or UO_1804 (O_1804,N_28319,N_27507);
or UO_1805 (O_1805,N_29083,N_26631);
or UO_1806 (O_1806,N_27177,N_27731);
nand UO_1807 (O_1807,N_25653,N_28698);
xnor UO_1808 (O_1808,N_28688,N_25322);
and UO_1809 (O_1809,N_29124,N_27534);
and UO_1810 (O_1810,N_24303,N_26765);
nor UO_1811 (O_1811,N_27913,N_28260);
nor UO_1812 (O_1812,N_26652,N_25171);
xor UO_1813 (O_1813,N_26218,N_25766);
or UO_1814 (O_1814,N_28882,N_28268);
nand UO_1815 (O_1815,N_25792,N_27279);
nand UO_1816 (O_1816,N_27515,N_27849);
nor UO_1817 (O_1817,N_26545,N_25416);
xnor UO_1818 (O_1818,N_25005,N_25395);
nand UO_1819 (O_1819,N_29097,N_29259);
nor UO_1820 (O_1820,N_27026,N_29139);
nor UO_1821 (O_1821,N_28713,N_29813);
nand UO_1822 (O_1822,N_27939,N_28179);
or UO_1823 (O_1823,N_29901,N_29396);
or UO_1824 (O_1824,N_25894,N_26230);
xnor UO_1825 (O_1825,N_27881,N_29261);
or UO_1826 (O_1826,N_24968,N_24962);
and UO_1827 (O_1827,N_27261,N_27263);
nand UO_1828 (O_1828,N_25251,N_28967);
nor UO_1829 (O_1829,N_26055,N_26212);
xnor UO_1830 (O_1830,N_24547,N_29799);
xor UO_1831 (O_1831,N_29674,N_24479);
nor UO_1832 (O_1832,N_29085,N_29543);
nor UO_1833 (O_1833,N_26388,N_27814);
xor UO_1834 (O_1834,N_29515,N_27410);
and UO_1835 (O_1835,N_28329,N_29145);
nand UO_1836 (O_1836,N_26355,N_29876);
xor UO_1837 (O_1837,N_24480,N_29792);
or UO_1838 (O_1838,N_28507,N_27459);
or UO_1839 (O_1839,N_26834,N_26049);
nand UO_1840 (O_1840,N_28542,N_28887);
and UO_1841 (O_1841,N_27630,N_26929);
xor UO_1842 (O_1842,N_29638,N_27589);
or UO_1843 (O_1843,N_26575,N_26060);
nand UO_1844 (O_1844,N_29588,N_29219);
xnor UO_1845 (O_1845,N_29963,N_25762);
nor UO_1846 (O_1846,N_28152,N_25753);
and UO_1847 (O_1847,N_26838,N_25874);
and UO_1848 (O_1848,N_27358,N_25464);
xnor UO_1849 (O_1849,N_25692,N_24182);
nand UO_1850 (O_1850,N_29216,N_28316);
nor UO_1851 (O_1851,N_25445,N_29811);
or UO_1852 (O_1852,N_25532,N_26551);
or UO_1853 (O_1853,N_25759,N_26566);
xnor UO_1854 (O_1854,N_27477,N_29451);
nor UO_1855 (O_1855,N_26863,N_25756);
xnor UO_1856 (O_1856,N_24042,N_27374);
xnor UO_1857 (O_1857,N_27088,N_29896);
or UO_1858 (O_1858,N_27674,N_27604);
nand UO_1859 (O_1859,N_29985,N_28450);
and UO_1860 (O_1860,N_29920,N_28500);
and UO_1861 (O_1861,N_28581,N_25770);
nor UO_1862 (O_1862,N_26031,N_24246);
and UO_1863 (O_1863,N_26808,N_26295);
xnor UO_1864 (O_1864,N_25288,N_29968);
or UO_1865 (O_1865,N_24605,N_26324);
or UO_1866 (O_1866,N_24441,N_29268);
or UO_1867 (O_1867,N_28891,N_24703);
nor UO_1868 (O_1868,N_26068,N_28361);
and UO_1869 (O_1869,N_28422,N_26675);
xnor UO_1870 (O_1870,N_26885,N_28974);
or UO_1871 (O_1871,N_28879,N_25842);
nand UO_1872 (O_1872,N_25751,N_29345);
nand UO_1873 (O_1873,N_25587,N_24675);
or UO_1874 (O_1874,N_27891,N_27677);
or UO_1875 (O_1875,N_29709,N_29201);
nand UO_1876 (O_1876,N_27055,N_29672);
and UO_1877 (O_1877,N_26580,N_24918);
nor UO_1878 (O_1878,N_25764,N_27886);
nand UO_1879 (O_1879,N_27799,N_24458);
nand UO_1880 (O_1880,N_28898,N_28752);
nand UO_1881 (O_1881,N_29723,N_29507);
nand UO_1882 (O_1882,N_27633,N_25620);
and UO_1883 (O_1883,N_27542,N_29070);
nor UO_1884 (O_1884,N_25220,N_25346);
and UO_1885 (O_1885,N_25181,N_29351);
or UO_1886 (O_1886,N_24279,N_28685);
or UO_1887 (O_1887,N_25528,N_27352);
nor UO_1888 (O_1888,N_24543,N_24216);
xor UO_1889 (O_1889,N_29380,N_28612);
xnor UO_1890 (O_1890,N_29273,N_28952);
or UO_1891 (O_1891,N_25077,N_24816);
nand UO_1892 (O_1892,N_26356,N_29319);
or UO_1893 (O_1893,N_27064,N_28421);
xor UO_1894 (O_1894,N_25689,N_25527);
nand UO_1895 (O_1895,N_28585,N_26116);
nand UO_1896 (O_1896,N_26955,N_29120);
nor UO_1897 (O_1897,N_26718,N_25079);
and UO_1898 (O_1898,N_29851,N_29767);
or UO_1899 (O_1899,N_26998,N_29350);
nand UO_1900 (O_1900,N_28557,N_26036);
xor UO_1901 (O_1901,N_26190,N_25396);
nor UO_1902 (O_1902,N_24994,N_25579);
nor UO_1903 (O_1903,N_24952,N_27973);
or UO_1904 (O_1904,N_26633,N_28774);
and UO_1905 (O_1905,N_28946,N_28716);
or UO_1906 (O_1906,N_24225,N_24313);
nand UO_1907 (O_1907,N_28313,N_24823);
or UO_1908 (O_1908,N_27779,N_28132);
and UO_1909 (O_1909,N_28827,N_26187);
nor UO_1910 (O_1910,N_26262,N_25502);
and UO_1911 (O_1911,N_25524,N_28455);
or UO_1912 (O_1912,N_27852,N_24713);
xor UO_1913 (O_1913,N_29476,N_27681);
nand UO_1914 (O_1914,N_24551,N_26991);
or UO_1915 (O_1915,N_25642,N_29922);
and UO_1916 (O_1916,N_25955,N_29701);
xor UO_1917 (O_1917,N_24139,N_26185);
nand UO_1918 (O_1918,N_24157,N_29402);
nor UO_1919 (O_1919,N_26086,N_24534);
nand UO_1920 (O_1920,N_29170,N_28954);
nand UO_1921 (O_1921,N_29725,N_28953);
nor UO_1922 (O_1922,N_24683,N_26317);
nand UO_1923 (O_1923,N_27565,N_29063);
xnor UO_1924 (O_1924,N_24957,N_27392);
or UO_1925 (O_1925,N_26723,N_25824);
and UO_1926 (O_1926,N_29770,N_27316);
and UO_1927 (O_1927,N_27946,N_27521);
nor UO_1928 (O_1928,N_27519,N_24274);
xor UO_1929 (O_1929,N_29030,N_26217);
xor UO_1930 (O_1930,N_28025,N_29660);
or UO_1931 (O_1931,N_28348,N_24483);
xor UO_1932 (O_1932,N_25461,N_29245);
and UO_1933 (O_1933,N_28582,N_26587);
nand UO_1934 (O_1934,N_25073,N_26156);
or UO_1935 (O_1935,N_29848,N_25594);
nand UO_1936 (O_1936,N_24459,N_29487);
xor UO_1937 (O_1937,N_28971,N_24981);
xnor UO_1938 (O_1938,N_26409,N_27246);
and UO_1939 (O_1939,N_26379,N_28706);
and UO_1940 (O_1940,N_27623,N_29326);
xor UO_1941 (O_1941,N_27841,N_27328);
and UO_1942 (O_1942,N_24275,N_27215);
and UO_1943 (O_1943,N_26435,N_24993);
xor UO_1944 (O_1944,N_26840,N_24433);
nor UO_1945 (O_1945,N_27120,N_24773);
nand UO_1946 (O_1946,N_27356,N_26363);
and UO_1947 (O_1947,N_24272,N_28095);
and UO_1948 (O_1948,N_28069,N_29806);
nor UO_1949 (O_1949,N_28665,N_25786);
or UO_1950 (O_1950,N_27688,N_24362);
xnor UO_1951 (O_1951,N_29153,N_27713);
and UO_1952 (O_1952,N_27895,N_28956);
nor UO_1953 (O_1953,N_26888,N_28883);
xnor UO_1954 (O_1954,N_24379,N_29579);
and UO_1955 (O_1955,N_24143,N_24335);
nor UO_1956 (O_1956,N_27654,N_26289);
nand UO_1957 (O_1957,N_29758,N_25050);
nand UO_1958 (O_1958,N_27922,N_28531);
nor UO_1959 (O_1959,N_29845,N_25219);
or UO_1960 (O_1960,N_26939,N_29223);
xor UO_1961 (O_1961,N_24960,N_24114);
or UO_1962 (O_1962,N_29119,N_27732);
xor UO_1963 (O_1963,N_27422,N_26868);
nor UO_1964 (O_1964,N_27634,N_28817);
or UO_1965 (O_1965,N_24397,N_26629);
xnor UO_1966 (O_1966,N_29277,N_24429);
and UO_1967 (O_1967,N_26220,N_28480);
nand UO_1968 (O_1968,N_28003,N_24314);
xnor UO_1969 (O_1969,N_24068,N_29425);
or UO_1970 (O_1970,N_25905,N_29441);
and UO_1971 (O_1971,N_25481,N_24835);
or UO_1972 (O_1972,N_29583,N_26896);
nor UO_1973 (O_1973,N_26923,N_29538);
and UO_1974 (O_1974,N_24638,N_24620);
and UO_1975 (O_1975,N_26866,N_29069);
or UO_1976 (O_1976,N_27880,N_24697);
or UO_1977 (O_1977,N_27406,N_28955);
or UO_1978 (O_1978,N_27377,N_26126);
nand UO_1979 (O_1979,N_25493,N_28067);
nand UO_1980 (O_1980,N_28634,N_27009);
and UO_1981 (O_1981,N_27875,N_28358);
or UO_1982 (O_1982,N_29559,N_24663);
nand UO_1983 (O_1983,N_29871,N_25324);
xnor UO_1984 (O_1984,N_28867,N_25957);
nor UO_1985 (O_1985,N_28409,N_26837);
nand UO_1986 (O_1986,N_27189,N_24666);
nor UO_1987 (O_1987,N_25355,N_25602);
and UO_1988 (O_1988,N_25629,N_29009);
nor UO_1989 (O_1989,N_25885,N_24798);
and UO_1990 (O_1990,N_28089,N_27454);
and UO_1991 (O_1991,N_28364,N_26733);
and UO_1992 (O_1992,N_24427,N_24419);
nor UO_1993 (O_1993,N_28392,N_29631);
nand UO_1994 (O_1994,N_27985,N_27819);
nand UO_1995 (O_1995,N_24554,N_26735);
nand UO_1996 (O_1996,N_28857,N_28046);
nor UO_1997 (O_1997,N_29000,N_25403);
nor UO_1998 (O_1998,N_27818,N_24526);
nand UO_1999 (O_1999,N_29234,N_25912);
nor UO_2000 (O_2000,N_26919,N_24052);
and UO_2001 (O_2001,N_28865,N_24859);
nand UO_2002 (O_2002,N_28901,N_29829);
xnor UO_2003 (O_2003,N_27714,N_25415);
nand UO_2004 (O_2004,N_24258,N_25746);
xor UO_2005 (O_2005,N_27438,N_26877);
xnor UO_2006 (O_2006,N_28499,N_29321);
or UO_2007 (O_2007,N_25083,N_26577);
or UO_2008 (O_2008,N_29466,N_27057);
nor UO_2009 (O_2009,N_29101,N_26537);
or UO_2010 (O_2010,N_27581,N_24159);
nand UO_2011 (O_2011,N_28679,N_24093);
and UO_2012 (O_2012,N_24524,N_29343);
nand UO_2013 (O_2013,N_28388,N_29026);
nand UO_2014 (O_2014,N_28536,N_26401);
or UO_2015 (O_2015,N_28873,N_25495);
nor UO_2016 (O_2016,N_28575,N_25482);
nor UO_2017 (O_2017,N_29196,N_29651);
nand UO_2018 (O_2018,N_24018,N_25715);
or UO_2019 (O_2019,N_25596,N_25902);
and UO_2020 (O_2020,N_25444,N_26915);
or UO_2021 (O_2021,N_29929,N_29472);
nor UO_2022 (O_2022,N_26052,N_29284);
and UO_2023 (O_2023,N_28453,N_29450);
nand UO_2024 (O_2024,N_28958,N_26592);
nor UO_2025 (O_2025,N_27066,N_27679);
or UO_2026 (O_2026,N_25152,N_29290);
nor UO_2027 (O_2027,N_24197,N_27602);
nand UO_2028 (O_2028,N_29150,N_24254);
nand UO_2029 (O_2029,N_25708,N_29332);
nor UO_2030 (O_2030,N_27887,N_24992);
nand UO_2031 (O_2031,N_28768,N_24455);
nor UO_2032 (O_2032,N_24975,N_24363);
and UO_2033 (O_2033,N_29605,N_29569);
nand UO_2034 (O_2034,N_29019,N_27965);
nor UO_2035 (O_2035,N_28705,N_27853);
and UO_2036 (O_2036,N_24575,N_28403);
or UO_2037 (O_2037,N_26096,N_28162);
nand UO_2038 (O_2038,N_29258,N_29942);
nand UO_2039 (O_2039,N_28540,N_24235);
nand UO_2040 (O_2040,N_27218,N_29493);
or UO_2041 (O_2041,N_28944,N_29618);
nor UO_2042 (O_2042,N_26335,N_27457);
xnor UO_2043 (O_2043,N_25257,N_26054);
nand UO_2044 (O_2044,N_27659,N_29465);
xnor UO_2045 (O_2045,N_26827,N_28290);
or UO_2046 (O_2046,N_26210,N_29662);
nand UO_2047 (O_2047,N_26861,N_26106);
and UO_2048 (O_2048,N_28144,N_28554);
xnor UO_2049 (O_2049,N_27931,N_25299);
xor UO_2050 (O_2050,N_28346,N_26597);
xnor UO_2051 (O_2051,N_24682,N_28535);
or UO_2052 (O_2052,N_24008,N_26203);
and UO_2053 (O_2053,N_28625,N_27320);
nand UO_2054 (O_2054,N_29545,N_28915);
nand UO_2055 (O_2055,N_28295,N_26763);
xnor UO_2056 (O_2056,N_24443,N_27235);
nand UO_2057 (O_2057,N_28390,N_25857);
or UO_2058 (O_2058,N_24334,N_26320);
nor UO_2059 (O_2059,N_26823,N_26398);
and UO_2060 (O_2060,N_27027,N_28680);
nor UO_2061 (O_2061,N_26649,N_28075);
or UO_2062 (O_2062,N_26347,N_27244);
or UO_2063 (O_2063,N_26950,N_29238);
nor UO_2064 (O_2064,N_27728,N_26377);
nor UO_2065 (O_2065,N_29312,N_29821);
nand UO_2066 (O_2066,N_25490,N_26746);
nand UO_2067 (O_2067,N_24827,N_24233);
and UO_2068 (O_2068,N_27361,N_28197);
and UO_2069 (O_2069,N_27417,N_26362);
and UO_2070 (O_2070,N_29093,N_29154);
nand UO_2071 (O_2071,N_26213,N_25656);
nand UO_2072 (O_2072,N_26796,N_28298);
nand UO_2073 (O_2073,N_26042,N_29080);
nand UO_2074 (O_2074,N_26527,N_28733);
nand UO_2075 (O_2075,N_28371,N_24566);
nand UO_2076 (O_2076,N_24230,N_28477);
xor UO_2077 (O_2077,N_24706,N_27470);
xor UO_2078 (O_2078,N_26313,N_28699);
nor UO_2079 (O_2079,N_27718,N_26216);
or UO_2080 (O_2080,N_28184,N_26848);
or UO_2081 (O_2081,N_24845,N_27540);
xnor UO_2082 (O_2082,N_25034,N_28485);
or UO_2083 (O_2083,N_29446,N_24596);
xnor UO_2084 (O_2084,N_29574,N_29971);
xnor UO_2085 (O_2085,N_29861,N_25256);
or UO_2086 (O_2086,N_29325,N_25061);
nand UO_2087 (O_2087,N_29903,N_27348);
xor UO_2088 (O_2088,N_24920,N_25196);
and UO_2089 (O_2089,N_27974,N_28223);
or UO_2090 (O_2090,N_25606,N_25710);
xor UO_2091 (O_2091,N_27301,N_29608);
nor UO_2092 (O_2092,N_24616,N_24148);
and UO_2093 (O_2093,N_29622,N_27428);
or UO_2094 (O_2094,N_26824,N_26158);
nor UO_2095 (O_2095,N_29535,N_27113);
nand UO_2096 (O_2096,N_25489,N_26238);
xnor UO_2097 (O_2097,N_26148,N_28555);
nor UO_2098 (O_2098,N_29361,N_28600);
nor UO_2099 (O_2099,N_28694,N_24921);
nand UO_2100 (O_2100,N_24494,N_29632);
xnor UO_2101 (O_2101,N_26992,N_28082);
or UO_2102 (O_2102,N_24116,N_25189);
and UO_2103 (O_2103,N_29328,N_28488);
and UO_2104 (O_2104,N_29354,N_24208);
nor UO_2105 (O_2105,N_26967,N_29337);
xnor UO_2106 (O_2106,N_27591,N_28807);
nor UO_2107 (O_2107,N_27433,N_25165);
nand UO_2108 (O_2108,N_27857,N_28235);
xnor UO_2109 (O_2109,N_24842,N_24207);
or UO_2110 (O_2110,N_28192,N_29578);
xnor UO_2111 (O_2111,N_24195,N_28889);
xor UO_2112 (O_2112,N_27954,N_28287);
or UO_2113 (O_2113,N_27582,N_24593);
nand UO_2114 (O_2114,N_25652,N_26191);
nand UO_2115 (O_2115,N_26658,N_26147);
or UO_2116 (O_2116,N_27270,N_25847);
nor UO_2117 (O_2117,N_25402,N_28942);
or UO_2118 (O_2118,N_29623,N_27725);
nor UO_2119 (O_2119,N_28475,N_24333);
nand UO_2120 (O_2120,N_24290,N_24654);
xor UO_2121 (O_2121,N_24411,N_28677);
nor UO_2122 (O_2122,N_26373,N_26312);
or UO_2123 (O_2123,N_25932,N_27268);
and UO_2124 (O_2124,N_26428,N_26995);
xnor UO_2125 (O_2125,N_28220,N_24851);
and UO_2126 (O_2126,N_28644,N_24847);
nand UO_2127 (O_2127,N_27149,N_29228);
or UO_2128 (O_2128,N_25778,N_25875);
and UO_2129 (O_2129,N_29648,N_28267);
nand UO_2130 (O_2130,N_26461,N_24786);
or UO_2131 (O_2131,N_27171,N_27010);
or UO_2132 (O_2132,N_24046,N_27309);
or UO_2133 (O_2133,N_25458,N_27898);
and UO_2134 (O_2134,N_25598,N_26381);
nor UO_2135 (O_2135,N_28449,N_26507);
xor UO_2136 (O_2136,N_25533,N_28823);
nor UO_2137 (O_2137,N_29781,N_24027);
or UO_2138 (O_2138,N_25140,N_25244);
or UO_2139 (O_2139,N_28831,N_29065);
or UO_2140 (O_2140,N_27360,N_27222);
nor UO_2141 (O_2141,N_29338,N_25989);
and UO_2142 (O_2142,N_24026,N_28158);
and UO_2143 (O_2143,N_26725,N_26080);
or UO_2144 (O_2144,N_29432,N_24515);
or UO_2145 (O_2145,N_27179,N_28935);
nand UO_2146 (O_2146,N_24354,N_26786);
or UO_2147 (O_2147,N_29542,N_25353);
or UO_2148 (O_2148,N_24615,N_27647);
nor UO_2149 (O_2149,N_24630,N_29779);
or UO_2150 (O_2150,N_28890,N_28818);
nand UO_2151 (O_2151,N_27690,N_29311);
or UO_2152 (O_2152,N_26131,N_24746);
nand UO_2153 (O_2153,N_27744,N_26567);
or UO_2154 (O_2154,N_25330,N_27184);
xor UO_2155 (O_2155,N_26351,N_27599);
or UO_2156 (O_2156,N_28021,N_27808);
and UO_2157 (O_2157,N_28798,N_26352);
nand UO_2158 (O_2158,N_24632,N_29969);
nand UO_2159 (O_2159,N_24015,N_28730);
nor UO_2160 (O_2160,N_29653,N_25906);
nor UO_2161 (O_2161,N_26418,N_27025);
and UO_2162 (O_2162,N_24573,N_27062);
nand UO_2163 (O_2163,N_26976,N_28800);
nand UO_2164 (O_2164,N_24447,N_26128);
xor UO_2165 (O_2165,N_29500,N_25321);
or UO_2166 (O_2166,N_26064,N_26439);
xnor UO_2167 (O_2167,N_27004,N_28068);
and UO_2168 (O_2168,N_25958,N_29843);
nor UO_2169 (O_2169,N_25117,N_25314);
and UO_2170 (O_2170,N_28893,N_27100);
or UO_2171 (O_2171,N_29526,N_26850);
or UO_2172 (O_2172,N_28837,N_26666);
nor UO_2173 (O_2173,N_26123,N_24548);
and UO_2174 (O_2174,N_28796,N_24115);
nor UO_2175 (O_2175,N_25133,N_29541);
or UO_2176 (O_2176,N_27860,N_26764);
or UO_2177 (O_2177,N_26757,N_29429);
nor UO_2178 (O_2178,N_28766,N_29853);
nand UO_2179 (O_2179,N_29468,N_27440);
or UO_2180 (O_2180,N_26903,N_28274);
and UO_2181 (O_2181,N_26114,N_28334);
and UO_2182 (O_2182,N_27444,N_27080);
nand UO_2183 (O_2183,N_25260,N_25252);
xnor UO_2184 (O_2184,N_28051,N_27236);
and UO_2185 (O_2185,N_27557,N_28262);
xor UO_2186 (O_2186,N_28762,N_28062);
or UO_2187 (O_2187,N_26095,N_28405);
and UO_2188 (O_2188,N_26532,N_26895);
nand UO_2189 (O_2189,N_28006,N_28465);
nor UO_2190 (O_2190,N_24924,N_25969);
or UO_2191 (O_2191,N_28895,N_26242);
nor UO_2192 (O_2192,N_28379,N_29986);
nand UO_2193 (O_2193,N_27746,N_29596);
and UO_2194 (O_2194,N_25424,N_28777);
nand UO_2195 (O_2195,N_29742,N_27997);
xor UO_2196 (O_2196,N_26548,N_26531);
nor UO_2197 (O_2197,N_24075,N_26913);
nor UO_2198 (O_2198,N_29809,N_28172);
and UO_2199 (O_2199,N_27230,N_25853);
nor UO_2200 (O_2200,N_26772,N_24370);
or UO_2201 (O_2201,N_28797,N_29383);
and UO_2202 (O_2202,N_24926,N_29696);
or UO_2203 (O_2203,N_27437,N_24722);
xor UO_2204 (O_2204,N_28044,N_29619);
or UO_2205 (O_2205,N_26280,N_24405);
nand UO_2206 (O_2206,N_25139,N_26807);
nand UO_2207 (O_2207,N_24131,N_24791);
xnor UO_2208 (O_2208,N_26977,N_29015);
xnor UO_2209 (O_2209,N_27335,N_29018);
or UO_2210 (O_2210,N_27803,N_28682);
nand UO_2211 (O_2211,N_28288,N_27628);
nand UO_2212 (O_2212,N_27264,N_25303);
nor UO_2213 (O_2213,N_25850,N_26506);
xor UO_2214 (O_2214,N_25327,N_28650);
and UO_2215 (O_2215,N_24716,N_29098);
nand UO_2216 (O_2216,N_28517,N_25676);
nor UO_2217 (O_2217,N_27924,N_27283);
xnor UO_2218 (O_2218,N_29612,N_28238);
nand UO_2219 (O_2219,N_28533,N_24866);
and UO_2220 (O_2220,N_25401,N_27138);
nand UO_2221 (O_2221,N_26711,N_24236);
or UO_2222 (O_2222,N_26470,N_26902);
or UO_2223 (O_2223,N_26809,N_27768);
or UO_2224 (O_2224,N_29900,N_24377);
xnor UO_2225 (O_2225,N_29276,N_25655);
nor UO_2226 (O_2226,N_27984,N_27548);
nand UO_2227 (O_2227,N_26433,N_28339);
xnor UO_2228 (O_2228,N_26206,N_24060);
xor UO_2229 (O_2229,N_25865,N_24136);
xor UO_2230 (O_2230,N_24829,N_24073);
xnor UO_2231 (O_2231,N_24887,N_27949);
nor UO_2232 (O_2232,N_29734,N_25356);
xnor UO_2233 (O_2233,N_26773,N_26949);
and UO_2234 (O_2234,N_26374,N_24431);
and UO_2235 (O_2235,N_29603,N_28722);
and UO_2236 (O_2236,N_25365,N_25698);
nor UO_2237 (O_2237,N_28710,N_25379);
or UO_2238 (O_2238,N_29523,N_24677);
xor UO_2239 (O_2239,N_28343,N_29681);
or UO_2240 (O_2240,N_25604,N_27926);
and UO_2241 (O_2241,N_27723,N_28143);
or UO_2242 (O_2242,N_26508,N_27938);
nand UO_2243 (O_2243,N_26632,N_29427);
nor UO_2244 (O_2244,N_24229,N_26070);
nand UO_2245 (O_2245,N_27777,N_29136);
xnor UO_2246 (O_2246,N_28054,N_27783);
nand UO_2247 (O_2247,N_24094,N_28795);
nand UO_2248 (O_2248,N_25625,N_25903);
nand UO_2249 (O_2249,N_27353,N_24780);
xnor UO_2250 (O_2250,N_28567,N_24346);
nand UO_2251 (O_2251,N_24610,N_28303);
nor UO_2252 (O_2252,N_25369,N_25963);
nand UO_2253 (O_2253,N_27056,N_29710);
nor UO_2254 (O_2254,N_27959,N_28900);
nor UO_2255 (O_2255,N_25693,N_28121);
xor UO_2256 (O_2256,N_25868,N_26595);
or UO_2257 (O_2257,N_29989,N_26669);
or UO_2258 (O_2258,N_25182,N_28529);
nor UO_2259 (O_2259,N_24467,N_29591);
or UO_2260 (O_2260,N_25086,N_27727);
or UO_2261 (O_2261,N_28254,N_24702);
or UO_2262 (O_2262,N_25779,N_28726);
xnor UO_2263 (O_2263,N_29644,N_24928);
nand UO_2264 (O_2264,N_28154,N_26975);
xnor UO_2265 (O_2265,N_24301,N_26301);
and UO_2266 (O_2266,N_27434,N_24792);
or UO_2267 (O_2267,N_24404,N_26078);
or UO_2268 (O_2268,N_26369,N_27237);
nand UO_2269 (O_2269,N_26232,N_26591);
or UO_2270 (O_2270,N_26139,N_26536);
nor UO_2271 (O_2271,N_28056,N_28246);
nor UO_2272 (O_2272,N_29102,N_28461);
nor UO_2273 (O_2273,N_28704,N_26460);
and UO_2274 (O_2274,N_27481,N_27040);
or UO_2275 (O_2275,N_26768,N_26978);
nand UO_2276 (O_2276,N_25377,N_24902);
and UO_2277 (O_2277,N_28354,N_27416);
xnor UO_2278 (O_2278,N_27888,N_27228);
and UO_2279 (O_2279,N_24240,N_26671);
or UO_2280 (O_2280,N_26348,N_24954);
nor UO_2281 (O_2281,N_25881,N_27551);
and UO_2282 (O_2282,N_26413,N_24733);
nand UO_2283 (O_2283,N_26951,N_29909);
nor UO_2284 (O_2284,N_25994,N_24428);
xnor UO_2285 (O_2285,N_26491,N_26432);
or UO_2286 (O_2286,N_24205,N_25116);
xor UO_2287 (O_2287,N_27105,N_29123);
or UO_2288 (O_2288,N_25510,N_27733);
nor UO_2289 (O_2289,N_28906,N_24878);
or UO_2290 (O_2290,N_25104,N_27509);
nor UO_2291 (O_2291,N_27831,N_27560);
nand UO_2292 (O_2292,N_24579,N_29818);
or UO_2293 (O_2293,N_25240,N_29159);
and UO_2294 (O_2294,N_24793,N_29654);
or UO_2295 (O_2295,N_26618,N_28081);
nor UO_2296 (O_2296,N_25057,N_29249);
nor UO_2297 (O_2297,N_28306,N_24237);
nor UO_2298 (O_2298,N_28019,N_25959);
xor UO_2299 (O_2299,N_24108,N_27608);
nor UO_2300 (O_2300,N_25126,N_25114);
and UO_2301 (O_2301,N_26415,N_24916);
or UO_2302 (O_2302,N_29006,N_29206);
xor UO_2303 (O_2303,N_29954,N_26249);
and UO_2304 (O_2304,N_24934,N_25907);
or UO_2305 (O_2305,N_25852,N_24761);
or UO_2306 (O_2306,N_26111,N_27622);
nand UO_2307 (O_2307,N_26641,N_26325);
nand UO_2308 (O_2308,N_27451,N_28972);
or UO_2309 (O_2309,N_25223,N_24645);
nand UO_2310 (O_2310,N_24452,N_25209);
xor UO_2311 (O_2311,N_28663,N_24412);
and UO_2312 (O_2312,N_26742,N_25965);
or UO_2313 (O_2313,N_26149,N_26627);
and UO_2314 (O_2314,N_25460,N_26088);
and UO_2315 (O_2315,N_24948,N_25108);
and UO_2316 (O_2316,N_27851,N_29358);
and UO_2317 (O_2317,N_29544,N_27048);
nand UO_2318 (O_2318,N_26968,N_25872);
nor UO_2319 (O_2319,N_24012,N_24544);
and UO_2320 (O_2320,N_24488,N_28058);
xor UO_2321 (O_2321,N_26117,N_29413);
or UO_2322 (O_2322,N_25060,N_29753);
and UO_2323 (O_2323,N_24013,N_27405);
xor UO_2324 (O_2324,N_24062,N_24065);
xnor UO_2325 (O_2325,N_29140,N_27288);
or UO_2326 (O_2326,N_25887,N_29247);
and UO_2327 (O_2327,N_25977,N_29057);
nand UO_2328 (O_2328,N_28881,N_27219);
or UO_2329 (O_2329,N_28040,N_27501);
xor UO_2330 (O_2330,N_25342,N_27685);
and UO_2331 (O_2331,N_25809,N_24388);
xor UO_2332 (O_2332,N_28451,N_27514);
or UO_2333 (O_2333,N_25940,N_26032);
nand UO_2334 (O_2334,N_24572,N_26141);
nor UO_2335 (O_2335,N_27497,N_26180);
or UO_2336 (O_2336,N_25155,N_26364);
xnor UO_2337 (O_2337,N_26228,N_28981);
or UO_2338 (O_2338,N_28411,N_26752);
or UO_2339 (O_2339,N_24132,N_24651);
nand UO_2340 (O_2340,N_26371,N_24760);
nand UO_2341 (O_2341,N_25831,N_26015);
nand UO_2342 (O_2342,N_27709,N_29126);
or UO_2343 (O_2343,N_27933,N_25884);
xor UO_2344 (O_2344,N_25072,N_28478);
and UO_2345 (O_2345,N_26125,N_28270);
and UO_2346 (O_2346,N_28902,N_28366);
or UO_2347 (O_2347,N_25237,N_27493);
nand UO_2348 (O_2348,N_28866,N_25878);
and UO_2349 (O_2349,N_28312,N_26043);
nand UO_2350 (O_2350,N_25951,N_27687);
nor UO_2351 (O_2351,N_28689,N_25262);
xnor UO_2352 (O_2352,N_24383,N_29698);
nand UO_2353 (O_2353,N_24107,N_27640);
and UO_2354 (O_2354,N_24732,N_25090);
nor UO_2355 (O_2355,N_27159,N_24462);
nor UO_2356 (O_2356,N_27274,N_28053);
and UO_2357 (O_2357,N_24521,N_28638);
nor UO_2358 (O_2358,N_24808,N_29071);
and UO_2359 (O_2359,N_26209,N_26655);
or UO_2360 (O_2360,N_27127,N_26936);
and UO_2361 (O_2361,N_27760,N_28910);
nand UO_2362 (O_2362,N_24089,N_28217);
nor UO_2363 (O_2363,N_27188,N_25595);
and UO_2364 (O_2364,N_29417,N_29727);
or UO_2365 (O_2365,N_25590,N_25931);
nor UO_2366 (O_2366,N_29602,N_24525);
or UO_2367 (O_2367,N_28997,N_26782);
or UO_2368 (O_2368,N_25880,N_26175);
and UO_2369 (O_2369,N_24529,N_24884);
or UO_2370 (O_2370,N_25106,N_25359);
nand UO_2371 (O_2371,N_27776,N_25581);
nor UO_2372 (O_2372,N_28849,N_25570);
or UO_2373 (O_2373,N_29315,N_25454);
xor UO_2374 (O_2374,N_29230,N_25222);
and UO_2375 (O_2375,N_24223,N_27618);
nor UO_2376 (O_2376,N_29997,N_27827);
xnor UO_2377 (O_2377,N_29056,N_25290);
or UO_2378 (O_2378,N_28538,N_27878);
xnor UO_2379 (O_2379,N_25988,N_28050);
or UO_2380 (O_2380,N_25383,N_26501);
xnor UO_2381 (O_2381,N_26270,N_29248);
or UO_2382 (O_2382,N_29947,N_24367);
nor UO_2383 (O_2383,N_24614,N_24297);
or UO_2384 (O_2384,N_29658,N_29445);
nand UO_2385 (O_2385,N_27793,N_28161);
and UO_2386 (O_2386,N_24539,N_26300);
or UO_2387 (O_2387,N_25463,N_25767);
nor UO_2388 (O_2388,N_29438,N_27252);
or UO_2389 (O_2389,N_25320,N_25275);
nand UO_2390 (O_2390,N_25128,N_25295);
or UO_2391 (O_2391,N_27306,N_27698);
xor UO_2392 (O_2392,N_26449,N_25561);
nor UO_2393 (O_2393,N_28277,N_27442);
or UO_2394 (O_2394,N_25858,N_24266);
xnor UO_2395 (O_2395,N_27813,N_25666);
and UO_2396 (O_2396,N_24930,N_27098);
nand UO_2397 (O_2397,N_24249,N_24696);
nand UO_2398 (O_2398,N_29121,N_27958);
nor UO_2399 (O_2399,N_27525,N_28813);
nand UO_2400 (O_2400,N_28690,N_28213);
nor UO_2401 (O_2401,N_28674,N_24590);
and UO_2402 (O_2402,N_28701,N_29517);
nand UO_2403 (O_2403,N_24797,N_27168);
xor UO_2404 (O_2404,N_25297,N_25825);
nor UO_2405 (O_2405,N_26172,N_29916);
xor UO_2406 (O_2406,N_29221,N_28514);
xnor UO_2407 (O_2407,N_25909,N_25388);
or UO_2408 (O_2408,N_26024,N_29855);
xnor UO_2409 (O_2409,N_29381,N_27128);
nand UO_2410 (O_2410,N_24245,N_27833);
or UO_2411 (O_2411,N_29034,N_27412);
nand UO_2412 (O_2412,N_29182,N_29379);
or UO_2413 (O_2413,N_28537,N_24848);
or UO_2414 (O_2414,N_26954,N_28750);
nor UO_2415 (O_2415,N_28394,N_29473);
nor UO_2416 (O_2416,N_24470,N_29780);
nor UO_2417 (O_2417,N_26514,N_26058);
nand UO_2418 (O_2418,N_28659,N_27151);
xor UO_2419 (O_2419,N_24711,N_24841);
xnor UO_2420 (O_2420,N_29611,N_28770);
or UO_2421 (O_2421,N_29774,N_25740);
or UO_2422 (O_2422,N_24024,N_25765);
or UO_2423 (O_2423,N_26549,N_26367);
and UO_2424 (O_2424,N_25094,N_29548);
nand UO_2425 (O_2425,N_28114,N_24528);
nand UO_2426 (O_2426,N_27873,N_26876);
and UO_2427 (O_2427,N_25525,N_26654);
xnor UO_2428 (O_2428,N_27124,N_28765);
xnor UO_2429 (O_2429,N_29301,N_27281);
or UO_2430 (O_2430,N_26504,N_27045);
nand UO_2431 (O_2431,N_29416,N_24417);
nor UO_2432 (O_2432,N_25608,N_27419);
xnor UO_2433 (O_2433,N_29814,N_24365);
nand UO_2434 (O_2434,N_27125,N_25942);
xnor UO_2435 (O_2435,N_28820,N_25075);
nor UO_2436 (O_2436,N_26688,N_29285);
xor UO_2437 (O_2437,N_27911,N_24647);
xnor UO_2438 (O_2438,N_27191,N_25343);
nand UO_2439 (O_2439,N_24569,N_26598);
nand UO_2440 (O_2440,N_29386,N_27533);
xnor UO_2441 (O_2441,N_27541,N_28180);
or UO_2442 (O_2442,N_24030,N_24940);
nand UO_2443 (O_2443,N_25357,N_27649);
nor UO_2444 (O_2444,N_25548,N_29458);
nand UO_2445 (O_2445,N_28205,N_28987);
xnor UO_2446 (O_2446,N_28973,N_26630);
and UO_2447 (O_2447,N_24378,N_28074);
xnor UO_2448 (O_2448,N_29297,N_29841);
nor UO_2449 (O_2449,N_25964,N_28066);
nand UO_2450 (O_2450,N_27307,N_24656);
xor UO_2451 (O_2451,N_29062,N_28926);
and UO_2452 (O_2452,N_29740,N_28047);
nand UO_2453 (O_2453,N_25367,N_29688);
nor UO_2454 (O_2454,N_25372,N_26361);
xnor UO_2455 (O_2455,N_26170,N_24726);
or UO_2456 (O_2456,N_24352,N_24300);
or UO_2457 (O_2457,N_24874,N_28760);
nor UO_2458 (O_2458,N_29313,N_25597);
or UO_2459 (O_2459,N_25286,N_26731);
or UO_2460 (O_2460,N_29682,N_26560);
or UO_2461 (O_2461,N_26161,N_25492);
nor UO_2462 (O_2462,N_25308,N_27885);
nand UO_2463 (O_2463,N_26478,N_25573);
nand UO_2464 (O_2464,N_29054,N_28558);
nor UO_2465 (O_2465,N_24051,N_26818);
xnor UO_2466 (O_2466,N_27139,N_24971);
or UO_2467 (O_2467,N_27319,N_24998);
nor UO_2468 (O_2468,N_28878,N_26020);
nand UO_2469 (O_2469,N_24735,N_27022);
xor UO_2470 (O_2470,N_26780,N_29974);
and UO_2471 (O_2471,N_25624,N_28851);
and UO_2472 (O_2472,N_29490,N_24913);
nor UO_2473 (O_2473,N_24850,N_29937);
or UO_2474 (O_2474,N_25276,N_26302);
and UO_2475 (O_2475,N_25103,N_29235);
nor UO_2476 (O_2476,N_25704,N_25771);
nor UO_2477 (O_2477,N_24982,N_25509);
nand UO_2478 (O_2478,N_24781,N_27903);
and UO_2479 (O_2479,N_25004,N_29408);
nand UO_2480 (O_2480,N_27854,N_27332);
nor UO_2481 (O_2481,N_28142,N_27842);
or UO_2482 (O_2482,N_27613,N_24609);
and UO_2483 (O_2483,N_25890,N_26559);
or UO_2484 (O_2484,N_27154,N_28323);
nor UO_2485 (O_2485,N_25800,N_24329);
xor UO_2486 (O_2486,N_29347,N_26920);
nand UO_2487 (O_2487,N_25168,N_29530);
or UO_2488 (O_2488,N_27755,N_29977);
nor UO_2489 (O_2489,N_27919,N_25479);
nand UO_2490 (O_2490,N_26315,N_25651);
or UO_2491 (O_2491,N_27280,N_28351);
nor UO_2492 (O_2492,N_28492,N_26258);
nor UO_2493 (O_2493,N_26667,N_27642);
and UO_2494 (O_2494,N_25081,N_27844);
nand UO_2495 (O_2495,N_26585,N_27767);
nand UO_2496 (O_2496,N_28734,N_26624);
nor UO_2497 (O_2497,N_26942,N_24966);
nor UO_2498 (O_2498,N_28497,N_25012);
nand UO_2499 (O_2499,N_27807,N_28511);
nor UO_2500 (O_2500,N_28892,N_25497);
and UO_2501 (O_2501,N_27559,N_29421);
nor UO_2502 (O_2502,N_27792,N_28253);
nor UO_2503 (O_2503,N_25803,N_28442);
or UO_2504 (O_2504,N_26985,N_28105);
xnor UO_2505 (O_2505,N_29728,N_26687);
and UO_2506 (O_2506,N_26722,N_26737);
and UO_2507 (O_2507,N_29506,N_25646);
and UO_2508 (O_2508,N_24674,N_28583);
and UO_2509 (O_2509,N_28527,N_25638);
or UO_2510 (O_2510,N_24776,N_25043);
or UO_2511 (O_2511,N_26864,N_24130);
xnor UO_2512 (O_2512,N_26322,N_24594);
nor UO_2513 (O_2513,N_28304,N_28092);
and UO_2514 (O_2514,N_25536,N_27797);
nand UO_2515 (O_2515,N_29776,N_24843);
nor UO_2516 (O_2516,N_26274,N_24324);
and UO_2517 (O_2517,N_24751,N_24678);
xnor UO_2518 (O_2518,N_27641,N_28995);
and UO_2519 (O_2519,N_26030,N_25521);
nor UO_2520 (O_2520,N_25616,N_26503);
and UO_2521 (O_2521,N_28368,N_27133);
xor UO_2522 (O_2522,N_25381,N_29966);
and UO_2523 (O_2523,N_27238,N_28330);
or UO_2524 (O_2524,N_25752,N_26079);
nor UO_2525 (O_2525,N_25859,N_26296);
nor UO_2526 (O_2526,N_27741,N_28992);
xnor UO_2527 (O_2527,N_25164,N_26804);
and UO_2528 (O_2528,N_27606,N_28410);
xnor UO_2529 (O_2529,N_28135,N_24839);
nand UO_2530 (O_2530,N_25728,N_29987);
nand UO_2531 (O_2531,N_29522,N_24049);
or UO_2532 (O_2532,N_24983,N_29562);
or UO_2533 (O_2533,N_25782,N_24077);
xnor UO_2534 (O_2534,N_27241,N_29278);
xor UO_2535 (O_2535,N_25575,N_24943);
xnor UO_2536 (O_2536,N_29768,N_29320);
nand UO_2537 (O_2537,N_26008,N_24111);
xnor UO_2538 (O_2538,N_24338,N_25225);
and UO_2539 (O_2539,N_25087,N_29637);
xor UO_2540 (O_2540,N_26344,N_29483);
nor UO_2541 (O_2541,N_24747,N_29299);
nand UO_2542 (O_2542,N_27114,N_25971);
and UO_2543 (O_2543,N_28649,N_26378);
and UO_2544 (O_2544,N_26023,N_25645);
or UO_2545 (O_2545,N_24693,N_24100);
nand UO_2546 (O_2546,N_28471,N_27295);
nor UO_2547 (O_2547,N_24813,N_27322);
or UO_2548 (O_2548,N_24045,N_25947);
xnor UO_2549 (O_2549,N_25428,N_29869);
nand UO_2550 (O_2550,N_29634,N_27964);
and UO_2551 (O_2551,N_28840,N_27180);
nand UO_2552 (O_2552,N_24893,N_27169);
or UO_2553 (O_2553,N_25835,N_27750);
and UO_2554 (O_2554,N_26832,N_29593);
and UO_2555 (O_2555,N_27865,N_25478);
and UO_2556 (O_2556,N_28784,N_25660);
or UO_2557 (O_2557,N_27766,N_26869);
xnor UO_2558 (O_2558,N_27134,N_28284);
or UO_2559 (O_2559,N_27981,N_28580);
xor UO_2560 (O_2560,N_25888,N_26485);
xor UO_2561 (O_2561,N_24110,N_24224);
or UO_2562 (O_2562,N_24867,N_28203);
nor UO_2563 (O_2563,N_26930,N_27282);
or UO_2564 (O_2564,N_26872,N_24778);
and UO_2565 (O_2565,N_25923,N_29816);
and UO_2566 (O_2566,N_26421,N_27753);
and UO_2567 (O_2567,N_29160,N_25064);
or UO_2568 (O_2568,N_24489,N_27778);
or UO_2569 (O_2569,N_26806,N_26943);
nand UO_2570 (O_2570,N_27552,N_26447);
xor UO_2571 (O_2571,N_29677,N_28963);
xor UO_2572 (O_2572,N_27195,N_24688);
nand UO_2573 (O_2573,N_27363,N_26635);
xor UO_2574 (O_2574,N_25292,N_29570);
nand UO_2575 (O_2575,N_27802,N_28541);
or UO_2576 (O_2576,N_24914,N_29670);
nor UO_2577 (O_2577,N_24743,N_27351);
nand UO_2578 (O_2578,N_29512,N_24796);
and UO_2579 (O_2579,N_24342,N_26215);
nand UO_2580 (O_2580,N_28065,N_29364);
or UO_2581 (O_2581,N_27245,N_28960);
xor UO_2582 (O_2582,N_25439,N_29976);
and UO_2583 (O_2583,N_27600,N_24629);
nand UO_2584 (O_2584,N_29755,N_29912);
and UO_2585 (O_2585,N_29886,N_27305);
xnor UO_2586 (O_2586,N_27272,N_28727);
or UO_2587 (O_2587,N_28509,N_29838);
or UO_2588 (O_2588,N_25661,N_29730);
xnor UO_2589 (O_2589,N_27809,N_29887);
nand UO_2590 (O_2590,N_28641,N_24200);
xor UO_2591 (O_2591,N_29636,N_24325);
xnor UO_2592 (O_2592,N_26339,N_28790);
nand UO_2593 (O_2593,N_27375,N_26948);
or UO_2594 (O_2594,N_24653,N_29748);
or UO_2595 (O_2595,N_27137,N_29208);
xnor UO_2596 (O_2596,N_26132,N_28107);
or UO_2597 (O_2597,N_26584,N_29766);
nor UO_2598 (O_2598,N_26419,N_29606);
nor UO_2599 (O_2599,N_24894,N_25123);
xnor UO_2600 (O_2600,N_27646,N_27231);
nand UO_2601 (O_2601,N_28101,N_29763);
and UO_2602 (O_2602,N_29046,N_28078);
nor UO_2603 (O_2603,N_29905,N_26164);
nand UO_2604 (O_2604,N_29128,N_25233);
nand UO_2605 (O_2605,N_28539,N_26269);
and UO_2606 (O_2606,N_29368,N_26474);
or UO_2607 (O_2607,N_28739,N_28208);
nor UO_2608 (O_2608,N_24401,N_26243);
nand UO_2609 (O_2609,N_29697,N_27119);
or UO_2610 (O_2610,N_28183,N_26963);
nand UO_2611 (O_2611,N_24478,N_24498);
xnor UO_2612 (O_2612,N_24889,N_24368);
or UO_2613 (O_2613,N_27675,N_29761);
xnor UO_2614 (O_2614,N_28391,N_29906);
nor UO_2615 (O_2615,N_25323,N_29384);
xor UO_2616 (O_2616,N_29142,N_29183);
nand UO_2617 (O_2617,N_28011,N_26908);
nand UO_2618 (O_2618,N_25851,N_28194);
xnor UO_2619 (O_2619,N_28393,N_28269);
or UO_2620 (O_2620,N_25586,N_24694);
xnor UO_2621 (O_2621,N_25750,N_24637);
xnor UO_2622 (O_2622,N_29031,N_25637);
and UO_2623 (O_2623,N_27068,N_28014);
and UO_2624 (O_2624,N_29099,N_24817);
nor UO_2625 (O_2625,N_28908,N_27812);
or UO_2626 (O_2626,N_29039,N_29798);
xor UO_2627 (O_2627,N_27165,N_26586);
or UO_2628 (O_2628,N_28225,N_26093);
and UO_2629 (O_2629,N_26129,N_28429);
xnor UO_2630 (O_2630,N_27960,N_24486);
nand UO_2631 (O_2631,N_25607,N_28620);
and UO_2632 (O_2632,N_26412,N_26171);
or UO_2633 (O_2633,N_29405,N_26290);
nand UO_2634 (O_2634,N_25662,N_27982);
or UO_2635 (O_2635,N_27953,N_24389);
nor UO_2636 (O_2636,N_25436,N_29398);
xor UO_2637 (O_2637,N_27834,N_26623);
xnor UO_2638 (O_2638,N_28714,N_26515);
xor UO_2639 (O_2639,N_29572,N_26056);
nand UO_2640 (O_2640,N_27758,N_26053);
or UO_2641 (O_2641,N_24742,N_25267);
and UO_2642 (O_2642,N_28070,N_27595);
nor UO_2643 (O_2643,N_24161,N_27828);
or UO_2644 (O_2644,N_25036,N_25055);
xnor UO_2645 (O_2645,N_29707,N_24880);
and UO_2646 (O_2646,N_26543,N_28349);
xor UO_2647 (O_2647,N_27970,N_28886);
or UO_2648 (O_2648,N_29552,N_27693);
xnor UO_2649 (O_2649,N_25159,N_28061);
nor UO_2650 (O_2650,N_29703,N_27995);
or UO_2651 (O_2651,N_27397,N_26663);
xnor UO_2652 (O_2652,N_26684,N_27018);
nand UO_2653 (O_2653,N_27694,N_29388);
or UO_2654 (O_2654,N_27624,N_27213);
nor UO_2655 (O_2655,N_24601,N_27503);
nor UO_2656 (O_2656,N_24061,N_24288);
nor UO_2657 (O_2657,N_26109,N_28181);
and UO_2658 (O_2658,N_27963,N_28314);
or UO_2659 (O_2659,N_26177,N_26707);
or UO_2660 (O_2660,N_28613,N_25995);
nor UO_2661 (O_2661,N_27743,N_29828);
and UO_2662 (O_2662,N_28129,N_24400);
or UO_2663 (O_2663,N_29597,N_25272);
and UO_2664 (O_2664,N_25941,N_25312);
or UO_2665 (O_2665,N_25259,N_25150);
nor UO_2666 (O_2666,N_27103,N_29392);
xnor UO_2667 (O_2667,N_25294,N_26316);
nand UO_2668 (O_2668,N_28945,N_25009);
nand UO_2669 (O_2669,N_26907,N_25016);
and UO_2670 (O_2670,N_25474,N_26784);
or UO_2671 (O_2671,N_27366,N_24612);
or UO_2672 (O_2672,N_29348,N_29524);
xnor UO_2673 (O_2673,N_24309,N_24676);
nor UO_2674 (O_2674,N_29979,N_28662);
xnor UO_2675 (O_2675,N_27918,N_25711);
or UO_2676 (O_2676,N_24347,N_24549);
and UO_2677 (O_2677,N_28215,N_24091);
and UO_2678 (O_2678,N_29582,N_27774);
or UO_2679 (O_2679,N_25927,N_25508);
nand UO_2680 (O_2680,N_24721,N_29892);
xnor UO_2681 (O_2681,N_26547,N_26390);
or UO_2682 (O_2682,N_28384,N_29613);
xnor UO_2683 (O_2683,N_27039,N_28377);
nand UO_2684 (O_2684,N_28318,N_29773);
or UO_2685 (O_2685,N_28015,N_25169);
or UO_2686 (O_2686,N_28424,N_25540);
nand UO_2687 (O_2687,N_25419,N_24504);
nor UO_2688 (O_2688,N_27388,N_26973);
nor UO_2689 (O_2689,N_28187,N_26730);
xor UO_2690 (O_2690,N_29443,N_24188);
xnor UO_2691 (O_2691,N_25713,N_25391);
nand UO_2692 (O_2692,N_27936,N_27118);
nor UO_2693 (O_2693,N_27126,N_26622);
nor UO_2694 (O_2694,N_28938,N_24206);
or UO_2695 (O_2695,N_25634,N_29984);
xor UO_2696 (O_2696,N_24938,N_28149);
nor UO_2697 (O_2697,N_29076,N_28512);
nor UO_2698 (O_2698,N_24564,N_25161);
and UO_2699 (O_2699,N_25442,N_25694);
xor UO_2700 (O_2700,N_26142,N_29272);
or UO_2701 (O_2701,N_29250,N_26286);
nor UO_2702 (O_2702,N_27083,N_28332);
nand UO_2703 (O_2703,N_26333,N_27861);
or UO_2704 (O_2704,N_25491,N_25386);
or UO_2705 (O_2705,N_26893,N_24899);
nand UO_2706 (O_2706,N_28309,N_25900);
nor UO_2707 (O_2707,N_25382,N_29371);
and UO_2708 (O_2708,N_24113,N_27214);
nand UO_2709 (O_2709,N_27635,N_25282);
and UO_2710 (O_2710,N_27204,N_29177);
and UO_2711 (O_2711,N_27086,N_29716);
nor UO_2712 (O_2712,N_26287,N_24987);
or UO_2713 (O_2713,N_29931,N_28928);
nand UO_2714 (O_2714,N_26273,N_28604);
or UO_2715 (O_2715,N_28802,N_29365);
nand UO_2716 (O_2716,N_27763,N_24897);
and UO_2717 (O_2717,N_26038,N_27378);
nand UO_2718 (O_2718,N_28299,N_25775);
and UO_2719 (O_2719,N_25632,N_29387);
xnor UO_2720 (O_2720,N_29178,N_26891);
and UO_2721 (O_2721,N_28401,N_28829);
xnor UO_2722 (O_2722,N_24284,N_26820);
or UO_2723 (O_2723,N_28224,N_25541);
nor UO_2724 (O_2724,N_27379,N_26518);
xnor UO_2725 (O_2725,N_27135,N_27596);
nor UO_2726 (O_2726,N_25100,N_25933);
and UO_2727 (O_2727,N_28950,N_29484);
nor UO_2728 (O_2728,N_26754,N_28399);
and UO_2729 (O_2729,N_28691,N_29983);
and UO_2730 (O_2730,N_28417,N_25400);
or UO_2731 (O_2731,N_24684,N_25721);
nand UO_2732 (O_2732,N_26011,N_25705);
nand UO_2733 (O_2733,N_26594,N_24740);
and UO_2734 (O_2734,N_28487,N_24949);
nor UO_2735 (O_2735,N_25146,N_28018);
xnor UO_2736 (O_2736,N_24832,N_28083);
nor UO_2737 (O_2737,N_26197,N_29551);
nand UO_2738 (O_2738,N_25919,N_28125);
nor UO_2739 (O_2739,N_25975,N_29577);
and UO_2740 (O_2740,N_29064,N_29156);
xnor UO_2741 (O_2741,N_28119,N_29812);
or UO_2742 (O_2742,N_27123,N_28252);
and UO_2743 (O_2743,N_26875,N_24580);
nor UO_2744 (O_2744,N_28671,N_25736);
and UO_2745 (O_2745,N_28042,N_25019);
or UO_2746 (O_2746,N_28483,N_29694);
nor UO_2747 (O_2747,N_28173,N_29214);
and UO_2748 (O_2748,N_28859,N_25437);
nor UO_2749 (O_2749,N_28806,N_28912);
and UO_2750 (O_2750,N_29680,N_26647);
nand UO_2751 (O_2751,N_24156,N_24005);
or UO_2752 (O_2752,N_24032,N_24002);
nor UO_2753 (O_2753,N_24306,N_28376);
nor UO_2754 (O_2754,N_26018,N_28148);
nand UO_2755 (O_2755,N_24357,N_28651);
nand UO_2756 (O_2756,N_28876,N_29044);
and UO_2757 (O_2757,N_27683,N_24503);
or UO_2758 (O_2758,N_26941,N_26399);
nor UO_2759 (O_2759,N_27967,N_28280);
and UO_2760 (O_2760,N_27160,N_25697);
nand UO_2761 (O_2761,N_26152,N_26553);
nand UO_2762 (O_2762,N_24545,N_29823);
and UO_2763 (O_2763,N_28448,N_24072);
nand UO_2764 (O_2764,N_27469,N_28362);
nor UO_2765 (O_2765,N_25266,N_28852);
or UO_2766 (O_2766,N_25832,N_24386);
nor UO_2767 (O_2767,N_27484,N_24410);
or UO_2768 (O_2768,N_25249,N_28398);
or UO_2769 (O_2769,N_26463,N_27572);
nand UO_2770 (O_2770,N_26240,N_26620);
or UO_2771 (O_2771,N_24671,N_27639);
or UO_2772 (O_2772,N_27321,N_28446);
and UO_2773 (O_2773,N_27517,N_24221);
nor UO_2774 (O_2774,N_25425,N_24067);
and UO_2775 (O_2775,N_25936,N_29801);
xor UO_2776 (O_2776,N_29207,N_26076);
xnor UO_2777 (O_2777,N_25610,N_29738);
and UO_2778 (O_2778,N_27664,N_28936);
nor UO_2779 (O_2779,N_25285,N_26244);
or UO_2780 (O_2780,N_28925,N_26265);
or UO_2781 (O_2781,N_28846,N_27843);
or UO_2782 (O_2782,N_29789,N_27429);
or UO_2783 (O_2783,N_28870,N_26845);
nor UO_2784 (O_2784,N_24393,N_24442);
xor UO_2785 (O_2785,N_25924,N_26179);
nor UO_2786 (O_2786,N_24802,N_29213);
nor UO_2787 (O_2787,N_29274,N_28808);
xnor UO_2788 (O_2788,N_25674,N_25743);
xor UO_2789 (O_2789,N_25059,N_28347);
or UO_2790 (O_2790,N_29237,N_28775);
nor UO_2791 (O_2791,N_27524,N_25983);
and UO_2792 (O_2792,N_24536,N_28607);
xor UO_2793 (O_2793,N_26186,N_28911);
or UO_2794 (O_2794,N_25309,N_26201);
or UO_2795 (O_2795,N_29902,N_27490);
or UO_2796 (O_2796,N_28033,N_29529);
or UO_2797 (O_2797,N_24669,N_26407);
and UO_2798 (O_2798,N_29777,N_25332);
or UO_2799 (O_2799,N_26640,N_26610);
nand UO_2800 (O_2800,N_26705,N_25922);
and UO_2801 (O_2801,N_29333,N_29584);
nand UO_2802 (O_2802,N_24361,N_25098);
nand UO_2803 (O_2803,N_25230,N_24640);
xnor UO_2804 (O_2804,N_26019,N_28548);
xnor UO_2805 (O_2805,N_24989,N_25421);
xor UO_2806 (O_2806,N_27669,N_26225);
or UO_2807 (O_2807,N_27645,N_27734);
nand UO_2808 (O_2808,N_27966,N_29190);
and UO_2809 (O_2809,N_25070,N_27285);
or UO_2810 (O_2810,N_25459,N_28201);
or UO_2811 (O_2811,N_29415,N_25216);
nand UO_2812 (O_2812,N_29135,N_26953);
and UO_2813 (O_2813,N_26787,N_26397);
nor UO_2814 (O_2814,N_24744,N_25035);
or UO_2815 (O_2815,N_25068,N_28414);
nor UO_2816 (O_2816,N_29822,N_24078);
xor UO_2817 (O_2817,N_25811,N_24896);
xnor UO_2818 (O_2818,N_26519,N_27977);
and UO_2819 (O_2819,N_24196,N_29263);
and UO_2820 (O_2820,N_28432,N_27996);
nor UO_2821 (O_2821,N_28365,N_24613);
and UO_2822 (O_2822,N_24840,N_28632);
nand UO_2823 (O_2823,N_29870,N_29435);
and UO_2824 (O_2824,N_29307,N_27001);
nand UO_2825 (O_2825,N_26855,N_25229);
and UO_2826 (O_2826,N_28408,N_24054);
and UO_2827 (O_2827,N_27770,N_27736);
xor UO_2828 (O_2828,N_29412,N_26760);
nor UO_2829 (O_2829,N_27874,N_29430);
nand UO_2830 (O_2830,N_24468,N_25760);
or UO_2831 (O_2831,N_24825,N_29231);
nand UO_2832 (O_2832,N_27820,N_27899);
or UO_2833 (O_2833,N_25631,N_29089);
xor UO_2834 (O_2834,N_29437,N_28922);
nor UO_2835 (O_2835,N_28240,N_29294);
xnor UO_2836 (O_2836,N_28122,N_25042);
nand UO_2837 (O_2837,N_27811,N_25972);
nor UO_2838 (O_2838,N_29820,N_27253);
and UO_2839 (O_2839,N_27920,N_25641);
nand UO_2840 (O_2840,N_26726,N_25619);
or UO_2841 (O_2841,N_28940,N_26715);
nand UO_2842 (O_2842,N_24407,N_28606);
nand UO_2843 (O_2843,N_24812,N_29378);
and UO_2844 (O_2844,N_24530,N_28037);
nor UO_2845 (O_2845,N_27962,N_26307);
nor UO_2846 (O_2846,N_24650,N_25351);
nor UO_2847 (O_2847,N_26701,N_28719);
nor UO_2848 (O_2848,N_27383,N_27612);
nor UO_2849 (O_2849,N_26599,N_25201);
and UO_2850 (O_2850,N_28404,N_27398);
xor UO_2851 (O_2851,N_29885,N_25387);
nand UO_2852 (O_2852,N_24319,N_29176);
or UO_2853 (O_2853,N_28885,N_28216);
xor UO_2854 (O_2854,N_29282,N_27003);
nor UO_2855 (O_2855,N_28563,N_24484);
xor UO_2856 (O_2856,N_28626,N_28202);
nor UO_2857 (O_2857,N_29375,N_27203);
nor UO_2858 (O_2858,N_25142,N_25018);
or UO_2859 (O_2859,N_28904,N_24826);
nand UO_2860 (O_2860,N_29146,N_24883);
nor UO_2861 (O_2861,N_29549,N_26406);
and UO_2862 (O_2862,N_24420,N_24056);
or UO_2863 (O_2863,N_26002,N_24487);
and UO_2864 (O_2864,N_29151,N_24120);
nand UO_2865 (O_2865,N_27211,N_24931);
xor UO_2866 (O_2866,N_24320,N_25854);
xor UO_2867 (O_2867,N_24000,N_26236);
xor UO_2868 (O_2868,N_26937,N_26889);
and UO_2869 (O_2869,N_28657,N_24917);
and UO_2870 (O_2870,N_27697,N_26385);
nor UO_2871 (O_2871,N_26558,N_24064);
nor UO_2872 (O_2872,N_27892,N_28748);
and UO_2873 (O_2873,N_27183,N_28236);
nand UO_2874 (O_2874,N_25613,N_24482);
nor UO_2875 (O_2875,N_29113,N_29646);
or UO_2876 (O_2876,N_27277,N_29669);
or UO_2877 (O_2877,N_27549,N_25440);
or UO_2878 (O_2878,N_24009,N_28457);
xnor UO_2879 (O_2879,N_24326,N_27046);
xor UO_2880 (O_2880,N_24364,N_29782);
and UO_2881 (O_2881,N_26483,N_28178);
nor UO_2882 (O_2882,N_24748,N_24888);
or UO_2883 (O_2883,N_27076,N_28725);
nand UO_2884 (O_2884,N_25569,N_24768);
nor UO_2885 (O_2885,N_27346,N_29547);
and UO_2886 (O_2886,N_27867,N_27074);
nand UO_2887 (O_2887,N_25826,N_27908);
xnor UO_2888 (O_2888,N_24500,N_29204);
xor UO_2889 (O_2889,N_26522,N_28920);
nor UO_2890 (O_2890,N_29765,N_25979);
nand UO_2891 (O_2891,N_28794,N_25287);
xnor UO_2892 (O_2892,N_26792,N_25815);
nor UO_2893 (O_2893,N_24126,N_26691);
nor UO_2894 (O_2894,N_27653,N_28242);
nand UO_2895 (O_2895,N_25487,N_27650);
and UO_2896 (O_2896,N_26358,N_24451);
nor UO_2897 (O_2897,N_24979,N_26498);
nor UO_2898 (O_2898,N_24328,N_27112);
nand UO_2899 (O_2899,N_27729,N_27476);
or UO_2900 (O_2900,N_25997,N_27901);
xnor UO_2901 (O_2901,N_27943,N_25901);
xnor UO_2902 (O_2902,N_25664,N_28340);
and UO_2903 (O_2903,N_24641,N_24034);
xor UO_2904 (O_2904,N_26897,N_24519);
nand UO_2905 (O_2905,N_28672,N_28345);
nor UO_2906 (O_2906,N_25572,N_29854);
and UO_2907 (O_2907,N_27350,N_27371);
nor UO_2908 (O_2908,N_26890,N_25293);
nor UO_2909 (O_2909,N_28601,N_27950);
or UO_2910 (O_2910,N_24584,N_28373);
nor UO_2911 (O_2911,N_24964,N_24454);
or UO_2912 (O_2912,N_28979,N_26856);
or UO_2913 (O_2913,N_24758,N_28147);
nand UO_2914 (O_2914,N_26484,N_28353);
or UO_2915 (O_2915,N_27505,N_26993);
xor UO_2916 (O_2916,N_25319,N_27627);
or UO_2917 (O_2917,N_24098,N_29840);
nor UO_2918 (O_2918,N_25802,N_24729);
or UO_2919 (O_2919,N_25696,N_29711);
or UO_2920 (O_2920,N_25950,N_24070);
and UO_2921 (O_2921,N_25733,N_26103);
and UO_2922 (O_2922,N_28285,N_26434);
or UO_2923 (O_2923,N_29884,N_26071);
nor UO_2924 (O_2924,N_26166,N_25151);
xnor UO_2925 (O_2925,N_29275,N_26077);
xor UO_2926 (O_2926,N_29209,N_26528);
nand UO_2927 (O_2927,N_25501,N_27916);
or UO_2928 (O_2928,N_24587,N_24289);
and UO_2929 (O_2929,N_24384,N_28821);
and UO_2930 (O_2930,N_27136,N_27178);
nand UO_2931 (O_2931,N_24658,N_29318);
or UO_2932 (O_2932,N_26755,N_25578);
nor UO_2933 (O_2933,N_24168,N_29511);
nor UO_2934 (O_2934,N_29363,N_24082);
and UO_2935 (O_2935,N_26775,N_29936);
or UO_2936 (O_2936,N_25560,N_26830);
or UO_2937 (O_2937,N_24175,N_26887);
nand UO_2938 (O_2938,N_28241,N_26429);
nor UO_2939 (O_2939,N_28102,N_28472);
and UO_2940 (O_2940,N_26101,N_24558);
or UO_2941 (O_2941,N_28970,N_27146);
or UO_2942 (O_2942,N_26860,N_29832);
and UO_2943 (O_2943,N_28586,N_29011);
nor UO_2944 (O_2944,N_26957,N_28508);
or UO_2945 (O_2945,N_24597,N_28123);
nand UO_2946 (O_2946,N_27987,N_28445);
and UO_2947 (O_2947,N_27658,N_28801);
or UO_2948 (O_2948,N_25961,N_28440);
and UO_2949 (O_2949,N_29460,N_27796);
and UO_2950 (O_2950,N_29692,N_27489);
nor UO_2951 (O_2951,N_28545,N_28611);
nand UO_2952 (O_2952,N_27715,N_27762);
or UO_2953 (O_2953,N_25526,N_24390);
and UO_2954 (O_2954,N_27452,N_29610);
nand UO_2955 (O_2955,N_27060,N_25724);
nor UO_2956 (O_2956,N_28661,N_24085);
xor UO_2957 (O_2957,N_26354,N_26900);
xnor UO_2958 (O_2958,N_25840,N_24932);
xor UO_2959 (O_2959,N_24855,N_26905);
nand UO_2960 (O_2960,N_28759,N_29875);
nand UO_2961 (O_2961,N_28639,N_28835);
and UO_2962 (O_2962,N_25571,N_29122);
nand UO_2963 (O_2963,N_24351,N_29166);
and UO_2964 (O_2964,N_26852,N_26940);
or UO_2965 (O_2965,N_25781,N_28550);
and UO_2966 (O_2966,N_24099,N_29744);
nor UO_2967 (O_2967,N_25904,N_27522);
nor UO_2968 (O_2968,N_24477,N_26282);
xor UO_2969 (O_2969,N_25991,N_26600);
or UO_2970 (O_2970,N_26781,N_28221);
or UO_2971 (O_2971,N_28467,N_29356);
nand UO_2972 (O_2972,N_28433,N_27170);
nand UO_2973 (O_2973,N_25101,N_29485);
xor UO_2974 (O_2974,N_29629,N_24173);
and UO_2975 (O_2975,N_26000,N_28008);
nor UO_2976 (O_2976,N_28617,N_26467);
nand UO_2977 (O_2977,N_28305,N_28126);
nand UO_2978 (O_2978,N_28341,N_29316);
nor UO_2979 (O_2979,N_27075,N_25839);
or UO_2980 (O_2980,N_28871,N_27166);
nor UO_2981 (O_2981,N_24922,N_27917);
and UO_2982 (O_2982,N_25772,N_25044);
and UO_2983 (O_2983,N_29834,N_25148);
xnor UO_2984 (O_2984,N_29571,N_28412);
xnor UO_2985 (O_2985,N_27990,N_26394);
or UO_2986 (O_2986,N_28504,N_25496);
and UO_2987 (O_2987,N_27432,N_28041);
or UO_2988 (O_2988,N_27772,N_26337);
nor UO_2989 (O_2989,N_27502,N_24995);
nor UO_2990 (O_2990,N_28841,N_24757);
xor UO_2991 (O_2991,N_28720,N_26759);
and UO_2992 (O_2992,N_24141,N_28010);
nand UO_2993 (O_2993,N_25446,N_29935);
nand UO_2994 (O_2994,N_27594,N_26426);
nand UO_2995 (O_2995,N_26100,N_27994);
and UO_2996 (O_2996,N_25301,N_27884);
nor UO_2997 (O_2997,N_28697,N_28188);
xor UO_2998 (O_2998,N_26516,N_28059);
and UO_2999 (O_2999,N_25618,N_27526);
and UO_3000 (O_3000,N_29617,N_26708);
xor UO_3001 (O_3001,N_24336,N_24746);
nand UO_3002 (O_3002,N_25713,N_29237);
xor UO_3003 (O_3003,N_29506,N_27815);
xnor UO_3004 (O_3004,N_28011,N_26843);
nand UO_3005 (O_3005,N_28294,N_27530);
or UO_3006 (O_3006,N_26335,N_24838);
and UO_3007 (O_3007,N_26839,N_27040);
nand UO_3008 (O_3008,N_27987,N_27168);
nor UO_3009 (O_3009,N_25622,N_27214);
xnor UO_3010 (O_3010,N_27248,N_25656);
and UO_3011 (O_3011,N_29890,N_28030);
nor UO_3012 (O_3012,N_26347,N_25062);
or UO_3013 (O_3013,N_25175,N_29710);
nand UO_3014 (O_3014,N_26049,N_24111);
xnor UO_3015 (O_3015,N_28555,N_26394);
nand UO_3016 (O_3016,N_26394,N_25631);
xor UO_3017 (O_3017,N_27771,N_26027);
xor UO_3018 (O_3018,N_25830,N_29923);
and UO_3019 (O_3019,N_24045,N_27819);
xnor UO_3020 (O_3020,N_27558,N_25027);
nor UO_3021 (O_3021,N_28016,N_27446);
xor UO_3022 (O_3022,N_25870,N_27148);
nand UO_3023 (O_3023,N_25618,N_25126);
or UO_3024 (O_3024,N_25337,N_24309);
nand UO_3025 (O_3025,N_24705,N_27968);
xor UO_3026 (O_3026,N_25892,N_27439);
xnor UO_3027 (O_3027,N_24602,N_28586);
nor UO_3028 (O_3028,N_24412,N_27525);
xnor UO_3029 (O_3029,N_24499,N_25235);
or UO_3030 (O_3030,N_29715,N_28588);
and UO_3031 (O_3031,N_28480,N_24687);
or UO_3032 (O_3032,N_29947,N_24637);
and UO_3033 (O_3033,N_29912,N_28864);
and UO_3034 (O_3034,N_29366,N_26016);
nor UO_3035 (O_3035,N_29206,N_26726);
xor UO_3036 (O_3036,N_25373,N_26044);
or UO_3037 (O_3037,N_24616,N_28376);
and UO_3038 (O_3038,N_28435,N_28315);
nor UO_3039 (O_3039,N_29667,N_25280);
and UO_3040 (O_3040,N_24931,N_29469);
nor UO_3041 (O_3041,N_25611,N_29979);
nand UO_3042 (O_3042,N_25585,N_27511);
nor UO_3043 (O_3043,N_24141,N_29152);
xnor UO_3044 (O_3044,N_25822,N_26115);
xnor UO_3045 (O_3045,N_28336,N_29148);
nor UO_3046 (O_3046,N_27703,N_27527);
nor UO_3047 (O_3047,N_27068,N_26416);
nand UO_3048 (O_3048,N_26897,N_28919);
xor UO_3049 (O_3049,N_24116,N_25863);
nor UO_3050 (O_3050,N_29887,N_27080);
or UO_3051 (O_3051,N_24892,N_28596);
nor UO_3052 (O_3052,N_29291,N_29559);
xnor UO_3053 (O_3053,N_27106,N_27703);
or UO_3054 (O_3054,N_26365,N_28189);
nand UO_3055 (O_3055,N_27264,N_27560);
nand UO_3056 (O_3056,N_25699,N_29624);
xnor UO_3057 (O_3057,N_28194,N_28230);
and UO_3058 (O_3058,N_24138,N_25704);
or UO_3059 (O_3059,N_26982,N_27360);
and UO_3060 (O_3060,N_28117,N_24767);
nor UO_3061 (O_3061,N_28137,N_28522);
nor UO_3062 (O_3062,N_26582,N_24658);
nand UO_3063 (O_3063,N_27075,N_29832);
nand UO_3064 (O_3064,N_29159,N_28365);
nand UO_3065 (O_3065,N_24730,N_25180);
nand UO_3066 (O_3066,N_26770,N_24055);
and UO_3067 (O_3067,N_29270,N_29763);
or UO_3068 (O_3068,N_24220,N_26911);
nor UO_3069 (O_3069,N_28201,N_27987);
nor UO_3070 (O_3070,N_28646,N_25081);
xor UO_3071 (O_3071,N_24342,N_25165);
and UO_3072 (O_3072,N_27395,N_25105);
or UO_3073 (O_3073,N_26968,N_24070);
xnor UO_3074 (O_3074,N_25861,N_29066);
and UO_3075 (O_3075,N_24334,N_26919);
nand UO_3076 (O_3076,N_29105,N_25212);
and UO_3077 (O_3077,N_25367,N_24293);
nand UO_3078 (O_3078,N_27671,N_28171);
nand UO_3079 (O_3079,N_29467,N_29789);
nand UO_3080 (O_3080,N_25073,N_25147);
nor UO_3081 (O_3081,N_28541,N_25828);
nor UO_3082 (O_3082,N_27710,N_29763);
xnor UO_3083 (O_3083,N_29173,N_28955);
nor UO_3084 (O_3084,N_24836,N_29777);
nand UO_3085 (O_3085,N_29586,N_28136);
xor UO_3086 (O_3086,N_24676,N_24870);
nor UO_3087 (O_3087,N_28074,N_26114);
and UO_3088 (O_3088,N_29021,N_28239);
nor UO_3089 (O_3089,N_27004,N_25757);
nor UO_3090 (O_3090,N_27583,N_25139);
xor UO_3091 (O_3091,N_25581,N_28352);
xor UO_3092 (O_3092,N_26238,N_26866);
or UO_3093 (O_3093,N_28173,N_27228);
or UO_3094 (O_3094,N_24846,N_29414);
nor UO_3095 (O_3095,N_25848,N_24705);
or UO_3096 (O_3096,N_26446,N_26618);
and UO_3097 (O_3097,N_26505,N_27092);
nor UO_3098 (O_3098,N_27864,N_28628);
nand UO_3099 (O_3099,N_27641,N_27322);
nor UO_3100 (O_3100,N_27897,N_24048);
xnor UO_3101 (O_3101,N_27334,N_27766);
or UO_3102 (O_3102,N_29126,N_24416);
nand UO_3103 (O_3103,N_27066,N_26115);
nor UO_3104 (O_3104,N_29575,N_26417);
and UO_3105 (O_3105,N_25666,N_26362);
nand UO_3106 (O_3106,N_25758,N_26468);
nor UO_3107 (O_3107,N_29201,N_27415);
or UO_3108 (O_3108,N_29154,N_24171);
nand UO_3109 (O_3109,N_28202,N_26590);
and UO_3110 (O_3110,N_24040,N_28029);
xor UO_3111 (O_3111,N_27893,N_29811);
nor UO_3112 (O_3112,N_25952,N_25269);
nor UO_3113 (O_3113,N_24807,N_29932);
xor UO_3114 (O_3114,N_29650,N_28436);
nor UO_3115 (O_3115,N_29477,N_24524);
or UO_3116 (O_3116,N_29635,N_24858);
or UO_3117 (O_3117,N_27422,N_28763);
nand UO_3118 (O_3118,N_24508,N_29816);
nand UO_3119 (O_3119,N_29376,N_26294);
nor UO_3120 (O_3120,N_29140,N_26969);
nand UO_3121 (O_3121,N_29990,N_25504);
nand UO_3122 (O_3122,N_25102,N_26438);
or UO_3123 (O_3123,N_24361,N_28057);
or UO_3124 (O_3124,N_28356,N_28847);
nor UO_3125 (O_3125,N_26614,N_25814);
or UO_3126 (O_3126,N_24560,N_28845);
and UO_3127 (O_3127,N_29671,N_27039);
xnor UO_3128 (O_3128,N_26778,N_29653);
and UO_3129 (O_3129,N_24929,N_27251);
and UO_3130 (O_3130,N_29900,N_29869);
nor UO_3131 (O_3131,N_27642,N_29527);
nand UO_3132 (O_3132,N_29875,N_25962);
nand UO_3133 (O_3133,N_27635,N_25131);
xor UO_3134 (O_3134,N_26302,N_29497);
and UO_3135 (O_3135,N_24196,N_28543);
or UO_3136 (O_3136,N_25839,N_26402);
nand UO_3137 (O_3137,N_27075,N_24924);
and UO_3138 (O_3138,N_26083,N_28007);
xnor UO_3139 (O_3139,N_25172,N_24294);
nand UO_3140 (O_3140,N_26790,N_27474);
or UO_3141 (O_3141,N_26817,N_29128);
or UO_3142 (O_3142,N_25843,N_27562);
or UO_3143 (O_3143,N_25985,N_28938);
or UO_3144 (O_3144,N_28026,N_27953);
xnor UO_3145 (O_3145,N_28212,N_27825);
nor UO_3146 (O_3146,N_29344,N_29857);
xor UO_3147 (O_3147,N_28501,N_24271);
and UO_3148 (O_3148,N_25191,N_25726);
and UO_3149 (O_3149,N_26755,N_25395);
nand UO_3150 (O_3150,N_26539,N_25880);
xnor UO_3151 (O_3151,N_27372,N_24558);
or UO_3152 (O_3152,N_27367,N_25267);
nor UO_3153 (O_3153,N_24556,N_27822);
and UO_3154 (O_3154,N_24456,N_27911);
and UO_3155 (O_3155,N_29568,N_24186);
and UO_3156 (O_3156,N_29911,N_27113);
xnor UO_3157 (O_3157,N_28386,N_26542);
nor UO_3158 (O_3158,N_24105,N_29308);
nand UO_3159 (O_3159,N_29229,N_28129);
and UO_3160 (O_3160,N_25895,N_24926);
nand UO_3161 (O_3161,N_24216,N_25928);
or UO_3162 (O_3162,N_24779,N_28864);
and UO_3163 (O_3163,N_26667,N_29623);
nor UO_3164 (O_3164,N_29839,N_29152);
xor UO_3165 (O_3165,N_28874,N_29804);
nor UO_3166 (O_3166,N_26468,N_29158);
or UO_3167 (O_3167,N_29489,N_26247);
nand UO_3168 (O_3168,N_24359,N_28883);
and UO_3169 (O_3169,N_28659,N_24617);
nand UO_3170 (O_3170,N_26942,N_24441);
nor UO_3171 (O_3171,N_27659,N_25784);
nand UO_3172 (O_3172,N_24092,N_25829);
or UO_3173 (O_3173,N_27663,N_27951);
or UO_3174 (O_3174,N_25085,N_28997);
xnor UO_3175 (O_3175,N_27042,N_25521);
nand UO_3176 (O_3176,N_24258,N_24074);
or UO_3177 (O_3177,N_25734,N_26914);
nand UO_3178 (O_3178,N_25171,N_25286);
nor UO_3179 (O_3179,N_27767,N_25238);
xor UO_3180 (O_3180,N_25704,N_26687);
nand UO_3181 (O_3181,N_25870,N_27457);
nand UO_3182 (O_3182,N_29924,N_24430);
and UO_3183 (O_3183,N_27263,N_27819);
nor UO_3184 (O_3184,N_27880,N_25872);
nand UO_3185 (O_3185,N_25232,N_27705);
and UO_3186 (O_3186,N_25430,N_28446);
or UO_3187 (O_3187,N_29345,N_27815);
nand UO_3188 (O_3188,N_24408,N_24958);
and UO_3189 (O_3189,N_29265,N_26472);
or UO_3190 (O_3190,N_27150,N_29409);
xor UO_3191 (O_3191,N_26916,N_26232);
or UO_3192 (O_3192,N_26856,N_24448);
nor UO_3193 (O_3193,N_24325,N_26390);
or UO_3194 (O_3194,N_26398,N_24136);
and UO_3195 (O_3195,N_25727,N_24731);
and UO_3196 (O_3196,N_29729,N_26734);
nand UO_3197 (O_3197,N_29654,N_27691);
xor UO_3198 (O_3198,N_29648,N_28700);
and UO_3199 (O_3199,N_25591,N_26751);
nor UO_3200 (O_3200,N_28527,N_29928);
nor UO_3201 (O_3201,N_27899,N_29015);
xor UO_3202 (O_3202,N_28423,N_28215);
xor UO_3203 (O_3203,N_29783,N_24879);
nor UO_3204 (O_3204,N_28049,N_29739);
nand UO_3205 (O_3205,N_27251,N_28552);
nor UO_3206 (O_3206,N_26683,N_28913);
or UO_3207 (O_3207,N_28873,N_27675);
xnor UO_3208 (O_3208,N_24209,N_29723);
or UO_3209 (O_3209,N_28493,N_28458);
or UO_3210 (O_3210,N_26538,N_26315);
nand UO_3211 (O_3211,N_25890,N_26776);
xor UO_3212 (O_3212,N_29414,N_29801);
nand UO_3213 (O_3213,N_29393,N_25441);
nand UO_3214 (O_3214,N_24883,N_29853);
or UO_3215 (O_3215,N_24358,N_28856);
and UO_3216 (O_3216,N_27845,N_28146);
xor UO_3217 (O_3217,N_29255,N_24012);
xnor UO_3218 (O_3218,N_28093,N_29057);
and UO_3219 (O_3219,N_28528,N_25813);
or UO_3220 (O_3220,N_27683,N_29974);
and UO_3221 (O_3221,N_26391,N_24978);
and UO_3222 (O_3222,N_29942,N_26649);
xnor UO_3223 (O_3223,N_25002,N_29723);
or UO_3224 (O_3224,N_26534,N_29817);
or UO_3225 (O_3225,N_25819,N_25059);
xnor UO_3226 (O_3226,N_27090,N_24553);
xnor UO_3227 (O_3227,N_24903,N_27998);
or UO_3228 (O_3228,N_24435,N_26078);
or UO_3229 (O_3229,N_26261,N_24882);
and UO_3230 (O_3230,N_26505,N_26859);
nor UO_3231 (O_3231,N_28497,N_24901);
nor UO_3232 (O_3232,N_26506,N_27457);
nand UO_3233 (O_3233,N_25164,N_26715);
xnor UO_3234 (O_3234,N_24211,N_27118);
or UO_3235 (O_3235,N_25507,N_29659);
nand UO_3236 (O_3236,N_28938,N_28437);
and UO_3237 (O_3237,N_24056,N_27569);
or UO_3238 (O_3238,N_28773,N_29129);
nand UO_3239 (O_3239,N_25827,N_29048);
nor UO_3240 (O_3240,N_25525,N_27290);
and UO_3241 (O_3241,N_28845,N_25167);
xnor UO_3242 (O_3242,N_26790,N_25293);
or UO_3243 (O_3243,N_24345,N_29358);
nor UO_3244 (O_3244,N_24914,N_27193);
nand UO_3245 (O_3245,N_25450,N_29781);
nor UO_3246 (O_3246,N_29064,N_26252);
nand UO_3247 (O_3247,N_24653,N_24804);
xnor UO_3248 (O_3248,N_25626,N_27339);
or UO_3249 (O_3249,N_27618,N_25804);
xor UO_3250 (O_3250,N_28364,N_25652);
nand UO_3251 (O_3251,N_25541,N_26323);
and UO_3252 (O_3252,N_29497,N_29595);
nand UO_3253 (O_3253,N_29374,N_29093);
and UO_3254 (O_3254,N_26061,N_25595);
xnor UO_3255 (O_3255,N_26077,N_28059);
xnor UO_3256 (O_3256,N_25472,N_28781);
and UO_3257 (O_3257,N_26727,N_26987);
or UO_3258 (O_3258,N_29538,N_27932);
or UO_3259 (O_3259,N_25196,N_29259);
nor UO_3260 (O_3260,N_24768,N_28392);
xnor UO_3261 (O_3261,N_29415,N_26536);
or UO_3262 (O_3262,N_29965,N_26108);
and UO_3263 (O_3263,N_26331,N_24530);
xor UO_3264 (O_3264,N_29258,N_29167);
or UO_3265 (O_3265,N_27882,N_26731);
and UO_3266 (O_3266,N_26376,N_27270);
nor UO_3267 (O_3267,N_25255,N_25484);
xnor UO_3268 (O_3268,N_27252,N_29390);
xnor UO_3269 (O_3269,N_28001,N_27784);
and UO_3270 (O_3270,N_24650,N_25224);
nor UO_3271 (O_3271,N_27559,N_26477);
xor UO_3272 (O_3272,N_28450,N_29194);
and UO_3273 (O_3273,N_26209,N_25855);
and UO_3274 (O_3274,N_26907,N_27615);
xnor UO_3275 (O_3275,N_26404,N_29306);
and UO_3276 (O_3276,N_29802,N_27280);
nand UO_3277 (O_3277,N_25229,N_28141);
nand UO_3278 (O_3278,N_24992,N_28969);
nor UO_3279 (O_3279,N_25628,N_24995);
or UO_3280 (O_3280,N_26296,N_25545);
nor UO_3281 (O_3281,N_26193,N_27197);
and UO_3282 (O_3282,N_24245,N_26156);
xor UO_3283 (O_3283,N_24363,N_25763);
nand UO_3284 (O_3284,N_28665,N_28196);
or UO_3285 (O_3285,N_28641,N_28482);
nor UO_3286 (O_3286,N_25452,N_28002);
and UO_3287 (O_3287,N_27074,N_25820);
nand UO_3288 (O_3288,N_28470,N_29244);
nand UO_3289 (O_3289,N_27564,N_28371);
xnor UO_3290 (O_3290,N_24402,N_24858);
nand UO_3291 (O_3291,N_25043,N_28070);
or UO_3292 (O_3292,N_29185,N_24445);
nor UO_3293 (O_3293,N_29589,N_29953);
nor UO_3294 (O_3294,N_28943,N_24913);
or UO_3295 (O_3295,N_26557,N_24850);
and UO_3296 (O_3296,N_26471,N_28596);
nor UO_3297 (O_3297,N_26177,N_26892);
xnor UO_3298 (O_3298,N_26237,N_29627);
nand UO_3299 (O_3299,N_25755,N_28214);
and UO_3300 (O_3300,N_29654,N_27662);
and UO_3301 (O_3301,N_25716,N_28487);
or UO_3302 (O_3302,N_28284,N_29159);
nand UO_3303 (O_3303,N_27006,N_29140);
or UO_3304 (O_3304,N_27275,N_27840);
or UO_3305 (O_3305,N_26200,N_26331);
xnor UO_3306 (O_3306,N_29950,N_29192);
nand UO_3307 (O_3307,N_29495,N_25411);
and UO_3308 (O_3308,N_26676,N_26595);
nand UO_3309 (O_3309,N_25206,N_28791);
nor UO_3310 (O_3310,N_28012,N_25415);
or UO_3311 (O_3311,N_28637,N_28909);
nor UO_3312 (O_3312,N_27344,N_25025);
nor UO_3313 (O_3313,N_29067,N_27815);
nand UO_3314 (O_3314,N_24294,N_28010);
or UO_3315 (O_3315,N_28497,N_27532);
nand UO_3316 (O_3316,N_27783,N_29676);
nor UO_3317 (O_3317,N_28080,N_29460);
or UO_3318 (O_3318,N_26455,N_27691);
nor UO_3319 (O_3319,N_25069,N_29807);
or UO_3320 (O_3320,N_24286,N_26887);
nand UO_3321 (O_3321,N_28543,N_26751);
nand UO_3322 (O_3322,N_24796,N_28469);
nand UO_3323 (O_3323,N_27565,N_28713);
nor UO_3324 (O_3324,N_27555,N_27488);
and UO_3325 (O_3325,N_26986,N_28792);
or UO_3326 (O_3326,N_26937,N_25913);
and UO_3327 (O_3327,N_29054,N_27832);
or UO_3328 (O_3328,N_24804,N_27434);
and UO_3329 (O_3329,N_28347,N_26136);
nor UO_3330 (O_3330,N_26839,N_29375);
xnor UO_3331 (O_3331,N_24627,N_25657);
nor UO_3332 (O_3332,N_24453,N_29791);
or UO_3333 (O_3333,N_29417,N_27019);
or UO_3334 (O_3334,N_29700,N_27862);
or UO_3335 (O_3335,N_28802,N_25612);
nor UO_3336 (O_3336,N_25709,N_27426);
and UO_3337 (O_3337,N_27614,N_27881);
xnor UO_3338 (O_3338,N_27218,N_26896);
and UO_3339 (O_3339,N_27487,N_27695);
or UO_3340 (O_3340,N_25047,N_28431);
xnor UO_3341 (O_3341,N_24367,N_25461);
nor UO_3342 (O_3342,N_26490,N_24945);
nor UO_3343 (O_3343,N_25475,N_29021);
nand UO_3344 (O_3344,N_28433,N_27522);
or UO_3345 (O_3345,N_29500,N_28102);
nand UO_3346 (O_3346,N_24620,N_28214);
or UO_3347 (O_3347,N_28601,N_29719);
or UO_3348 (O_3348,N_25746,N_25846);
and UO_3349 (O_3349,N_25649,N_29861);
and UO_3350 (O_3350,N_28924,N_27235);
xnor UO_3351 (O_3351,N_24429,N_24768);
nand UO_3352 (O_3352,N_26762,N_25334);
nor UO_3353 (O_3353,N_24553,N_26305);
xnor UO_3354 (O_3354,N_25879,N_26087);
nand UO_3355 (O_3355,N_28326,N_27659);
nor UO_3356 (O_3356,N_29676,N_26486);
or UO_3357 (O_3357,N_25453,N_29486);
nor UO_3358 (O_3358,N_27407,N_29830);
or UO_3359 (O_3359,N_27327,N_28926);
xor UO_3360 (O_3360,N_24618,N_28700);
or UO_3361 (O_3361,N_28182,N_27816);
xor UO_3362 (O_3362,N_25462,N_26958);
nand UO_3363 (O_3363,N_25560,N_26272);
and UO_3364 (O_3364,N_29539,N_26115);
xor UO_3365 (O_3365,N_28692,N_27642);
nand UO_3366 (O_3366,N_24945,N_27482);
nor UO_3367 (O_3367,N_26456,N_25814);
xor UO_3368 (O_3368,N_26169,N_27658);
and UO_3369 (O_3369,N_26764,N_25095);
nor UO_3370 (O_3370,N_26192,N_29549);
nand UO_3371 (O_3371,N_28243,N_29323);
or UO_3372 (O_3372,N_27322,N_24569);
nor UO_3373 (O_3373,N_26320,N_25076);
xor UO_3374 (O_3374,N_27177,N_26855);
nor UO_3375 (O_3375,N_25253,N_25189);
xnor UO_3376 (O_3376,N_25381,N_24580);
or UO_3377 (O_3377,N_24278,N_29418);
and UO_3378 (O_3378,N_28136,N_27322);
nor UO_3379 (O_3379,N_24718,N_26740);
xnor UO_3380 (O_3380,N_24664,N_24077);
or UO_3381 (O_3381,N_27406,N_28839);
nor UO_3382 (O_3382,N_28946,N_26241);
nor UO_3383 (O_3383,N_25331,N_27609);
or UO_3384 (O_3384,N_26319,N_26611);
nor UO_3385 (O_3385,N_26314,N_29842);
xor UO_3386 (O_3386,N_29682,N_26796);
nand UO_3387 (O_3387,N_26364,N_26648);
xor UO_3388 (O_3388,N_25348,N_25544);
and UO_3389 (O_3389,N_25364,N_29837);
nor UO_3390 (O_3390,N_24316,N_24925);
or UO_3391 (O_3391,N_26943,N_25702);
or UO_3392 (O_3392,N_25855,N_29257);
or UO_3393 (O_3393,N_26254,N_24552);
and UO_3394 (O_3394,N_27551,N_27411);
nand UO_3395 (O_3395,N_28498,N_24741);
nand UO_3396 (O_3396,N_28129,N_28043);
xor UO_3397 (O_3397,N_24332,N_25833);
nand UO_3398 (O_3398,N_25395,N_28505);
or UO_3399 (O_3399,N_25055,N_27929);
or UO_3400 (O_3400,N_25812,N_29264);
or UO_3401 (O_3401,N_25221,N_28393);
or UO_3402 (O_3402,N_28637,N_27021);
xnor UO_3403 (O_3403,N_27469,N_29825);
or UO_3404 (O_3404,N_29712,N_28990);
and UO_3405 (O_3405,N_27475,N_26382);
nor UO_3406 (O_3406,N_29017,N_29079);
xnor UO_3407 (O_3407,N_26334,N_29662);
xnor UO_3408 (O_3408,N_29970,N_24917);
nand UO_3409 (O_3409,N_24356,N_25876);
nor UO_3410 (O_3410,N_24805,N_25136);
nor UO_3411 (O_3411,N_26360,N_27843);
and UO_3412 (O_3412,N_24694,N_25430);
nand UO_3413 (O_3413,N_26432,N_26927);
and UO_3414 (O_3414,N_25735,N_29542);
nor UO_3415 (O_3415,N_24719,N_28142);
xor UO_3416 (O_3416,N_26710,N_29651);
nand UO_3417 (O_3417,N_27270,N_28878);
xor UO_3418 (O_3418,N_29051,N_27559);
xnor UO_3419 (O_3419,N_29147,N_29056);
xor UO_3420 (O_3420,N_25966,N_27755);
xnor UO_3421 (O_3421,N_25438,N_26627);
xnor UO_3422 (O_3422,N_28341,N_28707);
xor UO_3423 (O_3423,N_29303,N_27608);
xnor UO_3424 (O_3424,N_27695,N_26131);
nand UO_3425 (O_3425,N_29007,N_28781);
and UO_3426 (O_3426,N_28468,N_27269);
xor UO_3427 (O_3427,N_29294,N_28340);
nor UO_3428 (O_3428,N_25024,N_25615);
and UO_3429 (O_3429,N_24840,N_26641);
nor UO_3430 (O_3430,N_26480,N_25596);
or UO_3431 (O_3431,N_27536,N_26561);
and UO_3432 (O_3432,N_26283,N_27321);
nand UO_3433 (O_3433,N_29243,N_29821);
nand UO_3434 (O_3434,N_24748,N_28311);
xnor UO_3435 (O_3435,N_25016,N_29379);
nor UO_3436 (O_3436,N_27834,N_27905);
and UO_3437 (O_3437,N_24215,N_28048);
xnor UO_3438 (O_3438,N_26685,N_26340);
or UO_3439 (O_3439,N_27003,N_24406);
xor UO_3440 (O_3440,N_24940,N_28349);
nor UO_3441 (O_3441,N_28274,N_27234);
or UO_3442 (O_3442,N_25432,N_27280);
xor UO_3443 (O_3443,N_29427,N_29400);
or UO_3444 (O_3444,N_29279,N_29629);
nand UO_3445 (O_3445,N_29426,N_24283);
nor UO_3446 (O_3446,N_26005,N_27582);
or UO_3447 (O_3447,N_25993,N_27744);
nor UO_3448 (O_3448,N_29227,N_29209);
or UO_3449 (O_3449,N_25914,N_26057);
nor UO_3450 (O_3450,N_24304,N_29694);
xnor UO_3451 (O_3451,N_24373,N_25164);
nor UO_3452 (O_3452,N_26978,N_26587);
nor UO_3453 (O_3453,N_25640,N_27392);
or UO_3454 (O_3454,N_29448,N_27988);
nand UO_3455 (O_3455,N_26164,N_27176);
nor UO_3456 (O_3456,N_28474,N_28051);
xor UO_3457 (O_3457,N_29639,N_28769);
or UO_3458 (O_3458,N_27089,N_25586);
or UO_3459 (O_3459,N_29517,N_27927);
and UO_3460 (O_3460,N_24237,N_28478);
and UO_3461 (O_3461,N_26328,N_28734);
nand UO_3462 (O_3462,N_25808,N_26683);
or UO_3463 (O_3463,N_24988,N_29381);
xor UO_3464 (O_3464,N_26039,N_29720);
or UO_3465 (O_3465,N_28920,N_24122);
nor UO_3466 (O_3466,N_25693,N_26169);
and UO_3467 (O_3467,N_27991,N_25505);
and UO_3468 (O_3468,N_24844,N_26750);
xnor UO_3469 (O_3469,N_24080,N_29343);
and UO_3470 (O_3470,N_28084,N_27028);
and UO_3471 (O_3471,N_25401,N_26579);
and UO_3472 (O_3472,N_28786,N_24635);
xor UO_3473 (O_3473,N_24190,N_28004);
nand UO_3474 (O_3474,N_28232,N_25075);
xor UO_3475 (O_3475,N_24542,N_26379);
or UO_3476 (O_3476,N_29339,N_27238);
or UO_3477 (O_3477,N_28402,N_28456);
and UO_3478 (O_3478,N_29556,N_25548);
or UO_3479 (O_3479,N_29322,N_27669);
xnor UO_3480 (O_3480,N_29304,N_28519);
nor UO_3481 (O_3481,N_26948,N_28985);
and UO_3482 (O_3482,N_26853,N_26519);
or UO_3483 (O_3483,N_25321,N_24181);
nor UO_3484 (O_3484,N_29290,N_27272);
or UO_3485 (O_3485,N_29358,N_24330);
nand UO_3486 (O_3486,N_29682,N_29426);
nand UO_3487 (O_3487,N_28435,N_27445);
xnor UO_3488 (O_3488,N_28600,N_24752);
xor UO_3489 (O_3489,N_29265,N_28088);
nand UO_3490 (O_3490,N_29701,N_25881);
nor UO_3491 (O_3491,N_28625,N_26920);
nor UO_3492 (O_3492,N_24173,N_27807);
nor UO_3493 (O_3493,N_28388,N_26132);
nand UO_3494 (O_3494,N_25166,N_26555);
or UO_3495 (O_3495,N_24451,N_24494);
and UO_3496 (O_3496,N_24635,N_24250);
nor UO_3497 (O_3497,N_26269,N_26724);
xor UO_3498 (O_3498,N_28068,N_29404);
nor UO_3499 (O_3499,N_25213,N_26133);
endmodule