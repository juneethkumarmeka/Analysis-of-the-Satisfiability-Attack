module basic_500_3000_500_4_levels_2xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_352,In_203);
and U1 (N_1,In_291,In_226);
and U2 (N_2,In_403,In_234);
nand U3 (N_3,In_386,In_258);
nor U4 (N_4,In_330,In_428);
and U5 (N_5,In_444,In_223);
and U6 (N_6,In_96,In_20);
or U7 (N_7,In_70,In_237);
and U8 (N_8,In_365,In_450);
or U9 (N_9,In_212,In_174);
nor U10 (N_10,In_303,In_170);
nor U11 (N_11,In_209,In_60);
and U12 (N_12,In_111,In_16);
or U13 (N_13,In_133,In_270);
and U14 (N_14,In_77,In_24);
or U15 (N_15,In_478,In_231);
or U16 (N_16,In_85,In_221);
nand U17 (N_17,In_206,In_198);
and U18 (N_18,In_371,In_317);
nand U19 (N_19,In_287,In_192);
nor U20 (N_20,In_254,In_94);
or U21 (N_21,In_479,In_344);
nor U22 (N_22,In_440,In_361);
or U23 (N_23,In_435,In_416);
xor U24 (N_24,In_281,In_137);
and U25 (N_25,In_54,In_50);
and U26 (N_26,In_56,In_393);
or U27 (N_27,In_306,In_417);
nor U28 (N_28,In_342,In_454);
or U29 (N_29,In_229,In_296);
or U30 (N_30,In_114,In_484);
nor U31 (N_31,In_61,In_336);
xor U32 (N_32,In_405,In_482);
xor U33 (N_33,In_183,In_280);
and U34 (N_34,In_29,In_156);
nand U35 (N_35,In_489,In_272);
and U36 (N_36,In_49,In_292);
and U37 (N_37,In_164,In_193);
or U38 (N_38,In_414,In_463);
nor U39 (N_39,In_123,In_62);
nand U40 (N_40,In_278,In_112);
nand U41 (N_41,In_87,In_233);
nand U42 (N_42,In_172,In_390);
and U43 (N_43,In_9,In_260);
or U44 (N_44,In_468,In_238);
and U45 (N_45,In_487,In_132);
or U46 (N_46,In_73,In_201);
nand U47 (N_47,In_411,In_255);
xnor U48 (N_48,In_488,In_169);
nor U49 (N_49,In_316,In_297);
xor U50 (N_50,In_438,In_18);
or U51 (N_51,In_309,In_93);
or U52 (N_52,In_301,In_419);
and U53 (N_53,In_415,In_437);
or U54 (N_54,In_376,In_124);
and U55 (N_55,In_245,In_101);
and U56 (N_56,In_285,In_339);
nand U57 (N_57,In_40,In_109);
and U58 (N_58,In_353,In_471);
or U59 (N_59,In_293,In_145);
and U60 (N_60,In_214,In_436);
and U61 (N_61,In_65,In_88);
nor U62 (N_62,In_373,In_263);
nand U63 (N_63,In_240,In_89);
and U64 (N_64,In_474,In_10);
nand U65 (N_65,In_224,In_477);
or U66 (N_66,In_154,In_149);
and U67 (N_67,In_429,In_117);
or U68 (N_68,In_422,In_141);
nor U69 (N_69,In_208,In_199);
and U70 (N_70,In_322,In_462);
nand U71 (N_71,In_79,In_75);
nand U72 (N_72,In_74,In_467);
nor U73 (N_73,In_447,In_289);
and U74 (N_74,In_387,In_91);
nor U75 (N_75,In_381,In_290);
and U76 (N_76,In_497,In_485);
nand U77 (N_77,In_247,In_34);
nand U78 (N_78,In_37,In_396);
nor U79 (N_79,In_51,In_104);
and U80 (N_80,In_142,In_496);
or U81 (N_81,In_143,In_335);
xnor U82 (N_82,In_358,In_125);
nand U83 (N_83,In_299,In_446);
or U84 (N_84,In_7,In_211);
or U85 (N_85,In_173,In_312);
nor U86 (N_86,In_443,In_210);
nor U87 (N_87,In_399,In_98);
nor U88 (N_88,In_315,In_307);
or U89 (N_89,In_304,In_458);
or U90 (N_90,In_434,In_346);
nand U91 (N_91,In_266,In_4);
nand U92 (N_92,In_323,In_286);
and U93 (N_93,In_2,In_242);
and U94 (N_94,In_382,In_385);
nand U95 (N_95,In_194,In_432);
nand U96 (N_96,In_81,In_42);
or U97 (N_97,In_216,In_340);
or U98 (N_98,In_155,In_269);
and U99 (N_99,In_333,In_480);
or U100 (N_100,In_57,In_261);
nand U101 (N_101,In_159,In_179);
or U102 (N_102,In_107,In_384);
or U103 (N_103,In_433,In_134);
nand U104 (N_104,In_265,In_425);
nor U105 (N_105,In_113,In_118);
or U106 (N_106,In_59,In_162);
and U107 (N_107,In_197,In_354);
or U108 (N_108,In_310,In_64);
or U109 (N_109,In_185,In_146);
nand U110 (N_110,In_95,In_486);
nand U111 (N_111,In_383,In_439);
or U112 (N_112,In_102,In_465);
nand U113 (N_113,In_232,In_168);
or U114 (N_114,In_298,In_391);
nand U115 (N_115,In_115,In_319);
xor U116 (N_116,In_246,In_476);
nand U117 (N_117,In_327,In_41);
or U118 (N_118,In_110,In_69);
and U119 (N_119,In_348,In_318);
or U120 (N_120,In_122,In_239);
or U121 (N_121,In_460,In_218);
nand U122 (N_122,In_495,In_499);
nand U123 (N_123,In_464,In_11);
nand U124 (N_124,In_186,In_128);
and U125 (N_125,In_167,In_19);
and U126 (N_126,In_369,In_175);
nor U127 (N_127,In_15,In_267);
and U128 (N_128,In_82,In_288);
or U129 (N_129,In_99,In_401);
nand U130 (N_130,In_235,In_0);
nor U131 (N_131,In_47,In_129);
nand U132 (N_132,In_324,In_375);
nor U133 (N_133,In_135,In_320);
nand U134 (N_134,In_283,In_359);
nand U135 (N_135,In_308,In_31);
nand U136 (N_136,In_248,In_329);
nor U137 (N_137,In_53,In_470);
nand U138 (N_138,In_268,In_1);
or U139 (N_139,In_420,In_282);
and U140 (N_140,In_103,In_328);
or U141 (N_141,In_138,In_380);
nor U142 (N_142,In_48,In_427);
nor U143 (N_143,In_347,In_448);
and U144 (N_144,In_338,In_35);
nand U145 (N_145,In_400,In_230);
nand U146 (N_146,In_372,In_351);
or U147 (N_147,In_204,In_127);
nand U148 (N_148,In_84,In_368);
or U149 (N_149,In_55,In_356);
or U150 (N_150,In_38,In_334);
nor U151 (N_151,In_457,In_68);
or U152 (N_152,In_116,In_357);
nand U153 (N_153,In_426,In_161);
nand U154 (N_154,In_46,In_295);
or U155 (N_155,In_26,In_139);
nor U156 (N_156,In_219,In_189);
and U157 (N_157,In_452,In_475);
and U158 (N_158,In_313,In_314);
or U159 (N_159,In_473,In_466);
or U160 (N_160,In_350,In_195);
or U161 (N_161,In_408,In_120);
and U162 (N_162,In_6,In_3);
nand U163 (N_163,In_284,In_39);
or U164 (N_164,In_273,In_367);
nand U165 (N_165,In_58,In_152);
nor U166 (N_166,In_241,In_483);
nor U167 (N_167,In_166,In_196);
and U168 (N_168,In_184,In_147);
nor U169 (N_169,In_325,In_366);
and U170 (N_170,In_188,In_92);
nor U171 (N_171,In_126,In_459);
or U172 (N_172,In_326,In_8);
and U173 (N_173,In_407,In_72);
nor U174 (N_174,In_337,In_277);
or U175 (N_175,In_250,In_131);
or U176 (N_176,In_136,In_43);
xor U177 (N_177,In_63,In_52);
and U178 (N_178,In_395,In_181);
or U179 (N_179,In_397,In_345);
nand U180 (N_180,In_205,In_431);
or U181 (N_181,In_171,In_244);
and U182 (N_182,In_378,In_424);
nand U183 (N_183,In_341,In_22);
nor U184 (N_184,In_17,In_412);
nor U185 (N_185,In_418,In_76);
nor U186 (N_186,In_461,In_274);
or U187 (N_187,In_153,In_360);
and U188 (N_188,In_481,In_182);
and U189 (N_189,In_157,In_349);
or U190 (N_190,In_493,In_392);
nor U191 (N_191,In_388,In_30);
or U192 (N_192,In_236,In_5);
nor U193 (N_193,In_97,In_86);
and U194 (N_194,In_321,In_445);
nand U195 (N_195,In_449,In_442);
and U196 (N_196,In_33,In_302);
or U197 (N_197,In_222,In_413);
or U198 (N_198,In_90,In_121);
or U199 (N_199,In_25,In_264);
nand U200 (N_200,In_27,In_108);
and U201 (N_201,In_398,In_377);
nor U202 (N_202,In_472,In_28);
nand U203 (N_203,In_441,In_490);
nand U204 (N_204,In_191,In_67);
nand U205 (N_205,In_355,In_259);
nand U206 (N_206,In_176,In_410);
nand U207 (N_207,In_163,In_379);
and U208 (N_208,In_332,In_178);
nor U209 (N_209,In_256,In_374);
and U210 (N_210,In_225,In_343);
and U211 (N_211,In_331,In_144);
or U212 (N_212,In_491,In_311);
nand U213 (N_213,In_305,In_119);
nand U214 (N_214,In_430,In_423);
xnor U215 (N_215,In_220,In_498);
or U216 (N_216,In_249,In_421);
or U217 (N_217,In_370,In_217);
or U218 (N_218,In_300,In_409);
nor U219 (N_219,In_394,In_207);
nor U220 (N_220,In_213,In_243);
nor U221 (N_221,In_364,In_215);
nand U222 (N_222,In_228,In_100);
or U223 (N_223,In_12,In_23);
and U224 (N_224,In_494,In_252);
or U225 (N_225,In_80,In_389);
and U226 (N_226,In_492,In_202);
and U227 (N_227,In_177,In_151);
and U228 (N_228,In_13,In_251);
nor U229 (N_229,In_158,In_451);
and U230 (N_230,In_14,In_402);
nor U231 (N_231,In_190,In_130);
or U232 (N_232,In_83,In_406);
and U233 (N_233,In_404,In_456);
nor U234 (N_234,In_275,In_105);
or U235 (N_235,In_453,In_362);
and U236 (N_236,In_44,In_227);
nor U237 (N_237,In_21,In_36);
nor U238 (N_238,In_45,In_140);
nand U239 (N_239,In_148,In_262);
nor U240 (N_240,In_32,In_71);
nand U241 (N_241,In_279,In_150);
and U242 (N_242,In_106,In_271);
nor U243 (N_243,In_180,In_455);
nor U244 (N_244,In_187,In_253);
nor U245 (N_245,In_257,In_294);
xor U246 (N_246,In_469,In_66);
nand U247 (N_247,In_160,In_165);
or U248 (N_248,In_276,In_363);
or U249 (N_249,In_200,In_78);
or U250 (N_250,In_141,In_2);
and U251 (N_251,In_297,In_24);
nand U252 (N_252,In_114,In_166);
and U253 (N_253,In_67,In_293);
nand U254 (N_254,In_21,In_468);
and U255 (N_255,In_315,In_493);
or U256 (N_256,In_494,In_340);
nand U257 (N_257,In_415,In_281);
nand U258 (N_258,In_183,In_417);
nor U259 (N_259,In_321,In_150);
nor U260 (N_260,In_318,In_453);
nand U261 (N_261,In_121,In_326);
nand U262 (N_262,In_196,In_35);
and U263 (N_263,In_280,In_205);
nand U264 (N_264,In_184,In_74);
nor U265 (N_265,In_15,In_394);
nand U266 (N_266,In_170,In_240);
or U267 (N_267,In_212,In_73);
or U268 (N_268,In_236,In_225);
nand U269 (N_269,In_371,In_11);
or U270 (N_270,In_430,In_336);
and U271 (N_271,In_162,In_396);
nor U272 (N_272,In_200,In_287);
nand U273 (N_273,In_108,In_483);
or U274 (N_274,In_263,In_241);
nor U275 (N_275,In_375,In_480);
nand U276 (N_276,In_472,In_461);
or U277 (N_277,In_304,In_103);
and U278 (N_278,In_453,In_78);
nor U279 (N_279,In_243,In_54);
and U280 (N_280,In_10,In_236);
and U281 (N_281,In_161,In_29);
nand U282 (N_282,In_110,In_336);
xnor U283 (N_283,In_295,In_131);
and U284 (N_284,In_496,In_327);
nand U285 (N_285,In_114,In_314);
or U286 (N_286,In_11,In_204);
and U287 (N_287,In_436,In_321);
nor U288 (N_288,In_476,In_41);
and U289 (N_289,In_464,In_149);
nor U290 (N_290,In_477,In_345);
nor U291 (N_291,In_347,In_250);
nand U292 (N_292,In_102,In_63);
or U293 (N_293,In_207,In_434);
xnor U294 (N_294,In_281,In_59);
nor U295 (N_295,In_243,In_140);
and U296 (N_296,In_139,In_459);
nand U297 (N_297,In_453,In_293);
and U298 (N_298,In_32,In_110);
and U299 (N_299,In_360,In_216);
or U300 (N_300,In_59,In_239);
or U301 (N_301,In_28,In_157);
and U302 (N_302,In_351,In_211);
and U303 (N_303,In_41,In_111);
nor U304 (N_304,In_303,In_142);
or U305 (N_305,In_169,In_438);
nand U306 (N_306,In_323,In_183);
nand U307 (N_307,In_56,In_45);
and U308 (N_308,In_224,In_108);
or U309 (N_309,In_55,In_267);
nor U310 (N_310,In_318,In_75);
and U311 (N_311,In_286,In_220);
or U312 (N_312,In_116,In_478);
or U313 (N_313,In_61,In_280);
and U314 (N_314,In_140,In_40);
or U315 (N_315,In_149,In_333);
or U316 (N_316,In_362,In_356);
or U317 (N_317,In_244,In_37);
nand U318 (N_318,In_340,In_97);
nor U319 (N_319,In_378,In_318);
or U320 (N_320,In_498,In_301);
xor U321 (N_321,In_299,In_339);
and U322 (N_322,In_179,In_10);
nor U323 (N_323,In_53,In_371);
and U324 (N_324,In_363,In_129);
and U325 (N_325,In_382,In_374);
nor U326 (N_326,In_90,In_357);
nand U327 (N_327,In_391,In_357);
or U328 (N_328,In_312,In_46);
and U329 (N_329,In_423,In_288);
nand U330 (N_330,In_168,In_384);
nand U331 (N_331,In_80,In_353);
nor U332 (N_332,In_67,In_59);
nand U333 (N_333,In_481,In_132);
nor U334 (N_334,In_311,In_206);
nand U335 (N_335,In_350,In_398);
nand U336 (N_336,In_380,In_403);
nor U337 (N_337,In_446,In_448);
or U338 (N_338,In_278,In_232);
nand U339 (N_339,In_347,In_51);
or U340 (N_340,In_122,In_487);
or U341 (N_341,In_305,In_209);
nor U342 (N_342,In_438,In_2);
or U343 (N_343,In_132,In_189);
nor U344 (N_344,In_481,In_493);
nor U345 (N_345,In_203,In_407);
and U346 (N_346,In_484,In_266);
and U347 (N_347,In_399,In_247);
and U348 (N_348,In_212,In_204);
or U349 (N_349,In_132,In_383);
nand U350 (N_350,In_172,In_436);
nand U351 (N_351,In_206,In_425);
nand U352 (N_352,In_359,In_404);
and U353 (N_353,In_172,In_220);
nor U354 (N_354,In_326,In_181);
nor U355 (N_355,In_357,In_416);
nor U356 (N_356,In_70,In_6);
nor U357 (N_357,In_165,In_231);
nor U358 (N_358,In_361,In_64);
nand U359 (N_359,In_363,In_279);
xnor U360 (N_360,In_203,In_367);
and U361 (N_361,In_325,In_387);
and U362 (N_362,In_377,In_154);
nor U363 (N_363,In_167,In_468);
or U364 (N_364,In_406,In_159);
and U365 (N_365,In_152,In_91);
and U366 (N_366,In_56,In_441);
or U367 (N_367,In_265,In_419);
or U368 (N_368,In_410,In_15);
nor U369 (N_369,In_229,In_383);
nor U370 (N_370,In_452,In_300);
nor U371 (N_371,In_447,In_378);
xor U372 (N_372,In_484,In_130);
nor U373 (N_373,In_150,In_313);
nor U374 (N_374,In_413,In_111);
nand U375 (N_375,In_164,In_331);
nand U376 (N_376,In_300,In_285);
nand U377 (N_377,In_64,In_407);
and U378 (N_378,In_465,In_187);
nand U379 (N_379,In_174,In_315);
or U380 (N_380,In_398,In_267);
nor U381 (N_381,In_245,In_44);
or U382 (N_382,In_419,In_260);
nand U383 (N_383,In_443,In_128);
or U384 (N_384,In_78,In_302);
or U385 (N_385,In_156,In_112);
nor U386 (N_386,In_112,In_362);
nand U387 (N_387,In_415,In_215);
and U388 (N_388,In_496,In_385);
and U389 (N_389,In_176,In_412);
or U390 (N_390,In_292,In_148);
and U391 (N_391,In_33,In_232);
or U392 (N_392,In_61,In_84);
xor U393 (N_393,In_41,In_291);
nand U394 (N_394,In_452,In_388);
nand U395 (N_395,In_498,In_181);
nor U396 (N_396,In_248,In_499);
and U397 (N_397,In_387,In_132);
nand U398 (N_398,In_133,In_135);
or U399 (N_399,In_320,In_13);
and U400 (N_400,In_267,In_397);
and U401 (N_401,In_268,In_113);
or U402 (N_402,In_137,In_115);
nor U403 (N_403,In_444,In_148);
or U404 (N_404,In_489,In_216);
xor U405 (N_405,In_238,In_117);
nor U406 (N_406,In_486,In_48);
and U407 (N_407,In_0,In_444);
nor U408 (N_408,In_287,In_354);
nor U409 (N_409,In_141,In_307);
or U410 (N_410,In_146,In_281);
nor U411 (N_411,In_157,In_86);
nand U412 (N_412,In_84,In_40);
or U413 (N_413,In_393,In_64);
and U414 (N_414,In_420,In_312);
and U415 (N_415,In_452,In_376);
and U416 (N_416,In_106,In_378);
and U417 (N_417,In_383,In_282);
or U418 (N_418,In_467,In_85);
or U419 (N_419,In_92,In_65);
and U420 (N_420,In_15,In_149);
and U421 (N_421,In_56,In_347);
and U422 (N_422,In_34,In_58);
and U423 (N_423,In_296,In_286);
or U424 (N_424,In_217,In_469);
nor U425 (N_425,In_283,In_222);
nor U426 (N_426,In_347,In_271);
nand U427 (N_427,In_329,In_174);
nor U428 (N_428,In_251,In_189);
nor U429 (N_429,In_230,In_85);
or U430 (N_430,In_351,In_265);
nor U431 (N_431,In_44,In_204);
and U432 (N_432,In_63,In_196);
or U433 (N_433,In_43,In_317);
and U434 (N_434,In_40,In_227);
xor U435 (N_435,In_294,In_398);
or U436 (N_436,In_139,In_120);
nor U437 (N_437,In_481,In_306);
nand U438 (N_438,In_72,In_129);
nor U439 (N_439,In_236,In_80);
nand U440 (N_440,In_107,In_50);
nand U441 (N_441,In_137,In_97);
nor U442 (N_442,In_279,In_405);
or U443 (N_443,In_229,In_270);
xor U444 (N_444,In_247,In_102);
xor U445 (N_445,In_227,In_199);
and U446 (N_446,In_197,In_467);
or U447 (N_447,In_67,In_229);
nand U448 (N_448,In_366,In_209);
nor U449 (N_449,In_258,In_62);
or U450 (N_450,In_360,In_176);
nand U451 (N_451,In_332,In_31);
and U452 (N_452,In_265,In_481);
or U453 (N_453,In_172,In_121);
and U454 (N_454,In_351,In_0);
nand U455 (N_455,In_255,In_160);
and U456 (N_456,In_58,In_414);
xor U457 (N_457,In_349,In_50);
nand U458 (N_458,In_493,In_103);
or U459 (N_459,In_186,In_460);
nand U460 (N_460,In_237,In_67);
or U461 (N_461,In_285,In_484);
and U462 (N_462,In_156,In_6);
nand U463 (N_463,In_363,In_418);
nor U464 (N_464,In_288,In_334);
nand U465 (N_465,In_113,In_26);
nand U466 (N_466,In_161,In_160);
nand U467 (N_467,In_419,In_342);
or U468 (N_468,In_198,In_422);
and U469 (N_469,In_208,In_69);
and U470 (N_470,In_431,In_369);
and U471 (N_471,In_464,In_349);
or U472 (N_472,In_362,In_179);
nor U473 (N_473,In_164,In_362);
and U474 (N_474,In_398,In_91);
nand U475 (N_475,In_108,In_131);
xnor U476 (N_476,In_223,In_237);
nand U477 (N_477,In_19,In_97);
or U478 (N_478,In_242,In_73);
or U479 (N_479,In_124,In_63);
xor U480 (N_480,In_95,In_424);
nor U481 (N_481,In_8,In_192);
or U482 (N_482,In_270,In_286);
nand U483 (N_483,In_436,In_222);
and U484 (N_484,In_111,In_499);
nand U485 (N_485,In_417,In_292);
and U486 (N_486,In_50,In_65);
nor U487 (N_487,In_213,In_183);
nor U488 (N_488,In_316,In_403);
nor U489 (N_489,In_354,In_459);
nor U490 (N_490,In_415,In_204);
nand U491 (N_491,In_497,In_186);
or U492 (N_492,In_156,In_257);
or U493 (N_493,In_499,In_465);
nand U494 (N_494,In_197,In_31);
or U495 (N_495,In_328,In_195);
or U496 (N_496,In_270,In_136);
nor U497 (N_497,In_82,In_140);
and U498 (N_498,In_173,In_150);
and U499 (N_499,In_131,In_178);
nor U500 (N_500,In_400,In_177);
nor U501 (N_501,In_271,In_342);
or U502 (N_502,In_132,In_183);
nand U503 (N_503,In_219,In_272);
nor U504 (N_504,In_63,In_28);
or U505 (N_505,In_175,In_313);
or U506 (N_506,In_328,In_433);
or U507 (N_507,In_347,In_281);
nor U508 (N_508,In_244,In_450);
nand U509 (N_509,In_308,In_248);
and U510 (N_510,In_285,In_68);
and U511 (N_511,In_416,In_388);
and U512 (N_512,In_241,In_136);
nand U513 (N_513,In_300,In_442);
or U514 (N_514,In_392,In_322);
xor U515 (N_515,In_38,In_298);
nor U516 (N_516,In_212,In_317);
and U517 (N_517,In_307,In_191);
and U518 (N_518,In_128,In_87);
and U519 (N_519,In_440,In_359);
and U520 (N_520,In_442,In_17);
and U521 (N_521,In_2,In_313);
nand U522 (N_522,In_304,In_362);
or U523 (N_523,In_464,In_282);
and U524 (N_524,In_90,In_226);
and U525 (N_525,In_30,In_355);
and U526 (N_526,In_223,In_360);
and U527 (N_527,In_50,In_236);
or U528 (N_528,In_249,In_447);
nor U529 (N_529,In_405,In_445);
and U530 (N_530,In_104,In_27);
nand U531 (N_531,In_392,In_109);
nor U532 (N_532,In_6,In_271);
or U533 (N_533,In_466,In_102);
and U534 (N_534,In_13,In_228);
and U535 (N_535,In_359,In_103);
or U536 (N_536,In_75,In_222);
or U537 (N_537,In_429,In_332);
xnor U538 (N_538,In_399,In_429);
and U539 (N_539,In_283,In_298);
or U540 (N_540,In_402,In_87);
nor U541 (N_541,In_142,In_328);
or U542 (N_542,In_184,In_1);
and U543 (N_543,In_133,In_54);
nor U544 (N_544,In_240,In_325);
or U545 (N_545,In_185,In_460);
nand U546 (N_546,In_310,In_75);
or U547 (N_547,In_150,In_291);
or U548 (N_548,In_452,In_33);
nor U549 (N_549,In_42,In_79);
nor U550 (N_550,In_200,In_427);
nand U551 (N_551,In_363,In_431);
nand U552 (N_552,In_437,In_391);
and U553 (N_553,In_256,In_385);
nor U554 (N_554,In_254,In_380);
nand U555 (N_555,In_364,In_57);
nand U556 (N_556,In_210,In_368);
nor U557 (N_557,In_400,In_174);
and U558 (N_558,In_224,In_253);
and U559 (N_559,In_312,In_59);
or U560 (N_560,In_115,In_269);
nand U561 (N_561,In_15,In_269);
or U562 (N_562,In_181,In_388);
nor U563 (N_563,In_441,In_129);
nand U564 (N_564,In_364,In_359);
nand U565 (N_565,In_153,In_272);
and U566 (N_566,In_338,In_236);
nand U567 (N_567,In_224,In_393);
or U568 (N_568,In_414,In_8);
nor U569 (N_569,In_39,In_130);
and U570 (N_570,In_344,In_194);
and U571 (N_571,In_278,In_48);
and U572 (N_572,In_130,In_410);
nand U573 (N_573,In_224,In_390);
nor U574 (N_574,In_215,In_284);
nand U575 (N_575,In_471,In_309);
and U576 (N_576,In_358,In_351);
or U577 (N_577,In_261,In_288);
and U578 (N_578,In_370,In_110);
nor U579 (N_579,In_138,In_445);
nor U580 (N_580,In_67,In_31);
and U581 (N_581,In_109,In_182);
nand U582 (N_582,In_468,In_426);
or U583 (N_583,In_317,In_386);
nand U584 (N_584,In_11,In_52);
or U585 (N_585,In_34,In_35);
or U586 (N_586,In_133,In_349);
or U587 (N_587,In_407,In_417);
or U588 (N_588,In_83,In_442);
or U589 (N_589,In_469,In_410);
nor U590 (N_590,In_476,In_208);
nor U591 (N_591,In_272,In_216);
and U592 (N_592,In_422,In_54);
or U593 (N_593,In_434,In_59);
and U594 (N_594,In_281,In_205);
and U595 (N_595,In_450,In_397);
or U596 (N_596,In_499,In_264);
nand U597 (N_597,In_371,In_48);
or U598 (N_598,In_165,In_492);
and U599 (N_599,In_475,In_461);
nor U600 (N_600,In_428,In_376);
or U601 (N_601,In_250,In_143);
and U602 (N_602,In_129,In_285);
nand U603 (N_603,In_480,In_149);
or U604 (N_604,In_265,In_422);
or U605 (N_605,In_142,In_492);
nand U606 (N_606,In_98,In_190);
or U607 (N_607,In_104,In_209);
or U608 (N_608,In_354,In_12);
nor U609 (N_609,In_7,In_430);
and U610 (N_610,In_351,In_60);
nor U611 (N_611,In_326,In_85);
or U612 (N_612,In_250,In_9);
and U613 (N_613,In_304,In_376);
nand U614 (N_614,In_39,In_278);
nand U615 (N_615,In_11,In_286);
nor U616 (N_616,In_5,In_209);
or U617 (N_617,In_358,In_111);
nor U618 (N_618,In_410,In_482);
or U619 (N_619,In_104,In_303);
or U620 (N_620,In_447,In_179);
and U621 (N_621,In_134,In_369);
nor U622 (N_622,In_250,In_374);
or U623 (N_623,In_239,In_332);
nor U624 (N_624,In_58,In_269);
nor U625 (N_625,In_299,In_67);
nor U626 (N_626,In_155,In_25);
or U627 (N_627,In_318,In_476);
xor U628 (N_628,In_36,In_192);
nand U629 (N_629,In_130,In_411);
or U630 (N_630,In_434,In_125);
nor U631 (N_631,In_218,In_96);
and U632 (N_632,In_208,In_380);
or U633 (N_633,In_207,In_31);
nand U634 (N_634,In_160,In_208);
or U635 (N_635,In_199,In_469);
nor U636 (N_636,In_275,In_360);
and U637 (N_637,In_357,In_398);
or U638 (N_638,In_309,In_135);
nand U639 (N_639,In_426,In_203);
nor U640 (N_640,In_5,In_382);
or U641 (N_641,In_114,In_208);
nand U642 (N_642,In_385,In_86);
or U643 (N_643,In_11,In_330);
nor U644 (N_644,In_441,In_231);
nor U645 (N_645,In_420,In_83);
nand U646 (N_646,In_33,In_142);
or U647 (N_647,In_123,In_266);
nand U648 (N_648,In_186,In_239);
nand U649 (N_649,In_394,In_105);
or U650 (N_650,In_86,In_401);
nand U651 (N_651,In_336,In_287);
or U652 (N_652,In_399,In_218);
and U653 (N_653,In_271,In_368);
and U654 (N_654,In_138,In_347);
nand U655 (N_655,In_324,In_346);
or U656 (N_656,In_473,In_210);
nor U657 (N_657,In_69,In_374);
nand U658 (N_658,In_155,In_48);
nand U659 (N_659,In_433,In_256);
nand U660 (N_660,In_150,In_413);
or U661 (N_661,In_106,In_17);
or U662 (N_662,In_499,In_405);
and U663 (N_663,In_405,In_175);
and U664 (N_664,In_145,In_155);
nand U665 (N_665,In_346,In_235);
xnor U666 (N_666,In_392,In_6);
nor U667 (N_667,In_99,In_237);
nor U668 (N_668,In_457,In_469);
and U669 (N_669,In_210,In_304);
nor U670 (N_670,In_289,In_473);
nor U671 (N_671,In_40,In_306);
and U672 (N_672,In_226,In_456);
nor U673 (N_673,In_450,In_377);
nor U674 (N_674,In_211,In_269);
nor U675 (N_675,In_162,In_186);
or U676 (N_676,In_268,In_261);
nor U677 (N_677,In_61,In_342);
and U678 (N_678,In_378,In_328);
or U679 (N_679,In_196,In_57);
or U680 (N_680,In_170,In_103);
nand U681 (N_681,In_263,In_362);
xnor U682 (N_682,In_120,In_326);
or U683 (N_683,In_238,In_10);
nor U684 (N_684,In_464,In_77);
nand U685 (N_685,In_479,In_140);
nor U686 (N_686,In_445,In_290);
nor U687 (N_687,In_282,In_372);
or U688 (N_688,In_15,In_8);
or U689 (N_689,In_342,In_136);
and U690 (N_690,In_355,In_304);
and U691 (N_691,In_229,In_69);
nor U692 (N_692,In_78,In_193);
or U693 (N_693,In_429,In_191);
nor U694 (N_694,In_58,In_364);
and U695 (N_695,In_150,In_121);
xor U696 (N_696,In_483,In_224);
nand U697 (N_697,In_467,In_306);
and U698 (N_698,In_295,In_130);
nor U699 (N_699,In_437,In_461);
nor U700 (N_700,In_475,In_17);
nand U701 (N_701,In_33,In_278);
or U702 (N_702,In_296,In_278);
nand U703 (N_703,In_240,In_152);
or U704 (N_704,In_349,In_352);
nor U705 (N_705,In_356,In_188);
and U706 (N_706,In_96,In_466);
nand U707 (N_707,In_116,In_199);
or U708 (N_708,In_353,In_115);
nor U709 (N_709,In_267,In_152);
or U710 (N_710,In_443,In_248);
nand U711 (N_711,In_440,In_419);
nand U712 (N_712,In_225,In_147);
xnor U713 (N_713,In_346,In_313);
and U714 (N_714,In_356,In_464);
nor U715 (N_715,In_250,In_453);
and U716 (N_716,In_321,In_399);
nand U717 (N_717,In_440,In_110);
nand U718 (N_718,In_174,In_82);
nand U719 (N_719,In_158,In_129);
and U720 (N_720,In_130,In_442);
or U721 (N_721,In_311,In_5);
nand U722 (N_722,In_213,In_189);
and U723 (N_723,In_97,In_3);
nand U724 (N_724,In_437,In_427);
and U725 (N_725,In_427,In_246);
or U726 (N_726,In_88,In_29);
nand U727 (N_727,In_92,In_11);
nand U728 (N_728,In_85,In_349);
or U729 (N_729,In_231,In_249);
nand U730 (N_730,In_191,In_21);
and U731 (N_731,In_217,In_479);
nand U732 (N_732,In_482,In_325);
or U733 (N_733,In_108,In_207);
nor U734 (N_734,In_248,In_220);
and U735 (N_735,In_201,In_336);
nor U736 (N_736,In_488,In_111);
nor U737 (N_737,In_97,In_458);
nand U738 (N_738,In_157,In_490);
or U739 (N_739,In_144,In_481);
or U740 (N_740,In_434,In_286);
or U741 (N_741,In_271,In_144);
nor U742 (N_742,In_300,In_209);
and U743 (N_743,In_29,In_185);
nand U744 (N_744,In_46,In_304);
nand U745 (N_745,In_346,In_205);
and U746 (N_746,In_240,In_69);
nor U747 (N_747,In_419,In_105);
or U748 (N_748,In_135,In_102);
or U749 (N_749,In_1,In_122);
or U750 (N_750,N_221,N_238);
nor U751 (N_751,N_374,N_470);
and U752 (N_752,N_542,N_688);
xnor U753 (N_753,N_19,N_117);
nor U754 (N_754,N_497,N_725);
nor U755 (N_755,N_595,N_434);
nor U756 (N_756,N_426,N_367);
or U757 (N_757,N_586,N_445);
nand U758 (N_758,N_175,N_342);
or U759 (N_759,N_50,N_600);
nand U760 (N_760,N_546,N_483);
nor U761 (N_761,N_641,N_333);
nor U762 (N_762,N_89,N_160);
and U763 (N_763,N_745,N_419);
xnor U764 (N_764,N_505,N_601);
nand U765 (N_765,N_414,N_158);
and U766 (N_766,N_576,N_711);
or U767 (N_767,N_695,N_39);
or U768 (N_768,N_727,N_194);
or U769 (N_769,N_61,N_170);
or U770 (N_770,N_480,N_197);
or U771 (N_771,N_616,N_612);
nor U772 (N_772,N_569,N_491);
nor U773 (N_773,N_555,N_473);
nor U774 (N_774,N_114,N_351);
and U775 (N_775,N_326,N_495);
or U776 (N_776,N_732,N_359);
nor U777 (N_777,N_609,N_206);
or U778 (N_778,N_185,N_211);
nor U779 (N_779,N_412,N_369);
nand U780 (N_780,N_111,N_715);
nor U781 (N_781,N_734,N_566);
xor U782 (N_782,N_637,N_607);
and U783 (N_783,N_101,N_280);
xnor U784 (N_784,N_404,N_161);
nor U785 (N_785,N_335,N_10);
nand U786 (N_786,N_363,N_233);
or U787 (N_787,N_662,N_489);
and U788 (N_788,N_471,N_382);
nand U789 (N_789,N_630,N_676);
nor U790 (N_790,N_429,N_479);
or U791 (N_791,N_738,N_97);
nor U792 (N_792,N_431,N_449);
nand U793 (N_793,N_613,N_289);
nand U794 (N_794,N_273,N_106);
and U795 (N_795,N_443,N_344);
and U796 (N_796,N_2,N_693);
nor U797 (N_797,N_271,N_151);
nand U798 (N_798,N_452,N_340);
and U799 (N_799,N_82,N_583);
nor U800 (N_800,N_60,N_407);
or U801 (N_801,N_587,N_137);
nand U802 (N_802,N_604,N_26);
and U803 (N_803,N_509,N_679);
or U804 (N_804,N_104,N_598);
or U805 (N_805,N_490,N_400);
and U806 (N_806,N_269,N_716);
nand U807 (N_807,N_217,N_574);
nor U808 (N_808,N_384,N_469);
nand U809 (N_809,N_76,N_534);
nor U810 (N_810,N_124,N_308);
nor U811 (N_811,N_409,N_740);
nand U812 (N_812,N_183,N_385);
nor U813 (N_813,N_9,N_47);
and U814 (N_814,N_685,N_589);
nor U815 (N_815,N_648,N_731);
nand U816 (N_816,N_585,N_309);
nand U817 (N_817,N_401,N_665);
or U818 (N_818,N_748,N_41);
nand U819 (N_819,N_572,N_736);
nor U820 (N_820,N_168,N_533);
and U821 (N_821,N_180,N_427);
nor U822 (N_822,N_651,N_116);
nor U823 (N_823,N_262,N_307);
or U824 (N_824,N_159,N_654);
or U825 (N_825,N_261,N_515);
and U826 (N_826,N_163,N_355);
nor U827 (N_827,N_200,N_69);
or U828 (N_828,N_189,N_279);
nand U829 (N_829,N_712,N_84);
nand U830 (N_830,N_494,N_156);
nor U831 (N_831,N_442,N_121);
and U832 (N_832,N_455,N_678);
and U833 (N_833,N_27,N_242);
and U834 (N_834,N_146,N_173);
or U835 (N_835,N_222,N_257);
nor U836 (N_836,N_339,N_564);
nor U837 (N_837,N_424,N_380);
nor U838 (N_838,N_191,N_234);
nor U839 (N_839,N_324,N_499);
xor U840 (N_840,N_93,N_747);
or U841 (N_841,N_230,N_43);
nor U842 (N_842,N_235,N_256);
nor U843 (N_843,N_461,N_11);
and U844 (N_844,N_59,N_488);
and U845 (N_845,N_559,N_347);
or U846 (N_846,N_735,N_518);
and U847 (N_847,N_627,N_387);
and U848 (N_848,N_330,N_258);
and U849 (N_849,N_226,N_130);
or U850 (N_850,N_644,N_203);
and U851 (N_851,N_40,N_615);
nor U852 (N_852,N_171,N_742);
nand U853 (N_853,N_167,N_81);
and U854 (N_854,N_35,N_334);
nand U855 (N_855,N_579,N_208);
or U856 (N_856,N_193,N_558);
or U857 (N_857,N_366,N_95);
or U858 (N_858,N_336,N_502);
nand U859 (N_859,N_592,N_487);
or U860 (N_860,N_465,N_100);
or U861 (N_861,N_552,N_96);
nor U862 (N_862,N_90,N_724);
nand U863 (N_863,N_28,N_299);
nand U864 (N_864,N_51,N_632);
nor U865 (N_865,N_373,N_410);
and U866 (N_866,N_148,N_364);
and U867 (N_867,N_266,N_531);
and U868 (N_868,N_212,N_543);
and U869 (N_869,N_67,N_378);
nor U870 (N_870,N_204,N_128);
nand U871 (N_871,N_78,N_320);
nand U872 (N_872,N_147,N_105);
nor U873 (N_873,N_352,N_99);
or U874 (N_874,N_408,N_38);
nand U875 (N_875,N_686,N_567);
or U876 (N_876,N_162,N_232);
and U877 (N_877,N_671,N_165);
or U878 (N_878,N_45,N_444);
and U879 (N_879,N_746,N_687);
nand U880 (N_880,N_118,N_251);
nor U881 (N_881,N_597,N_492);
or U882 (N_882,N_525,N_12);
or U883 (N_883,N_649,N_125);
nor U884 (N_884,N_129,N_236);
nand U885 (N_885,N_64,N_594);
or U886 (N_886,N_31,N_275);
nor U887 (N_887,N_536,N_246);
nand U888 (N_888,N_126,N_88);
nor U889 (N_889,N_522,N_94);
nor U890 (N_890,N_628,N_143);
nor U891 (N_891,N_565,N_482);
nand U892 (N_892,N_79,N_523);
or U893 (N_893,N_227,N_353);
nor U894 (N_894,N_402,N_416);
and U895 (N_895,N_29,N_610);
or U896 (N_896,N_321,N_396);
nand U897 (N_897,N_220,N_729);
nand U898 (N_898,N_57,N_511);
or U899 (N_899,N_638,N_521);
nor U900 (N_900,N_317,N_300);
xor U901 (N_901,N_697,N_690);
nand U902 (N_902,N_605,N_643);
and U903 (N_903,N_288,N_292);
or U904 (N_904,N_207,N_535);
nand U905 (N_905,N_58,N_4);
and U906 (N_906,N_413,N_294);
nor U907 (N_907,N_358,N_13);
nor U908 (N_908,N_322,N_392);
nor U909 (N_909,N_153,N_0);
and U910 (N_910,N_655,N_377);
nor U911 (N_911,N_428,N_500);
nand U912 (N_912,N_721,N_30);
and U913 (N_913,N_606,N_403);
nand U914 (N_914,N_164,N_357);
and U915 (N_915,N_145,N_350);
nand U916 (N_916,N_17,N_477);
nand U917 (N_917,N_393,N_713);
nand U918 (N_918,N_98,N_225);
and U919 (N_919,N_278,N_692);
or U920 (N_920,N_91,N_584);
nand U921 (N_921,N_216,N_504);
nand U922 (N_922,N_512,N_318);
nand U923 (N_923,N_312,N_365);
nor U924 (N_924,N_142,N_135);
or U925 (N_925,N_458,N_18);
nand U926 (N_926,N_653,N_701);
or U927 (N_927,N_285,N_22);
xnor U928 (N_928,N_451,N_723);
nor U929 (N_929,N_626,N_672);
nand U930 (N_930,N_132,N_20);
nor U931 (N_931,N_42,N_141);
nor U932 (N_932,N_219,N_343);
nor U933 (N_933,N_629,N_120);
nand U934 (N_934,N_441,N_484);
nor U935 (N_935,N_507,N_381);
and U936 (N_936,N_25,N_707);
and U937 (N_937,N_5,N_647);
and U938 (N_938,N_157,N_631);
xor U939 (N_939,N_741,N_674);
nor U940 (N_940,N_291,N_37);
nand U941 (N_941,N_578,N_503);
and U942 (N_942,N_608,N_652);
nand U943 (N_943,N_14,N_744);
or U944 (N_944,N_136,N_250);
nand U945 (N_945,N_658,N_249);
or U946 (N_946,N_557,N_311);
and U947 (N_947,N_526,N_140);
and U948 (N_948,N_32,N_44);
nand U949 (N_949,N_622,N_706);
nand U950 (N_950,N_726,N_474);
or U951 (N_951,N_306,N_349);
nor U952 (N_952,N_667,N_370);
and U953 (N_953,N_176,N_625);
nand U954 (N_954,N_150,N_337);
or U955 (N_955,N_398,N_575);
xor U956 (N_956,N_749,N_541);
nor U957 (N_957,N_720,N_415);
or U958 (N_958,N_77,N_181);
nand U959 (N_959,N_421,N_178);
or U960 (N_960,N_664,N_259);
and U961 (N_961,N_301,N_72);
nor U962 (N_962,N_450,N_314);
or U963 (N_963,N_109,N_389);
nor U964 (N_964,N_528,N_463);
nor U965 (N_965,N_195,N_553);
and U966 (N_966,N_562,N_681);
or U967 (N_967,N_417,N_411);
nor U968 (N_968,N_54,N_3);
nor U969 (N_969,N_102,N_379);
and U970 (N_970,N_623,N_113);
xnor U971 (N_971,N_71,N_582);
nor U972 (N_972,N_538,N_694);
and U973 (N_973,N_677,N_544);
and U974 (N_974,N_593,N_149);
nor U975 (N_975,N_476,N_80);
nor U976 (N_976,N_34,N_172);
nor U977 (N_977,N_570,N_437);
nand U978 (N_978,N_702,N_532);
nand U979 (N_979,N_70,N_708);
nor U980 (N_980,N_1,N_272);
or U981 (N_981,N_399,N_619);
nand U982 (N_982,N_639,N_420);
and U983 (N_983,N_730,N_633);
and U984 (N_984,N_53,N_545);
or U985 (N_985,N_303,N_201);
or U986 (N_986,N_23,N_295);
or U987 (N_987,N_669,N_590);
nand U988 (N_988,N_739,N_154);
nor U989 (N_989,N_560,N_550);
nand U990 (N_990,N_86,N_620);
nor U991 (N_991,N_563,N_305);
nor U992 (N_992,N_663,N_122);
nor U993 (N_993,N_298,N_85);
and U994 (N_994,N_56,N_166);
nand U995 (N_995,N_733,N_656);
and U996 (N_996,N_395,N_467);
or U997 (N_997,N_313,N_673);
nand U998 (N_998,N_430,N_646);
nor U999 (N_999,N_268,N_635);
nor U1000 (N_1000,N_276,N_152);
xor U1001 (N_1001,N_63,N_284);
nand U1002 (N_1002,N_290,N_155);
or U1003 (N_1003,N_645,N_223);
or U1004 (N_1004,N_331,N_659);
and U1005 (N_1005,N_475,N_134);
nand U1006 (N_1006,N_325,N_698);
nor U1007 (N_1007,N_433,N_241);
or U1008 (N_1008,N_577,N_237);
or U1009 (N_1009,N_260,N_508);
nand U1010 (N_1010,N_718,N_425);
or U1011 (N_1011,N_107,N_372);
and U1012 (N_1012,N_177,N_253);
and U1013 (N_1013,N_556,N_354);
and U1014 (N_1014,N_383,N_516);
or U1015 (N_1015,N_714,N_517);
nand U1016 (N_1016,N_573,N_599);
xor U1017 (N_1017,N_368,N_498);
nor U1018 (N_1018,N_506,N_360);
nor U1019 (N_1019,N_440,N_213);
nor U1020 (N_1020,N_540,N_199);
or U1021 (N_1021,N_530,N_472);
or U1022 (N_1022,N_24,N_139);
and U1023 (N_1023,N_254,N_74);
nor U1024 (N_1024,N_537,N_561);
nand U1025 (N_1025,N_115,N_277);
nor U1026 (N_1026,N_496,N_8);
nand U1027 (N_1027,N_661,N_182);
xor U1028 (N_1028,N_524,N_478);
nand U1029 (N_1029,N_244,N_205);
nand U1030 (N_1030,N_239,N_689);
or U1031 (N_1031,N_581,N_493);
and U1032 (N_1032,N_700,N_650);
nor U1033 (N_1033,N_315,N_103);
nand U1034 (N_1034,N_660,N_388);
nand U1035 (N_1035,N_179,N_432);
or U1036 (N_1036,N_683,N_328);
nand U1037 (N_1037,N_423,N_580);
or U1038 (N_1038,N_252,N_68);
or U1039 (N_1039,N_187,N_287);
and U1040 (N_1040,N_636,N_722);
or U1041 (N_1041,N_243,N_481);
and U1042 (N_1042,N_709,N_348);
nor U1043 (N_1043,N_527,N_296);
and U1044 (N_1044,N_617,N_642);
nand U1045 (N_1045,N_510,N_319);
xor U1046 (N_1046,N_248,N_513);
nand U1047 (N_1047,N_209,N_293);
and U1048 (N_1048,N_62,N_55);
nand U1049 (N_1049,N_75,N_743);
and U1050 (N_1050,N_704,N_468);
and U1051 (N_1051,N_453,N_456);
or U1052 (N_1052,N_329,N_691);
or U1053 (N_1053,N_33,N_390);
nor U1054 (N_1054,N_274,N_666);
and U1055 (N_1055,N_131,N_133);
nor U1056 (N_1056,N_696,N_435);
nor U1057 (N_1057,N_112,N_341);
and U1058 (N_1058,N_264,N_459);
or U1059 (N_1059,N_682,N_640);
or U1060 (N_1060,N_514,N_188);
or U1061 (N_1061,N_46,N_231);
nor U1062 (N_1062,N_705,N_229);
or U1063 (N_1063,N_386,N_728);
nand U1064 (N_1064,N_202,N_323);
or U1065 (N_1065,N_36,N_611);
nor U1066 (N_1066,N_361,N_362);
and U1067 (N_1067,N_123,N_554);
and U1068 (N_1068,N_282,N_520);
and U1069 (N_1069,N_618,N_422);
nor U1070 (N_1070,N_405,N_548);
and U1071 (N_1071,N_356,N_447);
nor U1072 (N_1072,N_737,N_228);
and U1073 (N_1073,N_539,N_621);
xnor U1074 (N_1074,N_684,N_66);
nor U1075 (N_1075,N_265,N_87);
and U1076 (N_1076,N_210,N_65);
xor U1077 (N_1077,N_73,N_302);
nand U1078 (N_1078,N_169,N_699);
nor U1079 (N_1079,N_286,N_501);
and U1080 (N_1080,N_16,N_549);
nand U1081 (N_1081,N_7,N_371);
or U1082 (N_1082,N_591,N_418);
nor U1083 (N_1083,N_267,N_214);
nand U1084 (N_1084,N_192,N_327);
nand U1085 (N_1085,N_190,N_144);
and U1086 (N_1086,N_406,N_439);
nand U1087 (N_1087,N_448,N_119);
or U1088 (N_1088,N_247,N_376);
and U1089 (N_1089,N_184,N_680);
or U1090 (N_1090,N_255,N_316);
nor U1091 (N_1091,N_48,N_215);
and U1092 (N_1092,N_397,N_375);
nor U1093 (N_1093,N_454,N_391);
and U1094 (N_1094,N_52,N_670);
nor U1095 (N_1095,N_614,N_547);
nand U1096 (N_1096,N_92,N_332);
nor U1097 (N_1097,N_198,N_485);
nor U1098 (N_1098,N_283,N_568);
and U1099 (N_1099,N_281,N_310);
or U1100 (N_1100,N_446,N_345);
or U1101 (N_1101,N_466,N_486);
or U1102 (N_1102,N_464,N_657);
and U1103 (N_1103,N_719,N_529);
nand U1104 (N_1104,N_83,N_602);
and U1105 (N_1105,N_263,N_224);
or U1106 (N_1106,N_21,N_551);
or U1107 (N_1107,N_460,N_174);
nand U1108 (N_1108,N_127,N_436);
nor U1109 (N_1109,N_138,N_710);
or U1110 (N_1110,N_108,N_49);
nor U1111 (N_1111,N_462,N_394);
and U1112 (N_1112,N_675,N_218);
or U1113 (N_1113,N_703,N_603);
or U1114 (N_1114,N_338,N_438);
or U1115 (N_1115,N_110,N_624);
or U1116 (N_1116,N_304,N_270);
or U1117 (N_1117,N_588,N_571);
and U1118 (N_1118,N_297,N_15);
and U1119 (N_1119,N_596,N_186);
nand U1120 (N_1120,N_6,N_245);
nor U1121 (N_1121,N_240,N_346);
nor U1122 (N_1122,N_634,N_717);
or U1123 (N_1123,N_668,N_519);
nand U1124 (N_1124,N_457,N_196);
nand U1125 (N_1125,N_443,N_75);
or U1126 (N_1126,N_489,N_7);
or U1127 (N_1127,N_642,N_604);
and U1128 (N_1128,N_556,N_309);
and U1129 (N_1129,N_105,N_691);
or U1130 (N_1130,N_64,N_25);
nand U1131 (N_1131,N_250,N_337);
and U1132 (N_1132,N_290,N_696);
and U1133 (N_1133,N_611,N_396);
or U1134 (N_1134,N_529,N_332);
or U1135 (N_1135,N_633,N_483);
nor U1136 (N_1136,N_506,N_245);
nand U1137 (N_1137,N_73,N_37);
nor U1138 (N_1138,N_483,N_22);
or U1139 (N_1139,N_471,N_566);
nor U1140 (N_1140,N_633,N_212);
nor U1141 (N_1141,N_464,N_266);
nor U1142 (N_1142,N_586,N_493);
nor U1143 (N_1143,N_511,N_655);
nand U1144 (N_1144,N_476,N_260);
nor U1145 (N_1145,N_706,N_519);
or U1146 (N_1146,N_536,N_503);
or U1147 (N_1147,N_582,N_642);
and U1148 (N_1148,N_298,N_408);
nor U1149 (N_1149,N_84,N_231);
nand U1150 (N_1150,N_90,N_567);
and U1151 (N_1151,N_482,N_18);
and U1152 (N_1152,N_32,N_405);
nand U1153 (N_1153,N_18,N_501);
nand U1154 (N_1154,N_281,N_21);
or U1155 (N_1155,N_386,N_205);
nand U1156 (N_1156,N_424,N_402);
and U1157 (N_1157,N_167,N_270);
or U1158 (N_1158,N_519,N_505);
or U1159 (N_1159,N_170,N_607);
and U1160 (N_1160,N_463,N_348);
or U1161 (N_1161,N_371,N_639);
nor U1162 (N_1162,N_376,N_436);
or U1163 (N_1163,N_550,N_210);
nor U1164 (N_1164,N_458,N_11);
or U1165 (N_1165,N_276,N_561);
or U1166 (N_1166,N_66,N_346);
or U1167 (N_1167,N_673,N_732);
nand U1168 (N_1168,N_46,N_509);
or U1169 (N_1169,N_127,N_376);
or U1170 (N_1170,N_235,N_698);
and U1171 (N_1171,N_458,N_560);
nand U1172 (N_1172,N_313,N_407);
and U1173 (N_1173,N_556,N_685);
nor U1174 (N_1174,N_377,N_121);
nand U1175 (N_1175,N_380,N_370);
and U1176 (N_1176,N_274,N_366);
or U1177 (N_1177,N_138,N_521);
nor U1178 (N_1178,N_194,N_76);
nand U1179 (N_1179,N_268,N_38);
nand U1180 (N_1180,N_133,N_259);
nand U1181 (N_1181,N_316,N_438);
nor U1182 (N_1182,N_349,N_678);
and U1183 (N_1183,N_159,N_742);
nand U1184 (N_1184,N_344,N_169);
and U1185 (N_1185,N_612,N_374);
xnor U1186 (N_1186,N_83,N_297);
nand U1187 (N_1187,N_133,N_505);
or U1188 (N_1188,N_18,N_451);
and U1189 (N_1189,N_25,N_219);
nor U1190 (N_1190,N_47,N_35);
or U1191 (N_1191,N_457,N_218);
or U1192 (N_1192,N_279,N_483);
or U1193 (N_1193,N_140,N_527);
nand U1194 (N_1194,N_547,N_687);
or U1195 (N_1195,N_418,N_531);
or U1196 (N_1196,N_172,N_562);
xnor U1197 (N_1197,N_281,N_76);
nor U1198 (N_1198,N_446,N_748);
or U1199 (N_1199,N_589,N_740);
xnor U1200 (N_1200,N_585,N_215);
nor U1201 (N_1201,N_507,N_446);
and U1202 (N_1202,N_235,N_201);
xor U1203 (N_1203,N_604,N_410);
or U1204 (N_1204,N_159,N_240);
nor U1205 (N_1205,N_370,N_645);
and U1206 (N_1206,N_151,N_411);
nand U1207 (N_1207,N_527,N_206);
and U1208 (N_1208,N_453,N_346);
and U1209 (N_1209,N_176,N_116);
or U1210 (N_1210,N_76,N_536);
and U1211 (N_1211,N_501,N_526);
nand U1212 (N_1212,N_416,N_123);
or U1213 (N_1213,N_638,N_334);
and U1214 (N_1214,N_178,N_350);
nand U1215 (N_1215,N_185,N_560);
nand U1216 (N_1216,N_29,N_143);
and U1217 (N_1217,N_689,N_22);
or U1218 (N_1218,N_152,N_597);
nand U1219 (N_1219,N_369,N_110);
or U1220 (N_1220,N_136,N_365);
nor U1221 (N_1221,N_537,N_395);
nand U1222 (N_1222,N_688,N_9);
and U1223 (N_1223,N_40,N_505);
nand U1224 (N_1224,N_609,N_210);
nor U1225 (N_1225,N_154,N_372);
nand U1226 (N_1226,N_427,N_429);
nand U1227 (N_1227,N_199,N_283);
nor U1228 (N_1228,N_292,N_445);
or U1229 (N_1229,N_389,N_498);
xnor U1230 (N_1230,N_410,N_188);
or U1231 (N_1231,N_361,N_321);
nor U1232 (N_1232,N_697,N_429);
and U1233 (N_1233,N_41,N_500);
nor U1234 (N_1234,N_5,N_357);
nand U1235 (N_1235,N_252,N_639);
nor U1236 (N_1236,N_747,N_249);
xnor U1237 (N_1237,N_594,N_128);
nor U1238 (N_1238,N_157,N_74);
and U1239 (N_1239,N_226,N_582);
or U1240 (N_1240,N_296,N_129);
nand U1241 (N_1241,N_27,N_547);
nand U1242 (N_1242,N_558,N_742);
nor U1243 (N_1243,N_634,N_537);
and U1244 (N_1244,N_525,N_584);
nand U1245 (N_1245,N_551,N_30);
or U1246 (N_1246,N_306,N_415);
or U1247 (N_1247,N_197,N_99);
nand U1248 (N_1248,N_437,N_134);
nor U1249 (N_1249,N_180,N_303);
or U1250 (N_1250,N_17,N_363);
nand U1251 (N_1251,N_262,N_486);
nor U1252 (N_1252,N_715,N_112);
nand U1253 (N_1253,N_541,N_246);
or U1254 (N_1254,N_13,N_520);
or U1255 (N_1255,N_272,N_404);
nor U1256 (N_1256,N_263,N_19);
nor U1257 (N_1257,N_470,N_314);
nor U1258 (N_1258,N_8,N_384);
nand U1259 (N_1259,N_584,N_118);
nand U1260 (N_1260,N_202,N_442);
nand U1261 (N_1261,N_93,N_316);
nor U1262 (N_1262,N_747,N_333);
nor U1263 (N_1263,N_86,N_387);
or U1264 (N_1264,N_114,N_634);
or U1265 (N_1265,N_399,N_735);
and U1266 (N_1266,N_612,N_133);
and U1267 (N_1267,N_485,N_651);
nand U1268 (N_1268,N_584,N_635);
or U1269 (N_1269,N_685,N_645);
or U1270 (N_1270,N_576,N_630);
nor U1271 (N_1271,N_306,N_414);
and U1272 (N_1272,N_576,N_395);
nor U1273 (N_1273,N_239,N_536);
and U1274 (N_1274,N_607,N_734);
nor U1275 (N_1275,N_318,N_31);
or U1276 (N_1276,N_54,N_327);
nand U1277 (N_1277,N_228,N_659);
nor U1278 (N_1278,N_507,N_485);
nor U1279 (N_1279,N_465,N_193);
nor U1280 (N_1280,N_252,N_549);
xor U1281 (N_1281,N_470,N_143);
nor U1282 (N_1282,N_210,N_541);
or U1283 (N_1283,N_686,N_201);
nand U1284 (N_1284,N_564,N_106);
nand U1285 (N_1285,N_559,N_420);
nor U1286 (N_1286,N_685,N_729);
nor U1287 (N_1287,N_488,N_435);
nand U1288 (N_1288,N_712,N_609);
nand U1289 (N_1289,N_156,N_746);
nand U1290 (N_1290,N_317,N_485);
nand U1291 (N_1291,N_550,N_238);
nand U1292 (N_1292,N_375,N_4);
and U1293 (N_1293,N_96,N_437);
nor U1294 (N_1294,N_475,N_440);
nor U1295 (N_1295,N_502,N_297);
and U1296 (N_1296,N_289,N_216);
or U1297 (N_1297,N_597,N_510);
nand U1298 (N_1298,N_541,N_506);
nor U1299 (N_1299,N_709,N_514);
nand U1300 (N_1300,N_645,N_398);
nor U1301 (N_1301,N_540,N_455);
nand U1302 (N_1302,N_677,N_178);
and U1303 (N_1303,N_536,N_727);
and U1304 (N_1304,N_271,N_723);
or U1305 (N_1305,N_422,N_608);
and U1306 (N_1306,N_308,N_508);
nand U1307 (N_1307,N_54,N_655);
and U1308 (N_1308,N_314,N_363);
nor U1309 (N_1309,N_167,N_485);
and U1310 (N_1310,N_447,N_154);
or U1311 (N_1311,N_536,N_381);
and U1312 (N_1312,N_140,N_270);
nor U1313 (N_1313,N_253,N_516);
nor U1314 (N_1314,N_512,N_361);
nor U1315 (N_1315,N_463,N_605);
or U1316 (N_1316,N_230,N_720);
or U1317 (N_1317,N_596,N_71);
nand U1318 (N_1318,N_359,N_409);
or U1319 (N_1319,N_32,N_413);
and U1320 (N_1320,N_454,N_636);
nor U1321 (N_1321,N_681,N_120);
or U1322 (N_1322,N_519,N_538);
nand U1323 (N_1323,N_549,N_709);
nor U1324 (N_1324,N_65,N_336);
nand U1325 (N_1325,N_748,N_688);
and U1326 (N_1326,N_63,N_628);
nand U1327 (N_1327,N_28,N_82);
nor U1328 (N_1328,N_238,N_258);
nor U1329 (N_1329,N_590,N_369);
nand U1330 (N_1330,N_106,N_312);
or U1331 (N_1331,N_666,N_47);
nor U1332 (N_1332,N_70,N_3);
or U1333 (N_1333,N_29,N_471);
or U1334 (N_1334,N_163,N_427);
nor U1335 (N_1335,N_229,N_564);
and U1336 (N_1336,N_583,N_12);
or U1337 (N_1337,N_190,N_447);
and U1338 (N_1338,N_530,N_491);
nor U1339 (N_1339,N_631,N_535);
xor U1340 (N_1340,N_512,N_138);
nand U1341 (N_1341,N_232,N_618);
nand U1342 (N_1342,N_109,N_256);
or U1343 (N_1343,N_160,N_346);
or U1344 (N_1344,N_24,N_462);
nand U1345 (N_1345,N_301,N_209);
nor U1346 (N_1346,N_354,N_145);
nand U1347 (N_1347,N_508,N_352);
and U1348 (N_1348,N_353,N_168);
and U1349 (N_1349,N_447,N_88);
and U1350 (N_1350,N_186,N_615);
or U1351 (N_1351,N_490,N_439);
and U1352 (N_1352,N_342,N_66);
nor U1353 (N_1353,N_123,N_380);
nand U1354 (N_1354,N_167,N_654);
nand U1355 (N_1355,N_81,N_176);
and U1356 (N_1356,N_627,N_733);
xnor U1357 (N_1357,N_510,N_256);
nand U1358 (N_1358,N_197,N_484);
nor U1359 (N_1359,N_625,N_470);
and U1360 (N_1360,N_134,N_586);
or U1361 (N_1361,N_275,N_66);
and U1362 (N_1362,N_289,N_267);
nand U1363 (N_1363,N_670,N_333);
or U1364 (N_1364,N_104,N_274);
nand U1365 (N_1365,N_422,N_97);
nor U1366 (N_1366,N_396,N_506);
nor U1367 (N_1367,N_177,N_621);
or U1368 (N_1368,N_286,N_255);
or U1369 (N_1369,N_425,N_78);
and U1370 (N_1370,N_450,N_517);
nor U1371 (N_1371,N_715,N_96);
and U1372 (N_1372,N_9,N_605);
nor U1373 (N_1373,N_124,N_311);
or U1374 (N_1374,N_370,N_324);
nand U1375 (N_1375,N_539,N_675);
nor U1376 (N_1376,N_362,N_76);
nand U1377 (N_1377,N_342,N_97);
and U1378 (N_1378,N_347,N_402);
and U1379 (N_1379,N_554,N_715);
or U1380 (N_1380,N_551,N_618);
or U1381 (N_1381,N_665,N_162);
or U1382 (N_1382,N_70,N_428);
nor U1383 (N_1383,N_599,N_741);
and U1384 (N_1384,N_271,N_555);
or U1385 (N_1385,N_50,N_17);
nand U1386 (N_1386,N_581,N_659);
and U1387 (N_1387,N_87,N_445);
nand U1388 (N_1388,N_313,N_294);
nor U1389 (N_1389,N_631,N_441);
nor U1390 (N_1390,N_520,N_485);
nand U1391 (N_1391,N_297,N_41);
nor U1392 (N_1392,N_667,N_325);
nand U1393 (N_1393,N_365,N_729);
nor U1394 (N_1394,N_302,N_125);
nor U1395 (N_1395,N_547,N_101);
nor U1396 (N_1396,N_305,N_435);
and U1397 (N_1397,N_582,N_155);
nand U1398 (N_1398,N_21,N_122);
nand U1399 (N_1399,N_189,N_664);
nor U1400 (N_1400,N_474,N_543);
or U1401 (N_1401,N_327,N_8);
and U1402 (N_1402,N_609,N_452);
nor U1403 (N_1403,N_267,N_7);
nor U1404 (N_1404,N_380,N_701);
or U1405 (N_1405,N_515,N_68);
nor U1406 (N_1406,N_246,N_155);
and U1407 (N_1407,N_514,N_240);
and U1408 (N_1408,N_630,N_66);
xnor U1409 (N_1409,N_112,N_300);
nand U1410 (N_1410,N_11,N_514);
nor U1411 (N_1411,N_565,N_707);
nand U1412 (N_1412,N_586,N_514);
nand U1413 (N_1413,N_648,N_116);
nor U1414 (N_1414,N_103,N_316);
and U1415 (N_1415,N_395,N_99);
or U1416 (N_1416,N_540,N_575);
nor U1417 (N_1417,N_680,N_36);
or U1418 (N_1418,N_523,N_526);
and U1419 (N_1419,N_459,N_65);
and U1420 (N_1420,N_737,N_501);
nand U1421 (N_1421,N_409,N_646);
xnor U1422 (N_1422,N_205,N_231);
nor U1423 (N_1423,N_135,N_385);
or U1424 (N_1424,N_222,N_424);
nand U1425 (N_1425,N_15,N_96);
nor U1426 (N_1426,N_685,N_695);
and U1427 (N_1427,N_705,N_477);
or U1428 (N_1428,N_440,N_86);
or U1429 (N_1429,N_654,N_684);
and U1430 (N_1430,N_367,N_118);
nand U1431 (N_1431,N_166,N_217);
or U1432 (N_1432,N_400,N_621);
and U1433 (N_1433,N_682,N_333);
nor U1434 (N_1434,N_105,N_426);
xor U1435 (N_1435,N_437,N_728);
nand U1436 (N_1436,N_14,N_379);
nor U1437 (N_1437,N_34,N_659);
or U1438 (N_1438,N_641,N_166);
nor U1439 (N_1439,N_158,N_375);
nor U1440 (N_1440,N_195,N_683);
and U1441 (N_1441,N_11,N_84);
nor U1442 (N_1442,N_75,N_105);
nor U1443 (N_1443,N_303,N_456);
or U1444 (N_1444,N_637,N_162);
or U1445 (N_1445,N_29,N_114);
or U1446 (N_1446,N_143,N_158);
nor U1447 (N_1447,N_654,N_630);
or U1448 (N_1448,N_608,N_63);
or U1449 (N_1449,N_434,N_56);
and U1450 (N_1450,N_411,N_81);
and U1451 (N_1451,N_255,N_645);
nand U1452 (N_1452,N_529,N_139);
nand U1453 (N_1453,N_381,N_496);
and U1454 (N_1454,N_612,N_499);
or U1455 (N_1455,N_616,N_562);
and U1456 (N_1456,N_346,N_250);
xor U1457 (N_1457,N_345,N_306);
or U1458 (N_1458,N_637,N_719);
or U1459 (N_1459,N_428,N_287);
nand U1460 (N_1460,N_136,N_584);
nand U1461 (N_1461,N_14,N_554);
and U1462 (N_1462,N_330,N_371);
nor U1463 (N_1463,N_153,N_575);
nor U1464 (N_1464,N_465,N_604);
nand U1465 (N_1465,N_626,N_311);
nor U1466 (N_1466,N_370,N_541);
nor U1467 (N_1467,N_659,N_141);
nand U1468 (N_1468,N_540,N_687);
nor U1469 (N_1469,N_50,N_250);
nor U1470 (N_1470,N_673,N_360);
xnor U1471 (N_1471,N_405,N_547);
nand U1472 (N_1472,N_70,N_133);
nor U1473 (N_1473,N_361,N_463);
or U1474 (N_1474,N_188,N_606);
nor U1475 (N_1475,N_350,N_160);
nor U1476 (N_1476,N_451,N_356);
or U1477 (N_1477,N_82,N_382);
nand U1478 (N_1478,N_266,N_307);
nand U1479 (N_1479,N_108,N_635);
nand U1480 (N_1480,N_313,N_466);
and U1481 (N_1481,N_278,N_353);
nand U1482 (N_1482,N_629,N_201);
or U1483 (N_1483,N_98,N_652);
nand U1484 (N_1484,N_387,N_426);
nand U1485 (N_1485,N_84,N_718);
nand U1486 (N_1486,N_729,N_322);
and U1487 (N_1487,N_746,N_650);
and U1488 (N_1488,N_585,N_14);
nor U1489 (N_1489,N_164,N_598);
nor U1490 (N_1490,N_188,N_713);
nor U1491 (N_1491,N_348,N_189);
and U1492 (N_1492,N_270,N_467);
nand U1493 (N_1493,N_186,N_228);
and U1494 (N_1494,N_584,N_213);
nor U1495 (N_1495,N_158,N_269);
or U1496 (N_1496,N_691,N_508);
and U1497 (N_1497,N_368,N_314);
xnor U1498 (N_1498,N_429,N_238);
and U1499 (N_1499,N_128,N_259);
nand U1500 (N_1500,N_1318,N_1175);
and U1501 (N_1501,N_1430,N_847);
nor U1502 (N_1502,N_1121,N_1324);
and U1503 (N_1503,N_902,N_1282);
nor U1504 (N_1504,N_1106,N_898);
nor U1505 (N_1505,N_1073,N_1322);
nand U1506 (N_1506,N_766,N_1115);
nor U1507 (N_1507,N_939,N_1114);
nor U1508 (N_1508,N_1268,N_1427);
nand U1509 (N_1509,N_1257,N_997);
or U1510 (N_1510,N_1197,N_1043);
and U1511 (N_1511,N_1474,N_1097);
or U1512 (N_1512,N_968,N_1364);
and U1513 (N_1513,N_1065,N_1450);
or U1514 (N_1514,N_1206,N_1440);
nand U1515 (N_1515,N_770,N_909);
and U1516 (N_1516,N_1074,N_1300);
or U1517 (N_1517,N_1353,N_768);
or U1518 (N_1518,N_1159,N_1231);
nor U1519 (N_1519,N_1358,N_1188);
nor U1520 (N_1520,N_1029,N_925);
or U1521 (N_1521,N_1341,N_1251);
nor U1522 (N_1522,N_1140,N_1241);
nand U1523 (N_1523,N_781,N_981);
nand U1524 (N_1524,N_1262,N_944);
nand U1525 (N_1525,N_1299,N_1357);
nand U1526 (N_1526,N_1185,N_1352);
nor U1527 (N_1527,N_1199,N_1298);
and U1528 (N_1528,N_1165,N_963);
nor U1529 (N_1529,N_955,N_880);
nand U1530 (N_1530,N_1220,N_1442);
nor U1531 (N_1531,N_971,N_836);
or U1532 (N_1532,N_1174,N_1327);
and U1533 (N_1533,N_1328,N_864);
nor U1534 (N_1534,N_884,N_800);
and U1535 (N_1535,N_1494,N_1448);
nand U1536 (N_1536,N_1201,N_1177);
and U1537 (N_1537,N_848,N_1258);
or U1538 (N_1538,N_760,N_793);
nand U1539 (N_1539,N_761,N_1454);
nand U1540 (N_1540,N_1014,N_1006);
xor U1541 (N_1541,N_1271,N_1195);
nor U1542 (N_1542,N_775,N_1018);
nor U1543 (N_1543,N_1412,N_811);
nand U1544 (N_1544,N_1356,N_1212);
or U1545 (N_1545,N_1335,N_1062);
nand U1546 (N_1546,N_855,N_1064);
or U1547 (N_1547,N_1105,N_1210);
and U1548 (N_1548,N_1055,N_1048);
or U1549 (N_1549,N_1343,N_1375);
nor U1550 (N_1550,N_1093,N_846);
xnor U1551 (N_1551,N_818,N_1112);
nor U1552 (N_1552,N_1110,N_1484);
or U1553 (N_1553,N_1287,N_961);
and U1554 (N_1554,N_1173,N_1270);
and U1555 (N_1555,N_930,N_1422);
nor U1556 (N_1556,N_1168,N_1263);
and U1557 (N_1557,N_949,N_755);
or U1558 (N_1558,N_980,N_1451);
nand U1559 (N_1559,N_1303,N_1053);
nand U1560 (N_1560,N_1242,N_1128);
nand U1561 (N_1561,N_1002,N_1397);
nor U1562 (N_1562,N_1143,N_1475);
nand U1563 (N_1563,N_1331,N_1005);
nor U1564 (N_1564,N_1481,N_1330);
nand U1565 (N_1565,N_1379,N_1304);
nor U1566 (N_1566,N_1314,N_1041);
nor U1567 (N_1567,N_825,N_929);
or U1568 (N_1568,N_1090,N_1100);
and U1569 (N_1569,N_1408,N_1340);
nor U1570 (N_1570,N_1488,N_1189);
nand U1571 (N_1571,N_807,N_853);
nand U1572 (N_1572,N_1499,N_1286);
nand U1573 (N_1573,N_844,N_1207);
and U1574 (N_1574,N_1489,N_1040);
and U1575 (N_1575,N_915,N_1365);
or U1576 (N_1576,N_1030,N_897);
nor U1577 (N_1577,N_1204,N_1019);
nor U1578 (N_1578,N_865,N_1301);
nor U1579 (N_1579,N_1089,N_868);
or U1580 (N_1580,N_1393,N_1349);
nor U1581 (N_1581,N_1186,N_923);
xnor U1582 (N_1582,N_1034,N_808);
and U1583 (N_1583,N_866,N_769);
nand U1584 (N_1584,N_1493,N_838);
and U1585 (N_1585,N_1361,N_1081);
nor U1586 (N_1586,N_1443,N_788);
and U1587 (N_1587,N_860,N_1439);
nor U1588 (N_1588,N_916,N_1176);
or U1589 (N_1589,N_1059,N_1249);
or U1590 (N_1590,N_1339,N_794);
nor U1591 (N_1591,N_859,N_1142);
nand U1592 (N_1592,N_1109,N_888);
nor U1593 (N_1593,N_863,N_1329);
nor U1594 (N_1594,N_988,N_1264);
or U1595 (N_1595,N_1198,N_840);
or U1596 (N_1596,N_1461,N_1052);
and U1597 (N_1597,N_911,N_891);
nor U1598 (N_1598,N_1426,N_1056);
nor U1599 (N_1599,N_751,N_1103);
nor U1600 (N_1600,N_1369,N_1203);
nand U1601 (N_1601,N_1194,N_1421);
nor U1602 (N_1602,N_764,N_1205);
nand U1603 (N_1603,N_1462,N_1482);
or U1604 (N_1604,N_1266,N_1285);
nor U1605 (N_1605,N_1079,N_1162);
xnor U1606 (N_1606,N_1163,N_977);
or U1607 (N_1607,N_852,N_1191);
nor U1608 (N_1608,N_1274,N_932);
and U1609 (N_1609,N_1158,N_1181);
and U1610 (N_1610,N_1148,N_917);
and U1611 (N_1611,N_871,N_1178);
nand U1612 (N_1612,N_1269,N_990);
or U1613 (N_1613,N_1374,N_1061);
and U1614 (N_1614,N_934,N_1278);
or U1615 (N_1615,N_805,N_1072);
xnor U1616 (N_1616,N_833,N_1476);
or U1617 (N_1617,N_966,N_1399);
and U1618 (N_1618,N_970,N_1350);
nand U1619 (N_1619,N_1498,N_908);
nor U1620 (N_1620,N_850,N_1347);
nor U1621 (N_1621,N_1313,N_1233);
nand U1622 (N_1622,N_1311,N_992);
and U1623 (N_1623,N_1388,N_822);
nor U1624 (N_1624,N_1133,N_754);
nor U1625 (N_1625,N_842,N_1135);
nand U1626 (N_1626,N_841,N_1292);
nor U1627 (N_1627,N_1398,N_1360);
nand U1628 (N_1628,N_1382,N_1326);
and U1629 (N_1629,N_1230,N_1316);
and U1630 (N_1630,N_1453,N_1101);
nand U1631 (N_1631,N_1216,N_1245);
nand U1632 (N_1632,N_1338,N_1265);
xor U1633 (N_1633,N_1141,N_1460);
nand U1634 (N_1634,N_1359,N_1192);
or U1635 (N_1635,N_802,N_1363);
nor U1636 (N_1636,N_1348,N_1290);
or U1637 (N_1637,N_757,N_1256);
nor U1638 (N_1638,N_1319,N_1446);
or U1639 (N_1639,N_940,N_835);
or U1640 (N_1640,N_1490,N_1063);
and U1641 (N_1641,N_1208,N_1108);
nor U1642 (N_1642,N_830,N_1456);
nor U1643 (N_1643,N_782,N_994);
or U1644 (N_1644,N_1323,N_1305);
nand U1645 (N_1645,N_1077,N_879);
nand U1646 (N_1646,N_1126,N_964);
nand U1647 (N_1647,N_1116,N_1373);
or U1648 (N_1648,N_784,N_1229);
or U1649 (N_1649,N_1336,N_1050);
xor U1650 (N_1650,N_858,N_1325);
and U1651 (N_1651,N_1254,N_1289);
or U1652 (N_1652,N_1459,N_1051);
nand U1653 (N_1653,N_1409,N_806);
nand U1654 (N_1654,N_1084,N_1202);
nand U1655 (N_1655,N_1119,N_869);
nand U1656 (N_1656,N_1211,N_792);
and U1657 (N_1657,N_1279,N_1312);
nor U1658 (N_1658,N_1008,N_943);
and U1659 (N_1659,N_753,N_1144);
nor U1660 (N_1660,N_780,N_1013);
and U1661 (N_1661,N_1009,N_1280);
or U1662 (N_1662,N_881,N_877);
and U1663 (N_1663,N_1416,N_1130);
or U1664 (N_1664,N_1071,N_998);
nand U1665 (N_1665,N_1468,N_1376);
or U1666 (N_1666,N_803,N_1415);
nand U1667 (N_1667,N_1237,N_1337);
and U1668 (N_1668,N_1297,N_1020);
or U1669 (N_1669,N_893,N_1463);
nand U1670 (N_1670,N_845,N_1293);
nand U1671 (N_1671,N_1215,N_1378);
or U1672 (N_1672,N_1392,N_867);
nand U1673 (N_1673,N_756,N_758);
nor U1674 (N_1674,N_1272,N_1099);
or U1675 (N_1675,N_941,N_959);
nand U1676 (N_1676,N_1066,N_791);
nand U1677 (N_1677,N_1473,N_957);
and U1678 (N_1678,N_1445,N_1139);
and U1679 (N_1679,N_851,N_1486);
nor U1680 (N_1680,N_1492,N_1037);
and U1681 (N_1681,N_1068,N_989);
nand U1682 (N_1682,N_889,N_1044);
and U1683 (N_1683,N_839,N_759);
nor U1684 (N_1684,N_829,N_1138);
and U1685 (N_1685,N_827,N_899);
nand U1686 (N_1686,N_1088,N_797);
nand U1687 (N_1687,N_1153,N_1118);
or U1688 (N_1688,N_1320,N_920);
nand U1689 (N_1689,N_1067,N_1223);
nand U1690 (N_1690,N_1224,N_1228);
nand U1691 (N_1691,N_1385,N_798);
and U1692 (N_1692,N_922,N_783);
and U1693 (N_1693,N_1120,N_813);
nand U1694 (N_1694,N_1413,N_1469);
nor U1695 (N_1695,N_1342,N_1394);
or U1696 (N_1696,N_1387,N_857);
xnor U1697 (N_1697,N_772,N_1383);
nor U1698 (N_1698,N_804,N_826);
or U1699 (N_1699,N_1260,N_849);
or U1700 (N_1700,N_1437,N_823);
and U1701 (N_1701,N_876,N_1017);
nand U1702 (N_1702,N_1267,N_1087);
and U1703 (N_1703,N_837,N_1396);
nand U1704 (N_1704,N_862,N_935);
or U1705 (N_1705,N_778,N_1196);
or U1706 (N_1706,N_1367,N_1407);
xnor U1707 (N_1707,N_1244,N_1283);
or U1708 (N_1708,N_907,N_921);
nor U1709 (N_1709,N_1479,N_809);
or U1710 (N_1710,N_928,N_812);
and U1711 (N_1711,N_1240,N_1395);
nand U1712 (N_1712,N_962,N_1154);
nor U1713 (N_1713,N_1465,N_1418);
nor U1714 (N_1714,N_926,N_870);
or U1715 (N_1715,N_1021,N_1447);
nand U1716 (N_1716,N_1161,N_1302);
nor U1717 (N_1717,N_1047,N_1334);
nand U1718 (N_1718,N_901,N_1368);
or U1719 (N_1719,N_1317,N_1478);
nor U1720 (N_1720,N_1321,N_976);
and U1721 (N_1721,N_904,N_1222);
xnor U1722 (N_1722,N_1083,N_1184);
and U1723 (N_1723,N_1410,N_885);
nor U1724 (N_1724,N_982,N_1057);
and U1725 (N_1725,N_1149,N_1243);
nand U1726 (N_1726,N_1281,N_875);
nand U1727 (N_1727,N_1076,N_931);
or U1728 (N_1728,N_1370,N_1255);
nor U1729 (N_1729,N_767,N_1225);
and U1730 (N_1730,N_1273,N_1424);
nand U1731 (N_1731,N_882,N_1042);
xor U1732 (N_1732,N_906,N_1308);
nand U1733 (N_1733,N_1190,N_1155);
nand U1734 (N_1734,N_969,N_1169);
nand U1735 (N_1735,N_1086,N_1487);
nand U1736 (N_1736,N_912,N_1036);
nand U1737 (N_1737,N_1362,N_1069);
and U1738 (N_1738,N_820,N_1092);
or U1739 (N_1739,N_945,N_886);
nand U1740 (N_1740,N_938,N_771);
nand U1741 (N_1741,N_1193,N_1449);
and U1742 (N_1742,N_1252,N_965);
and U1743 (N_1743,N_1007,N_960);
xor U1744 (N_1744,N_953,N_834);
or U1745 (N_1745,N_1085,N_1035);
and U1746 (N_1746,N_786,N_1150);
or U1747 (N_1747,N_1124,N_1354);
and U1748 (N_1748,N_1384,N_1123);
nor U1749 (N_1749,N_1049,N_1038);
or U1750 (N_1750,N_1032,N_883);
nand U1751 (N_1751,N_856,N_1423);
nand U1752 (N_1752,N_1261,N_1315);
nor U1753 (N_1753,N_1111,N_1132);
and U1754 (N_1754,N_1003,N_1136);
nand U1755 (N_1755,N_1275,N_789);
nor U1756 (N_1756,N_1452,N_1200);
nor U1757 (N_1757,N_903,N_1219);
or U1758 (N_1758,N_1179,N_1152);
nand U1759 (N_1759,N_950,N_1010);
nor U1760 (N_1760,N_763,N_1167);
nand U1761 (N_1761,N_790,N_1247);
nor U1762 (N_1762,N_1250,N_918);
nor U1763 (N_1763,N_843,N_1259);
and U1764 (N_1764,N_817,N_1344);
and U1765 (N_1765,N_1022,N_1027);
nor U1766 (N_1766,N_1355,N_937);
nor U1767 (N_1767,N_1226,N_832);
xor U1768 (N_1768,N_913,N_890);
and U1769 (N_1769,N_1406,N_1058);
and U1770 (N_1770,N_1147,N_958);
or U1771 (N_1771,N_1480,N_1333);
nand U1772 (N_1772,N_1248,N_1496);
nor U1773 (N_1773,N_1172,N_896);
nand U1774 (N_1774,N_1171,N_821);
nor U1775 (N_1775,N_967,N_1217);
or U1776 (N_1776,N_1238,N_1221);
and U1777 (N_1777,N_1390,N_1471);
nand U1778 (N_1778,N_1346,N_1070);
nor U1779 (N_1779,N_1246,N_1411);
nor U1780 (N_1780,N_1428,N_995);
nor U1781 (N_1781,N_987,N_1026);
nand U1782 (N_1782,N_1157,N_1295);
or U1783 (N_1783,N_1082,N_974);
and U1784 (N_1784,N_1389,N_1386);
nor U1785 (N_1785,N_1284,N_774);
nor U1786 (N_1786,N_942,N_1011);
nor U1787 (N_1787,N_975,N_785);
and U1788 (N_1788,N_762,N_1405);
and U1789 (N_1789,N_1234,N_1094);
xor U1790 (N_1790,N_936,N_1458);
nor U1791 (N_1791,N_1483,N_1000);
and U1792 (N_1792,N_777,N_1080);
nand U1793 (N_1793,N_1146,N_1134);
nor U1794 (N_1794,N_1419,N_1232);
nand U1795 (N_1795,N_1276,N_927);
xnor U1796 (N_1796,N_1381,N_946);
or U1797 (N_1797,N_973,N_1425);
or U1798 (N_1798,N_1391,N_1431);
or U1799 (N_1799,N_1306,N_1031);
nand U1800 (N_1800,N_773,N_1156);
nor U1801 (N_1801,N_1277,N_854);
and U1802 (N_1802,N_983,N_1414);
nor U1803 (N_1803,N_991,N_1491);
and U1804 (N_1804,N_1060,N_819);
nor U1805 (N_1805,N_984,N_978);
nand U1806 (N_1806,N_952,N_986);
nor U1807 (N_1807,N_799,N_828);
nor U1808 (N_1808,N_993,N_1402);
nand U1809 (N_1809,N_1434,N_1025);
and U1810 (N_1810,N_895,N_1170);
and U1811 (N_1811,N_1429,N_1096);
nor U1812 (N_1812,N_1098,N_1296);
and U1813 (N_1813,N_1457,N_1001);
nor U1814 (N_1814,N_887,N_1127);
or U1815 (N_1815,N_1464,N_801);
and U1816 (N_1816,N_878,N_1166);
or U1817 (N_1817,N_1012,N_996);
nand U1818 (N_1818,N_1218,N_1023);
and U1819 (N_1819,N_1332,N_919);
or U1820 (N_1820,N_1209,N_1039);
or U1821 (N_1821,N_1444,N_1239);
xnor U1822 (N_1822,N_796,N_1294);
and U1823 (N_1823,N_1182,N_979);
xnor U1824 (N_1824,N_1436,N_1401);
nand U1825 (N_1825,N_1438,N_752);
and U1826 (N_1826,N_795,N_1472);
nor U1827 (N_1827,N_810,N_1016);
and U1828 (N_1828,N_1467,N_1420);
and U1829 (N_1829,N_815,N_1046);
and U1830 (N_1830,N_831,N_1131);
or U1831 (N_1831,N_905,N_1291);
nand U1832 (N_1832,N_750,N_1253);
and U1833 (N_1833,N_1433,N_1028);
or U1834 (N_1834,N_1227,N_873);
or U1835 (N_1835,N_1187,N_1078);
or U1836 (N_1836,N_999,N_1004);
nor U1837 (N_1837,N_900,N_1497);
nand U1838 (N_1838,N_776,N_1366);
nand U1839 (N_1839,N_1403,N_1470);
or U1840 (N_1840,N_1024,N_1307);
nor U1841 (N_1841,N_1091,N_1404);
or U1842 (N_1842,N_947,N_1372);
nand U1843 (N_1843,N_1435,N_1310);
nand U1844 (N_1844,N_1235,N_1380);
and U1845 (N_1845,N_1045,N_1183);
nor U1846 (N_1846,N_1129,N_910);
or U1847 (N_1847,N_1485,N_1345);
nand U1848 (N_1848,N_1400,N_872);
xnor U1849 (N_1849,N_1351,N_874);
xnor U1850 (N_1850,N_948,N_1214);
or U1851 (N_1851,N_1122,N_779);
and U1852 (N_1852,N_1377,N_1213);
nor U1853 (N_1853,N_1160,N_1477);
or U1854 (N_1854,N_1371,N_1015);
nor U1855 (N_1855,N_824,N_951);
nand U1856 (N_1856,N_1432,N_956);
nor U1857 (N_1857,N_1441,N_861);
or U1858 (N_1858,N_1095,N_954);
nand U1859 (N_1859,N_1102,N_1113);
nand U1860 (N_1860,N_816,N_1151);
nand U1861 (N_1861,N_933,N_1309);
and U1862 (N_1862,N_1137,N_985);
or U1863 (N_1863,N_1236,N_914);
nand U1864 (N_1864,N_1288,N_972);
nor U1865 (N_1865,N_1104,N_1455);
nand U1866 (N_1866,N_1125,N_787);
or U1867 (N_1867,N_1164,N_1180);
and U1868 (N_1868,N_892,N_1107);
and U1869 (N_1869,N_924,N_1075);
nor U1870 (N_1870,N_894,N_1417);
or U1871 (N_1871,N_1117,N_814);
nand U1872 (N_1872,N_765,N_1033);
xnor U1873 (N_1873,N_1466,N_1145);
and U1874 (N_1874,N_1495,N_1054);
or U1875 (N_1875,N_1280,N_863);
nand U1876 (N_1876,N_1357,N_1126);
nor U1877 (N_1877,N_1136,N_952);
and U1878 (N_1878,N_1047,N_1103);
nand U1879 (N_1879,N_830,N_1138);
and U1880 (N_1880,N_920,N_1401);
or U1881 (N_1881,N_852,N_1180);
and U1882 (N_1882,N_1085,N_1443);
and U1883 (N_1883,N_767,N_1326);
or U1884 (N_1884,N_1385,N_842);
nand U1885 (N_1885,N_1223,N_1304);
nand U1886 (N_1886,N_1312,N_1360);
or U1887 (N_1887,N_927,N_1357);
and U1888 (N_1888,N_1085,N_960);
nand U1889 (N_1889,N_1450,N_770);
nor U1890 (N_1890,N_1405,N_807);
nand U1891 (N_1891,N_1111,N_1059);
nor U1892 (N_1892,N_1267,N_921);
nor U1893 (N_1893,N_1064,N_864);
nor U1894 (N_1894,N_1015,N_881);
nor U1895 (N_1895,N_1472,N_902);
and U1896 (N_1896,N_995,N_921);
nand U1897 (N_1897,N_820,N_1238);
nand U1898 (N_1898,N_1138,N_750);
or U1899 (N_1899,N_838,N_1449);
xor U1900 (N_1900,N_1123,N_1291);
and U1901 (N_1901,N_1029,N_1439);
nor U1902 (N_1902,N_1497,N_1170);
or U1903 (N_1903,N_1465,N_1444);
nand U1904 (N_1904,N_1187,N_1476);
nand U1905 (N_1905,N_1293,N_834);
or U1906 (N_1906,N_903,N_1406);
and U1907 (N_1907,N_1034,N_1385);
and U1908 (N_1908,N_852,N_905);
and U1909 (N_1909,N_953,N_930);
and U1910 (N_1910,N_1053,N_918);
and U1911 (N_1911,N_780,N_817);
or U1912 (N_1912,N_931,N_1239);
nand U1913 (N_1913,N_1313,N_756);
or U1914 (N_1914,N_1366,N_1177);
nor U1915 (N_1915,N_1494,N_759);
nand U1916 (N_1916,N_1293,N_1092);
and U1917 (N_1917,N_1316,N_1237);
or U1918 (N_1918,N_786,N_1462);
or U1919 (N_1919,N_1191,N_854);
and U1920 (N_1920,N_945,N_872);
xnor U1921 (N_1921,N_1405,N_1083);
and U1922 (N_1922,N_1453,N_766);
and U1923 (N_1923,N_1381,N_894);
and U1924 (N_1924,N_1039,N_1273);
and U1925 (N_1925,N_1080,N_1434);
nand U1926 (N_1926,N_1227,N_1091);
nand U1927 (N_1927,N_1480,N_851);
and U1928 (N_1928,N_824,N_782);
or U1929 (N_1929,N_1037,N_1087);
nand U1930 (N_1930,N_1427,N_897);
nor U1931 (N_1931,N_1413,N_1176);
and U1932 (N_1932,N_1472,N_1135);
nand U1933 (N_1933,N_1267,N_913);
or U1934 (N_1934,N_909,N_1052);
and U1935 (N_1935,N_920,N_857);
and U1936 (N_1936,N_1134,N_1073);
nor U1937 (N_1937,N_872,N_1302);
and U1938 (N_1938,N_807,N_1225);
or U1939 (N_1939,N_1285,N_803);
or U1940 (N_1940,N_1472,N_1406);
and U1941 (N_1941,N_1468,N_1372);
nor U1942 (N_1942,N_1146,N_1170);
and U1943 (N_1943,N_794,N_795);
nand U1944 (N_1944,N_751,N_1167);
nand U1945 (N_1945,N_1189,N_908);
and U1946 (N_1946,N_1479,N_1240);
and U1947 (N_1947,N_811,N_771);
nand U1948 (N_1948,N_1350,N_1216);
nor U1949 (N_1949,N_1309,N_1312);
or U1950 (N_1950,N_1062,N_1282);
nand U1951 (N_1951,N_867,N_881);
nand U1952 (N_1952,N_1304,N_1005);
nor U1953 (N_1953,N_1370,N_1217);
xor U1954 (N_1954,N_812,N_1176);
and U1955 (N_1955,N_1208,N_1147);
or U1956 (N_1956,N_869,N_1427);
or U1957 (N_1957,N_1222,N_1259);
or U1958 (N_1958,N_831,N_1408);
nor U1959 (N_1959,N_1150,N_822);
nor U1960 (N_1960,N_1290,N_1380);
or U1961 (N_1961,N_1163,N_1349);
or U1962 (N_1962,N_1185,N_1290);
or U1963 (N_1963,N_883,N_1038);
nor U1964 (N_1964,N_800,N_1197);
nor U1965 (N_1965,N_1125,N_833);
or U1966 (N_1966,N_1205,N_1448);
nand U1967 (N_1967,N_1415,N_1463);
or U1968 (N_1968,N_1216,N_1494);
or U1969 (N_1969,N_1264,N_859);
nor U1970 (N_1970,N_1097,N_1475);
nand U1971 (N_1971,N_1417,N_854);
nand U1972 (N_1972,N_770,N_1441);
nor U1973 (N_1973,N_1368,N_1049);
and U1974 (N_1974,N_1124,N_1497);
nor U1975 (N_1975,N_1196,N_1060);
or U1976 (N_1976,N_1498,N_761);
nand U1977 (N_1977,N_1271,N_1327);
nor U1978 (N_1978,N_1124,N_1270);
or U1979 (N_1979,N_845,N_957);
nor U1980 (N_1980,N_1243,N_1194);
nand U1981 (N_1981,N_770,N_962);
or U1982 (N_1982,N_1441,N_1236);
nand U1983 (N_1983,N_1186,N_1038);
and U1984 (N_1984,N_1313,N_1074);
or U1985 (N_1985,N_889,N_829);
nor U1986 (N_1986,N_870,N_1046);
or U1987 (N_1987,N_1037,N_1340);
nand U1988 (N_1988,N_895,N_807);
and U1989 (N_1989,N_931,N_1170);
nand U1990 (N_1990,N_839,N_1340);
nor U1991 (N_1991,N_967,N_1039);
or U1992 (N_1992,N_1174,N_1065);
nand U1993 (N_1993,N_846,N_1340);
and U1994 (N_1994,N_1228,N_1399);
and U1995 (N_1995,N_1354,N_1236);
and U1996 (N_1996,N_1040,N_910);
nand U1997 (N_1997,N_1163,N_1420);
nand U1998 (N_1998,N_1057,N_1121);
nand U1999 (N_1999,N_1120,N_1328);
and U2000 (N_2000,N_764,N_1309);
and U2001 (N_2001,N_975,N_1117);
nand U2002 (N_2002,N_1013,N_1287);
nor U2003 (N_2003,N_1383,N_1107);
nand U2004 (N_2004,N_1182,N_1141);
xor U2005 (N_2005,N_871,N_796);
or U2006 (N_2006,N_792,N_1159);
nand U2007 (N_2007,N_1110,N_1280);
nor U2008 (N_2008,N_1282,N_832);
nor U2009 (N_2009,N_1147,N_772);
and U2010 (N_2010,N_987,N_771);
nand U2011 (N_2011,N_1062,N_786);
and U2012 (N_2012,N_1397,N_879);
nand U2013 (N_2013,N_1415,N_841);
or U2014 (N_2014,N_1117,N_1471);
or U2015 (N_2015,N_1082,N_956);
nand U2016 (N_2016,N_793,N_1020);
nand U2017 (N_2017,N_1007,N_1312);
or U2018 (N_2018,N_908,N_1329);
or U2019 (N_2019,N_1309,N_1299);
nor U2020 (N_2020,N_1385,N_992);
or U2021 (N_2021,N_948,N_1005);
or U2022 (N_2022,N_1066,N_1441);
or U2023 (N_2023,N_799,N_885);
nand U2024 (N_2024,N_1456,N_1267);
nor U2025 (N_2025,N_1141,N_1419);
nor U2026 (N_2026,N_1468,N_928);
nor U2027 (N_2027,N_1322,N_1135);
nand U2028 (N_2028,N_1351,N_936);
and U2029 (N_2029,N_1261,N_1012);
nand U2030 (N_2030,N_1329,N_919);
nand U2031 (N_2031,N_965,N_869);
or U2032 (N_2032,N_773,N_1343);
nor U2033 (N_2033,N_1013,N_1289);
or U2034 (N_2034,N_1250,N_1074);
or U2035 (N_2035,N_966,N_1298);
nor U2036 (N_2036,N_828,N_813);
nand U2037 (N_2037,N_867,N_1294);
nor U2038 (N_2038,N_780,N_1223);
nand U2039 (N_2039,N_1102,N_1132);
or U2040 (N_2040,N_826,N_1035);
and U2041 (N_2041,N_779,N_768);
nand U2042 (N_2042,N_1347,N_980);
nor U2043 (N_2043,N_881,N_1263);
and U2044 (N_2044,N_785,N_756);
nand U2045 (N_2045,N_1472,N_1102);
and U2046 (N_2046,N_800,N_1133);
nor U2047 (N_2047,N_982,N_865);
nor U2048 (N_2048,N_1209,N_1055);
and U2049 (N_2049,N_1496,N_1268);
or U2050 (N_2050,N_1348,N_1340);
or U2051 (N_2051,N_877,N_849);
nand U2052 (N_2052,N_835,N_1154);
and U2053 (N_2053,N_1205,N_837);
xnor U2054 (N_2054,N_1439,N_769);
nand U2055 (N_2055,N_1403,N_1205);
nor U2056 (N_2056,N_869,N_1074);
or U2057 (N_2057,N_903,N_1360);
or U2058 (N_2058,N_1022,N_1159);
nand U2059 (N_2059,N_946,N_898);
or U2060 (N_2060,N_764,N_785);
and U2061 (N_2061,N_1068,N_820);
or U2062 (N_2062,N_1050,N_1210);
and U2063 (N_2063,N_875,N_1100);
nand U2064 (N_2064,N_1167,N_821);
and U2065 (N_2065,N_1075,N_1250);
and U2066 (N_2066,N_1041,N_763);
nor U2067 (N_2067,N_919,N_805);
xor U2068 (N_2068,N_1486,N_1306);
nor U2069 (N_2069,N_818,N_1141);
and U2070 (N_2070,N_1400,N_1192);
or U2071 (N_2071,N_1303,N_1087);
nand U2072 (N_2072,N_946,N_782);
or U2073 (N_2073,N_1486,N_1112);
nand U2074 (N_2074,N_910,N_1378);
and U2075 (N_2075,N_915,N_1142);
nor U2076 (N_2076,N_1151,N_1291);
nor U2077 (N_2077,N_1027,N_815);
nand U2078 (N_2078,N_1474,N_898);
or U2079 (N_2079,N_1315,N_1140);
xor U2080 (N_2080,N_879,N_861);
or U2081 (N_2081,N_1026,N_1266);
nand U2082 (N_2082,N_1161,N_1332);
nor U2083 (N_2083,N_1313,N_1377);
nand U2084 (N_2084,N_1473,N_767);
and U2085 (N_2085,N_1475,N_1498);
nor U2086 (N_2086,N_1025,N_808);
or U2087 (N_2087,N_1185,N_1115);
nand U2088 (N_2088,N_1289,N_1351);
nand U2089 (N_2089,N_765,N_1339);
nor U2090 (N_2090,N_920,N_780);
nor U2091 (N_2091,N_887,N_943);
nor U2092 (N_2092,N_754,N_1156);
and U2093 (N_2093,N_1093,N_1234);
and U2094 (N_2094,N_1365,N_1457);
nor U2095 (N_2095,N_1389,N_1120);
or U2096 (N_2096,N_1441,N_863);
and U2097 (N_2097,N_882,N_1088);
nand U2098 (N_2098,N_1005,N_1092);
and U2099 (N_2099,N_1090,N_1320);
or U2100 (N_2100,N_1072,N_1403);
or U2101 (N_2101,N_1460,N_1021);
or U2102 (N_2102,N_1289,N_1337);
nor U2103 (N_2103,N_1045,N_1217);
nor U2104 (N_2104,N_1119,N_1147);
nand U2105 (N_2105,N_913,N_802);
nor U2106 (N_2106,N_1157,N_785);
or U2107 (N_2107,N_972,N_1243);
nor U2108 (N_2108,N_1082,N_1471);
xor U2109 (N_2109,N_1070,N_1158);
nand U2110 (N_2110,N_1444,N_1091);
or U2111 (N_2111,N_1086,N_1214);
nor U2112 (N_2112,N_1312,N_766);
nor U2113 (N_2113,N_1257,N_1348);
nand U2114 (N_2114,N_1468,N_1119);
or U2115 (N_2115,N_1451,N_1350);
and U2116 (N_2116,N_1380,N_1119);
nor U2117 (N_2117,N_860,N_1229);
or U2118 (N_2118,N_784,N_1002);
or U2119 (N_2119,N_771,N_836);
nand U2120 (N_2120,N_1031,N_889);
or U2121 (N_2121,N_800,N_879);
nor U2122 (N_2122,N_1108,N_1123);
and U2123 (N_2123,N_1390,N_1291);
and U2124 (N_2124,N_1431,N_855);
and U2125 (N_2125,N_874,N_1393);
and U2126 (N_2126,N_936,N_958);
nand U2127 (N_2127,N_1243,N_988);
and U2128 (N_2128,N_1065,N_1227);
nor U2129 (N_2129,N_984,N_1233);
and U2130 (N_2130,N_1306,N_1370);
nand U2131 (N_2131,N_760,N_1262);
and U2132 (N_2132,N_911,N_1440);
or U2133 (N_2133,N_1461,N_1253);
or U2134 (N_2134,N_1464,N_1439);
nor U2135 (N_2135,N_1226,N_1219);
and U2136 (N_2136,N_1040,N_1323);
nand U2137 (N_2137,N_780,N_752);
nand U2138 (N_2138,N_1463,N_1316);
nor U2139 (N_2139,N_1387,N_1375);
and U2140 (N_2140,N_1008,N_1336);
nor U2141 (N_2141,N_813,N_1246);
and U2142 (N_2142,N_1071,N_1386);
nand U2143 (N_2143,N_1222,N_1252);
and U2144 (N_2144,N_1208,N_1401);
nor U2145 (N_2145,N_872,N_1078);
nor U2146 (N_2146,N_759,N_1051);
nand U2147 (N_2147,N_828,N_1058);
nor U2148 (N_2148,N_1280,N_1126);
or U2149 (N_2149,N_1049,N_820);
nand U2150 (N_2150,N_1201,N_951);
nand U2151 (N_2151,N_1142,N_1358);
nand U2152 (N_2152,N_791,N_1198);
nor U2153 (N_2153,N_1491,N_800);
nor U2154 (N_2154,N_1478,N_1056);
or U2155 (N_2155,N_1255,N_1332);
or U2156 (N_2156,N_1227,N_1422);
and U2157 (N_2157,N_835,N_1069);
and U2158 (N_2158,N_922,N_921);
nand U2159 (N_2159,N_1496,N_1000);
or U2160 (N_2160,N_1262,N_1325);
or U2161 (N_2161,N_1083,N_1394);
and U2162 (N_2162,N_1284,N_1019);
and U2163 (N_2163,N_830,N_943);
nor U2164 (N_2164,N_1439,N_1417);
or U2165 (N_2165,N_1130,N_843);
or U2166 (N_2166,N_1428,N_802);
or U2167 (N_2167,N_1130,N_783);
or U2168 (N_2168,N_1278,N_1068);
or U2169 (N_2169,N_1424,N_1239);
or U2170 (N_2170,N_974,N_1483);
nand U2171 (N_2171,N_1153,N_864);
nand U2172 (N_2172,N_1143,N_1402);
or U2173 (N_2173,N_1483,N_1444);
nor U2174 (N_2174,N_1187,N_991);
or U2175 (N_2175,N_1202,N_836);
or U2176 (N_2176,N_1066,N_927);
nand U2177 (N_2177,N_1358,N_1391);
xor U2178 (N_2178,N_1430,N_1177);
or U2179 (N_2179,N_1098,N_1472);
nand U2180 (N_2180,N_1038,N_921);
nor U2181 (N_2181,N_1039,N_1281);
and U2182 (N_2182,N_1046,N_1226);
or U2183 (N_2183,N_1342,N_1087);
or U2184 (N_2184,N_1128,N_1131);
nor U2185 (N_2185,N_1120,N_1074);
nand U2186 (N_2186,N_1242,N_1438);
nand U2187 (N_2187,N_1478,N_1384);
and U2188 (N_2188,N_1485,N_1475);
and U2189 (N_2189,N_1233,N_1085);
nand U2190 (N_2190,N_1059,N_1077);
nor U2191 (N_2191,N_841,N_845);
and U2192 (N_2192,N_1113,N_1423);
nand U2193 (N_2193,N_827,N_1460);
or U2194 (N_2194,N_1338,N_1041);
or U2195 (N_2195,N_1191,N_1420);
or U2196 (N_2196,N_1236,N_918);
nand U2197 (N_2197,N_1367,N_1088);
nand U2198 (N_2198,N_982,N_1132);
and U2199 (N_2199,N_1148,N_1221);
and U2200 (N_2200,N_1142,N_1369);
and U2201 (N_2201,N_1368,N_1198);
nor U2202 (N_2202,N_1244,N_1464);
nor U2203 (N_2203,N_1182,N_1184);
nor U2204 (N_2204,N_1036,N_1086);
nor U2205 (N_2205,N_1339,N_1296);
and U2206 (N_2206,N_905,N_1417);
nand U2207 (N_2207,N_1303,N_1244);
nor U2208 (N_2208,N_867,N_860);
xor U2209 (N_2209,N_1463,N_1188);
nor U2210 (N_2210,N_1271,N_956);
nor U2211 (N_2211,N_908,N_1367);
nor U2212 (N_2212,N_1000,N_1256);
nand U2213 (N_2213,N_1421,N_833);
and U2214 (N_2214,N_1438,N_800);
or U2215 (N_2215,N_1089,N_1254);
xnor U2216 (N_2216,N_1488,N_1123);
nand U2217 (N_2217,N_796,N_1076);
nand U2218 (N_2218,N_1074,N_1178);
or U2219 (N_2219,N_960,N_959);
nor U2220 (N_2220,N_1085,N_1387);
or U2221 (N_2221,N_1282,N_1124);
nand U2222 (N_2222,N_933,N_1044);
nand U2223 (N_2223,N_1470,N_1182);
nor U2224 (N_2224,N_1448,N_829);
nand U2225 (N_2225,N_1385,N_1073);
nand U2226 (N_2226,N_797,N_1195);
or U2227 (N_2227,N_1391,N_1165);
nand U2228 (N_2228,N_767,N_1360);
nand U2229 (N_2229,N_816,N_822);
and U2230 (N_2230,N_803,N_830);
and U2231 (N_2231,N_1351,N_772);
or U2232 (N_2232,N_1454,N_1285);
or U2233 (N_2233,N_1214,N_1091);
or U2234 (N_2234,N_1422,N_1184);
nor U2235 (N_2235,N_1364,N_1046);
or U2236 (N_2236,N_1287,N_868);
nand U2237 (N_2237,N_1018,N_1495);
nor U2238 (N_2238,N_786,N_778);
nor U2239 (N_2239,N_1003,N_935);
or U2240 (N_2240,N_984,N_1062);
nand U2241 (N_2241,N_925,N_972);
or U2242 (N_2242,N_1339,N_871);
nor U2243 (N_2243,N_1421,N_1335);
or U2244 (N_2244,N_1309,N_816);
and U2245 (N_2245,N_1470,N_1218);
or U2246 (N_2246,N_795,N_1347);
nor U2247 (N_2247,N_1101,N_764);
or U2248 (N_2248,N_1369,N_1172);
xor U2249 (N_2249,N_845,N_760);
or U2250 (N_2250,N_2020,N_1928);
nand U2251 (N_2251,N_2206,N_1749);
nand U2252 (N_2252,N_1530,N_1876);
or U2253 (N_2253,N_2031,N_1835);
or U2254 (N_2254,N_1827,N_1939);
nor U2255 (N_2255,N_2017,N_1547);
nand U2256 (N_2256,N_2009,N_1762);
and U2257 (N_2257,N_1694,N_1802);
nand U2258 (N_2258,N_1846,N_2076);
and U2259 (N_2259,N_2142,N_1770);
and U2260 (N_2260,N_2063,N_2155);
and U2261 (N_2261,N_1851,N_1922);
and U2262 (N_2262,N_2146,N_1677);
nand U2263 (N_2263,N_2183,N_2164);
nor U2264 (N_2264,N_1648,N_1946);
or U2265 (N_2265,N_1535,N_1560);
xnor U2266 (N_2266,N_1572,N_2236);
nor U2267 (N_2267,N_2047,N_1746);
nor U2268 (N_2268,N_1951,N_1754);
and U2269 (N_2269,N_1532,N_1859);
nor U2270 (N_2270,N_1673,N_2062);
nor U2271 (N_2271,N_1760,N_1796);
and U2272 (N_2272,N_2098,N_2120);
nand U2273 (N_2273,N_1825,N_2054);
or U2274 (N_2274,N_2227,N_1515);
or U2275 (N_2275,N_1542,N_1929);
or U2276 (N_2276,N_1565,N_1660);
and U2277 (N_2277,N_1671,N_1863);
xor U2278 (N_2278,N_1892,N_1751);
nand U2279 (N_2279,N_2212,N_2088);
or U2280 (N_2280,N_1943,N_1785);
nor U2281 (N_2281,N_1653,N_2129);
and U2282 (N_2282,N_1901,N_1566);
nor U2283 (N_2283,N_1501,N_1799);
nor U2284 (N_2284,N_1812,N_2203);
nor U2285 (N_2285,N_2171,N_1744);
nor U2286 (N_2286,N_1644,N_2221);
or U2287 (N_2287,N_1878,N_2182);
nor U2288 (N_2288,N_1920,N_1781);
or U2289 (N_2289,N_2015,N_1769);
or U2290 (N_2290,N_1725,N_1557);
nor U2291 (N_2291,N_1521,N_1953);
or U2292 (N_2292,N_1803,N_1787);
and U2293 (N_2293,N_1964,N_2148);
nor U2294 (N_2294,N_1686,N_1674);
nand U2295 (N_2295,N_1693,N_1940);
nand U2296 (N_2296,N_2100,N_1767);
nand U2297 (N_2297,N_1942,N_1831);
or U2298 (N_2298,N_1748,N_1556);
nand U2299 (N_2299,N_1883,N_2166);
nor U2300 (N_2300,N_1675,N_2187);
or U2301 (N_2301,N_1524,N_2097);
nor U2302 (N_2302,N_1722,N_2083);
and U2303 (N_2303,N_1957,N_2176);
and U2304 (N_2304,N_2096,N_2213);
nand U2305 (N_2305,N_2133,N_1716);
nor U2306 (N_2306,N_2128,N_2215);
nor U2307 (N_2307,N_1982,N_1931);
and U2308 (N_2308,N_2150,N_2066);
and U2309 (N_2309,N_2030,N_1850);
or U2310 (N_2310,N_1585,N_1930);
nor U2311 (N_2311,N_1650,N_2130);
and U2312 (N_2312,N_2000,N_1840);
nor U2313 (N_2313,N_1807,N_1618);
nand U2314 (N_2314,N_2163,N_2021);
and U2315 (N_2315,N_1607,N_1571);
and U2316 (N_2316,N_1724,N_1527);
nand U2317 (N_2317,N_2121,N_2214);
nor U2318 (N_2318,N_1625,N_1670);
and U2319 (N_2319,N_1555,N_1634);
xor U2320 (N_2320,N_1509,N_1737);
and U2321 (N_2321,N_1741,N_1918);
nand U2322 (N_2322,N_2114,N_2105);
nand U2323 (N_2323,N_1913,N_2153);
nand U2324 (N_2324,N_1983,N_1643);
nand U2325 (N_2325,N_1981,N_1882);
or U2326 (N_2326,N_1755,N_1993);
nand U2327 (N_2327,N_2157,N_2209);
and U2328 (N_2328,N_1582,N_2075);
nand U2329 (N_2329,N_1632,N_2246);
xor U2330 (N_2330,N_2180,N_2074);
or U2331 (N_2331,N_1800,N_2044);
and U2332 (N_2332,N_1952,N_2177);
and U2333 (N_2333,N_1856,N_1868);
or U2334 (N_2334,N_1649,N_1717);
and U2335 (N_2335,N_2023,N_1646);
xnor U2336 (N_2336,N_1552,N_1534);
and U2337 (N_2337,N_1663,N_1962);
nor U2338 (N_2338,N_2041,N_2058);
or U2339 (N_2339,N_1814,N_1589);
and U2340 (N_2340,N_2011,N_1834);
and U2341 (N_2341,N_2205,N_1775);
or U2342 (N_2342,N_1742,N_1626);
or U2343 (N_2343,N_1898,N_1911);
nand U2344 (N_2344,N_1705,N_1645);
nand U2345 (N_2345,N_1761,N_2035);
nor U2346 (N_2346,N_1576,N_1688);
and U2347 (N_2347,N_1852,N_1699);
nor U2348 (N_2348,N_1975,N_2003);
nand U2349 (N_2349,N_2039,N_1786);
or U2350 (N_2350,N_2233,N_2081);
or U2351 (N_2351,N_2005,N_1641);
and U2352 (N_2352,N_1621,N_1619);
nor U2353 (N_2353,N_1804,N_1662);
nor U2354 (N_2354,N_2159,N_1906);
and U2355 (N_2355,N_2226,N_1638);
nand U2356 (N_2356,N_1847,N_1642);
and U2357 (N_2357,N_2043,N_2235);
or U2358 (N_2358,N_1551,N_2013);
nor U2359 (N_2359,N_1887,N_1733);
and U2360 (N_2360,N_2211,N_1708);
or U2361 (N_2361,N_1798,N_2022);
and U2362 (N_2362,N_2172,N_1895);
or U2363 (N_2363,N_2200,N_2190);
and U2364 (N_2364,N_1947,N_1777);
nor U2365 (N_2365,N_2145,N_1907);
nand U2366 (N_2366,N_2006,N_1541);
nand U2367 (N_2367,N_2012,N_1985);
nor U2368 (N_2368,N_1603,N_1558);
and U2369 (N_2369,N_1743,N_2199);
or U2370 (N_2370,N_2029,N_1941);
and U2371 (N_2371,N_1651,N_1680);
and U2372 (N_2372,N_2237,N_2124);
nand U2373 (N_2373,N_1845,N_1763);
or U2374 (N_2374,N_1961,N_1960);
nand U2375 (N_2375,N_2179,N_1602);
and U2376 (N_2376,N_1816,N_1734);
nor U2377 (N_2377,N_1606,N_2147);
and U2378 (N_2378,N_1806,N_1912);
and U2379 (N_2379,N_1706,N_1682);
and U2380 (N_2380,N_1696,N_1715);
nand U2381 (N_2381,N_2038,N_2077);
nand U2382 (N_2382,N_1658,N_1583);
nor U2383 (N_2383,N_1857,N_1996);
nand U2384 (N_2384,N_1932,N_1875);
nor U2385 (N_2385,N_2138,N_1709);
nand U2386 (N_2386,N_2067,N_1832);
or U2387 (N_2387,N_1844,N_2195);
or U2388 (N_2388,N_2061,N_1500);
or U2389 (N_2389,N_1679,N_1720);
nor U2390 (N_2390,N_1829,N_1639);
or U2391 (N_2391,N_1936,N_2109);
or U2392 (N_2392,N_2173,N_1593);
or U2393 (N_2393,N_2239,N_1885);
or U2394 (N_2394,N_1702,N_2104);
and U2395 (N_2395,N_1860,N_2079);
nor U2396 (N_2396,N_2089,N_2007);
nand U2397 (N_2397,N_1780,N_1504);
and U2398 (N_2398,N_1783,N_1886);
nor U2399 (N_2399,N_1672,N_1570);
nand U2400 (N_2400,N_1620,N_2071);
and U2401 (N_2401,N_1853,N_2135);
xor U2402 (N_2402,N_2117,N_1514);
and U2403 (N_2403,N_2032,N_1782);
or U2404 (N_2404,N_2095,N_1533);
nand U2405 (N_2405,N_2048,N_1976);
or U2406 (N_2406,N_2004,N_2132);
nand U2407 (N_2407,N_1575,N_1830);
nor U2408 (N_2408,N_1801,N_1977);
nand U2409 (N_2409,N_2119,N_2018);
nor U2410 (N_2410,N_1508,N_1869);
nand U2411 (N_2411,N_1897,N_2231);
and U2412 (N_2412,N_2094,N_2056);
and U2413 (N_2413,N_2069,N_2106);
nor U2414 (N_2414,N_1601,N_1750);
or U2415 (N_2415,N_2193,N_2181);
and U2416 (N_2416,N_2158,N_1959);
nand U2417 (N_2417,N_1854,N_2242);
nand U2418 (N_2418,N_1926,N_1788);
and U2419 (N_2419,N_1822,N_1537);
nor U2420 (N_2420,N_1948,N_1927);
and U2421 (N_2421,N_1910,N_2249);
nand U2422 (N_2422,N_1700,N_2191);
or U2423 (N_2423,N_1870,N_1721);
and U2424 (N_2424,N_1678,N_2188);
xnor U2425 (N_2425,N_1980,N_1969);
xor U2426 (N_2426,N_2101,N_2175);
nor U2427 (N_2427,N_1905,N_1924);
xnor U2428 (N_2428,N_1668,N_1810);
and U2429 (N_2429,N_1635,N_2168);
or U2430 (N_2430,N_2218,N_2025);
or U2431 (N_2431,N_2189,N_1880);
or U2432 (N_2432,N_2161,N_2238);
and U2433 (N_2433,N_2103,N_1609);
or U2434 (N_2434,N_1774,N_1684);
nand U2435 (N_2435,N_1992,N_2068);
or U2436 (N_2436,N_1776,N_1581);
nand U2437 (N_2437,N_2234,N_1511);
xor U2438 (N_2438,N_1838,N_2156);
or U2439 (N_2439,N_2241,N_1710);
or U2440 (N_2440,N_2049,N_2194);
nand U2441 (N_2441,N_1864,N_2116);
nand U2442 (N_2442,N_2202,N_2028);
xnor U2443 (N_2443,N_1934,N_1604);
and U2444 (N_2444,N_1937,N_1884);
nor U2445 (N_2445,N_1657,N_1974);
nor U2446 (N_2446,N_1998,N_2210);
nor U2447 (N_2447,N_1564,N_1797);
nor U2448 (N_2448,N_1595,N_1548);
or U2449 (N_2449,N_1971,N_1544);
nor U2450 (N_2450,N_2232,N_1756);
nand U2451 (N_2451,N_1766,N_2014);
nand U2452 (N_2452,N_1773,N_1656);
and U2453 (N_2453,N_2134,N_1888);
nand U2454 (N_2454,N_1889,N_2046);
nand U2455 (N_2455,N_1752,N_1711);
and U2456 (N_2456,N_1611,N_1861);
or U2457 (N_2457,N_2086,N_2151);
nand U2458 (N_2458,N_1768,N_1820);
nand U2459 (N_2459,N_1628,N_1567);
nand U2460 (N_2460,N_1669,N_1811);
and U2461 (N_2461,N_1818,N_1808);
or U2462 (N_2462,N_1989,N_1701);
nor U2463 (N_2463,N_1652,N_1622);
and U2464 (N_2464,N_2244,N_1784);
nand U2465 (N_2465,N_1554,N_1730);
nor U2466 (N_2466,N_2220,N_2092);
nand U2467 (N_2467,N_2186,N_2084);
or U2468 (N_2468,N_1970,N_1516);
nand U2469 (N_2469,N_2169,N_1624);
or U2470 (N_2470,N_1914,N_2115);
or U2471 (N_2471,N_1965,N_2126);
nand U2472 (N_2472,N_1938,N_1809);
and U2473 (N_2473,N_1915,N_2033);
nand U2474 (N_2474,N_2107,N_1614);
nand U2475 (N_2475,N_1713,N_1719);
and U2476 (N_2476,N_1950,N_1584);
and U2477 (N_2477,N_1600,N_2192);
or U2478 (N_2478,N_1654,N_1732);
or U2479 (N_2479,N_1529,N_2052);
nor U2480 (N_2480,N_2053,N_1973);
nand U2481 (N_2481,N_1902,N_1765);
nand U2482 (N_2482,N_1704,N_2051);
nor U2483 (N_2483,N_2162,N_2245);
xnor U2484 (N_2484,N_1823,N_1972);
nand U2485 (N_2485,N_1837,N_1740);
nor U2486 (N_2486,N_1608,N_1945);
and U2487 (N_2487,N_1828,N_1667);
nand U2488 (N_2488,N_1525,N_1685);
or U2489 (N_2489,N_2204,N_2174);
nor U2490 (N_2490,N_1877,N_2111);
and U2491 (N_2491,N_2059,N_2201);
and U2492 (N_2492,N_1518,N_2008);
or U2493 (N_2493,N_1712,N_1771);
or U2494 (N_2494,N_2170,N_2216);
and U2495 (N_2495,N_1545,N_1824);
and U2496 (N_2496,N_1731,N_1986);
nor U2497 (N_2497,N_2055,N_1736);
nor U2498 (N_2498,N_2152,N_2240);
nand U2499 (N_2499,N_1591,N_1687);
or U2500 (N_2500,N_1899,N_2073);
nor U2501 (N_2501,N_2167,N_2230);
nor U2502 (N_2502,N_1866,N_1578);
nand U2503 (N_2503,N_1563,N_1543);
or U2504 (N_2504,N_1935,N_1637);
or U2505 (N_2505,N_1689,N_1896);
nor U2506 (N_2506,N_2137,N_1963);
and U2507 (N_2507,N_1855,N_1862);
or U2508 (N_2508,N_1791,N_1598);
nand U2509 (N_2509,N_2144,N_1664);
nand U2510 (N_2510,N_1873,N_1903);
or U2511 (N_2511,N_2027,N_2208);
and U2512 (N_2512,N_1890,N_2110);
xnor U2513 (N_2513,N_2045,N_2184);
and U2514 (N_2514,N_1714,N_1954);
nand U2515 (N_2515,N_2198,N_1842);
nor U2516 (N_2516,N_1586,N_2091);
or U2517 (N_2517,N_1944,N_1617);
nor U2518 (N_2518,N_1958,N_1997);
and U2519 (N_2519,N_2225,N_1553);
or U2520 (N_2520,N_1596,N_1647);
and U2521 (N_2521,N_1549,N_2065);
nor U2522 (N_2522,N_1627,N_1655);
or U2523 (N_2523,N_1729,N_1728);
nor U2524 (N_2524,N_2219,N_2143);
and U2525 (N_2525,N_1753,N_1616);
nand U2526 (N_2526,N_1574,N_2136);
and U2527 (N_2527,N_1908,N_1718);
and U2528 (N_2528,N_1523,N_2016);
nor U2529 (N_2529,N_1605,N_1988);
and U2530 (N_2530,N_2248,N_2040);
and U2531 (N_2531,N_1629,N_1817);
or U2532 (N_2532,N_1921,N_2178);
nor U2533 (N_2533,N_1833,N_1550);
nand U2534 (N_2534,N_2222,N_1592);
and U2535 (N_2535,N_2064,N_2149);
nand U2536 (N_2536,N_2224,N_1949);
or U2537 (N_2537,N_1795,N_1841);
nor U2538 (N_2538,N_1539,N_1967);
nand U2539 (N_2539,N_1790,N_1610);
nor U2540 (N_2540,N_1821,N_2093);
or U2541 (N_2541,N_1999,N_1665);
nor U2542 (N_2542,N_2113,N_2122);
nor U2543 (N_2543,N_1568,N_2160);
nor U2544 (N_2544,N_1502,N_1994);
nand U2545 (N_2545,N_1612,N_1506);
nor U2546 (N_2546,N_1789,N_1503);
nor U2547 (N_2547,N_1893,N_1538);
or U2548 (N_2548,N_1698,N_1874);
nand U2549 (N_2549,N_1735,N_2154);
or U2550 (N_2550,N_1703,N_1917);
or U2551 (N_2551,N_1745,N_1633);
nand U2552 (N_2552,N_1546,N_1793);
or U2553 (N_2553,N_1759,N_2002);
nor U2554 (N_2554,N_1805,N_1848);
nor U2555 (N_2555,N_2197,N_2036);
nand U2556 (N_2556,N_1519,N_2141);
and U2557 (N_2557,N_1881,N_1562);
nand U2558 (N_2558,N_1978,N_1531);
or U2559 (N_2559,N_1956,N_1510);
or U2560 (N_2560,N_1692,N_1727);
nor U2561 (N_2561,N_1577,N_1738);
nor U2562 (N_2562,N_1758,N_1690);
nor U2563 (N_2563,N_1615,N_1858);
nor U2564 (N_2564,N_2217,N_1849);
and U2565 (N_2565,N_1826,N_1588);
or U2566 (N_2566,N_1879,N_1933);
xnor U2567 (N_2567,N_2024,N_1995);
or U2568 (N_2568,N_2034,N_1512);
nor U2569 (N_2569,N_1587,N_1630);
nor U2570 (N_2570,N_2223,N_2243);
nor U2571 (N_2571,N_1872,N_2050);
or U2572 (N_2572,N_2057,N_2125);
nand U2573 (N_2573,N_1517,N_1779);
nor U2574 (N_2574,N_1505,N_1909);
or U2575 (N_2575,N_2207,N_1815);
xor U2576 (N_2576,N_1526,N_2118);
nand U2577 (N_2577,N_1676,N_1636);
nand U2578 (N_2578,N_1867,N_2090);
nor U2579 (N_2579,N_1990,N_1987);
nor U2580 (N_2580,N_1661,N_1979);
and U2581 (N_2581,N_2072,N_1925);
nor U2582 (N_2582,N_1916,N_1561);
nor U2583 (N_2583,N_2087,N_1613);
and U2584 (N_2584,N_1747,N_1659);
or U2585 (N_2585,N_1772,N_1683);
nand U2586 (N_2586,N_1640,N_2010);
and U2587 (N_2587,N_1955,N_1697);
nor U2588 (N_2588,N_2112,N_1623);
and U2589 (N_2589,N_1792,N_2228);
nor U2590 (N_2590,N_1984,N_1764);
or U2591 (N_2591,N_1778,N_1968);
xnor U2592 (N_2592,N_2026,N_1739);
or U2593 (N_2593,N_2102,N_2140);
or U2594 (N_2594,N_2070,N_1569);
nor U2595 (N_2595,N_1707,N_1597);
or U2596 (N_2596,N_1666,N_1923);
nand U2597 (N_2597,N_2165,N_2080);
nor U2598 (N_2598,N_1559,N_1522);
or U2599 (N_2599,N_1580,N_2085);
and U2600 (N_2600,N_1599,N_2060);
nand U2601 (N_2601,N_1513,N_1894);
or U2602 (N_2602,N_1540,N_1966);
or U2603 (N_2603,N_1590,N_1594);
nor U2604 (N_2604,N_1726,N_1919);
nand U2605 (N_2605,N_1871,N_1839);
nor U2606 (N_2606,N_2127,N_2037);
nand U2607 (N_2607,N_1681,N_1813);
nand U2608 (N_2608,N_1900,N_1836);
nor U2609 (N_2609,N_1536,N_1757);
nor U2610 (N_2610,N_2123,N_2131);
nand U2611 (N_2611,N_2042,N_2108);
and U2612 (N_2612,N_1865,N_1507);
nor U2613 (N_2613,N_1723,N_2247);
nor U2614 (N_2614,N_2078,N_1579);
or U2615 (N_2615,N_2229,N_1794);
and U2616 (N_2616,N_1528,N_1819);
nand U2617 (N_2617,N_1691,N_2019);
nor U2618 (N_2618,N_1843,N_2185);
nand U2619 (N_2619,N_2082,N_1520);
nand U2620 (N_2620,N_1573,N_2196);
nand U2621 (N_2621,N_1695,N_1904);
nand U2622 (N_2622,N_2139,N_1891);
nor U2623 (N_2623,N_2001,N_2099);
xnor U2624 (N_2624,N_1991,N_1631);
xnor U2625 (N_2625,N_1742,N_1987);
nand U2626 (N_2626,N_1594,N_1608);
or U2627 (N_2627,N_2144,N_2038);
or U2628 (N_2628,N_1751,N_2153);
nor U2629 (N_2629,N_2109,N_1759);
and U2630 (N_2630,N_1508,N_2159);
nor U2631 (N_2631,N_1974,N_2183);
and U2632 (N_2632,N_1568,N_1958);
nor U2633 (N_2633,N_2053,N_2043);
nor U2634 (N_2634,N_1601,N_1549);
nor U2635 (N_2635,N_2122,N_1742);
nor U2636 (N_2636,N_2069,N_2052);
nor U2637 (N_2637,N_1659,N_1539);
and U2638 (N_2638,N_2098,N_2090);
nand U2639 (N_2639,N_1946,N_1728);
and U2640 (N_2640,N_1951,N_1864);
and U2641 (N_2641,N_2186,N_2236);
nor U2642 (N_2642,N_1591,N_2209);
nor U2643 (N_2643,N_2142,N_2017);
nor U2644 (N_2644,N_2100,N_1549);
nand U2645 (N_2645,N_1878,N_2163);
nand U2646 (N_2646,N_2065,N_1653);
or U2647 (N_2647,N_2036,N_1863);
nor U2648 (N_2648,N_2138,N_2202);
or U2649 (N_2649,N_1566,N_2116);
or U2650 (N_2650,N_1844,N_1747);
nor U2651 (N_2651,N_1581,N_2209);
nor U2652 (N_2652,N_1787,N_1579);
nor U2653 (N_2653,N_2051,N_1608);
nand U2654 (N_2654,N_1732,N_2127);
nand U2655 (N_2655,N_2245,N_2154);
nand U2656 (N_2656,N_2002,N_1590);
or U2657 (N_2657,N_1524,N_2112);
and U2658 (N_2658,N_1614,N_2081);
nor U2659 (N_2659,N_2199,N_1925);
and U2660 (N_2660,N_1544,N_2037);
or U2661 (N_2661,N_1691,N_2042);
nor U2662 (N_2662,N_1821,N_1889);
nand U2663 (N_2663,N_1790,N_1548);
nor U2664 (N_2664,N_1699,N_1715);
nand U2665 (N_2665,N_1541,N_1836);
and U2666 (N_2666,N_2228,N_2203);
nor U2667 (N_2667,N_1622,N_2055);
and U2668 (N_2668,N_2010,N_1866);
or U2669 (N_2669,N_1991,N_2017);
nand U2670 (N_2670,N_1532,N_1713);
nand U2671 (N_2671,N_1658,N_2071);
nand U2672 (N_2672,N_1773,N_2234);
nor U2673 (N_2673,N_1557,N_1747);
nor U2674 (N_2674,N_2178,N_1674);
nand U2675 (N_2675,N_1517,N_1847);
and U2676 (N_2676,N_2188,N_1877);
or U2677 (N_2677,N_1550,N_2089);
nor U2678 (N_2678,N_1515,N_1626);
and U2679 (N_2679,N_1978,N_2219);
nand U2680 (N_2680,N_1751,N_1780);
or U2681 (N_2681,N_2198,N_2019);
nand U2682 (N_2682,N_2090,N_1606);
nor U2683 (N_2683,N_2095,N_1609);
nand U2684 (N_2684,N_2201,N_2048);
nand U2685 (N_2685,N_1651,N_2042);
nor U2686 (N_2686,N_1958,N_2181);
and U2687 (N_2687,N_1879,N_1851);
nand U2688 (N_2688,N_2234,N_1766);
nand U2689 (N_2689,N_2100,N_1880);
nor U2690 (N_2690,N_1677,N_1553);
and U2691 (N_2691,N_1709,N_1549);
nand U2692 (N_2692,N_2005,N_2085);
or U2693 (N_2693,N_2009,N_1885);
or U2694 (N_2694,N_2126,N_1788);
or U2695 (N_2695,N_1710,N_2084);
nor U2696 (N_2696,N_2219,N_1827);
nand U2697 (N_2697,N_2153,N_2221);
or U2698 (N_2698,N_2007,N_1551);
nand U2699 (N_2699,N_1840,N_1521);
or U2700 (N_2700,N_2073,N_2099);
or U2701 (N_2701,N_2221,N_2216);
and U2702 (N_2702,N_1586,N_1868);
nor U2703 (N_2703,N_1814,N_1555);
xor U2704 (N_2704,N_1680,N_1996);
or U2705 (N_2705,N_1626,N_2131);
nor U2706 (N_2706,N_2163,N_1520);
nor U2707 (N_2707,N_1826,N_1531);
and U2708 (N_2708,N_1550,N_2243);
nor U2709 (N_2709,N_1820,N_2190);
or U2710 (N_2710,N_2072,N_1713);
or U2711 (N_2711,N_2064,N_1845);
or U2712 (N_2712,N_1838,N_1866);
nor U2713 (N_2713,N_1925,N_1602);
and U2714 (N_2714,N_1535,N_1980);
nor U2715 (N_2715,N_1735,N_1684);
nor U2716 (N_2716,N_1696,N_1571);
nand U2717 (N_2717,N_1636,N_1783);
nand U2718 (N_2718,N_2103,N_1635);
or U2719 (N_2719,N_1637,N_2017);
nand U2720 (N_2720,N_1967,N_1506);
nand U2721 (N_2721,N_1513,N_1929);
and U2722 (N_2722,N_2189,N_1779);
or U2723 (N_2723,N_2058,N_2228);
nor U2724 (N_2724,N_1591,N_1836);
nor U2725 (N_2725,N_1807,N_1690);
nor U2726 (N_2726,N_1961,N_2055);
nand U2727 (N_2727,N_1642,N_2219);
nand U2728 (N_2728,N_2044,N_1872);
nand U2729 (N_2729,N_1903,N_1939);
nor U2730 (N_2730,N_1726,N_2193);
and U2731 (N_2731,N_1603,N_2209);
nor U2732 (N_2732,N_1815,N_2054);
and U2733 (N_2733,N_1851,N_2066);
nand U2734 (N_2734,N_1852,N_1814);
and U2735 (N_2735,N_2168,N_1541);
nand U2736 (N_2736,N_1614,N_2171);
nand U2737 (N_2737,N_1673,N_1919);
and U2738 (N_2738,N_1954,N_1899);
nor U2739 (N_2739,N_2187,N_1897);
nor U2740 (N_2740,N_1505,N_1625);
nor U2741 (N_2741,N_1523,N_1780);
or U2742 (N_2742,N_1921,N_2018);
or U2743 (N_2743,N_1714,N_1524);
nor U2744 (N_2744,N_2088,N_1601);
nor U2745 (N_2745,N_2112,N_2217);
or U2746 (N_2746,N_1969,N_1849);
and U2747 (N_2747,N_1983,N_1602);
nor U2748 (N_2748,N_1512,N_2075);
nor U2749 (N_2749,N_1998,N_2091);
nor U2750 (N_2750,N_1953,N_1559);
and U2751 (N_2751,N_2146,N_1930);
nand U2752 (N_2752,N_1879,N_1548);
and U2753 (N_2753,N_2073,N_1721);
nor U2754 (N_2754,N_1545,N_1875);
xnor U2755 (N_2755,N_1550,N_1864);
or U2756 (N_2756,N_1760,N_1895);
and U2757 (N_2757,N_2058,N_1507);
nand U2758 (N_2758,N_1502,N_1911);
nor U2759 (N_2759,N_1635,N_2148);
xnor U2760 (N_2760,N_1990,N_2162);
nand U2761 (N_2761,N_1627,N_1978);
nor U2762 (N_2762,N_1627,N_2070);
or U2763 (N_2763,N_1599,N_1571);
and U2764 (N_2764,N_1935,N_1875);
or U2765 (N_2765,N_1844,N_2234);
nor U2766 (N_2766,N_2191,N_1972);
nor U2767 (N_2767,N_1506,N_1944);
or U2768 (N_2768,N_1994,N_2194);
or U2769 (N_2769,N_1983,N_2232);
nor U2770 (N_2770,N_2182,N_1680);
and U2771 (N_2771,N_1781,N_1778);
nand U2772 (N_2772,N_2097,N_1867);
nand U2773 (N_2773,N_1792,N_2085);
nor U2774 (N_2774,N_1574,N_1783);
nor U2775 (N_2775,N_1927,N_1589);
nand U2776 (N_2776,N_1769,N_1825);
nand U2777 (N_2777,N_1675,N_1819);
and U2778 (N_2778,N_1982,N_1600);
or U2779 (N_2779,N_1529,N_1881);
and U2780 (N_2780,N_1708,N_1659);
or U2781 (N_2781,N_1939,N_1720);
or U2782 (N_2782,N_1958,N_2136);
nor U2783 (N_2783,N_2157,N_2221);
nor U2784 (N_2784,N_1773,N_2188);
or U2785 (N_2785,N_1865,N_2012);
nand U2786 (N_2786,N_1942,N_1721);
nand U2787 (N_2787,N_1828,N_2137);
nor U2788 (N_2788,N_1777,N_1576);
and U2789 (N_2789,N_1935,N_1782);
and U2790 (N_2790,N_1596,N_1945);
xor U2791 (N_2791,N_2010,N_1868);
nor U2792 (N_2792,N_2018,N_2135);
nand U2793 (N_2793,N_1903,N_1579);
nand U2794 (N_2794,N_1584,N_2055);
nor U2795 (N_2795,N_1954,N_1692);
xnor U2796 (N_2796,N_1561,N_2164);
nand U2797 (N_2797,N_1978,N_1838);
nand U2798 (N_2798,N_1749,N_2143);
nand U2799 (N_2799,N_1641,N_1598);
or U2800 (N_2800,N_1555,N_1901);
nand U2801 (N_2801,N_1658,N_1969);
and U2802 (N_2802,N_2027,N_1507);
or U2803 (N_2803,N_2205,N_1807);
nand U2804 (N_2804,N_1540,N_2188);
or U2805 (N_2805,N_2212,N_1742);
and U2806 (N_2806,N_1971,N_1906);
and U2807 (N_2807,N_1798,N_2114);
and U2808 (N_2808,N_1965,N_2143);
or U2809 (N_2809,N_1724,N_1805);
and U2810 (N_2810,N_1918,N_1515);
nor U2811 (N_2811,N_2034,N_2132);
nor U2812 (N_2812,N_2125,N_1590);
xor U2813 (N_2813,N_2132,N_2085);
nor U2814 (N_2814,N_2072,N_1921);
or U2815 (N_2815,N_1585,N_1676);
nor U2816 (N_2816,N_1795,N_1567);
nor U2817 (N_2817,N_2199,N_1916);
or U2818 (N_2818,N_2187,N_1535);
or U2819 (N_2819,N_2105,N_1918);
or U2820 (N_2820,N_1694,N_1842);
and U2821 (N_2821,N_1990,N_1715);
or U2822 (N_2822,N_1666,N_1922);
nand U2823 (N_2823,N_1925,N_1771);
nand U2824 (N_2824,N_2029,N_1804);
and U2825 (N_2825,N_2116,N_1502);
nand U2826 (N_2826,N_2114,N_1822);
nor U2827 (N_2827,N_2161,N_1622);
nand U2828 (N_2828,N_1528,N_2045);
nand U2829 (N_2829,N_1831,N_1877);
nand U2830 (N_2830,N_2027,N_1885);
or U2831 (N_2831,N_2149,N_1830);
and U2832 (N_2832,N_2242,N_1669);
nand U2833 (N_2833,N_1614,N_2109);
or U2834 (N_2834,N_1778,N_1931);
nand U2835 (N_2835,N_1757,N_1878);
nand U2836 (N_2836,N_1659,N_1931);
nand U2837 (N_2837,N_1562,N_1874);
xnor U2838 (N_2838,N_2191,N_2241);
nand U2839 (N_2839,N_2005,N_2178);
nand U2840 (N_2840,N_1811,N_1553);
nand U2841 (N_2841,N_1538,N_1532);
nor U2842 (N_2842,N_2200,N_1909);
nor U2843 (N_2843,N_2189,N_2018);
xnor U2844 (N_2844,N_1810,N_2082);
and U2845 (N_2845,N_1679,N_1564);
nor U2846 (N_2846,N_2156,N_1571);
nor U2847 (N_2847,N_1894,N_2057);
nand U2848 (N_2848,N_2244,N_1544);
nor U2849 (N_2849,N_2137,N_1860);
and U2850 (N_2850,N_1817,N_1788);
or U2851 (N_2851,N_1694,N_1570);
or U2852 (N_2852,N_1507,N_1540);
nand U2853 (N_2853,N_1898,N_2044);
nand U2854 (N_2854,N_1768,N_1907);
nor U2855 (N_2855,N_1566,N_1932);
nand U2856 (N_2856,N_2125,N_1887);
nand U2857 (N_2857,N_2125,N_1731);
nand U2858 (N_2858,N_2003,N_1788);
nand U2859 (N_2859,N_2151,N_2019);
and U2860 (N_2860,N_1634,N_1874);
or U2861 (N_2861,N_1658,N_1736);
nand U2862 (N_2862,N_1712,N_1753);
and U2863 (N_2863,N_1952,N_1564);
and U2864 (N_2864,N_1617,N_2239);
and U2865 (N_2865,N_1616,N_1641);
and U2866 (N_2866,N_2227,N_1622);
or U2867 (N_2867,N_1556,N_2086);
nor U2868 (N_2868,N_1882,N_1800);
or U2869 (N_2869,N_1541,N_1748);
nor U2870 (N_2870,N_2061,N_1780);
and U2871 (N_2871,N_1858,N_1631);
or U2872 (N_2872,N_2198,N_1734);
and U2873 (N_2873,N_1642,N_1879);
nand U2874 (N_2874,N_1800,N_1781);
nand U2875 (N_2875,N_2011,N_1704);
nand U2876 (N_2876,N_2116,N_1774);
nor U2877 (N_2877,N_1679,N_1627);
or U2878 (N_2878,N_1712,N_1776);
nor U2879 (N_2879,N_1744,N_2017);
nor U2880 (N_2880,N_1758,N_1870);
nor U2881 (N_2881,N_2133,N_1635);
nand U2882 (N_2882,N_2103,N_1944);
nor U2883 (N_2883,N_2164,N_1694);
and U2884 (N_2884,N_2063,N_2123);
nand U2885 (N_2885,N_1630,N_2012);
and U2886 (N_2886,N_2201,N_2106);
and U2887 (N_2887,N_2171,N_1594);
nand U2888 (N_2888,N_1550,N_1881);
or U2889 (N_2889,N_1828,N_1940);
nor U2890 (N_2890,N_1941,N_2154);
nor U2891 (N_2891,N_1925,N_1596);
or U2892 (N_2892,N_1740,N_1994);
and U2893 (N_2893,N_1824,N_1663);
or U2894 (N_2894,N_2222,N_1923);
or U2895 (N_2895,N_2199,N_1761);
or U2896 (N_2896,N_1543,N_1634);
nand U2897 (N_2897,N_2118,N_1890);
nand U2898 (N_2898,N_1619,N_1797);
or U2899 (N_2899,N_2031,N_2085);
nand U2900 (N_2900,N_2153,N_2037);
nand U2901 (N_2901,N_2216,N_1976);
nand U2902 (N_2902,N_1504,N_1622);
and U2903 (N_2903,N_1976,N_1503);
nor U2904 (N_2904,N_1641,N_1758);
nor U2905 (N_2905,N_2004,N_1931);
nor U2906 (N_2906,N_2160,N_2081);
xnor U2907 (N_2907,N_1897,N_2013);
nor U2908 (N_2908,N_1567,N_2011);
and U2909 (N_2909,N_2138,N_2223);
nand U2910 (N_2910,N_1734,N_1866);
nand U2911 (N_2911,N_1828,N_2119);
and U2912 (N_2912,N_1516,N_1952);
and U2913 (N_2913,N_1758,N_2230);
or U2914 (N_2914,N_1784,N_1936);
nand U2915 (N_2915,N_2109,N_2128);
nand U2916 (N_2916,N_2072,N_2007);
nand U2917 (N_2917,N_2223,N_2014);
or U2918 (N_2918,N_2139,N_1790);
and U2919 (N_2919,N_1801,N_2202);
or U2920 (N_2920,N_2049,N_1977);
xnor U2921 (N_2921,N_1510,N_1606);
and U2922 (N_2922,N_2035,N_1537);
nand U2923 (N_2923,N_1984,N_2053);
nor U2924 (N_2924,N_1617,N_2079);
nand U2925 (N_2925,N_2235,N_1880);
xor U2926 (N_2926,N_2206,N_1907);
nand U2927 (N_2927,N_1739,N_1880);
nand U2928 (N_2928,N_1631,N_1565);
and U2929 (N_2929,N_2107,N_1568);
nor U2930 (N_2930,N_1536,N_1563);
nor U2931 (N_2931,N_2214,N_2100);
nor U2932 (N_2932,N_2229,N_1830);
nor U2933 (N_2933,N_1535,N_2074);
nand U2934 (N_2934,N_2031,N_1892);
or U2935 (N_2935,N_1953,N_2223);
nand U2936 (N_2936,N_1740,N_1724);
or U2937 (N_2937,N_1814,N_1697);
or U2938 (N_2938,N_2186,N_1696);
nor U2939 (N_2939,N_2007,N_2206);
nand U2940 (N_2940,N_1503,N_2042);
nand U2941 (N_2941,N_1651,N_1531);
or U2942 (N_2942,N_2135,N_2205);
or U2943 (N_2943,N_1953,N_2052);
or U2944 (N_2944,N_1622,N_2054);
and U2945 (N_2945,N_1869,N_1827);
or U2946 (N_2946,N_2159,N_1633);
and U2947 (N_2947,N_1785,N_2172);
nand U2948 (N_2948,N_2229,N_2078);
xnor U2949 (N_2949,N_1991,N_1866);
nand U2950 (N_2950,N_1651,N_1592);
and U2951 (N_2951,N_1758,N_1970);
nand U2952 (N_2952,N_2024,N_1975);
nand U2953 (N_2953,N_1565,N_2215);
nor U2954 (N_2954,N_2001,N_1968);
nand U2955 (N_2955,N_2129,N_2192);
nor U2956 (N_2956,N_1888,N_1765);
or U2957 (N_2957,N_1892,N_1635);
nor U2958 (N_2958,N_2180,N_1620);
and U2959 (N_2959,N_1718,N_1874);
or U2960 (N_2960,N_2240,N_1638);
or U2961 (N_2961,N_2146,N_1758);
nor U2962 (N_2962,N_1586,N_1598);
xnor U2963 (N_2963,N_2048,N_1986);
nor U2964 (N_2964,N_2093,N_1928);
or U2965 (N_2965,N_2020,N_1721);
nand U2966 (N_2966,N_1656,N_1673);
and U2967 (N_2967,N_2056,N_2049);
or U2968 (N_2968,N_1829,N_1684);
nor U2969 (N_2969,N_1802,N_2133);
xnor U2970 (N_2970,N_1564,N_2100);
and U2971 (N_2971,N_1859,N_2198);
nor U2972 (N_2972,N_1828,N_1880);
nor U2973 (N_2973,N_2108,N_1867);
or U2974 (N_2974,N_1873,N_1961);
xnor U2975 (N_2975,N_1949,N_2175);
nand U2976 (N_2976,N_2013,N_2222);
and U2977 (N_2977,N_1838,N_1518);
nor U2978 (N_2978,N_2045,N_1852);
and U2979 (N_2979,N_1820,N_1801);
and U2980 (N_2980,N_1580,N_1662);
nand U2981 (N_2981,N_1585,N_1870);
and U2982 (N_2982,N_1818,N_1813);
and U2983 (N_2983,N_2113,N_2204);
and U2984 (N_2984,N_1818,N_1851);
nor U2985 (N_2985,N_1705,N_1536);
nand U2986 (N_2986,N_1549,N_1894);
nand U2987 (N_2987,N_2056,N_1775);
or U2988 (N_2988,N_1919,N_2129);
nand U2989 (N_2989,N_2195,N_1986);
or U2990 (N_2990,N_2032,N_1855);
nand U2991 (N_2991,N_2233,N_1591);
nand U2992 (N_2992,N_2084,N_1642);
or U2993 (N_2993,N_1630,N_1774);
or U2994 (N_2994,N_1619,N_2154);
nand U2995 (N_2995,N_1991,N_1861);
and U2996 (N_2996,N_1677,N_2218);
and U2997 (N_2997,N_1612,N_1858);
xor U2998 (N_2998,N_2212,N_1640);
nand U2999 (N_2999,N_1738,N_2188);
and UO_0 (O_0,N_2882,N_2888);
nand UO_1 (O_1,N_2908,N_2275);
nor UO_2 (O_2,N_2490,N_2460);
or UO_3 (O_3,N_2293,N_2943);
nand UO_4 (O_4,N_2349,N_2594);
and UO_5 (O_5,N_2565,N_2622);
or UO_6 (O_6,N_2392,N_2376);
nand UO_7 (O_7,N_2590,N_2328);
or UO_8 (O_8,N_2385,N_2756);
nor UO_9 (O_9,N_2901,N_2654);
nand UO_10 (O_10,N_2833,N_2981);
or UO_11 (O_11,N_2386,N_2475);
or UO_12 (O_12,N_2874,N_2842);
nor UO_13 (O_13,N_2628,N_2303);
and UO_14 (O_14,N_2442,N_2387);
and UO_15 (O_15,N_2734,N_2689);
and UO_16 (O_16,N_2600,N_2671);
or UO_17 (O_17,N_2843,N_2714);
and UO_18 (O_18,N_2423,N_2481);
nor UO_19 (O_19,N_2408,N_2838);
nor UO_20 (O_20,N_2958,N_2320);
or UO_21 (O_21,N_2634,N_2496);
and UO_22 (O_22,N_2401,N_2782);
nor UO_23 (O_23,N_2538,N_2429);
or UO_24 (O_24,N_2798,N_2961);
or UO_25 (O_25,N_2934,N_2727);
and UO_26 (O_26,N_2873,N_2801);
or UO_27 (O_27,N_2891,N_2695);
nor UO_28 (O_28,N_2643,N_2662);
or UO_29 (O_29,N_2664,N_2911);
nand UO_30 (O_30,N_2732,N_2630);
and UO_31 (O_31,N_2862,N_2332);
or UO_32 (O_32,N_2399,N_2375);
or UO_33 (O_33,N_2347,N_2315);
nand UO_34 (O_34,N_2716,N_2489);
or UO_35 (O_35,N_2892,N_2825);
and UO_36 (O_36,N_2897,N_2517);
or UO_37 (O_37,N_2639,N_2933);
and UO_38 (O_38,N_2614,N_2415);
nor UO_39 (O_39,N_2729,N_2304);
nor UO_40 (O_40,N_2640,N_2356);
nand UO_41 (O_41,N_2661,N_2709);
xor UO_42 (O_42,N_2260,N_2972);
nand UO_43 (O_43,N_2635,N_2333);
nor UO_44 (O_44,N_2395,N_2780);
nand UO_45 (O_45,N_2866,N_2339);
nor UO_46 (O_46,N_2353,N_2667);
and UO_47 (O_47,N_2849,N_2301);
or UO_48 (O_48,N_2726,N_2769);
nand UO_49 (O_49,N_2510,N_2577);
or UO_50 (O_50,N_2827,N_2438);
nand UO_51 (O_51,N_2354,N_2850);
nor UO_52 (O_52,N_2751,N_2997);
or UO_53 (O_53,N_2610,N_2504);
or UO_54 (O_54,N_2644,N_2567);
and UO_55 (O_55,N_2281,N_2461);
and UO_56 (O_56,N_2425,N_2306);
and UO_57 (O_57,N_2403,N_2605);
nor UO_58 (O_58,N_2529,N_2291);
or UO_59 (O_59,N_2251,N_2717);
nor UO_60 (O_60,N_2578,N_2784);
or UO_61 (O_61,N_2521,N_2334);
nand UO_62 (O_62,N_2525,N_2995);
nor UO_63 (O_63,N_2559,N_2868);
nand UO_64 (O_64,N_2730,N_2791);
and UO_65 (O_65,N_2542,N_2712);
nand UO_66 (O_66,N_2816,N_2852);
and UO_67 (O_67,N_2450,N_2469);
or UO_68 (O_68,N_2571,N_2956);
or UO_69 (O_69,N_2651,N_2471);
nor UO_70 (O_70,N_2337,N_2417);
nor UO_71 (O_71,N_2487,N_2407);
nor UO_72 (O_72,N_2418,N_2276);
nor UO_73 (O_73,N_2267,N_2674);
and UO_74 (O_74,N_2338,N_2533);
and UO_75 (O_75,N_2938,N_2994);
and UO_76 (O_76,N_2677,N_2980);
nand UO_77 (O_77,N_2700,N_2327);
nand UO_78 (O_78,N_2885,N_2531);
or UO_79 (O_79,N_2715,N_2731);
and UO_80 (O_80,N_2269,N_2806);
and UO_81 (O_81,N_2768,N_2692);
or UO_82 (O_82,N_2587,N_2270);
nand UO_83 (O_83,N_2398,N_2394);
nand UO_84 (O_84,N_2422,N_2545);
nor UO_85 (O_85,N_2472,N_2457);
nand UO_86 (O_86,N_2553,N_2406);
or UO_87 (O_87,N_2840,N_2813);
or UO_88 (O_88,N_2859,N_2638);
nor UO_89 (O_89,N_2554,N_2973);
nor UO_90 (O_90,N_2591,N_2430);
or UO_91 (O_91,N_2286,N_2879);
nor UO_92 (O_92,N_2774,N_2632);
and UO_93 (O_93,N_2711,N_2397);
nor UO_94 (O_94,N_2528,N_2598);
nand UO_95 (O_95,N_2993,N_2645);
or UO_96 (O_96,N_2581,N_2812);
nand UO_97 (O_97,N_2513,N_2760);
nand UO_98 (O_98,N_2575,N_2777);
or UO_99 (O_99,N_2410,N_2904);
nand UO_100 (O_100,N_2705,N_2467);
nor UO_101 (O_101,N_2926,N_2984);
nor UO_102 (O_102,N_2996,N_2602);
or UO_103 (O_103,N_2435,N_2437);
and UO_104 (O_104,N_2748,N_2673);
and UO_105 (O_105,N_2881,N_2771);
and UO_106 (O_106,N_2382,N_2839);
nand UO_107 (O_107,N_2953,N_2987);
nand UO_108 (O_108,N_2823,N_2562);
nand UO_109 (O_109,N_2256,N_2935);
or UO_110 (O_110,N_2343,N_2274);
nor UO_111 (O_111,N_2696,N_2390);
nand UO_112 (O_112,N_2878,N_2814);
or UO_113 (O_113,N_2713,N_2316);
or UO_114 (O_114,N_2548,N_2648);
or UO_115 (O_115,N_2297,N_2668);
or UO_116 (O_116,N_2348,N_2788);
or UO_117 (O_117,N_2307,N_2379);
or UO_118 (O_118,N_2400,N_2787);
or UO_119 (O_119,N_2707,N_2362);
or UO_120 (O_120,N_2884,N_2723);
or UO_121 (O_121,N_2988,N_2255);
xor UO_122 (O_122,N_2856,N_2483);
or UO_123 (O_123,N_2826,N_2288);
nor UO_124 (O_124,N_2377,N_2913);
nor UO_125 (O_125,N_2273,N_2942);
nand UO_126 (O_126,N_2848,N_2757);
nor UO_127 (O_127,N_2350,N_2477);
or UO_128 (O_128,N_2580,N_2318);
nand UO_129 (O_129,N_2693,N_2268);
or UO_130 (O_130,N_2773,N_2424);
or UO_131 (O_131,N_2599,N_2684);
nand UO_132 (O_132,N_2380,N_2739);
or UO_133 (O_133,N_2595,N_2902);
nor UO_134 (O_134,N_2741,N_2770);
nand UO_135 (O_135,N_2719,N_2679);
or UO_136 (O_136,N_2371,N_2459);
nand UO_137 (O_137,N_2287,N_2660);
nand UO_138 (O_138,N_2434,N_2931);
or UO_139 (O_139,N_2448,N_2570);
nor UO_140 (O_140,N_2420,N_2828);
and UO_141 (O_141,N_2979,N_2793);
nor UO_142 (O_142,N_2396,N_2985);
and UO_143 (O_143,N_2657,N_2945);
nor UO_144 (O_144,N_2617,N_2710);
or UO_145 (O_145,N_2313,N_2498);
and UO_146 (O_146,N_2975,N_2703);
and UO_147 (O_147,N_2809,N_2309);
and UO_148 (O_148,N_2558,N_2758);
nor UO_149 (O_149,N_2670,N_2566);
or UO_150 (O_150,N_2957,N_2466);
or UO_151 (O_151,N_2519,N_2412);
or UO_152 (O_152,N_2607,N_2686);
xnor UO_153 (O_153,N_2861,N_2948);
or UO_154 (O_154,N_2968,N_2962);
or UO_155 (O_155,N_2701,N_2324);
and UO_156 (O_156,N_2322,N_2752);
or UO_157 (O_157,N_2294,N_2683);
and UO_158 (O_158,N_2573,N_2925);
and UO_159 (O_159,N_2363,N_2799);
nand UO_160 (O_160,N_2918,N_2786);
xor UO_161 (O_161,N_2261,N_2296);
and UO_162 (O_162,N_2724,N_2427);
nor UO_163 (O_163,N_2894,N_2503);
or UO_164 (O_164,N_2302,N_2906);
or UO_165 (O_165,N_2970,N_2432);
and UO_166 (O_166,N_2647,N_2821);
nand UO_167 (O_167,N_2688,N_2642);
nor UO_168 (O_168,N_2572,N_2761);
and UO_169 (O_169,N_2818,N_2971);
nand UO_170 (O_170,N_2568,N_2738);
or UO_171 (O_171,N_2305,N_2522);
or UO_172 (O_172,N_2608,N_2300);
and UO_173 (O_173,N_2944,N_2543);
and UO_174 (O_174,N_2555,N_2999);
nand UO_175 (O_175,N_2804,N_2764);
nand UO_176 (O_176,N_2772,N_2308);
and UO_177 (O_177,N_2669,N_2967);
nor UO_178 (O_178,N_2253,N_2659);
and UO_179 (O_179,N_2592,N_2783);
nor UO_180 (O_180,N_2704,N_2494);
nor UO_181 (O_181,N_2747,N_2516);
nor UO_182 (O_182,N_2523,N_2653);
or UO_183 (O_183,N_2830,N_2458);
and UO_184 (O_184,N_2615,N_2867);
nor UO_185 (O_185,N_2560,N_2927);
nor UO_186 (O_186,N_2829,N_2456);
nand UO_187 (O_187,N_2585,N_2920);
nand UO_188 (O_188,N_2890,N_2441);
and UO_189 (O_189,N_2845,N_2797);
nand UO_190 (O_190,N_2557,N_2323);
nand UO_191 (O_191,N_2507,N_2292);
and UO_192 (O_192,N_2853,N_2340);
nand UO_193 (O_193,N_2982,N_2373);
and UO_194 (O_194,N_2792,N_2737);
nand UO_195 (O_195,N_2986,N_2493);
or UO_196 (O_196,N_2750,N_2998);
and UO_197 (O_197,N_2807,N_2547);
nor UO_198 (O_198,N_2718,N_2453);
nand UO_199 (O_199,N_2983,N_2551);
or UO_200 (O_200,N_2621,N_2699);
nand UO_201 (O_201,N_2462,N_2636);
nand UO_202 (O_202,N_2279,N_2663);
nand UO_203 (O_203,N_2440,N_2298);
nand UO_204 (O_204,N_2672,N_2624);
nand UO_205 (O_205,N_2702,N_2841);
and UO_206 (O_206,N_2546,N_2433);
nand UO_207 (O_207,N_2781,N_2940);
or UO_208 (O_208,N_2616,N_2314);
nand UO_209 (O_209,N_2550,N_2949);
nor UO_210 (O_210,N_2312,N_2698);
or UO_211 (O_211,N_2665,N_2974);
nor UO_212 (O_212,N_2691,N_2589);
or UO_213 (O_213,N_2416,N_2351);
and UO_214 (O_214,N_2992,N_2870);
xor UO_215 (O_215,N_2626,N_2497);
nor UO_216 (O_216,N_2835,N_2685);
nor UO_217 (O_217,N_2910,N_2414);
nor UO_218 (O_218,N_2484,N_2335);
nor UO_219 (O_219,N_2488,N_2929);
nand UO_220 (O_220,N_2368,N_2413);
and UO_221 (O_221,N_2893,N_2619);
or UO_222 (O_222,N_2790,N_2864);
nor UO_223 (O_223,N_2597,N_2536);
nor UO_224 (O_224,N_2524,N_2733);
xnor UO_225 (O_225,N_2502,N_2532);
nor UO_226 (O_226,N_2745,N_2342);
or UO_227 (O_227,N_2563,N_2478);
or UO_228 (O_228,N_2837,N_2969);
or UO_229 (O_229,N_2832,N_2344);
nand UO_230 (O_230,N_2883,N_2574);
nand UO_231 (O_231,N_2916,N_2606);
and UO_232 (O_232,N_2922,N_2364);
and UO_233 (O_233,N_2795,N_2978);
or UO_234 (O_234,N_2947,N_2631);
or UO_235 (O_235,N_2742,N_2909);
nand UO_236 (O_236,N_2473,N_2796);
nand UO_237 (O_237,N_2552,N_2869);
and UO_238 (O_238,N_2954,N_2939);
and UO_239 (O_239,N_2655,N_2820);
and UO_240 (O_240,N_2889,N_2541);
and UO_241 (O_241,N_2544,N_2411);
and UO_242 (O_242,N_2612,N_2899);
nand UO_243 (O_243,N_2896,N_2346);
nor UO_244 (O_244,N_2766,N_2431);
nor UO_245 (O_245,N_2754,N_2930);
nor UO_246 (O_246,N_2778,N_2381);
and UO_247 (O_247,N_2360,N_2720);
or UO_248 (O_248,N_2326,N_2439);
and UO_249 (O_249,N_2900,N_2923);
nor UO_250 (O_250,N_2641,N_2914);
nand UO_251 (O_251,N_2384,N_2656);
nor UO_252 (O_252,N_2317,N_2404);
or UO_253 (O_253,N_2361,N_2649);
or UO_254 (O_254,N_2762,N_2875);
nor UO_255 (O_255,N_2556,N_2444);
xnor UO_256 (O_256,N_2370,N_2311);
and UO_257 (O_257,N_2378,N_2611);
nor UO_258 (O_258,N_2263,N_2325);
nand UO_259 (O_259,N_2675,N_2419);
and UO_260 (O_260,N_2250,N_2965);
and UO_261 (O_261,N_2321,N_2500);
nand UO_262 (O_262,N_2860,N_2508);
nor UO_263 (O_263,N_2932,N_2629);
nor UO_264 (O_264,N_2266,N_2846);
nand UO_265 (O_265,N_2736,N_2676);
and UO_266 (O_266,N_2357,N_2802);
and UO_267 (O_267,N_2603,N_2582);
nor UO_268 (O_268,N_2586,N_2960);
nor UO_269 (O_269,N_2445,N_2514);
and UO_270 (O_270,N_2627,N_2569);
or UO_271 (O_271,N_2252,N_2779);
and UO_272 (O_272,N_2601,N_2623);
and UO_273 (O_273,N_2271,N_2919);
nand UO_274 (O_274,N_2646,N_2800);
xnor UO_275 (O_275,N_2511,N_2690);
nand UO_276 (O_276,N_2989,N_2977);
nand UO_277 (O_277,N_2391,N_2805);
and UO_278 (O_278,N_2259,N_2620);
and UO_279 (O_279,N_2725,N_2789);
and UO_280 (O_280,N_2680,N_2682);
nor UO_281 (O_281,N_2449,N_2822);
and UO_282 (O_282,N_2990,N_2858);
and UO_283 (O_283,N_2609,N_2451);
or UO_284 (O_284,N_2658,N_2530);
nand UO_285 (O_285,N_2767,N_2785);
nand UO_286 (O_286,N_2936,N_2765);
or UO_287 (O_287,N_2393,N_2650);
nand UO_288 (O_288,N_2277,N_2755);
nand UO_289 (O_289,N_2898,N_2697);
and UO_290 (O_290,N_2358,N_2369);
and UO_291 (O_291,N_2265,N_2564);
nand UO_292 (O_292,N_2505,N_2759);
nand UO_293 (O_293,N_2290,N_2844);
nand UO_294 (O_294,N_2284,N_2775);
nor UO_295 (O_295,N_2464,N_2604);
and UO_296 (O_296,N_2588,N_2593);
or UO_297 (O_297,N_2468,N_2465);
or UO_298 (O_298,N_2877,N_2283);
or UO_299 (O_299,N_2506,N_2876);
or UO_300 (O_300,N_2625,N_2319);
nand UO_301 (O_301,N_2388,N_2289);
nand UO_302 (O_302,N_2652,N_2374);
and UO_303 (O_303,N_2855,N_2865);
nand UO_304 (O_304,N_2946,N_2409);
nand UO_305 (O_305,N_2366,N_2436);
and UO_306 (O_306,N_2561,N_2495);
nor UO_307 (O_307,N_2887,N_2753);
nand UO_308 (O_308,N_2479,N_2405);
or UO_309 (O_309,N_2421,N_2817);
or UO_310 (O_310,N_2743,N_2955);
and UO_311 (O_311,N_2959,N_2345);
nand UO_312 (O_312,N_2501,N_2474);
or UO_313 (O_313,N_2966,N_2584);
nand UO_314 (O_314,N_2367,N_2310);
or UO_315 (O_315,N_2295,N_2952);
nor UO_316 (O_316,N_2485,N_2518);
nand UO_317 (O_317,N_2583,N_2372);
nor UO_318 (O_318,N_2443,N_2637);
nor UO_319 (O_319,N_2499,N_2463);
nand UO_320 (O_320,N_2482,N_2526);
and UO_321 (O_321,N_2426,N_2912);
nand UO_322 (O_322,N_2596,N_2633);
or UO_323 (O_323,N_2428,N_2470);
nor UO_324 (O_324,N_2928,N_2491);
nand UO_325 (O_325,N_2834,N_2905);
nor UO_326 (O_326,N_2880,N_2383);
and UO_327 (O_327,N_2365,N_2282);
nor UO_328 (O_328,N_2871,N_2254);
nor UO_329 (O_329,N_2963,N_2831);
and UO_330 (O_330,N_2794,N_2666);
xor UO_331 (O_331,N_2847,N_2694);
or UO_332 (O_332,N_2540,N_2857);
nor UO_333 (O_333,N_2336,N_2476);
or UO_334 (O_334,N_2512,N_2854);
nand UO_335 (O_335,N_2903,N_2515);
nand UO_336 (O_336,N_2872,N_2687);
nor UO_337 (O_337,N_2721,N_2951);
or UO_338 (O_338,N_2746,N_2535);
nor UO_339 (O_339,N_2480,N_2895);
or UO_340 (O_340,N_2819,N_2613);
or UO_341 (O_341,N_2681,N_2886);
or UO_342 (O_342,N_2917,N_2257);
nand UO_343 (O_343,N_2492,N_2937);
or UO_344 (O_344,N_2446,N_2454);
and UO_345 (O_345,N_2976,N_2728);
and UO_346 (O_346,N_2964,N_2740);
or UO_347 (O_347,N_2389,N_2272);
nor UO_348 (O_348,N_2776,N_2285);
nand UO_349 (O_349,N_2258,N_2455);
nor UO_350 (O_350,N_2815,N_2539);
xor UO_351 (O_351,N_2402,N_2355);
and UO_352 (O_352,N_2708,N_2618);
nand UO_353 (O_353,N_2331,N_2549);
xor UO_354 (O_354,N_2744,N_2811);
nand UO_355 (O_355,N_2991,N_2810);
nand UO_356 (O_356,N_2520,N_2706);
or UO_357 (O_357,N_2447,N_2941);
nor UO_358 (O_358,N_2808,N_2527);
nand UO_359 (O_359,N_2735,N_2264);
or UO_360 (O_360,N_2329,N_2341);
nor UO_361 (O_361,N_2803,N_2299);
or UO_362 (O_362,N_2763,N_2722);
or UO_363 (O_363,N_2509,N_2824);
nand UO_364 (O_364,N_2924,N_2851);
nand UO_365 (O_365,N_2836,N_2678);
or UO_366 (O_366,N_2534,N_2278);
and UO_367 (O_367,N_2262,N_2452);
and UO_368 (O_368,N_2537,N_2576);
nand UO_369 (O_369,N_2863,N_2921);
nand UO_370 (O_370,N_2352,N_2330);
nor UO_371 (O_371,N_2579,N_2280);
or UO_372 (O_372,N_2907,N_2749);
nor UO_373 (O_373,N_2915,N_2359);
or UO_374 (O_374,N_2950,N_2486);
or UO_375 (O_375,N_2606,N_2555);
or UO_376 (O_376,N_2853,N_2670);
nor UO_377 (O_377,N_2799,N_2401);
nor UO_378 (O_378,N_2523,N_2691);
nand UO_379 (O_379,N_2268,N_2475);
or UO_380 (O_380,N_2732,N_2983);
or UO_381 (O_381,N_2338,N_2596);
nand UO_382 (O_382,N_2612,N_2429);
xor UO_383 (O_383,N_2712,N_2342);
or UO_384 (O_384,N_2352,N_2687);
nand UO_385 (O_385,N_2575,N_2546);
and UO_386 (O_386,N_2288,N_2901);
xor UO_387 (O_387,N_2298,N_2461);
and UO_388 (O_388,N_2270,N_2693);
nor UO_389 (O_389,N_2426,N_2838);
nor UO_390 (O_390,N_2702,N_2408);
or UO_391 (O_391,N_2876,N_2728);
nand UO_392 (O_392,N_2437,N_2773);
and UO_393 (O_393,N_2308,N_2791);
and UO_394 (O_394,N_2612,N_2621);
nor UO_395 (O_395,N_2625,N_2669);
and UO_396 (O_396,N_2677,N_2770);
or UO_397 (O_397,N_2505,N_2826);
nand UO_398 (O_398,N_2505,N_2655);
nor UO_399 (O_399,N_2254,N_2701);
nand UO_400 (O_400,N_2465,N_2902);
or UO_401 (O_401,N_2665,N_2583);
and UO_402 (O_402,N_2689,N_2909);
nand UO_403 (O_403,N_2625,N_2460);
nor UO_404 (O_404,N_2954,N_2633);
or UO_405 (O_405,N_2330,N_2627);
xor UO_406 (O_406,N_2828,N_2401);
nor UO_407 (O_407,N_2311,N_2827);
nand UO_408 (O_408,N_2744,N_2835);
and UO_409 (O_409,N_2509,N_2736);
and UO_410 (O_410,N_2554,N_2780);
nor UO_411 (O_411,N_2703,N_2470);
or UO_412 (O_412,N_2391,N_2903);
nand UO_413 (O_413,N_2277,N_2865);
nand UO_414 (O_414,N_2531,N_2586);
and UO_415 (O_415,N_2536,N_2442);
nor UO_416 (O_416,N_2887,N_2362);
or UO_417 (O_417,N_2258,N_2498);
nor UO_418 (O_418,N_2671,N_2927);
nor UO_419 (O_419,N_2484,N_2608);
nand UO_420 (O_420,N_2332,N_2736);
nand UO_421 (O_421,N_2662,N_2641);
and UO_422 (O_422,N_2602,N_2349);
nand UO_423 (O_423,N_2986,N_2587);
or UO_424 (O_424,N_2457,N_2749);
and UO_425 (O_425,N_2807,N_2379);
nand UO_426 (O_426,N_2804,N_2595);
xor UO_427 (O_427,N_2885,N_2285);
nor UO_428 (O_428,N_2340,N_2818);
and UO_429 (O_429,N_2641,N_2456);
nor UO_430 (O_430,N_2998,N_2485);
nor UO_431 (O_431,N_2806,N_2690);
xor UO_432 (O_432,N_2971,N_2503);
or UO_433 (O_433,N_2565,N_2768);
nand UO_434 (O_434,N_2676,N_2666);
or UO_435 (O_435,N_2460,N_2810);
nor UO_436 (O_436,N_2736,N_2886);
and UO_437 (O_437,N_2866,N_2755);
or UO_438 (O_438,N_2363,N_2681);
and UO_439 (O_439,N_2642,N_2991);
nor UO_440 (O_440,N_2415,N_2721);
nand UO_441 (O_441,N_2737,N_2445);
and UO_442 (O_442,N_2324,N_2863);
and UO_443 (O_443,N_2264,N_2704);
and UO_444 (O_444,N_2783,N_2525);
or UO_445 (O_445,N_2629,N_2319);
or UO_446 (O_446,N_2823,N_2774);
nand UO_447 (O_447,N_2392,N_2740);
nand UO_448 (O_448,N_2972,N_2422);
nor UO_449 (O_449,N_2911,N_2988);
and UO_450 (O_450,N_2505,N_2548);
nand UO_451 (O_451,N_2438,N_2672);
or UO_452 (O_452,N_2948,N_2455);
or UO_453 (O_453,N_2478,N_2770);
and UO_454 (O_454,N_2626,N_2654);
nor UO_455 (O_455,N_2755,N_2506);
xor UO_456 (O_456,N_2370,N_2889);
nand UO_457 (O_457,N_2864,N_2688);
and UO_458 (O_458,N_2349,N_2639);
nand UO_459 (O_459,N_2720,N_2282);
xnor UO_460 (O_460,N_2919,N_2424);
or UO_461 (O_461,N_2677,N_2782);
or UO_462 (O_462,N_2581,N_2663);
nor UO_463 (O_463,N_2374,N_2598);
nand UO_464 (O_464,N_2555,N_2369);
or UO_465 (O_465,N_2991,N_2297);
or UO_466 (O_466,N_2534,N_2274);
nand UO_467 (O_467,N_2588,N_2898);
nand UO_468 (O_468,N_2485,N_2856);
nand UO_469 (O_469,N_2732,N_2788);
nor UO_470 (O_470,N_2990,N_2403);
nand UO_471 (O_471,N_2300,N_2293);
nand UO_472 (O_472,N_2876,N_2723);
and UO_473 (O_473,N_2596,N_2279);
nor UO_474 (O_474,N_2966,N_2304);
nand UO_475 (O_475,N_2759,N_2436);
nand UO_476 (O_476,N_2798,N_2565);
nand UO_477 (O_477,N_2970,N_2285);
and UO_478 (O_478,N_2350,N_2418);
or UO_479 (O_479,N_2756,N_2548);
nor UO_480 (O_480,N_2484,N_2556);
nor UO_481 (O_481,N_2491,N_2356);
and UO_482 (O_482,N_2667,N_2745);
nor UO_483 (O_483,N_2272,N_2860);
or UO_484 (O_484,N_2540,N_2954);
nor UO_485 (O_485,N_2761,N_2667);
or UO_486 (O_486,N_2501,N_2718);
nand UO_487 (O_487,N_2312,N_2413);
or UO_488 (O_488,N_2447,N_2369);
nand UO_489 (O_489,N_2304,N_2712);
nand UO_490 (O_490,N_2419,N_2673);
and UO_491 (O_491,N_2524,N_2587);
or UO_492 (O_492,N_2440,N_2902);
nor UO_493 (O_493,N_2714,N_2672);
or UO_494 (O_494,N_2311,N_2632);
or UO_495 (O_495,N_2508,N_2611);
and UO_496 (O_496,N_2770,N_2347);
nand UO_497 (O_497,N_2955,N_2900);
or UO_498 (O_498,N_2483,N_2377);
nor UO_499 (O_499,N_2339,N_2891);
endmodule