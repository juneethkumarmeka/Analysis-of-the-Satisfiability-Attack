module basic_500_3000_500_3_levels_1xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_467,In_436);
nand U1 (N_1,In_236,In_67);
and U2 (N_2,In_109,In_128);
and U3 (N_3,In_16,In_246);
nand U4 (N_4,In_313,In_85);
or U5 (N_5,In_361,In_166);
nand U6 (N_6,In_421,In_244);
nor U7 (N_7,In_420,In_154);
or U8 (N_8,In_305,In_115);
or U9 (N_9,In_229,In_188);
and U10 (N_10,In_435,In_287);
nand U11 (N_11,In_369,In_151);
nor U12 (N_12,In_382,In_482);
and U13 (N_13,In_400,In_279);
and U14 (N_14,In_268,In_402);
nand U15 (N_15,In_104,In_23);
and U16 (N_16,In_392,In_479);
and U17 (N_17,In_300,In_350);
nor U18 (N_18,In_391,In_167);
nor U19 (N_19,In_256,In_240);
nor U20 (N_20,In_405,In_404);
nand U21 (N_21,In_301,In_428);
nand U22 (N_22,In_238,In_71);
and U23 (N_23,In_239,In_314);
and U24 (N_24,In_157,In_178);
nor U25 (N_25,In_267,In_231);
or U26 (N_26,In_389,In_53);
or U27 (N_27,In_211,In_273);
or U28 (N_28,In_378,In_70);
or U29 (N_29,In_9,In_312);
and U30 (N_30,In_164,In_2);
nor U31 (N_31,In_270,In_72);
nor U32 (N_32,In_106,In_340);
nor U33 (N_33,In_19,In_440);
or U34 (N_34,In_200,In_38);
nor U35 (N_35,In_387,In_245);
and U36 (N_36,In_176,In_429);
and U37 (N_37,In_186,In_39);
nand U38 (N_38,In_281,In_218);
and U39 (N_39,In_373,In_439);
and U40 (N_40,In_105,In_148);
or U41 (N_41,In_263,In_484);
nor U42 (N_42,In_49,In_78);
nand U43 (N_43,In_189,In_32);
and U44 (N_44,In_469,In_321);
or U45 (N_45,In_422,In_496);
or U46 (N_46,In_202,In_475);
nand U47 (N_47,In_185,In_88);
nor U48 (N_48,In_356,In_410);
nand U49 (N_49,In_360,In_359);
or U50 (N_50,In_187,In_180);
nand U51 (N_51,In_155,In_223);
nand U52 (N_52,In_205,In_36);
or U53 (N_53,In_61,In_383);
and U54 (N_54,In_81,In_96);
and U55 (N_55,In_393,In_217);
and U56 (N_56,In_12,In_437);
and U57 (N_57,In_492,In_499);
nor U58 (N_58,In_83,In_194);
and U59 (N_59,In_354,In_374);
or U60 (N_60,In_262,In_325);
or U61 (N_61,In_311,In_25);
and U62 (N_62,In_193,In_214);
nand U63 (N_63,In_206,In_134);
nor U64 (N_64,In_444,In_460);
nor U65 (N_65,In_168,In_427);
or U66 (N_66,In_198,In_355);
or U67 (N_67,In_441,In_65);
or U68 (N_68,In_418,In_261);
nand U69 (N_69,In_250,In_304);
or U70 (N_70,In_465,In_485);
nor U71 (N_71,In_282,In_170);
and U72 (N_72,In_116,In_107);
and U73 (N_73,In_323,In_99);
nand U74 (N_74,In_425,In_35);
nor U75 (N_75,In_183,In_114);
or U76 (N_76,In_409,In_137);
or U77 (N_77,In_288,In_324);
nand U78 (N_78,In_34,In_278);
nor U79 (N_79,In_433,In_364);
nor U80 (N_80,In_181,In_121);
or U81 (N_81,In_210,In_341);
and U82 (N_82,In_481,In_289);
nor U83 (N_83,In_495,In_269);
nand U84 (N_84,In_111,In_251);
or U85 (N_85,In_252,In_87);
or U86 (N_86,In_266,In_451);
or U87 (N_87,In_464,In_209);
nand U88 (N_88,In_489,In_490);
nor U89 (N_89,In_345,In_468);
nor U90 (N_90,In_342,In_126);
or U91 (N_91,In_259,In_358);
and U92 (N_92,In_172,In_57);
or U93 (N_93,In_29,In_58);
nand U94 (N_94,In_8,In_296);
nor U95 (N_95,In_474,In_20);
nand U96 (N_96,In_13,In_320);
or U97 (N_97,In_381,In_21);
nand U98 (N_98,In_276,In_163);
or U99 (N_99,In_362,In_280);
nand U100 (N_100,In_130,In_286);
or U101 (N_101,In_349,In_412);
or U102 (N_102,In_367,In_227);
or U103 (N_103,In_17,In_318);
or U104 (N_104,In_461,In_327);
nand U105 (N_105,In_366,In_123);
or U106 (N_106,In_315,In_306);
or U107 (N_107,In_284,In_64);
nor U108 (N_108,In_331,In_442);
or U109 (N_109,In_316,In_234);
and U110 (N_110,In_42,In_396);
or U111 (N_111,In_283,In_415);
nand U112 (N_112,In_368,In_86);
nor U113 (N_113,In_470,In_473);
nor U114 (N_114,In_132,In_445);
nand U115 (N_115,In_184,In_119);
or U116 (N_116,In_28,In_277);
nand U117 (N_117,In_149,In_357);
nor U118 (N_118,In_307,In_326);
and U119 (N_119,In_122,In_162);
nor U120 (N_120,In_254,In_472);
and U121 (N_121,In_448,In_7);
or U122 (N_122,In_253,In_417);
and U123 (N_123,In_450,In_295);
nand U124 (N_124,In_161,In_182);
and U125 (N_125,In_69,In_299);
and U126 (N_126,In_80,In_447);
and U127 (N_127,In_139,In_483);
and U128 (N_128,In_46,In_55);
nor U129 (N_129,In_466,In_95);
nor U130 (N_130,In_192,In_487);
nor U131 (N_131,In_265,In_379);
nor U132 (N_132,In_297,In_191);
nand U133 (N_133,In_232,In_416);
nor U134 (N_134,In_213,In_332);
nand U135 (N_135,In_177,In_197);
or U136 (N_136,In_335,In_138);
or U137 (N_137,In_249,In_478);
or U138 (N_138,In_174,In_201);
or U139 (N_139,In_76,In_41);
and U140 (N_140,In_219,In_91);
and U141 (N_141,In_411,In_140);
or U142 (N_142,In_131,In_66);
nor U143 (N_143,In_135,In_491);
and U144 (N_144,In_462,In_272);
nor U145 (N_145,In_463,In_363);
nor U146 (N_146,In_169,In_322);
nand U147 (N_147,In_243,In_47);
nor U148 (N_148,In_22,In_408);
nand U149 (N_149,In_113,In_380);
and U150 (N_150,In_255,In_5);
nand U151 (N_151,In_136,In_302);
or U152 (N_152,In_431,In_63);
or U153 (N_153,In_233,In_216);
nor U154 (N_154,In_127,In_260);
nand U155 (N_155,In_175,In_237);
nand U156 (N_156,In_377,In_203);
nand U157 (N_157,In_60,In_446);
nor U158 (N_158,In_212,In_334);
nor U159 (N_159,In_141,In_74);
and U160 (N_160,In_449,In_352);
and U161 (N_161,In_100,In_370);
nor U162 (N_162,In_31,In_292);
nand U163 (N_163,In_56,In_77);
nand U164 (N_164,In_3,In_376);
nor U165 (N_165,In_50,In_424);
and U166 (N_166,In_258,In_480);
or U167 (N_167,In_399,In_48);
or U168 (N_168,In_271,In_24);
nor U169 (N_169,In_10,In_336);
or U170 (N_170,In_458,In_27);
and U171 (N_171,In_26,In_153);
nor U172 (N_172,In_129,In_101);
and U173 (N_173,In_493,In_455);
nand U174 (N_174,In_110,In_147);
nand U175 (N_175,In_330,In_18);
nand U176 (N_176,In_353,In_52);
or U177 (N_177,In_92,In_90);
nor U178 (N_178,In_375,In_434);
or U179 (N_179,In_432,In_40);
nor U180 (N_180,In_30,In_328);
or U181 (N_181,In_208,In_275);
nand U182 (N_182,In_75,In_308);
and U183 (N_183,In_476,In_386);
nand U184 (N_184,In_365,In_257);
nand U185 (N_185,In_426,In_6);
and U186 (N_186,In_303,In_309);
or U187 (N_187,In_14,In_403);
nor U188 (N_188,In_388,In_497);
nor U189 (N_189,In_54,In_459);
and U190 (N_190,In_346,In_108);
nand U191 (N_191,In_339,In_471);
nand U192 (N_192,In_51,In_143);
nor U193 (N_193,In_241,In_125);
nand U194 (N_194,In_419,In_310);
nor U195 (N_195,In_156,In_220);
or U196 (N_196,In_344,In_68);
nor U197 (N_197,In_319,In_150);
nand U198 (N_198,In_222,In_406);
nor U199 (N_199,In_207,In_1);
nor U200 (N_200,In_371,In_199);
nand U201 (N_201,In_413,In_486);
and U202 (N_202,In_242,In_248);
and U203 (N_203,In_372,In_454);
nand U204 (N_204,In_133,In_204);
nand U205 (N_205,In_453,In_225);
and U206 (N_206,In_103,In_230);
and U207 (N_207,In_438,In_158);
nand U208 (N_208,In_494,In_15);
and U209 (N_209,In_73,In_452);
nand U210 (N_210,In_37,In_285);
or U211 (N_211,In_118,In_488);
nor U212 (N_212,In_112,In_290);
nand U213 (N_213,In_457,In_94);
nand U214 (N_214,In_401,In_394);
or U215 (N_215,In_79,In_298);
or U216 (N_216,In_443,In_343);
or U217 (N_217,In_117,In_62);
nand U218 (N_218,In_196,In_351);
nor U219 (N_219,In_385,In_171);
or U220 (N_220,In_190,In_159);
and U221 (N_221,In_93,In_4);
nor U222 (N_222,In_235,In_274);
and U223 (N_223,In_98,In_0);
and U224 (N_224,In_398,In_264);
or U225 (N_225,In_124,In_215);
or U226 (N_226,In_347,In_226);
nand U227 (N_227,In_146,In_152);
nor U228 (N_228,In_173,In_293);
or U229 (N_229,In_317,In_102);
nand U230 (N_230,In_44,In_82);
nor U231 (N_231,In_477,In_120);
nand U232 (N_232,In_160,In_228);
nand U233 (N_233,In_43,In_33);
nor U234 (N_234,In_414,In_329);
and U235 (N_235,In_337,In_395);
nand U236 (N_236,In_338,In_348);
nor U237 (N_237,In_144,In_179);
and U238 (N_238,In_145,In_384);
nor U239 (N_239,In_142,In_221);
and U240 (N_240,In_333,In_498);
nand U241 (N_241,In_224,In_165);
and U242 (N_242,In_247,In_11);
and U243 (N_243,In_89,In_423);
nor U244 (N_244,In_291,In_456);
nand U245 (N_245,In_397,In_294);
nor U246 (N_246,In_59,In_430);
and U247 (N_247,In_45,In_195);
nor U248 (N_248,In_390,In_84);
or U249 (N_249,In_407,In_97);
nand U250 (N_250,In_200,In_183);
and U251 (N_251,In_445,In_165);
or U252 (N_252,In_356,In_39);
or U253 (N_253,In_194,In_399);
nor U254 (N_254,In_406,In_250);
nand U255 (N_255,In_152,In_398);
and U256 (N_256,In_274,In_251);
xnor U257 (N_257,In_428,In_145);
and U258 (N_258,In_69,In_74);
or U259 (N_259,In_317,In_78);
nor U260 (N_260,In_94,In_174);
nor U261 (N_261,In_288,In_294);
and U262 (N_262,In_388,In_28);
or U263 (N_263,In_47,In_335);
or U264 (N_264,In_115,In_100);
nor U265 (N_265,In_300,In_96);
nor U266 (N_266,In_26,In_78);
nor U267 (N_267,In_236,In_465);
or U268 (N_268,In_81,In_291);
nand U269 (N_269,In_161,In_340);
nand U270 (N_270,In_369,In_147);
and U271 (N_271,In_337,In_318);
and U272 (N_272,In_499,In_35);
nand U273 (N_273,In_72,In_90);
or U274 (N_274,In_388,In_482);
nand U275 (N_275,In_171,In_215);
or U276 (N_276,In_346,In_102);
nor U277 (N_277,In_28,In_344);
and U278 (N_278,In_251,In_244);
nor U279 (N_279,In_288,In_252);
and U280 (N_280,In_411,In_233);
nor U281 (N_281,In_2,In_189);
nand U282 (N_282,In_190,In_112);
or U283 (N_283,In_382,In_259);
nand U284 (N_284,In_87,In_497);
and U285 (N_285,In_234,In_101);
or U286 (N_286,In_27,In_313);
or U287 (N_287,In_10,In_177);
or U288 (N_288,In_31,In_263);
and U289 (N_289,In_451,In_10);
nand U290 (N_290,In_22,In_139);
nor U291 (N_291,In_135,In_90);
nor U292 (N_292,In_424,In_311);
nor U293 (N_293,In_182,In_139);
nand U294 (N_294,In_96,In_310);
and U295 (N_295,In_6,In_72);
xor U296 (N_296,In_167,In_192);
or U297 (N_297,In_143,In_284);
or U298 (N_298,In_125,In_455);
nand U299 (N_299,In_139,In_493);
nand U300 (N_300,In_11,In_325);
nand U301 (N_301,In_344,In_91);
and U302 (N_302,In_147,In_431);
nand U303 (N_303,In_218,In_438);
or U304 (N_304,In_70,In_388);
nand U305 (N_305,In_303,In_111);
or U306 (N_306,In_113,In_49);
and U307 (N_307,In_337,In_42);
nand U308 (N_308,In_162,In_328);
nor U309 (N_309,In_175,In_181);
nor U310 (N_310,In_421,In_13);
or U311 (N_311,In_79,In_268);
and U312 (N_312,In_43,In_369);
or U313 (N_313,In_53,In_174);
or U314 (N_314,In_361,In_460);
nor U315 (N_315,In_321,In_419);
nand U316 (N_316,In_201,In_305);
nand U317 (N_317,In_170,In_148);
nor U318 (N_318,In_417,In_136);
nand U319 (N_319,In_332,In_414);
nor U320 (N_320,In_98,In_61);
xnor U321 (N_321,In_136,In_207);
nor U322 (N_322,In_435,In_319);
nand U323 (N_323,In_347,In_494);
or U324 (N_324,In_305,In_224);
or U325 (N_325,In_294,In_65);
nand U326 (N_326,In_373,In_92);
nor U327 (N_327,In_97,In_447);
and U328 (N_328,In_106,In_119);
nor U329 (N_329,In_248,In_285);
or U330 (N_330,In_164,In_477);
or U331 (N_331,In_406,In_243);
and U332 (N_332,In_499,In_480);
xnor U333 (N_333,In_369,In_458);
or U334 (N_334,In_398,In_333);
nand U335 (N_335,In_463,In_322);
nor U336 (N_336,In_149,In_383);
or U337 (N_337,In_445,In_387);
nor U338 (N_338,In_29,In_316);
nor U339 (N_339,In_99,In_133);
nor U340 (N_340,In_251,In_465);
or U341 (N_341,In_54,In_462);
and U342 (N_342,In_456,In_145);
or U343 (N_343,In_137,In_440);
nor U344 (N_344,In_118,In_392);
and U345 (N_345,In_382,In_231);
or U346 (N_346,In_360,In_210);
nand U347 (N_347,In_398,In_149);
nand U348 (N_348,In_153,In_478);
and U349 (N_349,In_69,In_294);
nand U350 (N_350,In_210,In_197);
nor U351 (N_351,In_199,In_251);
and U352 (N_352,In_284,In_93);
and U353 (N_353,In_336,In_255);
or U354 (N_354,In_308,In_427);
and U355 (N_355,In_19,In_368);
and U356 (N_356,In_365,In_139);
and U357 (N_357,In_475,In_399);
nor U358 (N_358,In_23,In_156);
nor U359 (N_359,In_84,In_36);
nor U360 (N_360,In_176,In_230);
and U361 (N_361,In_359,In_343);
and U362 (N_362,In_153,In_341);
or U363 (N_363,In_383,In_83);
and U364 (N_364,In_498,In_384);
and U365 (N_365,In_206,In_337);
and U366 (N_366,In_407,In_473);
nor U367 (N_367,In_212,In_197);
nand U368 (N_368,In_186,In_157);
or U369 (N_369,In_196,In_264);
nor U370 (N_370,In_455,In_190);
nor U371 (N_371,In_91,In_129);
or U372 (N_372,In_63,In_64);
nand U373 (N_373,In_242,In_160);
nor U374 (N_374,In_256,In_67);
nor U375 (N_375,In_257,In_284);
nor U376 (N_376,In_405,In_397);
or U377 (N_377,In_173,In_420);
nand U378 (N_378,In_450,In_269);
and U379 (N_379,In_120,In_405);
nor U380 (N_380,In_381,In_207);
nor U381 (N_381,In_116,In_467);
and U382 (N_382,In_301,In_297);
and U383 (N_383,In_253,In_493);
or U384 (N_384,In_122,In_367);
nor U385 (N_385,In_395,In_309);
or U386 (N_386,In_477,In_230);
and U387 (N_387,In_98,In_262);
nor U388 (N_388,In_273,In_278);
nand U389 (N_389,In_415,In_447);
and U390 (N_390,In_42,In_339);
nand U391 (N_391,In_67,In_384);
nand U392 (N_392,In_407,In_90);
nor U393 (N_393,In_269,In_117);
and U394 (N_394,In_20,In_492);
nor U395 (N_395,In_414,In_93);
or U396 (N_396,In_469,In_477);
nand U397 (N_397,In_337,In_436);
or U398 (N_398,In_43,In_69);
and U399 (N_399,In_172,In_427);
and U400 (N_400,In_312,In_496);
nand U401 (N_401,In_277,In_111);
nor U402 (N_402,In_184,In_227);
or U403 (N_403,In_439,In_294);
or U404 (N_404,In_416,In_316);
nand U405 (N_405,In_409,In_63);
nand U406 (N_406,In_16,In_37);
and U407 (N_407,In_352,In_457);
and U408 (N_408,In_167,In_94);
nor U409 (N_409,In_189,In_194);
or U410 (N_410,In_78,In_330);
or U411 (N_411,In_156,In_188);
or U412 (N_412,In_246,In_45);
xnor U413 (N_413,In_310,In_45);
or U414 (N_414,In_397,In_186);
or U415 (N_415,In_419,In_122);
nand U416 (N_416,In_297,In_351);
or U417 (N_417,In_35,In_18);
and U418 (N_418,In_432,In_23);
xor U419 (N_419,In_143,In_12);
or U420 (N_420,In_458,In_136);
nor U421 (N_421,In_19,In_103);
and U422 (N_422,In_133,In_131);
and U423 (N_423,In_92,In_417);
or U424 (N_424,In_29,In_377);
nand U425 (N_425,In_448,In_302);
nand U426 (N_426,In_94,In_132);
and U427 (N_427,In_48,In_251);
or U428 (N_428,In_37,In_48);
nor U429 (N_429,In_7,In_349);
nand U430 (N_430,In_193,In_199);
or U431 (N_431,In_16,In_394);
and U432 (N_432,In_135,In_94);
nand U433 (N_433,In_474,In_405);
nand U434 (N_434,In_429,In_93);
nor U435 (N_435,In_387,In_228);
nand U436 (N_436,In_301,In_234);
nor U437 (N_437,In_364,In_349);
or U438 (N_438,In_109,In_436);
or U439 (N_439,In_14,In_206);
nor U440 (N_440,In_43,In_480);
nand U441 (N_441,In_262,In_38);
and U442 (N_442,In_256,In_196);
nor U443 (N_443,In_270,In_177);
nand U444 (N_444,In_239,In_361);
or U445 (N_445,In_411,In_302);
nand U446 (N_446,In_433,In_291);
or U447 (N_447,In_93,In_452);
or U448 (N_448,In_155,In_416);
or U449 (N_449,In_428,In_249);
nand U450 (N_450,In_94,In_246);
nand U451 (N_451,In_137,In_252);
or U452 (N_452,In_79,In_230);
or U453 (N_453,In_323,In_406);
and U454 (N_454,In_114,In_432);
nand U455 (N_455,In_414,In_341);
nand U456 (N_456,In_431,In_321);
and U457 (N_457,In_95,In_381);
and U458 (N_458,In_201,In_111);
nor U459 (N_459,In_267,In_108);
nor U460 (N_460,In_227,In_132);
nand U461 (N_461,In_351,In_187);
nand U462 (N_462,In_287,In_116);
nand U463 (N_463,In_281,In_240);
and U464 (N_464,In_365,In_187);
nand U465 (N_465,In_312,In_316);
or U466 (N_466,In_280,In_4);
and U467 (N_467,In_264,In_424);
or U468 (N_468,In_225,In_372);
and U469 (N_469,In_288,In_232);
nor U470 (N_470,In_57,In_165);
nor U471 (N_471,In_344,In_476);
nor U472 (N_472,In_15,In_481);
nand U473 (N_473,In_139,In_246);
nand U474 (N_474,In_12,In_145);
nor U475 (N_475,In_394,In_61);
and U476 (N_476,In_281,In_67);
nor U477 (N_477,In_78,In_455);
nand U478 (N_478,In_193,In_447);
and U479 (N_479,In_133,In_173);
nor U480 (N_480,In_112,In_54);
nor U481 (N_481,In_305,In_270);
and U482 (N_482,In_152,In_207);
and U483 (N_483,In_436,In_58);
nand U484 (N_484,In_184,In_33);
nand U485 (N_485,In_76,In_255);
nor U486 (N_486,In_44,In_378);
and U487 (N_487,In_279,In_277);
or U488 (N_488,In_149,In_354);
or U489 (N_489,In_64,In_123);
or U490 (N_490,In_118,In_482);
or U491 (N_491,In_239,In_251);
and U492 (N_492,In_2,In_38);
and U493 (N_493,In_314,In_320);
nor U494 (N_494,In_457,In_475);
or U495 (N_495,In_400,In_441);
nor U496 (N_496,In_349,In_63);
and U497 (N_497,In_183,In_283);
nand U498 (N_498,In_136,In_445);
nor U499 (N_499,In_31,In_466);
nand U500 (N_500,In_159,In_470);
and U501 (N_501,In_19,In_4);
nand U502 (N_502,In_214,In_44);
and U503 (N_503,In_320,In_46);
nor U504 (N_504,In_9,In_280);
nor U505 (N_505,In_373,In_280);
or U506 (N_506,In_494,In_495);
or U507 (N_507,In_202,In_225);
nor U508 (N_508,In_264,In_484);
or U509 (N_509,In_146,In_289);
nand U510 (N_510,In_97,In_184);
nor U511 (N_511,In_89,In_382);
and U512 (N_512,In_79,In_378);
nor U513 (N_513,In_357,In_182);
and U514 (N_514,In_219,In_208);
nor U515 (N_515,In_481,In_338);
or U516 (N_516,In_152,In_233);
nor U517 (N_517,In_62,In_288);
or U518 (N_518,In_485,In_296);
nor U519 (N_519,In_294,In_252);
or U520 (N_520,In_28,In_495);
or U521 (N_521,In_139,In_215);
nor U522 (N_522,In_110,In_451);
nand U523 (N_523,In_405,In_43);
nor U524 (N_524,In_395,In_85);
nor U525 (N_525,In_308,In_416);
and U526 (N_526,In_77,In_398);
or U527 (N_527,In_321,In_191);
xnor U528 (N_528,In_318,In_259);
nand U529 (N_529,In_134,In_101);
and U530 (N_530,In_455,In_47);
or U531 (N_531,In_283,In_82);
nor U532 (N_532,In_74,In_275);
nand U533 (N_533,In_53,In_259);
or U534 (N_534,In_56,In_115);
or U535 (N_535,In_256,In_8);
nor U536 (N_536,In_289,In_242);
nor U537 (N_537,In_59,In_165);
nor U538 (N_538,In_94,In_270);
nand U539 (N_539,In_399,In_430);
and U540 (N_540,In_225,In_110);
nor U541 (N_541,In_234,In_42);
or U542 (N_542,In_282,In_1);
and U543 (N_543,In_171,In_491);
nor U544 (N_544,In_109,In_112);
nor U545 (N_545,In_366,In_178);
xnor U546 (N_546,In_322,In_49);
xnor U547 (N_547,In_75,In_361);
or U548 (N_548,In_415,In_190);
and U549 (N_549,In_274,In_469);
or U550 (N_550,In_27,In_87);
and U551 (N_551,In_206,In_379);
and U552 (N_552,In_254,In_328);
nor U553 (N_553,In_303,In_47);
nor U554 (N_554,In_340,In_253);
xnor U555 (N_555,In_144,In_241);
or U556 (N_556,In_307,In_329);
nand U557 (N_557,In_166,In_381);
or U558 (N_558,In_0,In_466);
or U559 (N_559,In_101,In_392);
nand U560 (N_560,In_303,In_274);
nand U561 (N_561,In_172,In_456);
nor U562 (N_562,In_401,In_471);
nor U563 (N_563,In_125,In_142);
nand U564 (N_564,In_133,In_388);
or U565 (N_565,In_10,In_174);
and U566 (N_566,In_318,In_49);
and U567 (N_567,In_25,In_82);
nand U568 (N_568,In_490,In_213);
nor U569 (N_569,In_462,In_344);
or U570 (N_570,In_372,In_360);
nand U571 (N_571,In_260,In_164);
or U572 (N_572,In_491,In_391);
nor U573 (N_573,In_207,In_61);
nor U574 (N_574,In_149,In_195);
nor U575 (N_575,In_400,In_56);
nand U576 (N_576,In_124,In_171);
and U577 (N_577,In_81,In_121);
and U578 (N_578,In_368,In_133);
nor U579 (N_579,In_464,In_460);
nor U580 (N_580,In_367,In_138);
or U581 (N_581,In_454,In_391);
or U582 (N_582,In_182,In_305);
or U583 (N_583,In_401,In_305);
nor U584 (N_584,In_96,In_106);
nor U585 (N_585,In_269,In_220);
or U586 (N_586,In_407,In_67);
nor U587 (N_587,In_362,In_252);
nand U588 (N_588,In_474,In_160);
nand U589 (N_589,In_281,In_180);
or U590 (N_590,In_269,In_389);
or U591 (N_591,In_37,In_44);
or U592 (N_592,In_284,In_10);
nor U593 (N_593,In_334,In_327);
and U594 (N_594,In_262,In_452);
nand U595 (N_595,In_77,In_90);
nand U596 (N_596,In_141,In_68);
or U597 (N_597,In_428,In_239);
or U598 (N_598,In_246,In_313);
nor U599 (N_599,In_109,In_479);
nor U600 (N_600,In_31,In_29);
and U601 (N_601,In_285,In_475);
nor U602 (N_602,In_16,In_53);
nor U603 (N_603,In_499,In_193);
nor U604 (N_604,In_461,In_49);
nand U605 (N_605,In_442,In_148);
nand U606 (N_606,In_140,In_42);
nor U607 (N_607,In_210,In_249);
and U608 (N_608,In_149,In_51);
or U609 (N_609,In_365,In_90);
xor U610 (N_610,In_117,In_148);
nand U611 (N_611,In_194,In_96);
nand U612 (N_612,In_188,In_298);
and U613 (N_613,In_67,In_264);
nor U614 (N_614,In_43,In_470);
nor U615 (N_615,In_29,In_275);
or U616 (N_616,In_83,In_347);
and U617 (N_617,In_149,In_110);
nand U618 (N_618,In_114,In_100);
and U619 (N_619,In_478,In_389);
or U620 (N_620,In_208,In_268);
or U621 (N_621,In_357,In_360);
nand U622 (N_622,In_123,In_432);
and U623 (N_623,In_253,In_88);
nand U624 (N_624,In_350,In_148);
and U625 (N_625,In_328,In_272);
or U626 (N_626,In_138,In_337);
and U627 (N_627,In_160,In_60);
and U628 (N_628,In_430,In_95);
or U629 (N_629,In_470,In_476);
nand U630 (N_630,In_350,In_485);
or U631 (N_631,In_88,In_487);
or U632 (N_632,In_492,In_21);
or U633 (N_633,In_420,In_364);
or U634 (N_634,In_19,In_68);
and U635 (N_635,In_469,In_284);
nand U636 (N_636,In_198,In_301);
nor U637 (N_637,In_388,In_315);
nor U638 (N_638,In_162,In_355);
or U639 (N_639,In_273,In_293);
nand U640 (N_640,In_25,In_105);
nand U641 (N_641,In_267,In_368);
and U642 (N_642,In_77,In_220);
nor U643 (N_643,In_98,In_229);
and U644 (N_644,In_468,In_64);
and U645 (N_645,In_268,In_374);
or U646 (N_646,In_184,In_139);
nand U647 (N_647,In_85,In_315);
nor U648 (N_648,In_283,In_195);
and U649 (N_649,In_259,In_119);
nor U650 (N_650,In_356,In_349);
or U651 (N_651,In_143,In_7);
or U652 (N_652,In_37,In_8);
or U653 (N_653,In_187,In_322);
or U654 (N_654,In_283,In_368);
and U655 (N_655,In_180,In_243);
or U656 (N_656,In_101,In_253);
and U657 (N_657,In_4,In_433);
and U658 (N_658,In_325,In_276);
nor U659 (N_659,In_76,In_206);
nand U660 (N_660,In_345,In_16);
nand U661 (N_661,In_438,In_55);
nand U662 (N_662,In_457,In_317);
or U663 (N_663,In_463,In_3);
and U664 (N_664,In_392,In_3);
and U665 (N_665,In_315,In_253);
and U666 (N_666,In_327,In_152);
nor U667 (N_667,In_240,In_372);
nor U668 (N_668,In_300,In_218);
and U669 (N_669,In_237,In_288);
or U670 (N_670,In_194,In_462);
nor U671 (N_671,In_115,In_41);
nand U672 (N_672,In_273,In_169);
and U673 (N_673,In_499,In_311);
nor U674 (N_674,In_482,In_39);
and U675 (N_675,In_310,In_459);
nand U676 (N_676,In_157,In_214);
nor U677 (N_677,In_478,In_73);
nand U678 (N_678,In_257,In_225);
nand U679 (N_679,In_167,In_483);
and U680 (N_680,In_315,In_157);
nand U681 (N_681,In_211,In_430);
and U682 (N_682,In_324,In_473);
and U683 (N_683,In_13,In_91);
or U684 (N_684,In_161,In_262);
nor U685 (N_685,In_295,In_470);
nand U686 (N_686,In_171,In_157);
and U687 (N_687,In_165,In_243);
nand U688 (N_688,In_83,In_11);
or U689 (N_689,In_315,In_136);
nor U690 (N_690,In_141,In_278);
nor U691 (N_691,In_392,In_400);
xor U692 (N_692,In_324,In_127);
nand U693 (N_693,In_180,In_312);
nor U694 (N_694,In_34,In_280);
and U695 (N_695,In_373,In_310);
nand U696 (N_696,In_135,In_383);
nor U697 (N_697,In_386,In_266);
nor U698 (N_698,In_124,In_221);
or U699 (N_699,In_285,In_136);
nand U700 (N_700,In_84,In_315);
nand U701 (N_701,In_442,In_102);
and U702 (N_702,In_196,In_2);
nor U703 (N_703,In_0,In_227);
nand U704 (N_704,In_394,In_62);
or U705 (N_705,In_39,In_353);
or U706 (N_706,In_58,In_11);
and U707 (N_707,In_178,In_378);
or U708 (N_708,In_219,In_267);
nand U709 (N_709,In_290,In_5);
nor U710 (N_710,In_157,In_458);
nor U711 (N_711,In_482,In_487);
or U712 (N_712,In_49,In_141);
and U713 (N_713,In_217,In_468);
nand U714 (N_714,In_228,In_203);
or U715 (N_715,In_222,In_94);
and U716 (N_716,In_318,In_86);
and U717 (N_717,In_138,In_415);
or U718 (N_718,In_50,In_498);
nand U719 (N_719,In_376,In_90);
nor U720 (N_720,In_426,In_422);
or U721 (N_721,In_132,In_71);
nor U722 (N_722,In_442,In_313);
and U723 (N_723,In_308,In_78);
nor U724 (N_724,In_208,In_34);
and U725 (N_725,In_378,In_60);
or U726 (N_726,In_89,In_352);
nor U727 (N_727,In_376,In_84);
and U728 (N_728,In_169,In_29);
or U729 (N_729,In_318,In_419);
nor U730 (N_730,In_49,In_28);
or U731 (N_731,In_314,In_493);
nor U732 (N_732,In_3,In_225);
nor U733 (N_733,In_247,In_176);
and U734 (N_734,In_112,In_363);
nand U735 (N_735,In_212,In_105);
nor U736 (N_736,In_290,In_44);
nor U737 (N_737,In_274,In_357);
and U738 (N_738,In_164,In_114);
nor U739 (N_739,In_223,In_340);
or U740 (N_740,In_443,In_300);
nand U741 (N_741,In_226,In_336);
nor U742 (N_742,In_166,In_319);
nor U743 (N_743,In_142,In_207);
and U744 (N_744,In_10,In_490);
and U745 (N_745,In_22,In_312);
nand U746 (N_746,In_172,In_155);
or U747 (N_747,In_152,In_494);
xnor U748 (N_748,In_352,In_450);
nand U749 (N_749,In_254,In_145);
nor U750 (N_750,In_358,In_159);
or U751 (N_751,In_317,In_420);
nand U752 (N_752,In_325,In_154);
or U753 (N_753,In_169,In_241);
nand U754 (N_754,In_30,In_97);
or U755 (N_755,In_53,In_38);
xnor U756 (N_756,In_227,In_450);
or U757 (N_757,In_276,In_448);
and U758 (N_758,In_343,In_31);
nor U759 (N_759,In_367,In_330);
nor U760 (N_760,In_222,In_491);
nand U761 (N_761,In_429,In_431);
and U762 (N_762,In_475,In_130);
nand U763 (N_763,In_156,In_357);
nand U764 (N_764,In_471,In_77);
nor U765 (N_765,In_477,In_72);
nor U766 (N_766,In_498,In_66);
nor U767 (N_767,In_486,In_37);
or U768 (N_768,In_488,In_208);
nand U769 (N_769,In_58,In_217);
nor U770 (N_770,In_46,In_285);
and U771 (N_771,In_233,In_496);
and U772 (N_772,In_288,In_317);
and U773 (N_773,In_176,In_78);
nor U774 (N_774,In_299,In_322);
and U775 (N_775,In_217,In_219);
or U776 (N_776,In_178,In_34);
and U777 (N_777,In_251,In_265);
nand U778 (N_778,In_485,In_163);
and U779 (N_779,In_119,In_26);
and U780 (N_780,In_96,In_401);
nor U781 (N_781,In_339,In_80);
nor U782 (N_782,In_115,In_1);
and U783 (N_783,In_117,In_175);
nor U784 (N_784,In_441,In_389);
nand U785 (N_785,In_275,In_407);
nor U786 (N_786,In_52,In_127);
nor U787 (N_787,In_59,In_427);
nand U788 (N_788,In_88,In_392);
or U789 (N_789,In_3,In_448);
or U790 (N_790,In_481,In_303);
or U791 (N_791,In_94,In_190);
or U792 (N_792,In_385,In_223);
and U793 (N_793,In_317,In_115);
nand U794 (N_794,In_112,In_375);
nor U795 (N_795,In_318,In_373);
nor U796 (N_796,In_299,In_298);
and U797 (N_797,In_462,In_432);
and U798 (N_798,In_209,In_439);
nor U799 (N_799,In_376,In_442);
and U800 (N_800,In_478,In_189);
nor U801 (N_801,In_255,In_345);
and U802 (N_802,In_2,In_124);
nor U803 (N_803,In_177,In_281);
or U804 (N_804,In_169,In_349);
nand U805 (N_805,In_68,In_471);
and U806 (N_806,In_123,In_358);
or U807 (N_807,In_246,In_212);
nand U808 (N_808,In_385,In_48);
nand U809 (N_809,In_130,In_165);
and U810 (N_810,In_335,In_150);
nand U811 (N_811,In_196,In_204);
nand U812 (N_812,In_308,In_128);
nor U813 (N_813,In_175,In_159);
nand U814 (N_814,In_341,In_188);
and U815 (N_815,In_388,In_313);
nand U816 (N_816,In_103,In_351);
nand U817 (N_817,In_466,In_212);
or U818 (N_818,In_295,In_413);
nor U819 (N_819,In_200,In_147);
and U820 (N_820,In_154,In_356);
nor U821 (N_821,In_17,In_421);
or U822 (N_822,In_266,In_174);
or U823 (N_823,In_396,In_235);
and U824 (N_824,In_174,In_189);
and U825 (N_825,In_278,In_271);
or U826 (N_826,In_77,In_422);
nor U827 (N_827,In_250,In_462);
or U828 (N_828,In_219,In_244);
or U829 (N_829,In_273,In_206);
nand U830 (N_830,In_486,In_193);
nand U831 (N_831,In_255,In_124);
or U832 (N_832,In_19,In_288);
nand U833 (N_833,In_159,In_50);
or U834 (N_834,In_390,In_196);
and U835 (N_835,In_247,In_162);
nand U836 (N_836,In_208,In_394);
and U837 (N_837,In_358,In_27);
nand U838 (N_838,In_70,In_454);
nand U839 (N_839,In_154,In_114);
and U840 (N_840,In_136,In_212);
nor U841 (N_841,In_352,In_452);
nand U842 (N_842,In_110,In_251);
nand U843 (N_843,In_389,In_249);
or U844 (N_844,In_226,In_107);
or U845 (N_845,In_150,In_451);
nor U846 (N_846,In_418,In_19);
nor U847 (N_847,In_395,In_366);
and U848 (N_848,In_235,In_295);
nor U849 (N_849,In_233,In_17);
nor U850 (N_850,In_474,In_65);
or U851 (N_851,In_376,In_356);
nand U852 (N_852,In_62,In_476);
nand U853 (N_853,In_41,In_72);
or U854 (N_854,In_36,In_183);
nand U855 (N_855,In_71,In_94);
nor U856 (N_856,In_211,In_184);
or U857 (N_857,In_375,In_86);
nor U858 (N_858,In_124,In_9);
xnor U859 (N_859,In_269,In_209);
nand U860 (N_860,In_20,In_365);
and U861 (N_861,In_330,In_272);
xnor U862 (N_862,In_277,In_109);
nor U863 (N_863,In_117,In_498);
nor U864 (N_864,In_334,In_467);
and U865 (N_865,In_144,In_422);
or U866 (N_866,In_177,In_86);
nor U867 (N_867,In_6,In_249);
nand U868 (N_868,In_134,In_157);
nor U869 (N_869,In_324,In_93);
nor U870 (N_870,In_370,In_176);
and U871 (N_871,In_134,In_222);
or U872 (N_872,In_39,In_384);
or U873 (N_873,In_73,In_489);
and U874 (N_874,In_325,In_132);
or U875 (N_875,In_389,In_43);
nor U876 (N_876,In_20,In_201);
and U877 (N_877,In_274,In_343);
nor U878 (N_878,In_463,In_424);
nor U879 (N_879,In_323,In_67);
and U880 (N_880,In_243,In_56);
nand U881 (N_881,In_112,In_240);
and U882 (N_882,In_331,In_130);
nand U883 (N_883,In_424,In_194);
nand U884 (N_884,In_450,In_322);
nor U885 (N_885,In_68,In_439);
and U886 (N_886,In_392,In_59);
nand U887 (N_887,In_10,In_25);
nand U888 (N_888,In_260,In_381);
nor U889 (N_889,In_70,In_288);
nor U890 (N_890,In_61,In_134);
and U891 (N_891,In_49,In_195);
nand U892 (N_892,In_192,In_422);
and U893 (N_893,In_209,In_300);
or U894 (N_894,In_162,In_445);
nor U895 (N_895,In_481,In_104);
nor U896 (N_896,In_328,In_112);
and U897 (N_897,In_241,In_86);
or U898 (N_898,In_312,In_402);
and U899 (N_899,In_183,In_65);
and U900 (N_900,In_479,In_262);
or U901 (N_901,In_18,In_389);
and U902 (N_902,In_313,In_306);
nor U903 (N_903,In_495,In_498);
nor U904 (N_904,In_108,In_438);
nand U905 (N_905,In_54,In_234);
or U906 (N_906,In_104,In_102);
or U907 (N_907,In_257,In_11);
or U908 (N_908,In_46,In_342);
nor U909 (N_909,In_329,In_112);
or U910 (N_910,In_227,In_105);
nand U911 (N_911,In_182,In_7);
or U912 (N_912,In_365,In_151);
or U913 (N_913,In_205,In_475);
or U914 (N_914,In_400,In_96);
nand U915 (N_915,In_265,In_151);
nor U916 (N_916,In_105,In_32);
and U917 (N_917,In_476,In_495);
or U918 (N_918,In_366,In_352);
and U919 (N_919,In_123,In_63);
or U920 (N_920,In_312,In_207);
nand U921 (N_921,In_310,In_495);
nor U922 (N_922,In_383,In_410);
nand U923 (N_923,In_136,In_151);
nand U924 (N_924,In_113,In_149);
and U925 (N_925,In_236,In_455);
or U926 (N_926,In_159,In_400);
and U927 (N_927,In_308,In_0);
nor U928 (N_928,In_385,In_173);
and U929 (N_929,In_401,In_93);
nor U930 (N_930,In_346,In_86);
and U931 (N_931,In_475,In_288);
and U932 (N_932,In_378,In_384);
and U933 (N_933,In_356,In_477);
nor U934 (N_934,In_270,In_258);
xor U935 (N_935,In_443,In_344);
or U936 (N_936,In_363,In_110);
nand U937 (N_937,In_293,In_251);
and U938 (N_938,In_145,In_81);
nor U939 (N_939,In_234,In_135);
or U940 (N_940,In_50,In_260);
and U941 (N_941,In_391,In_270);
nand U942 (N_942,In_279,In_122);
or U943 (N_943,In_170,In_107);
and U944 (N_944,In_231,In_431);
or U945 (N_945,In_145,In_320);
nor U946 (N_946,In_111,In_30);
nor U947 (N_947,In_165,In_292);
and U948 (N_948,In_286,In_225);
nand U949 (N_949,In_234,In_305);
nand U950 (N_950,In_296,In_169);
nor U951 (N_951,In_74,In_103);
and U952 (N_952,In_489,In_102);
nor U953 (N_953,In_465,In_34);
or U954 (N_954,In_200,In_83);
or U955 (N_955,In_396,In_65);
and U956 (N_956,In_42,In_463);
nor U957 (N_957,In_98,In_46);
nor U958 (N_958,In_279,In_244);
or U959 (N_959,In_178,In_493);
or U960 (N_960,In_430,In_13);
and U961 (N_961,In_92,In_354);
and U962 (N_962,In_4,In_52);
and U963 (N_963,In_214,In_472);
nor U964 (N_964,In_370,In_332);
nor U965 (N_965,In_380,In_450);
or U966 (N_966,In_137,In_301);
or U967 (N_967,In_37,In_216);
or U968 (N_968,In_471,In_61);
nand U969 (N_969,In_111,In_432);
and U970 (N_970,In_344,In_267);
nor U971 (N_971,In_142,In_304);
and U972 (N_972,In_6,In_173);
nand U973 (N_973,In_296,In_300);
or U974 (N_974,In_392,In_453);
or U975 (N_975,In_27,In_251);
nand U976 (N_976,In_244,In_348);
nand U977 (N_977,In_234,In_425);
nand U978 (N_978,In_458,In_182);
and U979 (N_979,In_296,In_425);
nand U980 (N_980,In_24,In_191);
or U981 (N_981,In_201,In_113);
and U982 (N_982,In_130,In_323);
and U983 (N_983,In_33,In_476);
or U984 (N_984,In_328,In_298);
or U985 (N_985,In_402,In_418);
and U986 (N_986,In_432,In_372);
nor U987 (N_987,In_299,In_303);
and U988 (N_988,In_231,In_211);
nand U989 (N_989,In_167,In_249);
nor U990 (N_990,In_202,In_329);
nand U991 (N_991,In_219,In_139);
and U992 (N_992,In_245,In_205);
nor U993 (N_993,In_412,In_287);
nor U994 (N_994,In_350,In_294);
nor U995 (N_995,In_134,In_288);
and U996 (N_996,In_41,In_356);
or U997 (N_997,In_304,In_31);
or U998 (N_998,In_260,In_60);
or U999 (N_999,In_14,In_135);
and U1000 (N_1000,N_120,N_417);
and U1001 (N_1001,N_205,N_565);
or U1002 (N_1002,N_840,N_960);
or U1003 (N_1003,N_548,N_515);
nand U1004 (N_1004,N_309,N_701);
nand U1005 (N_1005,N_106,N_697);
or U1006 (N_1006,N_787,N_43);
nand U1007 (N_1007,N_335,N_508);
nand U1008 (N_1008,N_892,N_645);
nor U1009 (N_1009,N_729,N_597);
or U1010 (N_1010,N_40,N_483);
nand U1011 (N_1011,N_285,N_741);
nand U1012 (N_1012,N_653,N_896);
nor U1013 (N_1013,N_372,N_656);
and U1014 (N_1014,N_466,N_222);
and U1015 (N_1015,N_608,N_428);
or U1016 (N_1016,N_540,N_368);
xor U1017 (N_1017,N_487,N_952);
nand U1018 (N_1018,N_983,N_533);
or U1019 (N_1019,N_180,N_255);
and U1020 (N_1020,N_611,N_676);
and U1021 (N_1021,N_659,N_705);
or U1022 (N_1022,N_855,N_674);
or U1023 (N_1023,N_410,N_901);
or U1024 (N_1024,N_273,N_332);
or U1025 (N_1025,N_196,N_346);
and U1026 (N_1026,N_987,N_152);
nor U1027 (N_1027,N_637,N_703);
nand U1028 (N_1028,N_61,N_31);
or U1029 (N_1029,N_799,N_329);
or U1030 (N_1030,N_925,N_225);
and U1031 (N_1031,N_795,N_53);
and U1032 (N_1032,N_234,N_903);
or U1033 (N_1033,N_721,N_405);
nand U1034 (N_1034,N_857,N_14);
nand U1035 (N_1035,N_917,N_238);
nand U1036 (N_1036,N_739,N_619);
nand U1037 (N_1037,N_157,N_360);
or U1038 (N_1038,N_74,N_162);
or U1039 (N_1039,N_570,N_700);
and U1040 (N_1040,N_810,N_35);
and U1041 (N_1041,N_291,N_861);
or U1042 (N_1042,N_618,N_376);
or U1043 (N_1043,N_782,N_842);
or U1044 (N_1044,N_272,N_558);
and U1045 (N_1045,N_2,N_937);
or U1046 (N_1046,N_140,N_947);
nor U1047 (N_1047,N_704,N_292);
and U1048 (N_1048,N_747,N_45);
or U1049 (N_1049,N_490,N_315);
or U1050 (N_1050,N_841,N_145);
nand U1051 (N_1051,N_698,N_848);
nor U1052 (N_1052,N_874,N_616);
nand U1053 (N_1053,N_679,N_362);
or U1054 (N_1054,N_274,N_334);
xor U1055 (N_1055,N_563,N_657);
and U1056 (N_1056,N_716,N_123);
or U1057 (N_1057,N_615,N_564);
nor U1058 (N_1058,N_582,N_149);
and U1059 (N_1059,N_764,N_21);
nor U1060 (N_1060,N_757,N_994);
nand U1061 (N_1061,N_265,N_885);
nand U1062 (N_1062,N_651,N_707);
and U1063 (N_1063,N_153,N_522);
nor U1064 (N_1064,N_312,N_424);
and U1065 (N_1065,N_509,N_601);
nand U1066 (N_1066,N_461,N_517);
nor U1067 (N_1067,N_497,N_37);
and U1068 (N_1068,N_210,N_830);
nor U1069 (N_1069,N_437,N_17);
and U1070 (N_1070,N_838,N_436);
nor U1071 (N_1071,N_480,N_792);
nor U1072 (N_1072,N_529,N_160);
nor U1073 (N_1073,N_804,N_101);
and U1074 (N_1074,N_696,N_228);
or U1075 (N_1075,N_536,N_96);
nand U1076 (N_1076,N_215,N_752);
or U1077 (N_1077,N_220,N_507);
and U1078 (N_1078,N_778,N_636);
or U1079 (N_1079,N_237,N_82);
or U1080 (N_1080,N_911,N_904);
nor U1081 (N_1081,N_866,N_849);
nor U1082 (N_1082,N_229,N_572);
or U1083 (N_1083,N_403,N_734);
and U1084 (N_1084,N_688,N_467);
or U1085 (N_1085,N_71,N_641);
nand U1086 (N_1086,N_279,N_539);
nor U1087 (N_1087,N_54,N_455);
or U1088 (N_1088,N_206,N_571);
nand U1089 (N_1089,N_389,N_643);
nand U1090 (N_1090,N_109,N_786);
nor U1091 (N_1091,N_769,N_800);
nand U1092 (N_1092,N_502,N_603);
nand U1093 (N_1093,N_468,N_452);
or U1094 (N_1094,N_982,N_107);
nor U1095 (N_1095,N_683,N_433);
nor U1096 (N_1096,N_882,N_669);
xnor U1097 (N_1097,N_811,N_457);
nor U1098 (N_1098,N_444,N_48);
and U1099 (N_1099,N_835,N_336);
or U1100 (N_1100,N_541,N_382);
nor U1101 (N_1101,N_358,N_95);
nor U1102 (N_1102,N_19,N_890);
or U1103 (N_1103,N_355,N_197);
nand U1104 (N_1104,N_257,N_246);
nor U1105 (N_1105,N_913,N_875);
or U1106 (N_1106,N_105,N_300);
nor U1107 (N_1107,N_387,N_143);
nor U1108 (N_1108,N_859,N_104);
and U1109 (N_1109,N_774,N_858);
nor U1110 (N_1110,N_22,N_469);
and U1111 (N_1111,N_673,N_780);
and U1112 (N_1112,N_844,N_204);
or U1113 (N_1113,N_131,N_116);
nand U1114 (N_1114,N_585,N_187);
nand U1115 (N_1115,N_141,N_744);
and U1116 (N_1116,N_494,N_422);
nor U1117 (N_1117,N_944,N_337);
or U1118 (N_1118,N_344,N_83);
nor U1119 (N_1119,N_612,N_532);
nor U1120 (N_1120,N_167,N_826);
and U1121 (N_1121,N_60,N_883);
or U1122 (N_1122,N_393,N_562);
or U1123 (N_1123,N_170,N_356);
and U1124 (N_1124,N_420,N_55);
and U1125 (N_1125,N_52,N_295);
nor U1126 (N_1126,N_535,N_284);
nor U1127 (N_1127,N_652,N_863);
or U1128 (N_1128,N_974,N_70);
and U1129 (N_1129,N_341,N_834);
and U1130 (N_1130,N_798,N_458);
nor U1131 (N_1131,N_9,N_333);
and U1132 (N_1132,N_137,N_640);
or U1133 (N_1133,N_134,N_650);
nand U1134 (N_1134,N_259,N_577);
nand U1135 (N_1135,N_302,N_998);
nand U1136 (N_1136,N_28,N_527);
and U1137 (N_1137,N_317,N_918);
nor U1138 (N_1138,N_520,N_796);
nand U1139 (N_1139,N_516,N_419);
or U1140 (N_1140,N_371,N_690);
or U1141 (N_1141,N_837,N_899);
or U1142 (N_1142,N_32,N_915);
nand U1143 (N_1143,N_51,N_794);
or U1144 (N_1144,N_7,N_489);
or U1145 (N_1145,N_477,N_230);
nand U1146 (N_1146,N_537,N_694);
nor U1147 (N_1147,N_59,N_260);
or U1148 (N_1148,N_130,N_755);
or U1149 (N_1149,N_10,N_610);
xnor U1150 (N_1150,N_921,N_808);
and U1151 (N_1151,N_756,N_631);
nor U1152 (N_1152,N_776,N_948);
and U1153 (N_1153,N_730,N_24);
or U1154 (N_1154,N_8,N_596);
or U1155 (N_1155,N_168,N_208);
or U1156 (N_1156,N_248,N_390);
nor U1157 (N_1157,N_593,N_661);
or U1158 (N_1158,N_606,N_972);
and U1159 (N_1159,N_303,N_126);
or U1160 (N_1160,N_414,N_607);
nand U1161 (N_1161,N_854,N_860);
and U1162 (N_1162,N_430,N_20);
or U1163 (N_1163,N_500,N_117);
or U1164 (N_1164,N_560,N_313);
nor U1165 (N_1165,N_938,N_154);
or U1166 (N_1166,N_240,N_587);
and U1167 (N_1167,N_87,N_267);
nand U1168 (N_1168,N_453,N_809);
or U1169 (N_1169,N_677,N_579);
nor U1170 (N_1170,N_634,N_289);
and U1171 (N_1171,N_16,N_110);
or U1172 (N_1172,N_602,N_488);
and U1173 (N_1173,N_3,N_797);
nand U1174 (N_1174,N_588,N_351);
or U1175 (N_1175,N_584,N_373);
nand U1176 (N_1176,N_250,N_667);
or U1177 (N_1177,N_977,N_962);
nor U1178 (N_1178,N_412,N_266);
or U1179 (N_1179,N_980,N_446);
and U1180 (N_1180,N_103,N_98);
nand U1181 (N_1181,N_299,N_802);
or U1182 (N_1182,N_544,N_714);
or U1183 (N_1183,N_114,N_280);
and U1184 (N_1184,N_252,N_906);
nand U1185 (N_1185,N_803,N_49);
nand U1186 (N_1186,N_297,N_672);
nand U1187 (N_1187,N_407,N_581);
and U1188 (N_1188,N_176,N_354);
or U1189 (N_1189,N_852,N_256);
xnor U1190 (N_1190,N_715,N_865);
and U1191 (N_1191,N_682,N_448);
and U1192 (N_1192,N_871,N_324);
nor U1193 (N_1193,N_594,N_148);
and U1194 (N_1194,N_833,N_326);
nand U1195 (N_1195,N_772,N_689);
nor U1196 (N_1196,N_819,N_945);
and U1197 (N_1197,N_484,N_818);
nor U1198 (N_1198,N_869,N_46);
and U1199 (N_1199,N_965,N_888);
or U1200 (N_1200,N_567,N_680);
and U1201 (N_1201,N_968,N_993);
nand U1202 (N_1202,N_68,N_831);
nand U1203 (N_1203,N_85,N_853);
nand U1204 (N_1204,N_415,N_200);
or U1205 (N_1205,N_304,N_970);
nor U1206 (N_1206,N_973,N_129);
nor U1207 (N_1207,N_666,N_505);
and U1208 (N_1208,N_323,N_367);
and U1209 (N_1209,N_749,N_374);
nand U1210 (N_1210,N_327,N_247);
nand U1211 (N_1211,N_216,N_50);
and U1212 (N_1212,N_307,N_348);
nor U1213 (N_1213,N_733,N_413);
and U1214 (N_1214,N_727,N_967);
nand U1215 (N_1215,N_771,N_203);
or U1216 (N_1216,N_894,N_660);
nor U1217 (N_1217,N_881,N_534);
nand U1218 (N_1218,N_406,N_271);
nor U1219 (N_1219,N_979,N_165);
nor U1220 (N_1220,N_194,N_243);
nand U1221 (N_1221,N_649,N_963);
and U1222 (N_1222,N_531,N_825);
or U1223 (N_1223,N_552,N_63);
nand U1224 (N_1224,N_270,N_732);
nand U1225 (N_1225,N_978,N_575);
nor U1226 (N_1226,N_112,N_648);
or U1227 (N_1227,N_202,N_832);
nor U1228 (N_1228,N_378,N_359);
or U1229 (N_1229,N_870,N_501);
nand U1230 (N_1230,N_627,N_876);
or U1231 (N_1231,N_791,N_182);
and U1232 (N_1232,N_905,N_454);
or U1233 (N_1233,N_64,N_261);
and U1234 (N_1234,N_958,N_122);
nor U1235 (N_1235,N_924,N_282);
or U1236 (N_1236,N_347,N_908);
nand U1237 (N_1237,N_545,N_161);
nand U1238 (N_1238,N_133,N_512);
nor U1239 (N_1239,N_159,N_298);
nor U1240 (N_1240,N_824,N_884);
nor U1241 (N_1241,N_635,N_1);
and U1242 (N_1242,N_15,N_604);
and U1243 (N_1243,N_275,N_817);
nor U1244 (N_1244,N_935,N_499);
nor U1245 (N_1245,N_693,N_766);
and U1246 (N_1246,N_249,N_986);
nor U1247 (N_1247,N_183,N_872);
or U1248 (N_1248,N_330,N_76);
nor U1249 (N_1249,N_592,N_42);
or U1250 (N_1250,N_151,N_318);
or U1251 (N_1251,N_4,N_177);
or U1252 (N_1252,N_801,N_418);
and U1253 (N_1253,N_268,N_614);
or U1254 (N_1254,N_773,N_370);
nand U1255 (N_1255,N_169,N_439);
or U1256 (N_1256,N_338,N_164);
nor U1257 (N_1257,N_97,N_877);
nand U1258 (N_1258,N_687,N_922);
nand U1259 (N_1259,N_878,N_495);
nand U1260 (N_1260,N_94,N_242);
nor U1261 (N_1261,N_699,N_868);
and U1262 (N_1262,N_235,N_57);
or U1263 (N_1263,N_451,N_75);
xnor U1264 (N_1264,N_902,N_224);
nor U1265 (N_1265,N_662,N_12);
and U1266 (N_1266,N_391,N_613);
nor U1267 (N_1267,N_599,N_538);
and U1268 (N_1268,N_294,N_511);
nand U1269 (N_1269,N_746,N_665);
or U1270 (N_1270,N_263,N_595);
nor U1271 (N_1271,N_339,N_984);
nor U1272 (N_1272,N_940,N_740);
nand U1273 (N_1273,N_171,N_524);
nand U1274 (N_1274,N_719,N_115);
or U1275 (N_1275,N_692,N_0);
nand U1276 (N_1276,N_325,N_462);
nand U1277 (N_1277,N_723,N_990);
or U1278 (N_1278,N_758,N_851);
and U1279 (N_1279,N_301,N_836);
nor U1280 (N_1280,N_961,N_231);
and U1281 (N_1281,N_530,N_743);
and U1282 (N_1282,N_873,N_191);
or U1283 (N_1283,N_314,N_828);
nand U1284 (N_1284,N_551,N_623);
or U1285 (N_1285,N_621,N_379);
or U1286 (N_1286,N_375,N_626);
and U1287 (N_1287,N_654,N_471);
and U1288 (N_1288,N_181,N_720);
or U1289 (N_1289,N_158,N_384);
nor U1290 (N_1290,N_258,N_793);
and U1291 (N_1291,N_113,N_65);
nor U1292 (N_1292,N_543,N_90);
nand U1293 (N_1293,N_125,N_638);
and U1294 (N_1294,N_342,N_118);
nand U1295 (N_1295,N_226,N_622);
nor U1296 (N_1296,N_431,N_717);
and U1297 (N_1297,N_556,N_67);
nor U1298 (N_1298,N_762,N_929);
and U1299 (N_1299,N_44,N_155);
nor U1300 (N_1300,N_789,N_434);
nor U1301 (N_1301,N_425,N_435);
nand U1302 (N_1302,N_449,N_144);
or U1303 (N_1303,N_456,N_775);
nor U1304 (N_1304,N_62,N_969);
xnor U1305 (N_1305,N_549,N_486);
nand U1306 (N_1306,N_528,N_427);
or U1307 (N_1307,N_846,N_566);
and U1308 (N_1308,N_179,N_710);
nand U1309 (N_1309,N_748,N_363);
and U1310 (N_1310,N_737,N_163);
nand U1311 (N_1311,N_349,N_440);
and U1312 (N_1312,N_718,N_573);
and U1313 (N_1313,N_394,N_568);
xor U1314 (N_1314,N_788,N_283);
and U1315 (N_1315,N_685,N_293);
and U1316 (N_1316,N_11,N_686);
or U1317 (N_1317,N_423,N_521);
nand U1318 (N_1318,N_630,N_898);
or U1319 (N_1319,N_438,N_353);
and U1320 (N_1320,N_172,N_555);
or U1321 (N_1321,N_777,N_121);
or U1322 (N_1322,N_930,N_681);
or U1323 (N_1323,N_56,N_966);
and U1324 (N_1324,N_829,N_580);
nor U1325 (N_1325,N_33,N_916);
and U1326 (N_1326,N_178,N_475);
or U1327 (N_1327,N_862,N_934);
and U1328 (N_1328,N_276,N_767);
or U1329 (N_1329,N_478,N_476);
and U1330 (N_1330,N_943,N_695);
nand U1331 (N_1331,N_557,N_702);
or U1332 (N_1332,N_350,N_311);
and U1333 (N_1333,N_957,N_269);
or U1334 (N_1334,N_23,N_496);
or U1335 (N_1335,N_946,N_262);
nor U1336 (N_1336,N_923,N_460);
or U1337 (N_1337,N_956,N_322);
and U1338 (N_1338,N_569,N_213);
or U1339 (N_1339,N_928,N_675);
nand U1340 (N_1340,N_561,N_736);
nor U1341 (N_1341,N_907,N_620);
or U1342 (N_1342,N_352,N_212);
nand U1343 (N_1343,N_542,N_815);
or U1344 (N_1344,N_84,N_482);
nor U1345 (N_1345,N_411,N_73);
nor U1346 (N_1346,N_910,N_678);
nor U1347 (N_1347,N_932,N_81);
and U1348 (N_1348,N_949,N_760);
and U1349 (N_1349,N_820,N_472);
nand U1350 (N_1350,N_429,N_396);
nand U1351 (N_1351,N_443,N_843);
or U1352 (N_1352,N_399,N_463);
and U1353 (N_1353,N_209,N_18);
nor U1354 (N_1354,N_119,N_217);
xnor U1355 (N_1355,N_731,N_976);
nand U1356 (N_1356,N_600,N_328);
nand U1357 (N_1357,N_559,N_554);
and U1358 (N_1358,N_442,N_670);
and U1359 (N_1359,N_574,N_290);
nand U1360 (N_1360,N_340,N_964);
or U1361 (N_1361,N_850,N_609);
nand U1362 (N_1362,N_72,N_278);
and U1363 (N_1363,N_813,N_343);
nand U1364 (N_1364,N_503,N_708);
nor U1365 (N_1365,N_807,N_211);
nor U1366 (N_1366,N_219,N_245);
and U1367 (N_1367,N_69,N_136);
nand U1368 (N_1368,N_821,N_790);
or U1369 (N_1369,N_847,N_646);
nor U1370 (N_1370,N_954,N_288);
and U1371 (N_1371,N_959,N_691);
and U1372 (N_1372,N_712,N_124);
nor U1373 (N_1373,N_995,N_805);
nor U1374 (N_1374,N_232,N_485);
nand U1375 (N_1375,N_989,N_498);
and U1376 (N_1376,N_753,N_199);
nor U1377 (N_1377,N_244,N_658);
xor U1378 (N_1378,N_895,N_195);
and U1379 (N_1379,N_184,N_421);
or U1380 (N_1380,N_839,N_447);
and U1381 (N_1381,N_981,N_492);
and U1382 (N_1382,N_320,N_632);
or U1383 (N_1383,N_404,N_951);
or U1384 (N_1384,N_950,N_47);
or U1385 (N_1385,N_39,N_6);
nand U1386 (N_1386,N_175,N_578);
or U1387 (N_1387,N_409,N_470);
and U1388 (N_1388,N_920,N_281);
nand U1389 (N_1389,N_138,N_189);
or U1390 (N_1390,N_201,N_926);
and U1391 (N_1391,N_441,N_759);
and U1392 (N_1392,N_254,N_763);
and U1393 (N_1393,N_400,N_893);
and U1394 (N_1394,N_806,N_814);
nand U1395 (N_1395,N_264,N_66);
and U1396 (N_1396,N_479,N_589);
and U1397 (N_1397,N_655,N_132);
or U1398 (N_1398,N_432,N_889);
nor U1399 (N_1399,N_416,N_519);
nor U1400 (N_1400,N_306,N_38);
nor U1401 (N_1401,N_971,N_150);
nand U1402 (N_1402,N_931,N_459);
and U1403 (N_1403,N_305,N_880);
nand U1404 (N_1404,N_985,N_642);
nor U1405 (N_1405,N_823,N_504);
and U1406 (N_1406,N_174,N_975);
nand U1407 (N_1407,N_91,N_768);
nor U1408 (N_1408,N_812,N_41);
or U1409 (N_1409,N_713,N_668);
and U1410 (N_1410,N_735,N_88);
and U1411 (N_1411,N_386,N_518);
nand U1412 (N_1412,N_754,N_464);
nand U1413 (N_1413,N_864,N_856);
nand U1414 (N_1414,N_991,N_36);
nand U1415 (N_1415,N_380,N_845);
or U1416 (N_1416,N_392,N_77);
nor U1417 (N_1417,N_583,N_722);
and U1418 (N_1418,N_357,N_779);
or U1419 (N_1419,N_398,N_385);
nand U1420 (N_1420,N_111,N_953);
and U1421 (N_1421,N_628,N_728);
nor U1422 (N_1422,N_383,N_625);
nor U1423 (N_1423,N_364,N_99);
and U1424 (N_1424,N_218,N_102);
and U1425 (N_1425,N_93,N_933);
and U1426 (N_1426,N_92,N_253);
or U1427 (N_1427,N_781,N_214);
and U1428 (N_1428,N_127,N_591);
nand U1429 (N_1429,N_879,N_726);
or U1430 (N_1430,N_891,N_108);
and U1431 (N_1431,N_605,N_887);
nand U1432 (N_1432,N_784,N_369);
nor U1433 (N_1433,N_550,N_445);
nor U1434 (N_1434,N_525,N_233);
or U1435 (N_1435,N_58,N_186);
nor U1436 (N_1436,N_664,N_867);
and U1437 (N_1437,N_185,N_277);
nor U1438 (N_1438,N_785,N_927);
nand U1439 (N_1439,N_395,N_709);
and U1440 (N_1440,N_745,N_365);
or U1441 (N_1441,N_331,N_761);
and U1442 (N_1442,N_78,N_955);
nor U1443 (N_1443,N_765,N_381);
and U1444 (N_1444,N_647,N_783);
or U1445 (N_1445,N_366,N_156);
nor U1446 (N_1446,N_724,N_912);
and U1447 (N_1447,N_34,N_514);
and U1448 (N_1448,N_308,N_465);
nor U1449 (N_1449,N_25,N_27);
nor U1450 (N_1450,N_361,N_816);
nor U1451 (N_1451,N_936,N_86);
nand U1452 (N_1452,N_706,N_79);
nand U1453 (N_1453,N_345,N_100);
nand U1454 (N_1454,N_506,N_128);
and U1455 (N_1455,N_629,N_473);
and U1456 (N_1456,N_992,N_377);
nor U1457 (N_1457,N_188,N_135);
nand U1458 (N_1458,N_13,N_236);
nor U1459 (N_1459,N_725,N_751);
or U1460 (N_1460,N_30,N_426);
or U1461 (N_1461,N_319,N_919);
nor U1462 (N_1462,N_474,N_547);
nor U1463 (N_1463,N_493,N_227);
and U1464 (N_1464,N_914,N_190);
nor U1465 (N_1465,N_146,N_553);
or U1466 (N_1466,N_296,N_142);
nand U1467 (N_1467,N_546,N_139);
nor U1468 (N_1468,N_909,N_822);
and U1469 (N_1469,N_147,N_239);
nor U1470 (N_1470,N_491,N_192);
and U1471 (N_1471,N_166,N_397);
nand U1472 (N_1472,N_941,N_316);
and U1473 (N_1473,N_193,N_173);
or U1474 (N_1474,N_996,N_5);
nand U1475 (N_1475,N_401,N_221);
nand U1476 (N_1476,N_576,N_663);
nor U1477 (N_1477,N_742,N_198);
nor U1478 (N_1478,N_639,N_598);
nand U1479 (N_1479,N_827,N_750);
and U1480 (N_1480,N_241,N_321);
and U1481 (N_1481,N_988,N_586);
nand U1482 (N_1482,N_207,N_510);
or U1483 (N_1483,N_624,N_388);
nor U1484 (N_1484,N_671,N_526);
or U1485 (N_1485,N_287,N_939);
and U1486 (N_1486,N_89,N_29);
nand U1487 (N_1487,N_26,N_997);
and U1488 (N_1488,N_738,N_617);
nor U1489 (N_1489,N_684,N_408);
nor U1490 (N_1490,N_223,N_450);
or U1491 (N_1491,N_402,N_770);
or U1492 (N_1492,N_942,N_633);
nor U1493 (N_1493,N_310,N_897);
and U1494 (N_1494,N_590,N_513);
nor U1495 (N_1495,N_80,N_481);
and U1496 (N_1496,N_886,N_999);
nor U1497 (N_1497,N_711,N_286);
nor U1498 (N_1498,N_644,N_523);
nor U1499 (N_1499,N_900,N_251);
or U1500 (N_1500,N_409,N_632);
nor U1501 (N_1501,N_746,N_21);
or U1502 (N_1502,N_847,N_566);
or U1503 (N_1503,N_13,N_465);
nand U1504 (N_1504,N_103,N_467);
and U1505 (N_1505,N_813,N_373);
nor U1506 (N_1506,N_35,N_969);
and U1507 (N_1507,N_899,N_214);
nand U1508 (N_1508,N_449,N_997);
nand U1509 (N_1509,N_94,N_278);
nand U1510 (N_1510,N_684,N_672);
nor U1511 (N_1511,N_912,N_507);
nand U1512 (N_1512,N_673,N_225);
and U1513 (N_1513,N_293,N_921);
nand U1514 (N_1514,N_35,N_499);
nor U1515 (N_1515,N_301,N_26);
nand U1516 (N_1516,N_614,N_217);
nand U1517 (N_1517,N_402,N_640);
and U1518 (N_1518,N_991,N_81);
nor U1519 (N_1519,N_120,N_480);
nand U1520 (N_1520,N_402,N_777);
nor U1521 (N_1521,N_236,N_389);
nand U1522 (N_1522,N_974,N_172);
or U1523 (N_1523,N_883,N_58);
and U1524 (N_1524,N_721,N_944);
nor U1525 (N_1525,N_9,N_358);
nand U1526 (N_1526,N_165,N_934);
and U1527 (N_1527,N_701,N_523);
nand U1528 (N_1528,N_194,N_276);
or U1529 (N_1529,N_627,N_443);
or U1530 (N_1530,N_595,N_203);
nor U1531 (N_1531,N_150,N_289);
nand U1532 (N_1532,N_487,N_550);
and U1533 (N_1533,N_611,N_979);
nor U1534 (N_1534,N_65,N_35);
nand U1535 (N_1535,N_789,N_504);
nor U1536 (N_1536,N_759,N_171);
nor U1537 (N_1537,N_205,N_949);
and U1538 (N_1538,N_469,N_123);
nand U1539 (N_1539,N_768,N_284);
or U1540 (N_1540,N_17,N_191);
nand U1541 (N_1541,N_674,N_530);
and U1542 (N_1542,N_70,N_439);
nor U1543 (N_1543,N_259,N_544);
nor U1544 (N_1544,N_322,N_96);
or U1545 (N_1545,N_235,N_896);
nand U1546 (N_1546,N_59,N_171);
or U1547 (N_1547,N_831,N_997);
and U1548 (N_1548,N_891,N_892);
or U1549 (N_1549,N_201,N_577);
nor U1550 (N_1550,N_624,N_849);
or U1551 (N_1551,N_798,N_752);
nand U1552 (N_1552,N_606,N_892);
or U1553 (N_1553,N_339,N_128);
and U1554 (N_1554,N_587,N_593);
nand U1555 (N_1555,N_937,N_843);
or U1556 (N_1556,N_226,N_390);
nor U1557 (N_1557,N_468,N_787);
and U1558 (N_1558,N_158,N_184);
nor U1559 (N_1559,N_42,N_538);
nor U1560 (N_1560,N_550,N_868);
and U1561 (N_1561,N_329,N_511);
or U1562 (N_1562,N_563,N_36);
and U1563 (N_1563,N_56,N_328);
nand U1564 (N_1564,N_880,N_524);
nor U1565 (N_1565,N_20,N_990);
and U1566 (N_1566,N_513,N_681);
or U1567 (N_1567,N_173,N_499);
nand U1568 (N_1568,N_890,N_687);
nand U1569 (N_1569,N_127,N_588);
nand U1570 (N_1570,N_190,N_346);
nor U1571 (N_1571,N_735,N_493);
nor U1572 (N_1572,N_194,N_794);
nor U1573 (N_1573,N_820,N_493);
nor U1574 (N_1574,N_418,N_303);
and U1575 (N_1575,N_209,N_590);
nor U1576 (N_1576,N_284,N_514);
nor U1577 (N_1577,N_54,N_57);
and U1578 (N_1578,N_491,N_399);
nand U1579 (N_1579,N_110,N_696);
or U1580 (N_1580,N_393,N_979);
nand U1581 (N_1581,N_76,N_209);
and U1582 (N_1582,N_319,N_477);
nand U1583 (N_1583,N_831,N_246);
nand U1584 (N_1584,N_366,N_136);
nor U1585 (N_1585,N_612,N_914);
and U1586 (N_1586,N_200,N_304);
nand U1587 (N_1587,N_53,N_47);
and U1588 (N_1588,N_126,N_793);
nor U1589 (N_1589,N_267,N_877);
nand U1590 (N_1590,N_821,N_831);
nand U1591 (N_1591,N_588,N_17);
nand U1592 (N_1592,N_877,N_650);
or U1593 (N_1593,N_494,N_852);
nand U1594 (N_1594,N_883,N_964);
or U1595 (N_1595,N_286,N_33);
and U1596 (N_1596,N_83,N_358);
nor U1597 (N_1597,N_151,N_870);
and U1598 (N_1598,N_713,N_313);
nor U1599 (N_1599,N_680,N_604);
nand U1600 (N_1600,N_785,N_486);
or U1601 (N_1601,N_608,N_582);
xnor U1602 (N_1602,N_584,N_963);
nand U1603 (N_1603,N_990,N_796);
or U1604 (N_1604,N_321,N_210);
and U1605 (N_1605,N_858,N_815);
nor U1606 (N_1606,N_96,N_702);
nand U1607 (N_1607,N_901,N_183);
or U1608 (N_1608,N_413,N_322);
and U1609 (N_1609,N_783,N_598);
xnor U1610 (N_1610,N_608,N_108);
nor U1611 (N_1611,N_313,N_847);
nand U1612 (N_1612,N_870,N_645);
nand U1613 (N_1613,N_234,N_810);
nand U1614 (N_1614,N_740,N_321);
nor U1615 (N_1615,N_856,N_80);
and U1616 (N_1616,N_78,N_49);
and U1617 (N_1617,N_765,N_66);
nand U1618 (N_1618,N_95,N_215);
nor U1619 (N_1619,N_353,N_993);
nor U1620 (N_1620,N_923,N_397);
or U1621 (N_1621,N_589,N_991);
nand U1622 (N_1622,N_471,N_502);
nor U1623 (N_1623,N_260,N_154);
or U1624 (N_1624,N_12,N_202);
or U1625 (N_1625,N_342,N_592);
and U1626 (N_1626,N_463,N_767);
nor U1627 (N_1627,N_296,N_783);
nand U1628 (N_1628,N_170,N_794);
or U1629 (N_1629,N_534,N_177);
nand U1630 (N_1630,N_237,N_753);
nor U1631 (N_1631,N_776,N_696);
and U1632 (N_1632,N_732,N_900);
or U1633 (N_1633,N_310,N_536);
and U1634 (N_1634,N_214,N_44);
nor U1635 (N_1635,N_547,N_341);
and U1636 (N_1636,N_978,N_880);
or U1637 (N_1637,N_918,N_994);
nand U1638 (N_1638,N_473,N_183);
nor U1639 (N_1639,N_170,N_746);
nand U1640 (N_1640,N_658,N_838);
nand U1641 (N_1641,N_304,N_272);
nand U1642 (N_1642,N_690,N_97);
nand U1643 (N_1643,N_840,N_874);
or U1644 (N_1644,N_217,N_482);
nor U1645 (N_1645,N_980,N_581);
nor U1646 (N_1646,N_76,N_146);
nor U1647 (N_1647,N_693,N_33);
and U1648 (N_1648,N_277,N_371);
nor U1649 (N_1649,N_954,N_864);
xor U1650 (N_1650,N_325,N_142);
and U1651 (N_1651,N_669,N_792);
nor U1652 (N_1652,N_502,N_494);
nand U1653 (N_1653,N_3,N_45);
and U1654 (N_1654,N_642,N_986);
nand U1655 (N_1655,N_495,N_20);
nor U1656 (N_1656,N_803,N_562);
nor U1657 (N_1657,N_582,N_698);
or U1658 (N_1658,N_711,N_586);
and U1659 (N_1659,N_607,N_642);
and U1660 (N_1660,N_277,N_157);
nor U1661 (N_1661,N_608,N_447);
nor U1662 (N_1662,N_596,N_621);
and U1663 (N_1663,N_932,N_357);
or U1664 (N_1664,N_710,N_83);
nor U1665 (N_1665,N_539,N_775);
nand U1666 (N_1666,N_75,N_370);
nor U1667 (N_1667,N_284,N_566);
and U1668 (N_1668,N_381,N_74);
or U1669 (N_1669,N_423,N_211);
or U1670 (N_1670,N_933,N_436);
and U1671 (N_1671,N_623,N_717);
and U1672 (N_1672,N_854,N_114);
nand U1673 (N_1673,N_906,N_468);
nand U1674 (N_1674,N_496,N_858);
nand U1675 (N_1675,N_369,N_956);
and U1676 (N_1676,N_69,N_430);
and U1677 (N_1677,N_558,N_649);
and U1678 (N_1678,N_493,N_580);
or U1679 (N_1679,N_347,N_778);
and U1680 (N_1680,N_910,N_251);
or U1681 (N_1681,N_795,N_820);
or U1682 (N_1682,N_833,N_619);
nand U1683 (N_1683,N_395,N_884);
or U1684 (N_1684,N_914,N_578);
or U1685 (N_1685,N_984,N_408);
and U1686 (N_1686,N_36,N_934);
or U1687 (N_1687,N_7,N_587);
and U1688 (N_1688,N_879,N_677);
and U1689 (N_1689,N_174,N_73);
or U1690 (N_1690,N_333,N_661);
or U1691 (N_1691,N_740,N_500);
and U1692 (N_1692,N_348,N_234);
and U1693 (N_1693,N_716,N_197);
nor U1694 (N_1694,N_98,N_622);
and U1695 (N_1695,N_603,N_91);
nor U1696 (N_1696,N_147,N_237);
and U1697 (N_1697,N_433,N_145);
nor U1698 (N_1698,N_69,N_414);
or U1699 (N_1699,N_337,N_196);
and U1700 (N_1700,N_509,N_415);
and U1701 (N_1701,N_249,N_0);
nand U1702 (N_1702,N_660,N_257);
and U1703 (N_1703,N_757,N_652);
and U1704 (N_1704,N_178,N_63);
nor U1705 (N_1705,N_39,N_602);
or U1706 (N_1706,N_752,N_976);
and U1707 (N_1707,N_376,N_846);
or U1708 (N_1708,N_343,N_67);
and U1709 (N_1709,N_757,N_402);
or U1710 (N_1710,N_52,N_225);
or U1711 (N_1711,N_251,N_814);
or U1712 (N_1712,N_724,N_548);
and U1713 (N_1713,N_49,N_448);
and U1714 (N_1714,N_732,N_765);
or U1715 (N_1715,N_825,N_696);
or U1716 (N_1716,N_430,N_763);
and U1717 (N_1717,N_528,N_758);
nor U1718 (N_1718,N_355,N_4);
and U1719 (N_1719,N_76,N_151);
nand U1720 (N_1720,N_149,N_177);
and U1721 (N_1721,N_257,N_569);
and U1722 (N_1722,N_168,N_963);
nand U1723 (N_1723,N_268,N_454);
nand U1724 (N_1724,N_811,N_128);
xnor U1725 (N_1725,N_740,N_267);
nor U1726 (N_1726,N_180,N_929);
and U1727 (N_1727,N_613,N_45);
or U1728 (N_1728,N_302,N_555);
or U1729 (N_1729,N_480,N_905);
nand U1730 (N_1730,N_310,N_972);
or U1731 (N_1731,N_846,N_201);
or U1732 (N_1732,N_865,N_521);
and U1733 (N_1733,N_224,N_518);
and U1734 (N_1734,N_744,N_337);
or U1735 (N_1735,N_771,N_657);
nand U1736 (N_1736,N_733,N_178);
nand U1737 (N_1737,N_137,N_799);
nand U1738 (N_1738,N_847,N_801);
nor U1739 (N_1739,N_354,N_168);
or U1740 (N_1740,N_694,N_691);
and U1741 (N_1741,N_698,N_563);
or U1742 (N_1742,N_501,N_858);
and U1743 (N_1743,N_99,N_337);
or U1744 (N_1744,N_512,N_115);
and U1745 (N_1745,N_217,N_814);
and U1746 (N_1746,N_997,N_274);
nor U1747 (N_1747,N_318,N_232);
or U1748 (N_1748,N_142,N_366);
nand U1749 (N_1749,N_660,N_867);
nand U1750 (N_1750,N_156,N_991);
nor U1751 (N_1751,N_581,N_487);
nor U1752 (N_1752,N_443,N_983);
or U1753 (N_1753,N_103,N_431);
nand U1754 (N_1754,N_803,N_97);
or U1755 (N_1755,N_592,N_638);
nand U1756 (N_1756,N_475,N_890);
nand U1757 (N_1757,N_2,N_839);
or U1758 (N_1758,N_589,N_573);
nor U1759 (N_1759,N_619,N_197);
nand U1760 (N_1760,N_509,N_822);
and U1761 (N_1761,N_634,N_112);
nor U1762 (N_1762,N_229,N_384);
xnor U1763 (N_1763,N_620,N_62);
nor U1764 (N_1764,N_461,N_58);
and U1765 (N_1765,N_359,N_257);
nor U1766 (N_1766,N_516,N_203);
or U1767 (N_1767,N_582,N_428);
or U1768 (N_1768,N_38,N_782);
nor U1769 (N_1769,N_444,N_239);
nand U1770 (N_1770,N_77,N_819);
or U1771 (N_1771,N_70,N_335);
or U1772 (N_1772,N_21,N_38);
nand U1773 (N_1773,N_499,N_850);
and U1774 (N_1774,N_903,N_89);
nor U1775 (N_1775,N_598,N_82);
and U1776 (N_1776,N_680,N_244);
and U1777 (N_1777,N_577,N_966);
nor U1778 (N_1778,N_774,N_767);
nand U1779 (N_1779,N_881,N_896);
nand U1780 (N_1780,N_873,N_879);
or U1781 (N_1781,N_219,N_420);
or U1782 (N_1782,N_253,N_577);
nor U1783 (N_1783,N_631,N_279);
nor U1784 (N_1784,N_783,N_87);
nor U1785 (N_1785,N_825,N_846);
nor U1786 (N_1786,N_799,N_484);
nor U1787 (N_1787,N_875,N_916);
nor U1788 (N_1788,N_698,N_990);
nor U1789 (N_1789,N_73,N_930);
or U1790 (N_1790,N_235,N_722);
nand U1791 (N_1791,N_396,N_792);
nor U1792 (N_1792,N_816,N_274);
nor U1793 (N_1793,N_290,N_502);
nor U1794 (N_1794,N_194,N_62);
nor U1795 (N_1795,N_90,N_568);
or U1796 (N_1796,N_222,N_755);
nand U1797 (N_1797,N_160,N_749);
or U1798 (N_1798,N_266,N_594);
nand U1799 (N_1799,N_926,N_410);
nand U1800 (N_1800,N_296,N_434);
or U1801 (N_1801,N_179,N_441);
nor U1802 (N_1802,N_881,N_907);
nor U1803 (N_1803,N_59,N_930);
or U1804 (N_1804,N_416,N_508);
or U1805 (N_1805,N_971,N_574);
nor U1806 (N_1806,N_385,N_809);
and U1807 (N_1807,N_765,N_763);
or U1808 (N_1808,N_817,N_581);
or U1809 (N_1809,N_827,N_358);
and U1810 (N_1810,N_114,N_588);
nand U1811 (N_1811,N_123,N_71);
nor U1812 (N_1812,N_610,N_438);
nor U1813 (N_1813,N_84,N_244);
or U1814 (N_1814,N_81,N_666);
and U1815 (N_1815,N_511,N_465);
and U1816 (N_1816,N_349,N_671);
or U1817 (N_1817,N_624,N_76);
nor U1818 (N_1818,N_333,N_853);
nor U1819 (N_1819,N_937,N_37);
nand U1820 (N_1820,N_810,N_938);
or U1821 (N_1821,N_491,N_699);
or U1822 (N_1822,N_287,N_406);
nand U1823 (N_1823,N_456,N_232);
and U1824 (N_1824,N_338,N_976);
and U1825 (N_1825,N_194,N_109);
and U1826 (N_1826,N_939,N_45);
nand U1827 (N_1827,N_268,N_206);
and U1828 (N_1828,N_993,N_22);
and U1829 (N_1829,N_753,N_288);
or U1830 (N_1830,N_809,N_816);
and U1831 (N_1831,N_507,N_756);
nor U1832 (N_1832,N_444,N_331);
and U1833 (N_1833,N_843,N_59);
or U1834 (N_1834,N_968,N_532);
or U1835 (N_1835,N_577,N_615);
or U1836 (N_1836,N_317,N_261);
nand U1837 (N_1837,N_795,N_619);
and U1838 (N_1838,N_555,N_585);
or U1839 (N_1839,N_649,N_11);
nor U1840 (N_1840,N_789,N_884);
nor U1841 (N_1841,N_777,N_269);
nand U1842 (N_1842,N_451,N_406);
nand U1843 (N_1843,N_145,N_451);
and U1844 (N_1844,N_834,N_410);
or U1845 (N_1845,N_255,N_909);
nand U1846 (N_1846,N_222,N_474);
nand U1847 (N_1847,N_657,N_886);
and U1848 (N_1848,N_838,N_6);
and U1849 (N_1849,N_194,N_985);
nand U1850 (N_1850,N_300,N_635);
or U1851 (N_1851,N_242,N_843);
or U1852 (N_1852,N_634,N_478);
and U1853 (N_1853,N_238,N_897);
nor U1854 (N_1854,N_221,N_704);
nor U1855 (N_1855,N_286,N_316);
nor U1856 (N_1856,N_401,N_492);
and U1857 (N_1857,N_95,N_450);
and U1858 (N_1858,N_572,N_499);
nand U1859 (N_1859,N_548,N_871);
nor U1860 (N_1860,N_313,N_821);
or U1861 (N_1861,N_428,N_167);
or U1862 (N_1862,N_245,N_470);
nand U1863 (N_1863,N_875,N_755);
nor U1864 (N_1864,N_569,N_880);
or U1865 (N_1865,N_393,N_806);
or U1866 (N_1866,N_579,N_865);
or U1867 (N_1867,N_918,N_663);
nand U1868 (N_1868,N_731,N_435);
or U1869 (N_1869,N_936,N_789);
nor U1870 (N_1870,N_861,N_775);
and U1871 (N_1871,N_161,N_707);
nor U1872 (N_1872,N_134,N_453);
and U1873 (N_1873,N_269,N_1);
or U1874 (N_1874,N_213,N_289);
and U1875 (N_1875,N_900,N_282);
and U1876 (N_1876,N_792,N_346);
or U1877 (N_1877,N_25,N_868);
nand U1878 (N_1878,N_566,N_404);
or U1879 (N_1879,N_243,N_735);
or U1880 (N_1880,N_952,N_461);
or U1881 (N_1881,N_811,N_932);
or U1882 (N_1882,N_461,N_13);
nand U1883 (N_1883,N_871,N_572);
and U1884 (N_1884,N_454,N_420);
or U1885 (N_1885,N_1,N_261);
and U1886 (N_1886,N_190,N_63);
and U1887 (N_1887,N_846,N_334);
and U1888 (N_1888,N_972,N_381);
or U1889 (N_1889,N_46,N_561);
nor U1890 (N_1890,N_945,N_982);
and U1891 (N_1891,N_649,N_341);
and U1892 (N_1892,N_90,N_723);
or U1893 (N_1893,N_636,N_221);
or U1894 (N_1894,N_326,N_486);
and U1895 (N_1895,N_443,N_602);
nor U1896 (N_1896,N_898,N_817);
or U1897 (N_1897,N_144,N_40);
or U1898 (N_1898,N_127,N_525);
nand U1899 (N_1899,N_60,N_482);
nand U1900 (N_1900,N_130,N_560);
nor U1901 (N_1901,N_782,N_387);
nand U1902 (N_1902,N_292,N_81);
nor U1903 (N_1903,N_739,N_855);
nor U1904 (N_1904,N_644,N_798);
and U1905 (N_1905,N_319,N_361);
or U1906 (N_1906,N_555,N_885);
nand U1907 (N_1907,N_523,N_769);
nor U1908 (N_1908,N_732,N_370);
nand U1909 (N_1909,N_962,N_853);
and U1910 (N_1910,N_215,N_387);
nor U1911 (N_1911,N_380,N_96);
or U1912 (N_1912,N_894,N_430);
and U1913 (N_1913,N_954,N_426);
nand U1914 (N_1914,N_398,N_652);
and U1915 (N_1915,N_626,N_77);
or U1916 (N_1916,N_711,N_119);
nor U1917 (N_1917,N_501,N_132);
or U1918 (N_1918,N_622,N_115);
or U1919 (N_1919,N_618,N_758);
nor U1920 (N_1920,N_649,N_989);
nor U1921 (N_1921,N_202,N_34);
and U1922 (N_1922,N_217,N_947);
nor U1923 (N_1923,N_694,N_875);
and U1924 (N_1924,N_642,N_193);
nor U1925 (N_1925,N_76,N_793);
nand U1926 (N_1926,N_597,N_881);
or U1927 (N_1927,N_745,N_545);
nand U1928 (N_1928,N_896,N_746);
nor U1929 (N_1929,N_302,N_211);
and U1930 (N_1930,N_571,N_857);
or U1931 (N_1931,N_886,N_170);
and U1932 (N_1932,N_932,N_472);
and U1933 (N_1933,N_359,N_350);
nor U1934 (N_1934,N_631,N_757);
nor U1935 (N_1935,N_243,N_971);
nand U1936 (N_1936,N_465,N_223);
nand U1937 (N_1937,N_296,N_650);
and U1938 (N_1938,N_611,N_87);
and U1939 (N_1939,N_115,N_770);
nand U1940 (N_1940,N_20,N_690);
or U1941 (N_1941,N_474,N_98);
or U1942 (N_1942,N_150,N_283);
nor U1943 (N_1943,N_869,N_748);
nand U1944 (N_1944,N_981,N_571);
or U1945 (N_1945,N_65,N_713);
nand U1946 (N_1946,N_903,N_377);
nor U1947 (N_1947,N_441,N_368);
or U1948 (N_1948,N_734,N_890);
nand U1949 (N_1949,N_563,N_691);
nor U1950 (N_1950,N_765,N_927);
or U1951 (N_1951,N_924,N_56);
nor U1952 (N_1952,N_89,N_144);
nor U1953 (N_1953,N_432,N_204);
nand U1954 (N_1954,N_967,N_864);
and U1955 (N_1955,N_592,N_170);
and U1956 (N_1956,N_971,N_230);
nor U1957 (N_1957,N_396,N_405);
nor U1958 (N_1958,N_611,N_448);
or U1959 (N_1959,N_759,N_731);
or U1960 (N_1960,N_120,N_664);
nand U1961 (N_1961,N_948,N_270);
nand U1962 (N_1962,N_100,N_432);
or U1963 (N_1963,N_250,N_779);
or U1964 (N_1964,N_254,N_120);
nor U1965 (N_1965,N_828,N_465);
nand U1966 (N_1966,N_796,N_627);
or U1967 (N_1967,N_359,N_292);
or U1968 (N_1968,N_993,N_29);
nand U1969 (N_1969,N_974,N_404);
or U1970 (N_1970,N_198,N_573);
nor U1971 (N_1971,N_543,N_22);
nand U1972 (N_1972,N_558,N_213);
or U1973 (N_1973,N_440,N_447);
nand U1974 (N_1974,N_398,N_775);
and U1975 (N_1975,N_902,N_900);
or U1976 (N_1976,N_566,N_637);
xor U1977 (N_1977,N_656,N_212);
nand U1978 (N_1978,N_362,N_919);
nand U1979 (N_1979,N_356,N_141);
or U1980 (N_1980,N_554,N_836);
nor U1981 (N_1981,N_706,N_185);
nor U1982 (N_1982,N_480,N_737);
and U1983 (N_1983,N_856,N_736);
or U1984 (N_1984,N_474,N_388);
nand U1985 (N_1985,N_152,N_955);
nor U1986 (N_1986,N_108,N_59);
nor U1987 (N_1987,N_879,N_392);
or U1988 (N_1988,N_761,N_495);
nor U1989 (N_1989,N_287,N_135);
or U1990 (N_1990,N_96,N_734);
nand U1991 (N_1991,N_698,N_268);
or U1992 (N_1992,N_996,N_16);
or U1993 (N_1993,N_9,N_487);
and U1994 (N_1994,N_606,N_714);
nand U1995 (N_1995,N_110,N_866);
or U1996 (N_1996,N_724,N_25);
or U1997 (N_1997,N_946,N_60);
and U1998 (N_1998,N_667,N_565);
and U1999 (N_1999,N_632,N_362);
or U2000 (N_2000,N_1244,N_1000);
nand U2001 (N_2001,N_1621,N_1345);
nor U2002 (N_2002,N_1236,N_1303);
xor U2003 (N_2003,N_1147,N_1466);
nor U2004 (N_2004,N_1554,N_1170);
nand U2005 (N_2005,N_1262,N_1094);
and U2006 (N_2006,N_1580,N_1652);
nand U2007 (N_2007,N_1898,N_1003);
nand U2008 (N_2008,N_1773,N_1548);
nor U2009 (N_2009,N_1245,N_1635);
or U2010 (N_2010,N_1662,N_1659);
nand U2011 (N_2011,N_1095,N_1622);
or U2012 (N_2012,N_1744,N_1311);
nor U2013 (N_2013,N_1098,N_1721);
and U2014 (N_2014,N_1775,N_1061);
nor U2015 (N_2015,N_1418,N_1038);
or U2016 (N_2016,N_1473,N_1544);
xnor U2017 (N_2017,N_1745,N_1588);
or U2018 (N_2018,N_1288,N_1162);
and U2019 (N_2019,N_1277,N_1546);
nand U2020 (N_2020,N_1292,N_1742);
or U2021 (N_2021,N_1612,N_1065);
or U2022 (N_2022,N_1282,N_1016);
or U2023 (N_2023,N_1856,N_1710);
and U2024 (N_2024,N_1354,N_1063);
nand U2025 (N_2025,N_1294,N_1753);
and U2026 (N_2026,N_1736,N_1519);
nor U2027 (N_2027,N_1238,N_1986);
and U2028 (N_2028,N_1416,N_1194);
xnor U2029 (N_2029,N_1728,N_1117);
or U2030 (N_2030,N_1924,N_1599);
nor U2031 (N_2031,N_1844,N_1078);
nor U2032 (N_2032,N_1070,N_1725);
nand U2033 (N_2033,N_1700,N_1112);
nand U2034 (N_2034,N_1819,N_1536);
or U2035 (N_2035,N_1730,N_1961);
or U2036 (N_2036,N_1571,N_1712);
or U2037 (N_2037,N_1793,N_1255);
or U2038 (N_2038,N_1584,N_1209);
or U2039 (N_2039,N_1709,N_1456);
and U2040 (N_2040,N_1022,N_1792);
nor U2041 (N_2041,N_1057,N_1796);
or U2042 (N_2042,N_1441,N_1368);
nor U2043 (N_2043,N_1115,N_1103);
nor U2044 (N_2044,N_1758,N_1278);
nand U2045 (N_2045,N_1422,N_1333);
and U2046 (N_2046,N_1099,N_1729);
or U2047 (N_2047,N_1188,N_1568);
and U2048 (N_2048,N_1026,N_1495);
nand U2049 (N_2049,N_1727,N_1297);
or U2050 (N_2050,N_1668,N_1577);
or U2051 (N_2051,N_1109,N_1910);
or U2052 (N_2052,N_1797,N_1380);
or U2053 (N_2053,N_1015,N_1781);
xor U2054 (N_2054,N_1952,N_1951);
or U2055 (N_2055,N_1020,N_1293);
and U2056 (N_2056,N_1077,N_1633);
and U2057 (N_2057,N_1152,N_1896);
or U2058 (N_2058,N_1769,N_1595);
nor U2059 (N_2059,N_1539,N_1248);
nor U2060 (N_2060,N_1252,N_1576);
nand U2061 (N_2061,N_1649,N_1053);
and U2062 (N_2062,N_1586,N_1686);
and U2063 (N_2063,N_1346,N_1446);
and U2064 (N_2064,N_1613,N_1179);
or U2065 (N_2065,N_1004,N_1861);
and U2066 (N_2066,N_1363,N_1189);
and U2067 (N_2067,N_1069,N_1153);
nor U2068 (N_2068,N_1562,N_1071);
or U2069 (N_2069,N_1629,N_1764);
nor U2070 (N_2070,N_1342,N_1934);
or U2071 (N_2071,N_1041,N_1430);
nand U2072 (N_2072,N_1178,N_1538);
nand U2073 (N_2073,N_1223,N_1500);
and U2074 (N_2074,N_1884,N_1999);
and U2075 (N_2075,N_1225,N_1645);
nand U2076 (N_2076,N_1677,N_1981);
and U2077 (N_2077,N_1206,N_1185);
nor U2078 (N_2078,N_1018,N_1085);
or U2079 (N_2079,N_1658,N_1062);
xnor U2080 (N_2080,N_1468,N_1828);
and U2081 (N_2081,N_1163,N_1589);
or U2082 (N_2082,N_1391,N_1770);
nor U2083 (N_2083,N_1478,N_1328);
nand U2084 (N_2084,N_1337,N_1143);
nand U2085 (N_2085,N_1883,N_1044);
and U2086 (N_2086,N_1506,N_1674);
and U2087 (N_2087,N_1798,N_1642);
nand U2088 (N_2088,N_1290,N_1196);
nor U2089 (N_2089,N_1955,N_1173);
nand U2090 (N_2090,N_1509,N_1265);
nand U2091 (N_2091,N_1033,N_1558);
or U2092 (N_2092,N_1937,N_1369);
or U2093 (N_2093,N_1208,N_1904);
or U2094 (N_2094,N_1240,N_1776);
and U2095 (N_2095,N_1315,N_1286);
nor U2096 (N_2096,N_1648,N_1512);
and U2097 (N_2097,N_1474,N_1624);
nor U2098 (N_2098,N_1203,N_1080);
and U2099 (N_2099,N_1481,N_1615);
and U2100 (N_2100,N_1911,N_1606);
or U2101 (N_2101,N_1372,N_1161);
and U2102 (N_2102,N_1426,N_1234);
or U2103 (N_2103,N_1281,N_1526);
nand U2104 (N_2104,N_1198,N_1367);
nand U2105 (N_2105,N_1988,N_1936);
and U2106 (N_2106,N_1148,N_1276);
nand U2107 (N_2107,N_1854,N_1992);
and U2108 (N_2108,N_1551,N_1533);
or U2109 (N_2109,N_1722,N_1912);
or U2110 (N_2110,N_1650,N_1582);
and U2111 (N_2111,N_1024,N_1905);
or U2112 (N_2112,N_1895,N_1157);
nor U2113 (N_2113,N_1267,N_1572);
or U2114 (N_2114,N_1154,N_1614);
nand U2115 (N_2115,N_1806,N_1717);
nor U2116 (N_2116,N_1435,N_1308);
nand U2117 (N_2117,N_1210,N_1687);
and U2118 (N_2118,N_1241,N_1738);
nor U2119 (N_2119,N_1860,N_1283);
nand U2120 (N_2120,N_1944,N_1480);
nor U2121 (N_2121,N_1270,N_1151);
and U2122 (N_2122,N_1406,N_1023);
and U2123 (N_2123,N_1839,N_1043);
and U2124 (N_2124,N_1908,N_1104);
and U2125 (N_2125,N_1397,N_1039);
and U2126 (N_2126,N_1857,N_1442);
nand U2127 (N_2127,N_1731,N_1461);
and U2128 (N_2128,N_1132,N_1974);
nor U2129 (N_2129,N_1953,N_1029);
and U2130 (N_2130,N_1697,N_1508);
nor U2131 (N_2131,N_1475,N_1213);
or U2132 (N_2132,N_1381,N_1131);
and U2133 (N_2133,N_1049,N_1619);
or U2134 (N_2134,N_1465,N_1723);
and U2135 (N_2135,N_1171,N_1802);
or U2136 (N_2136,N_1691,N_1079);
and U2137 (N_2137,N_1518,N_1529);
or U2138 (N_2138,N_1013,N_1880);
or U2139 (N_2139,N_1399,N_1682);
and U2140 (N_2140,N_1946,N_1176);
nor U2141 (N_2141,N_1761,N_1532);
and U2142 (N_2142,N_1027,N_1505);
or U2143 (N_2143,N_1829,N_1479);
and U2144 (N_2144,N_1256,N_1300);
and U2145 (N_2145,N_1611,N_1909);
or U2146 (N_2146,N_1317,N_1965);
nand U2147 (N_2147,N_1765,N_1984);
nand U2148 (N_2148,N_1754,N_1204);
or U2149 (N_2149,N_1125,N_1740);
nand U2150 (N_2150,N_1921,N_1821);
nand U2151 (N_2151,N_1343,N_1415);
or U2152 (N_2152,N_1216,N_1136);
nor U2153 (N_2153,N_1289,N_1597);
nor U2154 (N_2154,N_1890,N_1105);
and U2155 (N_2155,N_1864,N_1124);
nor U2156 (N_2156,N_1493,N_1340);
nand U2157 (N_2157,N_1195,N_1811);
nor U2158 (N_2158,N_1784,N_1219);
nor U2159 (N_2159,N_1634,N_1454);
and U2160 (N_2160,N_1871,N_1111);
nor U2161 (N_2161,N_1777,N_1523);
and U2162 (N_2162,N_1222,N_1110);
or U2163 (N_2163,N_1427,N_1149);
nor U2164 (N_2164,N_1230,N_1034);
and U2165 (N_2165,N_1824,N_1812);
nand U2166 (N_2166,N_1593,N_1200);
and U2167 (N_2167,N_1378,N_1836);
or U2168 (N_2168,N_1075,N_1675);
and U2169 (N_2169,N_1434,N_1226);
nor U2170 (N_2170,N_1414,N_1395);
and U2171 (N_2171,N_1128,N_1307);
and U2172 (N_2172,N_1967,N_1669);
and U2173 (N_2173,N_1835,N_1233);
and U2174 (N_2174,N_1167,N_1541);
and U2175 (N_2175,N_1032,N_1068);
nor U2176 (N_2176,N_1483,N_1302);
nor U2177 (N_2177,N_1771,N_1915);
and U2178 (N_2178,N_1334,N_1701);
nand U2179 (N_2179,N_1638,N_1684);
nand U2180 (N_2180,N_1849,N_1632);
nor U2181 (N_2181,N_1431,N_1888);
nand U2182 (N_2182,N_1799,N_1703);
nand U2183 (N_2183,N_1165,N_1366);
nor U2184 (N_2184,N_1177,N_1005);
and U2185 (N_2185,N_1371,N_1827);
or U2186 (N_2186,N_1779,N_1246);
nand U2187 (N_2187,N_1940,N_1833);
or U2188 (N_2188,N_1596,N_1263);
or U2189 (N_2189,N_1920,N_1386);
nand U2190 (N_2190,N_1808,N_1129);
and U2191 (N_2191,N_1834,N_1993);
and U2192 (N_2192,N_1467,N_1492);
nor U2193 (N_2193,N_1362,N_1159);
nand U2194 (N_2194,N_1756,N_1287);
nor U2195 (N_2195,N_1600,N_1045);
nor U2196 (N_2196,N_1983,N_1463);
and U2197 (N_2197,N_1377,N_1275);
and U2198 (N_2198,N_1997,N_1193);
or U2199 (N_2199,N_1818,N_1370);
nand U2200 (N_2200,N_1229,N_1978);
or U2201 (N_2201,N_1119,N_1690);
or U2202 (N_2202,N_1626,N_1011);
nand U2203 (N_2203,N_1862,N_1891);
nand U2204 (N_2204,N_1301,N_1810);
or U2205 (N_2205,N_1348,N_1349);
and U2206 (N_2206,N_1549,N_1733);
or U2207 (N_2207,N_1396,N_1579);
nand U2208 (N_2208,N_1212,N_1017);
nor U2209 (N_2209,N_1254,N_1585);
xnor U2210 (N_2210,N_1423,N_1329);
or U2211 (N_2211,N_1553,N_1943);
nand U2212 (N_2212,N_1323,N_1258);
and U2213 (N_2213,N_1875,N_1976);
nor U2214 (N_2214,N_1358,N_1498);
nand U2215 (N_2215,N_1928,N_1006);
or U2216 (N_2216,N_1139,N_1575);
and U2217 (N_2217,N_1106,N_1874);
nand U2218 (N_2218,N_1066,N_1172);
nand U2219 (N_2219,N_1059,N_1141);
or U2220 (N_2220,N_1168,N_1021);
nor U2221 (N_2221,N_1716,N_1628);
and U2222 (N_2222,N_1192,N_1557);
nand U2223 (N_2223,N_1429,N_1778);
nand U2224 (N_2224,N_1647,N_1605);
and U2225 (N_2225,N_1878,N_1393);
nor U2226 (N_2226,N_1900,N_1356);
nor U2227 (N_2227,N_1118,N_1948);
nor U2228 (N_2228,N_1001,N_1108);
or U2229 (N_2229,N_1930,N_1237);
or U2230 (N_2230,N_1607,N_1973);
and U2231 (N_2231,N_1931,N_1046);
nor U2232 (N_2232,N_1201,N_1299);
nand U2233 (N_2233,N_1664,N_1067);
nor U2234 (N_2234,N_1432,N_1603);
and U2235 (N_2235,N_1268,N_1653);
nand U2236 (N_2236,N_1504,N_1848);
and U2237 (N_2237,N_1766,N_1113);
nor U2238 (N_2238,N_1402,N_1250);
and U2239 (N_2239,N_1975,N_1608);
nand U2240 (N_2240,N_1350,N_1971);
or U2241 (N_2241,N_1452,N_1641);
nand U2242 (N_2242,N_1567,N_1962);
and U2243 (N_2243,N_1540,N_1130);
or U2244 (N_2244,N_1655,N_1637);
or U2245 (N_2245,N_1906,N_1590);
or U2246 (N_2246,N_1313,N_1954);
or U2247 (N_2247,N_1528,N_1747);
nor U2248 (N_2248,N_1511,N_1903);
nand U2249 (N_2249,N_1991,N_1403);
and U2250 (N_2250,N_1737,N_1138);
and U2251 (N_2251,N_1866,N_1160);
nand U2252 (N_2252,N_1760,N_1449);
or U2253 (N_2253,N_1321,N_1676);
and U2254 (N_2254,N_1251,N_1227);
nor U2255 (N_2255,N_1530,N_1873);
or U2256 (N_2256,N_1374,N_1566);
or U2257 (N_2257,N_1460,N_1385);
and U2258 (N_2258,N_1767,N_1521);
nand U2259 (N_2259,N_1060,N_1035);
nand U2260 (N_2260,N_1344,N_1469);
nor U2261 (N_2261,N_1056,N_1872);
nor U2262 (N_2262,N_1296,N_1715);
and U2263 (N_2263,N_1072,N_1081);
and U2264 (N_2264,N_1330,N_1096);
and U2265 (N_2265,N_1907,N_1837);
nor U2266 (N_2266,N_1899,N_1639);
or U2267 (N_2267,N_1054,N_1651);
nor U2268 (N_2268,N_1893,N_1145);
and U2269 (N_2269,N_1400,N_1092);
nor U2270 (N_2270,N_1507,N_1527);
nor U2271 (N_2271,N_1604,N_1887);
nand U2272 (N_2272,N_1671,N_1926);
and U2273 (N_2273,N_1394,N_1850);
xor U2274 (N_2274,N_1260,N_1089);
or U2275 (N_2275,N_1249,N_1324);
or U2276 (N_2276,N_1428,N_1123);
and U2277 (N_2277,N_1574,N_1869);
nand U2278 (N_2278,N_1643,N_1247);
nand U2279 (N_2279,N_1014,N_1679);
and U2280 (N_2280,N_1851,N_1790);
or U2281 (N_2281,N_1885,N_1542);
nand U2282 (N_2282,N_1718,N_1450);
nor U2283 (N_2283,N_1304,N_1365);
or U2284 (N_2284,N_1325,N_1996);
nor U2285 (N_2285,N_1922,N_1879);
or U2286 (N_2286,N_1413,N_1025);
or U2287 (N_2287,N_1318,N_1407);
or U2288 (N_2288,N_1217,N_1259);
nand U2289 (N_2289,N_1867,N_1815);
and U2290 (N_2290,N_1097,N_1735);
nor U2291 (N_2291,N_1338,N_1933);
and U2292 (N_2292,N_1578,N_1285);
nor U2293 (N_2293,N_1088,N_1444);
and U2294 (N_2294,N_1932,N_1617);
xor U2295 (N_2295,N_1694,N_1990);
nand U2296 (N_2296,N_1535,N_1257);
nand U2297 (N_2297,N_1140,N_1995);
or U2298 (N_2298,N_1487,N_1019);
and U2299 (N_2299,N_1826,N_1914);
or U2300 (N_2300,N_1295,N_1090);
nor U2301 (N_2301,N_1919,N_1424);
and U2302 (N_2302,N_1845,N_1670);
or U2303 (N_2303,N_1490,N_1312);
and U2304 (N_2304,N_1355,N_1859);
nor U2305 (N_2305,N_1620,N_1284);
or U2306 (N_2306,N_1524,N_1375);
nor U2307 (N_2307,N_1847,N_1726);
or U2308 (N_2308,N_1392,N_1142);
nor U2309 (N_2309,N_1306,N_1436);
nor U2310 (N_2310,N_1804,N_1009);
nand U2311 (N_2311,N_1925,N_1187);
nand U2312 (N_2312,N_1998,N_1309);
nor U2313 (N_2313,N_1618,N_1685);
nor U2314 (N_2314,N_1357,N_1447);
and U2315 (N_2315,N_1417,N_1264);
nand U2316 (N_2316,N_1387,N_1144);
nor U2317 (N_2317,N_1786,N_1291);
nor U2318 (N_2318,N_1752,N_1482);
nor U2319 (N_2319,N_1841,N_1221);
or U2320 (N_2320,N_1556,N_1616);
nand U2321 (N_2321,N_1977,N_1666);
and U2322 (N_2322,N_1445,N_1681);
nor U2323 (N_2323,N_1660,N_1379);
and U2324 (N_2324,N_1091,N_1352);
nand U2325 (N_2325,N_1947,N_1863);
nand U2326 (N_2326,N_1412,N_1842);
and U2327 (N_2327,N_1133,N_1084);
nor U2328 (N_2328,N_1763,N_1801);
and U2329 (N_2329,N_1074,N_1007);
nand U2330 (N_2330,N_1458,N_1831);
nand U2331 (N_2331,N_1114,N_1489);
nand U2332 (N_2332,N_1082,N_1843);
nor U2333 (N_2333,N_1601,N_1280);
nor U2334 (N_2334,N_1497,N_1002);
and U2335 (N_2335,N_1705,N_1031);
nor U2336 (N_2336,N_1503,N_1155);
and U2337 (N_2337,N_1499,N_1186);
or U2338 (N_2338,N_1076,N_1935);
or U2339 (N_2339,N_1332,N_1699);
or U2340 (N_2340,N_1419,N_1724);
nand U2341 (N_2341,N_1484,N_1064);
and U2342 (N_2342,N_1858,N_1459);
and U2343 (N_2343,N_1448,N_1987);
or U2344 (N_2344,N_1741,N_1273);
or U2345 (N_2345,N_1817,N_1772);
and U2346 (N_2346,N_1305,N_1120);
and U2347 (N_2347,N_1166,N_1689);
nor U2348 (N_2348,N_1134,N_1768);
nor U2349 (N_2349,N_1565,N_1780);
and U2350 (N_2350,N_1030,N_1774);
and U2351 (N_2351,N_1175,N_1037);
and U2352 (N_2352,N_1055,N_1814);
and U2353 (N_2353,N_1485,N_1762);
or U2354 (N_2354,N_1364,N_1347);
nand U2355 (N_2355,N_1877,N_1956);
nand U2356 (N_2356,N_1438,N_1457);
and U2357 (N_2357,N_1949,N_1488);
nor U2358 (N_2358,N_1972,N_1537);
nor U2359 (N_2359,N_1327,N_1587);
and U2360 (N_2360,N_1739,N_1361);
nor U2361 (N_2361,N_1522,N_1472);
or U2362 (N_2362,N_1502,N_1274);
and U2363 (N_2363,N_1516,N_1704);
nor U2364 (N_2364,N_1336,N_1547);
and U2365 (N_2365,N_1813,N_1146);
nand U2366 (N_2366,N_1389,N_1310);
or U2367 (N_2367,N_1950,N_1181);
or U2368 (N_2368,N_1594,N_1050);
or U2369 (N_2369,N_1693,N_1501);
nor U2370 (N_2370,N_1750,N_1960);
and U2371 (N_2371,N_1320,N_1359);
and U2372 (N_2372,N_1405,N_1868);
xor U2373 (N_2373,N_1470,N_1107);
or U2374 (N_2374,N_1202,N_1610);
nor U2375 (N_2375,N_1058,N_1443);
nand U2376 (N_2376,N_1351,N_1902);
nand U2377 (N_2377,N_1894,N_1360);
nand U2378 (N_2378,N_1205,N_1809);
nand U2379 (N_2379,N_1627,N_1116);
and U2380 (N_2380,N_1570,N_1787);
and U2381 (N_2381,N_1897,N_1698);
nor U2382 (N_2382,N_1794,N_1326);
nand U2383 (N_2383,N_1820,N_1901);
nand U2384 (N_2384,N_1654,N_1464);
nor U2385 (N_2385,N_1199,N_1609);
and U2386 (N_2386,N_1672,N_1550);
or U2387 (N_2387,N_1087,N_1411);
and U2388 (N_2388,N_1052,N_1822);
nor U2389 (N_2389,N_1319,N_1137);
or U2390 (N_2390,N_1958,N_1917);
or U2391 (N_2391,N_1425,N_1892);
nor U2392 (N_2392,N_1383,N_1959);
or U2393 (N_2393,N_1298,N_1939);
and U2394 (N_2394,N_1657,N_1086);
nand U2395 (N_2395,N_1243,N_1513);
and U2396 (N_2396,N_1942,N_1989);
nand U2397 (N_2397,N_1525,N_1266);
nor U2398 (N_2398,N_1782,N_1688);
or U2399 (N_2399,N_1376,N_1870);
or U2400 (N_2400,N_1830,N_1408);
nand U2401 (N_2401,N_1453,N_1047);
or U2402 (N_2402,N_1127,N_1569);
nor U2403 (N_2403,N_1184,N_1421);
and U2404 (N_2404,N_1439,N_1876);
or U2405 (N_2405,N_1966,N_1695);
and U2406 (N_2406,N_1591,N_1008);
and U2407 (N_2407,N_1390,N_1979);
or U2408 (N_2408,N_1656,N_1126);
and U2409 (N_2409,N_1732,N_1583);
nand U2410 (N_2410,N_1644,N_1825);
nor U2411 (N_2411,N_1331,N_1191);
and U2412 (N_2412,N_1881,N_1757);
and U2413 (N_2413,N_1335,N_1382);
nand U2414 (N_2414,N_1889,N_1759);
or U2415 (N_2415,N_1135,N_1169);
and U2416 (N_2416,N_1673,N_1555);
and U2417 (N_2417,N_1156,N_1713);
nor U2418 (N_2418,N_1783,N_1964);
or U2419 (N_2419,N_1028,N_1093);
or U2420 (N_2420,N_1231,N_1543);
or U2421 (N_2421,N_1945,N_1073);
nand U2422 (N_2422,N_1719,N_1122);
nor U2423 (N_2423,N_1625,N_1040);
or U2424 (N_2424,N_1218,N_1749);
and U2425 (N_2425,N_1755,N_1420);
nor U2426 (N_2426,N_1886,N_1968);
xor U2427 (N_2427,N_1788,N_1224);
or U2428 (N_2428,N_1409,N_1010);
and U2429 (N_2429,N_1846,N_1882);
xor U2430 (N_2430,N_1957,N_1440);
and U2431 (N_2431,N_1314,N_1515);
and U2432 (N_2432,N_1646,N_1197);
nor U2433 (N_2433,N_1471,N_1517);
nor U2434 (N_2434,N_1373,N_1678);
nor U2435 (N_2435,N_1623,N_1398);
or U2436 (N_2436,N_1272,N_1269);
or U2437 (N_2437,N_1228,N_1661);
or U2438 (N_2438,N_1803,N_1969);
nor U2439 (N_2439,N_1602,N_1051);
nor U2440 (N_2440,N_1994,N_1791);
nand U2441 (N_2441,N_1401,N_1707);
nand U2442 (N_2442,N_1663,N_1807);
nand U2443 (N_2443,N_1384,N_1271);
and U2444 (N_2444,N_1561,N_1036);
and U2445 (N_2445,N_1923,N_1496);
or U2446 (N_2446,N_1476,N_1261);
and U2447 (N_2447,N_1789,N_1805);
and U2448 (N_2448,N_1534,N_1491);
and U2449 (N_2449,N_1667,N_1795);
and U2450 (N_2450,N_1631,N_1164);
or U2451 (N_2451,N_1174,N_1215);
nand U2452 (N_2452,N_1980,N_1180);
xor U2453 (N_2453,N_1927,N_1190);
xnor U2454 (N_2454,N_1462,N_1564);
and U2455 (N_2455,N_1982,N_1559);
or U2456 (N_2456,N_1510,N_1838);
and U2457 (N_2457,N_1640,N_1183);
xor U2458 (N_2458,N_1630,N_1832);
or U2459 (N_2459,N_1552,N_1823);
nor U2460 (N_2460,N_1853,N_1816);
nor U2461 (N_2461,N_1865,N_1545);
or U2462 (N_2462,N_1477,N_1214);
xor U2463 (N_2463,N_1102,N_1437);
and U2464 (N_2464,N_1048,N_1692);
and U2465 (N_2465,N_1100,N_1182);
nand U2466 (N_2466,N_1665,N_1696);
nand U2467 (N_2467,N_1339,N_1598);
nand U2468 (N_2468,N_1242,N_1855);
or U2469 (N_2469,N_1388,N_1746);
or U2470 (N_2470,N_1220,N_1012);
nor U2471 (N_2471,N_1680,N_1239);
nand U2472 (N_2472,N_1840,N_1150);
nand U2473 (N_2473,N_1938,N_1232);
nand U2474 (N_2474,N_1573,N_1702);
or U2475 (N_2475,N_1279,N_1207);
nor U2476 (N_2476,N_1963,N_1751);
and U2477 (N_2477,N_1042,N_1520);
and U2478 (N_2478,N_1451,N_1785);
or U2479 (N_2479,N_1985,N_1734);
nand U2480 (N_2480,N_1800,N_1714);
nor U2481 (N_2481,N_1494,N_1711);
or U2482 (N_2482,N_1708,N_1341);
and U2483 (N_2483,N_1253,N_1852);
nand U2484 (N_2484,N_1410,N_1433);
or U2485 (N_2485,N_1211,N_1581);
nand U2486 (N_2486,N_1970,N_1592);
and U2487 (N_2487,N_1101,N_1706);
or U2488 (N_2488,N_1353,N_1560);
nor U2489 (N_2489,N_1913,N_1083);
and U2490 (N_2490,N_1929,N_1316);
nand U2491 (N_2491,N_1531,N_1235);
nand U2492 (N_2492,N_1748,N_1322);
or U2493 (N_2493,N_1720,N_1918);
or U2494 (N_2494,N_1743,N_1455);
nor U2495 (N_2495,N_1941,N_1636);
nor U2496 (N_2496,N_1916,N_1563);
or U2497 (N_2497,N_1514,N_1404);
nand U2498 (N_2498,N_1683,N_1158);
or U2499 (N_2499,N_1486,N_1121);
nand U2500 (N_2500,N_1248,N_1141);
and U2501 (N_2501,N_1677,N_1246);
or U2502 (N_2502,N_1732,N_1035);
and U2503 (N_2503,N_1963,N_1134);
nor U2504 (N_2504,N_1969,N_1570);
and U2505 (N_2505,N_1417,N_1632);
nand U2506 (N_2506,N_1696,N_1718);
and U2507 (N_2507,N_1331,N_1113);
or U2508 (N_2508,N_1242,N_1225);
and U2509 (N_2509,N_1986,N_1295);
nand U2510 (N_2510,N_1186,N_1068);
or U2511 (N_2511,N_1583,N_1669);
or U2512 (N_2512,N_1105,N_1863);
or U2513 (N_2513,N_1632,N_1788);
nor U2514 (N_2514,N_1169,N_1993);
or U2515 (N_2515,N_1333,N_1384);
or U2516 (N_2516,N_1165,N_1190);
nor U2517 (N_2517,N_1360,N_1229);
or U2518 (N_2518,N_1214,N_1603);
nand U2519 (N_2519,N_1258,N_1240);
or U2520 (N_2520,N_1425,N_1522);
and U2521 (N_2521,N_1859,N_1373);
nor U2522 (N_2522,N_1053,N_1595);
nand U2523 (N_2523,N_1032,N_1913);
nand U2524 (N_2524,N_1239,N_1178);
and U2525 (N_2525,N_1810,N_1127);
and U2526 (N_2526,N_1577,N_1952);
nand U2527 (N_2527,N_1805,N_1594);
and U2528 (N_2528,N_1227,N_1379);
nand U2529 (N_2529,N_1630,N_1567);
and U2530 (N_2530,N_1830,N_1406);
and U2531 (N_2531,N_1108,N_1840);
and U2532 (N_2532,N_1420,N_1900);
nor U2533 (N_2533,N_1471,N_1613);
nand U2534 (N_2534,N_1436,N_1655);
or U2535 (N_2535,N_1550,N_1842);
or U2536 (N_2536,N_1608,N_1770);
or U2537 (N_2537,N_1038,N_1397);
nor U2538 (N_2538,N_1090,N_1791);
and U2539 (N_2539,N_1553,N_1550);
and U2540 (N_2540,N_1986,N_1350);
nand U2541 (N_2541,N_1032,N_1668);
nor U2542 (N_2542,N_1323,N_1360);
and U2543 (N_2543,N_1717,N_1246);
or U2544 (N_2544,N_1983,N_1292);
xor U2545 (N_2545,N_1219,N_1338);
or U2546 (N_2546,N_1368,N_1627);
nand U2547 (N_2547,N_1984,N_1590);
nor U2548 (N_2548,N_1242,N_1337);
nor U2549 (N_2549,N_1156,N_1027);
nand U2550 (N_2550,N_1434,N_1053);
nand U2551 (N_2551,N_1544,N_1041);
or U2552 (N_2552,N_1004,N_1407);
nor U2553 (N_2553,N_1079,N_1942);
nand U2554 (N_2554,N_1915,N_1031);
and U2555 (N_2555,N_1171,N_1559);
nand U2556 (N_2556,N_1045,N_1616);
and U2557 (N_2557,N_1605,N_1928);
or U2558 (N_2558,N_1822,N_1781);
nor U2559 (N_2559,N_1628,N_1556);
nor U2560 (N_2560,N_1108,N_1392);
or U2561 (N_2561,N_1987,N_1425);
or U2562 (N_2562,N_1703,N_1213);
and U2563 (N_2563,N_1019,N_1395);
nor U2564 (N_2564,N_1773,N_1458);
nand U2565 (N_2565,N_1134,N_1522);
nand U2566 (N_2566,N_1776,N_1760);
nand U2567 (N_2567,N_1981,N_1970);
and U2568 (N_2568,N_1670,N_1074);
nand U2569 (N_2569,N_1409,N_1087);
and U2570 (N_2570,N_1179,N_1131);
and U2571 (N_2571,N_1739,N_1448);
nor U2572 (N_2572,N_1116,N_1664);
or U2573 (N_2573,N_1316,N_1486);
and U2574 (N_2574,N_1117,N_1883);
or U2575 (N_2575,N_1871,N_1617);
and U2576 (N_2576,N_1092,N_1387);
and U2577 (N_2577,N_1226,N_1814);
and U2578 (N_2578,N_1863,N_1152);
and U2579 (N_2579,N_1813,N_1235);
nor U2580 (N_2580,N_1898,N_1892);
nor U2581 (N_2581,N_1373,N_1978);
nor U2582 (N_2582,N_1148,N_1054);
nand U2583 (N_2583,N_1909,N_1683);
or U2584 (N_2584,N_1686,N_1247);
nand U2585 (N_2585,N_1306,N_1201);
nand U2586 (N_2586,N_1783,N_1527);
nor U2587 (N_2587,N_1687,N_1108);
nand U2588 (N_2588,N_1328,N_1798);
or U2589 (N_2589,N_1497,N_1321);
nand U2590 (N_2590,N_1426,N_1900);
or U2591 (N_2591,N_1083,N_1402);
nand U2592 (N_2592,N_1430,N_1724);
nand U2593 (N_2593,N_1772,N_1447);
and U2594 (N_2594,N_1669,N_1514);
or U2595 (N_2595,N_1143,N_1165);
and U2596 (N_2596,N_1852,N_1633);
or U2597 (N_2597,N_1291,N_1140);
nor U2598 (N_2598,N_1586,N_1524);
nand U2599 (N_2599,N_1886,N_1801);
or U2600 (N_2600,N_1135,N_1084);
or U2601 (N_2601,N_1287,N_1699);
nor U2602 (N_2602,N_1408,N_1215);
nor U2603 (N_2603,N_1229,N_1004);
nand U2604 (N_2604,N_1878,N_1177);
nor U2605 (N_2605,N_1773,N_1902);
and U2606 (N_2606,N_1691,N_1570);
and U2607 (N_2607,N_1442,N_1135);
or U2608 (N_2608,N_1037,N_1410);
nand U2609 (N_2609,N_1688,N_1027);
or U2610 (N_2610,N_1841,N_1616);
nor U2611 (N_2611,N_1664,N_1115);
nand U2612 (N_2612,N_1178,N_1313);
and U2613 (N_2613,N_1155,N_1464);
nand U2614 (N_2614,N_1258,N_1159);
nand U2615 (N_2615,N_1085,N_1463);
nand U2616 (N_2616,N_1055,N_1833);
nand U2617 (N_2617,N_1574,N_1175);
or U2618 (N_2618,N_1505,N_1800);
nand U2619 (N_2619,N_1668,N_1878);
nor U2620 (N_2620,N_1300,N_1463);
xor U2621 (N_2621,N_1295,N_1474);
nand U2622 (N_2622,N_1404,N_1888);
and U2623 (N_2623,N_1227,N_1212);
or U2624 (N_2624,N_1951,N_1905);
nand U2625 (N_2625,N_1499,N_1833);
nor U2626 (N_2626,N_1763,N_1532);
or U2627 (N_2627,N_1718,N_1548);
nor U2628 (N_2628,N_1481,N_1629);
nor U2629 (N_2629,N_1117,N_1247);
and U2630 (N_2630,N_1614,N_1551);
and U2631 (N_2631,N_1683,N_1137);
and U2632 (N_2632,N_1792,N_1721);
or U2633 (N_2633,N_1794,N_1725);
and U2634 (N_2634,N_1294,N_1325);
or U2635 (N_2635,N_1104,N_1075);
nand U2636 (N_2636,N_1086,N_1655);
nand U2637 (N_2637,N_1916,N_1974);
and U2638 (N_2638,N_1979,N_1523);
or U2639 (N_2639,N_1754,N_1543);
and U2640 (N_2640,N_1732,N_1067);
or U2641 (N_2641,N_1599,N_1253);
nor U2642 (N_2642,N_1606,N_1530);
or U2643 (N_2643,N_1454,N_1778);
or U2644 (N_2644,N_1587,N_1700);
nand U2645 (N_2645,N_1587,N_1869);
and U2646 (N_2646,N_1752,N_1578);
nand U2647 (N_2647,N_1043,N_1739);
or U2648 (N_2648,N_1144,N_1291);
and U2649 (N_2649,N_1012,N_1387);
nand U2650 (N_2650,N_1420,N_1748);
nor U2651 (N_2651,N_1836,N_1682);
and U2652 (N_2652,N_1134,N_1472);
nand U2653 (N_2653,N_1007,N_1292);
nand U2654 (N_2654,N_1069,N_1463);
or U2655 (N_2655,N_1056,N_1708);
nor U2656 (N_2656,N_1146,N_1179);
and U2657 (N_2657,N_1886,N_1134);
nand U2658 (N_2658,N_1371,N_1919);
nor U2659 (N_2659,N_1578,N_1083);
xor U2660 (N_2660,N_1027,N_1595);
nand U2661 (N_2661,N_1529,N_1115);
nand U2662 (N_2662,N_1154,N_1945);
nor U2663 (N_2663,N_1746,N_1099);
and U2664 (N_2664,N_1619,N_1985);
nand U2665 (N_2665,N_1700,N_1436);
nand U2666 (N_2666,N_1112,N_1500);
nor U2667 (N_2667,N_1104,N_1550);
nor U2668 (N_2668,N_1229,N_1127);
nand U2669 (N_2669,N_1102,N_1157);
and U2670 (N_2670,N_1888,N_1491);
and U2671 (N_2671,N_1032,N_1410);
nor U2672 (N_2672,N_1169,N_1195);
nor U2673 (N_2673,N_1611,N_1501);
and U2674 (N_2674,N_1358,N_1389);
or U2675 (N_2675,N_1611,N_1763);
nor U2676 (N_2676,N_1219,N_1242);
and U2677 (N_2677,N_1885,N_1764);
and U2678 (N_2678,N_1249,N_1836);
or U2679 (N_2679,N_1121,N_1043);
nand U2680 (N_2680,N_1163,N_1890);
or U2681 (N_2681,N_1637,N_1548);
and U2682 (N_2682,N_1818,N_1992);
and U2683 (N_2683,N_1086,N_1520);
nand U2684 (N_2684,N_1160,N_1754);
or U2685 (N_2685,N_1362,N_1781);
and U2686 (N_2686,N_1135,N_1944);
nand U2687 (N_2687,N_1234,N_1525);
and U2688 (N_2688,N_1362,N_1060);
nand U2689 (N_2689,N_1479,N_1495);
and U2690 (N_2690,N_1914,N_1891);
or U2691 (N_2691,N_1808,N_1452);
and U2692 (N_2692,N_1415,N_1761);
and U2693 (N_2693,N_1479,N_1036);
nand U2694 (N_2694,N_1303,N_1587);
nand U2695 (N_2695,N_1815,N_1206);
and U2696 (N_2696,N_1414,N_1734);
or U2697 (N_2697,N_1576,N_1741);
nor U2698 (N_2698,N_1500,N_1262);
nand U2699 (N_2699,N_1252,N_1346);
and U2700 (N_2700,N_1840,N_1967);
and U2701 (N_2701,N_1887,N_1006);
nor U2702 (N_2702,N_1835,N_1880);
and U2703 (N_2703,N_1584,N_1685);
and U2704 (N_2704,N_1836,N_1076);
nand U2705 (N_2705,N_1234,N_1991);
nor U2706 (N_2706,N_1276,N_1921);
nand U2707 (N_2707,N_1170,N_1241);
or U2708 (N_2708,N_1077,N_1726);
or U2709 (N_2709,N_1023,N_1674);
nand U2710 (N_2710,N_1799,N_1694);
and U2711 (N_2711,N_1486,N_1947);
or U2712 (N_2712,N_1553,N_1721);
nor U2713 (N_2713,N_1520,N_1108);
nor U2714 (N_2714,N_1118,N_1431);
or U2715 (N_2715,N_1650,N_1255);
nor U2716 (N_2716,N_1426,N_1710);
or U2717 (N_2717,N_1240,N_1792);
nand U2718 (N_2718,N_1528,N_1025);
and U2719 (N_2719,N_1661,N_1893);
or U2720 (N_2720,N_1292,N_1384);
and U2721 (N_2721,N_1972,N_1732);
nor U2722 (N_2722,N_1731,N_1824);
nor U2723 (N_2723,N_1469,N_1969);
or U2724 (N_2724,N_1813,N_1620);
nor U2725 (N_2725,N_1322,N_1902);
and U2726 (N_2726,N_1830,N_1966);
nand U2727 (N_2727,N_1762,N_1043);
nor U2728 (N_2728,N_1745,N_1894);
nor U2729 (N_2729,N_1256,N_1227);
nand U2730 (N_2730,N_1818,N_1283);
or U2731 (N_2731,N_1878,N_1479);
and U2732 (N_2732,N_1757,N_1347);
and U2733 (N_2733,N_1105,N_1697);
or U2734 (N_2734,N_1671,N_1566);
nand U2735 (N_2735,N_1669,N_1769);
or U2736 (N_2736,N_1391,N_1971);
or U2737 (N_2737,N_1854,N_1120);
or U2738 (N_2738,N_1713,N_1179);
and U2739 (N_2739,N_1702,N_1462);
nand U2740 (N_2740,N_1204,N_1670);
or U2741 (N_2741,N_1461,N_1849);
nor U2742 (N_2742,N_1227,N_1948);
and U2743 (N_2743,N_1326,N_1240);
nand U2744 (N_2744,N_1290,N_1915);
and U2745 (N_2745,N_1691,N_1102);
and U2746 (N_2746,N_1364,N_1831);
or U2747 (N_2747,N_1176,N_1081);
nor U2748 (N_2748,N_1050,N_1933);
and U2749 (N_2749,N_1911,N_1839);
or U2750 (N_2750,N_1844,N_1275);
nand U2751 (N_2751,N_1477,N_1229);
nor U2752 (N_2752,N_1557,N_1582);
nor U2753 (N_2753,N_1072,N_1216);
nand U2754 (N_2754,N_1039,N_1364);
or U2755 (N_2755,N_1801,N_1450);
and U2756 (N_2756,N_1851,N_1823);
nand U2757 (N_2757,N_1201,N_1966);
nor U2758 (N_2758,N_1559,N_1074);
or U2759 (N_2759,N_1141,N_1893);
nor U2760 (N_2760,N_1015,N_1123);
nor U2761 (N_2761,N_1012,N_1618);
and U2762 (N_2762,N_1416,N_1008);
nand U2763 (N_2763,N_1211,N_1374);
and U2764 (N_2764,N_1810,N_1314);
nand U2765 (N_2765,N_1494,N_1383);
nand U2766 (N_2766,N_1121,N_1024);
nor U2767 (N_2767,N_1539,N_1564);
nor U2768 (N_2768,N_1263,N_1637);
or U2769 (N_2769,N_1408,N_1065);
or U2770 (N_2770,N_1715,N_1834);
and U2771 (N_2771,N_1676,N_1417);
and U2772 (N_2772,N_1147,N_1612);
nand U2773 (N_2773,N_1185,N_1044);
and U2774 (N_2774,N_1379,N_1292);
or U2775 (N_2775,N_1424,N_1357);
nand U2776 (N_2776,N_1480,N_1821);
or U2777 (N_2777,N_1979,N_1233);
nand U2778 (N_2778,N_1922,N_1686);
and U2779 (N_2779,N_1421,N_1004);
or U2780 (N_2780,N_1595,N_1336);
nor U2781 (N_2781,N_1302,N_1123);
nand U2782 (N_2782,N_1652,N_1217);
and U2783 (N_2783,N_1399,N_1494);
or U2784 (N_2784,N_1117,N_1872);
and U2785 (N_2785,N_1230,N_1778);
and U2786 (N_2786,N_1387,N_1567);
nor U2787 (N_2787,N_1679,N_1295);
and U2788 (N_2788,N_1537,N_1936);
nand U2789 (N_2789,N_1912,N_1565);
nor U2790 (N_2790,N_1492,N_1898);
nand U2791 (N_2791,N_1671,N_1490);
and U2792 (N_2792,N_1893,N_1679);
nor U2793 (N_2793,N_1220,N_1974);
or U2794 (N_2794,N_1011,N_1015);
nor U2795 (N_2795,N_1752,N_1673);
or U2796 (N_2796,N_1213,N_1766);
nor U2797 (N_2797,N_1111,N_1594);
nor U2798 (N_2798,N_1768,N_1190);
nand U2799 (N_2799,N_1754,N_1130);
or U2800 (N_2800,N_1510,N_1748);
nand U2801 (N_2801,N_1686,N_1875);
nand U2802 (N_2802,N_1016,N_1084);
nor U2803 (N_2803,N_1402,N_1214);
and U2804 (N_2804,N_1232,N_1439);
or U2805 (N_2805,N_1518,N_1163);
and U2806 (N_2806,N_1040,N_1954);
nand U2807 (N_2807,N_1030,N_1407);
and U2808 (N_2808,N_1499,N_1382);
nor U2809 (N_2809,N_1085,N_1504);
nor U2810 (N_2810,N_1240,N_1356);
nand U2811 (N_2811,N_1605,N_1884);
or U2812 (N_2812,N_1216,N_1190);
and U2813 (N_2813,N_1641,N_1076);
and U2814 (N_2814,N_1496,N_1065);
and U2815 (N_2815,N_1106,N_1132);
or U2816 (N_2816,N_1148,N_1875);
and U2817 (N_2817,N_1752,N_1981);
nand U2818 (N_2818,N_1359,N_1188);
and U2819 (N_2819,N_1295,N_1550);
or U2820 (N_2820,N_1108,N_1667);
and U2821 (N_2821,N_1017,N_1297);
nand U2822 (N_2822,N_1051,N_1782);
or U2823 (N_2823,N_1374,N_1884);
nand U2824 (N_2824,N_1385,N_1725);
nand U2825 (N_2825,N_1912,N_1938);
or U2826 (N_2826,N_1675,N_1057);
nand U2827 (N_2827,N_1925,N_1823);
or U2828 (N_2828,N_1301,N_1615);
or U2829 (N_2829,N_1888,N_1017);
nand U2830 (N_2830,N_1700,N_1433);
nand U2831 (N_2831,N_1356,N_1514);
or U2832 (N_2832,N_1062,N_1242);
and U2833 (N_2833,N_1144,N_1718);
or U2834 (N_2834,N_1468,N_1833);
and U2835 (N_2835,N_1627,N_1730);
nand U2836 (N_2836,N_1098,N_1863);
nor U2837 (N_2837,N_1617,N_1995);
nand U2838 (N_2838,N_1864,N_1431);
nand U2839 (N_2839,N_1141,N_1979);
and U2840 (N_2840,N_1215,N_1411);
and U2841 (N_2841,N_1378,N_1483);
nand U2842 (N_2842,N_1067,N_1775);
and U2843 (N_2843,N_1863,N_1168);
nor U2844 (N_2844,N_1723,N_1757);
nand U2845 (N_2845,N_1692,N_1746);
and U2846 (N_2846,N_1737,N_1045);
and U2847 (N_2847,N_1171,N_1057);
and U2848 (N_2848,N_1213,N_1969);
nand U2849 (N_2849,N_1300,N_1241);
and U2850 (N_2850,N_1185,N_1506);
or U2851 (N_2851,N_1037,N_1931);
nand U2852 (N_2852,N_1941,N_1359);
and U2853 (N_2853,N_1830,N_1100);
nor U2854 (N_2854,N_1426,N_1502);
or U2855 (N_2855,N_1923,N_1724);
or U2856 (N_2856,N_1850,N_1984);
nor U2857 (N_2857,N_1141,N_1600);
or U2858 (N_2858,N_1683,N_1027);
nand U2859 (N_2859,N_1202,N_1689);
nand U2860 (N_2860,N_1825,N_1992);
or U2861 (N_2861,N_1730,N_1855);
nand U2862 (N_2862,N_1565,N_1511);
nand U2863 (N_2863,N_1954,N_1302);
xor U2864 (N_2864,N_1048,N_1155);
nor U2865 (N_2865,N_1428,N_1275);
nand U2866 (N_2866,N_1316,N_1362);
nor U2867 (N_2867,N_1553,N_1056);
or U2868 (N_2868,N_1018,N_1224);
and U2869 (N_2869,N_1676,N_1672);
nand U2870 (N_2870,N_1637,N_1319);
nand U2871 (N_2871,N_1493,N_1918);
nand U2872 (N_2872,N_1863,N_1917);
or U2873 (N_2873,N_1995,N_1877);
nand U2874 (N_2874,N_1625,N_1867);
or U2875 (N_2875,N_1942,N_1624);
nand U2876 (N_2876,N_1637,N_1908);
nand U2877 (N_2877,N_1125,N_1508);
nand U2878 (N_2878,N_1149,N_1344);
and U2879 (N_2879,N_1508,N_1205);
and U2880 (N_2880,N_1912,N_1028);
nand U2881 (N_2881,N_1853,N_1656);
nor U2882 (N_2882,N_1159,N_1240);
nor U2883 (N_2883,N_1338,N_1555);
nand U2884 (N_2884,N_1364,N_1705);
nand U2885 (N_2885,N_1303,N_1680);
or U2886 (N_2886,N_1608,N_1256);
nor U2887 (N_2887,N_1050,N_1473);
and U2888 (N_2888,N_1463,N_1502);
or U2889 (N_2889,N_1131,N_1969);
or U2890 (N_2890,N_1412,N_1651);
and U2891 (N_2891,N_1080,N_1515);
or U2892 (N_2892,N_1312,N_1540);
nand U2893 (N_2893,N_1717,N_1056);
nor U2894 (N_2894,N_1617,N_1726);
and U2895 (N_2895,N_1736,N_1949);
or U2896 (N_2896,N_1221,N_1775);
nor U2897 (N_2897,N_1493,N_1728);
or U2898 (N_2898,N_1163,N_1274);
nand U2899 (N_2899,N_1596,N_1954);
and U2900 (N_2900,N_1249,N_1562);
nor U2901 (N_2901,N_1659,N_1592);
nand U2902 (N_2902,N_1778,N_1409);
nor U2903 (N_2903,N_1088,N_1981);
nor U2904 (N_2904,N_1203,N_1513);
and U2905 (N_2905,N_1874,N_1777);
and U2906 (N_2906,N_1214,N_1312);
nand U2907 (N_2907,N_1414,N_1586);
and U2908 (N_2908,N_1856,N_1966);
and U2909 (N_2909,N_1620,N_1952);
nor U2910 (N_2910,N_1824,N_1496);
nand U2911 (N_2911,N_1186,N_1600);
or U2912 (N_2912,N_1665,N_1223);
or U2913 (N_2913,N_1639,N_1233);
or U2914 (N_2914,N_1544,N_1871);
nor U2915 (N_2915,N_1291,N_1364);
and U2916 (N_2916,N_1986,N_1121);
nand U2917 (N_2917,N_1643,N_1934);
and U2918 (N_2918,N_1175,N_1089);
and U2919 (N_2919,N_1177,N_1798);
or U2920 (N_2920,N_1305,N_1368);
nor U2921 (N_2921,N_1526,N_1159);
and U2922 (N_2922,N_1385,N_1522);
nand U2923 (N_2923,N_1526,N_1042);
and U2924 (N_2924,N_1524,N_1040);
nor U2925 (N_2925,N_1261,N_1466);
nand U2926 (N_2926,N_1392,N_1532);
and U2927 (N_2927,N_1849,N_1498);
nor U2928 (N_2928,N_1007,N_1793);
and U2929 (N_2929,N_1127,N_1750);
or U2930 (N_2930,N_1726,N_1387);
and U2931 (N_2931,N_1999,N_1422);
or U2932 (N_2932,N_1327,N_1713);
or U2933 (N_2933,N_1757,N_1776);
or U2934 (N_2934,N_1046,N_1929);
and U2935 (N_2935,N_1718,N_1545);
nor U2936 (N_2936,N_1524,N_1039);
or U2937 (N_2937,N_1941,N_1493);
and U2938 (N_2938,N_1455,N_1246);
nand U2939 (N_2939,N_1738,N_1079);
or U2940 (N_2940,N_1122,N_1444);
nor U2941 (N_2941,N_1044,N_1702);
or U2942 (N_2942,N_1659,N_1624);
or U2943 (N_2943,N_1970,N_1064);
or U2944 (N_2944,N_1453,N_1233);
nand U2945 (N_2945,N_1772,N_1585);
nand U2946 (N_2946,N_1215,N_1603);
or U2947 (N_2947,N_1940,N_1391);
or U2948 (N_2948,N_1817,N_1850);
nand U2949 (N_2949,N_1930,N_1657);
nand U2950 (N_2950,N_1143,N_1189);
nor U2951 (N_2951,N_1505,N_1588);
nand U2952 (N_2952,N_1612,N_1746);
and U2953 (N_2953,N_1231,N_1642);
and U2954 (N_2954,N_1930,N_1914);
nor U2955 (N_2955,N_1762,N_1661);
nand U2956 (N_2956,N_1744,N_1694);
nor U2957 (N_2957,N_1921,N_1948);
nand U2958 (N_2958,N_1136,N_1774);
nand U2959 (N_2959,N_1707,N_1813);
nand U2960 (N_2960,N_1466,N_1819);
or U2961 (N_2961,N_1973,N_1454);
or U2962 (N_2962,N_1044,N_1970);
nor U2963 (N_2963,N_1987,N_1252);
nand U2964 (N_2964,N_1989,N_1870);
or U2965 (N_2965,N_1791,N_1754);
and U2966 (N_2966,N_1685,N_1025);
nor U2967 (N_2967,N_1664,N_1246);
nor U2968 (N_2968,N_1203,N_1854);
and U2969 (N_2969,N_1187,N_1826);
nor U2970 (N_2970,N_1530,N_1510);
or U2971 (N_2971,N_1814,N_1598);
xnor U2972 (N_2972,N_1641,N_1942);
or U2973 (N_2973,N_1195,N_1304);
nor U2974 (N_2974,N_1716,N_1794);
or U2975 (N_2975,N_1225,N_1703);
nand U2976 (N_2976,N_1981,N_1886);
nand U2977 (N_2977,N_1186,N_1322);
nand U2978 (N_2978,N_1519,N_1496);
nor U2979 (N_2979,N_1953,N_1922);
nand U2980 (N_2980,N_1942,N_1372);
nor U2981 (N_2981,N_1097,N_1165);
nand U2982 (N_2982,N_1735,N_1448);
nand U2983 (N_2983,N_1537,N_1257);
nor U2984 (N_2984,N_1018,N_1299);
and U2985 (N_2985,N_1541,N_1746);
or U2986 (N_2986,N_1834,N_1618);
nor U2987 (N_2987,N_1179,N_1925);
nor U2988 (N_2988,N_1683,N_1510);
or U2989 (N_2989,N_1694,N_1042);
and U2990 (N_2990,N_1590,N_1472);
and U2991 (N_2991,N_1163,N_1990);
and U2992 (N_2992,N_1176,N_1048);
nor U2993 (N_2993,N_1801,N_1759);
or U2994 (N_2994,N_1723,N_1413);
nand U2995 (N_2995,N_1206,N_1322);
nand U2996 (N_2996,N_1899,N_1134);
or U2997 (N_2997,N_1793,N_1242);
nand U2998 (N_2998,N_1028,N_1114);
and U2999 (N_2999,N_1874,N_1639);
and UO_0 (O_0,N_2974,N_2506);
nor UO_1 (O_1,N_2234,N_2730);
or UO_2 (O_2,N_2806,N_2290);
nand UO_3 (O_3,N_2799,N_2649);
or UO_4 (O_4,N_2503,N_2460);
or UO_5 (O_5,N_2155,N_2393);
or UO_6 (O_6,N_2338,N_2851);
and UO_7 (O_7,N_2388,N_2544);
xnor UO_8 (O_8,N_2145,N_2299);
or UO_9 (O_9,N_2079,N_2275);
nand UO_10 (O_10,N_2431,N_2432);
nor UO_11 (O_11,N_2477,N_2747);
nor UO_12 (O_12,N_2762,N_2075);
nor UO_13 (O_13,N_2695,N_2436);
or UO_14 (O_14,N_2047,N_2426);
nand UO_15 (O_15,N_2434,N_2898);
nor UO_16 (O_16,N_2239,N_2727);
nand UO_17 (O_17,N_2895,N_2919);
nand UO_18 (O_18,N_2912,N_2813);
and UO_19 (O_19,N_2971,N_2441);
or UO_20 (O_20,N_2630,N_2067);
or UO_21 (O_21,N_2039,N_2716);
and UO_22 (O_22,N_2051,N_2328);
nor UO_23 (O_23,N_2597,N_2473);
nor UO_24 (O_24,N_2211,N_2420);
or UO_25 (O_25,N_2012,N_2086);
and UO_26 (O_26,N_2031,N_2395);
nand UO_27 (O_27,N_2190,N_2707);
nand UO_28 (O_28,N_2790,N_2748);
xnor UO_29 (O_29,N_2640,N_2585);
nand UO_30 (O_30,N_2939,N_2807);
or UO_31 (O_31,N_2524,N_2653);
and UO_32 (O_32,N_2107,N_2778);
nand UO_33 (O_33,N_2463,N_2046);
and UO_34 (O_34,N_2988,N_2365);
or UO_35 (O_35,N_2108,N_2595);
or UO_36 (O_36,N_2302,N_2602);
nand UO_37 (O_37,N_2651,N_2036);
or UO_38 (O_38,N_2952,N_2594);
and UO_39 (O_39,N_2427,N_2509);
nand UO_40 (O_40,N_2989,N_2829);
nor UO_41 (O_41,N_2025,N_2271);
and UO_42 (O_42,N_2871,N_2449);
and UO_43 (O_43,N_2179,N_2562);
and UO_44 (O_44,N_2852,N_2663);
nor UO_45 (O_45,N_2318,N_2744);
and UO_46 (O_46,N_2982,N_2618);
nand UO_47 (O_47,N_2557,N_2474);
nand UO_48 (O_48,N_2687,N_2932);
and UO_49 (O_49,N_2337,N_2158);
or UO_50 (O_50,N_2745,N_2720);
nand UO_51 (O_51,N_2887,N_2454);
nor UO_52 (O_52,N_2209,N_2811);
nand UO_53 (O_53,N_2896,N_2264);
and UO_54 (O_54,N_2515,N_2058);
nand UO_55 (O_55,N_2263,N_2537);
and UO_56 (O_56,N_2410,N_2044);
nor UO_57 (O_57,N_2733,N_2404);
or UO_58 (O_58,N_2776,N_2621);
nor UO_59 (O_59,N_2081,N_2493);
and UO_60 (O_60,N_2013,N_2225);
nand UO_61 (O_61,N_2043,N_2052);
nor UO_62 (O_62,N_2160,N_2576);
nor UO_63 (O_63,N_2294,N_2478);
nor UO_64 (O_64,N_2428,N_2001);
and UO_65 (O_65,N_2091,N_2827);
nand UO_66 (O_66,N_2169,N_2669);
or UO_67 (O_67,N_2507,N_2451);
or UO_68 (O_68,N_2379,N_2831);
or UO_69 (O_69,N_2459,N_2076);
nand UO_70 (O_70,N_2635,N_2125);
xor UO_71 (O_71,N_2516,N_2606);
or UO_72 (O_72,N_2942,N_2134);
nor UO_73 (O_73,N_2010,N_2953);
nand UO_74 (O_74,N_2380,N_2631);
nand UO_75 (O_75,N_2022,N_2986);
nand UO_76 (O_76,N_2425,N_2297);
or UO_77 (O_77,N_2386,N_2961);
nor UO_78 (O_78,N_2858,N_2998);
nor UO_79 (O_79,N_2705,N_2962);
and UO_80 (O_80,N_2166,N_2784);
nor UO_81 (O_81,N_2083,N_2540);
nand UO_82 (O_82,N_2118,N_2462);
and UO_83 (O_83,N_2583,N_2842);
nand UO_84 (O_84,N_2711,N_2140);
nand UO_85 (O_85,N_2609,N_2676);
or UO_86 (O_86,N_2893,N_2909);
and UO_87 (O_87,N_2770,N_2287);
or UO_88 (O_88,N_2468,N_2527);
or UO_89 (O_89,N_2743,N_2068);
nand UO_90 (O_90,N_2840,N_2274);
nand UO_91 (O_91,N_2485,N_2498);
or UO_92 (O_92,N_2200,N_2066);
nand UO_93 (O_93,N_2242,N_2384);
or UO_94 (O_94,N_2916,N_2149);
or UO_95 (O_95,N_2202,N_2715);
nand UO_96 (O_96,N_2526,N_2220);
nand UO_97 (O_97,N_2161,N_2728);
nor UO_98 (O_98,N_2453,N_2366);
or UO_99 (O_99,N_2890,N_2773);
nor UO_100 (O_100,N_2575,N_2628);
nand UO_101 (O_101,N_2456,N_2946);
and UO_102 (O_102,N_2276,N_2320);
nor UO_103 (O_103,N_2593,N_2972);
nand UO_104 (O_104,N_2882,N_2607);
or UO_105 (O_105,N_2963,N_2838);
nand UO_106 (O_106,N_2139,N_2258);
nor UO_107 (O_107,N_2689,N_2523);
xor UO_108 (O_108,N_2205,N_2159);
or UO_109 (O_109,N_2543,N_2339);
nor UO_110 (O_110,N_2448,N_2063);
or UO_111 (O_111,N_2880,N_2127);
or UO_112 (O_112,N_2027,N_2777);
nand UO_113 (O_113,N_2935,N_2009);
nor UO_114 (O_114,N_2930,N_2400);
and UO_115 (O_115,N_2056,N_2789);
nand UO_116 (O_116,N_2482,N_2574);
and UO_117 (O_117,N_2554,N_2119);
nor UO_118 (O_118,N_2708,N_2615);
or UO_119 (O_119,N_2530,N_2344);
or UO_120 (O_120,N_2977,N_2286);
nand UO_121 (O_121,N_2390,N_2280);
nor UO_122 (O_122,N_2800,N_2496);
nor UO_123 (O_123,N_2331,N_2250);
nand UO_124 (O_124,N_2182,N_2317);
or UO_125 (O_125,N_2661,N_2196);
nand UO_126 (O_126,N_2221,N_2110);
or UO_127 (O_127,N_2148,N_2112);
or UO_128 (O_128,N_2268,N_2579);
nand UO_129 (O_129,N_2472,N_2283);
nand UO_130 (O_130,N_2633,N_2752);
and UO_131 (O_131,N_2826,N_2756);
nand UO_132 (O_132,N_2521,N_2084);
nor UO_133 (O_133,N_2569,N_2124);
or UO_134 (O_134,N_2985,N_2105);
or UO_135 (O_135,N_2552,N_2195);
and UO_136 (O_136,N_2188,N_2539);
and UO_137 (O_137,N_2230,N_2017);
nor UO_138 (O_138,N_2656,N_2396);
nor UO_139 (O_139,N_2915,N_2954);
nand UO_140 (O_140,N_2817,N_2967);
and UO_141 (O_141,N_2500,N_2865);
and UO_142 (O_142,N_2003,N_2367);
and UO_143 (O_143,N_2435,N_2879);
and UO_144 (O_144,N_2550,N_2751);
or UO_145 (O_145,N_2361,N_2005);
and UO_146 (O_146,N_2674,N_2305);
nand UO_147 (O_147,N_2090,N_2513);
nand UO_148 (O_148,N_2164,N_2528);
nor UO_149 (O_149,N_2210,N_2995);
and UO_150 (O_150,N_2815,N_2313);
nor UO_151 (O_151,N_2658,N_2465);
and UO_152 (O_152,N_2872,N_2251);
and UO_153 (O_153,N_2444,N_2973);
nand UO_154 (O_154,N_2673,N_2901);
nor UO_155 (O_155,N_2095,N_2144);
or UO_156 (O_156,N_2399,N_2582);
or UO_157 (O_157,N_2937,N_2335);
or UO_158 (O_158,N_2345,N_2285);
or UO_159 (O_159,N_2497,N_2259);
nand UO_160 (O_160,N_2578,N_2522);
or UO_161 (O_161,N_2694,N_2494);
nand UO_162 (O_162,N_2011,N_2990);
and UO_163 (O_163,N_2545,N_2510);
or UO_164 (O_164,N_2358,N_2089);
and UO_165 (O_165,N_2682,N_2355);
and UO_166 (O_166,N_2308,N_2270);
or UO_167 (O_167,N_2941,N_2007);
nand UO_168 (O_168,N_2150,N_2353);
and UO_169 (O_169,N_2729,N_2814);
or UO_170 (O_170,N_2619,N_2841);
nor UO_171 (O_171,N_2376,N_2466);
or UO_172 (O_172,N_2731,N_2311);
or UO_173 (O_173,N_2843,N_2760);
and UO_174 (O_174,N_2306,N_2996);
nand UO_175 (O_175,N_2207,N_2677);
and UO_176 (O_176,N_2429,N_2710);
and UO_177 (O_177,N_2212,N_2678);
nor UO_178 (O_178,N_2352,N_2855);
nor UO_179 (O_179,N_2443,N_2152);
xor UO_180 (O_180,N_2596,N_2129);
nand UO_181 (O_181,N_2903,N_2757);
nor UO_182 (O_182,N_2934,N_2173);
or UO_183 (O_183,N_2162,N_2062);
nor UO_184 (O_184,N_2816,N_2269);
and UO_185 (O_185,N_2723,N_2726);
nor UO_186 (O_186,N_2120,N_2914);
nor UO_187 (O_187,N_2787,N_2892);
nand UO_188 (O_188,N_2214,N_2732);
or UO_189 (O_189,N_2644,N_2216);
or UO_190 (O_190,N_2796,N_2991);
and UO_191 (O_191,N_2020,N_2721);
nand UO_192 (O_192,N_2310,N_2712);
and UO_193 (O_193,N_2588,N_2284);
and UO_194 (O_194,N_2246,N_2714);
and UO_195 (O_195,N_2533,N_2944);
and UO_196 (O_196,N_2368,N_2016);
nand UO_197 (O_197,N_2303,N_2006);
and UO_198 (O_198,N_2755,N_2378);
nand UO_199 (O_199,N_2146,N_2080);
nand UO_200 (O_200,N_2072,N_2559);
and UO_201 (O_201,N_2795,N_2201);
nand UO_202 (O_202,N_2746,N_2725);
nor UO_203 (O_203,N_2761,N_2312);
or UO_204 (O_204,N_2680,N_2244);
and UO_205 (O_205,N_2542,N_2249);
nor UO_206 (O_206,N_2889,N_2958);
nand UO_207 (O_207,N_2048,N_2315);
nand UO_208 (O_208,N_2719,N_2423);
and UO_209 (O_209,N_2856,N_2359);
nor UO_210 (O_210,N_2419,N_2900);
nor UO_211 (O_211,N_2102,N_2165);
nand UO_212 (O_212,N_2739,N_2325);
and UO_213 (O_213,N_2861,N_2348);
and UO_214 (O_214,N_2867,N_2573);
and UO_215 (O_215,N_2098,N_2548);
and UO_216 (O_216,N_2405,N_2577);
nor UO_217 (O_217,N_2830,N_2183);
nand UO_218 (O_218,N_2553,N_2925);
and UO_219 (O_219,N_2490,N_2185);
nor UO_220 (O_220,N_2223,N_2877);
nor UO_221 (O_221,N_2863,N_2862);
and UO_222 (O_222,N_2955,N_2021);
or UO_223 (O_223,N_2910,N_2070);
and UO_224 (O_224,N_2458,N_2605);
nand UO_225 (O_225,N_2372,N_2032);
or UO_226 (O_226,N_2825,N_2130);
and UO_227 (O_227,N_2696,N_2277);
xor UO_228 (O_228,N_2520,N_2316);
nand UO_229 (O_229,N_2979,N_2194);
and UO_230 (O_230,N_2237,N_2413);
and UO_231 (O_231,N_2018,N_2753);
or UO_232 (O_232,N_2881,N_2002);
and UO_233 (O_233,N_2133,N_2298);
nor UO_234 (O_234,N_2422,N_2564);
and UO_235 (O_235,N_2671,N_2096);
or UO_236 (O_236,N_2004,N_2610);
nand UO_237 (O_237,N_2945,N_2397);
nand UO_238 (O_238,N_2163,N_2546);
nand UO_239 (O_239,N_2951,N_2672);
nand UO_240 (O_240,N_2301,N_2272);
nand UO_241 (O_241,N_2612,N_2532);
nor UO_242 (O_242,N_2929,N_2650);
and UO_243 (O_243,N_2099,N_2992);
nand UO_244 (O_244,N_2447,N_2904);
nor UO_245 (O_245,N_2467,N_2071);
nor UO_246 (O_246,N_2486,N_2864);
nor UO_247 (O_247,N_2906,N_2767);
or UO_248 (O_248,N_2886,N_2464);
nand UO_249 (O_249,N_2033,N_2783);
nand UO_250 (O_250,N_2768,N_2387);
or UO_251 (O_251,N_2804,N_2101);
and UO_252 (O_252,N_2781,N_2818);
nand UO_253 (O_253,N_2053,N_2803);
nand UO_254 (O_254,N_2808,N_2924);
or UO_255 (O_255,N_2421,N_2505);
or UO_256 (O_256,N_2853,N_2983);
and UO_257 (O_257,N_2383,N_2394);
or UO_258 (O_258,N_2774,N_2600);
nand UO_259 (O_259,N_2717,N_2476);
xor UO_260 (O_260,N_2495,N_2218);
or UO_261 (O_261,N_2117,N_2788);
nor UO_262 (O_262,N_2764,N_2975);
nand UO_263 (O_263,N_2997,N_2627);
and UO_264 (O_264,N_2055,N_2547);
and UO_265 (O_265,N_2085,N_2424);
nand UO_266 (O_266,N_2260,N_2920);
nor UO_267 (O_267,N_2178,N_2667);
or UO_268 (O_268,N_2180,N_2970);
nand UO_269 (O_269,N_2531,N_2391);
nand UO_270 (O_270,N_2833,N_2785);
and UO_271 (O_271,N_2568,N_2138);
nand UO_272 (O_272,N_2824,N_2686);
nand UO_273 (O_273,N_2965,N_2571);
or UO_274 (O_274,N_2253,N_2181);
or UO_275 (O_275,N_2135,N_2632);
or UO_276 (O_276,N_2878,N_2758);
or UO_277 (O_277,N_2293,N_2342);
nand UO_278 (O_278,N_2324,N_2199);
nand UO_279 (O_279,N_2374,N_2488);
nand UO_280 (O_280,N_2088,N_2481);
nor UO_281 (O_281,N_2549,N_2222);
or UO_282 (O_282,N_2791,N_2598);
and UO_283 (O_283,N_2812,N_2567);
nor UO_284 (O_284,N_2128,N_2587);
or UO_285 (O_285,N_2793,N_2534);
nor UO_286 (O_286,N_2452,N_2917);
or UO_287 (O_287,N_2837,N_2362);
nor UO_288 (O_288,N_2620,N_2614);
nand UO_289 (O_289,N_2763,N_2489);
nor UO_290 (O_290,N_2364,N_2082);
nand UO_291 (O_291,N_2077,N_2151);
nor UO_292 (O_292,N_2398,N_2450);
nor UO_293 (O_293,N_2646,N_2336);
nand UO_294 (O_294,N_2798,N_2535);
nand UO_295 (O_295,N_2832,N_2078);
or UO_296 (O_296,N_2279,N_2295);
nand UO_297 (O_297,N_2501,N_2153);
or UO_298 (O_298,N_2257,N_2690);
nor UO_299 (O_299,N_2839,N_2873);
nand UO_300 (O_300,N_2235,N_2045);
or UO_301 (O_301,N_2252,N_2330);
xnor UO_302 (O_302,N_2233,N_2377);
nand UO_303 (O_303,N_2304,N_2154);
nand UO_304 (O_304,N_2821,N_2885);
nor UO_305 (O_305,N_2603,N_2634);
and UO_306 (O_306,N_2688,N_2704);
and UO_307 (O_307,N_2766,N_2643);
nand UO_308 (O_308,N_2718,N_2581);
nor UO_309 (O_309,N_2802,N_2147);
nor UO_310 (O_310,N_2625,N_2430);
nand UO_311 (O_311,N_2191,N_2232);
or UO_312 (O_312,N_2541,N_2215);
or UO_313 (O_313,N_2623,N_2943);
nand UO_314 (O_314,N_2073,N_2256);
nand UO_315 (O_315,N_2104,N_2978);
or UO_316 (O_316,N_2291,N_2442);
and UO_317 (O_317,N_2357,N_2255);
nor UO_318 (O_318,N_2964,N_2484);
or UO_319 (O_319,N_2029,N_2103);
nand UO_320 (O_320,N_2340,N_2849);
nand UO_321 (O_321,N_2641,N_2229);
and UO_322 (O_322,N_2599,N_2470);
nand UO_323 (O_323,N_2122,N_2197);
or UO_324 (O_324,N_2994,N_2115);
nand UO_325 (O_325,N_2884,N_2775);
nand UO_326 (O_326,N_2735,N_2563);
or UO_327 (O_327,N_2848,N_2517);
nor UO_328 (O_328,N_2681,N_2868);
or UO_329 (O_329,N_2349,N_2565);
nand UO_330 (O_330,N_2536,N_2469);
and UO_331 (O_331,N_2859,N_2412);
xor UO_332 (O_332,N_2437,N_2957);
and UO_333 (O_333,N_2471,N_2350);
and UO_334 (O_334,N_2844,N_2969);
or UO_335 (O_335,N_2499,N_2809);
nor UO_336 (O_336,N_2854,N_2660);
or UO_337 (O_337,N_2480,N_2491);
nor UO_338 (O_338,N_2457,N_2401);
nor UO_339 (O_339,N_2409,N_2874);
and UO_340 (O_340,N_2243,N_2870);
nor UO_341 (O_341,N_2529,N_2888);
nand UO_342 (O_342,N_2823,N_2240);
or UO_343 (O_343,N_2512,N_2699);
nor UO_344 (O_344,N_2204,N_2341);
xor UO_345 (O_345,N_2759,N_2332);
nor UO_346 (O_346,N_2654,N_2950);
and UO_347 (O_347,N_2700,N_2741);
or UO_348 (O_348,N_2203,N_2172);
or UO_349 (O_349,N_2319,N_2736);
and UO_350 (O_350,N_2902,N_2966);
and UO_351 (O_351,N_2665,N_2248);
and UO_352 (O_352,N_2281,N_2604);
nor UO_353 (O_353,N_2267,N_2231);
or UO_354 (O_354,N_2956,N_2558);
nor UO_355 (O_355,N_2282,N_2241);
nor UO_356 (O_356,N_2168,N_2692);
or UO_357 (O_357,N_2525,N_2691);
nor UO_358 (O_358,N_2749,N_2309);
or UO_359 (O_359,N_2407,N_2703);
nand UO_360 (O_360,N_2213,N_2750);
or UO_361 (O_361,N_2948,N_2189);
and UO_362 (O_362,N_2415,N_2987);
nor UO_363 (O_363,N_2706,N_2176);
nor UO_364 (O_364,N_2296,N_2406);
nor UO_365 (O_365,N_2087,N_2132);
nand UO_366 (O_366,N_2265,N_2392);
nor UO_367 (O_367,N_2363,N_2822);
nand UO_368 (O_368,N_2502,N_2114);
nor UO_369 (O_369,N_2936,N_2740);
nor UO_370 (O_370,N_2670,N_2907);
nor UO_371 (O_371,N_2679,N_2926);
nor UO_372 (O_372,N_2794,N_2224);
or UO_373 (O_373,N_2551,N_2927);
nor UO_374 (O_374,N_2652,N_2984);
nand UO_375 (O_375,N_2883,N_2570);
nand UO_376 (O_376,N_2175,N_2369);
nor UO_377 (O_377,N_2590,N_2245);
and UO_378 (O_378,N_2608,N_2187);
and UO_379 (O_379,N_2779,N_2061);
or UO_380 (O_380,N_2734,N_2034);
nand UO_381 (O_381,N_2835,N_2254);
nand UO_382 (O_382,N_2142,N_2624);
and UO_383 (O_383,N_2684,N_2111);
and UO_384 (O_384,N_2184,N_2845);
nand UO_385 (O_385,N_2639,N_2024);
nand UO_386 (O_386,N_2617,N_2097);
or UO_387 (O_387,N_2492,N_2373);
nand UO_388 (O_388,N_2206,N_2461);
and UO_389 (O_389,N_2918,N_2050);
or UO_390 (O_390,N_2015,N_2026);
nand UO_391 (O_391,N_2266,N_2846);
and UO_392 (O_392,N_2504,N_2642);
nor UO_393 (O_393,N_2136,N_2780);
and UO_394 (O_394,N_2908,N_2698);
xnor UO_395 (O_395,N_2030,N_2177);
xnor UO_396 (O_396,N_2288,N_2314);
nor UO_397 (O_397,N_2064,N_2586);
or UO_398 (O_398,N_2333,N_2069);
nor UO_399 (O_399,N_2629,N_2611);
nor UO_400 (O_400,N_2968,N_2402);
nor UO_401 (O_401,N_2226,N_2518);
nand UO_402 (O_402,N_2113,N_2300);
or UO_403 (O_403,N_2126,N_2100);
nor UO_404 (O_404,N_2273,N_2561);
or UO_405 (O_405,N_2008,N_2913);
nand UO_406 (O_406,N_2307,N_2592);
and UO_407 (O_407,N_2123,N_2322);
or UO_408 (O_408,N_2143,N_2439);
and UO_409 (O_409,N_2662,N_2121);
nand UO_410 (O_410,N_2408,N_2261);
and UO_411 (O_411,N_2765,N_2041);
nand UO_412 (O_412,N_2616,N_2038);
and UO_413 (O_413,N_2580,N_2771);
and UO_414 (O_414,N_2836,N_2891);
and UO_415 (O_415,N_2054,N_2820);
or UO_416 (O_416,N_2327,N_2131);
and UO_417 (O_417,N_2106,N_2360);
nor UO_418 (O_418,N_2869,N_2343);
nand UO_419 (O_419,N_2389,N_2475);
xor UO_420 (O_420,N_2555,N_2828);
and UO_421 (O_421,N_2354,N_2219);
and UO_422 (O_422,N_2647,N_2049);
or UO_423 (O_423,N_2797,N_2446);
and UO_424 (O_424,N_2713,N_2514);
nor UO_425 (O_425,N_2170,N_2921);
nor UO_426 (O_426,N_2356,N_2247);
nand UO_427 (O_427,N_2782,N_2709);
nor UO_428 (O_428,N_2414,N_2724);
and UO_429 (O_429,N_2174,N_2483);
xnor UO_430 (O_430,N_2940,N_2192);
and UO_431 (O_431,N_2262,N_2487);
or UO_432 (O_432,N_2810,N_2928);
xor UO_433 (O_433,N_2742,N_2860);
and UO_434 (O_434,N_2959,N_2657);
nand UO_435 (O_435,N_2792,N_2278);
nor UO_436 (O_436,N_2613,N_2701);
or UO_437 (O_437,N_2385,N_2445);
nor UO_438 (O_438,N_2508,N_2065);
or UO_439 (O_439,N_2938,N_2238);
or UO_440 (O_440,N_2208,N_2923);
and UO_441 (O_441,N_2217,N_2511);
and UO_442 (O_442,N_2805,N_2976);
nor UO_443 (O_443,N_2664,N_2866);
and UO_444 (O_444,N_2014,N_2722);
nor UO_445 (O_445,N_2897,N_2371);
nor UO_446 (O_446,N_2351,N_2850);
nand UO_447 (O_447,N_2093,N_2993);
or UO_448 (O_448,N_2922,N_2334);
or UO_449 (O_449,N_2433,N_2772);
nor UO_450 (O_450,N_2193,N_2638);
xor UO_451 (O_451,N_2227,N_2572);
or UO_452 (O_452,N_2947,N_2659);
nand UO_453 (O_453,N_2933,N_2167);
or UO_454 (O_454,N_2801,N_2042);
nand UO_455 (O_455,N_2754,N_2949);
nand UO_456 (O_456,N_2438,N_2589);
or UO_457 (O_457,N_2876,N_2057);
or UO_458 (O_458,N_2019,N_2347);
and UO_459 (O_459,N_2556,N_2074);
nand UO_460 (O_460,N_2847,N_2834);
or UO_461 (O_461,N_2591,N_2668);
nand UO_462 (O_462,N_2769,N_2157);
and UO_463 (O_463,N_2819,N_2675);
nor UO_464 (O_464,N_2685,N_2228);
nor UO_465 (O_465,N_2584,N_2479);
nand UO_466 (O_466,N_2236,N_2693);
and UO_467 (O_467,N_2648,N_2137);
nor UO_468 (O_468,N_2786,N_2417);
nor UO_469 (O_469,N_2738,N_2116);
nand UO_470 (O_470,N_2329,N_2346);
nor UO_471 (O_471,N_2186,N_2403);
and UO_472 (O_472,N_2289,N_2875);
nor UO_473 (O_473,N_2416,N_2381);
nor UO_474 (O_474,N_2092,N_2198);
and UO_475 (O_475,N_2999,N_2899);
and UO_476 (O_476,N_2737,N_2519);
nor UO_477 (O_477,N_2911,N_2037);
and UO_478 (O_478,N_2326,N_2059);
and UO_479 (O_479,N_2683,N_2382);
or UO_480 (O_480,N_2455,N_2601);
nor UO_481 (O_481,N_2109,N_2411);
or UO_482 (O_482,N_2697,N_2035);
nand UO_483 (O_483,N_2566,N_2370);
or UO_484 (O_484,N_2171,N_2626);
nor UO_485 (O_485,N_2857,N_2156);
and UO_486 (O_486,N_2560,N_2094);
and UO_487 (O_487,N_2375,N_2023);
nor UO_488 (O_488,N_2418,N_2141);
nand UO_489 (O_489,N_2981,N_2655);
or UO_490 (O_490,N_2645,N_2292);
nand UO_491 (O_491,N_2538,N_2666);
or UO_492 (O_492,N_2636,N_2702);
nor UO_493 (O_493,N_2931,N_2980);
nand UO_494 (O_494,N_2960,N_2894);
nor UO_495 (O_495,N_2028,N_2060);
nor UO_496 (O_496,N_2637,N_2321);
or UO_497 (O_497,N_2000,N_2905);
nor UO_498 (O_498,N_2323,N_2622);
nand UO_499 (O_499,N_2440,N_2040);
endmodule