module basic_750_5000_1000_5_levels_2xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
nand U0 (N_0,In_511,In_217);
nor U1 (N_1,In_359,In_299);
nand U2 (N_2,In_683,In_218);
nand U3 (N_3,In_732,In_45);
nand U4 (N_4,In_625,In_428);
nor U5 (N_5,In_80,In_110);
nand U6 (N_6,In_214,In_573);
and U7 (N_7,In_11,In_333);
and U8 (N_8,In_220,In_698);
and U9 (N_9,In_709,In_326);
and U10 (N_10,In_638,In_649);
and U11 (N_11,In_191,In_648);
and U12 (N_12,In_463,In_387);
nor U13 (N_13,In_609,In_472);
nand U14 (N_14,In_377,In_79);
or U15 (N_15,In_200,In_340);
or U16 (N_16,In_584,In_636);
xnor U17 (N_17,In_249,In_597);
nand U18 (N_18,In_221,In_321);
xor U19 (N_19,In_152,In_660);
nor U20 (N_20,In_572,In_681);
and U21 (N_21,In_645,In_341);
or U22 (N_22,In_216,In_144);
nor U23 (N_23,In_274,In_189);
nor U24 (N_24,In_722,In_205);
nand U25 (N_25,In_153,In_251);
or U26 (N_26,In_442,In_529);
and U27 (N_27,In_320,In_92);
nand U28 (N_28,In_501,In_151);
nor U29 (N_29,In_52,In_165);
or U30 (N_30,In_420,In_48);
and U31 (N_31,In_739,In_591);
nand U32 (N_32,In_139,In_713);
nand U33 (N_33,In_395,In_237);
xor U34 (N_34,In_432,In_56);
nor U35 (N_35,In_479,In_720);
and U36 (N_36,In_381,In_230);
nand U37 (N_37,In_581,In_540);
nor U38 (N_38,In_673,In_714);
nor U39 (N_39,In_170,In_691);
or U40 (N_40,In_425,In_325);
nor U41 (N_41,In_113,In_568);
nand U42 (N_42,In_87,In_258);
or U43 (N_43,In_36,In_305);
and U44 (N_44,In_104,In_279);
nand U45 (N_45,In_630,In_357);
nand U46 (N_46,In_702,In_328);
xnor U47 (N_47,In_562,In_613);
or U48 (N_48,In_440,In_746);
or U49 (N_49,In_231,In_475);
or U50 (N_50,In_277,In_361);
nand U51 (N_51,In_253,In_372);
nor U52 (N_52,In_601,In_287);
and U53 (N_53,In_672,In_273);
or U54 (N_54,In_460,In_286);
xor U55 (N_55,In_524,In_336);
and U56 (N_56,In_350,In_384);
nor U57 (N_57,In_106,In_242);
nand U58 (N_58,In_76,In_243);
nor U59 (N_59,In_201,In_160);
and U60 (N_60,In_177,In_111);
nand U61 (N_61,In_682,In_268);
or U62 (N_62,In_347,In_539);
and U63 (N_63,In_364,In_495);
nor U64 (N_64,In_745,In_675);
and U65 (N_65,In_257,In_136);
and U66 (N_66,In_285,In_639);
nand U67 (N_67,In_606,In_203);
or U68 (N_68,In_541,In_657);
xnor U69 (N_69,In_626,In_598);
nand U70 (N_70,In_504,In_448);
or U71 (N_71,In_716,In_518);
nor U72 (N_72,In_138,In_267);
nor U73 (N_73,In_602,In_119);
or U74 (N_74,In_181,In_509);
or U75 (N_75,In_667,In_179);
nor U76 (N_76,In_150,In_409);
nand U77 (N_77,In_434,In_93);
or U78 (N_78,In_63,In_489);
xor U79 (N_79,In_309,In_345);
nor U80 (N_80,In_31,In_441);
or U81 (N_81,In_33,In_430);
nand U82 (N_82,In_17,In_629);
and U83 (N_83,In_346,In_133);
and U84 (N_84,In_417,In_500);
nand U85 (N_85,In_163,In_487);
and U86 (N_86,In_85,In_567);
or U87 (N_87,In_70,In_47);
and U88 (N_88,In_224,In_553);
and U89 (N_89,In_634,In_383);
nor U90 (N_90,In_679,In_736);
or U91 (N_91,In_588,In_414);
or U92 (N_92,In_307,In_450);
and U93 (N_93,In_664,In_248);
or U94 (N_94,In_456,In_9);
nand U95 (N_95,In_207,In_611);
or U96 (N_96,In_316,In_422);
xnor U97 (N_97,In_140,In_402);
and U98 (N_98,In_586,In_161);
nand U99 (N_99,In_652,In_507);
and U100 (N_100,In_526,In_519);
or U101 (N_101,In_656,In_536);
and U102 (N_102,In_491,In_356);
and U103 (N_103,In_143,In_368);
or U104 (N_104,In_585,In_329);
and U105 (N_105,In_729,In_98);
nand U106 (N_106,In_223,In_449);
nand U107 (N_107,In_15,In_2);
and U108 (N_108,In_738,In_544);
nor U109 (N_109,In_109,In_546);
or U110 (N_110,In_471,In_418);
and U111 (N_111,In_74,In_294);
nand U112 (N_112,In_677,In_49);
nand U113 (N_113,In_718,In_470);
and U114 (N_114,In_332,In_137);
nor U115 (N_115,In_727,In_592);
and U116 (N_116,In_228,In_50);
nor U117 (N_117,In_412,In_476);
and U118 (N_118,In_619,In_5);
nand U119 (N_119,In_662,In_292);
nand U120 (N_120,In_311,In_742);
nor U121 (N_121,In_306,In_114);
and U122 (N_122,In_229,In_705);
and U123 (N_123,In_580,In_353);
nand U124 (N_124,In_661,In_24);
or U125 (N_125,In_134,In_443);
and U126 (N_126,In_376,In_400);
nor U127 (N_127,In_454,In_78);
or U128 (N_128,In_465,In_30);
or U129 (N_129,In_25,In_275);
nand U130 (N_130,In_590,In_730);
or U131 (N_131,In_637,In_246);
nand U132 (N_132,In_342,In_528);
nand U133 (N_133,In_51,In_694);
or U134 (N_134,In_426,In_700);
or U135 (N_135,In_89,In_43);
or U136 (N_136,In_146,In_128);
nand U137 (N_137,In_498,In_20);
nand U138 (N_138,In_506,In_75);
or U139 (N_139,In_115,In_551);
nand U140 (N_140,In_65,In_123);
nand U141 (N_141,In_10,In_188);
nand U142 (N_142,In_262,In_499);
nand U143 (N_143,In_600,In_337);
nor U144 (N_144,In_125,In_545);
and U145 (N_145,In_535,In_445);
nor U146 (N_146,In_393,In_607);
xnor U147 (N_147,In_126,In_312);
nand U148 (N_148,In_360,In_438);
nand U149 (N_149,In_330,In_699);
nor U150 (N_150,In_178,In_452);
or U151 (N_151,In_180,In_122);
and U152 (N_152,In_505,In_704);
nor U153 (N_153,In_444,In_478);
nand U154 (N_154,In_559,In_141);
or U155 (N_155,In_627,In_530);
or U156 (N_156,In_41,In_644);
and U157 (N_157,In_38,In_236);
or U158 (N_158,In_735,In_105);
nand U159 (N_159,In_194,In_173);
nor U160 (N_160,In_354,In_521);
nor U161 (N_161,In_130,In_595);
and U162 (N_162,In_663,In_531);
nand U163 (N_163,In_685,In_620);
or U164 (N_164,In_62,In_351);
nor U165 (N_165,In_182,In_394);
or U166 (N_166,In_435,In_183);
nand U167 (N_167,In_254,In_339);
nand U168 (N_168,In_411,In_235);
nand U169 (N_169,In_338,In_255);
and U170 (N_170,In_54,In_579);
nor U171 (N_171,In_313,In_494);
and U172 (N_172,In_570,In_131);
and U173 (N_173,In_206,In_733);
nor U174 (N_174,In_523,In_94);
nand U175 (N_175,In_665,In_749);
or U176 (N_176,In_208,In_542);
nor U177 (N_177,In_238,In_296);
nor U178 (N_178,In_550,In_520);
and U179 (N_179,In_343,In_477);
and U180 (N_180,In_650,In_19);
nor U181 (N_181,In_697,In_482);
nand U182 (N_182,In_633,In_391);
or U183 (N_183,In_717,In_631);
or U184 (N_184,In_42,In_596);
nand U185 (N_185,In_34,In_149);
nor U186 (N_186,In_59,In_480);
nor U187 (N_187,In_226,In_158);
nand U188 (N_188,In_686,In_319);
nand U189 (N_189,In_747,In_508);
nand U190 (N_190,In_615,In_748);
nand U191 (N_191,In_40,In_587);
nor U192 (N_192,In_245,In_558);
nand U193 (N_193,In_233,In_513);
nand U194 (N_194,In_635,In_72);
nor U195 (N_195,In_622,In_583);
and U196 (N_196,In_564,In_647);
and U197 (N_197,In_28,In_453);
or U198 (N_198,In_29,In_616);
or U199 (N_199,In_68,In_678);
nand U200 (N_200,In_711,In_457);
and U201 (N_201,In_61,In_147);
nor U202 (N_202,In_405,In_403);
or U203 (N_203,In_710,In_614);
nor U204 (N_204,In_725,In_327);
nand U205 (N_205,In_646,In_58);
and U206 (N_206,In_431,In_186);
nor U207 (N_207,In_459,In_323);
nand U208 (N_208,In_537,In_576);
xnor U209 (N_209,In_632,In_458);
or U210 (N_210,In_563,In_240);
xor U211 (N_211,In_555,In_16);
nand U212 (N_212,In_703,In_348);
nand U213 (N_213,In_574,In_264);
nand U214 (N_214,In_538,In_198);
nand U215 (N_215,In_282,In_6);
nor U216 (N_216,In_96,In_250);
nor U217 (N_217,In_447,In_451);
and U218 (N_218,In_715,In_658);
nor U219 (N_219,In_669,In_304);
and U220 (N_220,In_145,In_116);
and U221 (N_221,In_227,In_302);
nand U222 (N_222,In_77,In_594);
nand U223 (N_223,In_159,In_278);
or U224 (N_224,In_514,In_166);
or U225 (N_225,In_532,In_696);
and U226 (N_226,In_388,In_196);
and U227 (N_227,In_209,In_569);
or U228 (N_228,In_32,In_175);
and U229 (N_229,In_389,In_604);
nor U230 (N_230,In_370,In_82);
nand U231 (N_231,In_516,In_399);
nand U232 (N_232,In_318,In_120);
nor U233 (N_233,In_561,In_0);
and U234 (N_234,In_190,In_643);
and U235 (N_235,In_118,In_8);
and U236 (N_236,In_14,In_192);
nor U237 (N_237,In_548,In_371);
nor U238 (N_238,In_35,In_334);
nand U239 (N_239,In_543,In_124);
and U240 (N_240,In_303,In_695);
nor U241 (N_241,In_565,In_464);
nand U242 (N_242,In_397,In_121);
nor U243 (N_243,In_301,In_618);
or U244 (N_244,In_427,In_651);
or U245 (N_245,In_628,In_69);
nor U246 (N_246,In_155,In_741);
nor U247 (N_247,In_44,In_467);
nor U248 (N_248,In_90,In_271);
and U249 (N_249,In_204,In_413);
nand U250 (N_250,In_743,In_676);
or U251 (N_251,In_724,In_112);
or U252 (N_252,In_88,In_640);
nand U253 (N_253,In_174,In_362);
xor U254 (N_254,In_210,In_571);
nand U255 (N_255,In_22,In_659);
or U256 (N_256,In_554,In_642);
nand U257 (N_257,In_502,In_534);
or U258 (N_258,In_55,In_97);
or U259 (N_259,In_53,In_252);
nand U260 (N_260,In_455,In_446);
and U261 (N_261,In_366,In_701);
nor U262 (N_262,In_27,In_382);
or U263 (N_263,In_64,In_212);
nor U264 (N_264,In_315,In_617);
and U265 (N_265,In_26,In_157);
and U266 (N_266,In_473,In_142);
and U267 (N_267,In_599,In_276);
and U268 (N_268,In_199,In_261);
or U269 (N_269,In_263,In_73);
or U270 (N_270,In_352,In_57);
and U271 (N_271,In_423,In_687);
nor U272 (N_272,In_1,In_67);
nand U273 (N_273,In_623,In_708);
nand U274 (N_274,In_222,In_726);
nor U275 (N_275,In_184,In_522);
or U276 (N_276,In_684,In_670);
nand U277 (N_277,In_462,In_439);
nand U278 (N_278,In_578,In_317);
nor U279 (N_279,In_99,In_39);
or U280 (N_280,In_84,In_466);
or U281 (N_281,In_13,In_290);
or U282 (N_282,In_515,In_300);
nand U283 (N_283,In_385,In_492);
and U284 (N_284,In_641,In_265);
nor U285 (N_285,In_232,In_269);
nor U286 (N_286,In_496,In_433);
xnor U287 (N_287,In_481,In_213);
nor U288 (N_288,In_483,In_162);
or U289 (N_289,In_4,In_612);
nand U290 (N_290,In_167,In_283);
xor U291 (N_291,In_168,In_712);
nand U292 (N_292,In_241,In_386);
nand U293 (N_293,In_171,In_101);
or U294 (N_294,In_624,In_398);
or U295 (N_295,In_197,In_270);
and U296 (N_296,In_510,In_666);
nand U297 (N_297,In_23,In_474);
nor U298 (N_298,In_549,In_259);
and U299 (N_299,In_176,In_37);
or U300 (N_300,In_533,In_298);
and U301 (N_301,In_429,In_488);
and U302 (N_302,In_740,In_557);
nor U303 (N_303,In_468,In_247);
or U304 (N_304,In_668,In_100);
nand U305 (N_305,In_415,In_117);
or U306 (N_306,In_373,In_202);
nor U307 (N_307,In_582,In_390);
or U308 (N_308,In_437,In_331);
nand U309 (N_309,In_215,In_421);
nor U310 (N_310,In_375,In_3);
or U311 (N_311,In_369,In_225);
and U312 (N_312,In_680,In_424);
and U313 (N_313,In_547,In_503);
nor U314 (N_314,In_575,In_83);
or U315 (N_315,In_719,In_436);
nand U316 (N_316,In_172,In_593);
nor U317 (N_317,In_310,In_653);
nor U318 (N_318,In_556,In_297);
xnor U319 (N_319,In_419,In_135);
nor U320 (N_320,In_156,In_367);
nor U321 (N_321,In_293,In_363);
or U322 (N_322,In_322,In_284);
and U323 (N_323,In_608,In_289);
or U324 (N_324,In_266,In_335);
or U325 (N_325,In_308,In_164);
and U326 (N_326,In_358,In_234);
nor U327 (N_327,In_107,In_517);
nand U328 (N_328,In_408,In_688);
or U329 (N_329,In_707,In_396);
nor U330 (N_330,In_281,In_512);
and U331 (N_331,In_86,In_21);
and U332 (N_332,In_239,In_654);
nor U333 (N_333,In_721,In_728);
nor U334 (N_334,In_60,In_244);
or U335 (N_335,In_621,In_469);
nand U336 (N_336,In_723,In_674);
nand U337 (N_337,In_66,In_671);
xnor U338 (N_338,In_527,In_102);
or U339 (N_339,In_731,In_392);
nand U340 (N_340,In_324,In_193);
nand U341 (N_341,In_280,In_187);
and U342 (N_342,In_195,In_560);
or U343 (N_343,In_103,In_404);
or U344 (N_344,In_355,In_81);
and U345 (N_345,In_12,In_493);
or U346 (N_346,In_154,In_401);
or U347 (N_347,In_132,In_374);
nand U348 (N_348,In_379,In_295);
and U349 (N_349,In_485,In_655);
nor U350 (N_350,In_461,In_589);
nand U351 (N_351,In_129,In_497);
and U352 (N_352,In_692,In_407);
nand U353 (N_353,In_71,In_380);
nand U354 (N_354,In_127,In_18);
and U355 (N_355,In_365,In_91);
nand U356 (N_356,In_706,In_490);
nand U357 (N_357,In_693,In_260);
nor U358 (N_358,In_577,In_349);
and U359 (N_359,In_219,In_737);
nand U360 (N_360,In_552,In_744);
nand U361 (N_361,In_610,In_689);
and U362 (N_362,In_288,In_169);
nor U363 (N_363,In_416,In_603);
or U364 (N_364,In_690,In_344);
nor U365 (N_365,In_46,In_108);
nand U366 (N_366,In_211,In_291);
or U367 (N_367,In_378,In_566);
nand U368 (N_368,In_95,In_185);
nor U369 (N_369,In_484,In_272);
and U370 (N_370,In_406,In_486);
nand U371 (N_371,In_148,In_256);
or U372 (N_372,In_314,In_410);
xnor U373 (N_373,In_734,In_525);
and U374 (N_374,In_605,In_7);
and U375 (N_375,In_566,In_30);
nor U376 (N_376,In_720,In_55);
or U377 (N_377,In_550,In_631);
or U378 (N_378,In_710,In_626);
nor U379 (N_379,In_102,In_710);
or U380 (N_380,In_86,In_164);
nand U381 (N_381,In_493,In_96);
nand U382 (N_382,In_166,In_542);
nor U383 (N_383,In_682,In_0);
or U384 (N_384,In_119,In_557);
and U385 (N_385,In_573,In_20);
nor U386 (N_386,In_0,In_228);
or U387 (N_387,In_712,In_243);
nand U388 (N_388,In_356,In_641);
or U389 (N_389,In_628,In_15);
xnor U390 (N_390,In_706,In_188);
nand U391 (N_391,In_702,In_574);
and U392 (N_392,In_537,In_217);
nor U393 (N_393,In_35,In_284);
nor U394 (N_394,In_230,In_151);
or U395 (N_395,In_659,In_153);
or U396 (N_396,In_82,In_689);
and U397 (N_397,In_226,In_302);
nand U398 (N_398,In_475,In_725);
and U399 (N_399,In_367,In_161);
or U400 (N_400,In_661,In_71);
nor U401 (N_401,In_35,In_248);
and U402 (N_402,In_1,In_292);
and U403 (N_403,In_50,In_711);
or U404 (N_404,In_449,In_149);
or U405 (N_405,In_442,In_645);
or U406 (N_406,In_424,In_318);
or U407 (N_407,In_716,In_465);
and U408 (N_408,In_219,In_2);
xnor U409 (N_409,In_77,In_566);
nand U410 (N_410,In_117,In_298);
nor U411 (N_411,In_504,In_317);
nand U412 (N_412,In_491,In_258);
nor U413 (N_413,In_672,In_567);
nand U414 (N_414,In_535,In_229);
nor U415 (N_415,In_329,In_601);
or U416 (N_416,In_516,In_540);
nand U417 (N_417,In_579,In_472);
and U418 (N_418,In_466,In_677);
and U419 (N_419,In_38,In_287);
and U420 (N_420,In_229,In_746);
and U421 (N_421,In_418,In_318);
and U422 (N_422,In_129,In_388);
nand U423 (N_423,In_125,In_715);
nand U424 (N_424,In_300,In_249);
nand U425 (N_425,In_353,In_571);
and U426 (N_426,In_710,In_318);
or U427 (N_427,In_126,In_340);
nand U428 (N_428,In_522,In_736);
nand U429 (N_429,In_585,In_641);
nand U430 (N_430,In_271,In_505);
nor U431 (N_431,In_511,In_118);
and U432 (N_432,In_552,In_22);
or U433 (N_433,In_200,In_515);
xnor U434 (N_434,In_294,In_565);
nor U435 (N_435,In_368,In_554);
nand U436 (N_436,In_465,In_422);
or U437 (N_437,In_729,In_261);
nand U438 (N_438,In_524,In_19);
xor U439 (N_439,In_473,In_688);
xor U440 (N_440,In_86,In_705);
nor U441 (N_441,In_140,In_173);
nor U442 (N_442,In_4,In_352);
and U443 (N_443,In_49,In_697);
or U444 (N_444,In_342,In_20);
nor U445 (N_445,In_223,In_549);
nand U446 (N_446,In_526,In_646);
nor U447 (N_447,In_171,In_335);
or U448 (N_448,In_46,In_555);
nand U449 (N_449,In_617,In_744);
or U450 (N_450,In_10,In_664);
and U451 (N_451,In_652,In_62);
or U452 (N_452,In_592,In_494);
and U453 (N_453,In_745,In_698);
nand U454 (N_454,In_671,In_665);
nor U455 (N_455,In_596,In_133);
nor U456 (N_456,In_260,In_409);
or U457 (N_457,In_573,In_418);
and U458 (N_458,In_124,In_638);
nand U459 (N_459,In_577,In_510);
or U460 (N_460,In_679,In_373);
nand U461 (N_461,In_115,In_457);
nand U462 (N_462,In_125,In_115);
nor U463 (N_463,In_711,In_512);
nor U464 (N_464,In_538,In_711);
and U465 (N_465,In_553,In_197);
xnor U466 (N_466,In_48,In_415);
and U467 (N_467,In_368,In_660);
nor U468 (N_468,In_745,In_411);
nand U469 (N_469,In_174,In_286);
or U470 (N_470,In_414,In_267);
nor U471 (N_471,In_539,In_366);
or U472 (N_472,In_115,In_150);
and U473 (N_473,In_436,In_517);
or U474 (N_474,In_505,In_721);
or U475 (N_475,In_535,In_722);
or U476 (N_476,In_571,In_416);
nand U477 (N_477,In_149,In_120);
and U478 (N_478,In_293,In_31);
nand U479 (N_479,In_27,In_302);
and U480 (N_480,In_319,In_499);
and U481 (N_481,In_70,In_397);
or U482 (N_482,In_317,In_599);
or U483 (N_483,In_520,In_564);
or U484 (N_484,In_21,In_627);
nor U485 (N_485,In_87,In_309);
or U486 (N_486,In_694,In_193);
nand U487 (N_487,In_428,In_373);
and U488 (N_488,In_369,In_524);
nor U489 (N_489,In_348,In_459);
or U490 (N_490,In_117,In_50);
and U491 (N_491,In_466,In_73);
xnor U492 (N_492,In_314,In_13);
and U493 (N_493,In_239,In_218);
and U494 (N_494,In_484,In_28);
nor U495 (N_495,In_81,In_578);
nor U496 (N_496,In_686,In_84);
and U497 (N_497,In_633,In_418);
or U498 (N_498,In_18,In_503);
nand U499 (N_499,In_652,In_359);
or U500 (N_500,In_363,In_261);
nor U501 (N_501,In_657,In_316);
and U502 (N_502,In_54,In_59);
nand U503 (N_503,In_599,In_422);
nor U504 (N_504,In_723,In_15);
nand U505 (N_505,In_510,In_65);
or U506 (N_506,In_569,In_36);
nor U507 (N_507,In_164,In_110);
nand U508 (N_508,In_389,In_739);
nand U509 (N_509,In_145,In_160);
nand U510 (N_510,In_46,In_381);
nor U511 (N_511,In_80,In_591);
xor U512 (N_512,In_332,In_418);
and U513 (N_513,In_554,In_218);
and U514 (N_514,In_280,In_490);
nor U515 (N_515,In_327,In_21);
nor U516 (N_516,In_566,In_32);
and U517 (N_517,In_519,In_125);
and U518 (N_518,In_85,In_405);
or U519 (N_519,In_723,In_661);
nor U520 (N_520,In_597,In_744);
or U521 (N_521,In_51,In_592);
and U522 (N_522,In_745,In_687);
or U523 (N_523,In_113,In_693);
and U524 (N_524,In_199,In_407);
nand U525 (N_525,In_97,In_607);
nor U526 (N_526,In_447,In_731);
and U527 (N_527,In_416,In_602);
or U528 (N_528,In_134,In_397);
and U529 (N_529,In_231,In_575);
and U530 (N_530,In_680,In_91);
nor U531 (N_531,In_422,In_122);
nor U532 (N_532,In_282,In_138);
or U533 (N_533,In_152,In_344);
and U534 (N_534,In_507,In_719);
nand U535 (N_535,In_481,In_629);
nor U536 (N_536,In_303,In_336);
nand U537 (N_537,In_665,In_233);
nor U538 (N_538,In_256,In_497);
nand U539 (N_539,In_89,In_37);
nand U540 (N_540,In_227,In_629);
nor U541 (N_541,In_375,In_472);
nand U542 (N_542,In_465,In_168);
nor U543 (N_543,In_115,In_67);
nor U544 (N_544,In_313,In_454);
nand U545 (N_545,In_558,In_680);
and U546 (N_546,In_20,In_350);
nor U547 (N_547,In_627,In_340);
and U548 (N_548,In_91,In_469);
nor U549 (N_549,In_381,In_698);
or U550 (N_550,In_587,In_353);
or U551 (N_551,In_731,In_280);
nor U552 (N_552,In_20,In_717);
nor U553 (N_553,In_460,In_112);
nor U554 (N_554,In_287,In_250);
nor U555 (N_555,In_637,In_330);
and U556 (N_556,In_377,In_528);
nor U557 (N_557,In_221,In_692);
or U558 (N_558,In_155,In_603);
and U559 (N_559,In_548,In_545);
nor U560 (N_560,In_613,In_439);
and U561 (N_561,In_10,In_494);
nand U562 (N_562,In_522,In_391);
nor U563 (N_563,In_719,In_35);
and U564 (N_564,In_519,In_102);
nand U565 (N_565,In_225,In_32);
nand U566 (N_566,In_603,In_263);
and U567 (N_567,In_404,In_295);
nand U568 (N_568,In_145,In_154);
or U569 (N_569,In_731,In_27);
nor U570 (N_570,In_322,In_10);
nor U571 (N_571,In_643,In_479);
and U572 (N_572,In_320,In_629);
nand U573 (N_573,In_425,In_496);
or U574 (N_574,In_269,In_78);
or U575 (N_575,In_680,In_312);
or U576 (N_576,In_731,In_611);
and U577 (N_577,In_255,In_115);
or U578 (N_578,In_219,In_572);
or U579 (N_579,In_641,In_304);
and U580 (N_580,In_289,In_668);
nor U581 (N_581,In_195,In_606);
and U582 (N_582,In_54,In_530);
nor U583 (N_583,In_393,In_119);
nand U584 (N_584,In_59,In_247);
or U585 (N_585,In_623,In_123);
or U586 (N_586,In_268,In_568);
nor U587 (N_587,In_377,In_720);
nor U588 (N_588,In_60,In_602);
and U589 (N_589,In_440,In_513);
nor U590 (N_590,In_32,In_160);
nand U591 (N_591,In_507,In_22);
nor U592 (N_592,In_126,In_210);
and U593 (N_593,In_553,In_398);
nand U594 (N_594,In_608,In_61);
and U595 (N_595,In_428,In_198);
and U596 (N_596,In_724,In_489);
nor U597 (N_597,In_437,In_241);
or U598 (N_598,In_334,In_84);
or U599 (N_599,In_398,In_637);
and U600 (N_600,In_262,In_150);
or U601 (N_601,In_219,In_471);
nand U602 (N_602,In_353,In_197);
or U603 (N_603,In_160,In_684);
or U604 (N_604,In_217,In_225);
nand U605 (N_605,In_164,In_230);
nand U606 (N_606,In_231,In_460);
nor U607 (N_607,In_631,In_495);
or U608 (N_608,In_623,In_400);
or U609 (N_609,In_258,In_379);
nor U610 (N_610,In_488,In_504);
and U611 (N_611,In_62,In_112);
nand U612 (N_612,In_565,In_231);
or U613 (N_613,In_738,In_87);
or U614 (N_614,In_681,In_629);
nand U615 (N_615,In_583,In_222);
and U616 (N_616,In_337,In_413);
or U617 (N_617,In_58,In_651);
nand U618 (N_618,In_579,In_58);
nand U619 (N_619,In_390,In_11);
nand U620 (N_620,In_240,In_48);
and U621 (N_621,In_413,In_472);
or U622 (N_622,In_151,In_331);
nor U623 (N_623,In_19,In_380);
nand U624 (N_624,In_1,In_722);
nand U625 (N_625,In_587,In_660);
nand U626 (N_626,In_449,In_366);
or U627 (N_627,In_220,In_660);
or U628 (N_628,In_66,In_96);
and U629 (N_629,In_607,In_330);
and U630 (N_630,In_305,In_232);
and U631 (N_631,In_75,In_127);
nand U632 (N_632,In_14,In_651);
and U633 (N_633,In_170,In_272);
or U634 (N_634,In_368,In_28);
and U635 (N_635,In_137,In_679);
and U636 (N_636,In_682,In_667);
nand U637 (N_637,In_353,In_412);
nand U638 (N_638,In_205,In_500);
or U639 (N_639,In_120,In_146);
and U640 (N_640,In_356,In_447);
and U641 (N_641,In_146,In_594);
or U642 (N_642,In_98,In_199);
or U643 (N_643,In_536,In_580);
and U644 (N_644,In_67,In_612);
nor U645 (N_645,In_535,In_162);
or U646 (N_646,In_170,In_620);
nand U647 (N_647,In_649,In_617);
or U648 (N_648,In_146,In_226);
nor U649 (N_649,In_443,In_27);
nor U650 (N_650,In_341,In_282);
nor U651 (N_651,In_26,In_748);
nand U652 (N_652,In_57,In_465);
and U653 (N_653,In_636,In_122);
nor U654 (N_654,In_211,In_186);
nor U655 (N_655,In_595,In_462);
or U656 (N_656,In_388,In_244);
and U657 (N_657,In_257,In_323);
or U658 (N_658,In_580,In_195);
nand U659 (N_659,In_75,In_184);
and U660 (N_660,In_731,In_256);
nor U661 (N_661,In_595,In_573);
or U662 (N_662,In_365,In_151);
nand U663 (N_663,In_428,In_553);
nand U664 (N_664,In_265,In_742);
nand U665 (N_665,In_116,In_164);
nor U666 (N_666,In_99,In_186);
xnor U667 (N_667,In_276,In_715);
or U668 (N_668,In_25,In_334);
nor U669 (N_669,In_38,In_74);
nand U670 (N_670,In_274,In_602);
nand U671 (N_671,In_181,In_467);
nand U672 (N_672,In_480,In_507);
nor U673 (N_673,In_481,In_181);
and U674 (N_674,In_442,In_341);
and U675 (N_675,In_690,In_555);
and U676 (N_676,In_645,In_343);
or U677 (N_677,In_748,In_709);
nor U678 (N_678,In_478,In_164);
xnor U679 (N_679,In_232,In_574);
nand U680 (N_680,In_592,In_700);
nand U681 (N_681,In_151,In_75);
nor U682 (N_682,In_106,In_456);
nand U683 (N_683,In_379,In_744);
and U684 (N_684,In_418,In_304);
nand U685 (N_685,In_251,In_310);
or U686 (N_686,In_726,In_599);
or U687 (N_687,In_31,In_713);
or U688 (N_688,In_740,In_554);
or U689 (N_689,In_64,In_245);
or U690 (N_690,In_47,In_48);
or U691 (N_691,In_480,In_301);
or U692 (N_692,In_383,In_626);
nor U693 (N_693,In_638,In_323);
nor U694 (N_694,In_75,In_571);
or U695 (N_695,In_179,In_312);
nand U696 (N_696,In_451,In_88);
or U697 (N_697,In_400,In_89);
nand U698 (N_698,In_455,In_519);
and U699 (N_699,In_40,In_674);
or U700 (N_700,In_154,In_175);
xor U701 (N_701,In_679,In_608);
and U702 (N_702,In_597,In_59);
and U703 (N_703,In_224,In_513);
and U704 (N_704,In_461,In_619);
or U705 (N_705,In_141,In_607);
and U706 (N_706,In_293,In_327);
nor U707 (N_707,In_706,In_422);
nor U708 (N_708,In_326,In_493);
nor U709 (N_709,In_744,In_172);
and U710 (N_710,In_432,In_375);
and U711 (N_711,In_672,In_461);
or U712 (N_712,In_410,In_22);
nand U713 (N_713,In_220,In_133);
and U714 (N_714,In_543,In_218);
nor U715 (N_715,In_194,In_522);
nor U716 (N_716,In_592,In_635);
nor U717 (N_717,In_110,In_234);
nor U718 (N_718,In_623,In_62);
nand U719 (N_719,In_584,In_10);
nor U720 (N_720,In_462,In_336);
xor U721 (N_721,In_8,In_116);
and U722 (N_722,In_25,In_242);
and U723 (N_723,In_624,In_322);
and U724 (N_724,In_661,In_576);
or U725 (N_725,In_265,In_686);
or U726 (N_726,In_61,In_155);
or U727 (N_727,In_735,In_553);
and U728 (N_728,In_364,In_66);
nor U729 (N_729,In_445,In_400);
and U730 (N_730,In_65,In_120);
xnor U731 (N_731,In_355,In_327);
or U732 (N_732,In_218,In_629);
or U733 (N_733,In_86,In_182);
nand U734 (N_734,In_647,In_650);
or U735 (N_735,In_443,In_433);
nor U736 (N_736,In_65,In_483);
nand U737 (N_737,In_193,In_236);
nor U738 (N_738,In_271,In_700);
nor U739 (N_739,In_488,In_661);
nor U740 (N_740,In_350,In_310);
and U741 (N_741,In_377,In_223);
xor U742 (N_742,In_409,In_625);
and U743 (N_743,In_21,In_737);
and U744 (N_744,In_266,In_536);
nor U745 (N_745,In_137,In_579);
nor U746 (N_746,In_689,In_504);
or U747 (N_747,In_498,In_87);
or U748 (N_748,In_743,In_40);
nor U749 (N_749,In_678,In_274);
or U750 (N_750,In_470,In_66);
nor U751 (N_751,In_659,In_654);
or U752 (N_752,In_527,In_703);
or U753 (N_753,In_268,In_329);
nor U754 (N_754,In_25,In_490);
nor U755 (N_755,In_310,In_449);
and U756 (N_756,In_212,In_472);
or U757 (N_757,In_310,In_334);
nand U758 (N_758,In_603,In_391);
nor U759 (N_759,In_23,In_67);
nand U760 (N_760,In_499,In_706);
nand U761 (N_761,In_168,In_71);
nor U762 (N_762,In_662,In_334);
nand U763 (N_763,In_585,In_552);
and U764 (N_764,In_419,In_351);
and U765 (N_765,In_514,In_466);
or U766 (N_766,In_169,In_258);
nand U767 (N_767,In_257,In_595);
or U768 (N_768,In_725,In_482);
and U769 (N_769,In_112,In_428);
nor U770 (N_770,In_385,In_741);
nor U771 (N_771,In_741,In_553);
or U772 (N_772,In_346,In_352);
or U773 (N_773,In_580,In_7);
and U774 (N_774,In_478,In_734);
and U775 (N_775,In_106,In_227);
nand U776 (N_776,In_344,In_260);
and U777 (N_777,In_66,In_31);
or U778 (N_778,In_216,In_358);
and U779 (N_779,In_680,In_700);
nand U780 (N_780,In_719,In_306);
or U781 (N_781,In_749,In_748);
nand U782 (N_782,In_746,In_182);
nand U783 (N_783,In_192,In_496);
or U784 (N_784,In_48,In_371);
and U785 (N_785,In_510,In_520);
or U786 (N_786,In_467,In_512);
nor U787 (N_787,In_261,In_611);
or U788 (N_788,In_224,In_418);
xnor U789 (N_789,In_285,In_294);
and U790 (N_790,In_75,In_138);
or U791 (N_791,In_561,In_569);
nor U792 (N_792,In_704,In_731);
nand U793 (N_793,In_670,In_81);
nor U794 (N_794,In_453,In_233);
or U795 (N_795,In_359,In_610);
nor U796 (N_796,In_68,In_634);
nor U797 (N_797,In_177,In_333);
and U798 (N_798,In_276,In_171);
nand U799 (N_799,In_241,In_567);
xor U800 (N_800,In_231,In_643);
nor U801 (N_801,In_591,In_475);
nor U802 (N_802,In_517,In_0);
or U803 (N_803,In_466,In_443);
or U804 (N_804,In_726,In_325);
and U805 (N_805,In_501,In_444);
or U806 (N_806,In_398,In_71);
and U807 (N_807,In_632,In_659);
nand U808 (N_808,In_480,In_4);
nand U809 (N_809,In_46,In_508);
nand U810 (N_810,In_82,In_192);
nand U811 (N_811,In_196,In_359);
nand U812 (N_812,In_524,In_430);
nor U813 (N_813,In_414,In_69);
nor U814 (N_814,In_690,In_708);
or U815 (N_815,In_162,In_449);
nand U816 (N_816,In_521,In_22);
and U817 (N_817,In_708,In_309);
nor U818 (N_818,In_471,In_316);
nand U819 (N_819,In_665,In_640);
or U820 (N_820,In_603,In_635);
and U821 (N_821,In_296,In_692);
and U822 (N_822,In_713,In_189);
and U823 (N_823,In_659,In_209);
and U824 (N_824,In_191,In_672);
or U825 (N_825,In_543,In_642);
xor U826 (N_826,In_415,In_216);
and U827 (N_827,In_206,In_0);
nand U828 (N_828,In_491,In_619);
and U829 (N_829,In_211,In_437);
or U830 (N_830,In_117,In_326);
and U831 (N_831,In_590,In_709);
and U832 (N_832,In_552,In_43);
or U833 (N_833,In_412,In_211);
nand U834 (N_834,In_486,In_177);
nand U835 (N_835,In_425,In_421);
nand U836 (N_836,In_19,In_512);
nor U837 (N_837,In_145,In_542);
nand U838 (N_838,In_581,In_626);
or U839 (N_839,In_259,In_499);
nor U840 (N_840,In_373,In_185);
nor U841 (N_841,In_450,In_320);
nor U842 (N_842,In_484,In_696);
nor U843 (N_843,In_103,In_504);
nor U844 (N_844,In_356,In_65);
nor U845 (N_845,In_413,In_24);
or U846 (N_846,In_314,In_135);
nand U847 (N_847,In_319,In_628);
nor U848 (N_848,In_247,In_507);
or U849 (N_849,In_644,In_87);
or U850 (N_850,In_343,In_638);
and U851 (N_851,In_658,In_597);
or U852 (N_852,In_528,In_293);
nand U853 (N_853,In_748,In_48);
nor U854 (N_854,In_301,In_634);
nand U855 (N_855,In_212,In_655);
or U856 (N_856,In_648,In_569);
nand U857 (N_857,In_642,In_129);
or U858 (N_858,In_611,In_268);
and U859 (N_859,In_103,In_499);
or U860 (N_860,In_270,In_721);
nand U861 (N_861,In_192,In_457);
and U862 (N_862,In_57,In_368);
nand U863 (N_863,In_8,In_653);
nand U864 (N_864,In_59,In_658);
or U865 (N_865,In_130,In_106);
or U866 (N_866,In_454,In_580);
or U867 (N_867,In_124,In_142);
nor U868 (N_868,In_344,In_114);
xnor U869 (N_869,In_3,In_0);
and U870 (N_870,In_737,In_387);
nor U871 (N_871,In_446,In_480);
nor U872 (N_872,In_28,In_138);
nor U873 (N_873,In_702,In_634);
nor U874 (N_874,In_480,In_468);
nand U875 (N_875,In_575,In_687);
nand U876 (N_876,In_455,In_498);
nor U877 (N_877,In_368,In_701);
and U878 (N_878,In_311,In_710);
and U879 (N_879,In_562,In_733);
or U880 (N_880,In_612,In_234);
or U881 (N_881,In_717,In_541);
and U882 (N_882,In_407,In_296);
nand U883 (N_883,In_243,In_567);
or U884 (N_884,In_491,In_462);
and U885 (N_885,In_735,In_497);
nor U886 (N_886,In_23,In_3);
nand U887 (N_887,In_550,In_48);
and U888 (N_888,In_293,In_445);
nor U889 (N_889,In_164,In_744);
nor U890 (N_890,In_48,In_430);
nand U891 (N_891,In_706,In_256);
or U892 (N_892,In_304,In_353);
and U893 (N_893,In_262,In_74);
or U894 (N_894,In_315,In_77);
and U895 (N_895,In_120,In_292);
nor U896 (N_896,In_602,In_7);
nor U897 (N_897,In_612,In_534);
or U898 (N_898,In_116,In_663);
nor U899 (N_899,In_703,In_672);
and U900 (N_900,In_51,In_468);
and U901 (N_901,In_204,In_182);
nor U902 (N_902,In_136,In_425);
or U903 (N_903,In_595,In_296);
or U904 (N_904,In_608,In_517);
or U905 (N_905,In_652,In_49);
nand U906 (N_906,In_409,In_502);
nand U907 (N_907,In_619,In_51);
nor U908 (N_908,In_346,In_53);
or U909 (N_909,In_466,In_661);
nor U910 (N_910,In_392,In_691);
nor U911 (N_911,In_490,In_257);
nand U912 (N_912,In_27,In_378);
nand U913 (N_913,In_475,In_366);
or U914 (N_914,In_2,In_154);
and U915 (N_915,In_194,In_481);
nand U916 (N_916,In_634,In_708);
and U917 (N_917,In_309,In_53);
or U918 (N_918,In_280,In_544);
nand U919 (N_919,In_133,In_341);
and U920 (N_920,In_191,In_249);
and U921 (N_921,In_620,In_624);
nand U922 (N_922,In_259,In_632);
or U923 (N_923,In_265,In_25);
or U924 (N_924,In_673,In_318);
nor U925 (N_925,In_13,In_492);
or U926 (N_926,In_576,In_78);
nand U927 (N_927,In_277,In_659);
and U928 (N_928,In_182,In_636);
nand U929 (N_929,In_724,In_723);
nand U930 (N_930,In_280,In_484);
and U931 (N_931,In_272,In_62);
or U932 (N_932,In_498,In_537);
nor U933 (N_933,In_441,In_749);
or U934 (N_934,In_351,In_94);
nor U935 (N_935,In_463,In_107);
nor U936 (N_936,In_515,In_482);
nand U937 (N_937,In_222,In_243);
and U938 (N_938,In_469,In_414);
and U939 (N_939,In_549,In_6);
and U940 (N_940,In_183,In_176);
and U941 (N_941,In_317,In_696);
nand U942 (N_942,In_486,In_163);
nor U943 (N_943,In_517,In_747);
and U944 (N_944,In_332,In_64);
nand U945 (N_945,In_423,In_85);
and U946 (N_946,In_8,In_641);
and U947 (N_947,In_261,In_250);
nand U948 (N_948,In_516,In_328);
nand U949 (N_949,In_106,In_407);
nand U950 (N_950,In_80,In_614);
nor U951 (N_951,In_266,In_556);
nand U952 (N_952,In_699,In_486);
nor U953 (N_953,In_492,In_306);
nor U954 (N_954,In_277,In_454);
nand U955 (N_955,In_110,In_91);
nand U956 (N_956,In_190,In_562);
and U957 (N_957,In_72,In_420);
and U958 (N_958,In_177,In_394);
or U959 (N_959,In_49,In_576);
xor U960 (N_960,In_639,In_278);
nor U961 (N_961,In_481,In_372);
and U962 (N_962,In_599,In_177);
or U963 (N_963,In_209,In_358);
or U964 (N_964,In_545,In_268);
and U965 (N_965,In_24,In_180);
or U966 (N_966,In_718,In_530);
nand U967 (N_967,In_176,In_651);
nor U968 (N_968,In_34,In_162);
and U969 (N_969,In_263,In_535);
and U970 (N_970,In_46,In_341);
nor U971 (N_971,In_10,In_646);
nand U972 (N_972,In_450,In_333);
and U973 (N_973,In_260,In_527);
nor U974 (N_974,In_85,In_184);
and U975 (N_975,In_5,In_688);
nor U976 (N_976,In_340,In_388);
nor U977 (N_977,In_22,In_394);
and U978 (N_978,In_679,In_416);
or U979 (N_979,In_303,In_84);
or U980 (N_980,In_1,In_721);
nand U981 (N_981,In_19,In_187);
and U982 (N_982,In_27,In_542);
and U983 (N_983,In_163,In_506);
nor U984 (N_984,In_314,In_101);
nand U985 (N_985,In_674,In_629);
nand U986 (N_986,In_538,In_73);
and U987 (N_987,In_126,In_526);
or U988 (N_988,In_281,In_494);
nand U989 (N_989,In_426,In_156);
and U990 (N_990,In_213,In_588);
or U991 (N_991,In_72,In_92);
nor U992 (N_992,In_690,In_194);
nor U993 (N_993,In_699,In_508);
and U994 (N_994,In_649,In_36);
nor U995 (N_995,In_433,In_28);
nand U996 (N_996,In_580,In_393);
nor U997 (N_997,In_152,In_279);
or U998 (N_998,In_689,In_409);
nand U999 (N_999,In_382,In_303);
nand U1000 (N_1000,N_925,N_50);
nor U1001 (N_1001,N_244,N_69);
or U1002 (N_1002,N_862,N_228);
nor U1003 (N_1003,N_717,N_676);
nand U1004 (N_1004,N_515,N_398);
nor U1005 (N_1005,N_437,N_268);
nand U1006 (N_1006,N_813,N_774);
or U1007 (N_1007,N_696,N_102);
xor U1008 (N_1008,N_903,N_242);
or U1009 (N_1009,N_38,N_389);
nor U1010 (N_1010,N_4,N_543);
or U1011 (N_1011,N_162,N_14);
nor U1012 (N_1012,N_538,N_475);
or U1013 (N_1013,N_189,N_37);
nor U1014 (N_1014,N_690,N_833);
and U1015 (N_1015,N_959,N_718);
and U1016 (N_1016,N_388,N_807);
or U1017 (N_1017,N_140,N_817);
nor U1018 (N_1018,N_122,N_53);
nor U1019 (N_1019,N_514,N_502);
nor U1020 (N_1020,N_148,N_697);
nand U1021 (N_1021,N_555,N_266);
and U1022 (N_1022,N_972,N_313);
and U1023 (N_1023,N_522,N_334);
and U1024 (N_1024,N_631,N_414);
nand U1025 (N_1025,N_84,N_853);
and U1026 (N_1026,N_963,N_33);
or U1027 (N_1027,N_846,N_897);
and U1028 (N_1028,N_149,N_188);
and U1029 (N_1029,N_982,N_308);
nor U1030 (N_1030,N_455,N_165);
nor U1031 (N_1031,N_156,N_668);
nor U1032 (N_1032,N_113,N_971);
nand U1033 (N_1033,N_863,N_539);
nand U1034 (N_1034,N_94,N_454);
or U1035 (N_1035,N_603,N_240);
or U1036 (N_1036,N_594,N_463);
nor U1037 (N_1037,N_536,N_91);
nand U1038 (N_1038,N_426,N_884);
nand U1039 (N_1039,N_915,N_800);
or U1040 (N_1040,N_418,N_721);
and U1041 (N_1041,N_493,N_312);
nand U1042 (N_1042,N_299,N_591);
nor U1043 (N_1043,N_753,N_190);
nor U1044 (N_1044,N_319,N_766);
and U1045 (N_1045,N_896,N_508);
and U1046 (N_1046,N_220,N_970);
and U1047 (N_1047,N_256,N_698);
nor U1048 (N_1048,N_986,N_910);
nand U1049 (N_1049,N_882,N_152);
or U1050 (N_1050,N_518,N_24);
nand U1051 (N_1051,N_890,N_318);
nand U1052 (N_1052,N_699,N_606);
and U1053 (N_1053,N_635,N_841);
nor U1054 (N_1054,N_874,N_615);
nor U1055 (N_1055,N_804,N_117);
nor U1056 (N_1056,N_627,N_579);
nor U1057 (N_1057,N_909,N_547);
nand U1058 (N_1058,N_684,N_99);
or U1059 (N_1059,N_253,N_366);
and U1060 (N_1060,N_649,N_586);
or U1061 (N_1061,N_767,N_947);
and U1062 (N_1062,N_981,N_505);
nand U1063 (N_1063,N_831,N_985);
nand U1064 (N_1064,N_404,N_533);
nor U1065 (N_1065,N_51,N_859);
and U1066 (N_1066,N_664,N_440);
and U1067 (N_1067,N_320,N_961);
and U1068 (N_1068,N_380,N_560);
and U1069 (N_1069,N_123,N_743);
nand U1070 (N_1070,N_783,N_154);
nor U1071 (N_1071,N_714,N_471);
and U1072 (N_1072,N_344,N_923);
or U1073 (N_1073,N_639,N_146);
and U1074 (N_1074,N_737,N_659);
or U1075 (N_1075,N_173,N_731);
nor U1076 (N_1076,N_520,N_584);
and U1077 (N_1077,N_693,N_453);
nor U1078 (N_1078,N_950,N_877);
or U1079 (N_1079,N_893,N_798);
or U1080 (N_1080,N_995,N_331);
nand U1081 (N_1081,N_292,N_397);
nand U1082 (N_1082,N_219,N_781);
nor U1083 (N_1083,N_270,N_337);
and U1084 (N_1084,N_566,N_793);
nor U1085 (N_1085,N_333,N_711);
nor U1086 (N_1086,N_55,N_561);
and U1087 (N_1087,N_772,N_21);
or U1088 (N_1088,N_104,N_726);
nor U1089 (N_1089,N_322,N_166);
nand U1090 (N_1090,N_234,N_215);
or U1091 (N_1091,N_734,N_20);
nor U1092 (N_1092,N_908,N_785);
nand U1093 (N_1093,N_430,N_392);
nor U1094 (N_1094,N_735,N_71);
nand U1095 (N_1095,N_498,N_329);
nand U1096 (N_1096,N_751,N_632);
nor U1097 (N_1097,N_89,N_445);
nor U1098 (N_1098,N_633,N_423);
or U1099 (N_1099,N_282,N_802);
or U1100 (N_1100,N_622,N_809);
nand U1101 (N_1101,N_490,N_439);
or U1102 (N_1102,N_376,N_400);
and U1103 (N_1103,N_938,N_487);
nand U1104 (N_1104,N_503,N_125);
and U1105 (N_1105,N_327,N_265);
nor U1106 (N_1106,N_429,N_980);
and U1107 (N_1107,N_279,N_665);
and U1108 (N_1108,N_480,N_132);
nand U1109 (N_1109,N_210,N_626);
nand U1110 (N_1110,N_250,N_485);
nand U1111 (N_1111,N_306,N_618);
nor U1112 (N_1112,N_760,N_685);
or U1113 (N_1113,N_209,N_629);
nor U1114 (N_1114,N_373,N_382);
or U1115 (N_1115,N_64,N_70);
nor U1116 (N_1116,N_724,N_93);
or U1117 (N_1117,N_174,N_211);
nand U1118 (N_1118,N_421,N_964);
and U1119 (N_1119,N_562,N_954);
and U1120 (N_1120,N_305,N_550);
or U1121 (N_1121,N_224,N_169);
nor U1122 (N_1122,N_596,N_467);
nand U1123 (N_1123,N_276,N_355);
or U1124 (N_1124,N_604,N_66);
and U1125 (N_1125,N_202,N_294);
and U1126 (N_1126,N_311,N_745);
nor U1127 (N_1127,N_630,N_967);
or U1128 (N_1128,N_221,N_9);
nand U1129 (N_1129,N_792,N_450);
and U1130 (N_1130,N_541,N_891);
and U1131 (N_1131,N_80,N_643);
and U1132 (N_1132,N_424,N_694);
and U1133 (N_1133,N_695,N_56);
nand U1134 (N_1134,N_43,N_571);
nand U1135 (N_1135,N_918,N_316);
or U1136 (N_1136,N_435,N_484);
nand U1137 (N_1137,N_624,N_110);
nand U1138 (N_1138,N_290,N_137);
nand U1139 (N_1139,N_275,N_406);
and U1140 (N_1140,N_778,N_675);
or U1141 (N_1141,N_992,N_991);
nand U1142 (N_1142,N_369,N_651);
nand U1143 (N_1143,N_363,N_326);
nand U1144 (N_1144,N_928,N_347);
nor U1145 (N_1145,N_849,N_597);
nor U1146 (N_1146,N_937,N_661);
nand U1147 (N_1147,N_432,N_818);
and U1148 (N_1148,N_246,N_235);
nand U1149 (N_1149,N_496,N_617);
nand U1150 (N_1150,N_76,N_956);
and U1151 (N_1151,N_323,N_481);
and U1152 (N_1152,N_177,N_838);
nor U1153 (N_1153,N_164,N_860);
and U1154 (N_1154,N_703,N_446);
and U1155 (N_1155,N_184,N_226);
or U1156 (N_1156,N_338,N_203);
or U1157 (N_1157,N_978,N_955);
and U1158 (N_1158,N_702,N_864);
or U1159 (N_1159,N_15,N_706);
nand U1160 (N_1160,N_222,N_887);
nor U1161 (N_1161,N_183,N_136);
nand U1162 (N_1162,N_387,N_269);
and U1163 (N_1163,N_569,N_636);
nor U1164 (N_1164,N_851,N_924);
nand U1165 (N_1165,N_207,N_260);
nand U1166 (N_1166,N_867,N_944);
nor U1167 (N_1167,N_18,N_713);
and U1168 (N_1168,N_172,N_705);
and U1169 (N_1169,N_663,N_523);
nor U1170 (N_1170,N_934,N_101);
or U1171 (N_1171,N_739,N_52);
nand U1172 (N_1172,N_88,N_477);
nor U1173 (N_1173,N_328,N_412);
nand U1174 (N_1174,N_29,N_712);
nand U1175 (N_1175,N_332,N_572);
nand U1176 (N_1176,N_150,N_997);
nor U1177 (N_1177,N_625,N_558);
nand U1178 (N_1178,N_36,N_607);
nor U1179 (N_1179,N_57,N_497);
nand U1180 (N_1180,N_286,N_921);
nand U1181 (N_1181,N_79,N_231);
nor U1182 (N_1182,N_720,N_285);
nor U1183 (N_1183,N_782,N_10);
xnor U1184 (N_1184,N_272,N_249);
nand U1185 (N_1185,N_855,N_763);
nor U1186 (N_1186,N_486,N_26);
xor U1187 (N_1187,N_899,N_686);
nand U1188 (N_1188,N_605,N_756);
or U1189 (N_1189,N_86,N_707);
nor U1190 (N_1190,N_92,N_820);
nand U1191 (N_1191,N_529,N_293);
or U1192 (N_1192,N_670,N_787);
or U1193 (N_1193,N_943,N_300);
xor U1194 (N_1194,N_59,N_535);
nor U1195 (N_1195,N_842,N_710);
or U1196 (N_1196,N_405,N_936);
or U1197 (N_1197,N_62,N_931);
and U1198 (N_1198,N_374,N_755);
nand U1199 (N_1199,N_834,N_570);
nand U1200 (N_1200,N_589,N_39);
nor U1201 (N_1201,N_461,N_628);
and U1202 (N_1202,N_768,N_510);
or U1203 (N_1203,N_302,N_794);
and U1204 (N_1204,N_193,N_109);
or U1205 (N_1205,N_602,N_297);
and U1206 (N_1206,N_108,N_100);
or U1207 (N_1207,N_977,N_142);
or U1208 (N_1208,N_213,N_672);
nand U1209 (N_1209,N_201,N_674);
nand U1210 (N_1210,N_314,N_170);
and U1211 (N_1211,N_919,N_770);
xor U1212 (N_1212,N_645,N_749);
nor U1213 (N_1213,N_621,N_677);
nor U1214 (N_1214,N_534,N_63);
nor U1215 (N_1215,N_574,N_390);
and U1216 (N_1216,N_564,N_230);
nor U1217 (N_1217,N_217,N_845);
nand U1218 (N_1218,N_837,N_530);
and U1219 (N_1219,N_35,N_216);
or U1220 (N_1220,N_557,N_524);
or U1221 (N_1221,N_658,N_460);
or U1222 (N_1222,N_264,N_727);
xor U1223 (N_1223,N_638,N_239);
nand U1224 (N_1224,N_957,N_163);
and U1225 (N_1225,N_233,N_948);
or U1226 (N_1226,N_839,N_556);
and U1227 (N_1227,N_719,N_178);
and U1228 (N_1228,N_2,N_462);
nor U1229 (N_1229,N_263,N_973);
and U1230 (N_1230,N_653,N_660);
and U1231 (N_1231,N_195,N_112);
nand U1232 (N_1232,N_124,N_254);
nor U1233 (N_1233,N_689,N_861);
nand U1234 (N_1234,N_22,N_715);
or U1235 (N_1235,N_669,N_31);
and U1236 (N_1236,N_7,N_612);
and U1237 (N_1237,N_277,N_941);
or U1238 (N_1238,N_468,N_879);
nor U1239 (N_1239,N_987,N_917);
nor U1240 (N_1240,N_823,N_17);
and U1241 (N_1241,N_451,N_280);
and U1242 (N_1242,N_443,N_349);
nor U1243 (N_1243,N_648,N_273);
nand U1244 (N_1244,N_546,N_854);
and U1245 (N_1245,N_87,N_67);
nor U1246 (N_1246,N_362,N_135);
nor U1247 (N_1247,N_105,N_114);
or U1248 (N_1248,N_930,N_548);
nor U1249 (N_1249,N_587,N_902);
nor U1250 (N_1250,N_824,N_509);
and U1251 (N_1251,N_262,N_175);
nor U1252 (N_1252,N_444,N_939);
nand U1253 (N_1253,N_161,N_598);
nand U1254 (N_1254,N_359,N_298);
nand U1255 (N_1255,N_351,N_532);
or U1256 (N_1256,N_403,N_168);
nand U1257 (N_1257,N_155,N_393);
nor U1258 (N_1258,N_916,N_284);
or U1259 (N_1259,N_447,N_383);
nand U1260 (N_1260,N_688,N_16);
nor U1261 (N_1261,N_321,N_197);
and U1262 (N_1262,N_700,N_492);
and U1263 (N_1263,N_881,N_223);
xnor U1264 (N_1264,N_866,N_3);
and U1265 (N_1265,N_339,N_478);
and U1266 (N_1266,N_654,N_788);
nand U1267 (N_1267,N_127,N_267);
nand U1268 (N_1268,N_377,N_777);
nand U1269 (N_1269,N_41,N_491);
and U1270 (N_1270,N_996,N_732);
and U1271 (N_1271,N_812,N_729);
or U1272 (N_1272,N_13,N_554);
or U1273 (N_1273,N_907,N_810);
or U1274 (N_1274,N_784,N_176);
and U1275 (N_1275,N_375,N_822);
nand U1276 (N_1276,N_869,N_620);
xnor U1277 (N_1277,N_611,N_682);
and U1278 (N_1278,N_34,N_708);
and U1279 (N_1279,N_360,N_501);
and U1280 (N_1280,N_245,N_370);
nand U1281 (N_1281,N_425,N_762);
nor U1282 (N_1282,N_979,N_358);
nand U1283 (N_1283,N_23,N_153);
nor U1284 (N_1284,N_367,N_214);
and U1285 (N_1285,N_722,N_678);
nand U1286 (N_1286,N_315,N_832);
nand U1287 (N_1287,N_307,N_900);
or U1288 (N_1288,N_691,N_962);
or U1289 (N_1289,N_805,N_776);
or U1290 (N_1290,N_552,N_898);
or U1291 (N_1291,N_927,N_906);
nor U1292 (N_1292,N_61,N_159);
or U1293 (N_1293,N_872,N_118);
and U1294 (N_1294,N_549,N_577);
and U1295 (N_1295,N_825,N_789);
nand U1296 (N_1296,N_45,N_870);
nand U1297 (N_1297,N_525,N_396);
nor U1298 (N_1298,N_850,N_773);
or U1299 (N_1299,N_976,N_346);
nor U1300 (N_1300,N_158,N_526);
nand U1301 (N_1301,N_98,N_513);
and U1302 (N_1302,N_160,N_85);
or U1303 (N_1303,N_616,N_73);
or U1304 (N_1304,N_856,N_865);
and U1305 (N_1305,N_126,N_911);
and U1306 (N_1306,N_920,N_575);
nor U1307 (N_1307,N_852,N_489);
or U1308 (N_1308,N_922,N_324);
nand U1309 (N_1309,N_399,N_474);
nand U1310 (N_1310,N_488,N_141);
or U1311 (N_1311,N_186,N_965);
and U1312 (N_1312,N_469,N_935);
or U1313 (N_1313,N_544,N_736);
or U1314 (N_1314,N_473,N_681);
nor U1315 (N_1315,N_457,N_143);
nor U1316 (N_1316,N_411,N_353);
and U1317 (N_1317,N_225,N_167);
nor U1318 (N_1318,N_551,N_452);
xnor U1319 (N_1319,N_95,N_634);
and U1320 (N_1320,N_641,N_261);
and U1321 (N_1321,N_769,N_565);
nor U1322 (N_1322,N_559,N_590);
and U1323 (N_1323,N_54,N_357);
xor U1324 (N_1324,N_229,N_236);
nor U1325 (N_1325,N_885,N_227);
nor U1326 (N_1326,N_932,N_342);
or U1327 (N_1327,N_880,N_106);
nand U1328 (N_1328,N_251,N_459);
and U1329 (N_1329,N_679,N_542);
nor U1330 (N_1330,N_512,N_198);
nand U1331 (N_1331,N_886,N_12);
nand U1332 (N_1332,N_287,N_740);
nand U1333 (N_1333,N_582,N_208);
nor U1334 (N_1334,N_945,N_111);
nand U1335 (N_1335,N_988,N_19);
nand U1336 (N_1336,N_790,N_563);
or U1337 (N_1337,N_704,N_379);
nor U1338 (N_1338,N_969,N_857);
nor U1339 (N_1339,N_128,N_402);
nor U1340 (N_1340,N_506,N_958);
nand U1341 (N_1341,N_199,N_901);
nor U1342 (N_1342,N_892,N_764);
nor U1343 (N_1343,N_642,N_44);
or U1344 (N_1344,N_65,N_181);
nor U1345 (N_1345,N_816,N_408);
nor U1346 (N_1346,N_68,N_519);
nand U1347 (N_1347,N_83,N_385);
and U1348 (N_1348,N_993,N_196);
or U1349 (N_1349,N_378,N_187);
and U1350 (N_1350,N_883,N_192);
nor U1351 (N_1351,N_814,N_431);
and U1352 (N_1352,N_657,N_139);
nor U1353 (N_1353,N_96,N_796);
nor U1354 (N_1354,N_465,N_449);
nand U1355 (N_1355,N_441,N_238);
or U1356 (N_1356,N_456,N_701);
and U1357 (N_1357,N_929,N_759);
and U1358 (N_1358,N_709,N_304);
or U1359 (N_1359,N_723,N_516);
and U1360 (N_1360,N_933,N_741);
and U1361 (N_1361,N_341,N_780);
nor U1362 (N_1362,N_687,N_966);
and U1363 (N_1363,N_655,N_576);
xnor U1364 (N_1364,N_32,N_619);
nand U1365 (N_1365,N_232,N_545);
nor U1366 (N_1366,N_115,N_103);
nand U1367 (N_1367,N_420,N_829);
and U1368 (N_1368,N_206,N_0);
nand U1369 (N_1369,N_666,N_82);
nand U1370 (N_1370,N_894,N_90);
and U1371 (N_1371,N_350,N_998);
or U1372 (N_1372,N_252,N_384);
nand U1373 (N_1373,N_953,N_650);
and U1374 (N_1374,N_47,N_464);
nand U1375 (N_1375,N_427,N_129);
nand U1376 (N_1376,N_335,N_815);
nand U1377 (N_1377,N_656,N_871);
nor U1378 (N_1378,N_42,N_81);
xor U1379 (N_1379,N_180,N_138);
nor U1380 (N_1380,N_354,N_826);
nor U1381 (N_1381,N_821,N_716);
nand U1382 (N_1382,N_801,N_567);
or U1383 (N_1383,N_278,N_364);
and U1384 (N_1384,N_25,N_483);
or U1385 (N_1385,N_835,N_40);
and U1386 (N_1386,N_588,N_243);
or U1387 (N_1387,N_309,N_553);
nor U1388 (N_1388,N_806,N_157);
or U1389 (N_1389,N_419,N_8);
or U1390 (N_1390,N_58,N_791);
nand U1391 (N_1391,N_975,N_728);
nand U1392 (N_1392,N_145,N_296);
nor U1393 (N_1393,N_733,N_614);
or U1394 (N_1394,N_391,N_325);
or U1395 (N_1395,N_761,N_212);
and U1396 (N_1396,N_983,N_301);
or U1397 (N_1397,N_905,N_585);
and U1398 (N_1398,N_466,N_799);
nor U1399 (N_1399,N_748,N_46);
or U1400 (N_1400,N_218,N_343);
nor U1401 (N_1401,N_795,N_78);
or U1402 (N_1402,N_171,N_904);
nand U1403 (N_1403,N_528,N_395);
nor U1404 (N_1404,N_878,N_537);
nand U1405 (N_1405,N_422,N_258);
nor U1406 (N_1406,N_680,N_599);
or U1407 (N_1407,N_797,N_6);
nand U1408 (N_1408,N_60,N_107);
nor U1409 (N_1409,N_194,N_786);
nor U1410 (N_1410,N_949,N_819);
nand U1411 (N_1411,N_984,N_990);
nand U1412 (N_1412,N_247,N_394);
nand U1413 (N_1413,N_131,N_595);
nor U1414 (N_1414,N_875,N_960);
nand U1415 (N_1415,N_416,N_578);
nand U1416 (N_1416,N_289,N_847);
and U1417 (N_1417,N_291,N_345);
and U1418 (N_1418,N_840,N_204);
nor U1419 (N_1419,N_951,N_182);
or U1420 (N_1420,N_237,N_310);
or U1421 (N_1421,N_281,N_30);
and U1422 (N_1422,N_803,N_744);
nor U1423 (N_1423,N_942,N_844);
and U1424 (N_1424,N_205,N_504);
or U1425 (N_1425,N_989,N_356);
and U1426 (N_1426,N_191,N_836);
nor U1427 (N_1427,N_144,N_592);
nor U1428 (N_1428,N_608,N_637);
or U1429 (N_1429,N_303,N_895);
nand U1430 (N_1430,N_259,N_527);
or U1431 (N_1431,N_147,N_74);
nand U1432 (N_1432,N_352,N_361);
or U1433 (N_1433,N_752,N_257);
and U1434 (N_1434,N_876,N_725);
nand U1435 (N_1435,N_601,N_1);
or U1436 (N_1436,N_49,N_476);
nand U1437 (N_1437,N_999,N_317);
nor U1438 (N_1438,N_531,N_583);
nand U1439 (N_1439,N_609,N_255);
and U1440 (N_1440,N_843,N_640);
nor U1441 (N_1441,N_433,N_381);
nor U1442 (N_1442,N_540,N_151);
nand U1443 (N_1443,N_288,N_771);
and U1444 (N_1444,N_808,N_200);
and U1445 (N_1445,N_926,N_610);
nor U1446 (N_1446,N_458,N_827);
nor U1447 (N_1447,N_858,N_482);
or U1448 (N_1448,N_365,N_48);
nor U1449 (N_1449,N_470,N_683);
or U1450 (N_1450,N_889,N_133);
nand U1451 (N_1451,N_241,N_652);
and U1452 (N_1452,N_644,N_494);
nor U1453 (N_1453,N_511,N_828);
nor U1454 (N_1454,N_673,N_368);
nand U1455 (N_1455,N_517,N_521);
nor U1456 (N_1456,N_742,N_888);
and U1457 (N_1457,N_479,N_775);
nand U1458 (N_1458,N_758,N_811);
and U1459 (N_1459,N_568,N_667);
nand U1460 (N_1460,N_116,N_507);
or U1461 (N_1461,N_747,N_994);
nand U1462 (N_1462,N_348,N_746);
nor U1463 (N_1463,N_500,N_401);
or U1464 (N_1464,N_952,N_692);
nor U1465 (N_1465,N_968,N_754);
or U1466 (N_1466,N_438,N_600);
nand U1467 (N_1467,N_946,N_77);
nand U1468 (N_1468,N_72,N_410);
nor U1469 (N_1469,N_671,N_120);
nand U1470 (N_1470,N_434,N_185);
nand U1471 (N_1471,N_738,N_340);
and U1472 (N_1472,N_662,N_646);
and U1473 (N_1473,N_407,N_613);
and U1474 (N_1474,N_830,N_130);
nor U1475 (N_1475,N_75,N_371);
and U1476 (N_1476,N_765,N_848);
nor U1477 (N_1477,N_573,N_868);
and U1478 (N_1478,N_580,N_271);
nor U1479 (N_1479,N_413,N_134);
nor U1480 (N_1480,N_409,N_121);
nor U1481 (N_1481,N_750,N_913);
nor U1482 (N_1482,N_623,N_779);
nand U1483 (N_1483,N_11,N_415);
nand U1484 (N_1484,N_442,N_914);
nand U1485 (N_1485,N_283,N_495);
nor U1486 (N_1486,N_436,N_428);
and U1487 (N_1487,N_97,N_472);
nand U1488 (N_1488,N_330,N_581);
nand U1489 (N_1489,N_912,N_5);
nand U1490 (N_1490,N_274,N_119);
and U1491 (N_1491,N_28,N_647);
nor U1492 (N_1492,N_27,N_974);
and U1493 (N_1493,N_295,N_372);
or U1494 (N_1494,N_179,N_873);
xnor U1495 (N_1495,N_593,N_248);
and U1496 (N_1496,N_417,N_730);
or U1497 (N_1497,N_336,N_499);
xor U1498 (N_1498,N_940,N_386);
nor U1499 (N_1499,N_757,N_448);
and U1500 (N_1500,N_949,N_445);
nand U1501 (N_1501,N_322,N_216);
and U1502 (N_1502,N_369,N_130);
nor U1503 (N_1503,N_983,N_774);
nor U1504 (N_1504,N_905,N_531);
nor U1505 (N_1505,N_751,N_999);
nor U1506 (N_1506,N_500,N_780);
nor U1507 (N_1507,N_557,N_836);
nand U1508 (N_1508,N_447,N_985);
nand U1509 (N_1509,N_233,N_37);
or U1510 (N_1510,N_264,N_119);
or U1511 (N_1511,N_731,N_733);
or U1512 (N_1512,N_285,N_37);
xnor U1513 (N_1513,N_147,N_901);
or U1514 (N_1514,N_992,N_826);
xnor U1515 (N_1515,N_181,N_866);
nor U1516 (N_1516,N_823,N_222);
nor U1517 (N_1517,N_776,N_10);
and U1518 (N_1518,N_58,N_713);
nor U1519 (N_1519,N_441,N_957);
and U1520 (N_1520,N_418,N_253);
or U1521 (N_1521,N_154,N_731);
nor U1522 (N_1522,N_537,N_296);
nand U1523 (N_1523,N_102,N_338);
nand U1524 (N_1524,N_315,N_841);
and U1525 (N_1525,N_524,N_767);
nor U1526 (N_1526,N_715,N_270);
nor U1527 (N_1527,N_41,N_314);
nor U1528 (N_1528,N_274,N_576);
nand U1529 (N_1529,N_25,N_848);
nor U1530 (N_1530,N_466,N_982);
nand U1531 (N_1531,N_123,N_514);
nand U1532 (N_1532,N_34,N_0);
nor U1533 (N_1533,N_758,N_72);
nand U1534 (N_1534,N_271,N_909);
or U1535 (N_1535,N_169,N_385);
nand U1536 (N_1536,N_490,N_953);
and U1537 (N_1537,N_825,N_673);
and U1538 (N_1538,N_936,N_611);
and U1539 (N_1539,N_294,N_949);
or U1540 (N_1540,N_758,N_55);
or U1541 (N_1541,N_979,N_549);
nor U1542 (N_1542,N_219,N_137);
or U1543 (N_1543,N_106,N_2);
and U1544 (N_1544,N_156,N_684);
and U1545 (N_1545,N_27,N_350);
and U1546 (N_1546,N_620,N_341);
or U1547 (N_1547,N_404,N_866);
or U1548 (N_1548,N_727,N_96);
nor U1549 (N_1549,N_488,N_611);
nand U1550 (N_1550,N_756,N_86);
and U1551 (N_1551,N_619,N_842);
nand U1552 (N_1552,N_554,N_459);
nand U1553 (N_1553,N_779,N_255);
and U1554 (N_1554,N_193,N_359);
or U1555 (N_1555,N_392,N_909);
and U1556 (N_1556,N_893,N_246);
and U1557 (N_1557,N_874,N_102);
nand U1558 (N_1558,N_834,N_116);
and U1559 (N_1559,N_735,N_524);
nand U1560 (N_1560,N_201,N_150);
and U1561 (N_1561,N_841,N_298);
nand U1562 (N_1562,N_377,N_803);
and U1563 (N_1563,N_92,N_793);
nand U1564 (N_1564,N_75,N_995);
or U1565 (N_1565,N_378,N_898);
nand U1566 (N_1566,N_361,N_614);
or U1567 (N_1567,N_876,N_742);
nor U1568 (N_1568,N_448,N_9);
nor U1569 (N_1569,N_663,N_436);
or U1570 (N_1570,N_159,N_989);
or U1571 (N_1571,N_572,N_220);
or U1572 (N_1572,N_32,N_162);
nor U1573 (N_1573,N_445,N_677);
nand U1574 (N_1574,N_344,N_996);
nor U1575 (N_1575,N_974,N_172);
nor U1576 (N_1576,N_871,N_246);
nor U1577 (N_1577,N_276,N_25);
nand U1578 (N_1578,N_260,N_309);
nor U1579 (N_1579,N_471,N_537);
nand U1580 (N_1580,N_761,N_683);
nor U1581 (N_1581,N_405,N_960);
and U1582 (N_1582,N_128,N_975);
nand U1583 (N_1583,N_302,N_990);
nor U1584 (N_1584,N_601,N_907);
or U1585 (N_1585,N_107,N_858);
nand U1586 (N_1586,N_832,N_859);
nor U1587 (N_1587,N_769,N_461);
nand U1588 (N_1588,N_613,N_807);
nand U1589 (N_1589,N_467,N_35);
and U1590 (N_1590,N_714,N_888);
and U1591 (N_1591,N_473,N_894);
and U1592 (N_1592,N_525,N_792);
or U1593 (N_1593,N_206,N_495);
or U1594 (N_1594,N_821,N_397);
nor U1595 (N_1595,N_207,N_57);
and U1596 (N_1596,N_321,N_758);
or U1597 (N_1597,N_870,N_361);
nor U1598 (N_1598,N_164,N_746);
and U1599 (N_1599,N_802,N_678);
nor U1600 (N_1600,N_356,N_479);
nand U1601 (N_1601,N_883,N_842);
and U1602 (N_1602,N_273,N_933);
or U1603 (N_1603,N_59,N_936);
nor U1604 (N_1604,N_46,N_205);
and U1605 (N_1605,N_626,N_971);
or U1606 (N_1606,N_108,N_314);
or U1607 (N_1607,N_495,N_603);
xnor U1608 (N_1608,N_592,N_380);
nand U1609 (N_1609,N_322,N_468);
nor U1610 (N_1610,N_678,N_438);
and U1611 (N_1611,N_794,N_570);
nand U1612 (N_1612,N_751,N_615);
nor U1613 (N_1613,N_741,N_632);
nand U1614 (N_1614,N_517,N_323);
and U1615 (N_1615,N_208,N_108);
or U1616 (N_1616,N_803,N_231);
nor U1617 (N_1617,N_791,N_191);
nand U1618 (N_1618,N_926,N_857);
nand U1619 (N_1619,N_798,N_814);
nand U1620 (N_1620,N_932,N_766);
or U1621 (N_1621,N_129,N_551);
or U1622 (N_1622,N_301,N_683);
and U1623 (N_1623,N_882,N_393);
nand U1624 (N_1624,N_808,N_238);
or U1625 (N_1625,N_754,N_912);
and U1626 (N_1626,N_83,N_785);
nand U1627 (N_1627,N_458,N_610);
and U1628 (N_1628,N_895,N_143);
or U1629 (N_1629,N_967,N_358);
and U1630 (N_1630,N_166,N_923);
nand U1631 (N_1631,N_394,N_799);
or U1632 (N_1632,N_128,N_644);
xnor U1633 (N_1633,N_739,N_109);
or U1634 (N_1634,N_751,N_705);
or U1635 (N_1635,N_760,N_448);
nor U1636 (N_1636,N_998,N_279);
and U1637 (N_1637,N_11,N_373);
nand U1638 (N_1638,N_802,N_482);
xor U1639 (N_1639,N_969,N_195);
nor U1640 (N_1640,N_54,N_245);
nand U1641 (N_1641,N_146,N_263);
and U1642 (N_1642,N_936,N_344);
nand U1643 (N_1643,N_313,N_513);
nand U1644 (N_1644,N_781,N_957);
nor U1645 (N_1645,N_234,N_656);
nand U1646 (N_1646,N_847,N_907);
or U1647 (N_1647,N_940,N_306);
nand U1648 (N_1648,N_10,N_278);
nor U1649 (N_1649,N_208,N_295);
and U1650 (N_1650,N_239,N_414);
and U1651 (N_1651,N_650,N_97);
xnor U1652 (N_1652,N_112,N_234);
or U1653 (N_1653,N_451,N_458);
and U1654 (N_1654,N_66,N_315);
and U1655 (N_1655,N_506,N_624);
nor U1656 (N_1656,N_854,N_474);
nand U1657 (N_1657,N_781,N_558);
or U1658 (N_1658,N_483,N_493);
or U1659 (N_1659,N_918,N_183);
nor U1660 (N_1660,N_871,N_592);
and U1661 (N_1661,N_974,N_797);
or U1662 (N_1662,N_778,N_730);
and U1663 (N_1663,N_71,N_354);
nand U1664 (N_1664,N_416,N_604);
and U1665 (N_1665,N_402,N_298);
and U1666 (N_1666,N_769,N_661);
nor U1667 (N_1667,N_391,N_168);
nand U1668 (N_1668,N_235,N_37);
xor U1669 (N_1669,N_967,N_686);
nor U1670 (N_1670,N_608,N_354);
nor U1671 (N_1671,N_788,N_325);
nand U1672 (N_1672,N_346,N_506);
nor U1673 (N_1673,N_416,N_654);
and U1674 (N_1674,N_377,N_792);
nand U1675 (N_1675,N_980,N_271);
or U1676 (N_1676,N_456,N_193);
nand U1677 (N_1677,N_127,N_340);
or U1678 (N_1678,N_412,N_529);
or U1679 (N_1679,N_384,N_616);
nand U1680 (N_1680,N_50,N_360);
and U1681 (N_1681,N_275,N_490);
or U1682 (N_1682,N_426,N_760);
and U1683 (N_1683,N_141,N_55);
or U1684 (N_1684,N_649,N_640);
nand U1685 (N_1685,N_198,N_104);
and U1686 (N_1686,N_800,N_60);
nand U1687 (N_1687,N_361,N_669);
or U1688 (N_1688,N_703,N_467);
and U1689 (N_1689,N_253,N_596);
nand U1690 (N_1690,N_126,N_4);
and U1691 (N_1691,N_123,N_71);
nor U1692 (N_1692,N_564,N_324);
nor U1693 (N_1693,N_714,N_391);
nand U1694 (N_1694,N_705,N_110);
nand U1695 (N_1695,N_123,N_853);
or U1696 (N_1696,N_460,N_784);
and U1697 (N_1697,N_619,N_938);
and U1698 (N_1698,N_633,N_762);
nand U1699 (N_1699,N_787,N_749);
or U1700 (N_1700,N_941,N_364);
nor U1701 (N_1701,N_947,N_56);
nand U1702 (N_1702,N_190,N_304);
nor U1703 (N_1703,N_708,N_112);
and U1704 (N_1704,N_125,N_186);
nand U1705 (N_1705,N_411,N_750);
and U1706 (N_1706,N_33,N_555);
nor U1707 (N_1707,N_355,N_516);
nor U1708 (N_1708,N_545,N_988);
nand U1709 (N_1709,N_941,N_102);
nor U1710 (N_1710,N_636,N_507);
and U1711 (N_1711,N_640,N_967);
and U1712 (N_1712,N_12,N_748);
or U1713 (N_1713,N_884,N_697);
and U1714 (N_1714,N_191,N_691);
and U1715 (N_1715,N_394,N_207);
nor U1716 (N_1716,N_222,N_6);
nor U1717 (N_1717,N_476,N_669);
or U1718 (N_1718,N_707,N_434);
nand U1719 (N_1719,N_901,N_368);
and U1720 (N_1720,N_410,N_170);
nand U1721 (N_1721,N_279,N_976);
or U1722 (N_1722,N_234,N_834);
or U1723 (N_1723,N_238,N_613);
nor U1724 (N_1724,N_833,N_372);
xnor U1725 (N_1725,N_89,N_342);
nand U1726 (N_1726,N_524,N_784);
or U1727 (N_1727,N_841,N_168);
and U1728 (N_1728,N_552,N_342);
or U1729 (N_1729,N_712,N_695);
nor U1730 (N_1730,N_855,N_837);
nor U1731 (N_1731,N_207,N_159);
nor U1732 (N_1732,N_776,N_896);
nor U1733 (N_1733,N_914,N_712);
nand U1734 (N_1734,N_979,N_657);
nor U1735 (N_1735,N_121,N_753);
nand U1736 (N_1736,N_712,N_164);
nor U1737 (N_1737,N_209,N_952);
and U1738 (N_1738,N_429,N_539);
nor U1739 (N_1739,N_157,N_798);
nand U1740 (N_1740,N_649,N_245);
nor U1741 (N_1741,N_90,N_684);
nor U1742 (N_1742,N_379,N_137);
nor U1743 (N_1743,N_642,N_255);
nand U1744 (N_1744,N_740,N_316);
or U1745 (N_1745,N_536,N_884);
and U1746 (N_1746,N_610,N_298);
or U1747 (N_1747,N_8,N_224);
nor U1748 (N_1748,N_691,N_497);
or U1749 (N_1749,N_419,N_496);
or U1750 (N_1750,N_191,N_250);
or U1751 (N_1751,N_536,N_472);
nand U1752 (N_1752,N_64,N_693);
nand U1753 (N_1753,N_891,N_393);
and U1754 (N_1754,N_760,N_456);
nor U1755 (N_1755,N_105,N_107);
or U1756 (N_1756,N_460,N_581);
nor U1757 (N_1757,N_891,N_285);
nand U1758 (N_1758,N_207,N_220);
or U1759 (N_1759,N_847,N_955);
nor U1760 (N_1760,N_515,N_28);
or U1761 (N_1761,N_219,N_22);
nand U1762 (N_1762,N_951,N_575);
nand U1763 (N_1763,N_966,N_404);
or U1764 (N_1764,N_85,N_122);
and U1765 (N_1765,N_807,N_443);
nor U1766 (N_1766,N_860,N_569);
nor U1767 (N_1767,N_872,N_110);
nand U1768 (N_1768,N_476,N_727);
nor U1769 (N_1769,N_357,N_398);
nand U1770 (N_1770,N_405,N_527);
or U1771 (N_1771,N_596,N_517);
nand U1772 (N_1772,N_867,N_624);
or U1773 (N_1773,N_865,N_693);
and U1774 (N_1774,N_288,N_793);
nor U1775 (N_1775,N_969,N_21);
nor U1776 (N_1776,N_101,N_441);
nor U1777 (N_1777,N_614,N_726);
nand U1778 (N_1778,N_122,N_292);
nor U1779 (N_1779,N_686,N_295);
nand U1780 (N_1780,N_176,N_439);
nor U1781 (N_1781,N_193,N_845);
or U1782 (N_1782,N_722,N_395);
nor U1783 (N_1783,N_993,N_911);
nand U1784 (N_1784,N_859,N_592);
nand U1785 (N_1785,N_583,N_516);
or U1786 (N_1786,N_462,N_621);
nand U1787 (N_1787,N_454,N_519);
or U1788 (N_1788,N_745,N_102);
and U1789 (N_1789,N_571,N_871);
nor U1790 (N_1790,N_506,N_447);
nand U1791 (N_1791,N_838,N_909);
nand U1792 (N_1792,N_466,N_680);
xor U1793 (N_1793,N_59,N_171);
nand U1794 (N_1794,N_885,N_925);
or U1795 (N_1795,N_914,N_918);
and U1796 (N_1796,N_970,N_677);
or U1797 (N_1797,N_870,N_830);
or U1798 (N_1798,N_210,N_49);
or U1799 (N_1799,N_929,N_977);
nor U1800 (N_1800,N_324,N_688);
xor U1801 (N_1801,N_498,N_891);
nor U1802 (N_1802,N_393,N_860);
and U1803 (N_1803,N_610,N_222);
and U1804 (N_1804,N_437,N_572);
or U1805 (N_1805,N_684,N_636);
and U1806 (N_1806,N_385,N_723);
xnor U1807 (N_1807,N_766,N_188);
or U1808 (N_1808,N_93,N_893);
and U1809 (N_1809,N_929,N_731);
nor U1810 (N_1810,N_596,N_890);
nand U1811 (N_1811,N_154,N_821);
nor U1812 (N_1812,N_549,N_509);
or U1813 (N_1813,N_712,N_924);
nand U1814 (N_1814,N_533,N_826);
or U1815 (N_1815,N_560,N_863);
nand U1816 (N_1816,N_418,N_4);
or U1817 (N_1817,N_95,N_231);
nand U1818 (N_1818,N_553,N_92);
xnor U1819 (N_1819,N_890,N_414);
or U1820 (N_1820,N_150,N_695);
or U1821 (N_1821,N_978,N_362);
and U1822 (N_1822,N_998,N_779);
nand U1823 (N_1823,N_431,N_227);
nand U1824 (N_1824,N_342,N_67);
or U1825 (N_1825,N_235,N_204);
nor U1826 (N_1826,N_252,N_623);
or U1827 (N_1827,N_622,N_350);
or U1828 (N_1828,N_672,N_569);
and U1829 (N_1829,N_866,N_325);
nand U1830 (N_1830,N_120,N_438);
xnor U1831 (N_1831,N_971,N_994);
or U1832 (N_1832,N_316,N_942);
and U1833 (N_1833,N_867,N_584);
nor U1834 (N_1834,N_981,N_879);
or U1835 (N_1835,N_572,N_856);
nand U1836 (N_1836,N_344,N_27);
or U1837 (N_1837,N_189,N_376);
and U1838 (N_1838,N_615,N_13);
or U1839 (N_1839,N_827,N_7);
nor U1840 (N_1840,N_349,N_398);
or U1841 (N_1841,N_899,N_935);
xnor U1842 (N_1842,N_318,N_865);
nand U1843 (N_1843,N_79,N_135);
or U1844 (N_1844,N_286,N_95);
nand U1845 (N_1845,N_160,N_748);
nand U1846 (N_1846,N_557,N_572);
nor U1847 (N_1847,N_942,N_902);
nand U1848 (N_1848,N_684,N_393);
or U1849 (N_1849,N_534,N_591);
and U1850 (N_1850,N_501,N_487);
nor U1851 (N_1851,N_765,N_48);
nand U1852 (N_1852,N_691,N_21);
nand U1853 (N_1853,N_840,N_620);
nand U1854 (N_1854,N_368,N_151);
and U1855 (N_1855,N_387,N_711);
nor U1856 (N_1856,N_948,N_294);
nand U1857 (N_1857,N_931,N_693);
or U1858 (N_1858,N_497,N_212);
or U1859 (N_1859,N_485,N_639);
or U1860 (N_1860,N_492,N_516);
nor U1861 (N_1861,N_43,N_906);
nor U1862 (N_1862,N_194,N_678);
and U1863 (N_1863,N_740,N_175);
or U1864 (N_1864,N_330,N_332);
and U1865 (N_1865,N_600,N_349);
nand U1866 (N_1866,N_899,N_27);
xor U1867 (N_1867,N_635,N_706);
nand U1868 (N_1868,N_575,N_684);
or U1869 (N_1869,N_983,N_636);
nor U1870 (N_1870,N_569,N_628);
nor U1871 (N_1871,N_770,N_716);
and U1872 (N_1872,N_770,N_56);
and U1873 (N_1873,N_752,N_459);
or U1874 (N_1874,N_203,N_238);
or U1875 (N_1875,N_111,N_20);
or U1876 (N_1876,N_245,N_929);
nor U1877 (N_1877,N_937,N_808);
or U1878 (N_1878,N_179,N_988);
nor U1879 (N_1879,N_101,N_424);
nor U1880 (N_1880,N_200,N_859);
nand U1881 (N_1881,N_861,N_541);
nor U1882 (N_1882,N_715,N_541);
nand U1883 (N_1883,N_510,N_366);
nand U1884 (N_1884,N_282,N_937);
nor U1885 (N_1885,N_980,N_77);
or U1886 (N_1886,N_618,N_928);
or U1887 (N_1887,N_33,N_185);
or U1888 (N_1888,N_63,N_847);
or U1889 (N_1889,N_761,N_503);
nor U1890 (N_1890,N_355,N_741);
or U1891 (N_1891,N_20,N_952);
or U1892 (N_1892,N_544,N_957);
and U1893 (N_1893,N_212,N_879);
nor U1894 (N_1894,N_852,N_234);
nor U1895 (N_1895,N_431,N_920);
nand U1896 (N_1896,N_309,N_430);
and U1897 (N_1897,N_195,N_933);
or U1898 (N_1898,N_430,N_336);
and U1899 (N_1899,N_134,N_816);
xor U1900 (N_1900,N_639,N_681);
nor U1901 (N_1901,N_985,N_943);
and U1902 (N_1902,N_177,N_148);
and U1903 (N_1903,N_832,N_766);
and U1904 (N_1904,N_633,N_829);
nor U1905 (N_1905,N_878,N_56);
nor U1906 (N_1906,N_106,N_23);
and U1907 (N_1907,N_201,N_774);
nor U1908 (N_1908,N_195,N_616);
and U1909 (N_1909,N_990,N_898);
nand U1910 (N_1910,N_763,N_901);
or U1911 (N_1911,N_244,N_574);
or U1912 (N_1912,N_160,N_661);
nor U1913 (N_1913,N_786,N_971);
or U1914 (N_1914,N_169,N_442);
nor U1915 (N_1915,N_854,N_446);
or U1916 (N_1916,N_448,N_870);
or U1917 (N_1917,N_617,N_329);
and U1918 (N_1918,N_174,N_267);
nand U1919 (N_1919,N_18,N_237);
or U1920 (N_1920,N_992,N_815);
and U1921 (N_1921,N_922,N_165);
nand U1922 (N_1922,N_292,N_910);
and U1923 (N_1923,N_359,N_21);
or U1924 (N_1924,N_196,N_490);
nor U1925 (N_1925,N_904,N_788);
and U1926 (N_1926,N_495,N_624);
or U1927 (N_1927,N_505,N_968);
nor U1928 (N_1928,N_37,N_107);
nand U1929 (N_1929,N_291,N_993);
or U1930 (N_1930,N_979,N_484);
nand U1931 (N_1931,N_295,N_991);
nor U1932 (N_1932,N_878,N_922);
and U1933 (N_1933,N_4,N_978);
nor U1934 (N_1934,N_625,N_668);
or U1935 (N_1935,N_121,N_177);
xnor U1936 (N_1936,N_72,N_218);
and U1937 (N_1937,N_634,N_363);
nand U1938 (N_1938,N_303,N_746);
nor U1939 (N_1939,N_508,N_411);
nor U1940 (N_1940,N_586,N_240);
and U1941 (N_1941,N_963,N_858);
xor U1942 (N_1942,N_829,N_765);
and U1943 (N_1943,N_372,N_639);
nand U1944 (N_1944,N_557,N_20);
nand U1945 (N_1945,N_766,N_390);
or U1946 (N_1946,N_673,N_335);
xor U1947 (N_1947,N_558,N_353);
nor U1948 (N_1948,N_937,N_591);
nor U1949 (N_1949,N_618,N_943);
or U1950 (N_1950,N_656,N_13);
and U1951 (N_1951,N_219,N_159);
or U1952 (N_1952,N_96,N_359);
nor U1953 (N_1953,N_260,N_972);
and U1954 (N_1954,N_941,N_772);
nor U1955 (N_1955,N_317,N_402);
or U1956 (N_1956,N_101,N_683);
or U1957 (N_1957,N_408,N_275);
nor U1958 (N_1958,N_288,N_986);
nand U1959 (N_1959,N_164,N_954);
nand U1960 (N_1960,N_990,N_380);
nor U1961 (N_1961,N_863,N_86);
nand U1962 (N_1962,N_914,N_520);
or U1963 (N_1963,N_983,N_257);
or U1964 (N_1964,N_400,N_6);
nand U1965 (N_1965,N_59,N_458);
nor U1966 (N_1966,N_637,N_309);
and U1967 (N_1967,N_690,N_276);
or U1968 (N_1968,N_970,N_370);
and U1969 (N_1969,N_414,N_323);
or U1970 (N_1970,N_967,N_485);
nor U1971 (N_1971,N_204,N_446);
xnor U1972 (N_1972,N_349,N_70);
xor U1973 (N_1973,N_633,N_129);
or U1974 (N_1974,N_538,N_89);
and U1975 (N_1975,N_572,N_650);
nand U1976 (N_1976,N_286,N_292);
nand U1977 (N_1977,N_716,N_371);
or U1978 (N_1978,N_693,N_446);
and U1979 (N_1979,N_977,N_828);
nand U1980 (N_1980,N_514,N_669);
nand U1981 (N_1981,N_215,N_352);
or U1982 (N_1982,N_156,N_543);
and U1983 (N_1983,N_959,N_441);
nand U1984 (N_1984,N_910,N_693);
and U1985 (N_1985,N_808,N_302);
or U1986 (N_1986,N_340,N_627);
nand U1987 (N_1987,N_33,N_706);
and U1988 (N_1988,N_799,N_118);
xor U1989 (N_1989,N_335,N_928);
or U1990 (N_1990,N_364,N_631);
nand U1991 (N_1991,N_103,N_404);
nand U1992 (N_1992,N_773,N_270);
nor U1993 (N_1993,N_818,N_938);
nand U1994 (N_1994,N_715,N_673);
nor U1995 (N_1995,N_660,N_547);
or U1996 (N_1996,N_850,N_957);
nor U1997 (N_1997,N_273,N_6);
and U1998 (N_1998,N_825,N_612);
nor U1999 (N_1999,N_720,N_715);
nor U2000 (N_2000,N_1356,N_1293);
or U2001 (N_2001,N_1942,N_1009);
nand U2002 (N_2002,N_1675,N_1700);
nor U2003 (N_2003,N_1708,N_1091);
nor U2004 (N_2004,N_1460,N_1059);
or U2005 (N_2005,N_1550,N_1053);
nor U2006 (N_2006,N_1449,N_1976);
nand U2007 (N_2007,N_1456,N_1487);
and U2008 (N_2008,N_1931,N_1027);
nor U2009 (N_2009,N_1219,N_1331);
and U2010 (N_2010,N_1162,N_1164);
and U2011 (N_2011,N_1485,N_1890);
and U2012 (N_2012,N_1187,N_1035);
and U2013 (N_2013,N_1384,N_1061);
nand U2014 (N_2014,N_1048,N_1596);
and U2015 (N_2015,N_1267,N_1787);
or U2016 (N_2016,N_1870,N_1818);
and U2017 (N_2017,N_1999,N_1711);
nor U2018 (N_2018,N_1945,N_1328);
and U2019 (N_2019,N_1809,N_1716);
nand U2020 (N_2020,N_1057,N_1691);
nor U2021 (N_2021,N_1914,N_1194);
nand U2022 (N_2022,N_1095,N_1515);
nand U2023 (N_2023,N_1011,N_1245);
nand U2024 (N_2024,N_1595,N_1520);
or U2025 (N_2025,N_1755,N_1078);
and U2026 (N_2026,N_1113,N_1569);
or U2027 (N_2027,N_1147,N_1758);
or U2028 (N_2028,N_1246,N_1026);
nor U2029 (N_2029,N_1768,N_1365);
nor U2030 (N_2030,N_1380,N_1020);
and U2031 (N_2031,N_1276,N_1070);
or U2032 (N_2032,N_1962,N_1547);
or U2033 (N_2033,N_1317,N_1014);
nor U2034 (N_2034,N_1626,N_1501);
nor U2035 (N_2035,N_1939,N_1851);
and U2036 (N_2036,N_1115,N_1021);
and U2037 (N_2037,N_1018,N_1660);
nand U2038 (N_2038,N_1629,N_1107);
and U2039 (N_2039,N_1714,N_1184);
and U2040 (N_2040,N_1412,N_1553);
or U2041 (N_2041,N_1154,N_1480);
or U2042 (N_2042,N_1320,N_1467);
nand U2043 (N_2043,N_1614,N_1774);
nand U2044 (N_2044,N_1438,N_1673);
and U2045 (N_2045,N_1453,N_1968);
or U2046 (N_2046,N_1486,N_1188);
and U2047 (N_2047,N_1579,N_1805);
and U2048 (N_2048,N_1208,N_1577);
or U2049 (N_2049,N_1712,N_1294);
nand U2050 (N_2050,N_1732,N_1340);
nand U2051 (N_2051,N_1559,N_1200);
nand U2052 (N_2052,N_1314,N_1977);
nor U2053 (N_2053,N_1685,N_1969);
nor U2054 (N_2054,N_1372,N_1475);
or U2055 (N_2055,N_1023,N_1257);
nor U2056 (N_2056,N_1802,N_1282);
nor U2057 (N_2057,N_1642,N_1135);
nor U2058 (N_2058,N_1876,N_1771);
and U2059 (N_2059,N_1672,N_1007);
or U2060 (N_2060,N_1610,N_1419);
and U2061 (N_2061,N_1721,N_1121);
or U2062 (N_2062,N_1473,N_1912);
nand U2063 (N_2063,N_1782,N_1592);
nand U2064 (N_2064,N_1959,N_1590);
or U2065 (N_2065,N_1929,N_1071);
nor U2066 (N_2066,N_1993,N_1639);
and U2067 (N_2067,N_1346,N_1854);
nand U2068 (N_2068,N_1288,N_1006);
or U2069 (N_2069,N_1043,N_1935);
nor U2070 (N_2070,N_1646,N_1278);
nor U2071 (N_2071,N_1253,N_1051);
nand U2072 (N_2072,N_1830,N_1069);
or U2073 (N_2073,N_1916,N_1047);
nor U2074 (N_2074,N_1989,N_1054);
nor U2075 (N_2075,N_1741,N_1540);
nor U2076 (N_2076,N_1795,N_1079);
and U2077 (N_2077,N_1676,N_1889);
nor U2078 (N_2078,N_1172,N_1546);
and U2079 (N_2079,N_1662,N_1322);
or U2080 (N_2080,N_1648,N_1155);
nand U2081 (N_2081,N_1376,N_1665);
or U2082 (N_2082,N_1954,N_1719);
nor U2083 (N_2083,N_1281,N_1955);
and U2084 (N_2084,N_1526,N_1283);
nand U2085 (N_2085,N_1607,N_1242);
and U2086 (N_2086,N_1858,N_1400);
and U2087 (N_2087,N_1883,N_1112);
or U2088 (N_2088,N_1213,N_1783);
and U2089 (N_2089,N_1826,N_1360);
and U2090 (N_2090,N_1171,N_1994);
nor U2091 (N_2091,N_1538,N_1810);
nand U2092 (N_2092,N_1867,N_1735);
nand U2093 (N_2093,N_1272,N_1630);
and U2094 (N_2094,N_1625,N_1581);
or U2095 (N_2095,N_1399,N_1508);
nor U2096 (N_2096,N_1899,N_1221);
and U2097 (N_2097,N_1841,N_1654);
nor U2098 (N_2098,N_1287,N_1562);
or U2099 (N_2099,N_1210,N_1106);
nor U2100 (N_2100,N_1203,N_1225);
nor U2101 (N_2101,N_1097,N_1045);
and U2102 (N_2102,N_1420,N_1313);
nand U2103 (N_2103,N_1726,N_1844);
and U2104 (N_2104,N_1584,N_1214);
nand U2105 (N_2105,N_1720,N_1872);
nor U2106 (N_2106,N_1146,N_1445);
nand U2107 (N_2107,N_1240,N_1885);
and U2108 (N_2108,N_1619,N_1457);
nor U2109 (N_2109,N_1689,N_1087);
and U2110 (N_2110,N_1759,N_1589);
nand U2111 (N_2111,N_1531,N_1522);
nand U2112 (N_2112,N_1388,N_1565);
nor U2113 (N_2113,N_1046,N_1695);
or U2114 (N_2114,N_1472,N_1754);
or U2115 (N_2115,N_1597,N_1973);
nand U2116 (N_2116,N_1049,N_1984);
and U2117 (N_2117,N_1866,N_1108);
and U2118 (N_2118,N_1205,N_1778);
and U2119 (N_2119,N_1183,N_1674);
or U2120 (N_2120,N_1650,N_1038);
nor U2121 (N_2121,N_1296,N_1692);
nor U2122 (N_2122,N_1568,N_1298);
or U2123 (N_2123,N_1111,N_1963);
nand U2124 (N_2124,N_1679,N_1443);
nor U2125 (N_2125,N_1943,N_1815);
nor U2126 (N_2126,N_1861,N_1848);
nor U2127 (N_2127,N_1458,N_1576);
or U2128 (N_2128,N_1825,N_1613);
nand U2129 (N_2129,N_1634,N_1258);
nand U2130 (N_2130,N_1000,N_1570);
and U2131 (N_2131,N_1284,N_1103);
and U2132 (N_2132,N_1279,N_1640);
nand U2133 (N_2133,N_1195,N_1292);
nand U2134 (N_2134,N_1838,N_1435);
nor U2135 (N_2135,N_1748,N_1381);
or U2136 (N_2136,N_1637,N_1093);
and U2137 (N_2137,N_1965,N_1554);
xor U2138 (N_2138,N_1996,N_1122);
or U2139 (N_2139,N_1667,N_1259);
and U2140 (N_2140,N_1131,N_1130);
nand U2141 (N_2141,N_1212,N_1713);
xnor U2142 (N_2142,N_1414,N_1418);
and U2143 (N_2143,N_1923,N_1436);
or U2144 (N_2144,N_1181,N_1940);
or U2145 (N_2145,N_1926,N_1133);
nor U2146 (N_2146,N_1289,N_1013);
or U2147 (N_2147,N_1505,N_1076);
or U2148 (N_2148,N_1316,N_1490);
nand U2149 (N_2149,N_1229,N_1652);
nand U2150 (N_2150,N_1509,N_1718);
and U2151 (N_2151,N_1392,N_1836);
nor U2152 (N_2152,N_1179,N_1439);
and U2153 (N_2153,N_1158,N_1028);
and U2154 (N_2154,N_1005,N_1189);
nor U2155 (N_2155,N_1469,N_1077);
and U2156 (N_2156,N_1752,N_1353);
and U2157 (N_2157,N_1792,N_1657);
and U2158 (N_2158,N_1333,N_1730);
nand U2159 (N_2159,N_1379,N_1961);
or U2160 (N_2160,N_1442,N_1539);
or U2161 (N_2161,N_1228,N_1015);
nand U2162 (N_2162,N_1575,N_1427);
nand U2163 (N_2163,N_1821,N_1390);
and U2164 (N_2164,N_1295,N_1285);
nand U2165 (N_2165,N_1177,N_1431);
or U2166 (N_2166,N_1717,N_1697);
and U2167 (N_2167,N_1850,N_1003);
nor U2168 (N_2168,N_1056,N_1555);
nor U2169 (N_2169,N_1124,N_1434);
nand U2170 (N_2170,N_1779,N_1823);
nor U2171 (N_2171,N_1928,N_1019);
and U2172 (N_2172,N_1297,N_1585);
xor U2173 (N_2173,N_1134,N_1081);
and U2174 (N_2174,N_1139,N_1303);
nor U2175 (N_2175,N_1724,N_1903);
xnor U2176 (N_2176,N_1886,N_1847);
nand U2177 (N_2177,N_1152,N_1970);
and U2178 (N_2178,N_1879,N_1310);
nand U2179 (N_2179,N_1141,N_1790);
nand U2180 (N_2180,N_1960,N_1643);
or U2181 (N_2181,N_1725,N_1966);
nand U2182 (N_2182,N_1033,N_1644);
or U2183 (N_2183,N_1710,N_1494);
and U2184 (N_2184,N_1729,N_1918);
and U2185 (N_2185,N_1857,N_1336);
nor U2186 (N_2186,N_1743,N_1041);
and U2187 (N_2187,N_1063,N_1558);
nand U2188 (N_2188,N_1483,N_1060);
nor U2189 (N_2189,N_1030,N_1136);
nand U2190 (N_2190,N_1196,N_1820);
and U2191 (N_2191,N_1512,N_1206);
or U2192 (N_2192,N_1271,N_1249);
and U2193 (N_2193,N_1243,N_1822);
nor U2194 (N_2194,N_1302,N_1341);
or U2195 (N_2195,N_1892,N_1776);
nor U2196 (N_2196,N_1801,N_1119);
or U2197 (N_2197,N_1173,N_1440);
or U2198 (N_2198,N_1426,N_1911);
nor U2199 (N_2199,N_1762,N_1266);
and U2200 (N_2200,N_1454,N_1393);
nand U2201 (N_2201,N_1819,N_1444);
or U2202 (N_2202,N_1425,N_1199);
nand U2203 (N_2203,N_1618,N_1044);
or U2204 (N_2204,N_1389,N_1615);
and U2205 (N_2205,N_1506,N_1153);
and U2206 (N_2206,N_1736,N_1017);
nand U2207 (N_2207,N_1764,N_1894);
or U2208 (N_2208,N_1367,N_1073);
nand U2209 (N_2209,N_1128,N_1739);
or U2210 (N_2210,N_1116,N_1941);
or U2211 (N_2211,N_1636,N_1991);
nor U2212 (N_2212,N_1319,N_1873);
and U2213 (N_2213,N_1471,N_1364);
and U2214 (N_2214,N_1268,N_1391);
nand U2215 (N_2215,N_1123,N_1495);
and U2216 (N_2216,N_1375,N_1734);
and U2217 (N_2217,N_1191,N_1798);
and U2218 (N_2218,N_1852,N_1747);
or U2219 (N_2219,N_1773,N_1525);
or U2220 (N_2220,N_1226,N_1120);
nor U2221 (N_2221,N_1042,N_1517);
nor U2222 (N_2222,N_1263,N_1148);
and U2223 (N_2223,N_1345,N_1036);
nand U2224 (N_2224,N_1410,N_1668);
nand U2225 (N_2225,N_1477,N_1080);
nor U2226 (N_2226,N_1706,N_1900);
nor U2227 (N_2227,N_1062,N_1990);
nand U2228 (N_2228,N_1432,N_1409);
nor U2229 (N_2229,N_1357,N_1447);
and U2230 (N_2230,N_1355,N_1658);
and U2231 (N_2231,N_1190,N_1016);
or U2232 (N_2232,N_1663,N_1533);
nor U2233 (N_2233,N_1324,N_1740);
xor U2234 (N_2234,N_1967,N_1757);
nand U2235 (N_2235,N_1745,N_1350);
or U2236 (N_2236,N_1863,N_1204);
nor U2237 (N_2237,N_1261,N_1702);
or U2238 (N_2238,N_1543,N_1144);
or U2239 (N_2239,N_1705,N_1549);
or U2240 (N_2240,N_1915,N_1157);
or U2241 (N_2241,N_1601,N_1193);
nand U2242 (N_2242,N_1829,N_1796);
and U2243 (N_2243,N_1544,N_1415);
nand U2244 (N_2244,N_1104,N_1982);
and U2245 (N_2245,N_1617,N_1402);
nand U2246 (N_2246,N_1680,N_1744);
or U2247 (N_2247,N_1012,N_1306);
or U2248 (N_2248,N_1898,N_1738);
nand U2249 (N_2249,N_1241,N_1881);
nor U2250 (N_2250,N_1766,N_1924);
nand U2251 (N_2251,N_1932,N_1140);
xor U2252 (N_2252,N_1653,N_1092);
xor U2253 (N_2253,N_1906,N_1305);
nor U2254 (N_2254,N_1383,N_1651);
nand U2255 (N_2255,N_1489,N_1156);
or U2256 (N_2256,N_1239,N_1039);
nand U2257 (N_2257,N_1430,N_1500);
and U2258 (N_2258,N_1574,N_1731);
nand U2259 (N_2259,N_1728,N_1269);
nor U2260 (N_2260,N_1358,N_1084);
and U2261 (N_2261,N_1611,N_1318);
nand U2262 (N_2262,N_1860,N_1519);
nand U2263 (N_2263,N_1169,N_1750);
nand U2264 (N_2264,N_1599,N_1274);
nand U2265 (N_2265,N_1834,N_1248);
and U2266 (N_2266,N_1799,N_1600);
or U2267 (N_2267,N_1608,N_1373);
nand U2268 (N_2268,N_1065,N_1224);
and U2269 (N_2269,N_1632,N_1416);
and U2270 (N_2270,N_1031,N_1493);
nand U2271 (N_2271,N_1952,N_1451);
xnor U2272 (N_2272,N_1405,N_1812);
and U2273 (N_2273,N_1234,N_1749);
nand U2274 (N_2274,N_1503,N_1270);
xnor U2275 (N_2275,N_1995,N_1704);
and U2276 (N_2276,N_1227,N_1609);
nand U2277 (N_2277,N_1201,N_1359);
nand U2278 (N_2278,N_1760,N_1507);
nor U2279 (N_2279,N_1542,N_1163);
or U2280 (N_2280,N_1623,N_1669);
and U2281 (N_2281,N_1315,N_1394);
nor U2282 (N_2282,N_1814,N_1192);
and U2283 (N_2283,N_1462,N_1265);
nand U2284 (N_2284,N_1050,N_1251);
or U2285 (N_2285,N_1448,N_1127);
nand U2286 (N_2286,N_1256,N_1304);
nand U2287 (N_2287,N_1536,N_1746);
or U2288 (N_2288,N_1987,N_1082);
nor U2289 (N_2289,N_1694,N_1450);
xnor U2290 (N_2290,N_1034,N_1602);
or U2291 (N_2291,N_1545,N_1429);
or U2292 (N_2292,N_1408,N_1833);
nand U2293 (N_2293,N_1105,N_1902);
and U2294 (N_2294,N_1645,N_1563);
and U2295 (N_2295,N_1344,N_1474);
and U2296 (N_2296,N_1789,N_1510);
and U2297 (N_2297,N_1933,N_1958);
nand U2298 (N_2298,N_1586,N_1803);
and U2299 (N_2299,N_1887,N_1780);
nand U2300 (N_2300,N_1465,N_1176);
nand U2301 (N_2301,N_1232,N_1572);
xnor U2302 (N_2302,N_1089,N_1484);
and U2303 (N_2303,N_1488,N_1185);
and U2304 (N_2304,N_1230,N_1482);
xor U2305 (N_2305,N_1403,N_1161);
or U2306 (N_2306,N_1529,N_1856);
xor U2307 (N_2307,N_1335,N_1594);
and U2308 (N_2308,N_1781,N_1004);
nand U2309 (N_2309,N_1511,N_1763);
or U2310 (N_2310,N_1964,N_1499);
nand U2311 (N_2311,N_1086,N_1291);
nor U2312 (N_2312,N_1580,N_1788);
nor U2313 (N_2313,N_1666,N_1875);
nand U2314 (N_2314,N_1913,N_1896);
or U2315 (N_2315,N_1514,N_1478);
nor U2316 (N_2316,N_1085,N_1715);
or U2317 (N_2317,N_1845,N_1138);
or U2318 (N_2318,N_1231,N_1557);
nor U2319 (N_2319,N_1010,N_1737);
or U2320 (N_2320,N_1659,N_1437);
or U2321 (N_2321,N_1423,N_1588);
or U2322 (N_2322,N_1351,N_1312);
nor U2323 (N_2323,N_1927,N_1534);
or U2324 (N_2324,N_1262,N_1180);
or U2325 (N_2325,N_1428,N_1215);
and U2326 (N_2326,N_1946,N_1684);
nand U2327 (N_2327,N_1216,N_1604);
and U2328 (N_2328,N_1603,N_1551);
xnor U2329 (N_2329,N_1068,N_1348);
and U2330 (N_2330,N_1733,N_1255);
and U2331 (N_2331,N_1223,N_1067);
nand U2332 (N_2332,N_1137,N_1635);
and U2333 (N_2333,N_1949,N_1524);
and U2334 (N_2334,N_1238,N_1701);
nand U2335 (N_2335,N_1150,N_1072);
or U2336 (N_2336,N_1260,N_1058);
nand U2337 (N_2337,N_1502,N_1907);
nor U2338 (N_2338,N_1598,N_1129);
or U2339 (N_2339,N_1905,N_1800);
nand U2340 (N_2340,N_1859,N_1530);
and U2341 (N_2341,N_1197,N_1693);
nor U2342 (N_2342,N_1002,N_1988);
nand U2343 (N_2343,N_1411,N_1828);
and U2344 (N_2344,N_1678,N_1661);
nor U2345 (N_2345,N_1877,N_1839);
or U2346 (N_2346,N_1853,N_1321);
nor U2347 (N_2347,N_1421,N_1981);
nor U2348 (N_2348,N_1908,N_1406);
and U2349 (N_2349,N_1871,N_1612);
or U2350 (N_2350,N_1688,N_1504);
and U2351 (N_2351,N_1094,N_1032);
and U2352 (N_2352,N_1290,N_1337);
and U2353 (N_2353,N_1541,N_1947);
and U2354 (N_2354,N_1207,N_1178);
nand U2355 (N_2355,N_1723,N_1948);
nand U2356 (N_2356,N_1466,N_1110);
nor U2357 (N_2357,N_1099,N_1564);
nor U2358 (N_2358,N_1864,N_1813);
xnor U2359 (N_2359,N_1143,N_1132);
or U2360 (N_2360,N_1978,N_1641);
and U2361 (N_2361,N_1109,N_1532);
nand U2362 (N_2362,N_1329,N_1793);
and U2363 (N_2363,N_1765,N_1024);
nand U2364 (N_2364,N_1647,N_1022);
nand U2365 (N_2365,N_1631,N_1218);
nand U2366 (N_2366,N_1950,N_1518);
and U2367 (N_2367,N_1649,N_1537);
nor U2368 (N_2368,N_1280,N_1835);
and U2369 (N_2369,N_1064,N_1244);
or U2370 (N_2370,N_1352,N_1953);
nor U2371 (N_2371,N_1951,N_1681);
or U2372 (N_2372,N_1347,N_1582);
or U2373 (N_2373,N_1627,N_1628);
and U2374 (N_2374,N_1126,N_1849);
and U2375 (N_2375,N_1250,N_1761);
nand U2376 (N_2376,N_1794,N_1492);
xnor U2377 (N_2377,N_1971,N_1186);
xor U2378 (N_2378,N_1535,N_1571);
nor U2379 (N_2379,N_1709,N_1118);
or U2380 (N_2380,N_1827,N_1247);
and U2381 (N_2381,N_1655,N_1997);
and U2382 (N_2382,N_1100,N_1893);
or U2383 (N_2383,N_1334,N_1880);
nor U2384 (N_2384,N_1904,N_1922);
nand U2385 (N_2385,N_1909,N_1166);
nand U2386 (N_2386,N_1433,N_1455);
or U2387 (N_2387,N_1497,N_1083);
nand U2388 (N_2388,N_1986,N_1481);
and U2389 (N_2389,N_1401,N_1377);
or U2390 (N_2390,N_1937,N_1622);
nor U2391 (N_2391,N_1677,N_1656);
xnor U2392 (N_2392,N_1784,N_1368);
and U2393 (N_2393,N_1621,N_1624);
nor U2394 (N_2394,N_1606,N_1374);
nor U2395 (N_2395,N_1891,N_1846);
and U2396 (N_2396,N_1101,N_1275);
nor U2397 (N_2397,N_1387,N_1682);
nor U2398 (N_2398,N_1727,N_1114);
or U2399 (N_2399,N_1742,N_1934);
nand U2400 (N_2400,N_1441,N_1868);
nand U2401 (N_2401,N_1327,N_1560);
or U2402 (N_2402,N_1753,N_1370);
or U2403 (N_2403,N_1308,N_1884);
or U2404 (N_2404,N_1025,N_1498);
nand U2405 (N_2405,N_1339,N_1664);
nand U2406 (N_2406,N_1386,N_1917);
or U2407 (N_2407,N_1371,N_1921);
nand U2408 (N_2408,N_1470,N_1865);
nand U2409 (N_2409,N_1527,N_1888);
nand U2410 (N_2410,N_1055,N_1556);
nand U2411 (N_2411,N_1985,N_1174);
or U2412 (N_2412,N_1040,N_1468);
and U2413 (N_2413,N_1362,N_1690);
nand U2414 (N_2414,N_1671,N_1452);
nor U2415 (N_2415,N_1417,N_1548);
or U2416 (N_2416,N_1722,N_1686);
and U2417 (N_2417,N_1307,N_1832);
xnor U2418 (N_2418,N_1300,N_1956);
or U2419 (N_2419,N_1895,N_1463);
or U2420 (N_2420,N_1378,N_1413);
nand U2421 (N_2421,N_1461,N_1252);
and U2422 (N_2422,N_1824,N_1422);
nor U2423 (N_2423,N_1366,N_1325);
nand U2424 (N_2424,N_1910,N_1175);
nor U2425 (N_2425,N_1775,N_1233);
and U2426 (N_2426,N_1616,N_1273);
and U2427 (N_2427,N_1573,N_1397);
and U2428 (N_2428,N_1756,N_1167);
nor U2429 (N_2429,N_1769,N_1395);
nand U2430 (N_2430,N_1361,N_1182);
and U2431 (N_2431,N_1168,N_1698);
nand U2432 (N_2432,N_1620,N_1385);
nand U2433 (N_2433,N_1840,N_1807);
nor U2434 (N_2434,N_1277,N_1332);
nor U2435 (N_2435,N_1811,N_1837);
nor U2436 (N_2436,N_1516,N_1343);
nor U2437 (N_2437,N_1102,N_1593);
nand U2438 (N_2438,N_1770,N_1633);
nand U2439 (N_2439,N_1299,N_1979);
or U2440 (N_2440,N_1831,N_1957);
nor U2441 (N_2441,N_1842,N_1008);
nor U2442 (N_2442,N_1683,N_1521);
nand U2443 (N_2443,N_1528,N_1919);
nand U2444 (N_2444,N_1699,N_1342);
and U2445 (N_2445,N_1791,N_1561);
nor U2446 (N_2446,N_1075,N_1786);
nor U2447 (N_2447,N_1424,N_1578);
or U2448 (N_2448,N_1670,N_1222);
and U2449 (N_2449,N_1817,N_1772);
nand U2450 (N_2450,N_1407,N_1160);
and U2451 (N_2451,N_1098,N_1382);
or U2452 (N_2452,N_1605,N_1808);
nor U2453 (N_2453,N_1235,N_1330);
nand U2454 (N_2454,N_1311,N_1349);
or U2455 (N_2455,N_1074,N_1944);
or U2456 (N_2456,N_1001,N_1117);
and U2457 (N_2457,N_1930,N_1090);
nand U2458 (N_2458,N_1198,N_1326);
or U2459 (N_2459,N_1843,N_1855);
or U2460 (N_2460,N_1096,N_1363);
or U2461 (N_2461,N_1125,N_1052);
and U2462 (N_2462,N_1088,N_1236);
or U2463 (N_2463,N_1446,N_1145);
nor U2464 (N_2464,N_1552,N_1587);
and U2465 (N_2465,N_1816,N_1513);
or U2466 (N_2466,N_1202,N_1479);
and U2467 (N_2467,N_1066,N_1217);
nor U2468 (N_2468,N_1211,N_1301);
nor U2469 (N_2469,N_1286,N_1785);
xor U2470 (N_2470,N_1767,N_1707);
or U2471 (N_2471,N_1925,N_1566);
and U2472 (N_2472,N_1583,N_1159);
nor U2473 (N_2473,N_1037,N_1309);
nor U2474 (N_2474,N_1974,N_1638);
nor U2475 (N_2475,N_1496,N_1237);
xnor U2476 (N_2476,N_1404,N_1874);
nand U2477 (N_2477,N_1264,N_1149);
or U2478 (N_2478,N_1878,N_1338);
nand U2479 (N_2479,N_1523,N_1696);
and U2480 (N_2480,N_1972,N_1459);
and U2481 (N_2481,N_1862,N_1464);
nor U2482 (N_2482,N_1806,N_1491);
nor U2483 (N_2483,N_1369,N_1777);
nor U2484 (N_2484,N_1920,N_1938);
or U2485 (N_2485,N_1897,N_1254);
nand U2486 (N_2486,N_1882,N_1687);
and U2487 (N_2487,N_1476,N_1804);
or U2488 (N_2488,N_1209,N_1029);
nor U2489 (N_2489,N_1151,N_1703);
and U2490 (N_2490,N_1751,N_1323);
nor U2491 (N_2491,N_1567,N_1901);
nor U2492 (N_2492,N_1797,N_1869);
nand U2493 (N_2493,N_1591,N_1936);
nor U2494 (N_2494,N_1396,N_1170);
nor U2495 (N_2495,N_1220,N_1165);
or U2496 (N_2496,N_1354,N_1983);
or U2497 (N_2497,N_1992,N_1980);
and U2498 (N_2498,N_1975,N_1398);
or U2499 (N_2499,N_1142,N_1998);
nor U2500 (N_2500,N_1447,N_1962);
nand U2501 (N_2501,N_1261,N_1965);
or U2502 (N_2502,N_1854,N_1847);
and U2503 (N_2503,N_1357,N_1334);
nor U2504 (N_2504,N_1723,N_1286);
and U2505 (N_2505,N_1805,N_1015);
nor U2506 (N_2506,N_1881,N_1457);
xor U2507 (N_2507,N_1656,N_1835);
and U2508 (N_2508,N_1875,N_1560);
and U2509 (N_2509,N_1318,N_1446);
and U2510 (N_2510,N_1133,N_1857);
nor U2511 (N_2511,N_1837,N_1602);
nor U2512 (N_2512,N_1415,N_1836);
and U2513 (N_2513,N_1862,N_1949);
and U2514 (N_2514,N_1251,N_1770);
nor U2515 (N_2515,N_1889,N_1430);
and U2516 (N_2516,N_1985,N_1163);
or U2517 (N_2517,N_1246,N_1942);
and U2518 (N_2518,N_1018,N_1940);
and U2519 (N_2519,N_1479,N_1236);
nor U2520 (N_2520,N_1550,N_1055);
nand U2521 (N_2521,N_1827,N_1276);
nand U2522 (N_2522,N_1053,N_1729);
nor U2523 (N_2523,N_1264,N_1215);
and U2524 (N_2524,N_1442,N_1743);
and U2525 (N_2525,N_1230,N_1685);
or U2526 (N_2526,N_1511,N_1474);
nor U2527 (N_2527,N_1592,N_1490);
and U2528 (N_2528,N_1733,N_1526);
or U2529 (N_2529,N_1529,N_1029);
or U2530 (N_2530,N_1752,N_1561);
nand U2531 (N_2531,N_1800,N_1987);
nor U2532 (N_2532,N_1749,N_1711);
nand U2533 (N_2533,N_1835,N_1607);
and U2534 (N_2534,N_1211,N_1447);
nand U2535 (N_2535,N_1808,N_1722);
or U2536 (N_2536,N_1485,N_1290);
and U2537 (N_2537,N_1509,N_1038);
or U2538 (N_2538,N_1120,N_1925);
nor U2539 (N_2539,N_1506,N_1002);
xor U2540 (N_2540,N_1595,N_1416);
and U2541 (N_2541,N_1995,N_1729);
or U2542 (N_2542,N_1349,N_1768);
nand U2543 (N_2543,N_1362,N_1993);
and U2544 (N_2544,N_1181,N_1521);
nand U2545 (N_2545,N_1589,N_1626);
nand U2546 (N_2546,N_1294,N_1945);
or U2547 (N_2547,N_1308,N_1755);
and U2548 (N_2548,N_1514,N_1812);
nand U2549 (N_2549,N_1710,N_1986);
or U2550 (N_2550,N_1357,N_1729);
or U2551 (N_2551,N_1966,N_1303);
xor U2552 (N_2552,N_1738,N_1493);
or U2553 (N_2553,N_1124,N_1905);
and U2554 (N_2554,N_1053,N_1334);
or U2555 (N_2555,N_1336,N_1207);
nand U2556 (N_2556,N_1784,N_1129);
and U2557 (N_2557,N_1003,N_1508);
nor U2558 (N_2558,N_1982,N_1203);
nor U2559 (N_2559,N_1763,N_1947);
nand U2560 (N_2560,N_1725,N_1930);
nor U2561 (N_2561,N_1640,N_1158);
and U2562 (N_2562,N_1880,N_1246);
or U2563 (N_2563,N_1056,N_1567);
or U2564 (N_2564,N_1046,N_1732);
nor U2565 (N_2565,N_1349,N_1456);
xnor U2566 (N_2566,N_1684,N_1156);
and U2567 (N_2567,N_1240,N_1584);
and U2568 (N_2568,N_1861,N_1342);
and U2569 (N_2569,N_1950,N_1301);
and U2570 (N_2570,N_1112,N_1157);
nor U2571 (N_2571,N_1097,N_1274);
nand U2572 (N_2572,N_1623,N_1522);
nand U2573 (N_2573,N_1255,N_1177);
or U2574 (N_2574,N_1373,N_1029);
nor U2575 (N_2575,N_1928,N_1190);
nand U2576 (N_2576,N_1390,N_1474);
or U2577 (N_2577,N_1629,N_1254);
nor U2578 (N_2578,N_1269,N_1097);
or U2579 (N_2579,N_1127,N_1412);
or U2580 (N_2580,N_1696,N_1817);
nor U2581 (N_2581,N_1487,N_1586);
nor U2582 (N_2582,N_1745,N_1524);
and U2583 (N_2583,N_1872,N_1657);
nand U2584 (N_2584,N_1757,N_1626);
nand U2585 (N_2585,N_1956,N_1302);
or U2586 (N_2586,N_1915,N_1601);
and U2587 (N_2587,N_1477,N_1664);
and U2588 (N_2588,N_1071,N_1817);
or U2589 (N_2589,N_1122,N_1091);
or U2590 (N_2590,N_1653,N_1233);
nor U2591 (N_2591,N_1453,N_1547);
nand U2592 (N_2592,N_1870,N_1905);
or U2593 (N_2593,N_1281,N_1345);
nor U2594 (N_2594,N_1650,N_1988);
and U2595 (N_2595,N_1025,N_1950);
nand U2596 (N_2596,N_1482,N_1181);
and U2597 (N_2597,N_1317,N_1877);
nor U2598 (N_2598,N_1337,N_1799);
or U2599 (N_2599,N_1020,N_1186);
nand U2600 (N_2600,N_1863,N_1124);
or U2601 (N_2601,N_1032,N_1375);
and U2602 (N_2602,N_1633,N_1719);
nor U2603 (N_2603,N_1917,N_1983);
nand U2604 (N_2604,N_1108,N_1336);
nand U2605 (N_2605,N_1229,N_1939);
nor U2606 (N_2606,N_1124,N_1911);
nand U2607 (N_2607,N_1459,N_1300);
nor U2608 (N_2608,N_1600,N_1066);
nand U2609 (N_2609,N_1219,N_1940);
nand U2610 (N_2610,N_1608,N_1824);
and U2611 (N_2611,N_1883,N_1365);
nand U2612 (N_2612,N_1470,N_1924);
nor U2613 (N_2613,N_1018,N_1081);
nor U2614 (N_2614,N_1100,N_1565);
or U2615 (N_2615,N_1365,N_1407);
and U2616 (N_2616,N_1027,N_1677);
nand U2617 (N_2617,N_1109,N_1584);
or U2618 (N_2618,N_1244,N_1267);
and U2619 (N_2619,N_1994,N_1467);
xnor U2620 (N_2620,N_1385,N_1168);
or U2621 (N_2621,N_1608,N_1296);
nor U2622 (N_2622,N_1901,N_1394);
nand U2623 (N_2623,N_1616,N_1093);
nand U2624 (N_2624,N_1004,N_1403);
and U2625 (N_2625,N_1649,N_1326);
nor U2626 (N_2626,N_1212,N_1083);
or U2627 (N_2627,N_1177,N_1895);
nor U2628 (N_2628,N_1914,N_1243);
or U2629 (N_2629,N_1729,N_1282);
nand U2630 (N_2630,N_1819,N_1686);
and U2631 (N_2631,N_1344,N_1737);
nor U2632 (N_2632,N_1530,N_1834);
nor U2633 (N_2633,N_1217,N_1616);
and U2634 (N_2634,N_1513,N_1000);
nand U2635 (N_2635,N_1901,N_1190);
nand U2636 (N_2636,N_1339,N_1235);
and U2637 (N_2637,N_1654,N_1100);
nor U2638 (N_2638,N_1406,N_1762);
and U2639 (N_2639,N_1794,N_1577);
nor U2640 (N_2640,N_1464,N_1448);
or U2641 (N_2641,N_1019,N_1806);
or U2642 (N_2642,N_1653,N_1747);
nor U2643 (N_2643,N_1345,N_1505);
and U2644 (N_2644,N_1833,N_1138);
nor U2645 (N_2645,N_1981,N_1858);
and U2646 (N_2646,N_1062,N_1576);
and U2647 (N_2647,N_1646,N_1097);
nand U2648 (N_2648,N_1119,N_1246);
nor U2649 (N_2649,N_1643,N_1441);
nand U2650 (N_2650,N_1432,N_1173);
or U2651 (N_2651,N_1199,N_1252);
nand U2652 (N_2652,N_1544,N_1848);
nand U2653 (N_2653,N_1407,N_1313);
nor U2654 (N_2654,N_1492,N_1681);
or U2655 (N_2655,N_1211,N_1939);
nand U2656 (N_2656,N_1631,N_1879);
and U2657 (N_2657,N_1522,N_1314);
and U2658 (N_2658,N_1710,N_1122);
xor U2659 (N_2659,N_1656,N_1359);
and U2660 (N_2660,N_1527,N_1733);
and U2661 (N_2661,N_1144,N_1014);
or U2662 (N_2662,N_1240,N_1090);
nor U2663 (N_2663,N_1139,N_1682);
and U2664 (N_2664,N_1206,N_1887);
nor U2665 (N_2665,N_1380,N_1228);
and U2666 (N_2666,N_1755,N_1062);
nand U2667 (N_2667,N_1092,N_1058);
or U2668 (N_2668,N_1718,N_1598);
or U2669 (N_2669,N_1777,N_1316);
nand U2670 (N_2670,N_1583,N_1360);
nand U2671 (N_2671,N_1019,N_1656);
or U2672 (N_2672,N_1941,N_1422);
or U2673 (N_2673,N_1424,N_1299);
and U2674 (N_2674,N_1179,N_1021);
or U2675 (N_2675,N_1229,N_1769);
or U2676 (N_2676,N_1984,N_1194);
nand U2677 (N_2677,N_1710,N_1453);
nor U2678 (N_2678,N_1644,N_1118);
or U2679 (N_2679,N_1816,N_1650);
nand U2680 (N_2680,N_1218,N_1378);
and U2681 (N_2681,N_1809,N_1885);
nor U2682 (N_2682,N_1850,N_1608);
or U2683 (N_2683,N_1032,N_1913);
nand U2684 (N_2684,N_1602,N_1003);
nor U2685 (N_2685,N_1417,N_1083);
nand U2686 (N_2686,N_1681,N_1659);
or U2687 (N_2687,N_1019,N_1565);
and U2688 (N_2688,N_1630,N_1769);
nand U2689 (N_2689,N_1311,N_1491);
and U2690 (N_2690,N_1366,N_1936);
nor U2691 (N_2691,N_1667,N_1907);
nor U2692 (N_2692,N_1407,N_1186);
or U2693 (N_2693,N_1764,N_1316);
nand U2694 (N_2694,N_1911,N_1707);
nand U2695 (N_2695,N_1897,N_1590);
and U2696 (N_2696,N_1115,N_1681);
and U2697 (N_2697,N_1244,N_1669);
or U2698 (N_2698,N_1915,N_1341);
nor U2699 (N_2699,N_1862,N_1733);
or U2700 (N_2700,N_1500,N_1696);
and U2701 (N_2701,N_1024,N_1966);
and U2702 (N_2702,N_1406,N_1939);
nor U2703 (N_2703,N_1684,N_1392);
and U2704 (N_2704,N_1614,N_1818);
nand U2705 (N_2705,N_1857,N_1607);
and U2706 (N_2706,N_1928,N_1844);
or U2707 (N_2707,N_1794,N_1006);
or U2708 (N_2708,N_1188,N_1105);
or U2709 (N_2709,N_1193,N_1920);
or U2710 (N_2710,N_1826,N_1192);
nand U2711 (N_2711,N_1683,N_1332);
nand U2712 (N_2712,N_1501,N_1620);
and U2713 (N_2713,N_1769,N_1904);
nor U2714 (N_2714,N_1431,N_1800);
nand U2715 (N_2715,N_1102,N_1710);
nand U2716 (N_2716,N_1911,N_1039);
and U2717 (N_2717,N_1863,N_1770);
and U2718 (N_2718,N_1236,N_1796);
nor U2719 (N_2719,N_1950,N_1160);
and U2720 (N_2720,N_1919,N_1834);
nand U2721 (N_2721,N_1057,N_1767);
nor U2722 (N_2722,N_1065,N_1246);
nor U2723 (N_2723,N_1167,N_1728);
nor U2724 (N_2724,N_1280,N_1880);
nand U2725 (N_2725,N_1331,N_1568);
nor U2726 (N_2726,N_1919,N_1492);
or U2727 (N_2727,N_1181,N_1573);
nand U2728 (N_2728,N_1589,N_1206);
or U2729 (N_2729,N_1218,N_1455);
or U2730 (N_2730,N_1214,N_1692);
or U2731 (N_2731,N_1999,N_1868);
or U2732 (N_2732,N_1501,N_1236);
nor U2733 (N_2733,N_1327,N_1303);
or U2734 (N_2734,N_1117,N_1926);
nor U2735 (N_2735,N_1917,N_1972);
nand U2736 (N_2736,N_1146,N_1326);
nor U2737 (N_2737,N_1497,N_1088);
nand U2738 (N_2738,N_1317,N_1353);
or U2739 (N_2739,N_1113,N_1517);
nor U2740 (N_2740,N_1340,N_1293);
nand U2741 (N_2741,N_1082,N_1443);
or U2742 (N_2742,N_1081,N_1468);
or U2743 (N_2743,N_1702,N_1219);
nor U2744 (N_2744,N_1956,N_1864);
or U2745 (N_2745,N_1921,N_1032);
and U2746 (N_2746,N_1067,N_1205);
or U2747 (N_2747,N_1980,N_1695);
or U2748 (N_2748,N_1172,N_1941);
xnor U2749 (N_2749,N_1007,N_1864);
nor U2750 (N_2750,N_1819,N_1591);
xor U2751 (N_2751,N_1318,N_1426);
nand U2752 (N_2752,N_1133,N_1002);
nor U2753 (N_2753,N_1848,N_1979);
nand U2754 (N_2754,N_1651,N_1868);
nor U2755 (N_2755,N_1779,N_1314);
or U2756 (N_2756,N_1640,N_1933);
nor U2757 (N_2757,N_1267,N_1721);
xnor U2758 (N_2758,N_1309,N_1663);
nand U2759 (N_2759,N_1121,N_1700);
nand U2760 (N_2760,N_1921,N_1933);
or U2761 (N_2761,N_1738,N_1674);
or U2762 (N_2762,N_1223,N_1852);
and U2763 (N_2763,N_1668,N_1034);
xor U2764 (N_2764,N_1361,N_1378);
or U2765 (N_2765,N_1499,N_1427);
and U2766 (N_2766,N_1836,N_1998);
or U2767 (N_2767,N_1621,N_1688);
nor U2768 (N_2768,N_1265,N_1970);
nor U2769 (N_2769,N_1372,N_1743);
and U2770 (N_2770,N_1563,N_1838);
nor U2771 (N_2771,N_1840,N_1255);
and U2772 (N_2772,N_1606,N_1206);
and U2773 (N_2773,N_1811,N_1939);
nand U2774 (N_2774,N_1340,N_1565);
or U2775 (N_2775,N_1420,N_1969);
and U2776 (N_2776,N_1966,N_1636);
nor U2777 (N_2777,N_1984,N_1985);
nor U2778 (N_2778,N_1124,N_1102);
nand U2779 (N_2779,N_1263,N_1074);
or U2780 (N_2780,N_1009,N_1199);
nand U2781 (N_2781,N_1319,N_1288);
and U2782 (N_2782,N_1183,N_1461);
nor U2783 (N_2783,N_1748,N_1307);
nor U2784 (N_2784,N_1553,N_1172);
nand U2785 (N_2785,N_1664,N_1376);
nand U2786 (N_2786,N_1279,N_1164);
nor U2787 (N_2787,N_1110,N_1831);
or U2788 (N_2788,N_1594,N_1384);
or U2789 (N_2789,N_1382,N_1312);
nor U2790 (N_2790,N_1345,N_1066);
nand U2791 (N_2791,N_1935,N_1133);
nor U2792 (N_2792,N_1662,N_1668);
nand U2793 (N_2793,N_1948,N_1070);
and U2794 (N_2794,N_1229,N_1464);
and U2795 (N_2795,N_1603,N_1878);
or U2796 (N_2796,N_1502,N_1895);
nand U2797 (N_2797,N_1777,N_1319);
nand U2798 (N_2798,N_1520,N_1044);
nor U2799 (N_2799,N_1950,N_1555);
and U2800 (N_2800,N_1711,N_1928);
or U2801 (N_2801,N_1675,N_1753);
nor U2802 (N_2802,N_1468,N_1421);
or U2803 (N_2803,N_1930,N_1289);
nand U2804 (N_2804,N_1891,N_1815);
and U2805 (N_2805,N_1288,N_1019);
and U2806 (N_2806,N_1099,N_1942);
xnor U2807 (N_2807,N_1954,N_1332);
nor U2808 (N_2808,N_1768,N_1038);
and U2809 (N_2809,N_1133,N_1439);
nand U2810 (N_2810,N_1488,N_1807);
or U2811 (N_2811,N_1091,N_1590);
nand U2812 (N_2812,N_1575,N_1125);
or U2813 (N_2813,N_1307,N_1709);
and U2814 (N_2814,N_1589,N_1280);
and U2815 (N_2815,N_1200,N_1531);
nor U2816 (N_2816,N_1069,N_1718);
nor U2817 (N_2817,N_1024,N_1648);
nor U2818 (N_2818,N_1929,N_1851);
and U2819 (N_2819,N_1660,N_1535);
or U2820 (N_2820,N_1189,N_1664);
or U2821 (N_2821,N_1845,N_1436);
and U2822 (N_2822,N_1405,N_1463);
nor U2823 (N_2823,N_1809,N_1729);
nor U2824 (N_2824,N_1845,N_1040);
and U2825 (N_2825,N_1511,N_1032);
nor U2826 (N_2826,N_1952,N_1080);
nand U2827 (N_2827,N_1946,N_1415);
and U2828 (N_2828,N_1030,N_1419);
nor U2829 (N_2829,N_1301,N_1327);
nor U2830 (N_2830,N_1715,N_1127);
nand U2831 (N_2831,N_1792,N_1696);
nor U2832 (N_2832,N_1284,N_1673);
or U2833 (N_2833,N_1363,N_1201);
nand U2834 (N_2834,N_1846,N_1603);
or U2835 (N_2835,N_1996,N_1886);
or U2836 (N_2836,N_1047,N_1337);
or U2837 (N_2837,N_1016,N_1220);
and U2838 (N_2838,N_1137,N_1022);
nand U2839 (N_2839,N_1464,N_1943);
and U2840 (N_2840,N_1172,N_1783);
nand U2841 (N_2841,N_1148,N_1407);
nor U2842 (N_2842,N_1998,N_1369);
or U2843 (N_2843,N_1314,N_1832);
or U2844 (N_2844,N_1658,N_1884);
nand U2845 (N_2845,N_1097,N_1903);
and U2846 (N_2846,N_1516,N_1639);
or U2847 (N_2847,N_1222,N_1470);
xor U2848 (N_2848,N_1934,N_1898);
or U2849 (N_2849,N_1301,N_1295);
and U2850 (N_2850,N_1753,N_1480);
and U2851 (N_2851,N_1529,N_1677);
or U2852 (N_2852,N_1403,N_1801);
or U2853 (N_2853,N_1478,N_1675);
nor U2854 (N_2854,N_1785,N_1263);
nor U2855 (N_2855,N_1523,N_1686);
or U2856 (N_2856,N_1604,N_1467);
and U2857 (N_2857,N_1718,N_1224);
and U2858 (N_2858,N_1409,N_1560);
or U2859 (N_2859,N_1168,N_1536);
xnor U2860 (N_2860,N_1186,N_1382);
nand U2861 (N_2861,N_1008,N_1925);
nand U2862 (N_2862,N_1992,N_1001);
nor U2863 (N_2863,N_1586,N_1485);
and U2864 (N_2864,N_1555,N_1847);
nand U2865 (N_2865,N_1098,N_1444);
and U2866 (N_2866,N_1789,N_1218);
nor U2867 (N_2867,N_1059,N_1366);
nor U2868 (N_2868,N_1010,N_1661);
and U2869 (N_2869,N_1179,N_1873);
nor U2870 (N_2870,N_1578,N_1915);
nor U2871 (N_2871,N_1020,N_1539);
nand U2872 (N_2872,N_1318,N_1458);
nor U2873 (N_2873,N_1988,N_1264);
and U2874 (N_2874,N_1101,N_1216);
nor U2875 (N_2875,N_1034,N_1527);
nor U2876 (N_2876,N_1117,N_1428);
nor U2877 (N_2877,N_1841,N_1320);
and U2878 (N_2878,N_1565,N_1213);
nor U2879 (N_2879,N_1213,N_1291);
nand U2880 (N_2880,N_1883,N_1670);
nand U2881 (N_2881,N_1618,N_1133);
nand U2882 (N_2882,N_1695,N_1901);
nor U2883 (N_2883,N_1965,N_1454);
nor U2884 (N_2884,N_1557,N_1345);
or U2885 (N_2885,N_1971,N_1055);
and U2886 (N_2886,N_1089,N_1576);
nor U2887 (N_2887,N_1491,N_1360);
or U2888 (N_2888,N_1401,N_1507);
or U2889 (N_2889,N_1231,N_1908);
and U2890 (N_2890,N_1982,N_1841);
and U2891 (N_2891,N_1061,N_1928);
and U2892 (N_2892,N_1648,N_1192);
or U2893 (N_2893,N_1488,N_1977);
or U2894 (N_2894,N_1627,N_1481);
nor U2895 (N_2895,N_1471,N_1758);
and U2896 (N_2896,N_1748,N_1040);
nor U2897 (N_2897,N_1998,N_1726);
nor U2898 (N_2898,N_1124,N_1041);
nand U2899 (N_2899,N_1955,N_1747);
and U2900 (N_2900,N_1638,N_1414);
or U2901 (N_2901,N_1571,N_1725);
and U2902 (N_2902,N_1208,N_1950);
nor U2903 (N_2903,N_1626,N_1047);
xor U2904 (N_2904,N_1076,N_1806);
and U2905 (N_2905,N_1203,N_1359);
nor U2906 (N_2906,N_1443,N_1439);
and U2907 (N_2907,N_1813,N_1833);
nand U2908 (N_2908,N_1315,N_1897);
nand U2909 (N_2909,N_1698,N_1697);
nand U2910 (N_2910,N_1350,N_1454);
or U2911 (N_2911,N_1885,N_1430);
nor U2912 (N_2912,N_1756,N_1487);
or U2913 (N_2913,N_1534,N_1310);
or U2914 (N_2914,N_1318,N_1730);
or U2915 (N_2915,N_1462,N_1571);
nand U2916 (N_2916,N_1789,N_1699);
nor U2917 (N_2917,N_1242,N_1573);
nor U2918 (N_2918,N_1696,N_1238);
and U2919 (N_2919,N_1309,N_1481);
nand U2920 (N_2920,N_1575,N_1495);
nor U2921 (N_2921,N_1153,N_1349);
nand U2922 (N_2922,N_1588,N_1348);
nor U2923 (N_2923,N_1462,N_1003);
nor U2924 (N_2924,N_1473,N_1880);
or U2925 (N_2925,N_1667,N_1775);
nand U2926 (N_2926,N_1976,N_1355);
nor U2927 (N_2927,N_1437,N_1527);
and U2928 (N_2928,N_1682,N_1350);
nor U2929 (N_2929,N_1791,N_1104);
or U2930 (N_2930,N_1420,N_1947);
nor U2931 (N_2931,N_1556,N_1962);
and U2932 (N_2932,N_1081,N_1832);
nor U2933 (N_2933,N_1046,N_1436);
and U2934 (N_2934,N_1253,N_1349);
or U2935 (N_2935,N_1286,N_1065);
nor U2936 (N_2936,N_1131,N_1171);
nand U2937 (N_2937,N_1358,N_1203);
or U2938 (N_2938,N_1859,N_1893);
or U2939 (N_2939,N_1013,N_1390);
and U2940 (N_2940,N_1010,N_1796);
and U2941 (N_2941,N_1479,N_1357);
nor U2942 (N_2942,N_1086,N_1054);
or U2943 (N_2943,N_1618,N_1086);
and U2944 (N_2944,N_1385,N_1057);
nor U2945 (N_2945,N_1471,N_1414);
nand U2946 (N_2946,N_1616,N_1816);
and U2947 (N_2947,N_1181,N_1041);
nand U2948 (N_2948,N_1346,N_1933);
and U2949 (N_2949,N_1339,N_1072);
nand U2950 (N_2950,N_1209,N_1664);
and U2951 (N_2951,N_1160,N_1636);
nand U2952 (N_2952,N_1340,N_1539);
or U2953 (N_2953,N_1702,N_1117);
nor U2954 (N_2954,N_1145,N_1386);
nor U2955 (N_2955,N_1706,N_1050);
or U2956 (N_2956,N_1516,N_1506);
xnor U2957 (N_2957,N_1899,N_1759);
nor U2958 (N_2958,N_1289,N_1381);
or U2959 (N_2959,N_1082,N_1682);
nor U2960 (N_2960,N_1110,N_1124);
nand U2961 (N_2961,N_1490,N_1952);
nand U2962 (N_2962,N_1322,N_1020);
nand U2963 (N_2963,N_1431,N_1200);
nor U2964 (N_2964,N_1298,N_1054);
xnor U2965 (N_2965,N_1538,N_1877);
nor U2966 (N_2966,N_1094,N_1150);
or U2967 (N_2967,N_1048,N_1880);
nand U2968 (N_2968,N_1459,N_1408);
and U2969 (N_2969,N_1753,N_1896);
nor U2970 (N_2970,N_1361,N_1031);
nand U2971 (N_2971,N_1827,N_1237);
nor U2972 (N_2972,N_1564,N_1937);
nor U2973 (N_2973,N_1323,N_1305);
nor U2974 (N_2974,N_1655,N_1492);
nand U2975 (N_2975,N_1529,N_1189);
nor U2976 (N_2976,N_1962,N_1718);
nand U2977 (N_2977,N_1882,N_1326);
nor U2978 (N_2978,N_1934,N_1377);
and U2979 (N_2979,N_1596,N_1887);
or U2980 (N_2980,N_1962,N_1651);
or U2981 (N_2981,N_1853,N_1619);
nand U2982 (N_2982,N_1130,N_1157);
nand U2983 (N_2983,N_1616,N_1052);
or U2984 (N_2984,N_1932,N_1441);
nand U2985 (N_2985,N_1417,N_1358);
or U2986 (N_2986,N_1529,N_1683);
and U2987 (N_2987,N_1308,N_1098);
nor U2988 (N_2988,N_1730,N_1449);
nand U2989 (N_2989,N_1014,N_1158);
nand U2990 (N_2990,N_1081,N_1238);
or U2991 (N_2991,N_1759,N_1939);
nand U2992 (N_2992,N_1506,N_1897);
nor U2993 (N_2993,N_1529,N_1272);
nor U2994 (N_2994,N_1145,N_1817);
nor U2995 (N_2995,N_1224,N_1849);
nand U2996 (N_2996,N_1680,N_1772);
nand U2997 (N_2997,N_1977,N_1354);
nand U2998 (N_2998,N_1998,N_1720);
or U2999 (N_2999,N_1510,N_1523);
nand U3000 (N_3000,N_2072,N_2765);
or U3001 (N_3001,N_2291,N_2273);
and U3002 (N_3002,N_2359,N_2536);
nand U3003 (N_3003,N_2325,N_2432);
nand U3004 (N_3004,N_2349,N_2414);
and U3005 (N_3005,N_2712,N_2292);
nand U3006 (N_3006,N_2129,N_2926);
and U3007 (N_3007,N_2831,N_2368);
or U3008 (N_3008,N_2340,N_2443);
nand U3009 (N_3009,N_2835,N_2295);
xnor U3010 (N_3010,N_2391,N_2800);
nand U3011 (N_3011,N_2724,N_2896);
nor U3012 (N_3012,N_2895,N_2616);
nor U3013 (N_3013,N_2269,N_2753);
xnor U3014 (N_3014,N_2634,N_2708);
nand U3015 (N_3015,N_2604,N_2675);
or U3016 (N_3016,N_2839,N_2646);
nand U3017 (N_3017,N_2271,N_2216);
nor U3018 (N_3018,N_2331,N_2783);
or U3019 (N_3019,N_2343,N_2672);
or U3020 (N_3020,N_2784,N_2163);
and U3021 (N_3021,N_2781,N_2294);
nor U3022 (N_3022,N_2931,N_2602);
nand U3023 (N_3023,N_2205,N_2068);
or U3024 (N_3024,N_2597,N_2300);
nor U3025 (N_3025,N_2780,N_2668);
nor U3026 (N_3026,N_2339,N_2716);
and U3027 (N_3027,N_2946,N_2524);
nor U3028 (N_3028,N_2215,N_2875);
nor U3029 (N_3029,N_2410,N_2983);
or U3030 (N_3030,N_2945,N_2416);
or U3031 (N_3031,N_2876,N_2282);
or U3032 (N_3032,N_2182,N_2375);
nor U3033 (N_3033,N_2454,N_2513);
nor U3034 (N_3034,N_2417,N_2326);
and U3035 (N_3035,N_2050,N_2250);
nand U3036 (N_3036,N_2165,N_2899);
or U3037 (N_3037,N_2310,N_2592);
and U3038 (N_3038,N_2030,N_2322);
nand U3039 (N_3039,N_2976,N_2575);
nor U3040 (N_3040,N_2409,N_2957);
and U3041 (N_3041,N_2860,N_2396);
or U3042 (N_3042,N_2230,N_2846);
and U3043 (N_3043,N_2123,N_2609);
nor U3044 (N_3044,N_2799,N_2483);
and U3045 (N_3045,N_2166,N_2670);
nor U3046 (N_3046,N_2499,N_2244);
nand U3047 (N_3047,N_2234,N_2491);
nor U3048 (N_3048,N_2460,N_2015);
nor U3049 (N_3049,N_2438,N_2071);
nor U3050 (N_3050,N_2116,N_2943);
nand U3051 (N_3051,N_2551,N_2120);
and U3052 (N_3052,N_2678,N_2545);
xnor U3053 (N_3053,N_2654,N_2971);
or U3054 (N_3054,N_2757,N_2445);
or U3055 (N_3055,N_2117,N_2917);
and U3056 (N_3056,N_2306,N_2963);
nor U3057 (N_3057,N_2266,N_2630);
nand U3058 (N_3058,N_2973,N_2397);
nor U3059 (N_3059,N_2452,N_2162);
nand U3060 (N_3060,N_2884,N_2225);
nand U3061 (N_3061,N_2841,N_2840);
or U3062 (N_3062,N_2956,N_2160);
nor U3063 (N_3063,N_2179,N_2703);
or U3064 (N_3064,N_2309,N_2156);
or U3065 (N_3065,N_2744,N_2580);
and U3066 (N_3066,N_2374,N_2878);
or U3067 (N_3067,N_2067,N_2605);
or U3068 (N_3068,N_2267,N_2212);
or U3069 (N_3069,N_2314,N_2958);
nand U3070 (N_3070,N_2241,N_2455);
nor U3071 (N_3071,N_2995,N_2132);
or U3072 (N_3072,N_2084,N_2679);
nor U3073 (N_3073,N_2587,N_2879);
or U3074 (N_3074,N_2770,N_2924);
xor U3075 (N_3075,N_2001,N_2194);
nor U3076 (N_3076,N_2694,N_2754);
or U3077 (N_3077,N_2504,N_2528);
and U3078 (N_3078,N_2131,N_2704);
nor U3079 (N_3079,N_2874,N_2407);
or U3080 (N_3080,N_2978,N_2832);
and U3081 (N_3081,N_2869,N_2111);
or U3082 (N_3082,N_2265,N_2425);
or U3083 (N_3083,N_2953,N_2382);
nor U3084 (N_3084,N_2110,N_2022);
or U3085 (N_3085,N_2099,N_2600);
xor U3086 (N_3086,N_2626,N_2013);
and U3087 (N_3087,N_2862,N_2993);
nor U3088 (N_3088,N_2458,N_2248);
or U3089 (N_3089,N_2548,N_2938);
nor U3090 (N_3090,N_2175,N_2210);
nor U3091 (N_3091,N_2803,N_2632);
nand U3092 (N_3092,N_2420,N_2774);
and U3093 (N_3093,N_2520,N_2151);
or U3094 (N_3094,N_2702,N_2222);
or U3095 (N_3095,N_2251,N_2968);
or U3096 (N_3096,N_2168,N_2974);
and U3097 (N_3097,N_2933,N_2402);
and U3098 (N_3098,N_2737,N_2886);
and U3099 (N_3099,N_2619,N_2719);
nand U3100 (N_3100,N_2429,N_2219);
nand U3101 (N_3101,N_2355,N_2611);
or U3102 (N_3102,N_2797,N_2764);
nor U3103 (N_3103,N_2544,N_2239);
and U3104 (N_3104,N_2915,N_2124);
nor U3105 (N_3105,N_2910,N_2440);
and U3106 (N_3106,N_2950,N_2979);
nor U3107 (N_3107,N_2469,N_2433);
and U3108 (N_3108,N_2809,N_2039);
and U3109 (N_3109,N_2649,N_2944);
xnor U3110 (N_3110,N_2334,N_2959);
nor U3111 (N_3111,N_2388,N_2237);
nand U3112 (N_3112,N_2141,N_2823);
or U3113 (N_3113,N_2725,N_2379);
nand U3114 (N_3114,N_2404,N_2061);
and U3115 (N_3115,N_2487,N_2361);
nor U3116 (N_3116,N_2105,N_2298);
nand U3117 (N_3117,N_2934,N_2509);
nand U3118 (N_3118,N_2169,N_2246);
and U3119 (N_3119,N_2090,N_2519);
or U3120 (N_3120,N_2181,N_2734);
nand U3121 (N_3121,N_2762,N_2387);
and U3122 (N_3122,N_2655,N_2590);
nor U3123 (N_3123,N_2512,N_2488);
or U3124 (N_3124,N_2383,N_2275);
or U3125 (N_3125,N_2289,N_2709);
xnor U3126 (N_3126,N_2844,N_2189);
xor U3127 (N_3127,N_2572,N_2629);
and U3128 (N_3128,N_2494,N_2500);
nor U3129 (N_3129,N_2645,N_2197);
and U3130 (N_3130,N_2647,N_2501);
or U3131 (N_3131,N_2190,N_2523);
and U3132 (N_3132,N_2150,N_2739);
nand U3133 (N_3133,N_2948,N_2585);
nand U3134 (N_3134,N_2919,N_2970);
nand U3135 (N_3135,N_2546,N_2569);
and U3136 (N_3136,N_2813,N_2601);
and U3137 (N_3137,N_2280,N_2456);
nand U3138 (N_3138,N_2008,N_2430);
nand U3139 (N_3139,N_2408,N_2082);
nand U3140 (N_3140,N_2108,N_2400);
nor U3141 (N_3141,N_2559,N_2053);
and U3142 (N_3142,N_2459,N_2665);
and U3143 (N_3143,N_2913,N_2961);
nor U3144 (N_3144,N_2279,N_2393);
and U3145 (N_3145,N_2522,N_2384);
nand U3146 (N_3146,N_2486,N_2054);
nor U3147 (N_3147,N_2637,N_2173);
or U3148 (N_3148,N_2617,N_2947);
nor U3149 (N_3149,N_2441,N_2386);
and U3150 (N_3150,N_2373,N_2228);
or U3151 (N_3151,N_2720,N_2932);
or U3152 (N_3152,N_2439,N_2960);
nor U3153 (N_3153,N_2718,N_2826);
or U3154 (N_3154,N_2989,N_2381);
nand U3155 (N_3155,N_2907,N_2444);
or U3156 (N_3156,N_2235,N_2422);
and U3157 (N_3157,N_2988,N_2911);
nand U3158 (N_3158,N_2263,N_2367);
nand U3159 (N_3159,N_2598,N_2866);
nand U3160 (N_3160,N_2855,N_2567);
or U3161 (N_3161,N_2745,N_2385);
or U3162 (N_3162,N_2196,N_2640);
nor U3163 (N_3163,N_2790,N_2557);
or U3164 (N_3164,N_2200,N_2043);
or U3165 (N_3165,N_2977,N_2994);
or U3166 (N_3166,N_2178,N_2999);
or U3167 (N_3167,N_2788,N_2330);
or U3168 (N_3168,N_2650,N_2871);
and U3169 (N_3169,N_2936,N_2207);
and U3170 (N_3170,N_2005,N_2159);
and U3171 (N_3171,N_2850,N_2152);
or U3172 (N_3172,N_2051,N_2514);
and U3173 (N_3173,N_2584,N_2170);
nand U3174 (N_3174,N_2479,N_2482);
nor U3175 (N_3175,N_2312,N_2324);
or U3176 (N_3176,N_2633,N_2258);
or U3177 (N_3177,N_2543,N_2673);
or U3178 (N_3178,N_2038,N_2881);
nand U3179 (N_3179,N_2106,N_2508);
nor U3180 (N_3180,N_2740,N_2816);
nor U3181 (N_3181,N_2636,N_2758);
and U3182 (N_3182,N_2603,N_2133);
nand U3183 (N_3183,N_2510,N_2927);
and U3184 (N_3184,N_2337,N_2025);
nor U3185 (N_3185,N_2270,N_2511);
nor U3186 (N_3186,N_2648,N_2807);
and U3187 (N_3187,N_2772,N_2589);
and U3188 (N_3188,N_2883,N_2113);
and U3189 (N_3189,N_2329,N_2136);
nor U3190 (N_3190,N_2097,N_2320);
and U3191 (N_3191,N_2204,N_2864);
nor U3192 (N_3192,N_2837,N_2036);
nor U3193 (N_3193,N_2849,N_2940);
nor U3194 (N_3194,N_2127,N_2538);
nor U3195 (N_3195,N_2254,N_2664);
and U3196 (N_3196,N_2748,N_2699);
or U3197 (N_3197,N_2437,N_2527);
and U3198 (N_3198,N_2233,N_2607);
and U3199 (N_3199,N_2683,N_2727);
and U3200 (N_3200,N_2560,N_2231);
nand U3201 (N_3201,N_2517,N_2307);
and U3202 (N_3202,N_2506,N_2089);
xnor U3203 (N_3203,N_2746,N_2614);
or U3204 (N_3204,N_2347,N_2966);
or U3205 (N_3205,N_2570,N_2568);
and U3206 (N_3206,N_2463,N_2466);
nand U3207 (N_3207,N_2092,N_2010);
nor U3208 (N_3208,N_2177,N_2714);
or U3209 (N_3209,N_2722,N_2473);
or U3210 (N_3210,N_2338,N_2149);
nand U3211 (N_3211,N_2490,N_2588);
or U3212 (N_3212,N_2660,N_2767);
or U3213 (N_3213,N_2122,N_2492);
nor U3214 (N_3214,N_2293,N_2087);
nor U3215 (N_3215,N_2109,N_2651);
or U3216 (N_3216,N_2776,N_2804);
and U3217 (N_3217,N_2362,N_2889);
nand U3218 (N_3218,N_2327,N_2260);
nor U3219 (N_3219,N_2192,N_2139);
nand U3220 (N_3220,N_2897,N_2747);
or U3221 (N_3221,N_2058,N_2556);
nor U3222 (N_3222,N_2134,N_2872);
and U3223 (N_3223,N_2211,N_2352);
nor U3224 (N_3224,N_2980,N_2771);
nor U3225 (N_3225,N_2315,N_2154);
or U3226 (N_3226,N_2606,N_2056);
nor U3227 (N_3227,N_2024,N_2208);
and U3228 (N_3228,N_2736,N_2047);
and U3229 (N_3229,N_2778,N_2112);
and U3230 (N_3230,N_2345,N_2688);
nand U3231 (N_3231,N_2903,N_2902);
nand U3232 (N_3232,N_2641,N_2566);
or U3233 (N_3233,N_2256,N_2795);
and U3234 (N_3234,N_2729,N_2255);
nor U3235 (N_3235,N_2922,N_2775);
and U3236 (N_3236,N_2153,N_2526);
nand U3237 (N_3237,N_2521,N_2287);
nor U3238 (N_3238,N_2591,N_2264);
and U3239 (N_3239,N_2411,N_2079);
and U3240 (N_3240,N_2518,N_2065);
and U3241 (N_3241,N_2595,N_2029);
nor U3242 (N_3242,N_2984,N_2579);
and U3243 (N_3243,N_2887,N_2462);
nand U3244 (N_3244,N_2401,N_2873);
or U3245 (N_3245,N_2446,N_2863);
or U3246 (N_3246,N_2405,N_2002);
or U3247 (N_3247,N_2257,N_2777);
nor U3248 (N_3248,N_2146,N_2666);
nand U3249 (N_3249,N_2893,N_2706);
or U3250 (N_3250,N_2842,N_2048);
or U3251 (N_3251,N_2485,N_2095);
nand U3252 (N_3252,N_2217,N_2531);
xnor U3253 (N_3253,N_2019,N_2652);
nand U3254 (N_3254,N_2990,N_2890);
nor U3255 (N_3255,N_2370,N_2532);
nand U3256 (N_3256,N_2667,N_2137);
nand U3257 (N_3257,N_2565,N_2717);
and U3258 (N_3258,N_2125,N_2007);
nand U3259 (N_3259,N_2692,N_2376);
or U3260 (N_3260,N_2794,N_2562);
nand U3261 (N_3261,N_2535,N_2020);
and U3262 (N_3262,N_2333,N_2898);
or U3263 (N_3263,N_2080,N_2624);
and U3264 (N_3264,N_2877,N_2623);
or U3265 (N_3265,N_2540,N_2833);
and U3266 (N_3266,N_2610,N_2817);
nor U3267 (N_3267,N_2870,N_2676);
and U3268 (N_3268,N_2245,N_2822);
and U3269 (N_3269,N_2918,N_2415);
and U3270 (N_3270,N_2348,N_2925);
or U3271 (N_3271,N_2495,N_2593);
and U3272 (N_3272,N_2243,N_2805);
and U3273 (N_3273,N_2700,N_2353);
nor U3274 (N_3274,N_2697,N_2360);
nand U3275 (N_3275,N_2052,N_2830);
and U3276 (N_3276,N_2226,N_2858);
or U3277 (N_3277,N_2721,N_2653);
nand U3278 (N_3278,N_2929,N_2827);
and U3279 (N_3279,N_2608,N_2909);
or U3280 (N_3280,N_2836,N_2098);
nand U3281 (N_3281,N_2213,N_2026);
nor U3282 (N_3282,N_2031,N_2996);
or U3283 (N_3283,N_2272,N_2582);
and U3284 (N_3284,N_2920,N_2693);
nand U3285 (N_3285,N_2313,N_2332);
or U3286 (N_3286,N_2144,N_2076);
and U3287 (N_3287,N_2969,N_2656);
nor U3288 (N_3288,N_2905,N_2759);
and U3289 (N_3289,N_2465,N_2316);
nand U3290 (N_3290,N_2581,N_2760);
or U3291 (N_3291,N_2147,N_2042);
nor U3292 (N_3292,N_2715,N_2371);
or U3293 (N_3293,N_2921,N_2319);
nand U3294 (N_3294,N_2768,N_2811);
or U3295 (N_3295,N_2372,N_2752);
xor U3296 (N_3296,N_2854,N_2576);
and U3297 (N_3297,N_2423,N_2094);
or U3298 (N_3298,N_2102,N_2421);
and U3299 (N_3299,N_2554,N_2145);
nand U3300 (N_3300,N_2203,N_2399);
and U3301 (N_3301,N_2023,N_2563);
nor U3302 (N_3302,N_2135,N_2288);
xor U3303 (N_3303,N_2639,N_2435);
nor U3304 (N_3304,N_2088,N_2075);
or U3305 (N_3305,N_2782,N_2659);
and U3306 (N_3306,N_2555,N_2419);
or U3307 (N_3307,N_2558,N_2100);
nand U3308 (N_3308,N_2573,N_2808);
nor U3309 (N_3309,N_2086,N_2478);
nand U3310 (N_3310,N_2148,N_2657);
nand U3311 (N_3311,N_2009,N_2003);
nor U3312 (N_3312,N_2480,N_2986);
and U3313 (N_3313,N_2350,N_2221);
and U3314 (N_3314,N_2062,N_2539);
or U3315 (N_3315,N_2227,N_2730);
nand U3316 (N_3316,N_2856,N_2069);
nor U3317 (N_3317,N_2982,N_2828);
nor U3318 (N_3318,N_2262,N_2199);
nand U3319 (N_3319,N_2176,N_2793);
nand U3320 (N_3320,N_2365,N_2952);
and U3321 (N_3321,N_2906,N_2077);
nand U3322 (N_3322,N_2928,N_2935);
nor U3323 (N_3323,N_2060,N_2766);
nand U3324 (N_3324,N_2912,N_2686);
or U3325 (N_3325,N_2115,N_2450);
or U3326 (N_3326,N_2644,N_2779);
nor U3327 (N_3327,N_2364,N_2378);
or U3328 (N_3328,N_2468,N_2413);
nand U3329 (N_3329,N_2594,N_2357);
nand U3330 (N_3330,N_2238,N_2427);
nand U3331 (N_3331,N_2232,N_2843);
and U3332 (N_3332,N_2628,N_2426);
nand U3333 (N_3333,N_2363,N_2119);
xnor U3334 (N_3334,N_2167,N_2302);
and U3335 (N_3335,N_2964,N_2281);
nor U3336 (N_3336,N_2369,N_2908);
nand U3337 (N_3337,N_2810,N_2188);
nand U3338 (N_3338,N_2091,N_2398);
and U3339 (N_3339,N_2882,N_2930);
or U3340 (N_3340,N_2412,N_2229);
nand U3341 (N_3341,N_2642,N_2276);
nor U3342 (N_3342,N_2202,N_2484);
nand U3343 (N_3343,N_2356,N_2880);
nand U3344 (N_3344,N_2096,N_2802);
nor U3345 (N_3345,N_2825,N_2796);
nor U3346 (N_3346,N_2277,N_2004);
or U3347 (N_3347,N_2161,N_2044);
xnor U3348 (N_3348,N_2516,N_2027);
and U3349 (N_3349,N_2489,N_2193);
and U3350 (N_3350,N_2972,N_2006);
nor U3351 (N_3351,N_2698,N_2761);
or U3352 (N_3352,N_2662,N_2738);
nand U3353 (N_3353,N_2049,N_2525);
nor U3354 (N_3354,N_2621,N_2138);
nand U3355 (N_3355,N_2171,N_2888);
and U3356 (N_3356,N_2868,N_2268);
or U3357 (N_3357,N_2701,N_2114);
nor U3358 (N_3358,N_2064,N_2997);
or U3359 (N_3359,N_2311,N_2157);
nand U3360 (N_3360,N_2852,N_2380);
and U3361 (N_3361,N_2472,N_2891);
and U3362 (N_3362,N_2583,N_2541);
xnor U3363 (N_3363,N_2829,N_2128);
and U3364 (N_3364,N_2627,N_2308);
or U3365 (N_3365,N_2820,N_2726);
or U3366 (N_3366,N_2174,N_2658);
nand U3367 (N_3367,N_2447,N_2418);
xnor U3368 (N_3368,N_2631,N_2493);
nor U3369 (N_3369,N_2034,N_2661);
and U3370 (N_3370,N_2596,N_2991);
nor U3371 (N_3371,N_2104,N_2622);
and U3372 (N_3372,N_2857,N_2434);
nand U3373 (N_3373,N_2121,N_2358);
nor U3374 (N_3374,N_2998,N_2962);
nand U3375 (N_3375,N_2424,N_2550);
nand U3376 (N_3376,N_2691,N_2261);
and U3377 (N_3377,N_2070,N_2253);
nor U3378 (N_3378,N_2290,N_2900);
nor U3379 (N_3379,N_2057,N_2564);
nor U3380 (N_3380,N_2059,N_2505);
and U3381 (N_3381,N_2477,N_2403);
nor U3382 (N_3382,N_2690,N_2140);
nor U3383 (N_3383,N_2464,N_2574);
nor U3384 (N_3384,N_2865,N_2707);
and U3385 (N_3385,N_2507,N_2283);
or U3386 (N_3386,N_2107,N_2949);
or U3387 (N_3387,N_2142,N_2769);
nand U3388 (N_3388,N_2939,N_2220);
xnor U3389 (N_3389,N_2126,N_2578);
or U3390 (N_3390,N_2756,N_2118);
nor U3391 (N_3391,N_2586,N_2249);
nand U3392 (N_3392,N_2818,N_2824);
or U3393 (N_3393,N_2806,N_2914);
or U3394 (N_3394,N_2981,N_2515);
nor U3395 (N_3395,N_2471,N_2083);
or U3396 (N_3396,N_2366,N_2209);
nor U3397 (N_3397,N_2011,N_2406);
nand U3398 (N_3398,N_2431,N_2728);
and U3399 (N_3399,N_2321,N_2130);
and U3400 (N_3400,N_2045,N_2242);
nor U3401 (N_3401,N_2821,N_2191);
nor U3402 (N_3402,N_2218,N_2763);
nand U3403 (N_3403,N_2335,N_2937);
nand U3404 (N_3404,N_2577,N_2467);
or U3405 (N_3405,N_2674,N_2014);
or U3406 (N_3406,N_2987,N_2143);
nor U3407 (N_3407,N_2663,N_2259);
or U3408 (N_3408,N_2336,N_2942);
nor U3409 (N_3409,N_2773,N_2682);
and U3410 (N_3410,N_2643,N_2377);
or U3411 (N_3411,N_2792,N_2055);
xnor U3412 (N_3412,N_2705,N_2449);
or U3413 (N_3413,N_2620,N_2063);
xnor U3414 (N_3414,N_2819,N_2967);
nand U3415 (N_3415,N_2812,N_2323);
nand U3416 (N_3416,N_2787,N_2503);
xor U3417 (N_3417,N_2530,N_2894);
nand U3418 (N_3418,N_2496,N_2814);
and U3419 (N_3419,N_2901,N_2041);
xnor U3420 (N_3420,N_2735,N_2285);
nand U3421 (N_3421,N_2187,N_2848);
nand U3422 (N_3422,N_2502,N_2695);
nor U3423 (N_3423,N_2696,N_2755);
nand U3424 (N_3424,N_2073,N_2954);
nand U3425 (N_3425,N_2461,N_2085);
and U3426 (N_3426,N_2750,N_2711);
nor U3427 (N_3427,N_2474,N_2028);
nor U3428 (N_3428,N_2498,N_2851);
nor U3429 (N_3429,N_2941,N_2681);
nor U3430 (N_3430,N_2457,N_2481);
or U3431 (N_3431,N_2297,N_2847);
nand U3432 (N_3432,N_2599,N_2158);
or U3433 (N_3433,N_2223,N_2284);
or U3434 (N_3434,N_2475,N_2389);
nand U3435 (N_3435,N_2328,N_2625);
nand U3436 (N_3436,N_2017,N_2299);
and U3437 (N_3437,N_2236,N_2751);
nor U3438 (N_3438,N_2186,N_2247);
nor U3439 (N_3439,N_2785,N_2021);
or U3440 (N_3440,N_2985,N_2671);
or U3441 (N_3441,N_2689,N_2224);
nand U3442 (N_3442,N_2497,N_2303);
nor U3443 (N_3443,N_2078,N_2000);
and U3444 (N_3444,N_2965,N_2687);
nand U3445 (N_3445,N_2892,N_2638);
or U3446 (N_3446,N_2669,N_2741);
nor U3447 (N_3447,N_2534,N_2046);
nor U3448 (N_3448,N_2561,N_2394);
or U3449 (N_3449,N_2035,N_2613);
and U3450 (N_3450,N_2615,N_2304);
and U3451 (N_3451,N_2206,N_2296);
and U3452 (N_3452,N_2834,N_2710);
nor U3453 (N_3453,N_2428,N_2164);
and U3454 (N_3454,N_2742,N_2448);
and U3455 (N_3455,N_2680,N_2571);
or U3456 (N_3456,N_2733,N_2786);
and U3457 (N_3457,N_2838,N_2180);
or U3458 (N_3458,N_2732,N_2533);
and U3459 (N_3459,N_2018,N_2552);
or U3460 (N_3460,N_2861,N_2185);
or U3461 (N_3461,N_2318,N_2723);
or U3462 (N_3462,N_2101,N_2395);
nand U3463 (N_3463,N_2252,N_2612);
nor U3464 (N_3464,N_2685,N_2904);
or U3465 (N_3465,N_2801,N_2081);
nand U3466 (N_3466,N_2214,N_2542);
and U3467 (N_3467,N_2183,N_2033);
and U3468 (N_3468,N_2286,N_2040);
or U3469 (N_3469,N_2074,N_2155);
and U3470 (N_3470,N_2351,N_2195);
nor U3471 (N_3471,N_2346,N_2037);
nor U3472 (N_3472,N_2618,N_2453);
nand U3473 (N_3473,N_2789,N_2436);
nand U3474 (N_3474,N_2278,N_2677);
nor U3475 (N_3475,N_2451,N_2815);
nor U3476 (N_3476,N_2341,N_2549);
or U3477 (N_3477,N_2093,N_2274);
nor U3478 (N_3478,N_2537,N_2390);
and U3479 (N_3479,N_2103,N_2553);
nor U3480 (N_3480,N_2442,N_2342);
and U3481 (N_3481,N_2798,N_2529);
nor U3482 (N_3482,N_2184,N_2867);
nand U3483 (N_3483,N_2317,N_2198);
and U3484 (N_3484,N_2547,N_2923);
and U3485 (N_3485,N_2392,N_2635);
nor U3486 (N_3486,N_2975,N_2201);
xor U3487 (N_3487,N_2470,N_2731);
or U3488 (N_3488,N_2016,N_2354);
and U3489 (N_3489,N_2916,N_2885);
or U3490 (N_3490,N_2032,N_2955);
nor U3491 (N_3491,N_2476,N_2791);
or U3492 (N_3492,N_2713,N_2240);
and U3493 (N_3493,N_2301,N_2684);
nor U3494 (N_3494,N_2749,N_2066);
or U3495 (N_3495,N_2845,N_2853);
and U3496 (N_3496,N_2951,N_2344);
nand U3497 (N_3497,N_2992,N_2743);
nor U3498 (N_3498,N_2305,N_2859);
nand U3499 (N_3499,N_2012,N_2172);
and U3500 (N_3500,N_2003,N_2877);
or U3501 (N_3501,N_2403,N_2125);
nand U3502 (N_3502,N_2216,N_2782);
or U3503 (N_3503,N_2577,N_2448);
nor U3504 (N_3504,N_2462,N_2263);
and U3505 (N_3505,N_2447,N_2471);
nand U3506 (N_3506,N_2922,N_2294);
nand U3507 (N_3507,N_2725,N_2499);
and U3508 (N_3508,N_2411,N_2918);
nand U3509 (N_3509,N_2644,N_2923);
nor U3510 (N_3510,N_2460,N_2181);
or U3511 (N_3511,N_2548,N_2913);
and U3512 (N_3512,N_2028,N_2180);
nor U3513 (N_3513,N_2857,N_2155);
and U3514 (N_3514,N_2086,N_2492);
or U3515 (N_3515,N_2145,N_2520);
nand U3516 (N_3516,N_2237,N_2521);
xor U3517 (N_3517,N_2254,N_2410);
and U3518 (N_3518,N_2668,N_2187);
or U3519 (N_3519,N_2015,N_2128);
nor U3520 (N_3520,N_2368,N_2281);
or U3521 (N_3521,N_2838,N_2368);
xor U3522 (N_3522,N_2271,N_2137);
nor U3523 (N_3523,N_2178,N_2473);
and U3524 (N_3524,N_2495,N_2641);
nand U3525 (N_3525,N_2268,N_2297);
nor U3526 (N_3526,N_2308,N_2448);
nand U3527 (N_3527,N_2180,N_2287);
nor U3528 (N_3528,N_2340,N_2595);
nand U3529 (N_3529,N_2947,N_2634);
or U3530 (N_3530,N_2256,N_2581);
and U3531 (N_3531,N_2142,N_2751);
nor U3532 (N_3532,N_2316,N_2120);
or U3533 (N_3533,N_2404,N_2496);
or U3534 (N_3534,N_2708,N_2507);
nor U3535 (N_3535,N_2488,N_2074);
nor U3536 (N_3536,N_2815,N_2723);
nand U3537 (N_3537,N_2242,N_2350);
and U3538 (N_3538,N_2092,N_2064);
or U3539 (N_3539,N_2999,N_2546);
and U3540 (N_3540,N_2960,N_2406);
nor U3541 (N_3541,N_2429,N_2601);
and U3542 (N_3542,N_2853,N_2253);
nor U3543 (N_3543,N_2146,N_2530);
and U3544 (N_3544,N_2013,N_2542);
nand U3545 (N_3545,N_2542,N_2202);
nor U3546 (N_3546,N_2423,N_2750);
nor U3547 (N_3547,N_2975,N_2487);
xnor U3548 (N_3548,N_2195,N_2597);
or U3549 (N_3549,N_2774,N_2725);
nor U3550 (N_3550,N_2240,N_2660);
and U3551 (N_3551,N_2673,N_2397);
and U3552 (N_3552,N_2672,N_2404);
nor U3553 (N_3553,N_2562,N_2989);
and U3554 (N_3554,N_2567,N_2680);
and U3555 (N_3555,N_2392,N_2752);
and U3556 (N_3556,N_2287,N_2516);
or U3557 (N_3557,N_2727,N_2405);
xor U3558 (N_3558,N_2165,N_2573);
and U3559 (N_3559,N_2480,N_2552);
nand U3560 (N_3560,N_2853,N_2448);
nand U3561 (N_3561,N_2162,N_2349);
nor U3562 (N_3562,N_2504,N_2327);
and U3563 (N_3563,N_2358,N_2430);
nor U3564 (N_3564,N_2591,N_2735);
nor U3565 (N_3565,N_2205,N_2985);
nor U3566 (N_3566,N_2196,N_2487);
nand U3567 (N_3567,N_2078,N_2438);
nor U3568 (N_3568,N_2912,N_2791);
nand U3569 (N_3569,N_2693,N_2667);
nand U3570 (N_3570,N_2387,N_2160);
nor U3571 (N_3571,N_2542,N_2824);
nor U3572 (N_3572,N_2425,N_2964);
nor U3573 (N_3573,N_2537,N_2508);
and U3574 (N_3574,N_2895,N_2693);
nand U3575 (N_3575,N_2412,N_2686);
and U3576 (N_3576,N_2058,N_2675);
nand U3577 (N_3577,N_2377,N_2177);
and U3578 (N_3578,N_2943,N_2070);
nor U3579 (N_3579,N_2128,N_2696);
nand U3580 (N_3580,N_2301,N_2049);
and U3581 (N_3581,N_2411,N_2785);
or U3582 (N_3582,N_2731,N_2193);
and U3583 (N_3583,N_2716,N_2824);
nor U3584 (N_3584,N_2494,N_2674);
or U3585 (N_3585,N_2405,N_2842);
or U3586 (N_3586,N_2292,N_2373);
or U3587 (N_3587,N_2262,N_2044);
and U3588 (N_3588,N_2202,N_2143);
nor U3589 (N_3589,N_2476,N_2688);
and U3590 (N_3590,N_2775,N_2376);
nand U3591 (N_3591,N_2675,N_2630);
and U3592 (N_3592,N_2625,N_2455);
or U3593 (N_3593,N_2615,N_2575);
or U3594 (N_3594,N_2467,N_2963);
and U3595 (N_3595,N_2485,N_2937);
or U3596 (N_3596,N_2767,N_2505);
or U3597 (N_3597,N_2191,N_2294);
nand U3598 (N_3598,N_2851,N_2260);
or U3599 (N_3599,N_2248,N_2216);
nand U3600 (N_3600,N_2567,N_2181);
nor U3601 (N_3601,N_2990,N_2851);
nor U3602 (N_3602,N_2323,N_2760);
nand U3603 (N_3603,N_2078,N_2952);
or U3604 (N_3604,N_2943,N_2815);
nand U3605 (N_3605,N_2327,N_2059);
or U3606 (N_3606,N_2045,N_2382);
or U3607 (N_3607,N_2308,N_2136);
nand U3608 (N_3608,N_2174,N_2154);
nor U3609 (N_3609,N_2787,N_2133);
nand U3610 (N_3610,N_2267,N_2925);
or U3611 (N_3611,N_2879,N_2455);
nor U3612 (N_3612,N_2488,N_2012);
nor U3613 (N_3613,N_2516,N_2974);
xnor U3614 (N_3614,N_2018,N_2410);
nand U3615 (N_3615,N_2215,N_2104);
nand U3616 (N_3616,N_2815,N_2953);
nor U3617 (N_3617,N_2099,N_2062);
and U3618 (N_3618,N_2656,N_2453);
or U3619 (N_3619,N_2151,N_2182);
or U3620 (N_3620,N_2975,N_2157);
xnor U3621 (N_3621,N_2362,N_2354);
or U3622 (N_3622,N_2339,N_2586);
and U3623 (N_3623,N_2723,N_2983);
nand U3624 (N_3624,N_2397,N_2487);
and U3625 (N_3625,N_2904,N_2772);
nand U3626 (N_3626,N_2890,N_2707);
or U3627 (N_3627,N_2207,N_2257);
or U3628 (N_3628,N_2413,N_2295);
and U3629 (N_3629,N_2148,N_2938);
nand U3630 (N_3630,N_2035,N_2686);
nand U3631 (N_3631,N_2453,N_2063);
nor U3632 (N_3632,N_2468,N_2301);
nand U3633 (N_3633,N_2806,N_2736);
and U3634 (N_3634,N_2427,N_2202);
and U3635 (N_3635,N_2941,N_2334);
nor U3636 (N_3636,N_2171,N_2419);
nand U3637 (N_3637,N_2312,N_2176);
nor U3638 (N_3638,N_2772,N_2631);
and U3639 (N_3639,N_2159,N_2422);
or U3640 (N_3640,N_2371,N_2551);
nand U3641 (N_3641,N_2386,N_2432);
nor U3642 (N_3642,N_2735,N_2458);
and U3643 (N_3643,N_2066,N_2318);
nand U3644 (N_3644,N_2503,N_2619);
nand U3645 (N_3645,N_2786,N_2811);
and U3646 (N_3646,N_2718,N_2283);
or U3647 (N_3647,N_2524,N_2709);
and U3648 (N_3648,N_2188,N_2842);
nor U3649 (N_3649,N_2833,N_2403);
nand U3650 (N_3650,N_2134,N_2249);
nor U3651 (N_3651,N_2446,N_2920);
nor U3652 (N_3652,N_2343,N_2383);
and U3653 (N_3653,N_2003,N_2472);
nand U3654 (N_3654,N_2985,N_2274);
xnor U3655 (N_3655,N_2164,N_2909);
nand U3656 (N_3656,N_2224,N_2324);
or U3657 (N_3657,N_2765,N_2964);
nor U3658 (N_3658,N_2247,N_2700);
nand U3659 (N_3659,N_2243,N_2612);
and U3660 (N_3660,N_2651,N_2553);
or U3661 (N_3661,N_2491,N_2294);
or U3662 (N_3662,N_2777,N_2194);
nor U3663 (N_3663,N_2316,N_2447);
and U3664 (N_3664,N_2062,N_2055);
nand U3665 (N_3665,N_2384,N_2041);
or U3666 (N_3666,N_2512,N_2834);
and U3667 (N_3667,N_2160,N_2580);
nor U3668 (N_3668,N_2491,N_2447);
nor U3669 (N_3669,N_2961,N_2351);
nand U3670 (N_3670,N_2075,N_2292);
nor U3671 (N_3671,N_2024,N_2390);
nor U3672 (N_3672,N_2669,N_2256);
nand U3673 (N_3673,N_2458,N_2893);
xnor U3674 (N_3674,N_2205,N_2242);
and U3675 (N_3675,N_2757,N_2114);
xnor U3676 (N_3676,N_2010,N_2233);
and U3677 (N_3677,N_2824,N_2258);
nand U3678 (N_3678,N_2457,N_2070);
nor U3679 (N_3679,N_2937,N_2216);
or U3680 (N_3680,N_2970,N_2078);
nor U3681 (N_3681,N_2698,N_2550);
nor U3682 (N_3682,N_2421,N_2346);
nand U3683 (N_3683,N_2417,N_2449);
nand U3684 (N_3684,N_2271,N_2953);
and U3685 (N_3685,N_2165,N_2121);
and U3686 (N_3686,N_2442,N_2511);
or U3687 (N_3687,N_2904,N_2566);
nand U3688 (N_3688,N_2800,N_2152);
and U3689 (N_3689,N_2797,N_2288);
or U3690 (N_3690,N_2913,N_2857);
nor U3691 (N_3691,N_2715,N_2481);
or U3692 (N_3692,N_2479,N_2314);
and U3693 (N_3693,N_2431,N_2392);
and U3694 (N_3694,N_2239,N_2060);
and U3695 (N_3695,N_2905,N_2201);
and U3696 (N_3696,N_2594,N_2423);
nand U3697 (N_3697,N_2737,N_2575);
nor U3698 (N_3698,N_2281,N_2287);
and U3699 (N_3699,N_2299,N_2933);
nand U3700 (N_3700,N_2517,N_2774);
and U3701 (N_3701,N_2221,N_2683);
and U3702 (N_3702,N_2349,N_2342);
and U3703 (N_3703,N_2749,N_2886);
or U3704 (N_3704,N_2916,N_2408);
and U3705 (N_3705,N_2477,N_2884);
or U3706 (N_3706,N_2937,N_2729);
nor U3707 (N_3707,N_2267,N_2579);
or U3708 (N_3708,N_2505,N_2711);
or U3709 (N_3709,N_2220,N_2326);
nor U3710 (N_3710,N_2755,N_2797);
nor U3711 (N_3711,N_2843,N_2281);
nand U3712 (N_3712,N_2964,N_2360);
nor U3713 (N_3713,N_2458,N_2581);
or U3714 (N_3714,N_2184,N_2974);
nand U3715 (N_3715,N_2178,N_2361);
nand U3716 (N_3716,N_2171,N_2173);
nor U3717 (N_3717,N_2454,N_2266);
nand U3718 (N_3718,N_2516,N_2682);
or U3719 (N_3719,N_2642,N_2998);
and U3720 (N_3720,N_2890,N_2515);
nor U3721 (N_3721,N_2488,N_2356);
or U3722 (N_3722,N_2888,N_2221);
nor U3723 (N_3723,N_2586,N_2014);
nor U3724 (N_3724,N_2019,N_2964);
and U3725 (N_3725,N_2980,N_2061);
nor U3726 (N_3726,N_2841,N_2469);
and U3727 (N_3727,N_2595,N_2451);
nor U3728 (N_3728,N_2043,N_2719);
and U3729 (N_3729,N_2704,N_2244);
and U3730 (N_3730,N_2733,N_2625);
nor U3731 (N_3731,N_2821,N_2333);
and U3732 (N_3732,N_2000,N_2090);
and U3733 (N_3733,N_2865,N_2444);
nand U3734 (N_3734,N_2697,N_2960);
nand U3735 (N_3735,N_2107,N_2064);
nand U3736 (N_3736,N_2805,N_2122);
or U3737 (N_3737,N_2064,N_2534);
and U3738 (N_3738,N_2203,N_2128);
and U3739 (N_3739,N_2374,N_2118);
nor U3740 (N_3740,N_2180,N_2899);
and U3741 (N_3741,N_2827,N_2948);
and U3742 (N_3742,N_2919,N_2336);
or U3743 (N_3743,N_2516,N_2450);
nand U3744 (N_3744,N_2890,N_2094);
nor U3745 (N_3745,N_2679,N_2030);
nor U3746 (N_3746,N_2910,N_2331);
or U3747 (N_3747,N_2894,N_2494);
nand U3748 (N_3748,N_2395,N_2585);
or U3749 (N_3749,N_2742,N_2287);
xnor U3750 (N_3750,N_2120,N_2820);
or U3751 (N_3751,N_2725,N_2039);
and U3752 (N_3752,N_2714,N_2402);
nand U3753 (N_3753,N_2884,N_2736);
or U3754 (N_3754,N_2454,N_2979);
or U3755 (N_3755,N_2404,N_2377);
xor U3756 (N_3756,N_2292,N_2011);
nand U3757 (N_3757,N_2732,N_2814);
nand U3758 (N_3758,N_2894,N_2681);
or U3759 (N_3759,N_2335,N_2704);
and U3760 (N_3760,N_2524,N_2909);
nor U3761 (N_3761,N_2586,N_2191);
nand U3762 (N_3762,N_2735,N_2551);
and U3763 (N_3763,N_2441,N_2606);
nand U3764 (N_3764,N_2921,N_2454);
or U3765 (N_3765,N_2528,N_2385);
or U3766 (N_3766,N_2606,N_2558);
nor U3767 (N_3767,N_2859,N_2932);
nor U3768 (N_3768,N_2669,N_2487);
nand U3769 (N_3769,N_2837,N_2639);
nor U3770 (N_3770,N_2952,N_2625);
nand U3771 (N_3771,N_2140,N_2854);
nor U3772 (N_3772,N_2563,N_2900);
or U3773 (N_3773,N_2135,N_2633);
nor U3774 (N_3774,N_2527,N_2100);
nand U3775 (N_3775,N_2689,N_2377);
or U3776 (N_3776,N_2560,N_2294);
or U3777 (N_3777,N_2589,N_2262);
or U3778 (N_3778,N_2587,N_2887);
and U3779 (N_3779,N_2734,N_2367);
or U3780 (N_3780,N_2670,N_2338);
xnor U3781 (N_3781,N_2894,N_2686);
or U3782 (N_3782,N_2318,N_2885);
or U3783 (N_3783,N_2230,N_2715);
or U3784 (N_3784,N_2313,N_2801);
nand U3785 (N_3785,N_2019,N_2359);
nand U3786 (N_3786,N_2169,N_2288);
and U3787 (N_3787,N_2847,N_2987);
nand U3788 (N_3788,N_2232,N_2887);
nor U3789 (N_3789,N_2525,N_2397);
and U3790 (N_3790,N_2481,N_2942);
and U3791 (N_3791,N_2783,N_2564);
nor U3792 (N_3792,N_2569,N_2533);
nor U3793 (N_3793,N_2912,N_2661);
or U3794 (N_3794,N_2080,N_2697);
xor U3795 (N_3795,N_2170,N_2285);
or U3796 (N_3796,N_2421,N_2127);
nand U3797 (N_3797,N_2592,N_2446);
xor U3798 (N_3798,N_2182,N_2525);
nand U3799 (N_3799,N_2809,N_2047);
nand U3800 (N_3800,N_2881,N_2096);
or U3801 (N_3801,N_2699,N_2548);
nor U3802 (N_3802,N_2633,N_2206);
and U3803 (N_3803,N_2307,N_2811);
nor U3804 (N_3804,N_2693,N_2584);
nor U3805 (N_3805,N_2611,N_2392);
nand U3806 (N_3806,N_2143,N_2927);
nor U3807 (N_3807,N_2017,N_2169);
nor U3808 (N_3808,N_2972,N_2733);
and U3809 (N_3809,N_2642,N_2886);
xnor U3810 (N_3810,N_2175,N_2162);
and U3811 (N_3811,N_2531,N_2684);
nand U3812 (N_3812,N_2889,N_2149);
nor U3813 (N_3813,N_2035,N_2869);
nor U3814 (N_3814,N_2869,N_2256);
nor U3815 (N_3815,N_2698,N_2764);
or U3816 (N_3816,N_2087,N_2111);
nor U3817 (N_3817,N_2407,N_2527);
or U3818 (N_3818,N_2726,N_2535);
nor U3819 (N_3819,N_2527,N_2006);
nand U3820 (N_3820,N_2525,N_2611);
xnor U3821 (N_3821,N_2323,N_2952);
nor U3822 (N_3822,N_2269,N_2666);
nand U3823 (N_3823,N_2414,N_2070);
nor U3824 (N_3824,N_2511,N_2152);
or U3825 (N_3825,N_2283,N_2697);
or U3826 (N_3826,N_2689,N_2854);
and U3827 (N_3827,N_2863,N_2511);
nand U3828 (N_3828,N_2153,N_2593);
or U3829 (N_3829,N_2525,N_2474);
or U3830 (N_3830,N_2981,N_2620);
and U3831 (N_3831,N_2978,N_2204);
and U3832 (N_3832,N_2910,N_2199);
or U3833 (N_3833,N_2140,N_2068);
or U3834 (N_3834,N_2103,N_2803);
nor U3835 (N_3835,N_2425,N_2765);
nand U3836 (N_3836,N_2867,N_2716);
nand U3837 (N_3837,N_2721,N_2032);
nor U3838 (N_3838,N_2374,N_2519);
nor U3839 (N_3839,N_2296,N_2271);
and U3840 (N_3840,N_2541,N_2693);
and U3841 (N_3841,N_2734,N_2713);
xnor U3842 (N_3842,N_2791,N_2245);
nor U3843 (N_3843,N_2745,N_2826);
and U3844 (N_3844,N_2988,N_2453);
xnor U3845 (N_3845,N_2083,N_2791);
or U3846 (N_3846,N_2613,N_2891);
and U3847 (N_3847,N_2949,N_2583);
nand U3848 (N_3848,N_2680,N_2206);
or U3849 (N_3849,N_2132,N_2242);
and U3850 (N_3850,N_2973,N_2304);
or U3851 (N_3851,N_2265,N_2574);
or U3852 (N_3852,N_2361,N_2414);
and U3853 (N_3853,N_2540,N_2604);
nor U3854 (N_3854,N_2025,N_2275);
or U3855 (N_3855,N_2103,N_2365);
nand U3856 (N_3856,N_2073,N_2423);
or U3857 (N_3857,N_2739,N_2978);
and U3858 (N_3858,N_2787,N_2650);
and U3859 (N_3859,N_2250,N_2133);
or U3860 (N_3860,N_2268,N_2432);
nand U3861 (N_3861,N_2085,N_2449);
nor U3862 (N_3862,N_2865,N_2073);
and U3863 (N_3863,N_2398,N_2343);
nor U3864 (N_3864,N_2842,N_2290);
nand U3865 (N_3865,N_2240,N_2181);
nor U3866 (N_3866,N_2215,N_2437);
nor U3867 (N_3867,N_2138,N_2243);
nor U3868 (N_3868,N_2114,N_2957);
nand U3869 (N_3869,N_2227,N_2708);
and U3870 (N_3870,N_2731,N_2547);
and U3871 (N_3871,N_2919,N_2564);
nand U3872 (N_3872,N_2279,N_2113);
nor U3873 (N_3873,N_2594,N_2360);
nand U3874 (N_3874,N_2913,N_2352);
xnor U3875 (N_3875,N_2102,N_2707);
and U3876 (N_3876,N_2538,N_2026);
nand U3877 (N_3877,N_2259,N_2714);
nor U3878 (N_3878,N_2527,N_2147);
and U3879 (N_3879,N_2652,N_2735);
or U3880 (N_3880,N_2615,N_2889);
nand U3881 (N_3881,N_2118,N_2110);
nand U3882 (N_3882,N_2362,N_2946);
or U3883 (N_3883,N_2121,N_2697);
and U3884 (N_3884,N_2015,N_2085);
nand U3885 (N_3885,N_2768,N_2163);
and U3886 (N_3886,N_2968,N_2641);
nor U3887 (N_3887,N_2769,N_2346);
nor U3888 (N_3888,N_2462,N_2858);
nand U3889 (N_3889,N_2120,N_2661);
nor U3890 (N_3890,N_2629,N_2335);
and U3891 (N_3891,N_2626,N_2579);
nand U3892 (N_3892,N_2353,N_2235);
and U3893 (N_3893,N_2975,N_2686);
and U3894 (N_3894,N_2513,N_2674);
and U3895 (N_3895,N_2180,N_2692);
nand U3896 (N_3896,N_2585,N_2189);
nand U3897 (N_3897,N_2127,N_2333);
or U3898 (N_3898,N_2691,N_2584);
or U3899 (N_3899,N_2495,N_2691);
nor U3900 (N_3900,N_2793,N_2261);
nor U3901 (N_3901,N_2701,N_2238);
nand U3902 (N_3902,N_2328,N_2520);
nor U3903 (N_3903,N_2079,N_2706);
or U3904 (N_3904,N_2674,N_2990);
or U3905 (N_3905,N_2104,N_2639);
nor U3906 (N_3906,N_2028,N_2458);
or U3907 (N_3907,N_2999,N_2860);
or U3908 (N_3908,N_2420,N_2482);
and U3909 (N_3909,N_2142,N_2430);
nand U3910 (N_3910,N_2020,N_2420);
xnor U3911 (N_3911,N_2482,N_2556);
nand U3912 (N_3912,N_2303,N_2387);
or U3913 (N_3913,N_2030,N_2330);
and U3914 (N_3914,N_2172,N_2744);
nor U3915 (N_3915,N_2958,N_2830);
nor U3916 (N_3916,N_2018,N_2654);
and U3917 (N_3917,N_2488,N_2665);
or U3918 (N_3918,N_2007,N_2635);
nand U3919 (N_3919,N_2694,N_2213);
nand U3920 (N_3920,N_2406,N_2804);
xnor U3921 (N_3921,N_2641,N_2570);
and U3922 (N_3922,N_2221,N_2789);
nor U3923 (N_3923,N_2913,N_2329);
nor U3924 (N_3924,N_2663,N_2166);
xnor U3925 (N_3925,N_2065,N_2102);
and U3926 (N_3926,N_2162,N_2384);
and U3927 (N_3927,N_2443,N_2514);
or U3928 (N_3928,N_2597,N_2407);
xor U3929 (N_3929,N_2800,N_2597);
xnor U3930 (N_3930,N_2509,N_2792);
nand U3931 (N_3931,N_2450,N_2578);
nor U3932 (N_3932,N_2813,N_2504);
and U3933 (N_3933,N_2319,N_2441);
nand U3934 (N_3934,N_2295,N_2859);
nor U3935 (N_3935,N_2749,N_2228);
nor U3936 (N_3936,N_2908,N_2440);
or U3937 (N_3937,N_2795,N_2050);
nor U3938 (N_3938,N_2964,N_2653);
nand U3939 (N_3939,N_2506,N_2550);
and U3940 (N_3940,N_2609,N_2734);
nor U3941 (N_3941,N_2339,N_2489);
and U3942 (N_3942,N_2520,N_2312);
and U3943 (N_3943,N_2027,N_2687);
or U3944 (N_3944,N_2212,N_2207);
or U3945 (N_3945,N_2379,N_2873);
or U3946 (N_3946,N_2649,N_2260);
or U3947 (N_3947,N_2391,N_2916);
nand U3948 (N_3948,N_2735,N_2679);
nand U3949 (N_3949,N_2114,N_2873);
and U3950 (N_3950,N_2509,N_2037);
xor U3951 (N_3951,N_2042,N_2946);
nor U3952 (N_3952,N_2573,N_2667);
and U3953 (N_3953,N_2551,N_2323);
nor U3954 (N_3954,N_2024,N_2055);
nand U3955 (N_3955,N_2822,N_2730);
nor U3956 (N_3956,N_2717,N_2870);
and U3957 (N_3957,N_2049,N_2371);
nand U3958 (N_3958,N_2886,N_2018);
nor U3959 (N_3959,N_2651,N_2980);
nand U3960 (N_3960,N_2042,N_2948);
or U3961 (N_3961,N_2450,N_2289);
xor U3962 (N_3962,N_2301,N_2484);
and U3963 (N_3963,N_2700,N_2305);
nand U3964 (N_3964,N_2882,N_2762);
xor U3965 (N_3965,N_2767,N_2990);
nand U3966 (N_3966,N_2582,N_2816);
xor U3967 (N_3967,N_2428,N_2322);
and U3968 (N_3968,N_2399,N_2522);
and U3969 (N_3969,N_2033,N_2358);
and U3970 (N_3970,N_2819,N_2552);
nand U3971 (N_3971,N_2246,N_2709);
nor U3972 (N_3972,N_2115,N_2891);
nor U3973 (N_3973,N_2817,N_2973);
or U3974 (N_3974,N_2483,N_2406);
nor U3975 (N_3975,N_2020,N_2533);
and U3976 (N_3976,N_2196,N_2111);
nand U3977 (N_3977,N_2203,N_2903);
nand U3978 (N_3978,N_2786,N_2382);
nor U3979 (N_3979,N_2379,N_2623);
and U3980 (N_3980,N_2185,N_2559);
or U3981 (N_3981,N_2029,N_2124);
nor U3982 (N_3982,N_2774,N_2205);
nor U3983 (N_3983,N_2882,N_2943);
nand U3984 (N_3984,N_2791,N_2007);
nor U3985 (N_3985,N_2915,N_2012);
and U3986 (N_3986,N_2906,N_2617);
or U3987 (N_3987,N_2237,N_2310);
and U3988 (N_3988,N_2484,N_2528);
and U3989 (N_3989,N_2105,N_2404);
nor U3990 (N_3990,N_2672,N_2482);
nand U3991 (N_3991,N_2375,N_2470);
and U3992 (N_3992,N_2214,N_2963);
and U3993 (N_3993,N_2798,N_2386);
nand U3994 (N_3994,N_2602,N_2654);
nand U3995 (N_3995,N_2557,N_2491);
and U3996 (N_3996,N_2966,N_2398);
or U3997 (N_3997,N_2510,N_2685);
and U3998 (N_3998,N_2274,N_2795);
nand U3999 (N_3999,N_2552,N_2131);
nor U4000 (N_4000,N_3178,N_3899);
or U4001 (N_4001,N_3932,N_3030);
or U4002 (N_4002,N_3065,N_3621);
nand U4003 (N_4003,N_3715,N_3979);
and U4004 (N_4004,N_3000,N_3414);
xor U4005 (N_4005,N_3796,N_3909);
and U4006 (N_4006,N_3207,N_3338);
or U4007 (N_4007,N_3163,N_3679);
nor U4008 (N_4008,N_3772,N_3939);
nand U4009 (N_4009,N_3795,N_3437);
or U4010 (N_4010,N_3730,N_3934);
and U4011 (N_4011,N_3937,N_3217);
and U4012 (N_4012,N_3131,N_3229);
or U4013 (N_4013,N_3494,N_3972);
or U4014 (N_4014,N_3875,N_3631);
nor U4015 (N_4015,N_3317,N_3246);
xnor U4016 (N_4016,N_3641,N_3614);
and U4017 (N_4017,N_3304,N_3223);
or U4018 (N_4018,N_3133,N_3467);
nor U4019 (N_4019,N_3056,N_3770);
xor U4020 (N_4020,N_3023,N_3896);
and U4021 (N_4021,N_3142,N_3067);
nor U4022 (N_4022,N_3855,N_3719);
and U4023 (N_4023,N_3793,N_3590);
nor U4024 (N_4024,N_3747,N_3559);
and U4025 (N_4025,N_3263,N_3589);
nand U4026 (N_4026,N_3552,N_3819);
nor U4027 (N_4027,N_3418,N_3569);
and U4028 (N_4028,N_3814,N_3813);
or U4029 (N_4029,N_3232,N_3392);
and U4030 (N_4030,N_3769,N_3202);
or U4031 (N_4031,N_3327,N_3568);
nor U4032 (N_4032,N_3637,N_3535);
or U4033 (N_4033,N_3493,N_3702);
or U4034 (N_4034,N_3235,N_3827);
nand U4035 (N_4035,N_3090,N_3815);
and U4036 (N_4036,N_3732,N_3809);
and U4037 (N_4037,N_3143,N_3300);
nor U4038 (N_4038,N_3593,N_3196);
and U4039 (N_4039,N_3149,N_3186);
and U4040 (N_4040,N_3669,N_3474);
nor U4041 (N_4041,N_3760,N_3876);
nor U4042 (N_4042,N_3975,N_3335);
and U4043 (N_4043,N_3581,N_3288);
and U4044 (N_4044,N_3870,N_3596);
and U4045 (N_4045,N_3943,N_3530);
and U4046 (N_4046,N_3622,N_3703);
nand U4047 (N_4047,N_3778,N_3215);
nand U4048 (N_4048,N_3691,N_3643);
nor U4049 (N_4049,N_3430,N_3992);
and U4050 (N_4050,N_3851,N_3499);
xor U4051 (N_4051,N_3836,N_3678);
nand U4052 (N_4052,N_3100,N_3889);
nand U4053 (N_4053,N_3856,N_3918);
nand U4054 (N_4054,N_3973,N_3490);
or U4055 (N_4055,N_3960,N_3152);
or U4056 (N_4056,N_3313,N_3192);
nor U4057 (N_4057,N_3160,N_3237);
xor U4058 (N_4058,N_3865,N_3952);
nor U4059 (N_4059,N_3005,N_3157);
and U4060 (N_4060,N_3253,N_3954);
or U4061 (N_4061,N_3416,N_3483);
nand U4062 (N_4062,N_3510,N_3228);
nor U4063 (N_4063,N_3900,N_3123);
or U4064 (N_4064,N_3653,N_3113);
or U4065 (N_4065,N_3132,N_3907);
nand U4066 (N_4066,N_3256,N_3517);
nor U4067 (N_4067,N_3551,N_3226);
nand U4068 (N_4068,N_3367,N_3096);
nor U4069 (N_4069,N_3369,N_3694);
nor U4070 (N_4070,N_3503,N_3574);
or U4071 (N_4071,N_3656,N_3766);
and U4072 (N_4072,N_3261,N_3696);
nor U4073 (N_4073,N_3060,N_3931);
nand U4074 (N_4074,N_3233,N_3668);
or U4075 (N_4075,N_3633,N_3013);
or U4076 (N_4076,N_3828,N_3540);
nor U4077 (N_4077,N_3842,N_3049);
nor U4078 (N_4078,N_3484,N_3071);
nor U4079 (N_4079,N_3447,N_3911);
nor U4080 (N_4080,N_3555,N_3472);
or U4081 (N_4081,N_3441,N_3455);
nor U4082 (N_4082,N_3940,N_3359);
nand U4083 (N_4083,N_3420,N_3741);
and U4084 (N_4084,N_3829,N_3846);
nand U4085 (N_4085,N_3761,N_3941);
or U4086 (N_4086,N_3356,N_3533);
or U4087 (N_4087,N_3029,N_3158);
or U4088 (N_4088,N_3379,N_3570);
nand U4089 (N_4089,N_3734,N_3166);
and U4090 (N_4090,N_3404,N_3859);
xor U4091 (N_4091,N_3337,N_3565);
nor U4092 (N_4092,N_3128,N_3269);
nand U4093 (N_4093,N_3955,N_3879);
or U4094 (N_4094,N_3638,N_3212);
nor U4095 (N_4095,N_3334,N_3620);
and U4096 (N_4096,N_3145,N_3150);
nand U4097 (N_4097,N_3002,N_3475);
nand U4098 (N_4098,N_3273,N_3124);
and U4099 (N_4099,N_3477,N_3936);
and U4100 (N_4100,N_3452,N_3072);
xor U4101 (N_4101,N_3713,N_3785);
nor U4102 (N_4102,N_3588,N_3466);
and U4103 (N_4103,N_3117,N_3343);
nor U4104 (N_4104,N_3767,N_3083);
nand U4105 (N_4105,N_3436,N_3502);
or U4106 (N_4106,N_3308,N_3504);
and U4107 (N_4107,N_3399,N_3492);
nor U4108 (N_4108,N_3208,N_3890);
nand U4109 (N_4109,N_3986,N_3670);
and U4110 (N_4110,N_3582,N_3381);
or U4111 (N_4111,N_3010,N_3634);
nor U4112 (N_4112,N_3409,N_3244);
and U4113 (N_4113,N_3262,N_3898);
or U4114 (N_4114,N_3460,N_3573);
nor U4115 (N_4115,N_3744,N_3545);
and U4116 (N_4116,N_3947,N_3561);
or U4117 (N_4117,N_3413,N_3473);
or U4118 (N_4118,N_3440,N_3996);
or U4119 (N_4119,N_3024,N_3649);
and U4120 (N_4120,N_3594,N_3443);
and U4121 (N_4121,N_3843,N_3862);
or U4122 (N_4122,N_3675,N_3967);
nor U4123 (N_4123,N_3182,N_3560);
nand U4124 (N_4124,N_3372,N_3821);
nand U4125 (N_4125,N_3945,N_3924);
nand U4126 (N_4126,N_3915,N_3839);
nor U4127 (N_4127,N_3841,N_3958);
and U4128 (N_4128,N_3286,N_3365);
or U4129 (N_4129,N_3174,N_3425);
or U4130 (N_4130,N_3004,N_3615);
nor U4131 (N_4131,N_3177,N_3252);
nor U4132 (N_4132,N_3609,N_3930);
and U4133 (N_4133,N_3092,N_3506);
and U4134 (N_4134,N_3251,N_3305);
nand U4135 (N_4135,N_3651,N_3347);
nand U4136 (N_4136,N_3961,N_3274);
nor U4137 (N_4137,N_3738,N_3726);
nand U4138 (N_4138,N_3716,N_3435);
nand U4139 (N_4139,N_3642,N_3240);
nor U4140 (N_4140,N_3611,N_3984);
nand U4141 (N_4141,N_3156,N_3037);
xnor U4142 (N_4142,N_3904,N_3102);
and U4143 (N_4143,N_3751,N_3033);
nand U4144 (N_4144,N_3923,N_3957);
or U4145 (N_4145,N_3429,N_3861);
or U4146 (N_4146,N_3784,N_3844);
nand U4147 (N_4147,N_3897,N_3075);
and U4148 (N_4148,N_3108,N_3978);
or U4149 (N_4149,N_3401,N_3777);
nand U4150 (N_4150,N_3797,N_3242);
or U4151 (N_4151,N_3737,N_3189);
or U4152 (N_4152,N_3034,N_3042);
nor U4153 (N_4153,N_3717,N_3028);
and U4154 (N_4154,N_3185,N_3360);
nor U4155 (N_4155,N_3362,N_3640);
or U4156 (N_4156,N_3892,N_3116);
and U4157 (N_4157,N_3903,N_3025);
nor U4158 (N_4158,N_3981,N_3558);
nand U4159 (N_4159,N_3771,N_3358);
or U4160 (N_4160,N_3564,N_3151);
nand U4161 (N_4161,N_3074,N_3197);
and U4162 (N_4162,N_3866,N_3276);
nor U4163 (N_4163,N_3720,N_3688);
nand U4164 (N_4164,N_3199,N_3345);
nor U4165 (N_4165,N_3194,N_3488);
and U4166 (N_4166,N_3598,N_3364);
or U4167 (N_4167,N_3714,N_3684);
nor U4168 (N_4168,N_3431,N_3370);
nor U4169 (N_4169,N_3674,N_3051);
nand U4170 (N_4170,N_3059,N_3549);
nand U4171 (N_4171,N_3439,N_3134);
and U4172 (N_4172,N_3883,N_3585);
or U4173 (N_4173,N_3445,N_3683);
nand U4174 (N_4174,N_3699,N_3873);
or U4175 (N_4175,N_3781,N_3706);
or U4176 (N_4176,N_3983,N_3032);
nor U4177 (N_4177,N_3129,N_3512);
nand U4178 (N_4178,N_3712,N_3069);
and U4179 (N_4179,N_3442,N_3292);
or U4180 (N_4180,N_3114,N_3001);
nand U4181 (N_4181,N_3799,N_3933);
and U4182 (N_4182,N_3718,N_3045);
nor U4183 (N_4183,N_3571,N_3057);
and U4184 (N_4184,N_3677,N_3221);
and U4185 (N_4185,N_3661,N_3135);
nand U4186 (N_4186,N_3423,N_3200);
and U4187 (N_4187,N_3608,N_3491);
or U4188 (N_4188,N_3127,N_3301);
nand U4189 (N_4189,N_3881,N_3736);
nand U4190 (N_4190,N_3852,N_3099);
nand U4191 (N_4191,N_3184,N_3657);
and U4192 (N_4192,N_3547,N_3011);
nor U4193 (N_4193,N_3016,N_3204);
nor U4194 (N_4194,N_3154,N_3600);
or U4195 (N_4195,N_3709,N_3603);
nor U4196 (N_4196,N_3146,N_3377);
nor U4197 (N_4197,N_3068,N_3525);
nand U4198 (N_4198,N_3735,N_3800);
nand U4199 (N_4199,N_3155,N_3104);
nor U4200 (N_4200,N_3554,N_3449);
or U4201 (N_4201,N_3780,N_3407);
nand U4202 (N_4202,N_3085,N_3239);
nand U4203 (N_4203,N_3697,N_3398);
and U4204 (N_4204,N_3518,N_3816);
nand U4205 (N_4205,N_3648,N_3058);
nor U4206 (N_4206,N_3991,N_3309);
nor U4207 (N_4207,N_3970,N_3089);
or U4208 (N_4208,N_3205,N_3371);
or U4209 (N_4209,N_3721,N_3663);
nand U4210 (N_4210,N_3774,N_3311);
and U4211 (N_4211,N_3987,N_3121);
or U4212 (N_4212,N_3055,N_3480);
nor U4213 (N_4213,N_3976,N_3066);
or U4214 (N_4214,N_3927,N_3546);
nor U4215 (N_4215,N_3378,N_3776);
nor U4216 (N_4216,N_3832,N_3461);
nand U4217 (N_4217,N_3938,N_3258);
nor U4218 (N_4218,N_3348,N_3126);
and U4219 (N_4219,N_3556,N_3339);
nand U4220 (N_4220,N_3740,N_3076);
and U4221 (N_4221,N_3148,N_3130);
nor U4222 (N_4222,N_3162,N_3968);
or U4223 (N_4223,N_3265,N_3476);
and U4224 (N_4224,N_3187,N_3840);
or U4225 (N_4225,N_3454,N_3755);
or U4226 (N_4226,N_3342,N_3022);
nor U4227 (N_4227,N_3681,N_3231);
nand U4228 (N_4228,N_3965,N_3765);
nand U4229 (N_4229,N_3950,N_3140);
nand U4230 (N_4230,N_3580,N_3733);
or U4231 (N_4231,N_3759,N_3385);
nand U4232 (N_4232,N_3341,N_3012);
nand U4233 (N_4233,N_3516,N_3479);
or U4234 (N_4234,N_3201,N_3562);
nor U4235 (N_4235,N_3336,N_3298);
nor U4236 (N_4236,N_3312,N_3974);
or U4237 (N_4237,N_3849,N_3354);
nor U4238 (N_4238,N_3424,N_3521);
or U4239 (N_4239,N_3181,N_3315);
nand U4240 (N_4240,N_3270,N_3387);
nor U4241 (N_4241,N_3528,N_3928);
nor U4242 (N_4242,N_3835,N_3944);
nor U4243 (N_4243,N_3153,N_3671);
nor U4244 (N_4244,N_3790,N_3906);
or U4245 (N_4245,N_3820,N_3410);
nand U4246 (N_4246,N_3858,N_3047);
and U4247 (N_4247,N_3542,N_3946);
and U4248 (N_4248,N_3527,N_3802);
xnor U4249 (N_4249,N_3434,N_3213);
and U4250 (N_4250,N_3014,N_3247);
or U4251 (N_4251,N_3159,N_3489);
and U4252 (N_4252,N_3321,N_3550);
and U4253 (N_4253,N_3523,N_3218);
nand U4254 (N_4254,N_3942,N_3700);
nand U4255 (N_4255,N_3526,N_3482);
nor U4256 (N_4256,N_3935,N_3188);
or U4257 (N_4257,N_3578,N_3260);
and U4258 (N_4258,N_3329,N_3064);
and U4259 (N_4259,N_3963,N_3872);
or U4260 (N_4260,N_3094,N_3623);
or U4261 (N_4261,N_3009,N_3122);
or U4262 (N_4262,N_3803,N_3757);
or U4263 (N_4263,N_3682,N_3500);
and U4264 (N_4264,N_3254,N_3962);
nand U4265 (N_4265,N_3557,N_3894);
and U4266 (N_4266,N_3805,N_3281);
and U4267 (N_4267,N_3210,N_3380);
or U4268 (N_4268,N_3639,N_3524);
nand U4269 (N_4269,N_3384,N_3421);
or U4270 (N_4270,N_3878,N_3912);
nand U4271 (N_4271,N_3754,N_3607);
and U4272 (N_4272,N_3664,N_3508);
xnor U4273 (N_4273,N_3850,N_3307);
and U4274 (N_4274,N_3914,N_3758);
or U4275 (N_4275,N_3318,N_3018);
nor U4276 (N_4276,N_3824,N_3902);
and U4277 (N_4277,N_3346,N_3823);
nor U4278 (N_4278,N_3344,N_3635);
and U4279 (N_4279,N_3169,N_3807);
nor U4280 (N_4280,N_3224,N_3515);
nor U4281 (N_4281,N_3806,N_3457);
or U4282 (N_4282,N_3278,N_3464);
nor U4283 (N_4283,N_3027,N_3999);
nor U4284 (N_4284,N_3395,N_3036);
or U4285 (N_4285,N_3328,N_3888);
or U4286 (N_4286,N_3990,N_3383);
nand U4287 (N_4287,N_3412,N_3616);
nor U4288 (N_4288,N_3655,N_3289);
or U4289 (N_4289,N_3501,N_3214);
nand U4290 (N_4290,N_3695,N_3350);
or U4291 (N_4291,N_3880,N_3481);
nand U4292 (N_4292,N_3138,N_3783);
nor U4293 (N_4293,N_3685,N_3020);
or U4294 (N_4294,N_3630,N_3125);
nand U4295 (N_4295,N_3349,N_3299);
or U4296 (N_4296,N_3427,N_3091);
or U4297 (N_4297,N_3959,N_3762);
nor U4298 (N_4298,N_3739,N_3908);
nand U4299 (N_4299,N_3019,N_3203);
nor U4300 (N_4300,N_3103,N_3486);
nor U4301 (N_4301,N_3507,N_3110);
nor U4302 (N_4302,N_3779,N_3749);
nand U4303 (N_4303,N_3763,N_3723);
nand U4304 (N_4304,N_3543,N_3164);
nor U4305 (N_4305,N_3804,N_3513);
nor U4306 (N_4306,N_3167,N_3078);
nor U4307 (N_4307,N_3711,N_3376);
nand U4308 (N_4308,N_3632,N_3993);
or U4309 (N_4309,N_3323,N_3921);
and U4310 (N_4310,N_3405,N_3511);
xor U4311 (N_4311,N_3705,N_3211);
and U4312 (N_4312,N_3495,N_3306);
and U4313 (N_4313,N_3120,N_3446);
nand U4314 (N_4314,N_3386,N_3698);
nand U4315 (N_4315,N_3264,N_3136);
nand U4316 (N_4316,N_3989,N_3920);
nor U4317 (N_4317,N_3929,N_3061);
or U4318 (N_4318,N_3003,N_3728);
nor U4319 (N_4319,N_3391,N_3853);
nand U4320 (N_4320,N_3595,N_3183);
nand U4321 (N_4321,N_3180,N_3786);
xnor U4322 (N_4322,N_3566,N_3817);
and U4323 (N_4323,N_3877,N_3161);
or U4324 (N_4324,N_3548,N_3082);
and U4325 (N_4325,N_3106,N_3172);
or U4326 (N_4326,N_3144,N_3704);
or U4327 (N_4327,N_3333,N_3812);
or U4328 (N_4328,N_3179,N_3792);
xor U4329 (N_4329,N_3165,N_3272);
and U4330 (N_4330,N_3388,N_3070);
nor U4331 (N_4331,N_3417,N_3271);
xor U4332 (N_4332,N_3801,N_3869);
nand U4333 (N_4333,N_3374,N_3026);
or U4334 (N_4334,N_3426,N_3687);
nor U4335 (N_4335,N_3956,N_3006);
and U4336 (N_4336,N_3206,N_3331);
or U4337 (N_4337,N_3913,N_3400);
or U4338 (N_4338,N_3982,N_3748);
nand U4339 (N_4339,N_3087,N_3433);
and U4340 (N_4340,N_3285,N_3248);
and U4341 (N_4341,N_3361,N_3077);
and U4342 (N_4342,N_3905,N_3686);
nand U4343 (N_4343,N_3279,N_3095);
and U4344 (N_4344,N_3326,N_3397);
nand U4345 (N_4345,N_3822,N_3266);
and U4346 (N_4346,N_3459,N_3833);
and U4347 (N_4347,N_3168,N_3864);
xor U4348 (N_4348,N_3408,N_3290);
xor U4349 (N_4349,N_3450,N_3296);
or U4350 (N_4350,N_3043,N_3411);
nand U4351 (N_4351,N_3357,N_3227);
or U4352 (N_4352,N_3176,N_3119);
nand U4353 (N_4353,N_3498,N_3531);
or U4354 (N_4354,N_3626,N_3764);
nor U4355 (N_4355,N_3216,N_3871);
nor U4356 (N_4356,N_3887,N_3662);
nor U4357 (N_4357,N_3743,N_3190);
nor U4358 (N_4358,N_3310,N_3041);
nor U4359 (N_4359,N_3137,N_3469);
nand U4360 (N_4360,N_3752,N_3363);
nand U4361 (N_4361,N_3282,N_3834);
or U4362 (N_4362,N_3599,N_3052);
nand U4363 (N_4363,N_3610,N_3791);
and U4364 (N_4364,N_3985,N_3617);
nor U4365 (N_4365,N_3319,N_3373);
nor U4366 (N_4366,N_3782,N_3468);
or U4367 (N_4367,N_3230,N_3977);
or U4368 (N_4368,N_3225,N_3463);
or U4369 (N_4369,N_3451,N_3330);
nor U4370 (N_4370,N_3756,N_3672);
or U4371 (N_4371,N_3857,N_3995);
nor U4372 (N_4372,N_3652,N_3953);
or U4373 (N_4373,N_3115,N_3406);
nand U4374 (N_4374,N_3831,N_3519);
nand U4375 (N_4375,N_3544,N_3838);
nand U4376 (N_4376,N_3567,N_3787);
nor U4377 (N_4377,N_3606,N_3522);
nand U4378 (N_4378,N_3040,N_3008);
nand U4379 (N_4379,N_3324,N_3654);
or U4380 (N_4380,N_3860,N_3293);
or U4381 (N_4381,N_3394,N_3725);
nand U4382 (N_4382,N_3539,N_3660);
xnor U4383 (N_4383,N_3646,N_3575);
nand U4384 (N_4384,N_3969,N_3093);
or U4385 (N_4385,N_3583,N_3746);
or U4386 (N_4386,N_3625,N_3415);
nor U4387 (N_4387,N_3845,N_3098);
nand U4388 (N_4388,N_3775,N_3922);
and U4389 (N_4389,N_3368,N_3673);
nand U4390 (N_4390,N_3084,N_3220);
xnor U4391 (N_4391,N_3275,N_3088);
or U4392 (N_4392,N_3462,N_3438);
nor U4393 (N_4393,N_3497,N_3366);
nor U4394 (N_4394,N_3268,N_3355);
and U4395 (N_4395,N_3287,N_3605);
nor U4396 (N_4396,N_3768,N_3742);
nand U4397 (N_4397,N_3448,N_3919);
nand U4398 (N_4398,N_3105,N_3825);
nand U4399 (N_4399,N_3062,N_3591);
xor U4400 (N_4400,N_3393,N_3017);
or U4401 (N_4401,N_3980,N_3925);
nor U4402 (N_4402,N_3666,N_3910);
nor U4403 (N_4403,N_3692,N_3303);
nor U4404 (N_4404,N_3496,N_3173);
or U4405 (N_4405,N_3283,N_3584);
nor U4406 (N_4406,N_3854,N_3044);
or U4407 (N_4407,N_3680,N_3403);
nand U4408 (N_4408,N_3389,N_3297);
and U4409 (N_4409,N_3826,N_3729);
nand U4410 (N_4410,N_3612,N_3322);
nor U4411 (N_4411,N_3808,N_3255);
nor U4412 (N_4412,N_3487,N_3419);
nand U4413 (N_4413,N_3478,N_3048);
nand U4414 (N_4414,N_3710,N_3624);
and U4415 (N_4415,N_3109,N_3867);
and U4416 (N_4416,N_3537,N_3209);
and U4417 (N_4417,N_3884,N_3753);
nor U4418 (N_4418,N_3284,N_3039);
nor U4419 (N_4419,N_3509,N_3097);
or U4420 (N_4420,N_3701,N_3994);
nor U4421 (N_4421,N_3332,N_3563);
or U4422 (N_4422,N_3788,N_3471);
nor U4423 (N_4423,N_3885,N_3794);
nand U4424 (N_4424,N_3021,N_3586);
nor U4425 (N_4425,N_3316,N_3080);
nand U4426 (N_4426,N_3745,N_3750);
xor U4427 (N_4427,N_3147,N_3170);
nand U4428 (N_4428,N_3353,N_3951);
nand U4429 (N_4429,N_3081,N_3249);
nor U4430 (N_4430,N_3277,N_3604);
or U4431 (N_4431,N_3601,N_3191);
nor U4432 (N_4432,N_3245,N_3219);
or U4433 (N_4433,N_3086,N_3665);
nor U4434 (N_4434,N_3243,N_3810);
and U4435 (N_4435,N_3597,N_3863);
or U4436 (N_4436,N_3241,N_3798);
or U4437 (N_4437,N_3302,N_3320);
nor U4438 (N_4438,N_3948,N_3727);
or U4439 (N_4439,N_3314,N_3830);
nand U4440 (N_4440,N_3390,N_3577);
nor U4441 (N_4441,N_3644,N_3667);
or U4442 (N_4442,N_3141,N_3053);
and U4443 (N_4443,N_3267,N_3916);
or U4444 (N_4444,N_3259,N_3453);
nand U4445 (N_4445,N_3236,N_3428);
nand U4446 (N_4446,N_3458,N_3485);
nand U4447 (N_4447,N_3971,N_3118);
or U4448 (N_4448,N_3514,N_3112);
and U4449 (N_4449,N_3811,N_3576);
or U4450 (N_4450,N_3536,N_3198);
xnor U4451 (N_4451,N_3351,N_3647);
or U4452 (N_4452,N_3534,N_3325);
nor U4453 (N_4453,N_3444,N_3139);
nor U4454 (N_4454,N_3587,N_3063);
or U4455 (N_4455,N_3352,N_3731);
or U4456 (N_4456,N_3658,N_3541);
nand U4457 (N_4457,N_3722,N_3789);
or U4458 (N_4458,N_3618,N_3046);
and U4459 (N_4459,N_3966,N_3520);
nand U4460 (N_4460,N_3619,N_3073);
xnor U4461 (N_4461,N_3988,N_3280);
or U4462 (N_4462,N_3847,N_3382);
or U4463 (N_4463,N_3690,N_3629);
nor U4464 (N_4464,N_3470,N_3529);
and U4465 (N_4465,N_3238,N_3874);
nor U4466 (N_4466,N_3538,N_3708);
nand U4467 (N_4467,N_3402,N_3689);
nor U4468 (N_4468,N_3456,N_3636);
nand U4469 (N_4469,N_3171,N_3949);
xor U4470 (N_4470,N_3572,N_3505);
and U4471 (N_4471,N_3234,N_3294);
nand U4472 (N_4472,N_3015,N_3193);
or U4473 (N_4473,N_3773,N_3257);
nor U4474 (N_4474,N_3901,N_3035);
and U4475 (N_4475,N_3659,N_3532);
nand U4476 (N_4476,N_3107,N_3848);
and U4477 (N_4477,N_3175,N_3882);
nand U4478 (N_4478,N_3613,N_3676);
nand U4479 (N_4479,N_3893,N_3926);
nor U4480 (N_4480,N_3396,N_3818);
nor U4481 (N_4481,N_3868,N_3054);
or U4482 (N_4482,N_3997,N_3465);
nor U4483 (N_4483,N_3964,N_3295);
nor U4484 (N_4484,N_3553,N_3650);
nor U4485 (N_4485,N_3222,N_3602);
and U4486 (N_4486,N_3340,N_3250);
and U4487 (N_4487,N_3837,N_3886);
nor U4488 (N_4488,N_3895,N_3592);
xnor U4489 (N_4489,N_3724,N_3579);
nand U4490 (N_4490,N_3195,N_3038);
and U4491 (N_4491,N_3101,N_3375);
nand U4492 (N_4492,N_3422,N_3031);
and U4493 (N_4493,N_3291,N_3079);
nor U4494 (N_4494,N_3891,N_3645);
and U4495 (N_4495,N_3917,N_3050);
nor U4496 (N_4496,N_3627,N_3998);
nor U4497 (N_4497,N_3707,N_3628);
and U4498 (N_4498,N_3007,N_3111);
and U4499 (N_4499,N_3693,N_3432);
or U4500 (N_4500,N_3268,N_3511);
nor U4501 (N_4501,N_3164,N_3205);
and U4502 (N_4502,N_3451,N_3444);
nand U4503 (N_4503,N_3613,N_3936);
nand U4504 (N_4504,N_3230,N_3705);
or U4505 (N_4505,N_3861,N_3243);
nand U4506 (N_4506,N_3310,N_3656);
nand U4507 (N_4507,N_3938,N_3057);
or U4508 (N_4508,N_3397,N_3436);
and U4509 (N_4509,N_3265,N_3137);
or U4510 (N_4510,N_3881,N_3898);
and U4511 (N_4511,N_3259,N_3219);
or U4512 (N_4512,N_3131,N_3737);
nor U4513 (N_4513,N_3930,N_3745);
nand U4514 (N_4514,N_3130,N_3822);
nor U4515 (N_4515,N_3724,N_3607);
nor U4516 (N_4516,N_3545,N_3998);
and U4517 (N_4517,N_3011,N_3152);
and U4518 (N_4518,N_3525,N_3107);
nand U4519 (N_4519,N_3285,N_3297);
nand U4520 (N_4520,N_3531,N_3039);
xor U4521 (N_4521,N_3745,N_3136);
and U4522 (N_4522,N_3784,N_3133);
nand U4523 (N_4523,N_3010,N_3785);
nor U4524 (N_4524,N_3423,N_3285);
or U4525 (N_4525,N_3521,N_3392);
and U4526 (N_4526,N_3921,N_3773);
nand U4527 (N_4527,N_3063,N_3829);
xor U4528 (N_4528,N_3845,N_3180);
and U4529 (N_4529,N_3221,N_3152);
nor U4530 (N_4530,N_3609,N_3099);
nand U4531 (N_4531,N_3804,N_3176);
nor U4532 (N_4532,N_3838,N_3982);
nand U4533 (N_4533,N_3787,N_3884);
nor U4534 (N_4534,N_3251,N_3599);
nand U4535 (N_4535,N_3105,N_3235);
or U4536 (N_4536,N_3873,N_3056);
or U4537 (N_4537,N_3420,N_3417);
and U4538 (N_4538,N_3967,N_3946);
nand U4539 (N_4539,N_3454,N_3768);
nor U4540 (N_4540,N_3196,N_3918);
nor U4541 (N_4541,N_3044,N_3978);
nor U4542 (N_4542,N_3457,N_3811);
or U4543 (N_4543,N_3839,N_3395);
nand U4544 (N_4544,N_3763,N_3324);
nand U4545 (N_4545,N_3183,N_3565);
xnor U4546 (N_4546,N_3357,N_3027);
nand U4547 (N_4547,N_3746,N_3806);
nor U4548 (N_4548,N_3254,N_3998);
nor U4549 (N_4549,N_3461,N_3662);
and U4550 (N_4550,N_3778,N_3510);
nor U4551 (N_4551,N_3541,N_3759);
and U4552 (N_4552,N_3361,N_3858);
and U4553 (N_4553,N_3962,N_3842);
nor U4554 (N_4554,N_3699,N_3006);
or U4555 (N_4555,N_3714,N_3656);
nor U4556 (N_4556,N_3247,N_3516);
and U4557 (N_4557,N_3660,N_3836);
nor U4558 (N_4558,N_3457,N_3435);
nand U4559 (N_4559,N_3740,N_3355);
or U4560 (N_4560,N_3963,N_3001);
nor U4561 (N_4561,N_3948,N_3033);
and U4562 (N_4562,N_3818,N_3102);
and U4563 (N_4563,N_3455,N_3926);
or U4564 (N_4564,N_3665,N_3746);
and U4565 (N_4565,N_3966,N_3016);
or U4566 (N_4566,N_3954,N_3574);
and U4567 (N_4567,N_3042,N_3702);
and U4568 (N_4568,N_3925,N_3276);
nand U4569 (N_4569,N_3056,N_3863);
nor U4570 (N_4570,N_3838,N_3153);
nand U4571 (N_4571,N_3651,N_3176);
nand U4572 (N_4572,N_3139,N_3735);
or U4573 (N_4573,N_3234,N_3836);
and U4574 (N_4574,N_3676,N_3481);
nand U4575 (N_4575,N_3688,N_3877);
nor U4576 (N_4576,N_3678,N_3107);
or U4577 (N_4577,N_3445,N_3409);
nor U4578 (N_4578,N_3488,N_3658);
nand U4579 (N_4579,N_3965,N_3988);
or U4580 (N_4580,N_3816,N_3862);
nand U4581 (N_4581,N_3584,N_3306);
nand U4582 (N_4582,N_3862,N_3516);
xor U4583 (N_4583,N_3154,N_3509);
nor U4584 (N_4584,N_3092,N_3481);
and U4585 (N_4585,N_3093,N_3388);
or U4586 (N_4586,N_3921,N_3611);
and U4587 (N_4587,N_3763,N_3497);
or U4588 (N_4588,N_3831,N_3263);
nand U4589 (N_4589,N_3819,N_3344);
nor U4590 (N_4590,N_3487,N_3769);
nor U4591 (N_4591,N_3819,N_3462);
nor U4592 (N_4592,N_3910,N_3570);
and U4593 (N_4593,N_3834,N_3829);
nor U4594 (N_4594,N_3144,N_3775);
nor U4595 (N_4595,N_3926,N_3471);
and U4596 (N_4596,N_3063,N_3799);
xor U4597 (N_4597,N_3996,N_3173);
nand U4598 (N_4598,N_3520,N_3481);
nand U4599 (N_4599,N_3731,N_3333);
nand U4600 (N_4600,N_3869,N_3506);
and U4601 (N_4601,N_3989,N_3094);
or U4602 (N_4602,N_3560,N_3304);
nor U4603 (N_4603,N_3573,N_3213);
or U4604 (N_4604,N_3535,N_3386);
and U4605 (N_4605,N_3665,N_3417);
and U4606 (N_4606,N_3482,N_3889);
or U4607 (N_4607,N_3058,N_3136);
and U4608 (N_4608,N_3108,N_3531);
and U4609 (N_4609,N_3661,N_3075);
nor U4610 (N_4610,N_3404,N_3949);
and U4611 (N_4611,N_3409,N_3321);
nand U4612 (N_4612,N_3910,N_3469);
nor U4613 (N_4613,N_3383,N_3348);
nand U4614 (N_4614,N_3604,N_3094);
and U4615 (N_4615,N_3777,N_3424);
nor U4616 (N_4616,N_3805,N_3838);
nor U4617 (N_4617,N_3342,N_3242);
nand U4618 (N_4618,N_3738,N_3811);
and U4619 (N_4619,N_3333,N_3831);
and U4620 (N_4620,N_3693,N_3231);
nor U4621 (N_4621,N_3381,N_3008);
nor U4622 (N_4622,N_3523,N_3545);
or U4623 (N_4623,N_3573,N_3729);
nor U4624 (N_4624,N_3181,N_3782);
and U4625 (N_4625,N_3078,N_3433);
or U4626 (N_4626,N_3481,N_3546);
nand U4627 (N_4627,N_3604,N_3926);
nand U4628 (N_4628,N_3868,N_3157);
nor U4629 (N_4629,N_3893,N_3656);
nand U4630 (N_4630,N_3214,N_3713);
nor U4631 (N_4631,N_3739,N_3495);
or U4632 (N_4632,N_3581,N_3481);
nor U4633 (N_4633,N_3736,N_3147);
and U4634 (N_4634,N_3783,N_3727);
or U4635 (N_4635,N_3933,N_3366);
nand U4636 (N_4636,N_3741,N_3082);
nor U4637 (N_4637,N_3584,N_3570);
or U4638 (N_4638,N_3205,N_3612);
or U4639 (N_4639,N_3034,N_3610);
and U4640 (N_4640,N_3152,N_3268);
nor U4641 (N_4641,N_3102,N_3615);
or U4642 (N_4642,N_3511,N_3062);
nor U4643 (N_4643,N_3717,N_3685);
or U4644 (N_4644,N_3803,N_3438);
nor U4645 (N_4645,N_3000,N_3265);
nand U4646 (N_4646,N_3067,N_3801);
or U4647 (N_4647,N_3176,N_3343);
nor U4648 (N_4648,N_3531,N_3461);
nor U4649 (N_4649,N_3782,N_3439);
or U4650 (N_4650,N_3903,N_3744);
or U4651 (N_4651,N_3996,N_3487);
or U4652 (N_4652,N_3162,N_3337);
nand U4653 (N_4653,N_3730,N_3122);
nor U4654 (N_4654,N_3156,N_3948);
or U4655 (N_4655,N_3379,N_3681);
nand U4656 (N_4656,N_3510,N_3796);
or U4657 (N_4657,N_3037,N_3193);
or U4658 (N_4658,N_3064,N_3370);
or U4659 (N_4659,N_3658,N_3328);
nor U4660 (N_4660,N_3061,N_3133);
nand U4661 (N_4661,N_3559,N_3331);
nand U4662 (N_4662,N_3157,N_3516);
and U4663 (N_4663,N_3846,N_3389);
xnor U4664 (N_4664,N_3556,N_3251);
or U4665 (N_4665,N_3597,N_3862);
nand U4666 (N_4666,N_3636,N_3961);
and U4667 (N_4667,N_3573,N_3313);
nand U4668 (N_4668,N_3221,N_3854);
nand U4669 (N_4669,N_3662,N_3888);
nand U4670 (N_4670,N_3992,N_3977);
nor U4671 (N_4671,N_3982,N_3317);
and U4672 (N_4672,N_3866,N_3516);
nand U4673 (N_4673,N_3711,N_3115);
nand U4674 (N_4674,N_3775,N_3060);
and U4675 (N_4675,N_3301,N_3407);
or U4676 (N_4676,N_3287,N_3214);
or U4677 (N_4677,N_3800,N_3593);
and U4678 (N_4678,N_3496,N_3712);
nand U4679 (N_4679,N_3940,N_3733);
nand U4680 (N_4680,N_3248,N_3613);
xnor U4681 (N_4681,N_3317,N_3802);
and U4682 (N_4682,N_3424,N_3991);
nand U4683 (N_4683,N_3151,N_3801);
and U4684 (N_4684,N_3703,N_3345);
or U4685 (N_4685,N_3793,N_3492);
nor U4686 (N_4686,N_3546,N_3420);
nor U4687 (N_4687,N_3261,N_3013);
and U4688 (N_4688,N_3626,N_3182);
and U4689 (N_4689,N_3979,N_3784);
or U4690 (N_4690,N_3942,N_3863);
or U4691 (N_4691,N_3872,N_3630);
xnor U4692 (N_4692,N_3642,N_3735);
nand U4693 (N_4693,N_3857,N_3722);
or U4694 (N_4694,N_3415,N_3168);
nand U4695 (N_4695,N_3153,N_3112);
nor U4696 (N_4696,N_3638,N_3849);
nand U4697 (N_4697,N_3267,N_3391);
nand U4698 (N_4698,N_3369,N_3256);
or U4699 (N_4699,N_3990,N_3099);
nor U4700 (N_4700,N_3956,N_3604);
nand U4701 (N_4701,N_3390,N_3322);
or U4702 (N_4702,N_3155,N_3583);
and U4703 (N_4703,N_3169,N_3173);
nand U4704 (N_4704,N_3923,N_3486);
nor U4705 (N_4705,N_3113,N_3257);
and U4706 (N_4706,N_3972,N_3473);
nor U4707 (N_4707,N_3626,N_3308);
or U4708 (N_4708,N_3784,N_3435);
nand U4709 (N_4709,N_3599,N_3735);
or U4710 (N_4710,N_3937,N_3459);
nand U4711 (N_4711,N_3932,N_3915);
and U4712 (N_4712,N_3225,N_3304);
or U4713 (N_4713,N_3530,N_3275);
nand U4714 (N_4714,N_3899,N_3298);
nand U4715 (N_4715,N_3956,N_3002);
nand U4716 (N_4716,N_3302,N_3154);
nand U4717 (N_4717,N_3747,N_3822);
and U4718 (N_4718,N_3476,N_3243);
nor U4719 (N_4719,N_3676,N_3079);
and U4720 (N_4720,N_3864,N_3677);
and U4721 (N_4721,N_3737,N_3661);
nor U4722 (N_4722,N_3387,N_3840);
and U4723 (N_4723,N_3074,N_3711);
and U4724 (N_4724,N_3772,N_3877);
nor U4725 (N_4725,N_3588,N_3229);
and U4726 (N_4726,N_3659,N_3998);
and U4727 (N_4727,N_3054,N_3429);
nor U4728 (N_4728,N_3346,N_3021);
and U4729 (N_4729,N_3929,N_3424);
nand U4730 (N_4730,N_3412,N_3674);
nor U4731 (N_4731,N_3481,N_3334);
nand U4732 (N_4732,N_3916,N_3683);
nand U4733 (N_4733,N_3978,N_3929);
nor U4734 (N_4734,N_3508,N_3321);
or U4735 (N_4735,N_3006,N_3803);
and U4736 (N_4736,N_3761,N_3755);
or U4737 (N_4737,N_3466,N_3508);
and U4738 (N_4738,N_3902,N_3052);
and U4739 (N_4739,N_3818,N_3580);
nand U4740 (N_4740,N_3563,N_3459);
and U4741 (N_4741,N_3033,N_3002);
nand U4742 (N_4742,N_3010,N_3149);
nor U4743 (N_4743,N_3640,N_3848);
nor U4744 (N_4744,N_3146,N_3587);
nand U4745 (N_4745,N_3120,N_3471);
nor U4746 (N_4746,N_3082,N_3571);
nor U4747 (N_4747,N_3265,N_3621);
or U4748 (N_4748,N_3468,N_3505);
and U4749 (N_4749,N_3893,N_3923);
and U4750 (N_4750,N_3485,N_3895);
nor U4751 (N_4751,N_3852,N_3496);
and U4752 (N_4752,N_3810,N_3837);
or U4753 (N_4753,N_3252,N_3006);
and U4754 (N_4754,N_3220,N_3790);
nand U4755 (N_4755,N_3125,N_3740);
nor U4756 (N_4756,N_3516,N_3336);
nor U4757 (N_4757,N_3567,N_3317);
or U4758 (N_4758,N_3681,N_3167);
nand U4759 (N_4759,N_3771,N_3070);
nor U4760 (N_4760,N_3448,N_3512);
nand U4761 (N_4761,N_3437,N_3121);
and U4762 (N_4762,N_3395,N_3622);
or U4763 (N_4763,N_3959,N_3790);
or U4764 (N_4764,N_3028,N_3466);
nor U4765 (N_4765,N_3976,N_3131);
nand U4766 (N_4766,N_3220,N_3900);
or U4767 (N_4767,N_3092,N_3709);
or U4768 (N_4768,N_3140,N_3915);
nor U4769 (N_4769,N_3905,N_3583);
or U4770 (N_4770,N_3546,N_3013);
and U4771 (N_4771,N_3455,N_3966);
nor U4772 (N_4772,N_3507,N_3418);
nand U4773 (N_4773,N_3418,N_3855);
nor U4774 (N_4774,N_3111,N_3547);
nor U4775 (N_4775,N_3489,N_3058);
xor U4776 (N_4776,N_3211,N_3202);
or U4777 (N_4777,N_3631,N_3031);
or U4778 (N_4778,N_3090,N_3208);
and U4779 (N_4779,N_3211,N_3521);
nand U4780 (N_4780,N_3927,N_3127);
and U4781 (N_4781,N_3046,N_3904);
nor U4782 (N_4782,N_3929,N_3694);
nand U4783 (N_4783,N_3032,N_3071);
and U4784 (N_4784,N_3650,N_3783);
nor U4785 (N_4785,N_3825,N_3497);
xor U4786 (N_4786,N_3646,N_3104);
nor U4787 (N_4787,N_3193,N_3511);
nor U4788 (N_4788,N_3194,N_3063);
and U4789 (N_4789,N_3109,N_3026);
nand U4790 (N_4790,N_3720,N_3839);
nor U4791 (N_4791,N_3660,N_3418);
nor U4792 (N_4792,N_3745,N_3620);
nor U4793 (N_4793,N_3778,N_3170);
nand U4794 (N_4794,N_3801,N_3939);
or U4795 (N_4795,N_3732,N_3170);
nor U4796 (N_4796,N_3803,N_3237);
nor U4797 (N_4797,N_3570,N_3475);
or U4798 (N_4798,N_3594,N_3866);
or U4799 (N_4799,N_3460,N_3648);
or U4800 (N_4800,N_3228,N_3696);
nand U4801 (N_4801,N_3368,N_3375);
or U4802 (N_4802,N_3887,N_3995);
and U4803 (N_4803,N_3569,N_3176);
and U4804 (N_4804,N_3177,N_3925);
and U4805 (N_4805,N_3875,N_3462);
and U4806 (N_4806,N_3823,N_3707);
nand U4807 (N_4807,N_3440,N_3088);
nor U4808 (N_4808,N_3229,N_3893);
nand U4809 (N_4809,N_3265,N_3540);
and U4810 (N_4810,N_3481,N_3133);
or U4811 (N_4811,N_3865,N_3152);
nor U4812 (N_4812,N_3155,N_3677);
and U4813 (N_4813,N_3118,N_3089);
nor U4814 (N_4814,N_3594,N_3389);
nand U4815 (N_4815,N_3534,N_3520);
and U4816 (N_4816,N_3239,N_3694);
nand U4817 (N_4817,N_3276,N_3758);
nor U4818 (N_4818,N_3610,N_3720);
nor U4819 (N_4819,N_3823,N_3080);
and U4820 (N_4820,N_3330,N_3708);
nand U4821 (N_4821,N_3758,N_3511);
and U4822 (N_4822,N_3810,N_3550);
xnor U4823 (N_4823,N_3219,N_3752);
or U4824 (N_4824,N_3716,N_3363);
nand U4825 (N_4825,N_3627,N_3727);
nand U4826 (N_4826,N_3627,N_3752);
xor U4827 (N_4827,N_3943,N_3317);
nand U4828 (N_4828,N_3526,N_3842);
and U4829 (N_4829,N_3455,N_3726);
and U4830 (N_4830,N_3051,N_3611);
or U4831 (N_4831,N_3413,N_3232);
nor U4832 (N_4832,N_3331,N_3974);
and U4833 (N_4833,N_3327,N_3241);
and U4834 (N_4834,N_3952,N_3405);
nor U4835 (N_4835,N_3792,N_3661);
and U4836 (N_4836,N_3425,N_3095);
nand U4837 (N_4837,N_3818,N_3948);
xor U4838 (N_4838,N_3038,N_3431);
or U4839 (N_4839,N_3642,N_3997);
or U4840 (N_4840,N_3076,N_3013);
or U4841 (N_4841,N_3217,N_3891);
nor U4842 (N_4842,N_3420,N_3758);
nand U4843 (N_4843,N_3228,N_3741);
xor U4844 (N_4844,N_3026,N_3680);
nor U4845 (N_4845,N_3002,N_3274);
and U4846 (N_4846,N_3527,N_3119);
nand U4847 (N_4847,N_3512,N_3804);
or U4848 (N_4848,N_3213,N_3215);
nand U4849 (N_4849,N_3167,N_3830);
nor U4850 (N_4850,N_3190,N_3754);
and U4851 (N_4851,N_3446,N_3494);
and U4852 (N_4852,N_3646,N_3847);
nand U4853 (N_4853,N_3682,N_3819);
nor U4854 (N_4854,N_3200,N_3260);
and U4855 (N_4855,N_3941,N_3298);
nand U4856 (N_4856,N_3832,N_3205);
or U4857 (N_4857,N_3997,N_3014);
xor U4858 (N_4858,N_3948,N_3419);
or U4859 (N_4859,N_3145,N_3044);
nand U4860 (N_4860,N_3054,N_3995);
nor U4861 (N_4861,N_3696,N_3637);
nor U4862 (N_4862,N_3461,N_3414);
nand U4863 (N_4863,N_3787,N_3407);
nor U4864 (N_4864,N_3019,N_3839);
nand U4865 (N_4865,N_3609,N_3452);
or U4866 (N_4866,N_3200,N_3760);
nor U4867 (N_4867,N_3288,N_3609);
nor U4868 (N_4868,N_3435,N_3474);
or U4869 (N_4869,N_3303,N_3600);
nand U4870 (N_4870,N_3425,N_3991);
nor U4871 (N_4871,N_3368,N_3920);
nand U4872 (N_4872,N_3691,N_3803);
nand U4873 (N_4873,N_3022,N_3685);
nand U4874 (N_4874,N_3162,N_3419);
or U4875 (N_4875,N_3248,N_3321);
nor U4876 (N_4876,N_3161,N_3727);
nand U4877 (N_4877,N_3293,N_3637);
and U4878 (N_4878,N_3110,N_3059);
and U4879 (N_4879,N_3550,N_3071);
nor U4880 (N_4880,N_3326,N_3604);
and U4881 (N_4881,N_3704,N_3111);
nor U4882 (N_4882,N_3511,N_3731);
nor U4883 (N_4883,N_3409,N_3846);
nand U4884 (N_4884,N_3963,N_3241);
and U4885 (N_4885,N_3828,N_3231);
and U4886 (N_4886,N_3152,N_3742);
nand U4887 (N_4887,N_3864,N_3020);
or U4888 (N_4888,N_3282,N_3809);
and U4889 (N_4889,N_3763,N_3596);
nand U4890 (N_4890,N_3682,N_3940);
or U4891 (N_4891,N_3295,N_3659);
nor U4892 (N_4892,N_3432,N_3902);
and U4893 (N_4893,N_3468,N_3340);
nor U4894 (N_4894,N_3271,N_3107);
and U4895 (N_4895,N_3312,N_3240);
or U4896 (N_4896,N_3899,N_3002);
or U4897 (N_4897,N_3874,N_3704);
nor U4898 (N_4898,N_3028,N_3300);
or U4899 (N_4899,N_3514,N_3854);
or U4900 (N_4900,N_3389,N_3448);
nand U4901 (N_4901,N_3342,N_3180);
nand U4902 (N_4902,N_3962,N_3055);
nand U4903 (N_4903,N_3631,N_3533);
xor U4904 (N_4904,N_3531,N_3183);
and U4905 (N_4905,N_3344,N_3215);
and U4906 (N_4906,N_3935,N_3340);
nor U4907 (N_4907,N_3259,N_3789);
and U4908 (N_4908,N_3954,N_3599);
nor U4909 (N_4909,N_3721,N_3896);
and U4910 (N_4910,N_3537,N_3530);
and U4911 (N_4911,N_3771,N_3502);
and U4912 (N_4912,N_3922,N_3397);
and U4913 (N_4913,N_3272,N_3362);
or U4914 (N_4914,N_3010,N_3547);
nor U4915 (N_4915,N_3330,N_3402);
nand U4916 (N_4916,N_3863,N_3908);
and U4917 (N_4917,N_3871,N_3803);
or U4918 (N_4918,N_3585,N_3598);
and U4919 (N_4919,N_3550,N_3880);
and U4920 (N_4920,N_3302,N_3926);
nand U4921 (N_4921,N_3490,N_3270);
nand U4922 (N_4922,N_3598,N_3541);
and U4923 (N_4923,N_3809,N_3074);
nor U4924 (N_4924,N_3224,N_3828);
or U4925 (N_4925,N_3521,N_3138);
nor U4926 (N_4926,N_3614,N_3545);
and U4927 (N_4927,N_3975,N_3399);
nand U4928 (N_4928,N_3830,N_3679);
nor U4929 (N_4929,N_3849,N_3054);
and U4930 (N_4930,N_3444,N_3094);
nand U4931 (N_4931,N_3138,N_3529);
nor U4932 (N_4932,N_3865,N_3288);
nor U4933 (N_4933,N_3845,N_3371);
or U4934 (N_4934,N_3604,N_3716);
nor U4935 (N_4935,N_3074,N_3167);
or U4936 (N_4936,N_3183,N_3604);
nor U4937 (N_4937,N_3707,N_3175);
or U4938 (N_4938,N_3690,N_3380);
and U4939 (N_4939,N_3153,N_3562);
and U4940 (N_4940,N_3610,N_3020);
or U4941 (N_4941,N_3806,N_3831);
xor U4942 (N_4942,N_3744,N_3713);
and U4943 (N_4943,N_3303,N_3946);
and U4944 (N_4944,N_3605,N_3757);
or U4945 (N_4945,N_3212,N_3620);
or U4946 (N_4946,N_3163,N_3347);
nor U4947 (N_4947,N_3740,N_3954);
xor U4948 (N_4948,N_3591,N_3934);
or U4949 (N_4949,N_3586,N_3513);
nor U4950 (N_4950,N_3870,N_3475);
and U4951 (N_4951,N_3674,N_3000);
or U4952 (N_4952,N_3346,N_3899);
nand U4953 (N_4953,N_3382,N_3025);
nor U4954 (N_4954,N_3933,N_3113);
nand U4955 (N_4955,N_3603,N_3209);
and U4956 (N_4956,N_3363,N_3443);
nand U4957 (N_4957,N_3498,N_3073);
nor U4958 (N_4958,N_3568,N_3957);
and U4959 (N_4959,N_3415,N_3038);
nand U4960 (N_4960,N_3351,N_3369);
or U4961 (N_4961,N_3477,N_3453);
nor U4962 (N_4962,N_3935,N_3336);
nor U4963 (N_4963,N_3208,N_3777);
nor U4964 (N_4964,N_3234,N_3240);
nand U4965 (N_4965,N_3459,N_3424);
or U4966 (N_4966,N_3571,N_3450);
nand U4967 (N_4967,N_3993,N_3838);
or U4968 (N_4968,N_3930,N_3469);
and U4969 (N_4969,N_3649,N_3884);
and U4970 (N_4970,N_3361,N_3718);
nand U4971 (N_4971,N_3854,N_3580);
and U4972 (N_4972,N_3848,N_3556);
or U4973 (N_4973,N_3385,N_3566);
or U4974 (N_4974,N_3283,N_3655);
nand U4975 (N_4975,N_3285,N_3495);
or U4976 (N_4976,N_3347,N_3855);
xor U4977 (N_4977,N_3043,N_3875);
nand U4978 (N_4978,N_3412,N_3212);
nor U4979 (N_4979,N_3409,N_3525);
and U4980 (N_4980,N_3885,N_3415);
and U4981 (N_4981,N_3347,N_3042);
and U4982 (N_4982,N_3280,N_3620);
nand U4983 (N_4983,N_3159,N_3624);
or U4984 (N_4984,N_3420,N_3707);
nand U4985 (N_4985,N_3057,N_3537);
and U4986 (N_4986,N_3002,N_3298);
nand U4987 (N_4987,N_3504,N_3264);
nand U4988 (N_4988,N_3815,N_3501);
xnor U4989 (N_4989,N_3386,N_3733);
nand U4990 (N_4990,N_3207,N_3284);
nor U4991 (N_4991,N_3618,N_3488);
or U4992 (N_4992,N_3009,N_3341);
and U4993 (N_4993,N_3143,N_3751);
and U4994 (N_4994,N_3234,N_3164);
or U4995 (N_4995,N_3559,N_3418);
nor U4996 (N_4996,N_3582,N_3121);
and U4997 (N_4997,N_3453,N_3313);
or U4998 (N_4998,N_3288,N_3406);
or U4999 (N_4999,N_3762,N_3490);
nor UO_0 (O_0,N_4656,N_4147);
nand UO_1 (O_1,N_4315,N_4751);
nand UO_2 (O_2,N_4082,N_4094);
and UO_3 (O_3,N_4199,N_4237);
xor UO_4 (O_4,N_4570,N_4612);
nor UO_5 (O_5,N_4418,N_4731);
and UO_6 (O_6,N_4009,N_4867);
and UO_7 (O_7,N_4224,N_4872);
or UO_8 (O_8,N_4606,N_4104);
or UO_9 (O_9,N_4963,N_4496);
nand UO_10 (O_10,N_4578,N_4412);
or UO_11 (O_11,N_4300,N_4893);
and UO_12 (O_12,N_4248,N_4782);
or UO_13 (O_13,N_4194,N_4351);
or UO_14 (O_14,N_4938,N_4477);
nor UO_15 (O_15,N_4512,N_4688);
and UO_16 (O_16,N_4952,N_4352);
or UO_17 (O_17,N_4895,N_4202);
nand UO_18 (O_18,N_4400,N_4310);
nand UO_19 (O_19,N_4918,N_4288);
nor UO_20 (O_20,N_4627,N_4028);
or UO_21 (O_21,N_4281,N_4522);
nor UO_22 (O_22,N_4760,N_4915);
nor UO_23 (O_23,N_4831,N_4291);
or UO_24 (O_24,N_4255,N_4883);
nor UO_25 (O_25,N_4748,N_4107);
nor UO_26 (O_26,N_4457,N_4221);
nand UO_27 (O_27,N_4419,N_4478);
and UO_28 (O_28,N_4120,N_4102);
and UO_29 (O_29,N_4302,N_4700);
nand UO_30 (O_30,N_4758,N_4163);
nor UO_31 (O_31,N_4912,N_4474);
or UO_32 (O_32,N_4131,N_4565);
nand UO_33 (O_33,N_4220,N_4200);
nor UO_34 (O_34,N_4738,N_4601);
nor UO_35 (O_35,N_4123,N_4402);
and UO_36 (O_36,N_4567,N_4353);
and UO_37 (O_37,N_4811,N_4820);
and UO_38 (O_38,N_4002,N_4337);
nand UO_39 (O_39,N_4066,N_4156);
nand UO_40 (O_40,N_4257,N_4509);
and UO_41 (O_41,N_4306,N_4985);
and UO_42 (O_42,N_4296,N_4781);
nor UO_43 (O_43,N_4650,N_4260);
or UO_44 (O_44,N_4371,N_4339);
or UO_45 (O_45,N_4961,N_4940);
nand UO_46 (O_46,N_4110,N_4857);
xnor UO_47 (O_47,N_4114,N_4662);
and UO_48 (O_48,N_4953,N_4747);
and UO_49 (O_49,N_4446,N_4794);
and UO_50 (O_50,N_4385,N_4757);
and UO_51 (O_51,N_4463,N_4362);
nand UO_52 (O_52,N_4792,N_4099);
and UO_53 (O_53,N_4798,N_4005);
nor UO_54 (O_54,N_4648,N_4668);
nand UO_55 (O_55,N_4242,N_4313);
nand UO_56 (O_56,N_4414,N_4868);
nand UO_57 (O_57,N_4319,N_4946);
nand UO_58 (O_58,N_4990,N_4611);
or UO_59 (O_59,N_4112,N_4462);
nor UO_60 (O_60,N_4910,N_4455);
nor UO_61 (O_61,N_4238,N_4020);
nor UO_62 (O_62,N_4908,N_4592);
or UO_63 (O_63,N_4886,N_4435);
nor UO_64 (O_64,N_4962,N_4773);
or UO_65 (O_65,N_4537,N_4774);
nor UO_66 (O_66,N_4994,N_4479);
and UO_67 (O_67,N_4433,N_4027);
nand UO_68 (O_68,N_4041,N_4396);
and UO_69 (O_69,N_4776,N_4192);
and UO_70 (O_70,N_4620,N_4877);
nor UO_71 (O_71,N_4771,N_4837);
nor UO_72 (O_72,N_4763,N_4989);
nor UO_73 (O_73,N_4326,N_4491);
and UO_74 (O_74,N_4060,N_4923);
nand UO_75 (O_75,N_4888,N_4614);
and UO_76 (O_76,N_4906,N_4514);
and UO_77 (O_77,N_4501,N_4165);
nand UO_78 (O_78,N_4182,N_4866);
nand UO_79 (O_79,N_4884,N_4719);
nand UO_80 (O_80,N_4960,N_4919);
nand UO_81 (O_81,N_4451,N_4206);
and UO_82 (O_82,N_4393,N_4417);
nor UO_83 (O_83,N_4954,N_4164);
nand UO_84 (O_84,N_4880,N_4708);
nand UO_85 (O_85,N_4991,N_4711);
nor UO_86 (O_86,N_4768,N_4690);
or UO_87 (O_87,N_4588,N_4368);
or UO_88 (O_88,N_4964,N_4226);
nand UO_89 (O_89,N_4955,N_4997);
or UO_90 (O_90,N_4864,N_4272);
or UO_91 (O_91,N_4299,N_4812);
nand UO_92 (O_92,N_4784,N_4977);
or UO_93 (O_93,N_4373,N_4907);
nand UO_94 (O_94,N_4370,N_4610);
nand UO_95 (O_95,N_4116,N_4609);
and UO_96 (O_96,N_4580,N_4324);
xor UO_97 (O_97,N_4191,N_4593);
and UO_98 (O_98,N_4484,N_4127);
nor UO_99 (O_99,N_4138,N_4905);
and UO_100 (O_100,N_4208,N_4314);
or UO_101 (O_101,N_4615,N_4141);
or UO_102 (O_102,N_4383,N_4978);
nor UO_103 (O_103,N_4063,N_4322);
nand UO_104 (O_104,N_4848,N_4635);
xor UO_105 (O_105,N_4694,N_4456);
nor UO_106 (O_106,N_4675,N_4759);
nor UO_107 (O_107,N_4466,N_4480);
and UO_108 (O_108,N_4413,N_4925);
nand UO_109 (O_109,N_4619,N_4563);
and UO_110 (O_110,N_4641,N_4591);
nor UO_111 (O_111,N_4967,N_4956);
nor UO_112 (O_112,N_4388,N_4840);
xor UO_113 (O_113,N_4506,N_4723);
or UO_114 (O_114,N_4196,N_4111);
nor UO_115 (O_115,N_4295,N_4323);
and UO_116 (O_116,N_4770,N_4485);
nor UO_117 (O_117,N_4354,N_4423);
or UO_118 (O_118,N_4439,N_4232);
nor UO_119 (O_119,N_4437,N_4034);
or UO_120 (O_120,N_4924,N_4394);
or UO_121 (O_121,N_4608,N_4448);
and UO_122 (O_122,N_4330,N_4073);
nand UO_123 (O_123,N_4449,N_4160);
or UO_124 (O_124,N_4205,N_4011);
nand UO_125 (O_125,N_4079,N_4974);
nor UO_126 (O_126,N_4741,N_4654);
nor UO_127 (O_127,N_4465,N_4247);
nand UO_128 (O_128,N_4613,N_4420);
nand UO_129 (O_129,N_4280,N_4287);
nand UO_130 (O_130,N_4790,N_4950);
and UO_131 (O_131,N_4416,N_4637);
nor UO_132 (O_132,N_4630,N_4096);
or UO_133 (O_133,N_4498,N_4704);
or UO_134 (O_134,N_4007,N_4922);
or UO_135 (O_135,N_4495,N_4970);
or UO_136 (O_136,N_4148,N_4429);
nand UO_137 (O_137,N_4555,N_4017);
nor UO_138 (O_138,N_4019,N_4483);
and UO_139 (O_139,N_4469,N_4746);
xor UO_140 (O_140,N_4062,N_4810);
nor UO_141 (O_141,N_4240,N_4834);
or UO_142 (O_142,N_4603,N_4730);
and UO_143 (O_143,N_4827,N_4887);
and UO_144 (O_144,N_4292,N_4705);
or UO_145 (O_145,N_4742,N_4273);
or UO_146 (O_146,N_4604,N_4461);
nor UO_147 (O_147,N_4693,N_4438);
nor UO_148 (O_148,N_4006,N_4231);
nand UO_149 (O_149,N_4854,N_4153);
or UO_150 (O_150,N_4431,N_4799);
nor UO_151 (O_151,N_4345,N_4329);
and UO_152 (O_152,N_4734,N_4442);
or UO_153 (O_153,N_4210,N_4266);
or UO_154 (O_154,N_4245,N_4766);
or UO_155 (O_155,N_4744,N_4142);
or UO_156 (O_156,N_4765,N_4059);
and UO_157 (O_157,N_4197,N_4707);
nand UO_158 (O_158,N_4830,N_4670);
and UO_159 (O_159,N_4179,N_4216);
or UO_160 (O_160,N_4189,N_4167);
or UO_161 (O_161,N_4589,N_4284);
or UO_162 (O_162,N_4904,N_4494);
xnor UO_163 (O_163,N_4012,N_4607);
or UO_164 (O_164,N_4862,N_4988);
and UO_165 (O_165,N_4499,N_4724);
and UO_166 (O_166,N_4044,N_4460);
or UO_167 (O_167,N_4486,N_4516);
and UO_168 (O_168,N_4346,N_4936);
or UO_169 (O_169,N_4204,N_4926);
nand UO_170 (O_170,N_4290,N_4367);
xnor UO_171 (O_171,N_4865,N_4118);
and UO_172 (O_172,N_4969,N_4301);
or UO_173 (O_173,N_4548,N_4203);
or UO_174 (O_174,N_4685,N_4298);
nand UO_175 (O_175,N_4721,N_4228);
nor UO_176 (O_176,N_4600,N_4889);
nand UO_177 (O_177,N_4035,N_4045);
or UO_178 (O_178,N_4382,N_4038);
xor UO_179 (O_179,N_4691,N_4334);
or UO_180 (O_180,N_4677,N_4689);
or UO_181 (O_181,N_4745,N_4750);
or UO_182 (O_182,N_4876,N_4428);
nor UO_183 (O_183,N_4086,N_4069);
and UO_184 (O_184,N_4958,N_4106);
nand UO_185 (O_185,N_4159,N_4360);
and UO_186 (O_186,N_4676,N_4528);
nand UO_187 (O_187,N_4836,N_4649);
nor UO_188 (O_188,N_4183,N_4276);
and UO_189 (O_189,N_4024,N_4875);
and UO_190 (O_190,N_4594,N_4572);
and UO_191 (O_191,N_4560,N_4942);
or UO_192 (O_192,N_4717,N_4444);
and UO_193 (O_193,N_4190,N_4134);
nand UO_194 (O_194,N_4934,N_4532);
or UO_195 (O_195,N_4775,N_4874);
or UO_196 (O_196,N_4472,N_4643);
nand UO_197 (O_197,N_4666,N_4481);
nor UO_198 (O_198,N_4155,N_4586);
or UO_199 (O_199,N_4490,N_4651);
nand UO_200 (O_200,N_4454,N_4125);
nor UO_201 (O_201,N_4263,N_4340);
and UO_202 (O_202,N_4638,N_4652);
and UO_203 (O_203,N_4380,N_4778);
or UO_204 (O_204,N_4316,N_4406);
nand UO_205 (O_205,N_4470,N_4253);
nor UO_206 (O_206,N_4171,N_4262);
and UO_207 (O_207,N_4780,N_4679);
and UO_208 (O_208,N_4361,N_4434);
nor UO_209 (O_209,N_4879,N_4686);
nand UO_210 (O_210,N_4050,N_4993);
and UO_211 (O_211,N_4937,N_4071);
xor UO_212 (O_212,N_4569,N_4551);
and UO_213 (O_213,N_4392,N_4184);
or UO_214 (O_214,N_4043,N_4795);
or UO_215 (O_215,N_4849,N_4832);
nor UO_216 (O_216,N_4185,N_4343);
xor UO_217 (O_217,N_4229,N_4278);
nand UO_218 (O_218,N_4508,N_4100);
or UO_219 (O_219,N_4188,N_4577);
or UO_220 (O_220,N_4140,N_4386);
nor UO_221 (O_221,N_4450,N_4500);
nor UO_222 (O_222,N_4935,N_4039);
nor UO_223 (O_223,N_4277,N_4732);
nor UO_224 (O_224,N_4986,N_4256);
and UO_225 (O_225,N_4640,N_4384);
or UO_226 (O_226,N_4422,N_4729);
and UO_227 (O_227,N_4198,N_4207);
and UO_228 (O_228,N_4574,N_4822);
nand UO_229 (O_229,N_4233,N_4624);
and UO_230 (O_230,N_4236,N_4356);
and UO_231 (O_231,N_4549,N_4909);
and UO_232 (O_232,N_4187,N_4254);
nor UO_233 (O_233,N_4535,N_4597);
and UO_234 (O_234,N_4796,N_4036);
nor UO_235 (O_235,N_4124,N_4149);
nand UO_236 (O_236,N_4128,N_4344);
and UO_237 (O_237,N_4014,N_4702);
nand UO_238 (O_238,N_4695,N_4896);
nor UO_239 (O_239,N_4475,N_4293);
nor UO_240 (O_240,N_4657,N_4787);
or UO_241 (O_241,N_4068,N_4720);
and UO_242 (O_242,N_4057,N_4755);
or UO_243 (O_243,N_4659,N_4716);
and UO_244 (O_244,N_4561,N_4871);
nand UO_245 (O_245,N_4425,N_4928);
or UO_246 (O_246,N_4852,N_4303);
nor UO_247 (O_247,N_4078,N_4180);
nand UO_248 (O_248,N_4021,N_4816);
or UO_249 (O_249,N_4992,N_4404);
nand UO_250 (O_250,N_4342,N_4008);
or UO_251 (O_251,N_4618,N_4056);
or UO_252 (O_252,N_4097,N_4312);
nor UO_253 (O_253,N_4636,N_4982);
nand UO_254 (O_254,N_4898,N_4000);
nor UO_255 (O_255,N_4283,N_4381);
or UO_256 (O_256,N_4582,N_4137);
or UO_257 (O_257,N_4553,N_4631);
nand UO_258 (O_258,N_4333,N_4803);
nand UO_259 (O_259,N_4602,N_4366);
and UO_260 (O_260,N_4825,N_4980);
nor UO_261 (O_261,N_4217,N_4983);
nor UO_262 (O_262,N_4921,N_4949);
or UO_263 (O_263,N_4540,N_4987);
and UO_264 (O_264,N_4003,N_4440);
nand UO_265 (O_265,N_4674,N_4025);
nor UO_266 (O_266,N_4842,N_4529);
nand UO_267 (O_267,N_4471,N_4850);
nand UO_268 (O_268,N_4855,N_4916);
nor UO_269 (O_269,N_4029,N_4347);
and UO_270 (O_270,N_4145,N_4075);
and UO_271 (O_271,N_4869,N_4927);
and UO_272 (O_272,N_4596,N_4870);
nand UO_273 (O_273,N_4289,N_4241);
nor UO_274 (O_274,N_4793,N_4336);
and UO_275 (O_275,N_4839,N_4943);
nor UO_276 (O_276,N_4350,N_4327);
nor UO_277 (O_277,N_4445,N_4274);
nor UO_278 (O_278,N_4115,N_4843);
xnor UO_279 (O_279,N_4511,N_4095);
and UO_280 (O_280,N_4890,N_4201);
or UO_281 (O_281,N_4806,N_4453);
nor UO_282 (O_282,N_4584,N_4265);
nand UO_283 (O_283,N_4359,N_4999);
or UO_284 (O_284,N_4430,N_4951);
nand UO_285 (O_285,N_4101,N_4546);
or UO_286 (O_286,N_4332,N_4170);
nor UO_287 (O_287,N_4441,N_4568);
nand UO_288 (O_288,N_4252,N_4995);
or UO_289 (O_289,N_4209,N_4157);
or UO_290 (O_290,N_4130,N_4258);
and UO_291 (O_291,N_4519,N_4785);
nand UO_292 (O_292,N_4534,N_4143);
nand UO_293 (O_293,N_4084,N_4894);
nor UO_294 (O_294,N_4432,N_4856);
and UO_295 (O_295,N_4223,N_4847);
nor UO_296 (O_296,N_4911,N_4733);
nand UO_297 (O_297,N_4311,N_4436);
or UO_298 (O_298,N_4320,N_4712);
nor UO_299 (O_299,N_4325,N_4348);
or UO_300 (O_300,N_4531,N_4452);
nand UO_301 (O_301,N_4234,N_4338);
nor UO_302 (O_302,N_4813,N_4358);
nor UO_303 (O_303,N_4317,N_4845);
and UO_304 (O_304,N_4105,N_4735);
nand UO_305 (O_305,N_4736,N_4562);
and UO_306 (O_306,N_4777,N_4341);
nand UO_307 (O_307,N_4851,N_4178);
and UO_308 (O_308,N_4395,N_4998);
xnor UO_309 (O_309,N_4004,N_4573);
or UO_310 (O_310,N_4091,N_4972);
xnor UO_311 (O_311,N_4761,N_4049);
and UO_312 (O_312,N_4053,N_4808);
nor UO_313 (O_313,N_4858,N_4575);
nor UO_314 (O_314,N_4030,N_4515);
or UO_315 (O_315,N_4931,N_4074);
or UO_316 (O_316,N_4052,N_4645);
nor UO_317 (O_317,N_4633,N_4559);
or UO_318 (O_318,N_4513,N_4647);
and UO_319 (O_319,N_4605,N_4818);
nor UO_320 (O_320,N_4524,N_4214);
or UO_321 (O_321,N_4215,N_4117);
nand UO_322 (O_322,N_4622,N_4061);
nor UO_323 (O_323,N_4459,N_4833);
and UO_324 (O_324,N_4681,N_4261);
or UO_325 (O_325,N_4558,N_4487);
nor UO_326 (O_326,N_4979,N_4505);
or UO_327 (O_327,N_4482,N_4133);
and UO_328 (O_328,N_4318,N_4375);
nor UO_329 (O_329,N_4841,N_4975);
and UO_330 (O_330,N_4800,N_4389);
nor UO_331 (O_331,N_4089,N_4718);
or UO_332 (O_332,N_4947,N_4634);
and UO_333 (O_333,N_4526,N_4722);
nand UO_334 (O_334,N_4920,N_4706);
nand UO_335 (O_335,N_4426,N_4616);
nor UO_336 (O_336,N_4873,N_4598);
nor UO_337 (O_337,N_4814,N_4655);
nand UO_338 (O_338,N_4407,N_4268);
nand UO_339 (O_339,N_4151,N_4398);
and UO_340 (O_340,N_4081,N_4587);
and UO_341 (O_341,N_4269,N_4779);
nor UO_342 (O_342,N_4109,N_4715);
nor UO_343 (O_343,N_4520,N_4828);
or UO_344 (O_344,N_4108,N_4881);
and UO_345 (O_345,N_4791,N_4365);
or UO_346 (O_346,N_4682,N_4166);
xnor UO_347 (O_347,N_4016,N_4427);
and UO_348 (O_348,N_4139,N_4663);
nand UO_349 (O_349,N_4379,N_4270);
nand UO_350 (O_350,N_4965,N_4701);
xor UO_351 (O_351,N_4222,N_4458);
nand UO_352 (O_352,N_4709,N_4807);
or UO_353 (O_353,N_4042,N_4897);
and UO_354 (O_354,N_4853,N_4421);
xor UO_355 (O_355,N_4948,N_4403);
nor UO_356 (O_356,N_4193,N_4687);
nor UO_357 (O_357,N_4692,N_4571);
or UO_358 (O_358,N_4113,N_4743);
and UO_359 (O_359,N_4121,N_4279);
nor UO_360 (O_360,N_4697,N_4901);
and UO_361 (O_361,N_4390,N_4251);
and UO_362 (O_362,N_4754,N_4521);
and UO_363 (O_363,N_4699,N_4067);
nor UO_364 (O_364,N_4369,N_4829);
nor UO_365 (O_365,N_4737,N_4054);
nand UO_366 (O_366,N_4399,N_4710);
nand UO_367 (O_367,N_4195,N_4579);
or UO_368 (O_368,N_4502,N_4328);
or UO_369 (O_369,N_4135,N_4860);
or UO_370 (O_370,N_4493,N_4671);
nor UO_371 (O_371,N_4617,N_4639);
and UO_372 (O_372,N_4981,N_4169);
or UO_373 (O_373,N_4377,N_4543);
nor UO_374 (O_374,N_4098,N_4032);
or UO_375 (O_375,N_4026,N_4557);
and UO_376 (O_376,N_4250,N_4518);
nand UO_377 (O_377,N_4667,N_4443);
and UO_378 (O_378,N_4249,N_4259);
nor UO_379 (O_379,N_4467,N_4891);
or UO_380 (O_380,N_4815,N_4271);
or UO_381 (O_381,N_4176,N_4103);
and UO_382 (O_382,N_4510,N_4387);
and UO_383 (O_383,N_4285,N_4173);
and UO_384 (O_384,N_4971,N_4294);
nor UO_385 (O_385,N_4243,N_4673);
nand UO_386 (O_386,N_4725,N_4933);
or UO_387 (O_387,N_4968,N_4168);
and UO_388 (O_388,N_4821,N_4401);
or UO_389 (O_389,N_4626,N_4186);
nand UO_390 (O_390,N_4536,N_4653);
nand UO_391 (O_391,N_4684,N_4033);
nor UO_392 (O_392,N_4181,N_4503);
and UO_393 (O_393,N_4929,N_4959);
nor UO_394 (O_394,N_4397,N_4882);
and UO_395 (O_395,N_4824,N_4917);
nand UO_396 (O_396,N_4488,N_4581);
or UO_397 (O_397,N_4903,N_4797);
or UO_398 (O_398,N_4899,N_4556);
nor UO_399 (O_399,N_4984,N_4661);
nor UO_400 (O_400,N_4885,N_4703);
nor UO_401 (O_401,N_4092,N_4542);
or UO_402 (O_402,N_4048,N_4805);
and UO_403 (O_403,N_4576,N_4018);
nor UO_404 (O_404,N_4835,N_4621);
nor UO_405 (O_405,N_4309,N_4658);
and UO_406 (O_406,N_4861,N_4599);
and UO_407 (O_407,N_4629,N_4683);
nand UO_408 (O_408,N_4788,N_4093);
or UO_409 (O_409,N_4065,N_4539);
xnor UO_410 (O_410,N_4468,N_4554);
or UO_411 (O_411,N_4212,N_4146);
or UO_412 (O_412,N_4878,N_4859);
and UO_413 (O_413,N_4070,N_4804);
nand UO_414 (O_414,N_4838,N_4447);
nand UO_415 (O_415,N_4809,N_4364);
nand UO_416 (O_416,N_4492,N_4001);
nand UO_417 (O_417,N_4150,N_4010);
or UO_418 (O_418,N_4900,N_4801);
or UO_419 (O_419,N_4530,N_4678);
nand UO_420 (O_420,N_4225,N_4304);
nand UO_421 (O_421,N_4585,N_4783);
or UO_422 (O_422,N_4307,N_4162);
or UO_423 (O_423,N_4698,N_4372);
nand UO_424 (O_424,N_4957,N_4246);
or UO_425 (O_425,N_4022,N_4739);
nand UO_426 (O_426,N_4424,N_4764);
or UO_427 (O_427,N_4726,N_4672);
or UO_428 (O_428,N_4538,N_4055);
nor UO_429 (O_429,N_4590,N_4772);
and UO_430 (O_430,N_4409,N_4632);
or UO_431 (O_431,N_4625,N_4126);
nand UO_432 (O_432,N_4660,N_4844);
nor UO_433 (O_433,N_4786,N_4665);
or UO_434 (O_434,N_4282,N_4154);
and UO_435 (O_435,N_4713,N_4239);
or UO_436 (O_436,N_4286,N_4267);
nand UO_437 (O_437,N_4525,N_4211);
or UO_438 (O_438,N_4378,N_4945);
nand UO_439 (O_439,N_4357,N_4642);
nand UO_440 (O_440,N_4595,N_4863);
and UO_441 (O_441,N_4727,N_4680);
nand UO_442 (O_442,N_4072,N_4664);
and UO_443 (O_443,N_4355,N_4083);
or UO_444 (O_444,N_4823,N_4077);
and UO_445 (O_445,N_4628,N_4058);
and UO_446 (O_446,N_4335,N_4892);
and UO_447 (O_447,N_4219,N_4297);
and UO_448 (O_448,N_4913,N_4464);
nand UO_449 (O_449,N_4013,N_4939);
and UO_450 (O_450,N_4545,N_4227);
or UO_451 (O_451,N_4122,N_4826);
and UO_452 (O_452,N_4161,N_4119);
and UO_453 (O_453,N_4047,N_4076);
nor UO_454 (O_454,N_4244,N_4762);
or UO_455 (O_455,N_4172,N_4973);
nand UO_456 (O_456,N_4177,N_4363);
or UO_457 (O_457,N_4550,N_4374);
nand UO_458 (O_458,N_4037,N_4753);
or UO_459 (O_459,N_4714,N_4415);
nor UO_460 (O_460,N_4473,N_4174);
or UO_461 (O_461,N_4802,N_4175);
or UO_462 (O_462,N_4566,N_4646);
xor UO_463 (O_463,N_4517,N_4489);
and UO_464 (O_464,N_4411,N_4015);
and UO_465 (O_465,N_4144,N_4976);
nand UO_466 (O_466,N_4547,N_4669);
nand UO_467 (O_467,N_4564,N_4902);
nor UO_468 (O_468,N_4046,N_4583);
and UO_469 (O_469,N_4264,N_4051);
and UO_470 (O_470,N_4749,N_4152);
nor UO_471 (O_471,N_4533,N_4944);
nor UO_472 (O_472,N_4230,N_4789);
nand UO_473 (O_473,N_4080,N_4349);
nor UO_474 (O_474,N_4235,N_4497);
nand UO_475 (O_475,N_4136,N_4476);
nand UO_476 (O_476,N_4331,N_4819);
and UO_477 (O_477,N_4321,N_4767);
and UO_478 (O_478,N_4090,N_4408);
nor UO_479 (O_479,N_4085,N_4064);
and UO_480 (O_480,N_4644,N_4930);
and UO_481 (O_481,N_4218,N_4305);
nand UO_482 (O_482,N_4376,N_4040);
nor UO_483 (O_483,N_4405,N_4527);
or UO_484 (O_484,N_4523,N_4756);
nor UO_485 (O_485,N_4728,N_4696);
or UO_486 (O_486,N_4087,N_4817);
or UO_487 (O_487,N_4504,N_4129);
or UO_488 (O_488,N_4023,N_4507);
and UO_489 (O_489,N_4941,N_4391);
and UO_490 (O_490,N_4213,N_4752);
nand UO_491 (O_491,N_4996,N_4275);
nand UO_492 (O_492,N_4932,N_4031);
nor UO_493 (O_493,N_4088,N_4158);
nor UO_494 (O_494,N_4544,N_4769);
or UO_495 (O_495,N_4132,N_4410);
or UO_496 (O_496,N_4740,N_4966);
nor UO_497 (O_497,N_4541,N_4552);
and UO_498 (O_498,N_4623,N_4308);
nand UO_499 (O_499,N_4846,N_4914);
and UO_500 (O_500,N_4680,N_4684);
nor UO_501 (O_501,N_4738,N_4482);
and UO_502 (O_502,N_4776,N_4570);
nand UO_503 (O_503,N_4115,N_4106);
and UO_504 (O_504,N_4686,N_4656);
or UO_505 (O_505,N_4807,N_4170);
nand UO_506 (O_506,N_4840,N_4544);
nor UO_507 (O_507,N_4482,N_4790);
and UO_508 (O_508,N_4697,N_4124);
nand UO_509 (O_509,N_4637,N_4874);
or UO_510 (O_510,N_4611,N_4403);
nand UO_511 (O_511,N_4312,N_4218);
nand UO_512 (O_512,N_4495,N_4674);
or UO_513 (O_513,N_4939,N_4948);
nand UO_514 (O_514,N_4985,N_4019);
nand UO_515 (O_515,N_4892,N_4116);
nand UO_516 (O_516,N_4543,N_4846);
and UO_517 (O_517,N_4966,N_4340);
nand UO_518 (O_518,N_4898,N_4400);
and UO_519 (O_519,N_4928,N_4470);
nor UO_520 (O_520,N_4349,N_4932);
and UO_521 (O_521,N_4514,N_4878);
or UO_522 (O_522,N_4041,N_4000);
and UO_523 (O_523,N_4418,N_4249);
nor UO_524 (O_524,N_4680,N_4153);
nor UO_525 (O_525,N_4380,N_4709);
nor UO_526 (O_526,N_4482,N_4094);
nor UO_527 (O_527,N_4719,N_4272);
and UO_528 (O_528,N_4618,N_4846);
or UO_529 (O_529,N_4182,N_4003);
and UO_530 (O_530,N_4564,N_4188);
and UO_531 (O_531,N_4729,N_4295);
nor UO_532 (O_532,N_4358,N_4324);
and UO_533 (O_533,N_4767,N_4184);
nand UO_534 (O_534,N_4688,N_4435);
and UO_535 (O_535,N_4546,N_4704);
nand UO_536 (O_536,N_4643,N_4666);
nor UO_537 (O_537,N_4972,N_4279);
and UO_538 (O_538,N_4365,N_4287);
nor UO_539 (O_539,N_4955,N_4529);
and UO_540 (O_540,N_4924,N_4384);
nor UO_541 (O_541,N_4127,N_4029);
or UO_542 (O_542,N_4279,N_4932);
or UO_543 (O_543,N_4370,N_4474);
nor UO_544 (O_544,N_4263,N_4014);
or UO_545 (O_545,N_4932,N_4351);
nor UO_546 (O_546,N_4696,N_4763);
nor UO_547 (O_547,N_4963,N_4888);
and UO_548 (O_548,N_4749,N_4172);
and UO_549 (O_549,N_4567,N_4077);
nor UO_550 (O_550,N_4282,N_4015);
xnor UO_551 (O_551,N_4792,N_4449);
nor UO_552 (O_552,N_4486,N_4041);
nor UO_553 (O_553,N_4617,N_4989);
and UO_554 (O_554,N_4845,N_4351);
nor UO_555 (O_555,N_4034,N_4095);
nand UO_556 (O_556,N_4626,N_4517);
nand UO_557 (O_557,N_4777,N_4216);
nand UO_558 (O_558,N_4602,N_4627);
and UO_559 (O_559,N_4740,N_4245);
and UO_560 (O_560,N_4847,N_4242);
or UO_561 (O_561,N_4163,N_4210);
and UO_562 (O_562,N_4150,N_4337);
or UO_563 (O_563,N_4317,N_4135);
nor UO_564 (O_564,N_4941,N_4226);
nor UO_565 (O_565,N_4534,N_4461);
and UO_566 (O_566,N_4317,N_4754);
or UO_567 (O_567,N_4213,N_4715);
or UO_568 (O_568,N_4902,N_4822);
nor UO_569 (O_569,N_4083,N_4097);
and UO_570 (O_570,N_4246,N_4670);
nand UO_571 (O_571,N_4580,N_4091);
nor UO_572 (O_572,N_4560,N_4268);
nor UO_573 (O_573,N_4506,N_4580);
or UO_574 (O_574,N_4645,N_4341);
nand UO_575 (O_575,N_4475,N_4633);
nand UO_576 (O_576,N_4957,N_4980);
nor UO_577 (O_577,N_4440,N_4778);
nand UO_578 (O_578,N_4845,N_4303);
xnor UO_579 (O_579,N_4127,N_4860);
nor UO_580 (O_580,N_4245,N_4089);
nand UO_581 (O_581,N_4603,N_4884);
nand UO_582 (O_582,N_4372,N_4699);
nand UO_583 (O_583,N_4407,N_4976);
nand UO_584 (O_584,N_4667,N_4717);
and UO_585 (O_585,N_4122,N_4231);
and UO_586 (O_586,N_4068,N_4628);
nor UO_587 (O_587,N_4566,N_4930);
nand UO_588 (O_588,N_4926,N_4670);
and UO_589 (O_589,N_4654,N_4217);
or UO_590 (O_590,N_4468,N_4376);
nor UO_591 (O_591,N_4738,N_4206);
nand UO_592 (O_592,N_4302,N_4584);
and UO_593 (O_593,N_4894,N_4473);
xor UO_594 (O_594,N_4407,N_4631);
xor UO_595 (O_595,N_4685,N_4866);
nand UO_596 (O_596,N_4437,N_4416);
or UO_597 (O_597,N_4396,N_4146);
nor UO_598 (O_598,N_4081,N_4483);
and UO_599 (O_599,N_4427,N_4126);
xnor UO_600 (O_600,N_4702,N_4063);
nor UO_601 (O_601,N_4481,N_4397);
nand UO_602 (O_602,N_4444,N_4258);
and UO_603 (O_603,N_4058,N_4957);
or UO_604 (O_604,N_4347,N_4513);
or UO_605 (O_605,N_4502,N_4778);
nor UO_606 (O_606,N_4611,N_4365);
and UO_607 (O_607,N_4924,N_4529);
nand UO_608 (O_608,N_4948,N_4958);
nor UO_609 (O_609,N_4861,N_4822);
nor UO_610 (O_610,N_4193,N_4379);
or UO_611 (O_611,N_4634,N_4544);
and UO_612 (O_612,N_4821,N_4956);
xor UO_613 (O_613,N_4827,N_4112);
and UO_614 (O_614,N_4175,N_4530);
nor UO_615 (O_615,N_4035,N_4596);
and UO_616 (O_616,N_4573,N_4565);
nor UO_617 (O_617,N_4616,N_4524);
nand UO_618 (O_618,N_4878,N_4208);
and UO_619 (O_619,N_4880,N_4108);
and UO_620 (O_620,N_4920,N_4077);
nand UO_621 (O_621,N_4925,N_4147);
and UO_622 (O_622,N_4753,N_4334);
nor UO_623 (O_623,N_4241,N_4532);
xor UO_624 (O_624,N_4527,N_4996);
xnor UO_625 (O_625,N_4337,N_4932);
xnor UO_626 (O_626,N_4074,N_4070);
and UO_627 (O_627,N_4259,N_4715);
nand UO_628 (O_628,N_4246,N_4242);
nand UO_629 (O_629,N_4992,N_4415);
nor UO_630 (O_630,N_4273,N_4004);
or UO_631 (O_631,N_4976,N_4575);
and UO_632 (O_632,N_4994,N_4168);
or UO_633 (O_633,N_4464,N_4223);
and UO_634 (O_634,N_4636,N_4927);
xnor UO_635 (O_635,N_4355,N_4787);
nand UO_636 (O_636,N_4774,N_4790);
nand UO_637 (O_637,N_4599,N_4786);
or UO_638 (O_638,N_4581,N_4853);
nand UO_639 (O_639,N_4869,N_4735);
nand UO_640 (O_640,N_4608,N_4773);
and UO_641 (O_641,N_4807,N_4087);
and UO_642 (O_642,N_4369,N_4931);
nor UO_643 (O_643,N_4507,N_4225);
and UO_644 (O_644,N_4374,N_4963);
nand UO_645 (O_645,N_4135,N_4912);
and UO_646 (O_646,N_4917,N_4894);
nand UO_647 (O_647,N_4115,N_4834);
and UO_648 (O_648,N_4622,N_4410);
nand UO_649 (O_649,N_4265,N_4764);
nor UO_650 (O_650,N_4013,N_4623);
or UO_651 (O_651,N_4566,N_4126);
nor UO_652 (O_652,N_4146,N_4361);
xnor UO_653 (O_653,N_4363,N_4130);
nand UO_654 (O_654,N_4975,N_4840);
and UO_655 (O_655,N_4843,N_4786);
and UO_656 (O_656,N_4380,N_4023);
nand UO_657 (O_657,N_4329,N_4171);
nor UO_658 (O_658,N_4793,N_4007);
nand UO_659 (O_659,N_4550,N_4412);
and UO_660 (O_660,N_4758,N_4431);
nand UO_661 (O_661,N_4986,N_4331);
nor UO_662 (O_662,N_4967,N_4537);
or UO_663 (O_663,N_4281,N_4096);
and UO_664 (O_664,N_4310,N_4962);
nor UO_665 (O_665,N_4288,N_4275);
or UO_666 (O_666,N_4529,N_4216);
nor UO_667 (O_667,N_4727,N_4484);
nand UO_668 (O_668,N_4474,N_4094);
or UO_669 (O_669,N_4717,N_4453);
nand UO_670 (O_670,N_4523,N_4596);
nand UO_671 (O_671,N_4462,N_4455);
nand UO_672 (O_672,N_4664,N_4108);
and UO_673 (O_673,N_4237,N_4052);
nand UO_674 (O_674,N_4625,N_4421);
or UO_675 (O_675,N_4298,N_4234);
nor UO_676 (O_676,N_4257,N_4073);
or UO_677 (O_677,N_4944,N_4585);
nand UO_678 (O_678,N_4058,N_4453);
or UO_679 (O_679,N_4969,N_4872);
nor UO_680 (O_680,N_4404,N_4555);
nand UO_681 (O_681,N_4074,N_4292);
and UO_682 (O_682,N_4479,N_4141);
nand UO_683 (O_683,N_4598,N_4688);
or UO_684 (O_684,N_4470,N_4971);
or UO_685 (O_685,N_4107,N_4230);
nor UO_686 (O_686,N_4651,N_4883);
nand UO_687 (O_687,N_4004,N_4319);
nor UO_688 (O_688,N_4931,N_4508);
nor UO_689 (O_689,N_4414,N_4707);
nor UO_690 (O_690,N_4943,N_4571);
nand UO_691 (O_691,N_4503,N_4364);
or UO_692 (O_692,N_4950,N_4219);
nor UO_693 (O_693,N_4714,N_4874);
and UO_694 (O_694,N_4562,N_4415);
and UO_695 (O_695,N_4407,N_4899);
or UO_696 (O_696,N_4255,N_4630);
and UO_697 (O_697,N_4953,N_4766);
and UO_698 (O_698,N_4018,N_4805);
or UO_699 (O_699,N_4902,N_4047);
nor UO_700 (O_700,N_4995,N_4795);
nand UO_701 (O_701,N_4478,N_4900);
and UO_702 (O_702,N_4280,N_4079);
nor UO_703 (O_703,N_4922,N_4288);
nor UO_704 (O_704,N_4668,N_4947);
and UO_705 (O_705,N_4608,N_4613);
nor UO_706 (O_706,N_4799,N_4783);
nor UO_707 (O_707,N_4509,N_4626);
nor UO_708 (O_708,N_4710,N_4920);
nand UO_709 (O_709,N_4379,N_4609);
nand UO_710 (O_710,N_4911,N_4141);
and UO_711 (O_711,N_4473,N_4731);
and UO_712 (O_712,N_4499,N_4457);
or UO_713 (O_713,N_4470,N_4478);
and UO_714 (O_714,N_4995,N_4984);
nand UO_715 (O_715,N_4822,N_4166);
or UO_716 (O_716,N_4299,N_4782);
and UO_717 (O_717,N_4841,N_4210);
or UO_718 (O_718,N_4634,N_4007);
or UO_719 (O_719,N_4569,N_4579);
and UO_720 (O_720,N_4725,N_4184);
and UO_721 (O_721,N_4867,N_4335);
and UO_722 (O_722,N_4155,N_4595);
and UO_723 (O_723,N_4326,N_4877);
and UO_724 (O_724,N_4279,N_4366);
and UO_725 (O_725,N_4786,N_4893);
nand UO_726 (O_726,N_4383,N_4507);
or UO_727 (O_727,N_4937,N_4997);
nand UO_728 (O_728,N_4025,N_4087);
or UO_729 (O_729,N_4189,N_4842);
nor UO_730 (O_730,N_4980,N_4994);
and UO_731 (O_731,N_4455,N_4498);
and UO_732 (O_732,N_4689,N_4224);
and UO_733 (O_733,N_4056,N_4280);
nor UO_734 (O_734,N_4681,N_4495);
nor UO_735 (O_735,N_4821,N_4913);
or UO_736 (O_736,N_4171,N_4020);
or UO_737 (O_737,N_4134,N_4728);
and UO_738 (O_738,N_4615,N_4941);
nor UO_739 (O_739,N_4177,N_4151);
or UO_740 (O_740,N_4932,N_4161);
and UO_741 (O_741,N_4695,N_4402);
nand UO_742 (O_742,N_4966,N_4370);
and UO_743 (O_743,N_4259,N_4413);
nand UO_744 (O_744,N_4865,N_4438);
nor UO_745 (O_745,N_4296,N_4104);
nand UO_746 (O_746,N_4849,N_4021);
or UO_747 (O_747,N_4871,N_4949);
or UO_748 (O_748,N_4693,N_4678);
nand UO_749 (O_749,N_4479,N_4269);
and UO_750 (O_750,N_4903,N_4007);
or UO_751 (O_751,N_4788,N_4935);
nand UO_752 (O_752,N_4908,N_4711);
or UO_753 (O_753,N_4566,N_4829);
nand UO_754 (O_754,N_4353,N_4864);
nand UO_755 (O_755,N_4010,N_4209);
or UO_756 (O_756,N_4498,N_4935);
and UO_757 (O_757,N_4553,N_4166);
nand UO_758 (O_758,N_4466,N_4168);
nand UO_759 (O_759,N_4315,N_4300);
nor UO_760 (O_760,N_4758,N_4039);
nand UO_761 (O_761,N_4606,N_4893);
and UO_762 (O_762,N_4338,N_4658);
nand UO_763 (O_763,N_4436,N_4112);
and UO_764 (O_764,N_4866,N_4698);
nor UO_765 (O_765,N_4757,N_4827);
or UO_766 (O_766,N_4542,N_4086);
or UO_767 (O_767,N_4826,N_4724);
and UO_768 (O_768,N_4471,N_4860);
and UO_769 (O_769,N_4721,N_4536);
and UO_770 (O_770,N_4466,N_4107);
or UO_771 (O_771,N_4532,N_4700);
and UO_772 (O_772,N_4508,N_4780);
and UO_773 (O_773,N_4344,N_4857);
or UO_774 (O_774,N_4931,N_4269);
and UO_775 (O_775,N_4013,N_4456);
and UO_776 (O_776,N_4881,N_4947);
or UO_777 (O_777,N_4866,N_4760);
or UO_778 (O_778,N_4487,N_4238);
and UO_779 (O_779,N_4298,N_4360);
nand UO_780 (O_780,N_4092,N_4577);
nor UO_781 (O_781,N_4082,N_4665);
and UO_782 (O_782,N_4949,N_4387);
nor UO_783 (O_783,N_4841,N_4823);
and UO_784 (O_784,N_4990,N_4702);
nand UO_785 (O_785,N_4866,N_4396);
or UO_786 (O_786,N_4698,N_4299);
nor UO_787 (O_787,N_4716,N_4857);
or UO_788 (O_788,N_4345,N_4069);
nand UO_789 (O_789,N_4222,N_4860);
nand UO_790 (O_790,N_4333,N_4337);
and UO_791 (O_791,N_4955,N_4316);
or UO_792 (O_792,N_4802,N_4914);
nor UO_793 (O_793,N_4346,N_4756);
and UO_794 (O_794,N_4360,N_4632);
and UO_795 (O_795,N_4940,N_4546);
nor UO_796 (O_796,N_4155,N_4946);
nor UO_797 (O_797,N_4873,N_4379);
and UO_798 (O_798,N_4204,N_4674);
or UO_799 (O_799,N_4401,N_4429);
nor UO_800 (O_800,N_4933,N_4294);
or UO_801 (O_801,N_4505,N_4813);
nor UO_802 (O_802,N_4937,N_4569);
xor UO_803 (O_803,N_4725,N_4462);
nand UO_804 (O_804,N_4556,N_4851);
or UO_805 (O_805,N_4709,N_4799);
and UO_806 (O_806,N_4878,N_4305);
or UO_807 (O_807,N_4338,N_4486);
and UO_808 (O_808,N_4134,N_4983);
nand UO_809 (O_809,N_4597,N_4322);
nand UO_810 (O_810,N_4337,N_4809);
nor UO_811 (O_811,N_4154,N_4956);
nor UO_812 (O_812,N_4890,N_4120);
nand UO_813 (O_813,N_4897,N_4774);
or UO_814 (O_814,N_4704,N_4448);
nand UO_815 (O_815,N_4194,N_4859);
and UO_816 (O_816,N_4617,N_4518);
nand UO_817 (O_817,N_4364,N_4859);
and UO_818 (O_818,N_4197,N_4094);
or UO_819 (O_819,N_4386,N_4115);
or UO_820 (O_820,N_4959,N_4096);
or UO_821 (O_821,N_4315,N_4948);
nor UO_822 (O_822,N_4196,N_4079);
nand UO_823 (O_823,N_4503,N_4164);
and UO_824 (O_824,N_4445,N_4977);
nand UO_825 (O_825,N_4079,N_4183);
or UO_826 (O_826,N_4802,N_4186);
and UO_827 (O_827,N_4503,N_4672);
or UO_828 (O_828,N_4634,N_4669);
and UO_829 (O_829,N_4124,N_4104);
nor UO_830 (O_830,N_4846,N_4683);
xor UO_831 (O_831,N_4070,N_4115);
or UO_832 (O_832,N_4658,N_4618);
and UO_833 (O_833,N_4024,N_4993);
or UO_834 (O_834,N_4596,N_4285);
or UO_835 (O_835,N_4788,N_4293);
or UO_836 (O_836,N_4695,N_4314);
and UO_837 (O_837,N_4423,N_4499);
nand UO_838 (O_838,N_4617,N_4324);
nand UO_839 (O_839,N_4495,N_4060);
and UO_840 (O_840,N_4269,N_4809);
or UO_841 (O_841,N_4029,N_4878);
or UO_842 (O_842,N_4641,N_4186);
nand UO_843 (O_843,N_4965,N_4714);
and UO_844 (O_844,N_4155,N_4486);
nor UO_845 (O_845,N_4122,N_4336);
nand UO_846 (O_846,N_4477,N_4221);
xor UO_847 (O_847,N_4544,N_4904);
nor UO_848 (O_848,N_4956,N_4331);
and UO_849 (O_849,N_4332,N_4227);
nand UO_850 (O_850,N_4668,N_4828);
and UO_851 (O_851,N_4381,N_4595);
nand UO_852 (O_852,N_4235,N_4291);
nand UO_853 (O_853,N_4785,N_4411);
and UO_854 (O_854,N_4053,N_4878);
nand UO_855 (O_855,N_4917,N_4854);
and UO_856 (O_856,N_4855,N_4447);
nor UO_857 (O_857,N_4301,N_4160);
nor UO_858 (O_858,N_4580,N_4386);
nand UO_859 (O_859,N_4493,N_4112);
nor UO_860 (O_860,N_4833,N_4370);
or UO_861 (O_861,N_4291,N_4991);
nor UO_862 (O_862,N_4175,N_4882);
or UO_863 (O_863,N_4028,N_4725);
nand UO_864 (O_864,N_4236,N_4262);
nand UO_865 (O_865,N_4666,N_4590);
or UO_866 (O_866,N_4747,N_4612);
nand UO_867 (O_867,N_4191,N_4489);
nand UO_868 (O_868,N_4566,N_4975);
or UO_869 (O_869,N_4185,N_4100);
nand UO_870 (O_870,N_4925,N_4776);
nand UO_871 (O_871,N_4257,N_4325);
and UO_872 (O_872,N_4205,N_4492);
and UO_873 (O_873,N_4143,N_4855);
nand UO_874 (O_874,N_4560,N_4259);
and UO_875 (O_875,N_4336,N_4818);
or UO_876 (O_876,N_4964,N_4663);
nor UO_877 (O_877,N_4146,N_4867);
nor UO_878 (O_878,N_4819,N_4496);
or UO_879 (O_879,N_4302,N_4390);
nand UO_880 (O_880,N_4189,N_4100);
nor UO_881 (O_881,N_4263,N_4022);
nor UO_882 (O_882,N_4365,N_4716);
nand UO_883 (O_883,N_4735,N_4935);
or UO_884 (O_884,N_4593,N_4435);
nand UO_885 (O_885,N_4016,N_4261);
or UO_886 (O_886,N_4011,N_4556);
xnor UO_887 (O_887,N_4642,N_4588);
nor UO_888 (O_888,N_4036,N_4965);
and UO_889 (O_889,N_4793,N_4820);
nand UO_890 (O_890,N_4638,N_4859);
nand UO_891 (O_891,N_4131,N_4197);
nor UO_892 (O_892,N_4478,N_4195);
or UO_893 (O_893,N_4821,N_4703);
xor UO_894 (O_894,N_4750,N_4037);
nor UO_895 (O_895,N_4235,N_4212);
or UO_896 (O_896,N_4656,N_4060);
and UO_897 (O_897,N_4438,N_4268);
nand UO_898 (O_898,N_4166,N_4698);
nand UO_899 (O_899,N_4719,N_4287);
nand UO_900 (O_900,N_4884,N_4521);
nor UO_901 (O_901,N_4968,N_4367);
xor UO_902 (O_902,N_4976,N_4310);
nor UO_903 (O_903,N_4317,N_4797);
nand UO_904 (O_904,N_4283,N_4757);
or UO_905 (O_905,N_4921,N_4241);
and UO_906 (O_906,N_4689,N_4682);
or UO_907 (O_907,N_4031,N_4195);
nand UO_908 (O_908,N_4606,N_4200);
nor UO_909 (O_909,N_4019,N_4085);
nor UO_910 (O_910,N_4529,N_4011);
or UO_911 (O_911,N_4402,N_4844);
nor UO_912 (O_912,N_4656,N_4445);
xnor UO_913 (O_913,N_4909,N_4078);
or UO_914 (O_914,N_4151,N_4330);
or UO_915 (O_915,N_4910,N_4890);
or UO_916 (O_916,N_4012,N_4796);
nor UO_917 (O_917,N_4591,N_4854);
nand UO_918 (O_918,N_4129,N_4340);
or UO_919 (O_919,N_4253,N_4145);
and UO_920 (O_920,N_4882,N_4701);
nor UO_921 (O_921,N_4985,N_4493);
or UO_922 (O_922,N_4637,N_4712);
and UO_923 (O_923,N_4428,N_4619);
nor UO_924 (O_924,N_4704,N_4762);
or UO_925 (O_925,N_4032,N_4609);
or UO_926 (O_926,N_4874,N_4744);
nor UO_927 (O_927,N_4560,N_4475);
or UO_928 (O_928,N_4666,N_4152);
nand UO_929 (O_929,N_4121,N_4387);
nand UO_930 (O_930,N_4107,N_4259);
nor UO_931 (O_931,N_4046,N_4037);
or UO_932 (O_932,N_4523,N_4359);
nor UO_933 (O_933,N_4790,N_4656);
nor UO_934 (O_934,N_4021,N_4332);
xnor UO_935 (O_935,N_4694,N_4642);
nor UO_936 (O_936,N_4601,N_4201);
or UO_937 (O_937,N_4673,N_4478);
nor UO_938 (O_938,N_4502,N_4423);
nand UO_939 (O_939,N_4728,N_4717);
xnor UO_940 (O_940,N_4431,N_4003);
nand UO_941 (O_941,N_4266,N_4592);
nand UO_942 (O_942,N_4389,N_4684);
nor UO_943 (O_943,N_4741,N_4214);
or UO_944 (O_944,N_4703,N_4380);
nand UO_945 (O_945,N_4187,N_4431);
or UO_946 (O_946,N_4869,N_4754);
and UO_947 (O_947,N_4860,N_4278);
nand UO_948 (O_948,N_4440,N_4953);
xor UO_949 (O_949,N_4526,N_4130);
nand UO_950 (O_950,N_4173,N_4231);
xnor UO_951 (O_951,N_4312,N_4563);
nor UO_952 (O_952,N_4968,N_4842);
nor UO_953 (O_953,N_4502,N_4819);
nand UO_954 (O_954,N_4905,N_4299);
nand UO_955 (O_955,N_4026,N_4578);
nand UO_956 (O_956,N_4194,N_4078);
nor UO_957 (O_957,N_4429,N_4711);
nand UO_958 (O_958,N_4529,N_4956);
or UO_959 (O_959,N_4729,N_4769);
or UO_960 (O_960,N_4484,N_4697);
xor UO_961 (O_961,N_4268,N_4562);
nor UO_962 (O_962,N_4738,N_4554);
or UO_963 (O_963,N_4877,N_4560);
and UO_964 (O_964,N_4518,N_4419);
nand UO_965 (O_965,N_4607,N_4006);
or UO_966 (O_966,N_4543,N_4513);
and UO_967 (O_967,N_4461,N_4040);
nand UO_968 (O_968,N_4192,N_4828);
nor UO_969 (O_969,N_4852,N_4249);
nor UO_970 (O_970,N_4876,N_4980);
or UO_971 (O_971,N_4739,N_4612);
nand UO_972 (O_972,N_4898,N_4925);
nand UO_973 (O_973,N_4802,N_4439);
nand UO_974 (O_974,N_4764,N_4035);
and UO_975 (O_975,N_4682,N_4345);
and UO_976 (O_976,N_4052,N_4164);
and UO_977 (O_977,N_4035,N_4362);
nor UO_978 (O_978,N_4891,N_4687);
nor UO_979 (O_979,N_4843,N_4994);
or UO_980 (O_980,N_4920,N_4722);
nor UO_981 (O_981,N_4617,N_4353);
or UO_982 (O_982,N_4366,N_4791);
nand UO_983 (O_983,N_4606,N_4790);
nor UO_984 (O_984,N_4857,N_4934);
xor UO_985 (O_985,N_4435,N_4367);
and UO_986 (O_986,N_4997,N_4981);
or UO_987 (O_987,N_4840,N_4972);
or UO_988 (O_988,N_4684,N_4721);
nand UO_989 (O_989,N_4228,N_4778);
nand UO_990 (O_990,N_4916,N_4441);
nand UO_991 (O_991,N_4031,N_4898);
nor UO_992 (O_992,N_4368,N_4323);
or UO_993 (O_993,N_4935,N_4642);
or UO_994 (O_994,N_4648,N_4650);
and UO_995 (O_995,N_4606,N_4684);
xor UO_996 (O_996,N_4270,N_4271);
or UO_997 (O_997,N_4520,N_4395);
or UO_998 (O_998,N_4302,N_4595);
nor UO_999 (O_999,N_4400,N_4890);
endmodule