module basic_500_3000_500_40_levels_1xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
and U0 (N_0,In_404,In_136);
or U1 (N_1,In_383,In_348);
and U2 (N_2,In_426,In_328);
nand U3 (N_3,In_83,In_364);
xor U4 (N_4,In_467,In_266);
xnor U5 (N_5,In_300,In_373);
nor U6 (N_6,In_209,In_332);
nand U7 (N_7,In_156,In_189);
or U8 (N_8,In_476,In_429);
or U9 (N_9,In_427,In_295);
or U10 (N_10,In_66,In_301);
nand U11 (N_11,In_269,In_468);
or U12 (N_12,In_402,In_433);
and U13 (N_13,In_327,In_163);
or U14 (N_14,In_461,In_321);
nor U15 (N_15,In_59,In_56);
and U16 (N_16,In_47,In_244);
and U17 (N_17,In_121,In_462);
nand U18 (N_18,In_202,In_330);
nand U19 (N_19,In_357,In_132);
nor U20 (N_20,In_389,In_148);
nand U21 (N_21,In_331,In_337);
or U22 (N_22,In_343,In_406);
and U23 (N_23,In_256,In_259);
nand U24 (N_24,In_355,In_217);
or U25 (N_25,In_480,In_495);
or U26 (N_26,In_65,In_82);
nand U27 (N_27,In_19,In_214);
or U28 (N_28,In_419,In_274);
nand U29 (N_29,In_395,In_161);
and U30 (N_30,In_282,In_442);
nand U31 (N_31,In_252,In_186);
nand U32 (N_32,In_339,In_428);
or U33 (N_33,In_31,In_104);
nand U34 (N_34,In_175,In_93);
nor U35 (N_35,In_72,In_415);
nand U36 (N_36,In_248,In_469);
nor U37 (N_37,In_306,In_2);
or U38 (N_38,In_483,In_363);
or U39 (N_39,In_127,In_255);
nand U40 (N_40,In_386,In_113);
nand U41 (N_41,In_110,In_228);
nand U42 (N_42,In_422,In_281);
or U43 (N_43,In_216,In_87);
nand U44 (N_44,In_459,In_311);
and U45 (N_45,In_173,In_275);
or U46 (N_46,In_102,In_24);
and U47 (N_47,In_124,In_448);
or U48 (N_48,In_211,In_40);
nor U49 (N_49,In_445,In_184);
and U50 (N_50,In_142,In_400);
nor U51 (N_51,In_162,In_125);
nand U52 (N_52,In_117,In_218);
nor U53 (N_53,In_188,In_116);
nand U54 (N_54,In_329,In_20);
nand U55 (N_55,In_303,In_70);
and U56 (N_56,In_78,In_335);
nor U57 (N_57,In_487,In_322);
and U58 (N_58,In_481,In_149);
nor U59 (N_59,In_69,In_361);
nand U60 (N_60,In_100,In_139);
nor U61 (N_61,In_420,In_405);
nand U62 (N_62,In_128,In_51);
nor U63 (N_63,In_308,In_73);
nor U64 (N_64,In_131,In_388);
nand U65 (N_65,In_285,In_22);
or U66 (N_66,In_470,In_181);
and U67 (N_67,In_397,In_342);
xor U68 (N_68,In_450,In_50);
nand U69 (N_69,In_243,In_224);
or U70 (N_70,In_287,In_62);
and U71 (N_71,In_166,In_263);
and U72 (N_72,In_246,In_257);
and U73 (N_73,In_151,In_354);
nand U74 (N_74,In_140,In_353);
and U75 (N_75,In_57,In_283);
and U76 (N_76,In_43,In_486);
nor U77 (N_77,In_253,In_196);
or U78 (N_78,In_201,In_367);
nor U79 (N_79,In_250,In_307);
nand U80 (N_80,In_169,In_356);
nand U81 (N_81,In_58,N_23);
nor U82 (N_82,N_53,In_118);
nor U83 (N_83,In_26,In_302);
xor U84 (N_84,In_61,In_114);
and U85 (N_85,In_314,In_28);
or U86 (N_86,In_371,In_492);
nor U87 (N_87,N_11,In_122);
nor U88 (N_88,In_413,In_23);
or U89 (N_89,In_230,In_475);
nor U90 (N_90,In_138,N_73);
nor U91 (N_91,In_309,In_418);
and U92 (N_92,In_394,In_130);
nand U93 (N_93,In_158,In_53);
nand U94 (N_94,In_238,In_458);
nand U95 (N_95,N_8,In_316);
xor U96 (N_96,In_349,N_58);
nor U97 (N_97,In_171,In_310);
nand U98 (N_98,In_203,N_35);
or U99 (N_99,In_251,In_152);
nand U100 (N_100,In_264,In_170);
and U101 (N_101,In_272,In_242);
and U102 (N_102,In_190,In_312);
or U103 (N_103,N_19,In_345);
nor U104 (N_104,N_14,In_240);
and U105 (N_105,In_111,In_176);
and U106 (N_106,In_466,In_150);
nor U107 (N_107,In_258,N_71);
xnor U108 (N_108,In_378,In_261);
or U109 (N_109,N_4,In_135);
nand U110 (N_110,In_412,In_103);
or U111 (N_111,In_374,In_236);
nand U112 (N_112,In_9,In_390);
nor U113 (N_113,In_319,In_408);
xor U114 (N_114,In_351,In_18);
nor U115 (N_115,In_120,In_325);
or U116 (N_116,N_18,In_197);
nand U117 (N_117,N_9,In_200);
nand U118 (N_118,In_67,N_52);
nand U119 (N_119,In_154,In_449);
or U120 (N_120,In_231,N_43);
or U121 (N_121,In_372,In_455);
nand U122 (N_122,N_32,In_447);
nand U123 (N_123,N_56,In_35);
nor U124 (N_124,In_381,N_7);
or U125 (N_125,In_365,In_71);
nor U126 (N_126,In_14,In_99);
nor U127 (N_127,In_168,In_155);
nor U128 (N_128,In_284,In_223);
and U129 (N_129,In_153,In_32);
nand U130 (N_130,In_64,In_89);
or U131 (N_131,In_401,In_334);
nand U132 (N_132,In_431,In_299);
nor U133 (N_133,In_289,N_24);
nand U134 (N_134,In_472,N_27);
and U135 (N_135,In_206,In_17);
and U136 (N_136,N_54,In_38);
and U137 (N_137,In_5,In_453);
nand U138 (N_138,In_396,In_235);
nand U139 (N_139,In_55,N_46);
or U140 (N_140,In_85,In_344);
nor U141 (N_141,In_368,In_254);
and U142 (N_142,In_317,In_474);
nor U143 (N_143,In_160,In_423);
or U144 (N_144,In_493,In_129);
or U145 (N_145,In_141,In_430);
nand U146 (N_146,In_8,In_48);
and U147 (N_147,In_421,In_465);
or U148 (N_148,In_333,In_277);
or U149 (N_149,In_477,In_393);
nand U150 (N_150,N_64,In_68);
and U151 (N_151,N_20,N_78);
or U152 (N_152,N_15,N_127);
nor U153 (N_153,In_375,In_6);
nor U154 (N_154,N_126,In_112);
or U155 (N_155,N_104,In_52);
and U156 (N_156,N_77,In_320);
and U157 (N_157,N_75,N_84);
nand U158 (N_158,N_69,In_249);
nor U159 (N_159,In_210,In_145);
and U160 (N_160,N_100,In_471);
and U161 (N_161,In_498,In_494);
nor U162 (N_162,N_128,In_460);
and U163 (N_163,N_115,In_366);
or U164 (N_164,In_376,In_96);
nand U165 (N_165,In_119,N_29);
xor U166 (N_166,In_382,N_137);
nor U167 (N_167,In_499,In_215);
nand U168 (N_168,In_425,N_31);
nand U169 (N_169,In_446,N_25);
nor U170 (N_170,In_90,In_391);
and U171 (N_171,N_61,In_340);
or U172 (N_172,In_358,N_85);
or U173 (N_173,In_268,N_90);
xor U174 (N_174,In_42,N_65);
nand U175 (N_175,In_74,N_107);
and U176 (N_176,N_44,In_414);
and U177 (N_177,In_434,In_225);
or U178 (N_178,In_290,N_33);
nand U179 (N_179,In_179,In_157);
and U180 (N_180,In_276,In_193);
and U181 (N_181,In_262,N_114);
nand U182 (N_182,In_199,N_95);
nor U183 (N_183,In_180,In_379);
nand U184 (N_184,In_398,N_89);
or U185 (N_185,N_118,In_399);
nor U186 (N_186,N_42,In_7);
and U187 (N_187,N_130,In_226);
or U188 (N_188,N_5,N_116);
and U189 (N_189,In_60,N_79);
and U190 (N_190,In_237,In_12);
nor U191 (N_191,N_146,In_313);
or U192 (N_192,N_139,In_457);
or U193 (N_193,In_437,N_68);
and U194 (N_194,In_270,N_120);
nor U195 (N_195,In_288,In_338);
nand U196 (N_196,In_232,In_488);
or U197 (N_197,In_15,In_443);
nor U198 (N_198,In_91,In_194);
nor U199 (N_199,N_124,In_241);
and U200 (N_200,N_74,N_94);
and U201 (N_201,N_105,N_10);
and U202 (N_202,In_95,N_28);
and U203 (N_203,N_37,N_45);
or U204 (N_204,In_220,N_135);
and U205 (N_205,N_55,In_101);
or U206 (N_206,N_113,In_123);
nand U207 (N_207,N_1,N_91);
nand U208 (N_208,N_12,In_165);
or U209 (N_209,In_185,In_92);
and U210 (N_210,In_37,In_410);
and U211 (N_211,In_305,N_63);
and U212 (N_212,In_403,In_369);
nor U213 (N_213,In_41,N_119);
nor U214 (N_214,In_16,N_38);
or U215 (N_215,In_234,In_229);
or U216 (N_216,N_49,N_96);
or U217 (N_217,In_167,In_177);
nor U218 (N_218,In_46,N_39);
nor U219 (N_219,In_267,In_473);
or U220 (N_220,In_451,In_39);
and U221 (N_221,In_456,In_435);
or U222 (N_222,N_66,In_341);
nand U223 (N_223,N_3,In_81);
nor U224 (N_224,In_279,In_392);
or U225 (N_225,N_216,In_294);
or U226 (N_226,In_298,N_0);
nand U227 (N_227,In_86,N_181);
nor U228 (N_228,N_161,In_45);
or U229 (N_229,N_17,In_49);
or U230 (N_230,In_192,N_83);
nor U231 (N_231,N_111,In_94);
nand U232 (N_232,N_189,N_175);
or U233 (N_233,N_98,In_296);
or U234 (N_234,In_260,In_159);
and U235 (N_235,In_172,N_172);
nor U236 (N_236,In_359,N_82);
and U237 (N_237,In_452,N_123);
nand U238 (N_238,In_291,N_99);
nand U239 (N_239,N_214,In_33);
and U240 (N_240,N_36,In_370);
nand U241 (N_241,In_3,N_129);
or U242 (N_242,N_51,In_10);
nor U243 (N_243,N_148,N_193);
nor U244 (N_244,N_155,N_81);
nand U245 (N_245,N_70,In_213);
and U246 (N_246,N_162,In_271);
xnor U247 (N_247,In_227,N_183);
or U248 (N_248,In_387,N_182);
and U249 (N_249,N_219,In_221);
and U250 (N_250,N_131,N_190);
nand U251 (N_251,In_384,In_496);
and U252 (N_252,N_62,In_324);
nor U253 (N_253,N_122,N_207);
or U254 (N_254,In_417,In_107);
nor U255 (N_255,In_377,In_79);
xnor U256 (N_256,N_169,N_170);
nand U257 (N_257,N_47,N_198);
and U258 (N_258,In_77,In_115);
nand U259 (N_259,N_48,In_143);
and U260 (N_260,In_0,In_346);
nor U261 (N_261,N_106,In_315);
and U262 (N_262,In_205,N_168);
nand U263 (N_263,N_194,In_146);
or U264 (N_264,In_164,In_497);
and U265 (N_265,N_125,In_144);
or U266 (N_266,N_2,In_105);
nor U267 (N_267,N_203,N_176);
and U268 (N_268,In_323,N_140);
nor U269 (N_269,In_97,In_484);
nor U270 (N_270,N_212,N_167);
nor U271 (N_271,N_13,In_207);
nor U272 (N_272,N_185,N_209);
and U273 (N_273,N_171,N_30);
nand U274 (N_274,In_191,In_347);
nor U275 (N_275,N_204,N_188);
nor U276 (N_276,In_88,In_198);
nor U277 (N_277,In_350,N_142);
nor U278 (N_278,In_482,N_213);
nand U279 (N_279,N_166,N_97);
or U280 (N_280,In_293,In_36);
nand U281 (N_281,N_40,In_336);
nor U282 (N_282,N_60,N_138);
nor U283 (N_283,In_27,In_432);
and U284 (N_284,N_196,In_239);
nand U285 (N_285,In_416,N_136);
or U286 (N_286,N_159,In_362);
and U287 (N_287,N_153,N_218);
and U288 (N_288,N_57,N_149);
nor U289 (N_289,In_436,N_88);
or U290 (N_290,In_489,N_217);
nand U291 (N_291,In_360,In_464);
or U292 (N_292,In_304,N_200);
and U293 (N_293,N_26,N_22);
nor U294 (N_294,In_63,In_195);
nor U295 (N_295,In_208,In_233);
or U296 (N_296,N_59,In_54);
and U297 (N_297,N_6,N_154);
nor U298 (N_298,N_186,In_44);
and U299 (N_299,N_141,N_178);
nand U300 (N_300,N_267,N_277);
and U301 (N_301,In_11,N_227);
and U302 (N_302,N_229,N_86);
nor U303 (N_303,N_163,N_156);
nor U304 (N_304,N_164,N_187);
nand U305 (N_305,N_278,N_67);
nand U306 (N_306,In_29,N_197);
nor U307 (N_307,In_280,In_222);
and U308 (N_308,N_246,N_110);
or U309 (N_309,N_103,N_180);
nand U310 (N_310,In_106,In_245);
nand U311 (N_311,N_282,N_232);
nor U312 (N_312,In_133,N_16);
nand U313 (N_313,N_291,N_221);
or U314 (N_314,In_174,In_352);
nand U315 (N_315,N_226,N_223);
and U316 (N_316,N_280,In_444);
nand U317 (N_317,N_262,N_260);
nand U318 (N_318,N_151,In_385);
nand U319 (N_319,N_179,In_424);
nand U320 (N_320,N_144,In_108);
nand U321 (N_321,N_150,In_479);
and U322 (N_322,N_108,N_132);
nand U323 (N_323,N_143,N_244);
xor U324 (N_324,N_275,N_249);
and U325 (N_325,N_255,In_318);
or U326 (N_326,N_276,N_257);
and U327 (N_327,In_278,N_174);
or U328 (N_328,N_250,In_134);
nor U329 (N_329,N_253,N_133);
and U330 (N_330,N_112,N_286);
nand U331 (N_331,N_76,In_21);
or U332 (N_332,N_147,In_1);
nand U333 (N_333,N_252,N_184);
or U334 (N_334,In_326,N_205);
nand U335 (N_335,In_13,N_265);
nand U336 (N_336,N_72,N_293);
nor U337 (N_337,N_289,In_147);
nand U338 (N_338,In_438,In_178);
nor U339 (N_339,N_243,N_238);
nand U340 (N_340,N_80,In_485);
and U341 (N_341,N_297,N_199);
nand U342 (N_342,In_187,In_182);
and U343 (N_343,N_220,In_84);
nor U344 (N_344,N_145,In_204);
nand U345 (N_345,In_98,N_87);
nand U346 (N_346,N_208,In_454);
and U347 (N_347,N_225,N_274);
or U348 (N_348,N_230,In_490);
and U349 (N_349,N_264,In_30);
nor U350 (N_350,N_228,N_152);
and U351 (N_351,N_222,N_160);
and U352 (N_352,N_235,N_191);
nand U353 (N_353,N_215,N_206);
xnor U354 (N_354,N_283,N_263);
or U355 (N_355,N_231,In_440);
nand U356 (N_356,N_245,N_102);
and U357 (N_357,N_173,In_247);
nor U358 (N_358,In_491,In_4);
and U359 (N_359,In_273,N_210);
or U360 (N_360,N_202,N_259);
nand U361 (N_361,N_269,N_34);
and U362 (N_362,In_478,N_242);
nand U363 (N_363,N_287,N_258);
and U364 (N_364,In_25,N_288);
nor U365 (N_365,In_439,N_158);
nand U366 (N_366,N_157,N_281);
nor U367 (N_367,N_284,In_212);
nor U368 (N_368,N_273,N_247);
and U369 (N_369,N_121,N_248);
nand U370 (N_370,N_296,N_256);
nand U371 (N_371,In_34,N_298);
nor U372 (N_372,In_126,In_407);
nor U373 (N_373,In_109,In_409);
nand U374 (N_374,N_279,N_254);
and U375 (N_375,N_341,N_306);
nand U376 (N_376,In_292,N_236);
nor U377 (N_377,In_183,N_233);
and U378 (N_378,N_312,N_330);
nor U379 (N_379,N_303,N_332);
nor U380 (N_380,N_309,N_354);
or U381 (N_381,N_299,In_80);
and U382 (N_382,N_333,N_360);
nor U383 (N_383,N_367,N_294);
and U384 (N_384,N_319,N_109);
or U385 (N_385,N_192,N_325);
and U386 (N_386,N_348,In_380);
nand U387 (N_387,N_285,N_272);
and U388 (N_388,N_343,N_373);
or U389 (N_389,N_318,N_352);
or U390 (N_390,N_351,N_311);
and U391 (N_391,N_320,In_463);
or U392 (N_392,N_41,N_101);
nor U393 (N_393,N_336,N_369);
nand U394 (N_394,N_334,In_219);
or U395 (N_395,N_240,N_326);
nor U396 (N_396,N_324,N_372);
nor U397 (N_397,N_304,N_177);
or U398 (N_398,N_358,N_355);
or U399 (N_399,N_329,N_314);
nand U400 (N_400,N_308,In_411);
nor U401 (N_401,N_370,N_335);
and U402 (N_402,In_297,N_328);
nor U403 (N_403,N_315,N_371);
nand U404 (N_404,N_346,N_251);
and U405 (N_405,N_338,N_366);
nor U406 (N_406,In_137,N_201);
and U407 (N_407,N_165,N_339);
and U408 (N_408,N_357,N_321);
nand U409 (N_409,N_239,N_195);
or U410 (N_410,N_317,N_347);
nor U411 (N_411,In_265,In_75);
nor U412 (N_412,N_307,N_323);
or U413 (N_413,N_305,N_362);
nor U414 (N_414,N_327,N_313);
nor U415 (N_415,N_337,N_134);
and U416 (N_416,N_295,N_93);
nand U417 (N_417,N_374,N_302);
or U418 (N_418,N_92,N_271);
nand U419 (N_419,N_331,N_211);
nand U420 (N_420,N_21,N_301);
and U421 (N_421,In_286,N_344);
nand U422 (N_422,N_364,N_356);
nand U423 (N_423,N_310,N_322);
or U424 (N_424,N_316,N_241);
nand U425 (N_425,N_345,N_268);
and U426 (N_426,N_224,N_350);
nand U427 (N_427,N_50,N_368);
nand U428 (N_428,N_342,N_290);
and U429 (N_429,N_349,N_365);
and U430 (N_430,N_266,N_361);
nand U431 (N_431,In_76,N_234);
and U432 (N_432,N_261,N_359);
and U433 (N_433,N_300,N_363);
and U434 (N_434,N_270,N_340);
and U435 (N_435,In_441,N_237);
nand U436 (N_436,N_353,N_117);
nor U437 (N_437,N_292,N_340);
nand U438 (N_438,In_80,N_352);
nand U439 (N_439,N_192,N_301);
and U440 (N_440,N_237,N_312);
or U441 (N_441,N_334,N_300);
nor U442 (N_442,N_362,N_290);
nand U443 (N_443,In_292,N_331);
or U444 (N_444,N_355,N_332);
xnor U445 (N_445,N_331,N_359);
and U446 (N_446,In_80,N_365);
nand U447 (N_447,N_336,N_299);
nand U448 (N_448,In_219,N_339);
nand U449 (N_449,N_358,N_353);
nand U450 (N_450,N_386,N_384);
nor U451 (N_451,N_391,N_408);
nand U452 (N_452,N_429,N_412);
nor U453 (N_453,N_427,N_398);
nand U454 (N_454,N_376,N_422);
and U455 (N_455,N_387,N_414);
nand U456 (N_456,N_444,N_438);
nor U457 (N_457,N_388,N_390);
nor U458 (N_458,N_436,N_418);
nand U459 (N_459,N_403,N_400);
nand U460 (N_460,N_421,N_405);
nand U461 (N_461,N_396,N_382);
nand U462 (N_462,N_389,N_420);
and U463 (N_463,N_392,N_432);
nand U464 (N_464,N_445,N_423);
or U465 (N_465,N_449,N_406);
and U466 (N_466,N_385,N_433);
nor U467 (N_467,N_393,N_447);
xor U468 (N_468,N_407,N_424);
or U469 (N_469,N_439,N_380);
nand U470 (N_470,N_411,N_375);
nor U471 (N_471,N_430,N_397);
and U472 (N_472,N_383,N_413);
nand U473 (N_473,N_416,N_448);
nand U474 (N_474,N_443,N_415);
and U475 (N_475,N_426,N_419);
nor U476 (N_476,N_379,N_410);
or U477 (N_477,N_378,N_431);
nand U478 (N_478,N_425,N_394);
and U479 (N_479,N_440,N_434);
nor U480 (N_480,N_402,N_428);
or U481 (N_481,N_381,N_442);
or U482 (N_482,N_399,N_437);
xor U483 (N_483,N_417,N_409);
nor U484 (N_484,N_377,N_401);
nand U485 (N_485,N_395,N_446);
or U486 (N_486,N_435,N_404);
and U487 (N_487,N_441,N_443);
nor U488 (N_488,N_394,N_414);
nand U489 (N_489,N_409,N_399);
or U490 (N_490,N_442,N_426);
or U491 (N_491,N_439,N_411);
nor U492 (N_492,N_402,N_404);
nor U493 (N_493,N_414,N_401);
and U494 (N_494,N_421,N_404);
or U495 (N_495,N_429,N_435);
nand U496 (N_496,N_447,N_388);
and U497 (N_497,N_431,N_440);
nor U498 (N_498,N_426,N_423);
nor U499 (N_499,N_424,N_412);
or U500 (N_500,N_380,N_418);
and U501 (N_501,N_435,N_427);
or U502 (N_502,N_379,N_436);
and U503 (N_503,N_376,N_387);
or U504 (N_504,N_440,N_438);
nand U505 (N_505,N_409,N_428);
and U506 (N_506,N_396,N_432);
or U507 (N_507,N_440,N_379);
or U508 (N_508,N_429,N_421);
nand U509 (N_509,N_441,N_444);
nor U510 (N_510,N_380,N_441);
and U511 (N_511,N_437,N_433);
nor U512 (N_512,N_417,N_436);
and U513 (N_513,N_427,N_422);
nand U514 (N_514,N_412,N_397);
or U515 (N_515,N_402,N_382);
nor U516 (N_516,N_387,N_422);
and U517 (N_517,N_391,N_392);
nand U518 (N_518,N_416,N_420);
nor U519 (N_519,N_392,N_412);
or U520 (N_520,N_403,N_410);
nor U521 (N_521,N_435,N_396);
nand U522 (N_522,N_412,N_446);
or U523 (N_523,N_389,N_429);
nor U524 (N_524,N_439,N_447);
or U525 (N_525,N_487,N_519);
nor U526 (N_526,N_507,N_450);
and U527 (N_527,N_473,N_491);
or U528 (N_528,N_521,N_454);
nor U529 (N_529,N_512,N_509);
and U530 (N_530,N_467,N_468);
or U531 (N_531,N_499,N_469);
and U532 (N_532,N_497,N_516);
nor U533 (N_533,N_482,N_472);
or U534 (N_534,N_474,N_490);
nand U535 (N_535,N_523,N_502);
or U536 (N_536,N_496,N_455);
nor U537 (N_537,N_505,N_503);
nand U538 (N_538,N_460,N_470);
and U539 (N_539,N_518,N_451);
nand U540 (N_540,N_504,N_495);
nor U541 (N_541,N_511,N_464);
or U542 (N_542,N_488,N_522);
nor U543 (N_543,N_486,N_506);
or U544 (N_544,N_517,N_475);
and U545 (N_545,N_510,N_508);
and U546 (N_546,N_461,N_462);
nor U547 (N_547,N_471,N_478);
nand U548 (N_548,N_484,N_483);
and U549 (N_549,N_520,N_524);
or U550 (N_550,N_476,N_494);
or U551 (N_551,N_480,N_477);
nor U552 (N_552,N_456,N_513);
or U553 (N_553,N_479,N_452);
and U554 (N_554,N_466,N_498);
and U555 (N_555,N_485,N_465);
nor U556 (N_556,N_489,N_500);
nand U557 (N_557,N_457,N_458);
and U558 (N_558,N_514,N_501);
nand U559 (N_559,N_492,N_493);
and U560 (N_560,N_481,N_453);
or U561 (N_561,N_459,N_463);
or U562 (N_562,N_515,N_488);
or U563 (N_563,N_459,N_488);
nor U564 (N_564,N_488,N_473);
nand U565 (N_565,N_478,N_469);
or U566 (N_566,N_518,N_513);
and U567 (N_567,N_520,N_487);
and U568 (N_568,N_450,N_480);
nor U569 (N_569,N_489,N_506);
nor U570 (N_570,N_468,N_494);
and U571 (N_571,N_458,N_473);
nand U572 (N_572,N_507,N_477);
nand U573 (N_573,N_516,N_475);
nand U574 (N_574,N_464,N_468);
or U575 (N_575,N_484,N_490);
xnor U576 (N_576,N_459,N_465);
and U577 (N_577,N_478,N_458);
or U578 (N_578,N_499,N_501);
nand U579 (N_579,N_497,N_509);
nor U580 (N_580,N_509,N_459);
nand U581 (N_581,N_480,N_504);
or U582 (N_582,N_510,N_506);
and U583 (N_583,N_506,N_453);
or U584 (N_584,N_468,N_488);
or U585 (N_585,N_464,N_506);
and U586 (N_586,N_469,N_483);
nor U587 (N_587,N_521,N_497);
nand U588 (N_588,N_495,N_452);
nor U589 (N_589,N_455,N_464);
nor U590 (N_590,N_504,N_494);
nand U591 (N_591,N_484,N_505);
nand U592 (N_592,N_457,N_490);
nor U593 (N_593,N_453,N_498);
nand U594 (N_594,N_507,N_464);
and U595 (N_595,N_513,N_470);
nor U596 (N_596,N_518,N_475);
nor U597 (N_597,N_470,N_483);
nand U598 (N_598,N_510,N_516);
or U599 (N_599,N_487,N_468);
and U600 (N_600,N_541,N_526);
nand U601 (N_601,N_560,N_575);
nand U602 (N_602,N_528,N_590);
nor U603 (N_603,N_543,N_545);
and U604 (N_604,N_554,N_591);
nand U605 (N_605,N_572,N_585);
or U606 (N_606,N_540,N_565);
nand U607 (N_607,N_547,N_525);
nor U608 (N_608,N_531,N_563);
nor U609 (N_609,N_548,N_594);
nand U610 (N_610,N_534,N_544);
nor U611 (N_611,N_588,N_532);
nand U612 (N_612,N_576,N_550);
nand U613 (N_613,N_582,N_529);
and U614 (N_614,N_537,N_578);
nand U615 (N_615,N_559,N_552);
nor U616 (N_616,N_542,N_562);
and U617 (N_617,N_595,N_577);
nand U618 (N_618,N_527,N_583);
nand U619 (N_619,N_574,N_555);
and U620 (N_620,N_596,N_573);
or U621 (N_621,N_569,N_566);
and U622 (N_622,N_570,N_551);
nand U623 (N_623,N_597,N_553);
and U624 (N_624,N_533,N_584);
or U625 (N_625,N_558,N_581);
or U626 (N_626,N_589,N_561);
and U627 (N_627,N_536,N_586);
nand U628 (N_628,N_530,N_535);
nand U629 (N_629,N_593,N_538);
or U630 (N_630,N_568,N_557);
and U631 (N_631,N_571,N_579);
or U632 (N_632,N_564,N_598);
and U633 (N_633,N_539,N_556);
or U634 (N_634,N_592,N_549);
nand U635 (N_635,N_580,N_587);
nor U636 (N_636,N_567,N_546);
nand U637 (N_637,N_599,N_546);
and U638 (N_638,N_593,N_569);
or U639 (N_639,N_579,N_572);
and U640 (N_640,N_543,N_590);
nand U641 (N_641,N_553,N_591);
or U642 (N_642,N_599,N_525);
or U643 (N_643,N_596,N_548);
nor U644 (N_644,N_533,N_545);
nor U645 (N_645,N_598,N_525);
nand U646 (N_646,N_551,N_599);
and U647 (N_647,N_566,N_560);
or U648 (N_648,N_554,N_548);
or U649 (N_649,N_567,N_562);
nand U650 (N_650,N_529,N_568);
and U651 (N_651,N_550,N_567);
nand U652 (N_652,N_557,N_528);
xnor U653 (N_653,N_579,N_570);
nand U654 (N_654,N_542,N_593);
or U655 (N_655,N_571,N_545);
and U656 (N_656,N_596,N_583);
and U657 (N_657,N_537,N_548);
nand U658 (N_658,N_532,N_596);
nand U659 (N_659,N_532,N_595);
or U660 (N_660,N_536,N_587);
nor U661 (N_661,N_565,N_532);
nor U662 (N_662,N_534,N_550);
nor U663 (N_663,N_560,N_572);
nor U664 (N_664,N_538,N_579);
nor U665 (N_665,N_581,N_564);
or U666 (N_666,N_570,N_593);
nor U667 (N_667,N_589,N_577);
and U668 (N_668,N_577,N_583);
and U669 (N_669,N_559,N_566);
or U670 (N_670,N_580,N_567);
and U671 (N_671,N_592,N_573);
and U672 (N_672,N_561,N_539);
and U673 (N_673,N_564,N_575);
nand U674 (N_674,N_538,N_544);
or U675 (N_675,N_667,N_625);
and U676 (N_676,N_624,N_661);
or U677 (N_677,N_656,N_647);
and U678 (N_678,N_631,N_638);
nand U679 (N_679,N_640,N_628);
and U680 (N_680,N_602,N_655);
or U681 (N_681,N_621,N_660);
or U682 (N_682,N_635,N_618);
and U683 (N_683,N_620,N_673);
nor U684 (N_684,N_611,N_629);
or U685 (N_685,N_612,N_616);
or U686 (N_686,N_619,N_666);
nor U687 (N_687,N_615,N_604);
and U688 (N_688,N_609,N_634);
nand U689 (N_689,N_658,N_650);
and U690 (N_690,N_643,N_636);
nor U691 (N_691,N_659,N_603);
or U692 (N_692,N_665,N_670);
and U693 (N_693,N_668,N_606);
and U694 (N_694,N_605,N_601);
or U695 (N_695,N_648,N_600);
nand U696 (N_696,N_663,N_657);
nor U697 (N_697,N_608,N_639);
or U698 (N_698,N_632,N_613);
nand U699 (N_699,N_637,N_644);
or U700 (N_700,N_630,N_674);
nor U701 (N_701,N_614,N_626);
nand U702 (N_702,N_646,N_669);
and U703 (N_703,N_651,N_627);
and U704 (N_704,N_610,N_664);
or U705 (N_705,N_633,N_623);
nor U706 (N_706,N_653,N_645);
or U707 (N_707,N_652,N_642);
nand U708 (N_708,N_607,N_617);
nor U709 (N_709,N_672,N_671);
or U710 (N_710,N_622,N_641);
nor U711 (N_711,N_649,N_654);
nand U712 (N_712,N_662,N_644);
nand U713 (N_713,N_664,N_648);
nand U714 (N_714,N_607,N_606);
or U715 (N_715,N_605,N_602);
and U716 (N_716,N_656,N_622);
nand U717 (N_717,N_610,N_631);
and U718 (N_718,N_661,N_628);
nor U719 (N_719,N_616,N_613);
and U720 (N_720,N_613,N_610);
or U721 (N_721,N_651,N_613);
or U722 (N_722,N_667,N_662);
and U723 (N_723,N_658,N_635);
nand U724 (N_724,N_643,N_671);
nor U725 (N_725,N_624,N_614);
nor U726 (N_726,N_673,N_646);
nand U727 (N_727,N_636,N_611);
nor U728 (N_728,N_624,N_654);
or U729 (N_729,N_609,N_611);
or U730 (N_730,N_651,N_644);
nor U731 (N_731,N_670,N_619);
nor U732 (N_732,N_602,N_603);
nand U733 (N_733,N_615,N_651);
and U734 (N_734,N_631,N_624);
and U735 (N_735,N_601,N_604);
xnor U736 (N_736,N_601,N_612);
nand U737 (N_737,N_601,N_665);
or U738 (N_738,N_656,N_605);
or U739 (N_739,N_658,N_667);
nand U740 (N_740,N_664,N_614);
nor U741 (N_741,N_645,N_615);
or U742 (N_742,N_608,N_614);
nand U743 (N_743,N_665,N_648);
or U744 (N_744,N_630,N_672);
or U745 (N_745,N_636,N_632);
nand U746 (N_746,N_614,N_647);
and U747 (N_747,N_636,N_652);
nor U748 (N_748,N_638,N_616);
nand U749 (N_749,N_636,N_612);
nand U750 (N_750,N_745,N_682);
nand U751 (N_751,N_680,N_715);
nor U752 (N_752,N_726,N_736);
nand U753 (N_753,N_710,N_676);
or U754 (N_754,N_749,N_734);
nand U755 (N_755,N_737,N_675);
nand U756 (N_756,N_716,N_742);
nand U757 (N_757,N_727,N_683);
or U758 (N_758,N_679,N_691);
and U759 (N_759,N_740,N_695);
or U760 (N_760,N_693,N_678);
or U761 (N_761,N_719,N_718);
or U762 (N_762,N_744,N_722);
nand U763 (N_763,N_735,N_690);
or U764 (N_764,N_701,N_699);
and U765 (N_765,N_739,N_709);
and U766 (N_766,N_686,N_697);
nand U767 (N_767,N_730,N_684);
or U768 (N_768,N_723,N_746);
nand U769 (N_769,N_748,N_741);
or U770 (N_770,N_729,N_692);
and U771 (N_771,N_694,N_717);
or U772 (N_772,N_720,N_721);
or U773 (N_773,N_685,N_731);
and U774 (N_774,N_702,N_711);
and U775 (N_775,N_698,N_708);
or U776 (N_776,N_714,N_724);
or U777 (N_777,N_738,N_696);
and U778 (N_778,N_733,N_705);
nand U779 (N_779,N_712,N_700);
nor U780 (N_780,N_747,N_707);
and U781 (N_781,N_687,N_681);
or U782 (N_782,N_677,N_728);
nand U783 (N_783,N_703,N_704);
nor U784 (N_784,N_732,N_725);
or U785 (N_785,N_688,N_689);
nand U786 (N_786,N_713,N_743);
nor U787 (N_787,N_706,N_720);
or U788 (N_788,N_682,N_721);
nand U789 (N_789,N_713,N_683);
or U790 (N_790,N_725,N_736);
nand U791 (N_791,N_749,N_717);
nor U792 (N_792,N_678,N_724);
and U793 (N_793,N_693,N_705);
nand U794 (N_794,N_733,N_748);
and U795 (N_795,N_698,N_721);
and U796 (N_796,N_677,N_685);
nor U797 (N_797,N_696,N_704);
nand U798 (N_798,N_742,N_740);
nor U799 (N_799,N_736,N_688);
or U800 (N_800,N_701,N_723);
and U801 (N_801,N_739,N_749);
nor U802 (N_802,N_680,N_709);
nand U803 (N_803,N_738,N_678);
and U804 (N_804,N_737,N_713);
or U805 (N_805,N_738,N_732);
nand U806 (N_806,N_744,N_686);
and U807 (N_807,N_734,N_743);
and U808 (N_808,N_727,N_688);
nand U809 (N_809,N_697,N_739);
nand U810 (N_810,N_730,N_733);
and U811 (N_811,N_730,N_739);
and U812 (N_812,N_736,N_692);
nand U813 (N_813,N_740,N_728);
or U814 (N_814,N_707,N_699);
or U815 (N_815,N_732,N_683);
or U816 (N_816,N_681,N_678);
nand U817 (N_817,N_741,N_717);
or U818 (N_818,N_708,N_706);
and U819 (N_819,N_715,N_703);
or U820 (N_820,N_723,N_717);
nand U821 (N_821,N_727,N_713);
or U822 (N_822,N_690,N_711);
and U823 (N_823,N_720,N_713);
or U824 (N_824,N_679,N_694);
nand U825 (N_825,N_802,N_767);
or U826 (N_826,N_766,N_815);
nor U827 (N_827,N_768,N_757);
or U828 (N_828,N_770,N_794);
nand U829 (N_829,N_761,N_782);
or U830 (N_830,N_824,N_792);
nand U831 (N_831,N_818,N_760);
or U832 (N_832,N_758,N_788);
nand U833 (N_833,N_810,N_807);
nor U834 (N_834,N_786,N_808);
xor U835 (N_835,N_772,N_819);
nor U836 (N_836,N_804,N_812);
and U837 (N_837,N_769,N_823);
or U838 (N_838,N_800,N_811);
and U839 (N_839,N_777,N_776);
and U840 (N_840,N_778,N_803);
and U841 (N_841,N_799,N_783);
nor U842 (N_842,N_806,N_784);
and U843 (N_843,N_781,N_759);
nand U844 (N_844,N_797,N_785);
xnor U845 (N_845,N_773,N_791);
and U846 (N_846,N_820,N_752);
nand U847 (N_847,N_821,N_753);
nor U848 (N_848,N_751,N_796);
and U849 (N_849,N_795,N_764);
nor U850 (N_850,N_754,N_790);
and U851 (N_851,N_755,N_775);
and U852 (N_852,N_816,N_765);
and U853 (N_853,N_774,N_779);
nor U854 (N_854,N_817,N_813);
nand U855 (N_855,N_814,N_756);
or U856 (N_856,N_805,N_763);
or U857 (N_857,N_789,N_798);
nor U858 (N_858,N_787,N_771);
and U859 (N_859,N_809,N_780);
nor U860 (N_860,N_750,N_793);
and U861 (N_861,N_762,N_822);
nand U862 (N_862,N_801,N_770);
and U863 (N_863,N_811,N_753);
and U864 (N_864,N_750,N_778);
nand U865 (N_865,N_772,N_784);
and U866 (N_866,N_801,N_750);
nor U867 (N_867,N_781,N_773);
nor U868 (N_868,N_755,N_754);
or U869 (N_869,N_766,N_810);
or U870 (N_870,N_755,N_788);
nand U871 (N_871,N_763,N_792);
or U872 (N_872,N_774,N_822);
or U873 (N_873,N_814,N_775);
or U874 (N_874,N_782,N_796);
and U875 (N_875,N_791,N_795);
nand U876 (N_876,N_786,N_810);
and U877 (N_877,N_778,N_807);
nand U878 (N_878,N_753,N_824);
xor U879 (N_879,N_773,N_775);
nand U880 (N_880,N_804,N_818);
and U881 (N_881,N_824,N_769);
and U882 (N_882,N_768,N_788);
and U883 (N_883,N_792,N_802);
or U884 (N_884,N_788,N_769);
and U885 (N_885,N_770,N_780);
and U886 (N_886,N_763,N_781);
nand U887 (N_887,N_810,N_816);
or U888 (N_888,N_763,N_766);
xnor U889 (N_889,N_787,N_820);
nand U890 (N_890,N_806,N_819);
nand U891 (N_891,N_817,N_766);
and U892 (N_892,N_781,N_772);
nor U893 (N_893,N_800,N_768);
nand U894 (N_894,N_773,N_780);
or U895 (N_895,N_785,N_757);
and U896 (N_896,N_810,N_814);
or U897 (N_897,N_803,N_769);
nand U898 (N_898,N_823,N_787);
nand U899 (N_899,N_819,N_774);
nand U900 (N_900,N_841,N_825);
and U901 (N_901,N_829,N_899);
and U902 (N_902,N_894,N_848);
nand U903 (N_903,N_844,N_884);
and U904 (N_904,N_885,N_846);
and U905 (N_905,N_874,N_881);
or U906 (N_906,N_831,N_862);
or U907 (N_907,N_871,N_861);
nor U908 (N_908,N_858,N_843);
nand U909 (N_909,N_868,N_875);
and U910 (N_910,N_859,N_886);
and U911 (N_911,N_828,N_890);
nor U912 (N_912,N_855,N_865);
nor U913 (N_913,N_834,N_840);
nand U914 (N_914,N_863,N_833);
nor U915 (N_915,N_878,N_851);
and U916 (N_916,N_896,N_852);
or U917 (N_917,N_836,N_888);
nor U918 (N_918,N_839,N_853);
nor U919 (N_919,N_830,N_850);
or U920 (N_920,N_869,N_892);
or U921 (N_921,N_891,N_872);
nand U922 (N_922,N_849,N_887);
or U923 (N_923,N_895,N_898);
nor U924 (N_924,N_837,N_857);
or U925 (N_925,N_842,N_832);
nor U926 (N_926,N_883,N_864);
and U927 (N_927,N_867,N_889);
and U928 (N_928,N_826,N_893);
nor U929 (N_929,N_870,N_847);
or U930 (N_930,N_845,N_827);
and U931 (N_931,N_880,N_876);
nor U932 (N_932,N_877,N_873);
nand U933 (N_933,N_897,N_854);
and U934 (N_934,N_879,N_856);
or U935 (N_935,N_860,N_882);
or U936 (N_936,N_866,N_838);
nand U937 (N_937,N_835,N_868);
or U938 (N_938,N_877,N_864);
nor U939 (N_939,N_854,N_837);
nor U940 (N_940,N_833,N_896);
nor U941 (N_941,N_855,N_827);
nor U942 (N_942,N_889,N_876);
and U943 (N_943,N_838,N_848);
and U944 (N_944,N_897,N_873);
or U945 (N_945,N_885,N_855);
nand U946 (N_946,N_859,N_841);
xnor U947 (N_947,N_854,N_886);
or U948 (N_948,N_860,N_897);
nor U949 (N_949,N_871,N_848);
nor U950 (N_950,N_854,N_893);
or U951 (N_951,N_899,N_865);
xor U952 (N_952,N_870,N_879);
or U953 (N_953,N_857,N_882);
and U954 (N_954,N_866,N_865);
or U955 (N_955,N_860,N_894);
nor U956 (N_956,N_885,N_892);
nand U957 (N_957,N_830,N_837);
nand U958 (N_958,N_873,N_874);
nor U959 (N_959,N_877,N_833);
and U960 (N_960,N_876,N_857);
nand U961 (N_961,N_855,N_869);
nor U962 (N_962,N_871,N_837);
nand U963 (N_963,N_871,N_832);
nand U964 (N_964,N_857,N_878);
nand U965 (N_965,N_878,N_889);
nand U966 (N_966,N_874,N_894);
nand U967 (N_967,N_839,N_881);
nand U968 (N_968,N_892,N_886);
or U969 (N_969,N_897,N_895);
nor U970 (N_970,N_843,N_893);
nand U971 (N_971,N_897,N_871);
nand U972 (N_972,N_851,N_890);
nor U973 (N_973,N_884,N_834);
nor U974 (N_974,N_845,N_852);
and U975 (N_975,N_909,N_939);
nor U976 (N_976,N_946,N_922);
nor U977 (N_977,N_917,N_953);
and U978 (N_978,N_918,N_964);
and U979 (N_979,N_940,N_910);
and U980 (N_980,N_923,N_961);
and U981 (N_981,N_904,N_958);
nand U982 (N_982,N_973,N_954);
nand U983 (N_983,N_934,N_941);
or U984 (N_984,N_960,N_949);
nor U985 (N_985,N_901,N_932);
and U986 (N_986,N_927,N_938);
and U987 (N_987,N_957,N_931);
and U988 (N_988,N_970,N_933);
or U989 (N_989,N_914,N_962);
nand U990 (N_990,N_921,N_928);
nand U991 (N_991,N_908,N_930);
or U992 (N_992,N_920,N_916);
nor U993 (N_993,N_965,N_900);
and U994 (N_994,N_935,N_903);
and U995 (N_995,N_956,N_974);
nor U996 (N_996,N_924,N_937);
or U997 (N_997,N_967,N_906);
or U998 (N_998,N_971,N_929);
nor U999 (N_999,N_936,N_951);
and U1000 (N_1000,N_911,N_972);
or U1001 (N_1001,N_905,N_942);
nor U1002 (N_1002,N_966,N_950);
nand U1003 (N_1003,N_959,N_926);
or U1004 (N_1004,N_943,N_947);
and U1005 (N_1005,N_919,N_952);
and U1006 (N_1006,N_913,N_955);
nand U1007 (N_1007,N_963,N_902);
nor U1008 (N_1008,N_925,N_945);
or U1009 (N_1009,N_907,N_912);
nand U1010 (N_1010,N_948,N_968);
nor U1011 (N_1011,N_944,N_915);
and U1012 (N_1012,N_969,N_918);
nand U1013 (N_1013,N_936,N_906);
and U1014 (N_1014,N_946,N_948);
nor U1015 (N_1015,N_947,N_932);
nor U1016 (N_1016,N_966,N_968);
nand U1017 (N_1017,N_969,N_913);
and U1018 (N_1018,N_955,N_942);
and U1019 (N_1019,N_942,N_912);
nand U1020 (N_1020,N_911,N_916);
nand U1021 (N_1021,N_906,N_958);
nand U1022 (N_1022,N_915,N_961);
or U1023 (N_1023,N_961,N_962);
nor U1024 (N_1024,N_916,N_923);
or U1025 (N_1025,N_935,N_929);
and U1026 (N_1026,N_970,N_956);
nor U1027 (N_1027,N_923,N_942);
or U1028 (N_1028,N_953,N_948);
nor U1029 (N_1029,N_970,N_946);
nand U1030 (N_1030,N_919,N_955);
nand U1031 (N_1031,N_911,N_959);
nand U1032 (N_1032,N_921,N_932);
nand U1033 (N_1033,N_905,N_967);
or U1034 (N_1034,N_912,N_961);
or U1035 (N_1035,N_947,N_962);
or U1036 (N_1036,N_913,N_962);
or U1037 (N_1037,N_901,N_924);
nor U1038 (N_1038,N_957,N_923);
nand U1039 (N_1039,N_919,N_970);
or U1040 (N_1040,N_969,N_967);
nor U1041 (N_1041,N_934,N_930);
nand U1042 (N_1042,N_940,N_905);
or U1043 (N_1043,N_934,N_903);
nand U1044 (N_1044,N_966,N_955);
or U1045 (N_1045,N_941,N_965);
or U1046 (N_1046,N_960,N_956);
nand U1047 (N_1047,N_964,N_930);
and U1048 (N_1048,N_934,N_927);
or U1049 (N_1049,N_927,N_948);
or U1050 (N_1050,N_990,N_1018);
nand U1051 (N_1051,N_1019,N_1012);
and U1052 (N_1052,N_1032,N_994);
and U1053 (N_1053,N_1003,N_1027);
or U1054 (N_1054,N_978,N_1004);
nor U1055 (N_1055,N_1011,N_982);
nand U1056 (N_1056,N_1008,N_980);
or U1057 (N_1057,N_998,N_1041);
nand U1058 (N_1058,N_1029,N_1006);
nor U1059 (N_1059,N_1015,N_1007);
and U1060 (N_1060,N_996,N_1013);
nor U1061 (N_1061,N_1024,N_981);
nor U1062 (N_1062,N_1047,N_993);
nor U1063 (N_1063,N_1000,N_1017);
xnor U1064 (N_1064,N_986,N_1028);
nand U1065 (N_1065,N_1002,N_987);
nand U1066 (N_1066,N_975,N_1040);
nor U1067 (N_1067,N_1045,N_995);
nand U1068 (N_1068,N_1014,N_1031);
nor U1069 (N_1069,N_1049,N_1001);
nand U1070 (N_1070,N_1034,N_1020);
or U1071 (N_1071,N_1036,N_1044);
or U1072 (N_1072,N_1038,N_985);
and U1073 (N_1073,N_1025,N_1039);
nor U1074 (N_1074,N_1035,N_1021);
or U1075 (N_1075,N_979,N_977);
or U1076 (N_1076,N_976,N_983);
nor U1077 (N_1077,N_984,N_1042);
or U1078 (N_1078,N_1048,N_992);
xor U1079 (N_1079,N_997,N_1010);
nand U1080 (N_1080,N_1046,N_991);
or U1081 (N_1081,N_999,N_1016);
nand U1082 (N_1082,N_1026,N_1037);
nor U1083 (N_1083,N_1022,N_1033);
or U1084 (N_1084,N_1005,N_1043);
nor U1085 (N_1085,N_1030,N_988);
or U1086 (N_1086,N_1023,N_1009);
nand U1087 (N_1087,N_989,N_1012);
nor U1088 (N_1088,N_1039,N_1045);
nor U1089 (N_1089,N_1015,N_988);
and U1090 (N_1090,N_1011,N_1047);
nor U1091 (N_1091,N_992,N_999);
nand U1092 (N_1092,N_1044,N_1019);
nand U1093 (N_1093,N_1041,N_1001);
and U1094 (N_1094,N_988,N_1028);
nand U1095 (N_1095,N_994,N_997);
nor U1096 (N_1096,N_976,N_1041);
and U1097 (N_1097,N_1029,N_1018);
and U1098 (N_1098,N_1033,N_1016);
and U1099 (N_1099,N_1025,N_1006);
and U1100 (N_1100,N_1043,N_996);
and U1101 (N_1101,N_994,N_976);
and U1102 (N_1102,N_988,N_1044);
nand U1103 (N_1103,N_1021,N_1048);
nor U1104 (N_1104,N_1008,N_1035);
and U1105 (N_1105,N_1012,N_1040);
and U1106 (N_1106,N_984,N_1019);
or U1107 (N_1107,N_1020,N_980);
nor U1108 (N_1108,N_1015,N_1028);
or U1109 (N_1109,N_1047,N_1032);
nand U1110 (N_1110,N_1019,N_991);
and U1111 (N_1111,N_1003,N_1034);
and U1112 (N_1112,N_1024,N_1034);
or U1113 (N_1113,N_977,N_992);
or U1114 (N_1114,N_1003,N_1028);
and U1115 (N_1115,N_992,N_981);
or U1116 (N_1116,N_1020,N_1015);
nor U1117 (N_1117,N_980,N_1027);
nor U1118 (N_1118,N_995,N_1046);
and U1119 (N_1119,N_1014,N_1005);
or U1120 (N_1120,N_1025,N_1009);
nand U1121 (N_1121,N_1047,N_1039);
or U1122 (N_1122,N_988,N_985);
or U1123 (N_1123,N_1049,N_985);
or U1124 (N_1124,N_994,N_1027);
nand U1125 (N_1125,N_1077,N_1088);
nand U1126 (N_1126,N_1124,N_1083);
and U1127 (N_1127,N_1116,N_1059);
and U1128 (N_1128,N_1056,N_1078);
nor U1129 (N_1129,N_1084,N_1118);
or U1130 (N_1130,N_1080,N_1066);
nor U1131 (N_1131,N_1121,N_1098);
nor U1132 (N_1132,N_1096,N_1061);
or U1133 (N_1133,N_1095,N_1090);
and U1134 (N_1134,N_1115,N_1107);
nand U1135 (N_1135,N_1091,N_1105);
nand U1136 (N_1136,N_1109,N_1120);
xnor U1137 (N_1137,N_1071,N_1075);
nand U1138 (N_1138,N_1073,N_1064);
or U1139 (N_1139,N_1108,N_1093);
or U1140 (N_1140,N_1122,N_1060);
nand U1141 (N_1141,N_1070,N_1099);
or U1142 (N_1142,N_1103,N_1062);
nand U1143 (N_1143,N_1111,N_1112);
and U1144 (N_1144,N_1089,N_1113);
and U1145 (N_1145,N_1097,N_1068);
nand U1146 (N_1146,N_1110,N_1094);
nor U1147 (N_1147,N_1058,N_1119);
or U1148 (N_1148,N_1052,N_1123);
nor U1149 (N_1149,N_1079,N_1072);
nand U1150 (N_1150,N_1102,N_1063);
or U1151 (N_1151,N_1067,N_1054);
or U1152 (N_1152,N_1114,N_1055);
nand U1153 (N_1153,N_1100,N_1117);
nor U1154 (N_1154,N_1082,N_1057);
nand U1155 (N_1155,N_1087,N_1081);
nand U1156 (N_1156,N_1053,N_1085);
and U1157 (N_1157,N_1050,N_1106);
or U1158 (N_1158,N_1086,N_1076);
and U1159 (N_1159,N_1104,N_1074);
and U1160 (N_1160,N_1065,N_1069);
and U1161 (N_1161,N_1051,N_1101);
nand U1162 (N_1162,N_1092,N_1117);
or U1163 (N_1163,N_1075,N_1123);
nor U1164 (N_1164,N_1114,N_1085);
or U1165 (N_1165,N_1096,N_1056);
and U1166 (N_1166,N_1052,N_1106);
and U1167 (N_1167,N_1072,N_1086);
nand U1168 (N_1168,N_1096,N_1121);
or U1169 (N_1169,N_1058,N_1107);
and U1170 (N_1170,N_1102,N_1099);
or U1171 (N_1171,N_1114,N_1086);
nand U1172 (N_1172,N_1112,N_1077);
nor U1173 (N_1173,N_1109,N_1071);
or U1174 (N_1174,N_1108,N_1110);
and U1175 (N_1175,N_1094,N_1073);
nand U1176 (N_1176,N_1120,N_1118);
nor U1177 (N_1177,N_1082,N_1121);
or U1178 (N_1178,N_1100,N_1082);
and U1179 (N_1179,N_1104,N_1089);
nand U1180 (N_1180,N_1070,N_1088);
or U1181 (N_1181,N_1066,N_1099);
and U1182 (N_1182,N_1087,N_1113);
or U1183 (N_1183,N_1077,N_1058);
nand U1184 (N_1184,N_1050,N_1081);
nand U1185 (N_1185,N_1065,N_1123);
or U1186 (N_1186,N_1101,N_1056);
and U1187 (N_1187,N_1064,N_1059);
nor U1188 (N_1188,N_1116,N_1120);
nand U1189 (N_1189,N_1122,N_1123);
nand U1190 (N_1190,N_1114,N_1084);
or U1191 (N_1191,N_1102,N_1070);
or U1192 (N_1192,N_1120,N_1110);
nor U1193 (N_1193,N_1067,N_1119);
nor U1194 (N_1194,N_1107,N_1117);
and U1195 (N_1195,N_1097,N_1073);
nor U1196 (N_1196,N_1096,N_1106);
nand U1197 (N_1197,N_1058,N_1078);
nand U1198 (N_1198,N_1123,N_1083);
nor U1199 (N_1199,N_1069,N_1057);
and U1200 (N_1200,N_1138,N_1145);
or U1201 (N_1201,N_1181,N_1152);
nor U1202 (N_1202,N_1158,N_1188);
and U1203 (N_1203,N_1160,N_1132);
or U1204 (N_1204,N_1161,N_1169);
and U1205 (N_1205,N_1146,N_1148);
or U1206 (N_1206,N_1156,N_1190);
nor U1207 (N_1207,N_1177,N_1143);
and U1208 (N_1208,N_1186,N_1163);
nand U1209 (N_1209,N_1151,N_1194);
nor U1210 (N_1210,N_1159,N_1171);
or U1211 (N_1211,N_1153,N_1135);
xor U1212 (N_1212,N_1165,N_1162);
nor U1213 (N_1213,N_1195,N_1166);
nor U1214 (N_1214,N_1189,N_1142);
and U1215 (N_1215,N_1140,N_1196);
and U1216 (N_1216,N_1136,N_1149);
and U1217 (N_1217,N_1179,N_1180);
nor U1218 (N_1218,N_1167,N_1150);
nor U1219 (N_1219,N_1198,N_1131);
and U1220 (N_1220,N_1176,N_1182);
and U1221 (N_1221,N_1178,N_1191);
nor U1222 (N_1222,N_1129,N_1141);
nand U1223 (N_1223,N_1187,N_1173);
and U1224 (N_1224,N_1168,N_1170);
xnor U1225 (N_1225,N_1175,N_1125);
nand U1226 (N_1226,N_1199,N_1185);
and U1227 (N_1227,N_1134,N_1126);
or U1228 (N_1228,N_1155,N_1192);
nand U1229 (N_1229,N_1197,N_1184);
or U1230 (N_1230,N_1157,N_1147);
nor U1231 (N_1231,N_1174,N_1139);
nand U1232 (N_1232,N_1154,N_1164);
nor U1233 (N_1233,N_1137,N_1127);
nand U1234 (N_1234,N_1128,N_1133);
nand U1235 (N_1235,N_1172,N_1193);
or U1236 (N_1236,N_1144,N_1130);
nor U1237 (N_1237,N_1183,N_1154);
or U1238 (N_1238,N_1182,N_1148);
nand U1239 (N_1239,N_1128,N_1146);
nand U1240 (N_1240,N_1128,N_1167);
and U1241 (N_1241,N_1139,N_1186);
nor U1242 (N_1242,N_1197,N_1165);
nand U1243 (N_1243,N_1150,N_1153);
nand U1244 (N_1244,N_1197,N_1178);
nor U1245 (N_1245,N_1197,N_1196);
nor U1246 (N_1246,N_1197,N_1170);
and U1247 (N_1247,N_1139,N_1160);
nand U1248 (N_1248,N_1131,N_1194);
nand U1249 (N_1249,N_1160,N_1190);
nor U1250 (N_1250,N_1195,N_1147);
nor U1251 (N_1251,N_1134,N_1142);
or U1252 (N_1252,N_1189,N_1187);
nor U1253 (N_1253,N_1135,N_1173);
nand U1254 (N_1254,N_1143,N_1154);
and U1255 (N_1255,N_1166,N_1158);
nand U1256 (N_1256,N_1170,N_1163);
or U1257 (N_1257,N_1154,N_1189);
and U1258 (N_1258,N_1158,N_1128);
nor U1259 (N_1259,N_1174,N_1170);
nor U1260 (N_1260,N_1126,N_1189);
nor U1261 (N_1261,N_1165,N_1138);
or U1262 (N_1262,N_1183,N_1174);
nand U1263 (N_1263,N_1186,N_1134);
nor U1264 (N_1264,N_1191,N_1190);
or U1265 (N_1265,N_1158,N_1195);
and U1266 (N_1266,N_1192,N_1199);
and U1267 (N_1267,N_1127,N_1167);
nor U1268 (N_1268,N_1196,N_1143);
nor U1269 (N_1269,N_1174,N_1176);
or U1270 (N_1270,N_1181,N_1172);
nand U1271 (N_1271,N_1173,N_1162);
or U1272 (N_1272,N_1152,N_1170);
nor U1273 (N_1273,N_1125,N_1156);
xor U1274 (N_1274,N_1154,N_1153);
and U1275 (N_1275,N_1204,N_1241);
nand U1276 (N_1276,N_1260,N_1229);
nor U1277 (N_1277,N_1265,N_1225);
nand U1278 (N_1278,N_1242,N_1267);
nand U1279 (N_1279,N_1201,N_1264);
or U1280 (N_1280,N_1254,N_1253);
and U1281 (N_1281,N_1250,N_1271);
xnor U1282 (N_1282,N_1247,N_1219);
and U1283 (N_1283,N_1212,N_1243);
and U1284 (N_1284,N_1262,N_1263);
nor U1285 (N_1285,N_1234,N_1266);
nor U1286 (N_1286,N_1249,N_1226);
nor U1287 (N_1287,N_1220,N_1270);
and U1288 (N_1288,N_1211,N_1223);
xnor U1289 (N_1289,N_1258,N_1269);
or U1290 (N_1290,N_1209,N_1235);
and U1291 (N_1291,N_1228,N_1206);
nand U1292 (N_1292,N_1213,N_1268);
nand U1293 (N_1293,N_1240,N_1200);
nor U1294 (N_1294,N_1214,N_1256);
and U1295 (N_1295,N_1272,N_1218);
nor U1296 (N_1296,N_1224,N_1216);
nand U1297 (N_1297,N_1274,N_1207);
nor U1298 (N_1298,N_1248,N_1205);
or U1299 (N_1299,N_1221,N_1233);
nand U1300 (N_1300,N_1230,N_1255);
nand U1301 (N_1301,N_1239,N_1244);
and U1302 (N_1302,N_1232,N_1208);
nor U1303 (N_1303,N_1217,N_1257);
nand U1304 (N_1304,N_1203,N_1210);
nor U1305 (N_1305,N_1259,N_1238);
nor U1306 (N_1306,N_1227,N_1222);
nor U1307 (N_1307,N_1261,N_1202);
nand U1308 (N_1308,N_1231,N_1237);
xnor U1309 (N_1309,N_1246,N_1251);
nor U1310 (N_1310,N_1245,N_1252);
or U1311 (N_1311,N_1215,N_1236);
or U1312 (N_1312,N_1273,N_1203);
and U1313 (N_1313,N_1257,N_1249);
nor U1314 (N_1314,N_1255,N_1221);
nor U1315 (N_1315,N_1242,N_1248);
nor U1316 (N_1316,N_1274,N_1243);
and U1317 (N_1317,N_1263,N_1261);
or U1318 (N_1318,N_1242,N_1230);
and U1319 (N_1319,N_1230,N_1221);
and U1320 (N_1320,N_1222,N_1217);
nor U1321 (N_1321,N_1223,N_1234);
nand U1322 (N_1322,N_1264,N_1257);
nor U1323 (N_1323,N_1237,N_1267);
nand U1324 (N_1324,N_1245,N_1214);
or U1325 (N_1325,N_1205,N_1245);
and U1326 (N_1326,N_1234,N_1256);
nand U1327 (N_1327,N_1271,N_1213);
and U1328 (N_1328,N_1253,N_1274);
nor U1329 (N_1329,N_1258,N_1219);
and U1330 (N_1330,N_1230,N_1234);
nand U1331 (N_1331,N_1248,N_1240);
nand U1332 (N_1332,N_1236,N_1214);
nand U1333 (N_1333,N_1207,N_1263);
or U1334 (N_1334,N_1258,N_1206);
nor U1335 (N_1335,N_1263,N_1238);
or U1336 (N_1336,N_1212,N_1248);
and U1337 (N_1337,N_1224,N_1239);
and U1338 (N_1338,N_1239,N_1241);
nand U1339 (N_1339,N_1268,N_1226);
and U1340 (N_1340,N_1231,N_1258);
and U1341 (N_1341,N_1207,N_1258);
and U1342 (N_1342,N_1233,N_1246);
and U1343 (N_1343,N_1261,N_1255);
nand U1344 (N_1344,N_1234,N_1219);
nor U1345 (N_1345,N_1239,N_1247);
or U1346 (N_1346,N_1207,N_1245);
nor U1347 (N_1347,N_1205,N_1214);
or U1348 (N_1348,N_1205,N_1250);
nand U1349 (N_1349,N_1239,N_1267);
and U1350 (N_1350,N_1306,N_1305);
nand U1351 (N_1351,N_1283,N_1320);
or U1352 (N_1352,N_1293,N_1318);
nand U1353 (N_1353,N_1280,N_1289);
nand U1354 (N_1354,N_1323,N_1346);
nand U1355 (N_1355,N_1331,N_1281);
or U1356 (N_1356,N_1297,N_1302);
nor U1357 (N_1357,N_1304,N_1348);
or U1358 (N_1358,N_1300,N_1335);
nor U1359 (N_1359,N_1326,N_1285);
or U1360 (N_1360,N_1347,N_1310);
or U1361 (N_1361,N_1311,N_1340);
and U1362 (N_1362,N_1288,N_1343);
nor U1363 (N_1363,N_1315,N_1301);
nand U1364 (N_1364,N_1322,N_1278);
nor U1365 (N_1365,N_1342,N_1345);
nand U1366 (N_1366,N_1336,N_1314);
and U1367 (N_1367,N_1286,N_1308);
and U1368 (N_1368,N_1282,N_1338);
nand U1369 (N_1369,N_1333,N_1287);
and U1370 (N_1370,N_1324,N_1341);
nor U1371 (N_1371,N_1316,N_1313);
or U1372 (N_1372,N_1344,N_1327);
or U1373 (N_1373,N_1298,N_1339);
nor U1374 (N_1374,N_1312,N_1307);
nor U1375 (N_1375,N_1334,N_1309);
nand U1376 (N_1376,N_1329,N_1317);
or U1377 (N_1377,N_1290,N_1294);
or U1378 (N_1378,N_1279,N_1330);
or U1379 (N_1379,N_1277,N_1284);
xnor U1380 (N_1380,N_1325,N_1295);
or U1381 (N_1381,N_1328,N_1349);
nand U1382 (N_1382,N_1332,N_1303);
or U1383 (N_1383,N_1296,N_1291);
and U1384 (N_1384,N_1337,N_1299);
or U1385 (N_1385,N_1276,N_1275);
nor U1386 (N_1386,N_1321,N_1292);
nor U1387 (N_1387,N_1319,N_1315);
nor U1388 (N_1388,N_1339,N_1303);
nand U1389 (N_1389,N_1343,N_1345);
xor U1390 (N_1390,N_1296,N_1323);
and U1391 (N_1391,N_1302,N_1325);
nand U1392 (N_1392,N_1305,N_1341);
and U1393 (N_1393,N_1282,N_1281);
nor U1394 (N_1394,N_1275,N_1306);
or U1395 (N_1395,N_1313,N_1320);
nand U1396 (N_1396,N_1340,N_1278);
nor U1397 (N_1397,N_1275,N_1322);
and U1398 (N_1398,N_1333,N_1275);
nand U1399 (N_1399,N_1348,N_1335);
xnor U1400 (N_1400,N_1348,N_1334);
nor U1401 (N_1401,N_1347,N_1281);
and U1402 (N_1402,N_1313,N_1327);
or U1403 (N_1403,N_1334,N_1320);
or U1404 (N_1404,N_1348,N_1276);
or U1405 (N_1405,N_1334,N_1340);
and U1406 (N_1406,N_1302,N_1282);
or U1407 (N_1407,N_1284,N_1288);
nor U1408 (N_1408,N_1305,N_1321);
and U1409 (N_1409,N_1298,N_1284);
nand U1410 (N_1410,N_1297,N_1296);
nor U1411 (N_1411,N_1309,N_1281);
and U1412 (N_1412,N_1305,N_1340);
nand U1413 (N_1413,N_1343,N_1281);
nor U1414 (N_1414,N_1297,N_1279);
nand U1415 (N_1415,N_1344,N_1296);
and U1416 (N_1416,N_1348,N_1337);
and U1417 (N_1417,N_1292,N_1286);
nor U1418 (N_1418,N_1284,N_1330);
nor U1419 (N_1419,N_1314,N_1285);
nor U1420 (N_1420,N_1307,N_1339);
or U1421 (N_1421,N_1326,N_1279);
and U1422 (N_1422,N_1287,N_1324);
and U1423 (N_1423,N_1282,N_1291);
nor U1424 (N_1424,N_1349,N_1325);
and U1425 (N_1425,N_1356,N_1397);
and U1426 (N_1426,N_1355,N_1422);
nor U1427 (N_1427,N_1391,N_1409);
nand U1428 (N_1428,N_1367,N_1423);
nor U1429 (N_1429,N_1373,N_1402);
and U1430 (N_1430,N_1384,N_1410);
or U1431 (N_1431,N_1379,N_1383);
or U1432 (N_1432,N_1357,N_1366);
nor U1433 (N_1433,N_1370,N_1380);
and U1434 (N_1434,N_1351,N_1418);
nand U1435 (N_1435,N_1419,N_1407);
nand U1436 (N_1436,N_1360,N_1396);
nor U1437 (N_1437,N_1361,N_1414);
nand U1438 (N_1438,N_1395,N_1353);
or U1439 (N_1439,N_1392,N_1421);
and U1440 (N_1440,N_1389,N_1401);
nor U1441 (N_1441,N_1404,N_1381);
xnor U1442 (N_1442,N_1376,N_1374);
or U1443 (N_1443,N_1385,N_1413);
or U1444 (N_1444,N_1406,N_1368);
or U1445 (N_1445,N_1375,N_1350);
nor U1446 (N_1446,N_1371,N_1382);
nor U1447 (N_1447,N_1387,N_1352);
and U1448 (N_1448,N_1363,N_1393);
or U1449 (N_1449,N_1359,N_1369);
nand U1450 (N_1450,N_1394,N_1354);
and U1451 (N_1451,N_1411,N_1417);
and U1452 (N_1452,N_1388,N_1378);
and U1453 (N_1453,N_1358,N_1424);
nand U1454 (N_1454,N_1364,N_1412);
nand U1455 (N_1455,N_1400,N_1365);
or U1456 (N_1456,N_1390,N_1405);
nor U1457 (N_1457,N_1420,N_1386);
nand U1458 (N_1458,N_1408,N_1416);
nor U1459 (N_1459,N_1398,N_1415);
nand U1460 (N_1460,N_1372,N_1362);
or U1461 (N_1461,N_1377,N_1399);
or U1462 (N_1462,N_1403,N_1376);
and U1463 (N_1463,N_1359,N_1384);
or U1464 (N_1464,N_1413,N_1350);
or U1465 (N_1465,N_1397,N_1382);
or U1466 (N_1466,N_1397,N_1369);
or U1467 (N_1467,N_1374,N_1359);
nor U1468 (N_1468,N_1394,N_1403);
nor U1469 (N_1469,N_1386,N_1378);
xor U1470 (N_1470,N_1415,N_1411);
nand U1471 (N_1471,N_1382,N_1357);
nor U1472 (N_1472,N_1365,N_1383);
and U1473 (N_1473,N_1413,N_1352);
or U1474 (N_1474,N_1350,N_1354);
nor U1475 (N_1475,N_1356,N_1423);
nand U1476 (N_1476,N_1402,N_1390);
nand U1477 (N_1477,N_1376,N_1413);
or U1478 (N_1478,N_1409,N_1376);
or U1479 (N_1479,N_1417,N_1373);
nand U1480 (N_1480,N_1381,N_1396);
or U1481 (N_1481,N_1353,N_1396);
nor U1482 (N_1482,N_1407,N_1406);
and U1483 (N_1483,N_1372,N_1398);
nand U1484 (N_1484,N_1385,N_1424);
and U1485 (N_1485,N_1420,N_1413);
nor U1486 (N_1486,N_1356,N_1374);
nand U1487 (N_1487,N_1382,N_1360);
and U1488 (N_1488,N_1362,N_1350);
or U1489 (N_1489,N_1351,N_1353);
or U1490 (N_1490,N_1355,N_1382);
nand U1491 (N_1491,N_1366,N_1352);
nand U1492 (N_1492,N_1403,N_1395);
nand U1493 (N_1493,N_1391,N_1358);
nand U1494 (N_1494,N_1408,N_1411);
or U1495 (N_1495,N_1353,N_1414);
nor U1496 (N_1496,N_1391,N_1381);
nand U1497 (N_1497,N_1392,N_1397);
or U1498 (N_1498,N_1353,N_1400);
or U1499 (N_1499,N_1371,N_1402);
nand U1500 (N_1500,N_1499,N_1463);
and U1501 (N_1501,N_1455,N_1437);
and U1502 (N_1502,N_1473,N_1439);
xnor U1503 (N_1503,N_1445,N_1426);
nand U1504 (N_1504,N_1496,N_1497);
or U1505 (N_1505,N_1476,N_1478);
or U1506 (N_1506,N_1470,N_1468);
nand U1507 (N_1507,N_1480,N_1490);
nor U1508 (N_1508,N_1438,N_1488);
and U1509 (N_1509,N_1435,N_1475);
and U1510 (N_1510,N_1450,N_1456);
or U1511 (N_1511,N_1493,N_1431);
xnor U1512 (N_1512,N_1447,N_1443);
and U1513 (N_1513,N_1494,N_1440);
and U1514 (N_1514,N_1451,N_1489);
nand U1515 (N_1515,N_1425,N_1474);
and U1516 (N_1516,N_1472,N_1464);
or U1517 (N_1517,N_1477,N_1481);
nor U1518 (N_1518,N_1498,N_1457);
nand U1519 (N_1519,N_1479,N_1466);
nor U1520 (N_1520,N_1449,N_1429);
or U1521 (N_1521,N_1492,N_1483);
nand U1522 (N_1522,N_1487,N_1486);
nor U1523 (N_1523,N_1465,N_1441);
and U1524 (N_1524,N_1458,N_1471);
nand U1525 (N_1525,N_1461,N_1467);
or U1526 (N_1526,N_1448,N_1446);
nand U1527 (N_1527,N_1460,N_1442);
and U1528 (N_1528,N_1469,N_1453);
nor U1529 (N_1529,N_1427,N_1482);
and U1530 (N_1530,N_1454,N_1495);
and U1531 (N_1531,N_1452,N_1459);
nor U1532 (N_1532,N_1484,N_1485);
nor U1533 (N_1533,N_1430,N_1436);
and U1534 (N_1534,N_1433,N_1428);
and U1535 (N_1535,N_1462,N_1444);
or U1536 (N_1536,N_1432,N_1491);
nor U1537 (N_1537,N_1434,N_1459);
and U1538 (N_1538,N_1472,N_1435);
nor U1539 (N_1539,N_1438,N_1485);
nor U1540 (N_1540,N_1495,N_1460);
and U1541 (N_1541,N_1426,N_1478);
nand U1542 (N_1542,N_1450,N_1499);
nor U1543 (N_1543,N_1428,N_1472);
xor U1544 (N_1544,N_1470,N_1464);
nand U1545 (N_1545,N_1457,N_1443);
and U1546 (N_1546,N_1476,N_1446);
or U1547 (N_1547,N_1469,N_1495);
nand U1548 (N_1548,N_1428,N_1477);
nor U1549 (N_1549,N_1425,N_1484);
nand U1550 (N_1550,N_1463,N_1467);
nor U1551 (N_1551,N_1497,N_1472);
and U1552 (N_1552,N_1465,N_1449);
or U1553 (N_1553,N_1432,N_1486);
or U1554 (N_1554,N_1481,N_1475);
or U1555 (N_1555,N_1489,N_1452);
or U1556 (N_1556,N_1425,N_1497);
nor U1557 (N_1557,N_1456,N_1490);
nand U1558 (N_1558,N_1445,N_1483);
xnor U1559 (N_1559,N_1448,N_1440);
nor U1560 (N_1560,N_1466,N_1477);
or U1561 (N_1561,N_1462,N_1450);
and U1562 (N_1562,N_1464,N_1484);
nand U1563 (N_1563,N_1481,N_1461);
xor U1564 (N_1564,N_1429,N_1478);
or U1565 (N_1565,N_1494,N_1450);
and U1566 (N_1566,N_1482,N_1462);
xor U1567 (N_1567,N_1430,N_1460);
nor U1568 (N_1568,N_1478,N_1450);
and U1569 (N_1569,N_1466,N_1446);
xor U1570 (N_1570,N_1465,N_1491);
nand U1571 (N_1571,N_1499,N_1490);
and U1572 (N_1572,N_1491,N_1445);
nand U1573 (N_1573,N_1472,N_1481);
nor U1574 (N_1574,N_1454,N_1496);
or U1575 (N_1575,N_1539,N_1518);
nor U1576 (N_1576,N_1541,N_1546);
nor U1577 (N_1577,N_1528,N_1517);
nand U1578 (N_1578,N_1505,N_1534);
nor U1579 (N_1579,N_1562,N_1551);
or U1580 (N_1580,N_1511,N_1557);
or U1581 (N_1581,N_1533,N_1535);
nor U1582 (N_1582,N_1516,N_1508);
xor U1583 (N_1583,N_1564,N_1553);
and U1584 (N_1584,N_1544,N_1568);
and U1585 (N_1585,N_1526,N_1566);
and U1586 (N_1586,N_1567,N_1554);
and U1587 (N_1587,N_1561,N_1545);
or U1588 (N_1588,N_1525,N_1565);
xnor U1589 (N_1589,N_1530,N_1513);
or U1590 (N_1590,N_1570,N_1512);
xor U1591 (N_1591,N_1569,N_1572);
xnor U1592 (N_1592,N_1522,N_1531);
and U1593 (N_1593,N_1515,N_1571);
or U1594 (N_1594,N_1519,N_1556);
nor U1595 (N_1595,N_1560,N_1559);
nor U1596 (N_1596,N_1550,N_1547);
or U1597 (N_1597,N_1548,N_1521);
and U1598 (N_1598,N_1563,N_1523);
nand U1599 (N_1599,N_1574,N_1501);
and U1600 (N_1600,N_1507,N_1543);
nor U1601 (N_1601,N_1527,N_1573);
xnor U1602 (N_1602,N_1500,N_1558);
nor U1603 (N_1603,N_1509,N_1542);
nor U1604 (N_1604,N_1552,N_1524);
nor U1605 (N_1605,N_1538,N_1514);
or U1606 (N_1606,N_1504,N_1529);
and U1607 (N_1607,N_1532,N_1540);
nor U1608 (N_1608,N_1502,N_1520);
nor U1609 (N_1609,N_1549,N_1537);
and U1610 (N_1610,N_1555,N_1536);
nand U1611 (N_1611,N_1506,N_1510);
and U1612 (N_1612,N_1503,N_1513);
and U1613 (N_1613,N_1519,N_1512);
or U1614 (N_1614,N_1521,N_1507);
and U1615 (N_1615,N_1539,N_1542);
or U1616 (N_1616,N_1555,N_1521);
or U1617 (N_1617,N_1563,N_1507);
nand U1618 (N_1618,N_1502,N_1551);
and U1619 (N_1619,N_1574,N_1548);
nand U1620 (N_1620,N_1570,N_1566);
or U1621 (N_1621,N_1566,N_1517);
and U1622 (N_1622,N_1547,N_1563);
nor U1623 (N_1623,N_1566,N_1500);
or U1624 (N_1624,N_1535,N_1551);
nor U1625 (N_1625,N_1537,N_1553);
or U1626 (N_1626,N_1559,N_1572);
or U1627 (N_1627,N_1508,N_1529);
and U1628 (N_1628,N_1553,N_1522);
or U1629 (N_1629,N_1573,N_1502);
nor U1630 (N_1630,N_1529,N_1546);
or U1631 (N_1631,N_1536,N_1551);
nor U1632 (N_1632,N_1527,N_1507);
and U1633 (N_1633,N_1538,N_1574);
or U1634 (N_1634,N_1550,N_1509);
nor U1635 (N_1635,N_1521,N_1516);
or U1636 (N_1636,N_1574,N_1530);
nor U1637 (N_1637,N_1540,N_1553);
nand U1638 (N_1638,N_1504,N_1525);
and U1639 (N_1639,N_1518,N_1543);
and U1640 (N_1640,N_1531,N_1501);
or U1641 (N_1641,N_1537,N_1539);
nand U1642 (N_1642,N_1549,N_1554);
nand U1643 (N_1643,N_1528,N_1500);
and U1644 (N_1644,N_1502,N_1544);
nand U1645 (N_1645,N_1573,N_1532);
and U1646 (N_1646,N_1527,N_1520);
nor U1647 (N_1647,N_1562,N_1508);
nor U1648 (N_1648,N_1565,N_1514);
nand U1649 (N_1649,N_1543,N_1521);
nand U1650 (N_1650,N_1631,N_1577);
xor U1651 (N_1651,N_1600,N_1592);
nand U1652 (N_1652,N_1637,N_1638);
nor U1653 (N_1653,N_1587,N_1628);
and U1654 (N_1654,N_1601,N_1616);
and U1655 (N_1655,N_1639,N_1581);
nand U1656 (N_1656,N_1645,N_1619);
and U1657 (N_1657,N_1585,N_1648);
and U1658 (N_1658,N_1591,N_1612);
or U1659 (N_1659,N_1609,N_1580);
nor U1660 (N_1660,N_1633,N_1644);
nand U1661 (N_1661,N_1588,N_1596);
nand U1662 (N_1662,N_1636,N_1625);
or U1663 (N_1663,N_1576,N_1590);
nand U1664 (N_1664,N_1640,N_1621);
or U1665 (N_1665,N_1603,N_1589);
or U1666 (N_1666,N_1606,N_1630);
and U1667 (N_1667,N_1643,N_1626);
or U1668 (N_1668,N_1594,N_1623);
nand U1669 (N_1669,N_1614,N_1624);
and U1670 (N_1670,N_1646,N_1611);
and U1671 (N_1671,N_1610,N_1598);
and U1672 (N_1672,N_1613,N_1632);
nand U1673 (N_1673,N_1647,N_1575);
nor U1674 (N_1674,N_1583,N_1627);
and U1675 (N_1675,N_1617,N_1602);
nand U1676 (N_1676,N_1641,N_1642);
and U1677 (N_1677,N_1615,N_1620);
nor U1678 (N_1678,N_1599,N_1579);
nor U1679 (N_1679,N_1593,N_1586);
and U1680 (N_1680,N_1635,N_1595);
nor U1681 (N_1681,N_1629,N_1604);
nor U1682 (N_1682,N_1608,N_1584);
or U1683 (N_1683,N_1582,N_1634);
or U1684 (N_1684,N_1618,N_1597);
or U1685 (N_1685,N_1578,N_1622);
or U1686 (N_1686,N_1649,N_1605);
and U1687 (N_1687,N_1607,N_1595);
nor U1688 (N_1688,N_1605,N_1599);
nor U1689 (N_1689,N_1628,N_1593);
and U1690 (N_1690,N_1620,N_1604);
nand U1691 (N_1691,N_1598,N_1618);
and U1692 (N_1692,N_1594,N_1622);
nand U1693 (N_1693,N_1615,N_1604);
nand U1694 (N_1694,N_1614,N_1587);
or U1695 (N_1695,N_1639,N_1629);
nor U1696 (N_1696,N_1593,N_1594);
or U1697 (N_1697,N_1599,N_1587);
nand U1698 (N_1698,N_1622,N_1586);
or U1699 (N_1699,N_1643,N_1625);
and U1700 (N_1700,N_1583,N_1643);
nor U1701 (N_1701,N_1584,N_1648);
nor U1702 (N_1702,N_1647,N_1593);
nand U1703 (N_1703,N_1628,N_1627);
nor U1704 (N_1704,N_1631,N_1639);
and U1705 (N_1705,N_1580,N_1590);
nor U1706 (N_1706,N_1640,N_1636);
nand U1707 (N_1707,N_1636,N_1577);
and U1708 (N_1708,N_1583,N_1617);
or U1709 (N_1709,N_1609,N_1642);
or U1710 (N_1710,N_1576,N_1597);
nor U1711 (N_1711,N_1632,N_1584);
and U1712 (N_1712,N_1639,N_1628);
nor U1713 (N_1713,N_1609,N_1634);
or U1714 (N_1714,N_1576,N_1621);
and U1715 (N_1715,N_1592,N_1638);
nand U1716 (N_1716,N_1644,N_1608);
xor U1717 (N_1717,N_1645,N_1626);
nand U1718 (N_1718,N_1597,N_1610);
or U1719 (N_1719,N_1630,N_1600);
nand U1720 (N_1720,N_1629,N_1615);
nor U1721 (N_1721,N_1628,N_1624);
nand U1722 (N_1722,N_1586,N_1641);
nand U1723 (N_1723,N_1629,N_1575);
and U1724 (N_1724,N_1644,N_1647);
and U1725 (N_1725,N_1659,N_1658);
or U1726 (N_1726,N_1720,N_1655);
nor U1727 (N_1727,N_1722,N_1666);
nand U1728 (N_1728,N_1709,N_1690);
or U1729 (N_1729,N_1676,N_1703);
or U1730 (N_1730,N_1686,N_1724);
nor U1731 (N_1731,N_1717,N_1693);
nor U1732 (N_1732,N_1670,N_1669);
or U1733 (N_1733,N_1654,N_1691);
xor U1734 (N_1734,N_1663,N_1678);
and U1735 (N_1735,N_1701,N_1680);
nand U1736 (N_1736,N_1721,N_1697);
nor U1737 (N_1737,N_1675,N_1651);
nand U1738 (N_1738,N_1660,N_1707);
and U1739 (N_1739,N_1662,N_1677);
nor U1740 (N_1740,N_1711,N_1712);
and U1741 (N_1741,N_1705,N_1661);
or U1742 (N_1742,N_1664,N_1653);
nor U1743 (N_1743,N_1665,N_1679);
nand U1744 (N_1744,N_1708,N_1650);
or U1745 (N_1745,N_1674,N_1683);
nor U1746 (N_1746,N_1723,N_1699);
and U1747 (N_1747,N_1704,N_1688);
and U1748 (N_1748,N_1713,N_1682);
and U1749 (N_1749,N_1718,N_1716);
xor U1750 (N_1750,N_1698,N_1692);
and U1751 (N_1751,N_1710,N_1694);
or U1752 (N_1752,N_1700,N_1652);
nand U1753 (N_1753,N_1673,N_1685);
nor U1754 (N_1754,N_1696,N_1719);
or U1755 (N_1755,N_1715,N_1702);
or U1756 (N_1756,N_1687,N_1681);
or U1757 (N_1757,N_1689,N_1668);
nand U1758 (N_1758,N_1667,N_1656);
nor U1759 (N_1759,N_1684,N_1714);
nor U1760 (N_1760,N_1657,N_1695);
and U1761 (N_1761,N_1672,N_1706);
nand U1762 (N_1762,N_1671,N_1657);
and U1763 (N_1763,N_1722,N_1711);
nor U1764 (N_1764,N_1677,N_1703);
and U1765 (N_1765,N_1679,N_1690);
and U1766 (N_1766,N_1721,N_1656);
and U1767 (N_1767,N_1724,N_1675);
nand U1768 (N_1768,N_1668,N_1654);
xor U1769 (N_1769,N_1665,N_1689);
or U1770 (N_1770,N_1713,N_1673);
and U1771 (N_1771,N_1703,N_1717);
nor U1772 (N_1772,N_1680,N_1677);
and U1773 (N_1773,N_1694,N_1697);
or U1774 (N_1774,N_1692,N_1697);
or U1775 (N_1775,N_1672,N_1693);
and U1776 (N_1776,N_1650,N_1694);
or U1777 (N_1777,N_1678,N_1667);
or U1778 (N_1778,N_1655,N_1694);
or U1779 (N_1779,N_1685,N_1680);
or U1780 (N_1780,N_1697,N_1706);
nand U1781 (N_1781,N_1723,N_1703);
nand U1782 (N_1782,N_1688,N_1717);
and U1783 (N_1783,N_1666,N_1673);
and U1784 (N_1784,N_1674,N_1671);
nand U1785 (N_1785,N_1711,N_1671);
nor U1786 (N_1786,N_1695,N_1668);
and U1787 (N_1787,N_1701,N_1679);
nor U1788 (N_1788,N_1699,N_1703);
nand U1789 (N_1789,N_1710,N_1684);
nor U1790 (N_1790,N_1683,N_1669);
nand U1791 (N_1791,N_1721,N_1676);
xnor U1792 (N_1792,N_1683,N_1670);
and U1793 (N_1793,N_1670,N_1664);
nand U1794 (N_1794,N_1694,N_1671);
nor U1795 (N_1795,N_1715,N_1720);
nor U1796 (N_1796,N_1681,N_1704);
nor U1797 (N_1797,N_1682,N_1708);
and U1798 (N_1798,N_1682,N_1691);
nor U1799 (N_1799,N_1708,N_1674);
nand U1800 (N_1800,N_1739,N_1783);
or U1801 (N_1801,N_1795,N_1777);
nor U1802 (N_1802,N_1779,N_1760);
or U1803 (N_1803,N_1749,N_1794);
nor U1804 (N_1804,N_1731,N_1727);
or U1805 (N_1805,N_1754,N_1756);
and U1806 (N_1806,N_1791,N_1757);
nor U1807 (N_1807,N_1736,N_1730);
nand U1808 (N_1808,N_1781,N_1780);
or U1809 (N_1809,N_1776,N_1796);
nand U1810 (N_1810,N_1774,N_1744);
nand U1811 (N_1811,N_1798,N_1759);
nand U1812 (N_1812,N_1789,N_1747);
and U1813 (N_1813,N_1799,N_1743);
and U1814 (N_1814,N_1786,N_1793);
nor U1815 (N_1815,N_1742,N_1770);
nor U1816 (N_1816,N_1792,N_1761);
and U1817 (N_1817,N_1773,N_1766);
or U1818 (N_1818,N_1729,N_1772);
or U1819 (N_1819,N_1763,N_1734);
and U1820 (N_1820,N_1737,N_1728);
nor U1821 (N_1821,N_1725,N_1765);
or U1822 (N_1822,N_1769,N_1785);
nand U1823 (N_1823,N_1788,N_1751);
and U1824 (N_1824,N_1745,N_1775);
or U1825 (N_1825,N_1735,N_1771);
nand U1826 (N_1826,N_1738,N_1748);
nand U1827 (N_1827,N_1746,N_1733);
or U1828 (N_1828,N_1732,N_1782);
nor U1829 (N_1829,N_1740,N_1750);
nand U1830 (N_1830,N_1768,N_1778);
nand U1831 (N_1831,N_1758,N_1741);
nor U1832 (N_1832,N_1755,N_1753);
or U1833 (N_1833,N_1752,N_1784);
nor U1834 (N_1834,N_1762,N_1726);
or U1835 (N_1835,N_1790,N_1764);
nand U1836 (N_1836,N_1797,N_1787);
and U1837 (N_1837,N_1767,N_1784);
nand U1838 (N_1838,N_1767,N_1799);
nor U1839 (N_1839,N_1741,N_1779);
or U1840 (N_1840,N_1789,N_1777);
or U1841 (N_1841,N_1775,N_1748);
nand U1842 (N_1842,N_1763,N_1768);
nand U1843 (N_1843,N_1755,N_1763);
or U1844 (N_1844,N_1741,N_1797);
or U1845 (N_1845,N_1769,N_1743);
nand U1846 (N_1846,N_1742,N_1732);
nor U1847 (N_1847,N_1799,N_1779);
nor U1848 (N_1848,N_1743,N_1747);
or U1849 (N_1849,N_1733,N_1743);
nand U1850 (N_1850,N_1788,N_1768);
nand U1851 (N_1851,N_1763,N_1775);
or U1852 (N_1852,N_1766,N_1738);
and U1853 (N_1853,N_1784,N_1759);
nor U1854 (N_1854,N_1778,N_1747);
or U1855 (N_1855,N_1753,N_1779);
nand U1856 (N_1856,N_1751,N_1767);
and U1857 (N_1857,N_1751,N_1781);
or U1858 (N_1858,N_1743,N_1744);
and U1859 (N_1859,N_1771,N_1744);
and U1860 (N_1860,N_1735,N_1763);
or U1861 (N_1861,N_1748,N_1729);
and U1862 (N_1862,N_1738,N_1759);
nand U1863 (N_1863,N_1751,N_1735);
nand U1864 (N_1864,N_1748,N_1733);
nor U1865 (N_1865,N_1790,N_1786);
nand U1866 (N_1866,N_1753,N_1730);
nand U1867 (N_1867,N_1780,N_1774);
nand U1868 (N_1868,N_1740,N_1749);
nor U1869 (N_1869,N_1770,N_1767);
nand U1870 (N_1870,N_1747,N_1728);
nor U1871 (N_1871,N_1792,N_1791);
nand U1872 (N_1872,N_1798,N_1784);
nor U1873 (N_1873,N_1771,N_1784);
or U1874 (N_1874,N_1783,N_1766);
or U1875 (N_1875,N_1863,N_1872);
and U1876 (N_1876,N_1827,N_1823);
or U1877 (N_1877,N_1836,N_1853);
nand U1878 (N_1878,N_1818,N_1860);
and U1879 (N_1879,N_1847,N_1832);
nand U1880 (N_1880,N_1819,N_1870);
and U1881 (N_1881,N_1825,N_1810);
nand U1882 (N_1882,N_1854,N_1817);
and U1883 (N_1883,N_1822,N_1816);
nor U1884 (N_1884,N_1852,N_1844);
nor U1885 (N_1885,N_1857,N_1862);
or U1886 (N_1886,N_1807,N_1831);
nand U1887 (N_1887,N_1874,N_1843);
nor U1888 (N_1888,N_1841,N_1855);
or U1889 (N_1889,N_1833,N_1806);
or U1890 (N_1890,N_1829,N_1835);
nor U1891 (N_1891,N_1856,N_1808);
or U1892 (N_1892,N_1842,N_1809);
and U1893 (N_1893,N_1820,N_1802);
nor U1894 (N_1894,N_1858,N_1848);
or U1895 (N_1895,N_1826,N_1830);
and U1896 (N_1896,N_1851,N_1850);
nand U1897 (N_1897,N_1867,N_1821);
nand U1898 (N_1898,N_1804,N_1800);
nand U1899 (N_1899,N_1846,N_1861);
nor U1900 (N_1900,N_1837,N_1801);
or U1901 (N_1901,N_1840,N_1813);
and U1902 (N_1902,N_1871,N_1811);
or U1903 (N_1903,N_1812,N_1834);
nand U1904 (N_1904,N_1849,N_1828);
and U1905 (N_1905,N_1814,N_1865);
and U1906 (N_1906,N_1815,N_1803);
nand U1907 (N_1907,N_1868,N_1805);
nor U1908 (N_1908,N_1866,N_1839);
nor U1909 (N_1909,N_1845,N_1838);
nor U1910 (N_1910,N_1869,N_1859);
or U1911 (N_1911,N_1864,N_1824);
or U1912 (N_1912,N_1873,N_1854);
and U1913 (N_1913,N_1818,N_1816);
and U1914 (N_1914,N_1805,N_1870);
or U1915 (N_1915,N_1830,N_1813);
and U1916 (N_1916,N_1852,N_1861);
or U1917 (N_1917,N_1823,N_1836);
nor U1918 (N_1918,N_1855,N_1838);
xor U1919 (N_1919,N_1826,N_1848);
nor U1920 (N_1920,N_1841,N_1808);
nand U1921 (N_1921,N_1872,N_1805);
nand U1922 (N_1922,N_1836,N_1818);
and U1923 (N_1923,N_1829,N_1810);
and U1924 (N_1924,N_1863,N_1822);
nor U1925 (N_1925,N_1834,N_1804);
nor U1926 (N_1926,N_1858,N_1821);
and U1927 (N_1927,N_1849,N_1873);
nor U1928 (N_1928,N_1873,N_1830);
nand U1929 (N_1929,N_1811,N_1870);
and U1930 (N_1930,N_1807,N_1862);
or U1931 (N_1931,N_1840,N_1873);
nand U1932 (N_1932,N_1801,N_1817);
nand U1933 (N_1933,N_1829,N_1825);
nand U1934 (N_1934,N_1872,N_1865);
or U1935 (N_1935,N_1872,N_1821);
and U1936 (N_1936,N_1870,N_1845);
or U1937 (N_1937,N_1847,N_1803);
nand U1938 (N_1938,N_1822,N_1866);
or U1939 (N_1939,N_1818,N_1849);
or U1940 (N_1940,N_1860,N_1840);
and U1941 (N_1941,N_1809,N_1872);
or U1942 (N_1942,N_1801,N_1847);
nor U1943 (N_1943,N_1800,N_1835);
and U1944 (N_1944,N_1805,N_1828);
nand U1945 (N_1945,N_1815,N_1874);
nand U1946 (N_1946,N_1831,N_1852);
and U1947 (N_1947,N_1849,N_1832);
nor U1948 (N_1948,N_1805,N_1837);
and U1949 (N_1949,N_1820,N_1825);
or U1950 (N_1950,N_1886,N_1919);
or U1951 (N_1951,N_1883,N_1945);
and U1952 (N_1952,N_1941,N_1903);
nand U1953 (N_1953,N_1890,N_1936);
nand U1954 (N_1954,N_1915,N_1884);
or U1955 (N_1955,N_1892,N_1911);
or U1956 (N_1956,N_1897,N_1885);
or U1957 (N_1957,N_1940,N_1927);
nor U1958 (N_1958,N_1893,N_1924);
nand U1959 (N_1959,N_1902,N_1944);
or U1960 (N_1960,N_1877,N_1889);
nand U1961 (N_1961,N_1914,N_1904);
nand U1962 (N_1962,N_1882,N_1878);
nand U1963 (N_1963,N_1926,N_1896);
or U1964 (N_1964,N_1925,N_1908);
and U1965 (N_1965,N_1916,N_1929);
nor U1966 (N_1966,N_1906,N_1879);
nor U1967 (N_1967,N_1923,N_1933);
and U1968 (N_1968,N_1900,N_1947);
nand U1969 (N_1969,N_1939,N_1876);
and U1970 (N_1970,N_1918,N_1912);
nand U1971 (N_1971,N_1907,N_1921);
or U1972 (N_1972,N_1905,N_1948);
and U1973 (N_1973,N_1922,N_1917);
and U1974 (N_1974,N_1895,N_1899);
and U1975 (N_1975,N_1913,N_1938);
and U1976 (N_1976,N_1898,N_1920);
or U1977 (N_1977,N_1935,N_1949);
and U1978 (N_1978,N_1891,N_1942);
nor U1979 (N_1979,N_1932,N_1946);
and U1980 (N_1980,N_1928,N_1894);
and U1981 (N_1981,N_1888,N_1909);
nor U1982 (N_1982,N_1943,N_1880);
nor U1983 (N_1983,N_1875,N_1910);
or U1984 (N_1984,N_1881,N_1901);
or U1985 (N_1985,N_1934,N_1887);
nand U1986 (N_1986,N_1930,N_1937);
and U1987 (N_1987,N_1931,N_1875);
nor U1988 (N_1988,N_1910,N_1923);
nand U1989 (N_1989,N_1930,N_1911);
and U1990 (N_1990,N_1899,N_1903);
nand U1991 (N_1991,N_1878,N_1934);
nor U1992 (N_1992,N_1906,N_1893);
nand U1993 (N_1993,N_1919,N_1894);
nand U1994 (N_1994,N_1902,N_1896);
and U1995 (N_1995,N_1922,N_1929);
and U1996 (N_1996,N_1895,N_1936);
and U1997 (N_1997,N_1948,N_1914);
nand U1998 (N_1998,N_1916,N_1889);
and U1999 (N_1999,N_1877,N_1880);
nand U2000 (N_2000,N_1905,N_1877);
nor U2001 (N_2001,N_1900,N_1894);
and U2002 (N_2002,N_1904,N_1915);
nor U2003 (N_2003,N_1876,N_1881);
and U2004 (N_2004,N_1877,N_1930);
and U2005 (N_2005,N_1911,N_1926);
nand U2006 (N_2006,N_1930,N_1901);
nor U2007 (N_2007,N_1883,N_1910);
and U2008 (N_2008,N_1895,N_1916);
nor U2009 (N_2009,N_1888,N_1882);
nor U2010 (N_2010,N_1891,N_1933);
or U2011 (N_2011,N_1948,N_1887);
or U2012 (N_2012,N_1914,N_1930);
nor U2013 (N_2013,N_1942,N_1913);
nor U2014 (N_2014,N_1875,N_1890);
nand U2015 (N_2015,N_1914,N_1919);
or U2016 (N_2016,N_1942,N_1944);
and U2017 (N_2017,N_1902,N_1884);
or U2018 (N_2018,N_1908,N_1936);
nor U2019 (N_2019,N_1894,N_1914);
nor U2020 (N_2020,N_1898,N_1888);
nor U2021 (N_2021,N_1909,N_1887);
and U2022 (N_2022,N_1921,N_1926);
nand U2023 (N_2023,N_1897,N_1948);
or U2024 (N_2024,N_1923,N_1918);
nand U2025 (N_2025,N_2014,N_1968);
nand U2026 (N_2026,N_1977,N_1997);
nand U2027 (N_2027,N_1983,N_1986);
and U2028 (N_2028,N_1976,N_2001);
or U2029 (N_2029,N_2022,N_1993);
nor U2030 (N_2030,N_1959,N_1967);
and U2031 (N_2031,N_1951,N_2024);
and U2032 (N_2032,N_1988,N_1969);
nor U2033 (N_2033,N_1956,N_1972);
nand U2034 (N_2034,N_2008,N_1990);
or U2035 (N_2035,N_2004,N_2018);
nor U2036 (N_2036,N_2011,N_2021);
or U2037 (N_2037,N_1966,N_1974);
and U2038 (N_2038,N_1953,N_2023);
nand U2039 (N_2039,N_2009,N_1991);
or U2040 (N_2040,N_1965,N_1998);
and U2041 (N_2041,N_1955,N_1992);
or U2042 (N_2042,N_1985,N_1980);
nand U2043 (N_2043,N_1982,N_2010);
nor U2044 (N_2044,N_2006,N_1950);
nor U2045 (N_2045,N_1984,N_1958);
nor U2046 (N_2046,N_1960,N_1964);
nor U2047 (N_2047,N_1978,N_2019);
and U2048 (N_2048,N_2007,N_1954);
or U2049 (N_2049,N_1994,N_1970);
and U2050 (N_2050,N_1957,N_2005);
nor U2051 (N_2051,N_1979,N_1995);
and U2052 (N_2052,N_1963,N_2020);
nand U2053 (N_2053,N_2002,N_1952);
nor U2054 (N_2054,N_2012,N_1996);
and U2055 (N_2055,N_1961,N_1971);
or U2056 (N_2056,N_1975,N_1999);
nor U2057 (N_2057,N_2013,N_1962);
nor U2058 (N_2058,N_2017,N_2015);
nand U2059 (N_2059,N_1987,N_1973);
nor U2060 (N_2060,N_1989,N_1981);
or U2061 (N_2061,N_2003,N_2000);
nand U2062 (N_2062,N_2016,N_1975);
nand U2063 (N_2063,N_1957,N_2006);
nand U2064 (N_2064,N_1953,N_1974);
and U2065 (N_2065,N_1990,N_2015);
nor U2066 (N_2066,N_1976,N_1961);
or U2067 (N_2067,N_2017,N_2024);
nor U2068 (N_2068,N_2005,N_2020);
nand U2069 (N_2069,N_1993,N_1999);
nand U2070 (N_2070,N_1960,N_1967);
nor U2071 (N_2071,N_1981,N_2015);
or U2072 (N_2072,N_2008,N_1958);
xnor U2073 (N_2073,N_1965,N_1966);
and U2074 (N_2074,N_1954,N_2024);
nor U2075 (N_2075,N_1954,N_1965);
or U2076 (N_2076,N_2002,N_1975);
and U2077 (N_2077,N_1988,N_1987);
or U2078 (N_2078,N_2010,N_2012);
and U2079 (N_2079,N_1958,N_1999);
and U2080 (N_2080,N_1967,N_1996);
and U2081 (N_2081,N_1995,N_1998);
nor U2082 (N_2082,N_1969,N_2018);
or U2083 (N_2083,N_2014,N_1975);
and U2084 (N_2084,N_1985,N_1955);
nor U2085 (N_2085,N_1983,N_2019);
or U2086 (N_2086,N_2021,N_2003);
and U2087 (N_2087,N_1958,N_1966);
and U2088 (N_2088,N_2002,N_1973);
or U2089 (N_2089,N_2012,N_1978);
or U2090 (N_2090,N_1968,N_1989);
nand U2091 (N_2091,N_1995,N_1974);
and U2092 (N_2092,N_1987,N_2005);
nand U2093 (N_2093,N_2009,N_1970);
or U2094 (N_2094,N_2002,N_1957);
or U2095 (N_2095,N_2022,N_2007);
and U2096 (N_2096,N_1986,N_1984);
or U2097 (N_2097,N_1979,N_2023);
and U2098 (N_2098,N_1968,N_1954);
and U2099 (N_2099,N_1998,N_1984);
or U2100 (N_2100,N_2064,N_2054);
or U2101 (N_2101,N_2092,N_2031);
and U2102 (N_2102,N_2090,N_2068);
and U2103 (N_2103,N_2087,N_2027);
or U2104 (N_2104,N_2085,N_2036);
nand U2105 (N_2105,N_2080,N_2061);
and U2106 (N_2106,N_2040,N_2071);
and U2107 (N_2107,N_2091,N_2098);
nand U2108 (N_2108,N_2069,N_2079);
or U2109 (N_2109,N_2051,N_2066);
nand U2110 (N_2110,N_2094,N_2035);
nor U2111 (N_2111,N_2032,N_2057);
nor U2112 (N_2112,N_2074,N_2041);
nor U2113 (N_2113,N_2063,N_2060);
nand U2114 (N_2114,N_2025,N_2026);
nor U2115 (N_2115,N_2045,N_2034);
or U2116 (N_2116,N_2062,N_2050);
nor U2117 (N_2117,N_2077,N_2056);
nand U2118 (N_2118,N_2078,N_2048);
or U2119 (N_2119,N_2039,N_2082);
or U2120 (N_2120,N_2099,N_2049);
nor U2121 (N_2121,N_2058,N_2029);
and U2122 (N_2122,N_2088,N_2047);
nand U2123 (N_2123,N_2073,N_2038);
nand U2124 (N_2124,N_2059,N_2033);
or U2125 (N_2125,N_2096,N_2075);
and U2126 (N_2126,N_2043,N_2052);
or U2127 (N_2127,N_2053,N_2044);
or U2128 (N_2128,N_2076,N_2028);
and U2129 (N_2129,N_2081,N_2089);
nand U2130 (N_2130,N_2083,N_2093);
and U2131 (N_2131,N_2067,N_2065);
nand U2132 (N_2132,N_2046,N_2086);
nor U2133 (N_2133,N_2055,N_2037);
nand U2134 (N_2134,N_2030,N_2072);
or U2135 (N_2135,N_2095,N_2042);
and U2136 (N_2136,N_2070,N_2084);
nor U2137 (N_2137,N_2097,N_2081);
and U2138 (N_2138,N_2091,N_2032);
nor U2139 (N_2139,N_2059,N_2041);
nor U2140 (N_2140,N_2068,N_2083);
nand U2141 (N_2141,N_2055,N_2035);
nor U2142 (N_2142,N_2088,N_2053);
and U2143 (N_2143,N_2065,N_2061);
or U2144 (N_2144,N_2029,N_2052);
nand U2145 (N_2145,N_2061,N_2069);
nand U2146 (N_2146,N_2076,N_2056);
and U2147 (N_2147,N_2029,N_2046);
and U2148 (N_2148,N_2086,N_2085);
and U2149 (N_2149,N_2073,N_2056);
xnor U2150 (N_2150,N_2057,N_2028);
xnor U2151 (N_2151,N_2059,N_2058);
and U2152 (N_2152,N_2030,N_2085);
or U2153 (N_2153,N_2057,N_2029);
nor U2154 (N_2154,N_2034,N_2063);
and U2155 (N_2155,N_2061,N_2032);
or U2156 (N_2156,N_2027,N_2094);
or U2157 (N_2157,N_2047,N_2093);
and U2158 (N_2158,N_2055,N_2075);
nand U2159 (N_2159,N_2097,N_2040);
and U2160 (N_2160,N_2054,N_2047);
nor U2161 (N_2161,N_2048,N_2073);
nand U2162 (N_2162,N_2078,N_2043);
and U2163 (N_2163,N_2095,N_2090);
xor U2164 (N_2164,N_2036,N_2080);
and U2165 (N_2165,N_2068,N_2040);
or U2166 (N_2166,N_2070,N_2066);
or U2167 (N_2167,N_2088,N_2066);
nor U2168 (N_2168,N_2059,N_2077);
nor U2169 (N_2169,N_2057,N_2077);
and U2170 (N_2170,N_2030,N_2050);
nand U2171 (N_2171,N_2037,N_2064);
and U2172 (N_2172,N_2064,N_2056);
or U2173 (N_2173,N_2025,N_2088);
and U2174 (N_2174,N_2080,N_2060);
nor U2175 (N_2175,N_2165,N_2163);
nor U2176 (N_2176,N_2105,N_2162);
nor U2177 (N_2177,N_2103,N_2125);
and U2178 (N_2178,N_2155,N_2171);
nand U2179 (N_2179,N_2116,N_2158);
or U2180 (N_2180,N_2149,N_2143);
nand U2181 (N_2181,N_2140,N_2131);
nand U2182 (N_2182,N_2111,N_2102);
nand U2183 (N_2183,N_2139,N_2134);
nor U2184 (N_2184,N_2124,N_2108);
nor U2185 (N_2185,N_2122,N_2164);
and U2186 (N_2186,N_2117,N_2109);
xnor U2187 (N_2187,N_2129,N_2156);
nor U2188 (N_2188,N_2144,N_2120);
nand U2189 (N_2189,N_2148,N_2160);
nor U2190 (N_2190,N_2142,N_2150);
and U2191 (N_2191,N_2167,N_2113);
and U2192 (N_2192,N_2157,N_2174);
or U2193 (N_2193,N_2118,N_2151);
or U2194 (N_2194,N_2133,N_2110);
nor U2195 (N_2195,N_2166,N_2137);
nor U2196 (N_2196,N_2153,N_2173);
or U2197 (N_2197,N_2172,N_2115);
nor U2198 (N_2198,N_2126,N_2104);
nor U2199 (N_2199,N_2121,N_2138);
nor U2200 (N_2200,N_2170,N_2135);
or U2201 (N_2201,N_2152,N_2119);
nor U2202 (N_2202,N_2106,N_2101);
nand U2203 (N_2203,N_2112,N_2132);
nand U2204 (N_2204,N_2136,N_2107);
and U2205 (N_2205,N_2127,N_2154);
or U2206 (N_2206,N_2128,N_2161);
nor U2207 (N_2207,N_2145,N_2130);
nor U2208 (N_2208,N_2100,N_2123);
or U2209 (N_2209,N_2169,N_2159);
or U2210 (N_2210,N_2146,N_2141);
and U2211 (N_2211,N_2114,N_2168);
or U2212 (N_2212,N_2147,N_2107);
and U2213 (N_2213,N_2119,N_2174);
or U2214 (N_2214,N_2107,N_2168);
and U2215 (N_2215,N_2145,N_2174);
and U2216 (N_2216,N_2152,N_2109);
nand U2217 (N_2217,N_2169,N_2132);
nor U2218 (N_2218,N_2137,N_2134);
nand U2219 (N_2219,N_2169,N_2156);
nor U2220 (N_2220,N_2165,N_2130);
or U2221 (N_2221,N_2139,N_2142);
xnor U2222 (N_2222,N_2153,N_2140);
nor U2223 (N_2223,N_2124,N_2163);
nand U2224 (N_2224,N_2120,N_2173);
and U2225 (N_2225,N_2174,N_2111);
nand U2226 (N_2226,N_2157,N_2147);
and U2227 (N_2227,N_2171,N_2121);
nand U2228 (N_2228,N_2173,N_2143);
nand U2229 (N_2229,N_2122,N_2132);
nand U2230 (N_2230,N_2103,N_2106);
or U2231 (N_2231,N_2121,N_2152);
nand U2232 (N_2232,N_2108,N_2147);
nor U2233 (N_2233,N_2167,N_2121);
nand U2234 (N_2234,N_2125,N_2114);
nor U2235 (N_2235,N_2100,N_2169);
or U2236 (N_2236,N_2148,N_2102);
nand U2237 (N_2237,N_2155,N_2142);
nand U2238 (N_2238,N_2140,N_2116);
nor U2239 (N_2239,N_2109,N_2156);
and U2240 (N_2240,N_2103,N_2115);
or U2241 (N_2241,N_2131,N_2143);
or U2242 (N_2242,N_2168,N_2113);
nand U2243 (N_2243,N_2169,N_2120);
and U2244 (N_2244,N_2151,N_2105);
nor U2245 (N_2245,N_2107,N_2103);
or U2246 (N_2246,N_2166,N_2157);
and U2247 (N_2247,N_2144,N_2164);
or U2248 (N_2248,N_2157,N_2108);
nand U2249 (N_2249,N_2127,N_2129);
nor U2250 (N_2250,N_2179,N_2190);
and U2251 (N_2251,N_2249,N_2230);
and U2252 (N_2252,N_2237,N_2178);
and U2253 (N_2253,N_2233,N_2236);
and U2254 (N_2254,N_2188,N_2248);
and U2255 (N_2255,N_2238,N_2219);
and U2256 (N_2256,N_2184,N_2222);
nand U2257 (N_2257,N_2208,N_2185);
nand U2258 (N_2258,N_2195,N_2244);
nor U2259 (N_2259,N_2241,N_2183);
nand U2260 (N_2260,N_2239,N_2200);
or U2261 (N_2261,N_2211,N_2187);
or U2262 (N_2262,N_2216,N_2206);
and U2263 (N_2263,N_2181,N_2182);
nor U2264 (N_2264,N_2205,N_2226);
nor U2265 (N_2265,N_2207,N_2192);
or U2266 (N_2266,N_2240,N_2189);
and U2267 (N_2267,N_2217,N_2193);
nand U2268 (N_2268,N_2212,N_2180);
nor U2269 (N_2269,N_2210,N_2229);
and U2270 (N_2270,N_2214,N_2175);
nor U2271 (N_2271,N_2223,N_2231);
and U2272 (N_2272,N_2232,N_2215);
nor U2273 (N_2273,N_2201,N_2235);
and U2274 (N_2274,N_2243,N_2247);
or U2275 (N_2275,N_2242,N_2245);
nand U2276 (N_2276,N_2225,N_2176);
or U2277 (N_2277,N_2209,N_2194);
nand U2278 (N_2278,N_2227,N_2234);
nand U2279 (N_2279,N_2224,N_2191);
or U2280 (N_2280,N_2177,N_2204);
nor U2281 (N_2281,N_2203,N_2228);
and U2282 (N_2282,N_2220,N_2213);
or U2283 (N_2283,N_2246,N_2218);
nand U2284 (N_2284,N_2186,N_2197);
and U2285 (N_2285,N_2221,N_2198);
or U2286 (N_2286,N_2202,N_2199);
nand U2287 (N_2287,N_2196,N_2236);
nand U2288 (N_2288,N_2249,N_2241);
and U2289 (N_2289,N_2240,N_2196);
nor U2290 (N_2290,N_2185,N_2194);
and U2291 (N_2291,N_2182,N_2238);
and U2292 (N_2292,N_2187,N_2196);
nor U2293 (N_2293,N_2246,N_2230);
or U2294 (N_2294,N_2208,N_2193);
and U2295 (N_2295,N_2232,N_2196);
and U2296 (N_2296,N_2185,N_2191);
nor U2297 (N_2297,N_2198,N_2249);
nor U2298 (N_2298,N_2218,N_2223);
or U2299 (N_2299,N_2247,N_2200);
nand U2300 (N_2300,N_2189,N_2198);
nand U2301 (N_2301,N_2200,N_2185);
nor U2302 (N_2302,N_2217,N_2225);
nand U2303 (N_2303,N_2215,N_2224);
nand U2304 (N_2304,N_2220,N_2197);
and U2305 (N_2305,N_2229,N_2221);
or U2306 (N_2306,N_2214,N_2208);
nand U2307 (N_2307,N_2224,N_2208);
and U2308 (N_2308,N_2179,N_2181);
nor U2309 (N_2309,N_2218,N_2243);
nor U2310 (N_2310,N_2218,N_2207);
nand U2311 (N_2311,N_2213,N_2216);
or U2312 (N_2312,N_2187,N_2222);
nand U2313 (N_2313,N_2195,N_2183);
nor U2314 (N_2314,N_2180,N_2207);
or U2315 (N_2315,N_2237,N_2225);
nand U2316 (N_2316,N_2219,N_2247);
nor U2317 (N_2317,N_2228,N_2196);
nor U2318 (N_2318,N_2181,N_2189);
or U2319 (N_2319,N_2180,N_2214);
and U2320 (N_2320,N_2203,N_2181);
or U2321 (N_2321,N_2177,N_2226);
and U2322 (N_2322,N_2192,N_2228);
or U2323 (N_2323,N_2222,N_2234);
nor U2324 (N_2324,N_2224,N_2185);
nand U2325 (N_2325,N_2288,N_2318);
or U2326 (N_2326,N_2315,N_2269);
or U2327 (N_2327,N_2262,N_2293);
and U2328 (N_2328,N_2284,N_2309);
nor U2329 (N_2329,N_2319,N_2277);
nor U2330 (N_2330,N_2285,N_2290);
nand U2331 (N_2331,N_2296,N_2260);
nor U2332 (N_2332,N_2280,N_2324);
nor U2333 (N_2333,N_2321,N_2303);
and U2334 (N_2334,N_2250,N_2304);
nor U2335 (N_2335,N_2317,N_2255);
nor U2336 (N_2336,N_2271,N_2266);
and U2337 (N_2337,N_2306,N_2256);
nand U2338 (N_2338,N_2261,N_2279);
or U2339 (N_2339,N_2263,N_2265);
and U2340 (N_2340,N_2322,N_2289);
nand U2341 (N_2341,N_2308,N_2276);
nor U2342 (N_2342,N_2267,N_2272);
and U2343 (N_2343,N_2258,N_2283);
nand U2344 (N_2344,N_2302,N_2287);
and U2345 (N_2345,N_2305,N_2275);
nor U2346 (N_2346,N_2320,N_2300);
or U2347 (N_2347,N_2253,N_2316);
and U2348 (N_2348,N_2264,N_2292);
or U2349 (N_2349,N_2274,N_2286);
and U2350 (N_2350,N_2257,N_2254);
or U2351 (N_2351,N_2259,N_2268);
or U2352 (N_2352,N_2301,N_2291);
and U2353 (N_2353,N_2295,N_2313);
nor U2354 (N_2354,N_2294,N_2314);
and U2355 (N_2355,N_2273,N_2281);
nor U2356 (N_2356,N_2298,N_2282);
or U2357 (N_2357,N_2251,N_2307);
or U2358 (N_2358,N_2312,N_2270);
nand U2359 (N_2359,N_2323,N_2311);
and U2360 (N_2360,N_2278,N_2299);
nand U2361 (N_2361,N_2252,N_2297);
nand U2362 (N_2362,N_2310,N_2275);
and U2363 (N_2363,N_2302,N_2251);
and U2364 (N_2364,N_2313,N_2307);
and U2365 (N_2365,N_2313,N_2304);
and U2366 (N_2366,N_2308,N_2322);
nand U2367 (N_2367,N_2279,N_2281);
nand U2368 (N_2368,N_2251,N_2298);
nand U2369 (N_2369,N_2267,N_2251);
or U2370 (N_2370,N_2307,N_2277);
nand U2371 (N_2371,N_2318,N_2308);
nand U2372 (N_2372,N_2307,N_2309);
and U2373 (N_2373,N_2302,N_2318);
nand U2374 (N_2374,N_2307,N_2316);
or U2375 (N_2375,N_2265,N_2301);
and U2376 (N_2376,N_2264,N_2257);
nand U2377 (N_2377,N_2265,N_2269);
nor U2378 (N_2378,N_2285,N_2269);
and U2379 (N_2379,N_2253,N_2269);
or U2380 (N_2380,N_2294,N_2307);
or U2381 (N_2381,N_2286,N_2305);
nand U2382 (N_2382,N_2265,N_2271);
or U2383 (N_2383,N_2275,N_2294);
or U2384 (N_2384,N_2253,N_2277);
or U2385 (N_2385,N_2308,N_2293);
nand U2386 (N_2386,N_2297,N_2288);
and U2387 (N_2387,N_2323,N_2291);
or U2388 (N_2388,N_2268,N_2287);
and U2389 (N_2389,N_2283,N_2295);
and U2390 (N_2390,N_2322,N_2300);
and U2391 (N_2391,N_2276,N_2313);
or U2392 (N_2392,N_2250,N_2270);
nor U2393 (N_2393,N_2291,N_2285);
or U2394 (N_2394,N_2310,N_2321);
nor U2395 (N_2395,N_2297,N_2274);
and U2396 (N_2396,N_2316,N_2308);
and U2397 (N_2397,N_2301,N_2299);
nand U2398 (N_2398,N_2255,N_2308);
and U2399 (N_2399,N_2315,N_2278);
nand U2400 (N_2400,N_2375,N_2385);
nand U2401 (N_2401,N_2363,N_2372);
and U2402 (N_2402,N_2373,N_2335);
or U2403 (N_2403,N_2395,N_2355);
or U2404 (N_2404,N_2329,N_2331);
nor U2405 (N_2405,N_2338,N_2368);
or U2406 (N_2406,N_2383,N_2330);
nor U2407 (N_2407,N_2392,N_2396);
or U2408 (N_2408,N_2371,N_2387);
nor U2409 (N_2409,N_2339,N_2348);
or U2410 (N_2410,N_2378,N_2386);
nor U2411 (N_2411,N_2340,N_2353);
nor U2412 (N_2412,N_2398,N_2364);
nor U2413 (N_2413,N_2334,N_2337);
or U2414 (N_2414,N_2388,N_2345);
and U2415 (N_2415,N_2326,N_2360);
nand U2416 (N_2416,N_2389,N_2358);
nor U2417 (N_2417,N_2349,N_2343);
or U2418 (N_2418,N_2381,N_2347);
nand U2419 (N_2419,N_2367,N_2362);
or U2420 (N_2420,N_2351,N_2342);
or U2421 (N_2421,N_2379,N_2361);
nor U2422 (N_2422,N_2391,N_2341);
nor U2423 (N_2423,N_2352,N_2357);
or U2424 (N_2424,N_2397,N_2354);
or U2425 (N_2425,N_2374,N_2346);
and U2426 (N_2426,N_2332,N_2366);
nand U2427 (N_2427,N_2333,N_2370);
or U2428 (N_2428,N_2365,N_2369);
nor U2429 (N_2429,N_2336,N_2356);
or U2430 (N_2430,N_2344,N_2376);
nand U2431 (N_2431,N_2327,N_2390);
and U2432 (N_2432,N_2382,N_2328);
nand U2433 (N_2433,N_2359,N_2393);
nor U2434 (N_2434,N_2380,N_2399);
nor U2435 (N_2435,N_2350,N_2325);
and U2436 (N_2436,N_2394,N_2384);
nor U2437 (N_2437,N_2377,N_2337);
nand U2438 (N_2438,N_2378,N_2342);
nand U2439 (N_2439,N_2387,N_2334);
and U2440 (N_2440,N_2387,N_2347);
and U2441 (N_2441,N_2335,N_2359);
nand U2442 (N_2442,N_2380,N_2340);
or U2443 (N_2443,N_2399,N_2390);
and U2444 (N_2444,N_2356,N_2355);
nand U2445 (N_2445,N_2358,N_2388);
nor U2446 (N_2446,N_2377,N_2363);
nand U2447 (N_2447,N_2351,N_2343);
or U2448 (N_2448,N_2399,N_2371);
or U2449 (N_2449,N_2350,N_2339);
nand U2450 (N_2450,N_2372,N_2353);
and U2451 (N_2451,N_2333,N_2394);
nand U2452 (N_2452,N_2375,N_2371);
nand U2453 (N_2453,N_2336,N_2389);
nand U2454 (N_2454,N_2375,N_2332);
and U2455 (N_2455,N_2329,N_2387);
xor U2456 (N_2456,N_2338,N_2385);
nand U2457 (N_2457,N_2325,N_2359);
nand U2458 (N_2458,N_2347,N_2332);
or U2459 (N_2459,N_2373,N_2360);
and U2460 (N_2460,N_2332,N_2326);
and U2461 (N_2461,N_2339,N_2392);
and U2462 (N_2462,N_2385,N_2372);
nand U2463 (N_2463,N_2346,N_2399);
nand U2464 (N_2464,N_2398,N_2355);
xor U2465 (N_2465,N_2378,N_2385);
and U2466 (N_2466,N_2356,N_2341);
or U2467 (N_2467,N_2382,N_2399);
nor U2468 (N_2468,N_2330,N_2374);
or U2469 (N_2469,N_2380,N_2343);
nor U2470 (N_2470,N_2379,N_2390);
and U2471 (N_2471,N_2326,N_2376);
or U2472 (N_2472,N_2399,N_2344);
nor U2473 (N_2473,N_2364,N_2333);
nor U2474 (N_2474,N_2354,N_2335);
or U2475 (N_2475,N_2451,N_2417);
or U2476 (N_2476,N_2407,N_2432);
and U2477 (N_2477,N_2406,N_2418);
nor U2478 (N_2478,N_2463,N_2440);
or U2479 (N_2479,N_2466,N_2439);
nand U2480 (N_2480,N_2459,N_2436);
or U2481 (N_2481,N_2472,N_2410);
or U2482 (N_2482,N_2401,N_2424);
nand U2483 (N_2483,N_2444,N_2400);
nor U2484 (N_2484,N_2448,N_2468);
nor U2485 (N_2485,N_2414,N_2469);
nor U2486 (N_2486,N_2471,N_2438);
nand U2487 (N_2487,N_2458,N_2452);
nand U2488 (N_2488,N_2433,N_2456);
nor U2489 (N_2489,N_2421,N_2419);
and U2490 (N_2490,N_2420,N_2408);
nor U2491 (N_2491,N_2445,N_2470);
nand U2492 (N_2492,N_2437,N_2409);
nand U2493 (N_2493,N_2460,N_2453);
or U2494 (N_2494,N_2467,N_2404);
nor U2495 (N_2495,N_2461,N_2415);
nor U2496 (N_2496,N_2413,N_2425);
nand U2497 (N_2497,N_2427,N_2411);
or U2498 (N_2498,N_2446,N_2441);
or U2499 (N_2499,N_2454,N_2473);
nor U2500 (N_2500,N_2422,N_2430);
and U2501 (N_2501,N_2423,N_2431);
nor U2502 (N_2502,N_2402,N_2442);
and U2503 (N_2503,N_2405,N_2462);
nor U2504 (N_2504,N_2435,N_2412);
or U2505 (N_2505,N_2416,N_2447);
nor U2506 (N_2506,N_2403,N_2465);
and U2507 (N_2507,N_2443,N_2450);
and U2508 (N_2508,N_2464,N_2434);
nand U2509 (N_2509,N_2449,N_2426);
and U2510 (N_2510,N_2457,N_2474);
nand U2511 (N_2511,N_2429,N_2428);
or U2512 (N_2512,N_2455,N_2433);
nand U2513 (N_2513,N_2450,N_2470);
and U2514 (N_2514,N_2436,N_2448);
nand U2515 (N_2515,N_2415,N_2421);
nand U2516 (N_2516,N_2474,N_2464);
and U2517 (N_2517,N_2400,N_2469);
nand U2518 (N_2518,N_2438,N_2408);
nor U2519 (N_2519,N_2463,N_2406);
nand U2520 (N_2520,N_2411,N_2462);
and U2521 (N_2521,N_2413,N_2433);
nor U2522 (N_2522,N_2404,N_2412);
nand U2523 (N_2523,N_2471,N_2445);
nor U2524 (N_2524,N_2427,N_2446);
and U2525 (N_2525,N_2457,N_2473);
nor U2526 (N_2526,N_2447,N_2428);
nand U2527 (N_2527,N_2464,N_2403);
and U2528 (N_2528,N_2438,N_2435);
nor U2529 (N_2529,N_2467,N_2459);
nor U2530 (N_2530,N_2403,N_2410);
nand U2531 (N_2531,N_2411,N_2436);
nand U2532 (N_2532,N_2446,N_2420);
or U2533 (N_2533,N_2459,N_2462);
and U2534 (N_2534,N_2453,N_2437);
and U2535 (N_2535,N_2401,N_2443);
nand U2536 (N_2536,N_2443,N_2422);
nand U2537 (N_2537,N_2461,N_2427);
nor U2538 (N_2538,N_2431,N_2442);
or U2539 (N_2539,N_2425,N_2439);
or U2540 (N_2540,N_2474,N_2461);
and U2541 (N_2541,N_2459,N_2411);
nand U2542 (N_2542,N_2433,N_2409);
or U2543 (N_2543,N_2422,N_2435);
nor U2544 (N_2544,N_2423,N_2422);
and U2545 (N_2545,N_2414,N_2439);
and U2546 (N_2546,N_2448,N_2418);
and U2547 (N_2547,N_2436,N_2421);
nand U2548 (N_2548,N_2405,N_2415);
or U2549 (N_2549,N_2436,N_2451);
or U2550 (N_2550,N_2513,N_2540);
nor U2551 (N_2551,N_2477,N_2548);
or U2552 (N_2552,N_2529,N_2492);
nand U2553 (N_2553,N_2484,N_2543);
or U2554 (N_2554,N_2503,N_2545);
nor U2555 (N_2555,N_2524,N_2536);
nand U2556 (N_2556,N_2510,N_2502);
nor U2557 (N_2557,N_2495,N_2481);
and U2558 (N_2558,N_2531,N_2526);
nand U2559 (N_2559,N_2487,N_2514);
nand U2560 (N_2560,N_2506,N_2496);
nand U2561 (N_2561,N_2505,N_2507);
or U2562 (N_2562,N_2516,N_2479);
and U2563 (N_2563,N_2497,N_2493);
nor U2564 (N_2564,N_2485,N_2518);
and U2565 (N_2565,N_2541,N_2494);
nand U2566 (N_2566,N_2483,N_2509);
nand U2567 (N_2567,N_2532,N_2482);
xor U2568 (N_2568,N_2517,N_2533);
xor U2569 (N_2569,N_2547,N_2489);
nand U2570 (N_2570,N_2504,N_2476);
or U2571 (N_2571,N_2508,N_2528);
and U2572 (N_2572,N_2525,N_2521);
nand U2573 (N_2573,N_2512,N_2539);
and U2574 (N_2574,N_2491,N_2544);
and U2575 (N_2575,N_2542,N_2499);
nand U2576 (N_2576,N_2535,N_2523);
xor U2577 (N_2577,N_2488,N_2537);
or U2578 (N_2578,N_2511,N_2527);
and U2579 (N_2579,N_2546,N_2490);
or U2580 (N_2580,N_2549,N_2475);
or U2581 (N_2581,N_2486,N_2538);
and U2582 (N_2582,N_2500,N_2519);
nor U2583 (N_2583,N_2522,N_2501);
or U2584 (N_2584,N_2478,N_2534);
and U2585 (N_2585,N_2530,N_2520);
nor U2586 (N_2586,N_2498,N_2515);
nand U2587 (N_2587,N_2480,N_2492);
and U2588 (N_2588,N_2537,N_2509);
or U2589 (N_2589,N_2496,N_2517);
nor U2590 (N_2590,N_2548,N_2527);
or U2591 (N_2591,N_2479,N_2524);
nand U2592 (N_2592,N_2486,N_2537);
nand U2593 (N_2593,N_2498,N_2509);
and U2594 (N_2594,N_2507,N_2516);
or U2595 (N_2595,N_2477,N_2545);
nor U2596 (N_2596,N_2535,N_2500);
nor U2597 (N_2597,N_2482,N_2512);
nand U2598 (N_2598,N_2549,N_2500);
nor U2599 (N_2599,N_2534,N_2529);
nand U2600 (N_2600,N_2507,N_2517);
or U2601 (N_2601,N_2486,N_2490);
or U2602 (N_2602,N_2522,N_2529);
and U2603 (N_2603,N_2478,N_2483);
nand U2604 (N_2604,N_2534,N_2492);
xnor U2605 (N_2605,N_2538,N_2494);
or U2606 (N_2606,N_2540,N_2478);
or U2607 (N_2607,N_2476,N_2520);
and U2608 (N_2608,N_2549,N_2526);
and U2609 (N_2609,N_2476,N_2519);
nor U2610 (N_2610,N_2519,N_2480);
or U2611 (N_2611,N_2527,N_2517);
nor U2612 (N_2612,N_2486,N_2528);
and U2613 (N_2613,N_2476,N_2502);
and U2614 (N_2614,N_2536,N_2541);
nor U2615 (N_2615,N_2504,N_2547);
or U2616 (N_2616,N_2484,N_2513);
or U2617 (N_2617,N_2523,N_2524);
nor U2618 (N_2618,N_2492,N_2517);
and U2619 (N_2619,N_2481,N_2490);
nor U2620 (N_2620,N_2479,N_2534);
nand U2621 (N_2621,N_2494,N_2546);
nand U2622 (N_2622,N_2509,N_2543);
and U2623 (N_2623,N_2507,N_2515);
or U2624 (N_2624,N_2522,N_2531);
nand U2625 (N_2625,N_2619,N_2578);
nor U2626 (N_2626,N_2551,N_2558);
and U2627 (N_2627,N_2585,N_2616);
nand U2628 (N_2628,N_2608,N_2579);
or U2629 (N_2629,N_2573,N_2565);
nor U2630 (N_2630,N_2593,N_2600);
nand U2631 (N_2631,N_2617,N_2607);
nor U2632 (N_2632,N_2562,N_2621);
and U2633 (N_2633,N_2587,N_2580);
or U2634 (N_2634,N_2623,N_2595);
nor U2635 (N_2635,N_2564,N_2599);
nor U2636 (N_2636,N_2589,N_2605);
nor U2637 (N_2637,N_2563,N_2612);
nor U2638 (N_2638,N_2552,N_2556);
and U2639 (N_2639,N_2609,N_2604);
nor U2640 (N_2640,N_2590,N_2574);
nand U2641 (N_2641,N_2560,N_2559);
nand U2642 (N_2642,N_2568,N_2572);
nor U2643 (N_2643,N_2601,N_2586);
or U2644 (N_2644,N_2581,N_2618);
or U2645 (N_2645,N_2575,N_2570);
nand U2646 (N_2646,N_2598,N_2571);
or U2647 (N_2647,N_2583,N_2550);
or U2648 (N_2648,N_2611,N_2566);
or U2649 (N_2649,N_2594,N_2576);
or U2650 (N_2650,N_2602,N_2615);
or U2651 (N_2651,N_2584,N_2596);
or U2652 (N_2652,N_2577,N_2610);
nand U2653 (N_2653,N_2603,N_2561);
and U2654 (N_2654,N_2553,N_2614);
or U2655 (N_2655,N_2624,N_2620);
and U2656 (N_2656,N_2557,N_2554);
nand U2657 (N_2657,N_2591,N_2613);
and U2658 (N_2658,N_2582,N_2597);
or U2659 (N_2659,N_2622,N_2592);
or U2660 (N_2660,N_2555,N_2567);
and U2661 (N_2661,N_2606,N_2569);
nand U2662 (N_2662,N_2588,N_2557);
or U2663 (N_2663,N_2587,N_2553);
nor U2664 (N_2664,N_2573,N_2581);
and U2665 (N_2665,N_2577,N_2568);
nand U2666 (N_2666,N_2613,N_2610);
nand U2667 (N_2667,N_2610,N_2622);
or U2668 (N_2668,N_2571,N_2560);
or U2669 (N_2669,N_2555,N_2575);
nand U2670 (N_2670,N_2573,N_2556);
or U2671 (N_2671,N_2558,N_2550);
nand U2672 (N_2672,N_2585,N_2596);
nand U2673 (N_2673,N_2573,N_2569);
or U2674 (N_2674,N_2605,N_2606);
nand U2675 (N_2675,N_2576,N_2619);
nand U2676 (N_2676,N_2623,N_2555);
nor U2677 (N_2677,N_2555,N_2550);
nor U2678 (N_2678,N_2620,N_2558);
nor U2679 (N_2679,N_2561,N_2580);
nand U2680 (N_2680,N_2559,N_2601);
or U2681 (N_2681,N_2610,N_2604);
or U2682 (N_2682,N_2608,N_2569);
nor U2683 (N_2683,N_2593,N_2557);
nand U2684 (N_2684,N_2617,N_2558);
or U2685 (N_2685,N_2604,N_2591);
nand U2686 (N_2686,N_2589,N_2565);
and U2687 (N_2687,N_2559,N_2596);
or U2688 (N_2688,N_2602,N_2581);
nand U2689 (N_2689,N_2585,N_2611);
nand U2690 (N_2690,N_2598,N_2574);
nand U2691 (N_2691,N_2586,N_2595);
nand U2692 (N_2692,N_2601,N_2608);
nor U2693 (N_2693,N_2555,N_2573);
nand U2694 (N_2694,N_2617,N_2581);
nor U2695 (N_2695,N_2590,N_2575);
nand U2696 (N_2696,N_2565,N_2605);
nor U2697 (N_2697,N_2606,N_2568);
or U2698 (N_2698,N_2550,N_2618);
nor U2699 (N_2699,N_2557,N_2550);
and U2700 (N_2700,N_2668,N_2695);
nand U2701 (N_2701,N_2660,N_2680);
nand U2702 (N_2702,N_2666,N_2634);
and U2703 (N_2703,N_2697,N_2667);
nand U2704 (N_2704,N_2682,N_2674);
and U2705 (N_2705,N_2625,N_2681);
or U2706 (N_2706,N_2669,N_2643);
and U2707 (N_2707,N_2646,N_2665);
nor U2708 (N_2708,N_2685,N_2690);
nand U2709 (N_2709,N_2655,N_2676);
nor U2710 (N_2710,N_2640,N_2657);
and U2711 (N_2711,N_2658,N_2654);
nand U2712 (N_2712,N_2636,N_2678);
nor U2713 (N_2713,N_2670,N_2627);
nand U2714 (N_2714,N_2637,N_2663);
or U2715 (N_2715,N_2652,N_2691);
nor U2716 (N_2716,N_2653,N_2650);
nor U2717 (N_2717,N_2642,N_2687);
nand U2718 (N_2718,N_2628,N_2664);
nand U2719 (N_2719,N_2692,N_2632);
and U2720 (N_2720,N_2696,N_2659);
or U2721 (N_2721,N_2626,N_2698);
nand U2722 (N_2722,N_2662,N_2694);
nor U2723 (N_2723,N_2688,N_2638);
nand U2724 (N_2724,N_2656,N_2648);
nand U2725 (N_2725,N_2629,N_2672);
or U2726 (N_2726,N_2651,N_2644);
and U2727 (N_2727,N_2661,N_2645);
nor U2728 (N_2728,N_2633,N_2686);
or U2729 (N_2729,N_2635,N_2673);
and U2730 (N_2730,N_2630,N_2699);
or U2731 (N_2731,N_2684,N_2675);
nor U2732 (N_2732,N_2679,N_2649);
or U2733 (N_2733,N_2677,N_2671);
and U2734 (N_2734,N_2641,N_2683);
nor U2735 (N_2735,N_2689,N_2647);
or U2736 (N_2736,N_2693,N_2639);
nor U2737 (N_2737,N_2631,N_2683);
or U2738 (N_2738,N_2645,N_2695);
nor U2739 (N_2739,N_2682,N_2689);
and U2740 (N_2740,N_2695,N_2682);
nor U2741 (N_2741,N_2651,N_2695);
and U2742 (N_2742,N_2673,N_2659);
nor U2743 (N_2743,N_2656,N_2639);
nand U2744 (N_2744,N_2627,N_2695);
nand U2745 (N_2745,N_2695,N_2659);
or U2746 (N_2746,N_2654,N_2697);
nor U2747 (N_2747,N_2685,N_2634);
and U2748 (N_2748,N_2651,N_2666);
nand U2749 (N_2749,N_2697,N_2698);
or U2750 (N_2750,N_2660,N_2669);
or U2751 (N_2751,N_2639,N_2637);
nand U2752 (N_2752,N_2632,N_2675);
nor U2753 (N_2753,N_2675,N_2659);
nor U2754 (N_2754,N_2636,N_2641);
nand U2755 (N_2755,N_2661,N_2692);
nor U2756 (N_2756,N_2672,N_2692);
and U2757 (N_2757,N_2696,N_2635);
or U2758 (N_2758,N_2638,N_2689);
or U2759 (N_2759,N_2667,N_2672);
nand U2760 (N_2760,N_2693,N_2671);
nand U2761 (N_2761,N_2651,N_2628);
nor U2762 (N_2762,N_2662,N_2632);
and U2763 (N_2763,N_2645,N_2665);
and U2764 (N_2764,N_2643,N_2639);
nor U2765 (N_2765,N_2678,N_2675);
nand U2766 (N_2766,N_2629,N_2668);
nand U2767 (N_2767,N_2673,N_2680);
nand U2768 (N_2768,N_2684,N_2637);
or U2769 (N_2769,N_2692,N_2654);
nor U2770 (N_2770,N_2633,N_2690);
and U2771 (N_2771,N_2632,N_2688);
or U2772 (N_2772,N_2647,N_2677);
nor U2773 (N_2773,N_2655,N_2688);
nor U2774 (N_2774,N_2674,N_2681);
or U2775 (N_2775,N_2758,N_2749);
or U2776 (N_2776,N_2764,N_2735);
nor U2777 (N_2777,N_2713,N_2753);
nand U2778 (N_2778,N_2748,N_2719);
nor U2779 (N_2779,N_2770,N_2733);
nand U2780 (N_2780,N_2766,N_2701);
and U2781 (N_2781,N_2761,N_2714);
nor U2782 (N_2782,N_2712,N_2732);
and U2783 (N_2783,N_2741,N_2710);
nand U2784 (N_2784,N_2752,N_2718);
and U2785 (N_2785,N_2774,N_2754);
or U2786 (N_2786,N_2769,N_2702);
nand U2787 (N_2787,N_2734,N_2747);
and U2788 (N_2788,N_2728,N_2756);
or U2789 (N_2789,N_2711,N_2737);
nor U2790 (N_2790,N_2725,N_2722);
and U2791 (N_2791,N_2730,N_2731);
nor U2792 (N_2792,N_2771,N_2729);
nor U2793 (N_2793,N_2759,N_2708);
nor U2794 (N_2794,N_2727,N_2745);
and U2795 (N_2795,N_2738,N_2715);
or U2796 (N_2796,N_2768,N_2773);
nand U2797 (N_2797,N_2720,N_2716);
and U2798 (N_2798,N_2706,N_2723);
nand U2799 (N_2799,N_2709,N_2765);
nand U2800 (N_2800,N_2707,N_2744);
nor U2801 (N_2801,N_2724,N_2700);
nand U2802 (N_2802,N_2736,N_2762);
or U2803 (N_2803,N_2760,N_2740);
or U2804 (N_2804,N_2746,N_2755);
xnor U2805 (N_2805,N_2703,N_2742);
or U2806 (N_2806,N_2721,N_2717);
and U2807 (N_2807,N_2726,N_2757);
and U2808 (N_2808,N_2767,N_2743);
nand U2809 (N_2809,N_2772,N_2763);
xnor U2810 (N_2810,N_2705,N_2751);
and U2811 (N_2811,N_2750,N_2704);
or U2812 (N_2812,N_2739,N_2771);
nand U2813 (N_2813,N_2761,N_2722);
or U2814 (N_2814,N_2743,N_2766);
nor U2815 (N_2815,N_2750,N_2720);
or U2816 (N_2816,N_2736,N_2714);
nor U2817 (N_2817,N_2720,N_2724);
nor U2818 (N_2818,N_2757,N_2714);
or U2819 (N_2819,N_2702,N_2760);
xnor U2820 (N_2820,N_2739,N_2725);
nand U2821 (N_2821,N_2727,N_2728);
or U2822 (N_2822,N_2719,N_2734);
nand U2823 (N_2823,N_2700,N_2746);
or U2824 (N_2824,N_2718,N_2735);
or U2825 (N_2825,N_2742,N_2769);
or U2826 (N_2826,N_2736,N_2702);
or U2827 (N_2827,N_2727,N_2750);
nor U2828 (N_2828,N_2713,N_2738);
or U2829 (N_2829,N_2706,N_2757);
and U2830 (N_2830,N_2740,N_2766);
or U2831 (N_2831,N_2701,N_2753);
and U2832 (N_2832,N_2753,N_2710);
and U2833 (N_2833,N_2749,N_2726);
nor U2834 (N_2834,N_2728,N_2760);
and U2835 (N_2835,N_2751,N_2700);
nor U2836 (N_2836,N_2736,N_2769);
and U2837 (N_2837,N_2734,N_2772);
nor U2838 (N_2838,N_2744,N_2725);
and U2839 (N_2839,N_2713,N_2736);
and U2840 (N_2840,N_2719,N_2715);
or U2841 (N_2841,N_2739,N_2704);
or U2842 (N_2842,N_2716,N_2769);
nor U2843 (N_2843,N_2733,N_2753);
or U2844 (N_2844,N_2771,N_2769);
or U2845 (N_2845,N_2758,N_2733);
or U2846 (N_2846,N_2707,N_2756);
nor U2847 (N_2847,N_2726,N_2753);
and U2848 (N_2848,N_2763,N_2755);
nand U2849 (N_2849,N_2772,N_2745);
and U2850 (N_2850,N_2799,N_2789);
or U2851 (N_2851,N_2777,N_2781);
nand U2852 (N_2852,N_2791,N_2845);
nand U2853 (N_2853,N_2847,N_2782);
nand U2854 (N_2854,N_2838,N_2839);
and U2855 (N_2855,N_2843,N_2797);
and U2856 (N_2856,N_2842,N_2800);
and U2857 (N_2857,N_2780,N_2844);
and U2858 (N_2858,N_2819,N_2836);
and U2859 (N_2859,N_2809,N_2846);
nor U2860 (N_2860,N_2841,N_2787);
and U2861 (N_2861,N_2805,N_2822);
nand U2862 (N_2862,N_2785,N_2824);
or U2863 (N_2863,N_2828,N_2806);
xor U2864 (N_2864,N_2823,N_2775);
or U2865 (N_2865,N_2788,N_2830);
and U2866 (N_2866,N_2812,N_2811);
xnor U2867 (N_2867,N_2783,N_2820);
and U2868 (N_2868,N_2849,N_2817);
nand U2869 (N_2869,N_2829,N_2804);
nor U2870 (N_2870,N_2821,N_2796);
nor U2871 (N_2871,N_2814,N_2810);
nand U2872 (N_2872,N_2832,N_2801);
nor U2873 (N_2873,N_2833,N_2776);
nand U2874 (N_2874,N_2778,N_2786);
nor U2875 (N_2875,N_2793,N_2808);
xor U2876 (N_2876,N_2802,N_2790);
or U2877 (N_2877,N_2815,N_2798);
and U2878 (N_2878,N_2835,N_2779);
and U2879 (N_2879,N_2813,N_2831);
nand U2880 (N_2880,N_2818,N_2834);
nand U2881 (N_2881,N_2827,N_2848);
and U2882 (N_2882,N_2837,N_2792);
nor U2883 (N_2883,N_2825,N_2803);
or U2884 (N_2884,N_2795,N_2840);
and U2885 (N_2885,N_2807,N_2784);
or U2886 (N_2886,N_2794,N_2816);
or U2887 (N_2887,N_2826,N_2804);
nand U2888 (N_2888,N_2832,N_2827);
and U2889 (N_2889,N_2798,N_2778);
nand U2890 (N_2890,N_2831,N_2826);
or U2891 (N_2891,N_2835,N_2815);
or U2892 (N_2892,N_2778,N_2783);
or U2893 (N_2893,N_2808,N_2781);
nor U2894 (N_2894,N_2787,N_2783);
nor U2895 (N_2895,N_2784,N_2845);
and U2896 (N_2896,N_2805,N_2787);
and U2897 (N_2897,N_2775,N_2847);
and U2898 (N_2898,N_2818,N_2778);
nand U2899 (N_2899,N_2801,N_2819);
nor U2900 (N_2900,N_2831,N_2801);
nor U2901 (N_2901,N_2788,N_2791);
or U2902 (N_2902,N_2829,N_2777);
or U2903 (N_2903,N_2843,N_2818);
nand U2904 (N_2904,N_2827,N_2802);
nor U2905 (N_2905,N_2779,N_2787);
nor U2906 (N_2906,N_2811,N_2823);
or U2907 (N_2907,N_2840,N_2839);
nand U2908 (N_2908,N_2834,N_2825);
nor U2909 (N_2909,N_2812,N_2808);
and U2910 (N_2910,N_2820,N_2828);
nor U2911 (N_2911,N_2844,N_2797);
nor U2912 (N_2912,N_2802,N_2848);
or U2913 (N_2913,N_2786,N_2849);
or U2914 (N_2914,N_2806,N_2783);
nor U2915 (N_2915,N_2786,N_2815);
and U2916 (N_2916,N_2832,N_2830);
or U2917 (N_2917,N_2792,N_2827);
nand U2918 (N_2918,N_2840,N_2846);
or U2919 (N_2919,N_2816,N_2806);
xnor U2920 (N_2920,N_2794,N_2804);
and U2921 (N_2921,N_2834,N_2823);
nor U2922 (N_2922,N_2779,N_2810);
nand U2923 (N_2923,N_2816,N_2781);
or U2924 (N_2924,N_2785,N_2777);
and U2925 (N_2925,N_2872,N_2860);
nor U2926 (N_2926,N_2909,N_2854);
and U2927 (N_2927,N_2907,N_2919);
and U2928 (N_2928,N_2921,N_2863);
nor U2929 (N_2929,N_2920,N_2904);
and U2930 (N_2930,N_2851,N_2890);
or U2931 (N_2931,N_2876,N_2855);
nor U2932 (N_2932,N_2862,N_2866);
and U2933 (N_2933,N_2885,N_2911);
or U2934 (N_2934,N_2883,N_2880);
nand U2935 (N_2935,N_2916,N_2858);
nor U2936 (N_2936,N_2886,N_2850);
nor U2937 (N_2937,N_2870,N_2912);
and U2938 (N_2938,N_2888,N_2899);
or U2939 (N_2939,N_2887,N_2877);
or U2940 (N_2940,N_2853,N_2895);
nand U2941 (N_2941,N_2868,N_2898);
nor U2942 (N_2942,N_2859,N_2881);
nand U2943 (N_2943,N_2918,N_2871);
nand U2944 (N_2944,N_2917,N_2852);
and U2945 (N_2945,N_2900,N_2891);
nor U2946 (N_2946,N_2924,N_2865);
nand U2947 (N_2947,N_2897,N_2857);
or U2948 (N_2948,N_2856,N_2915);
nor U2949 (N_2949,N_2882,N_2910);
nand U2950 (N_2950,N_2901,N_2878);
and U2951 (N_2951,N_2873,N_2923);
nand U2952 (N_2952,N_2908,N_2893);
or U2953 (N_2953,N_2913,N_2864);
nand U2954 (N_2954,N_2861,N_2906);
nand U2955 (N_2955,N_2867,N_2892);
nor U2956 (N_2956,N_2874,N_2903);
or U2957 (N_2957,N_2914,N_2879);
nor U2958 (N_2958,N_2884,N_2922);
nor U2959 (N_2959,N_2905,N_2896);
or U2960 (N_2960,N_2875,N_2902);
nand U2961 (N_2961,N_2894,N_2869);
and U2962 (N_2962,N_2889,N_2884);
and U2963 (N_2963,N_2922,N_2887);
and U2964 (N_2964,N_2907,N_2864);
or U2965 (N_2965,N_2851,N_2904);
nor U2966 (N_2966,N_2876,N_2901);
nor U2967 (N_2967,N_2912,N_2882);
or U2968 (N_2968,N_2912,N_2888);
nor U2969 (N_2969,N_2890,N_2886);
nand U2970 (N_2970,N_2872,N_2891);
nor U2971 (N_2971,N_2851,N_2874);
or U2972 (N_2972,N_2850,N_2882);
or U2973 (N_2973,N_2863,N_2882);
nor U2974 (N_2974,N_2900,N_2922);
and U2975 (N_2975,N_2921,N_2911);
nand U2976 (N_2976,N_2868,N_2897);
and U2977 (N_2977,N_2867,N_2873);
nor U2978 (N_2978,N_2898,N_2852);
nor U2979 (N_2979,N_2883,N_2858);
and U2980 (N_2980,N_2882,N_2885);
and U2981 (N_2981,N_2893,N_2903);
nor U2982 (N_2982,N_2864,N_2911);
xor U2983 (N_2983,N_2924,N_2852);
nand U2984 (N_2984,N_2863,N_2903);
and U2985 (N_2985,N_2883,N_2857);
nor U2986 (N_2986,N_2921,N_2876);
nor U2987 (N_2987,N_2923,N_2892);
nand U2988 (N_2988,N_2872,N_2868);
or U2989 (N_2989,N_2892,N_2857);
nand U2990 (N_2990,N_2883,N_2861);
and U2991 (N_2991,N_2859,N_2889);
and U2992 (N_2992,N_2924,N_2886);
xor U2993 (N_2993,N_2877,N_2867);
or U2994 (N_2994,N_2852,N_2921);
nor U2995 (N_2995,N_2905,N_2914);
nand U2996 (N_2996,N_2866,N_2857);
or U2997 (N_2997,N_2881,N_2874);
or U2998 (N_2998,N_2880,N_2918);
nand U2999 (N_2999,N_2922,N_2892);
or UO_0 (O_0,N_2973,N_2976);
nor UO_1 (O_1,N_2982,N_2943);
nor UO_2 (O_2,N_2977,N_2999);
nand UO_3 (O_3,N_2980,N_2989);
and UO_4 (O_4,N_2926,N_2964);
nand UO_5 (O_5,N_2928,N_2930);
or UO_6 (O_6,N_2998,N_2933);
and UO_7 (O_7,N_2953,N_2979);
and UO_8 (O_8,N_2972,N_2994);
nor UO_9 (O_9,N_2981,N_2946);
or UO_10 (O_10,N_2934,N_2968);
nand UO_11 (O_11,N_2945,N_2931);
nand UO_12 (O_12,N_2988,N_2938);
nor UO_13 (O_13,N_2960,N_2978);
nor UO_14 (O_14,N_2942,N_2944);
nand UO_15 (O_15,N_2986,N_2975);
or UO_16 (O_16,N_2995,N_2990);
nand UO_17 (O_17,N_2935,N_2993);
nor UO_18 (O_18,N_2961,N_2932);
nand UO_19 (O_19,N_2937,N_2957);
xnor UO_20 (O_20,N_2984,N_2970);
and UO_21 (O_21,N_2940,N_2992);
and UO_22 (O_22,N_2963,N_2971);
nand UO_23 (O_23,N_2983,N_2997);
or UO_24 (O_24,N_2991,N_2947);
nand UO_25 (O_25,N_2985,N_2951);
nor UO_26 (O_26,N_2996,N_2958);
and UO_27 (O_27,N_2954,N_2962);
or UO_28 (O_28,N_2967,N_2929);
and UO_29 (O_29,N_2966,N_2955);
or UO_30 (O_30,N_2927,N_2974);
and UO_31 (O_31,N_2941,N_2952);
nand UO_32 (O_32,N_2925,N_2949);
and UO_33 (O_33,N_2959,N_2987);
nand UO_34 (O_34,N_2969,N_2965);
nand UO_35 (O_35,N_2950,N_2936);
or UO_36 (O_36,N_2956,N_2948);
nand UO_37 (O_37,N_2939,N_2992);
or UO_38 (O_38,N_2944,N_2945);
or UO_39 (O_39,N_2992,N_2933);
or UO_40 (O_40,N_2958,N_2991);
and UO_41 (O_41,N_2939,N_2965);
nand UO_42 (O_42,N_2971,N_2947);
nand UO_43 (O_43,N_2963,N_2968);
and UO_44 (O_44,N_2984,N_2991);
and UO_45 (O_45,N_2975,N_2944);
and UO_46 (O_46,N_2950,N_2978);
nor UO_47 (O_47,N_2979,N_2942);
nor UO_48 (O_48,N_2925,N_2957);
xor UO_49 (O_49,N_2976,N_2965);
nor UO_50 (O_50,N_2954,N_2990);
and UO_51 (O_51,N_2969,N_2993);
and UO_52 (O_52,N_2929,N_2927);
or UO_53 (O_53,N_2938,N_2987);
and UO_54 (O_54,N_2963,N_2980);
nor UO_55 (O_55,N_2993,N_2980);
or UO_56 (O_56,N_2971,N_2982);
or UO_57 (O_57,N_2984,N_2948);
and UO_58 (O_58,N_2930,N_2963);
or UO_59 (O_59,N_2986,N_2941);
and UO_60 (O_60,N_2944,N_2984);
nor UO_61 (O_61,N_2963,N_2975);
and UO_62 (O_62,N_2975,N_2925);
nor UO_63 (O_63,N_2947,N_2976);
or UO_64 (O_64,N_2968,N_2975);
nor UO_65 (O_65,N_2966,N_2927);
xnor UO_66 (O_66,N_2931,N_2983);
or UO_67 (O_67,N_2950,N_2984);
and UO_68 (O_68,N_2956,N_2985);
and UO_69 (O_69,N_2969,N_2992);
nor UO_70 (O_70,N_2952,N_2999);
and UO_71 (O_71,N_2986,N_2971);
nand UO_72 (O_72,N_2976,N_2945);
nand UO_73 (O_73,N_2971,N_2925);
nor UO_74 (O_74,N_2940,N_2979);
nor UO_75 (O_75,N_2981,N_2998);
and UO_76 (O_76,N_2950,N_2925);
and UO_77 (O_77,N_2927,N_2942);
nand UO_78 (O_78,N_2986,N_2943);
and UO_79 (O_79,N_2951,N_2989);
nor UO_80 (O_80,N_2937,N_2941);
or UO_81 (O_81,N_2999,N_2936);
or UO_82 (O_82,N_2945,N_2996);
nor UO_83 (O_83,N_2929,N_2935);
xor UO_84 (O_84,N_2934,N_2963);
or UO_85 (O_85,N_2926,N_2976);
nor UO_86 (O_86,N_2951,N_2963);
nor UO_87 (O_87,N_2956,N_2935);
xor UO_88 (O_88,N_2958,N_2973);
nor UO_89 (O_89,N_2928,N_2948);
or UO_90 (O_90,N_2973,N_2943);
nand UO_91 (O_91,N_2981,N_2925);
nand UO_92 (O_92,N_2928,N_2962);
nand UO_93 (O_93,N_2925,N_2948);
and UO_94 (O_94,N_2949,N_2963);
or UO_95 (O_95,N_2942,N_2954);
nand UO_96 (O_96,N_2931,N_2960);
and UO_97 (O_97,N_2976,N_2970);
nor UO_98 (O_98,N_2992,N_2991);
nand UO_99 (O_99,N_2977,N_2935);
or UO_100 (O_100,N_2976,N_2937);
nor UO_101 (O_101,N_2930,N_2960);
or UO_102 (O_102,N_2982,N_2944);
nand UO_103 (O_103,N_2955,N_2940);
nor UO_104 (O_104,N_2955,N_2954);
and UO_105 (O_105,N_2958,N_2940);
and UO_106 (O_106,N_2951,N_2990);
and UO_107 (O_107,N_2944,N_2928);
and UO_108 (O_108,N_2927,N_2938);
and UO_109 (O_109,N_2992,N_2966);
nor UO_110 (O_110,N_2931,N_2981);
nand UO_111 (O_111,N_2982,N_2992);
nand UO_112 (O_112,N_2926,N_2995);
or UO_113 (O_113,N_2956,N_2969);
nand UO_114 (O_114,N_2989,N_2969);
nor UO_115 (O_115,N_2929,N_2943);
nor UO_116 (O_116,N_2965,N_2954);
nand UO_117 (O_117,N_2965,N_2949);
or UO_118 (O_118,N_2936,N_2947);
nand UO_119 (O_119,N_2963,N_2973);
or UO_120 (O_120,N_2953,N_2958);
and UO_121 (O_121,N_2975,N_2993);
and UO_122 (O_122,N_2981,N_2960);
nand UO_123 (O_123,N_2928,N_2987);
and UO_124 (O_124,N_2941,N_2995);
and UO_125 (O_125,N_2947,N_2984);
and UO_126 (O_126,N_2948,N_2932);
nor UO_127 (O_127,N_2961,N_2934);
or UO_128 (O_128,N_2928,N_2999);
nor UO_129 (O_129,N_2984,N_2971);
or UO_130 (O_130,N_2939,N_2972);
and UO_131 (O_131,N_2982,N_2994);
nor UO_132 (O_132,N_2948,N_2988);
and UO_133 (O_133,N_2951,N_2925);
or UO_134 (O_134,N_2996,N_2935);
and UO_135 (O_135,N_2936,N_2963);
nor UO_136 (O_136,N_2960,N_2945);
nand UO_137 (O_137,N_2957,N_2993);
nand UO_138 (O_138,N_2945,N_2952);
and UO_139 (O_139,N_2928,N_2925);
nor UO_140 (O_140,N_2997,N_2960);
or UO_141 (O_141,N_2931,N_2975);
or UO_142 (O_142,N_2932,N_2974);
and UO_143 (O_143,N_2937,N_2999);
nor UO_144 (O_144,N_2927,N_2932);
nand UO_145 (O_145,N_2953,N_2945);
nand UO_146 (O_146,N_2945,N_2946);
nand UO_147 (O_147,N_2939,N_2925);
or UO_148 (O_148,N_2991,N_2986);
and UO_149 (O_149,N_2946,N_2971);
nor UO_150 (O_150,N_2953,N_2997);
and UO_151 (O_151,N_2996,N_2973);
nand UO_152 (O_152,N_2967,N_2926);
nor UO_153 (O_153,N_2978,N_2957);
nor UO_154 (O_154,N_2929,N_2930);
nor UO_155 (O_155,N_2985,N_2941);
and UO_156 (O_156,N_2992,N_2964);
nor UO_157 (O_157,N_2980,N_2929);
and UO_158 (O_158,N_2987,N_2949);
nand UO_159 (O_159,N_2987,N_2948);
or UO_160 (O_160,N_2971,N_2936);
nand UO_161 (O_161,N_2994,N_2934);
nand UO_162 (O_162,N_2971,N_2977);
and UO_163 (O_163,N_2934,N_2943);
nand UO_164 (O_164,N_2980,N_2965);
or UO_165 (O_165,N_2949,N_2955);
nand UO_166 (O_166,N_2960,N_2987);
nand UO_167 (O_167,N_2934,N_2997);
and UO_168 (O_168,N_2985,N_2961);
and UO_169 (O_169,N_2927,N_2954);
or UO_170 (O_170,N_2948,N_2976);
or UO_171 (O_171,N_2950,N_2981);
nor UO_172 (O_172,N_2955,N_2973);
nor UO_173 (O_173,N_2970,N_2977);
and UO_174 (O_174,N_2956,N_2931);
nand UO_175 (O_175,N_2943,N_2968);
nand UO_176 (O_176,N_2958,N_2976);
and UO_177 (O_177,N_2988,N_2978);
nor UO_178 (O_178,N_2965,N_2955);
xnor UO_179 (O_179,N_2976,N_2990);
nand UO_180 (O_180,N_2949,N_2977);
and UO_181 (O_181,N_2962,N_2972);
and UO_182 (O_182,N_2999,N_2997);
nor UO_183 (O_183,N_2928,N_2974);
nand UO_184 (O_184,N_2926,N_2993);
or UO_185 (O_185,N_2928,N_2984);
and UO_186 (O_186,N_2965,N_2958);
or UO_187 (O_187,N_2948,N_2944);
nor UO_188 (O_188,N_2960,N_2975);
nor UO_189 (O_189,N_2928,N_2966);
or UO_190 (O_190,N_2949,N_2992);
nor UO_191 (O_191,N_2990,N_2966);
nor UO_192 (O_192,N_2994,N_2954);
nor UO_193 (O_193,N_2973,N_2928);
and UO_194 (O_194,N_2997,N_2954);
or UO_195 (O_195,N_2958,N_2931);
or UO_196 (O_196,N_2936,N_2980);
or UO_197 (O_197,N_2987,N_2995);
xnor UO_198 (O_198,N_2957,N_2934);
nor UO_199 (O_199,N_2996,N_2964);
or UO_200 (O_200,N_2948,N_2982);
and UO_201 (O_201,N_2973,N_2977);
and UO_202 (O_202,N_2975,N_2936);
and UO_203 (O_203,N_2964,N_2999);
nand UO_204 (O_204,N_2927,N_2953);
nor UO_205 (O_205,N_2935,N_2967);
nand UO_206 (O_206,N_2996,N_2959);
and UO_207 (O_207,N_2937,N_2950);
and UO_208 (O_208,N_2978,N_2972);
or UO_209 (O_209,N_2976,N_2998);
nand UO_210 (O_210,N_2990,N_2950);
or UO_211 (O_211,N_2987,N_2976);
nor UO_212 (O_212,N_2967,N_2941);
and UO_213 (O_213,N_2961,N_2981);
nor UO_214 (O_214,N_2950,N_2953);
nor UO_215 (O_215,N_2965,N_2935);
and UO_216 (O_216,N_2962,N_2946);
nand UO_217 (O_217,N_2963,N_2974);
nand UO_218 (O_218,N_2990,N_2989);
nand UO_219 (O_219,N_2954,N_2993);
and UO_220 (O_220,N_2950,N_2964);
and UO_221 (O_221,N_2931,N_2952);
nor UO_222 (O_222,N_2963,N_2982);
nor UO_223 (O_223,N_2940,N_2941);
and UO_224 (O_224,N_2952,N_2927);
nor UO_225 (O_225,N_2989,N_2943);
nand UO_226 (O_226,N_2977,N_2939);
nor UO_227 (O_227,N_2988,N_2983);
or UO_228 (O_228,N_2974,N_2945);
nand UO_229 (O_229,N_2997,N_2985);
and UO_230 (O_230,N_2967,N_2934);
nor UO_231 (O_231,N_2940,N_2948);
or UO_232 (O_232,N_2999,N_2985);
nand UO_233 (O_233,N_2930,N_2992);
and UO_234 (O_234,N_2974,N_2997);
nand UO_235 (O_235,N_2945,N_2933);
or UO_236 (O_236,N_2967,N_2943);
nor UO_237 (O_237,N_2987,N_2997);
nand UO_238 (O_238,N_2982,N_2986);
nand UO_239 (O_239,N_2996,N_2954);
nand UO_240 (O_240,N_2980,N_2948);
nor UO_241 (O_241,N_2964,N_2930);
or UO_242 (O_242,N_2935,N_2926);
nand UO_243 (O_243,N_2993,N_2932);
nor UO_244 (O_244,N_2996,N_2927);
or UO_245 (O_245,N_2964,N_2928);
or UO_246 (O_246,N_2950,N_2965);
nand UO_247 (O_247,N_2983,N_2952);
nand UO_248 (O_248,N_2925,N_2970);
nand UO_249 (O_249,N_2978,N_2984);
and UO_250 (O_250,N_2946,N_2970);
and UO_251 (O_251,N_2928,N_2954);
nand UO_252 (O_252,N_2966,N_2947);
and UO_253 (O_253,N_2973,N_2934);
nand UO_254 (O_254,N_2970,N_2926);
and UO_255 (O_255,N_2930,N_2941);
or UO_256 (O_256,N_2936,N_2976);
nor UO_257 (O_257,N_2936,N_2937);
nor UO_258 (O_258,N_2948,N_2963);
nand UO_259 (O_259,N_2936,N_2995);
nand UO_260 (O_260,N_2991,N_2961);
xnor UO_261 (O_261,N_2954,N_2941);
and UO_262 (O_262,N_2937,N_2986);
or UO_263 (O_263,N_2961,N_2931);
and UO_264 (O_264,N_2939,N_2987);
nor UO_265 (O_265,N_2993,N_2972);
and UO_266 (O_266,N_2932,N_2981);
or UO_267 (O_267,N_2931,N_2947);
and UO_268 (O_268,N_2997,N_2939);
nand UO_269 (O_269,N_2964,N_2981);
nor UO_270 (O_270,N_2945,N_2994);
and UO_271 (O_271,N_2982,N_2952);
or UO_272 (O_272,N_2993,N_2962);
nor UO_273 (O_273,N_2994,N_2974);
and UO_274 (O_274,N_2992,N_2980);
and UO_275 (O_275,N_2940,N_2986);
or UO_276 (O_276,N_2956,N_2939);
or UO_277 (O_277,N_2925,N_2977);
and UO_278 (O_278,N_2937,N_2935);
nor UO_279 (O_279,N_2994,N_2955);
and UO_280 (O_280,N_2948,N_2986);
and UO_281 (O_281,N_2931,N_2943);
or UO_282 (O_282,N_2949,N_2968);
nor UO_283 (O_283,N_2962,N_2938);
and UO_284 (O_284,N_2968,N_2933);
or UO_285 (O_285,N_2996,N_2948);
and UO_286 (O_286,N_2928,N_2957);
and UO_287 (O_287,N_2995,N_2986);
or UO_288 (O_288,N_2968,N_2996);
and UO_289 (O_289,N_2968,N_2928);
and UO_290 (O_290,N_2989,N_2971);
or UO_291 (O_291,N_2970,N_2968);
or UO_292 (O_292,N_2950,N_2989);
and UO_293 (O_293,N_2932,N_2956);
nor UO_294 (O_294,N_2976,N_2959);
or UO_295 (O_295,N_2927,N_2965);
nand UO_296 (O_296,N_2971,N_2991);
nand UO_297 (O_297,N_2968,N_2936);
or UO_298 (O_298,N_2975,N_2979);
nor UO_299 (O_299,N_2934,N_2956);
nor UO_300 (O_300,N_2926,N_2929);
or UO_301 (O_301,N_2990,N_2934);
nor UO_302 (O_302,N_2960,N_2926);
or UO_303 (O_303,N_2999,N_2953);
nor UO_304 (O_304,N_2971,N_2987);
or UO_305 (O_305,N_2967,N_2996);
nand UO_306 (O_306,N_2967,N_2972);
and UO_307 (O_307,N_2926,N_2941);
or UO_308 (O_308,N_2929,N_2944);
nor UO_309 (O_309,N_2953,N_2955);
or UO_310 (O_310,N_2976,N_2928);
and UO_311 (O_311,N_2943,N_2974);
nand UO_312 (O_312,N_2994,N_2995);
nor UO_313 (O_313,N_2945,N_2997);
nand UO_314 (O_314,N_2977,N_2933);
nor UO_315 (O_315,N_2964,N_2937);
nor UO_316 (O_316,N_2987,N_2990);
or UO_317 (O_317,N_2957,N_2941);
nor UO_318 (O_318,N_2975,N_2991);
nor UO_319 (O_319,N_2999,N_2965);
or UO_320 (O_320,N_2966,N_2942);
nand UO_321 (O_321,N_2985,N_2970);
nand UO_322 (O_322,N_2951,N_2971);
and UO_323 (O_323,N_2956,N_2984);
nor UO_324 (O_324,N_2954,N_2972);
nor UO_325 (O_325,N_2950,N_2985);
or UO_326 (O_326,N_2946,N_2956);
nand UO_327 (O_327,N_2987,N_2983);
nand UO_328 (O_328,N_2948,N_2992);
nand UO_329 (O_329,N_2983,N_2951);
nand UO_330 (O_330,N_2957,N_2979);
nor UO_331 (O_331,N_2938,N_2943);
nor UO_332 (O_332,N_2926,N_2966);
or UO_333 (O_333,N_2949,N_2966);
nor UO_334 (O_334,N_2957,N_2964);
nor UO_335 (O_335,N_2996,N_2941);
nand UO_336 (O_336,N_2948,N_2926);
or UO_337 (O_337,N_2984,N_2939);
nor UO_338 (O_338,N_2994,N_2973);
or UO_339 (O_339,N_2943,N_2925);
or UO_340 (O_340,N_2977,N_2958);
and UO_341 (O_341,N_2933,N_2972);
nand UO_342 (O_342,N_2992,N_2932);
nand UO_343 (O_343,N_2933,N_2983);
nor UO_344 (O_344,N_2981,N_2984);
or UO_345 (O_345,N_2965,N_2996);
nor UO_346 (O_346,N_2975,N_2985);
and UO_347 (O_347,N_2964,N_2929);
nor UO_348 (O_348,N_2933,N_2938);
and UO_349 (O_349,N_2932,N_2930);
and UO_350 (O_350,N_2962,N_2990);
nand UO_351 (O_351,N_2934,N_2995);
nor UO_352 (O_352,N_2988,N_2968);
or UO_353 (O_353,N_2964,N_2931);
or UO_354 (O_354,N_2930,N_2994);
nor UO_355 (O_355,N_2980,N_2927);
nor UO_356 (O_356,N_2961,N_2959);
nand UO_357 (O_357,N_2932,N_2933);
or UO_358 (O_358,N_2974,N_2929);
nand UO_359 (O_359,N_2979,N_2956);
nand UO_360 (O_360,N_2950,N_2973);
and UO_361 (O_361,N_2941,N_2955);
and UO_362 (O_362,N_2936,N_2988);
or UO_363 (O_363,N_2957,N_2963);
nand UO_364 (O_364,N_2969,N_2952);
and UO_365 (O_365,N_2997,N_2996);
and UO_366 (O_366,N_2972,N_2970);
and UO_367 (O_367,N_2946,N_2987);
and UO_368 (O_368,N_2936,N_2970);
nand UO_369 (O_369,N_2961,N_2949);
or UO_370 (O_370,N_2975,N_2939);
or UO_371 (O_371,N_2957,N_2951);
nor UO_372 (O_372,N_2932,N_2971);
nor UO_373 (O_373,N_2972,N_2979);
nor UO_374 (O_374,N_2928,N_2980);
and UO_375 (O_375,N_2964,N_2993);
nor UO_376 (O_376,N_2985,N_2982);
nor UO_377 (O_377,N_2938,N_2966);
nand UO_378 (O_378,N_2990,N_2980);
nor UO_379 (O_379,N_2980,N_2935);
nand UO_380 (O_380,N_2936,N_2974);
nor UO_381 (O_381,N_2930,N_2993);
or UO_382 (O_382,N_2929,N_2956);
and UO_383 (O_383,N_2985,N_2934);
nor UO_384 (O_384,N_2984,N_2968);
nor UO_385 (O_385,N_2932,N_2991);
or UO_386 (O_386,N_2979,N_2961);
and UO_387 (O_387,N_2950,N_2983);
nor UO_388 (O_388,N_2978,N_2929);
nor UO_389 (O_389,N_2988,N_2970);
nor UO_390 (O_390,N_2997,N_2937);
and UO_391 (O_391,N_2995,N_2930);
xor UO_392 (O_392,N_2987,N_2957);
nor UO_393 (O_393,N_2968,N_2927);
and UO_394 (O_394,N_2944,N_2978);
and UO_395 (O_395,N_2945,N_2947);
nor UO_396 (O_396,N_2979,N_2936);
nor UO_397 (O_397,N_2958,N_2961);
nor UO_398 (O_398,N_2959,N_2934);
and UO_399 (O_399,N_2937,N_2963);
or UO_400 (O_400,N_2930,N_2979);
nand UO_401 (O_401,N_2925,N_2953);
and UO_402 (O_402,N_2956,N_2959);
and UO_403 (O_403,N_2974,N_2982);
and UO_404 (O_404,N_2990,N_2933);
nor UO_405 (O_405,N_2953,N_2957);
nand UO_406 (O_406,N_2996,N_2966);
or UO_407 (O_407,N_2972,N_2997);
nand UO_408 (O_408,N_2944,N_2964);
nand UO_409 (O_409,N_2939,N_2991);
and UO_410 (O_410,N_2929,N_2985);
and UO_411 (O_411,N_2938,N_2940);
xnor UO_412 (O_412,N_2994,N_2950);
and UO_413 (O_413,N_2998,N_2966);
nor UO_414 (O_414,N_2930,N_2954);
or UO_415 (O_415,N_2925,N_2927);
nor UO_416 (O_416,N_2946,N_2926);
nor UO_417 (O_417,N_2930,N_2949);
or UO_418 (O_418,N_2942,N_2996);
and UO_419 (O_419,N_2949,N_2985);
and UO_420 (O_420,N_2933,N_2981);
or UO_421 (O_421,N_2983,N_2967);
nor UO_422 (O_422,N_2968,N_2954);
nor UO_423 (O_423,N_2970,N_2932);
nand UO_424 (O_424,N_2972,N_2926);
nor UO_425 (O_425,N_2962,N_2932);
or UO_426 (O_426,N_2935,N_2987);
and UO_427 (O_427,N_2931,N_2969);
nor UO_428 (O_428,N_2983,N_2937);
or UO_429 (O_429,N_2942,N_2974);
nor UO_430 (O_430,N_2945,N_2990);
nand UO_431 (O_431,N_2983,N_2998);
or UO_432 (O_432,N_2948,N_2971);
nor UO_433 (O_433,N_2972,N_2928);
nor UO_434 (O_434,N_2932,N_2986);
nor UO_435 (O_435,N_2959,N_2969);
nand UO_436 (O_436,N_2979,N_2996);
nor UO_437 (O_437,N_2944,N_2991);
nor UO_438 (O_438,N_2979,N_2964);
and UO_439 (O_439,N_2988,N_2994);
or UO_440 (O_440,N_2978,N_2975);
or UO_441 (O_441,N_2997,N_2958);
and UO_442 (O_442,N_2963,N_2994);
and UO_443 (O_443,N_2965,N_2979);
nand UO_444 (O_444,N_2999,N_2995);
and UO_445 (O_445,N_2957,N_2948);
and UO_446 (O_446,N_2956,N_2933);
or UO_447 (O_447,N_2978,N_2947);
or UO_448 (O_448,N_2979,N_2932);
and UO_449 (O_449,N_2999,N_2932);
nand UO_450 (O_450,N_2951,N_2977);
nand UO_451 (O_451,N_2931,N_2977);
or UO_452 (O_452,N_2976,N_2981);
nand UO_453 (O_453,N_2943,N_2951);
nand UO_454 (O_454,N_2973,N_2992);
or UO_455 (O_455,N_2991,N_2968);
and UO_456 (O_456,N_2979,N_2962);
and UO_457 (O_457,N_2926,N_2950);
and UO_458 (O_458,N_2959,N_2950);
nor UO_459 (O_459,N_2973,N_2941);
nand UO_460 (O_460,N_2932,N_2998);
nand UO_461 (O_461,N_2997,N_2952);
nor UO_462 (O_462,N_2988,N_2950);
nand UO_463 (O_463,N_2970,N_2993);
nand UO_464 (O_464,N_2976,N_2964);
xor UO_465 (O_465,N_2956,N_2994);
or UO_466 (O_466,N_2988,N_2944);
xor UO_467 (O_467,N_2931,N_2996);
or UO_468 (O_468,N_2995,N_2957);
nand UO_469 (O_469,N_2969,N_2967);
or UO_470 (O_470,N_2992,N_2975);
and UO_471 (O_471,N_2930,N_2968);
nand UO_472 (O_472,N_2925,N_2959);
and UO_473 (O_473,N_2941,N_2945);
or UO_474 (O_474,N_2983,N_2962);
or UO_475 (O_475,N_2939,N_2994);
nor UO_476 (O_476,N_2954,N_2989);
nand UO_477 (O_477,N_2962,N_2953);
nor UO_478 (O_478,N_2957,N_2962);
or UO_479 (O_479,N_2958,N_2959);
nand UO_480 (O_480,N_2935,N_2963);
and UO_481 (O_481,N_2998,N_2988);
and UO_482 (O_482,N_2972,N_2929);
nand UO_483 (O_483,N_2986,N_2930);
and UO_484 (O_484,N_2929,N_2928);
or UO_485 (O_485,N_2932,N_2984);
nand UO_486 (O_486,N_2953,N_2972);
nor UO_487 (O_487,N_2957,N_2933);
and UO_488 (O_488,N_2982,N_2954);
or UO_489 (O_489,N_2952,N_2951);
nor UO_490 (O_490,N_2955,N_2958);
or UO_491 (O_491,N_2946,N_2938);
and UO_492 (O_492,N_2996,N_2998);
nand UO_493 (O_493,N_2930,N_2944);
and UO_494 (O_494,N_2992,N_2944);
nor UO_495 (O_495,N_2927,N_2973);
nand UO_496 (O_496,N_2983,N_2947);
nand UO_497 (O_497,N_2986,N_2993);
nor UO_498 (O_498,N_2968,N_2955);
and UO_499 (O_499,N_2925,N_2962);
endmodule