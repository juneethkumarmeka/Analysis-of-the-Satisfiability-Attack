module basic_500_3000_500_5_levels_1xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_375,In_420);
nor U1 (N_1,In_171,In_157);
and U2 (N_2,In_142,In_319);
nor U3 (N_3,In_5,In_206);
nor U4 (N_4,In_355,In_159);
and U5 (N_5,In_62,In_86);
nand U6 (N_6,In_230,In_228);
nand U7 (N_7,In_468,In_361);
or U8 (N_8,In_457,In_426);
nand U9 (N_9,In_97,In_282);
and U10 (N_10,In_397,In_11);
or U11 (N_11,In_132,In_41);
or U12 (N_12,In_493,In_446);
nand U13 (N_13,In_209,In_290);
or U14 (N_14,In_150,In_182);
nor U15 (N_15,In_491,In_227);
and U16 (N_16,In_357,In_197);
nand U17 (N_17,In_279,In_35);
and U18 (N_18,In_73,In_237);
nand U19 (N_19,In_429,In_168);
and U20 (N_20,In_211,In_494);
nor U21 (N_21,In_193,In_336);
or U22 (N_22,In_274,In_323);
nand U23 (N_23,In_466,In_87);
or U24 (N_24,In_471,In_320);
nor U25 (N_25,In_344,In_31);
and U26 (N_26,In_307,In_124);
nand U27 (N_27,In_376,In_149);
and U28 (N_28,In_378,In_358);
nor U29 (N_29,In_176,In_184);
nor U30 (N_30,In_219,In_160);
nor U31 (N_31,In_127,In_377);
nand U32 (N_32,In_49,In_218);
and U33 (N_33,In_202,In_349);
nand U34 (N_34,In_164,In_108);
and U35 (N_35,In_96,In_327);
or U36 (N_36,In_386,In_194);
nor U37 (N_37,In_295,In_45);
or U38 (N_38,In_431,In_204);
nand U39 (N_39,In_186,In_247);
nor U40 (N_40,In_101,In_205);
nor U41 (N_41,In_146,In_153);
and U42 (N_42,In_210,In_367);
nor U43 (N_43,In_165,In_396);
nand U44 (N_44,In_94,In_67);
or U45 (N_45,In_434,In_325);
or U46 (N_46,In_14,In_221);
nand U47 (N_47,In_53,In_419);
or U48 (N_48,In_269,In_328);
or U49 (N_49,In_423,In_347);
nand U50 (N_50,In_388,In_170);
nand U51 (N_51,In_499,In_65);
nor U52 (N_52,In_185,In_178);
and U53 (N_53,In_331,In_403);
nand U54 (N_54,In_453,In_270);
nand U55 (N_55,In_283,In_58);
and U56 (N_56,In_253,In_255);
nor U57 (N_57,In_389,In_278);
nor U58 (N_58,In_63,In_179);
nor U59 (N_59,In_425,In_314);
or U60 (N_60,In_46,In_445);
nor U61 (N_61,In_217,In_112);
or U62 (N_62,In_43,In_66);
and U63 (N_63,In_360,In_381);
nor U64 (N_64,In_29,In_435);
and U65 (N_65,In_267,In_414);
nand U66 (N_66,In_24,In_48);
and U67 (N_67,In_92,In_301);
and U68 (N_68,In_313,In_248);
nor U69 (N_69,In_346,In_464);
nand U70 (N_70,In_384,In_369);
nand U71 (N_71,In_289,In_229);
or U72 (N_72,In_47,In_405);
and U73 (N_73,In_291,In_447);
or U74 (N_74,In_42,In_226);
or U75 (N_75,In_415,In_359);
nor U76 (N_76,In_3,In_98);
nor U77 (N_77,In_44,In_37);
or U78 (N_78,In_286,In_133);
or U79 (N_79,In_469,In_104);
and U80 (N_80,In_141,In_497);
and U81 (N_81,In_490,In_382);
nand U82 (N_82,In_456,In_27);
nand U83 (N_83,In_222,In_401);
nand U84 (N_84,In_161,In_277);
nand U85 (N_85,In_77,In_348);
and U86 (N_86,In_474,In_352);
and U87 (N_87,In_343,In_433);
or U88 (N_88,In_341,In_231);
and U89 (N_89,In_135,In_76);
nand U90 (N_90,In_380,In_488);
nor U91 (N_91,In_191,In_241);
nand U92 (N_92,In_353,In_345);
and U93 (N_93,In_110,In_311);
nand U94 (N_94,In_310,In_308);
and U95 (N_95,In_467,In_64);
and U96 (N_96,In_485,In_363);
nor U97 (N_97,In_462,In_100);
nand U98 (N_98,In_402,In_252);
xor U99 (N_99,In_69,In_472);
and U100 (N_100,In_299,In_16);
nand U101 (N_101,In_298,In_81);
and U102 (N_102,In_59,In_15);
nor U103 (N_103,In_71,In_495);
or U104 (N_104,In_317,In_262);
or U105 (N_105,In_326,In_392);
and U106 (N_106,In_4,In_215);
or U107 (N_107,In_188,In_276);
or U108 (N_108,In_232,In_409);
xnor U109 (N_109,In_154,In_373);
nor U110 (N_110,In_196,In_366);
and U111 (N_111,In_421,In_492);
nor U112 (N_112,In_408,In_128);
nand U113 (N_113,In_280,In_8);
and U114 (N_114,In_356,In_121);
nand U115 (N_115,In_138,In_334);
nand U116 (N_116,In_13,In_103);
and U117 (N_117,In_312,In_254);
nor U118 (N_118,In_246,In_6);
and U119 (N_119,In_195,In_236);
or U120 (N_120,In_477,In_12);
nor U121 (N_121,In_166,In_427);
and U122 (N_122,In_249,In_234);
xor U123 (N_123,In_83,In_105);
and U124 (N_124,In_258,In_264);
nor U125 (N_125,In_123,In_39);
nor U126 (N_126,In_259,In_296);
or U127 (N_127,In_23,In_18);
nor U128 (N_128,In_385,In_281);
nand U129 (N_129,In_309,In_461);
nor U130 (N_130,In_126,In_163);
or U131 (N_131,In_52,In_338);
or U132 (N_132,In_424,In_368);
and U133 (N_133,In_330,In_131);
nand U134 (N_134,In_441,In_432);
and U135 (N_135,In_25,In_362);
or U136 (N_136,In_339,In_20);
nand U137 (N_137,In_198,In_407);
or U138 (N_138,In_463,In_240);
nand U139 (N_139,In_272,In_379);
or U140 (N_140,In_129,In_275);
nand U141 (N_141,In_238,In_201);
and U142 (N_142,In_90,In_213);
nor U143 (N_143,In_475,In_111);
nand U144 (N_144,In_273,In_383);
xnor U145 (N_145,In_140,In_89);
and U146 (N_146,In_413,In_174);
and U147 (N_147,In_487,In_235);
or U148 (N_148,In_93,In_0);
and U149 (N_149,In_478,In_75);
nor U150 (N_150,In_95,In_333);
nor U151 (N_151,In_51,In_340);
nor U152 (N_152,In_102,In_114);
or U153 (N_153,In_483,In_61);
nand U154 (N_154,In_411,In_189);
and U155 (N_155,In_137,In_329);
nand U156 (N_156,In_1,In_162);
or U157 (N_157,In_297,In_106);
or U158 (N_158,In_79,In_448);
nor U159 (N_159,In_26,In_122);
nor U160 (N_160,In_91,In_422);
nand U161 (N_161,In_167,In_315);
or U162 (N_162,In_294,In_38);
or U163 (N_163,In_451,In_199);
nand U164 (N_164,In_117,In_34);
or U165 (N_165,In_9,In_173);
or U166 (N_166,In_155,In_410);
nor U167 (N_167,In_465,In_350);
and U168 (N_168,In_30,In_486);
or U169 (N_169,In_261,In_233);
or U170 (N_170,In_216,In_481);
nand U171 (N_171,In_21,In_36);
nor U172 (N_172,In_460,In_351);
and U173 (N_173,In_130,In_212);
or U174 (N_174,In_187,In_342);
nor U175 (N_175,In_439,In_444);
nor U176 (N_176,In_285,In_119);
and U177 (N_177,In_84,In_250);
and U178 (N_178,In_391,In_374);
nand U179 (N_179,In_256,In_223);
nor U180 (N_180,In_145,In_387);
and U181 (N_181,In_74,In_482);
nand U182 (N_182,In_136,In_85);
nand U183 (N_183,In_109,In_316);
nand U184 (N_184,In_293,In_395);
or U185 (N_185,In_496,In_55);
nand U186 (N_186,In_57,In_239);
nor U187 (N_187,In_364,In_152);
and U188 (N_188,In_354,In_337);
or U189 (N_189,In_470,In_225);
nor U190 (N_190,In_263,In_372);
or U191 (N_191,In_390,In_332);
and U192 (N_192,In_2,In_175);
and U193 (N_193,In_72,In_300);
nand U194 (N_194,In_17,In_207);
xor U195 (N_195,In_268,In_371);
and U196 (N_196,In_134,In_214);
nor U197 (N_197,In_302,In_416);
nor U198 (N_198,In_60,In_139);
and U199 (N_199,In_208,In_116);
or U200 (N_200,In_7,In_406);
or U201 (N_201,In_107,In_394);
and U202 (N_202,In_455,In_220);
and U203 (N_203,In_148,In_260);
and U204 (N_204,In_177,In_143);
and U205 (N_205,In_480,In_144);
and U206 (N_206,In_284,In_292);
nand U207 (N_207,In_266,In_365);
or U208 (N_208,In_430,In_113);
nand U209 (N_209,In_56,In_476);
and U210 (N_210,In_479,In_442);
and U211 (N_211,In_172,In_489);
and U212 (N_212,In_404,In_440);
nor U213 (N_213,In_70,In_203);
and U214 (N_214,In_125,In_370);
and U215 (N_215,In_183,In_473);
nand U216 (N_216,In_245,In_417);
and U217 (N_217,In_54,In_78);
or U218 (N_218,In_484,In_412);
and U219 (N_219,In_303,In_288);
or U220 (N_220,In_318,In_443);
nor U221 (N_221,In_190,In_257);
nand U222 (N_222,In_393,In_19);
or U223 (N_223,In_305,In_99);
nor U224 (N_224,In_271,In_82);
and U225 (N_225,In_287,In_321);
and U226 (N_226,In_28,In_398);
and U227 (N_227,In_243,In_147);
and U228 (N_228,In_68,In_242);
nor U229 (N_229,In_498,In_251);
nand U230 (N_230,In_88,In_22);
nor U231 (N_231,In_458,In_400);
nand U232 (N_232,In_169,In_459);
or U233 (N_233,In_80,In_306);
and U234 (N_234,In_438,In_437);
nand U235 (N_235,In_151,In_50);
nor U236 (N_236,In_10,In_33);
or U237 (N_237,In_156,In_265);
and U238 (N_238,In_120,In_428);
or U239 (N_239,In_118,In_324);
or U240 (N_240,In_192,In_436);
nand U241 (N_241,In_224,In_335);
nand U242 (N_242,In_115,In_304);
and U243 (N_243,In_450,In_244);
nand U244 (N_244,In_454,In_452);
nor U245 (N_245,In_32,In_449);
nand U246 (N_246,In_200,In_158);
and U247 (N_247,In_399,In_180);
and U248 (N_248,In_418,In_322);
nor U249 (N_249,In_181,In_40);
nand U250 (N_250,In_401,In_32);
and U251 (N_251,In_203,In_167);
nand U252 (N_252,In_220,In_215);
nand U253 (N_253,In_401,In_301);
nor U254 (N_254,In_89,In_300);
or U255 (N_255,In_46,In_252);
and U256 (N_256,In_497,In_475);
and U257 (N_257,In_98,In_188);
or U258 (N_258,In_95,In_303);
nor U259 (N_259,In_442,In_269);
or U260 (N_260,In_115,In_491);
nor U261 (N_261,In_316,In_423);
nor U262 (N_262,In_349,In_168);
and U263 (N_263,In_199,In_446);
nand U264 (N_264,In_30,In_109);
and U265 (N_265,In_254,In_13);
and U266 (N_266,In_486,In_264);
or U267 (N_267,In_462,In_31);
nand U268 (N_268,In_42,In_218);
nor U269 (N_269,In_101,In_337);
and U270 (N_270,In_176,In_365);
or U271 (N_271,In_141,In_177);
xnor U272 (N_272,In_62,In_172);
and U273 (N_273,In_203,In_357);
or U274 (N_274,In_412,In_471);
or U275 (N_275,In_48,In_364);
nand U276 (N_276,In_4,In_327);
nand U277 (N_277,In_107,In_100);
and U278 (N_278,In_364,In_0);
and U279 (N_279,In_481,In_96);
nor U280 (N_280,In_451,In_267);
or U281 (N_281,In_430,In_334);
or U282 (N_282,In_382,In_478);
or U283 (N_283,In_194,In_442);
nor U284 (N_284,In_239,In_232);
nand U285 (N_285,In_45,In_137);
nand U286 (N_286,In_192,In_61);
or U287 (N_287,In_319,In_155);
or U288 (N_288,In_172,In_101);
nor U289 (N_289,In_50,In_45);
nand U290 (N_290,In_397,In_364);
or U291 (N_291,In_132,In_6);
nor U292 (N_292,In_296,In_484);
and U293 (N_293,In_135,In_139);
nand U294 (N_294,In_353,In_288);
nor U295 (N_295,In_466,In_153);
nor U296 (N_296,In_183,In_52);
or U297 (N_297,In_451,In_205);
and U298 (N_298,In_477,In_460);
or U299 (N_299,In_445,In_146);
nor U300 (N_300,In_462,In_211);
nor U301 (N_301,In_142,In_257);
nand U302 (N_302,In_395,In_472);
nor U303 (N_303,In_239,In_496);
and U304 (N_304,In_257,In_0);
nor U305 (N_305,In_477,In_231);
or U306 (N_306,In_33,In_205);
or U307 (N_307,In_134,In_311);
or U308 (N_308,In_187,In_193);
nor U309 (N_309,In_476,In_59);
or U310 (N_310,In_381,In_296);
nor U311 (N_311,In_203,In_143);
or U312 (N_312,In_162,In_32);
or U313 (N_313,In_75,In_315);
and U314 (N_314,In_283,In_170);
nor U315 (N_315,In_5,In_106);
nor U316 (N_316,In_368,In_402);
and U317 (N_317,In_13,In_24);
or U318 (N_318,In_291,In_303);
or U319 (N_319,In_268,In_161);
nand U320 (N_320,In_329,In_262);
and U321 (N_321,In_456,In_44);
and U322 (N_322,In_333,In_283);
or U323 (N_323,In_177,In_65);
nor U324 (N_324,In_85,In_322);
nand U325 (N_325,In_330,In_465);
nand U326 (N_326,In_206,In_109);
nor U327 (N_327,In_420,In_153);
nor U328 (N_328,In_361,In_222);
nor U329 (N_329,In_116,In_300);
nand U330 (N_330,In_443,In_460);
or U331 (N_331,In_365,In_77);
nor U332 (N_332,In_178,In_3);
nor U333 (N_333,In_335,In_274);
or U334 (N_334,In_171,In_16);
or U335 (N_335,In_241,In_290);
or U336 (N_336,In_365,In_339);
and U337 (N_337,In_127,In_239);
nand U338 (N_338,In_300,In_125);
and U339 (N_339,In_258,In_471);
nand U340 (N_340,In_170,In_158);
nand U341 (N_341,In_48,In_346);
or U342 (N_342,In_398,In_157);
nor U343 (N_343,In_157,In_230);
nor U344 (N_344,In_465,In_294);
and U345 (N_345,In_164,In_434);
or U346 (N_346,In_448,In_158);
and U347 (N_347,In_472,In_57);
or U348 (N_348,In_386,In_458);
nand U349 (N_349,In_195,In_175);
and U350 (N_350,In_193,In_298);
or U351 (N_351,In_140,In_47);
or U352 (N_352,In_233,In_405);
nor U353 (N_353,In_86,In_214);
and U354 (N_354,In_157,In_85);
nand U355 (N_355,In_98,In_221);
nor U356 (N_356,In_133,In_220);
and U357 (N_357,In_442,In_1);
nor U358 (N_358,In_482,In_157);
nand U359 (N_359,In_322,In_215);
nand U360 (N_360,In_497,In_364);
and U361 (N_361,In_279,In_8);
nand U362 (N_362,In_354,In_436);
nand U363 (N_363,In_420,In_277);
nor U364 (N_364,In_415,In_165);
nor U365 (N_365,In_424,In_413);
or U366 (N_366,In_40,In_321);
or U367 (N_367,In_460,In_57);
or U368 (N_368,In_498,In_467);
nand U369 (N_369,In_69,In_325);
nand U370 (N_370,In_118,In_354);
nand U371 (N_371,In_229,In_255);
nand U372 (N_372,In_274,In_217);
nand U373 (N_373,In_360,In_479);
and U374 (N_374,In_489,In_275);
nand U375 (N_375,In_317,In_388);
and U376 (N_376,In_435,In_337);
nand U377 (N_377,In_215,In_353);
nand U378 (N_378,In_184,In_362);
xor U379 (N_379,In_375,In_86);
or U380 (N_380,In_386,In_360);
and U381 (N_381,In_475,In_45);
nand U382 (N_382,In_392,In_76);
nor U383 (N_383,In_176,In_108);
and U384 (N_384,In_177,In_448);
or U385 (N_385,In_242,In_12);
nor U386 (N_386,In_289,In_78);
and U387 (N_387,In_240,In_182);
nand U388 (N_388,In_393,In_234);
and U389 (N_389,In_397,In_79);
nand U390 (N_390,In_204,In_250);
and U391 (N_391,In_191,In_6);
nor U392 (N_392,In_68,In_71);
or U393 (N_393,In_355,In_184);
or U394 (N_394,In_253,In_466);
nor U395 (N_395,In_244,In_409);
and U396 (N_396,In_215,In_42);
and U397 (N_397,In_203,In_417);
and U398 (N_398,In_246,In_304);
nor U399 (N_399,In_91,In_84);
and U400 (N_400,In_295,In_64);
or U401 (N_401,In_233,In_332);
or U402 (N_402,In_305,In_215);
nor U403 (N_403,In_431,In_393);
or U404 (N_404,In_334,In_344);
nor U405 (N_405,In_441,In_268);
nand U406 (N_406,In_290,In_159);
and U407 (N_407,In_452,In_216);
nor U408 (N_408,In_65,In_92);
nand U409 (N_409,In_213,In_216);
and U410 (N_410,In_472,In_81);
and U411 (N_411,In_224,In_52);
nand U412 (N_412,In_158,In_452);
nor U413 (N_413,In_189,In_32);
nor U414 (N_414,In_312,In_390);
and U415 (N_415,In_296,In_433);
or U416 (N_416,In_120,In_485);
and U417 (N_417,In_25,In_256);
nor U418 (N_418,In_29,In_96);
and U419 (N_419,In_290,In_119);
nor U420 (N_420,In_78,In_480);
and U421 (N_421,In_50,In_302);
nand U422 (N_422,In_444,In_3);
nand U423 (N_423,In_36,In_260);
nor U424 (N_424,In_267,In_310);
nand U425 (N_425,In_281,In_74);
nand U426 (N_426,In_22,In_248);
and U427 (N_427,In_97,In_65);
and U428 (N_428,In_204,In_261);
and U429 (N_429,In_115,In_371);
nor U430 (N_430,In_346,In_215);
nand U431 (N_431,In_241,In_460);
or U432 (N_432,In_315,In_404);
or U433 (N_433,In_356,In_409);
or U434 (N_434,In_222,In_212);
nor U435 (N_435,In_54,In_52);
and U436 (N_436,In_410,In_143);
nor U437 (N_437,In_344,In_447);
nand U438 (N_438,In_437,In_159);
or U439 (N_439,In_100,In_19);
nor U440 (N_440,In_258,In_475);
and U441 (N_441,In_127,In_120);
nand U442 (N_442,In_111,In_444);
nor U443 (N_443,In_280,In_91);
or U444 (N_444,In_433,In_325);
and U445 (N_445,In_179,In_110);
or U446 (N_446,In_451,In_417);
or U447 (N_447,In_399,In_135);
nor U448 (N_448,In_191,In_313);
nor U449 (N_449,In_393,In_139);
and U450 (N_450,In_103,In_139);
and U451 (N_451,In_213,In_269);
or U452 (N_452,In_456,In_145);
and U453 (N_453,In_61,In_281);
nor U454 (N_454,In_303,In_267);
nand U455 (N_455,In_239,In_314);
nor U456 (N_456,In_267,In_387);
and U457 (N_457,In_447,In_269);
nand U458 (N_458,In_33,In_104);
and U459 (N_459,In_69,In_414);
nor U460 (N_460,In_86,In_41);
nand U461 (N_461,In_229,In_364);
nand U462 (N_462,In_159,In_288);
or U463 (N_463,In_64,In_493);
nand U464 (N_464,In_112,In_462);
and U465 (N_465,In_95,In_368);
or U466 (N_466,In_443,In_283);
and U467 (N_467,In_251,In_162);
nor U468 (N_468,In_52,In_371);
nand U469 (N_469,In_468,In_20);
nor U470 (N_470,In_196,In_7);
nor U471 (N_471,In_304,In_336);
and U472 (N_472,In_231,In_58);
and U473 (N_473,In_155,In_27);
xor U474 (N_474,In_13,In_166);
or U475 (N_475,In_5,In_32);
or U476 (N_476,In_377,In_351);
nand U477 (N_477,In_396,In_212);
nor U478 (N_478,In_316,In_493);
or U479 (N_479,In_348,In_105);
nor U480 (N_480,In_362,In_48);
nor U481 (N_481,In_220,In_285);
and U482 (N_482,In_104,In_417);
nor U483 (N_483,In_354,In_479);
or U484 (N_484,In_125,In_407);
nand U485 (N_485,In_138,In_9);
nor U486 (N_486,In_385,In_341);
nor U487 (N_487,In_314,In_269);
nor U488 (N_488,In_384,In_101);
nor U489 (N_489,In_270,In_460);
nand U490 (N_490,In_305,In_131);
and U491 (N_491,In_134,In_356);
or U492 (N_492,In_493,In_20);
nor U493 (N_493,In_92,In_331);
nand U494 (N_494,In_362,In_176);
and U495 (N_495,In_402,In_164);
or U496 (N_496,In_151,In_441);
nand U497 (N_497,In_156,In_137);
nor U498 (N_498,In_455,In_145);
and U499 (N_499,In_272,In_406);
and U500 (N_500,In_352,In_158);
or U501 (N_501,In_141,In_205);
or U502 (N_502,In_149,In_122);
nand U503 (N_503,In_403,In_443);
and U504 (N_504,In_198,In_20);
nor U505 (N_505,In_229,In_138);
nor U506 (N_506,In_51,In_174);
nand U507 (N_507,In_498,In_439);
and U508 (N_508,In_347,In_475);
or U509 (N_509,In_0,In_401);
or U510 (N_510,In_355,In_95);
nor U511 (N_511,In_204,In_164);
nand U512 (N_512,In_414,In_165);
nor U513 (N_513,In_169,In_411);
nor U514 (N_514,In_300,In_360);
nor U515 (N_515,In_199,In_407);
or U516 (N_516,In_323,In_309);
or U517 (N_517,In_475,In_333);
nand U518 (N_518,In_383,In_385);
and U519 (N_519,In_281,In_108);
and U520 (N_520,In_334,In_84);
nor U521 (N_521,In_50,In_346);
nor U522 (N_522,In_249,In_364);
and U523 (N_523,In_290,In_491);
nor U524 (N_524,In_332,In_295);
and U525 (N_525,In_442,In_391);
nand U526 (N_526,In_232,In_68);
nand U527 (N_527,In_66,In_98);
or U528 (N_528,In_223,In_283);
and U529 (N_529,In_253,In_432);
and U530 (N_530,In_255,In_366);
nor U531 (N_531,In_235,In_408);
or U532 (N_532,In_473,In_467);
nand U533 (N_533,In_231,In_422);
or U534 (N_534,In_434,In_165);
and U535 (N_535,In_358,In_80);
or U536 (N_536,In_104,In_31);
or U537 (N_537,In_158,In_172);
nand U538 (N_538,In_144,In_199);
xnor U539 (N_539,In_19,In_66);
nor U540 (N_540,In_300,In_491);
nor U541 (N_541,In_453,In_259);
nor U542 (N_542,In_370,In_452);
and U543 (N_543,In_413,In_442);
nand U544 (N_544,In_168,In_222);
and U545 (N_545,In_316,In_302);
and U546 (N_546,In_474,In_398);
and U547 (N_547,In_149,In_330);
nor U548 (N_548,In_76,In_295);
nor U549 (N_549,In_305,In_413);
or U550 (N_550,In_326,In_144);
or U551 (N_551,In_346,In_399);
nor U552 (N_552,In_177,In_1);
or U553 (N_553,In_341,In_428);
nand U554 (N_554,In_281,In_439);
nor U555 (N_555,In_178,In_344);
nand U556 (N_556,In_82,In_220);
nor U557 (N_557,In_447,In_411);
or U558 (N_558,In_399,In_361);
or U559 (N_559,In_201,In_20);
nand U560 (N_560,In_76,In_486);
or U561 (N_561,In_289,In_82);
nand U562 (N_562,In_403,In_258);
nand U563 (N_563,In_345,In_331);
and U564 (N_564,In_359,In_465);
and U565 (N_565,In_122,In_312);
xnor U566 (N_566,In_67,In_119);
nor U567 (N_567,In_436,In_209);
nor U568 (N_568,In_256,In_261);
nor U569 (N_569,In_161,In_246);
or U570 (N_570,In_201,In_121);
nand U571 (N_571,In_109,In_468);
nand U572 (N_572,In_400,In_424);
nand U573 (N_573,In_225,In_477);
and U574 (N_574,In_306,In_142);
nand U575 (N_575,In_68,In_170);
xnor U576 (N_576,In_131,In_286);
nand U577 (N_577,In_298,In_459);
or U578 (N_578,In_143,In_197);
nand U579 (N_579,In_471,In_326);
or U580 (N_580,In_64,In_355);
nand U581 (N_581,In_315,In_431);
nand U582 (N_582,In_336,In_92);
or U583 (N_583,In_343,In_14);
or U584 (N_584,In_12,In_312);
nor U585 (N_585,In_108,In_438);
nand U586 (N_586,In_2,In_12);
and U587 (N_587,In_229,In_133);
and U588 (N_588,In_263,In_21);
and U589 (N_589,In_491,In_221);
and U590 (N_590,In_313,In_268);
nor U591 (N_591,In_223,In_207);
or U592 (N_592,In_477,In_154);
and U593 (N_593,In_354,In_313);
and U594 (N_594,In_39,In_470);
nor U595 (N_595,In_438,In_379);
nand U596 (N_596,In_122,In_116);
or U597 (N_597,In_43,In_0);
and U598 (N_598,In_341,In_469);
nand U599 (N_599,In_131,In_316);
and U600 (N_600,N_318,N_227);
or U601 (N_601,N_384,N_412);
or U602 (N_602,N_365,N_552);
and U603 (N_603,N_126,N_25);
or U604 (N_604,N_89,N_91);
nand U605 (N_605,N_498,N_307);
nand U606 (N_606,N_296,N_24);
and U607 (N_607,N_175,N_110);
and U608 (N_608,N_234,N_94);
and U609 (N_609,N_397,N_53);
nand U610 (N_610,N_285,N_288);
nor U611 (N_611,N_414,N_97);
nand U612 (N_612,N_541,N_270);
nand U613 (N_613,N_119,N_28);
nor U614 (N_614,N_494,N_261);
or U615 (N_615,N_579,N_586);
nor U616 (N_616,N_484,N_395);
or U617 (N_617,N_294,N_396);
or U618 (N_618,N_135,N_338);
nand U619 (N_619,N_56,N_420);
nand U620 (N_620,N_247,N_316);
and U621 (N_621,N_473,N_352);
nand U622 (N_622,N_4,N_324);
nand U623 (N_623,N_60,N_444);
nor U624 (N_624,N_581,N_5);
and U625 (N_625,N_140,N_597);
nand U626 (N_626,N_272,N_82);
nor U627 (N_627,N_8,N_78);
or U628 (N_628,N_287,N_172);
nand U629 (N_629,N_81,N_15);
nand U630 (N_630,N_171,N_204);
or U631 (N_631,N_495,N_464);
nand U632 (N_632,N_73,N_353);
and U633 (N_633,N_465,N_402);
and U634 (N_634,N_167,N_523);
nor U635 (N_635,N_563,N_404);
nor U636 (N_636,N_400,N_540);
nor U637 (N_637,N_301,N_569);
nor U638 (N_638,N_197,N_374);
or U639 (N_639,N_79,N_302);
nor U640 (N_640,N_339,N_36);
nor U641 (N_641,N_105,N_405);
or U642 (N_642,N_159,N_551);
nand U643 (N_643,N_263,N_330);
and U644 (N_644,N_107,N_511);
xnor U645 (N_645,N_170,N_253);
and U646 (N_646,N_526,N_411);
or U647 (N_647,N_276,N_350);
nor U648 (N_648,N_446,N_92);
and U649 (N_649,N_65,N_554);
nor U650 (N_650,N_249,N_327);
nor U651 (N_651,N_516,N_162);
and U652 (N_652,N_359,N_435);
or U653 (N_653,N_96,N_328);
and U654 (N_654,N_485,N_478);
nor U655 (N_655,N_363,N_326);
nor U656 (N_656,N_510,N_504);
and U657 (N_657,N_205,N_262);
and U658 (N_658,N_35,N_341);
nand U659 (N_659,N_113,N_593);
and U660 (N_660,N_539,N_144);
and U661 (N_661,N_174,N_546);
or U662 (N_662,N_450,N_3);
and U663 (N_663,N_203,N_386);
and U664 (N_664,N_37,N_588);
or U665 (N_665,N_553,N_34);
nand U666 (N_666,N_325,N_310);
nor U667 (N_667,N_189,N_467);
or U668 (N_668,N_9,N_461);
nand U669 (N_669,N_472,N_27);
nor U670 (N_670,N_116,N_256);
nand U671 (N_671,N_442,N_124);
and U672 (N_672,N_88,N_535);
nor U673 (N_673,N_257,N_19);
or U674 (N_674,N_576,N_429);
or U675 (N_675,N_466,N_422);
nor U676 (N_676,N_136,N_533);
nor U677 (N_677,N_245,N_419);
or U678 (N_678,N_337,N_240);
nor U679 (N_679,N_59,N_375);
or U680 (N_680,N_232,N_154);
or U681 (N_681,N_222,N_399);
nand U682 (N_682,N_90,N_560);
nor U683 (N_683,N_229,N_164);
and U684 (N_684,N_574,N_371);
or U685 (N_685,N_50,N_572);
nor U686 (N_686,N_438,N_474);
nor U687 (N_687,N_483,N_317);
and U688 (N_688,N_499,N_190);
nor U689 (N_689,N_457,N_543);
nor U690 (N_690,N_566,N_520);
nand U691 (N_691,N_85,N_304);
nor U692 (N_692,N_214,N_7);
nand U693 (N_693,N_347,N_517);
or U694 (N_694,N_66,N_482);
nand U695 (N_695,N_244,N_246);
and U696 (N_696,N_226,N_127);
nand U697 (N_697,N_69,N_598);
or U698 (N_698,N_455,N_106);
nor U699 (N_699,N_391,N_254);
nor U700 (N_700,N_387,N_198);
nand U701 (N_701,N_131,N_344);
or U702 (N_702,N_236,N_80);
or U703 (N_703,N_208,N_538);
or U704 (N_704,N_441,N_114);
or U705 (N_705,N_202,N_258);
and U706 (N_706,N_133,N_280);
and U707 (N_707,N_292,N_480);
nand U708 (N_708,N_440,N_383);
nor U709 (N_709,N_549,N_217);
or U710 (N_710,N_173,N_282);
nand U711 (N_711,N_231,N_152);
nand U712 (N_712,N_587,N_77);
nand U713 (N_713,N_537,N_143);
nand U714 (N_714,N_416,N_401);
nor U715 (N_715,N_295,N_306);
or U716 (N_716,N_515,N_380);
xnor U717 (N_717,N_93,N_122);
nand U718 (N_718,N_260,N_489);
nand U719 (N_719,N_346,N_463);
or U720 (N_720,N_309,N_18);
nand U721 (N_721,N_477,N_321);
nand U722 (N_722,N_1,N_577);
nand U723 (N_723,N_595,N_468);
and U724 (N_724,N_233,N_486);
or U725 (N_725,N_241,N_536);
and U726 (N_726,N_142,N_385);
nand U727 (N_727,N_487,N_454);
nand U728 (N_728,N_445,N_108);
or U729 (N_729,N_392,N_443);
or U730 (N_730,N_458,N_248);
nor U731 (N_731,N_319,N_447);
xnor U732 (N_732,N_426,N_599);
nand U733 (N_733,N_590,N_503);
or U734 (N_734,N_51,N_218);
nand U735 (N_735,N_207,N_75);
nand U736 (N_736,N_67,N_462);
nor U737 (N_737,N_111,N_573);
nand U738 (N_738,N_571,N_531);
or U739 (N_739,N_421,N_264);
nand U740 (N_740,N_284,N_428);
nor U741 (N_741,N_354,N_83);
or U742 (N_742,N_112,N_196);
or U743 (N_743,N_14,N_373);
nor U744 (N_744,N_524,N_74);
nor U745 (N_745,N_239,N_379);
nor U746 (N_746,N_409,N_289);
or U747 (N_747,N_475,N_86);
and U748 (N_748,N_559,N_448);
and U749 (N_749,N_48,N_283);
or U750 (N_750,N_519,N_84);
or U751 (N_751,N_439,N_160);
nand U752 (N_752,N_95,N_130);
xnor U753 (N_753,N_456,N_49);
nand U754 (N_754,N_575,N_192);
or U755 (N_755,N_161,N_123);
or U756 (N_756,N_431,N_490);
and U757 (N_757,N_23,N_179);
nand U758 (N_758,N_413,N_230);
or U759 (N_759,N_155,N_206);
nor U760 (N_760,N_11,N_407);
nand U761 (N_761,N_237,N_532);
nand U762 (N_762,N_87,N_64);
nand U763 (N_763,N_471,N_449);
nand U764 (N_764,N_265,N_147);
nand U765 (N_765,N_313,N_393);
nor U766 (N_766,N_46,N_382);
and U767 (N_767,N_44,N_225);
or U768 (N_768,N_219,N_479);
and U769 (N_769,N_589,N_290);
nand U770 (N_770,N_323,N_216);
and U771 (N_771,N_340,N_32);
or U772 (N_772,N_279,N_33);
and U773 (N_773,N_369,N_388);
nand U774 (N_774,N_72,N_334);
nor U775 (N_775,N_26,N_176);
and U776 (N_776,N_180,N_286);
and U777 (N_777,N_492,N_356);
and U778 (N_778,N_355,N_527);
nand U779 (N_779,N_224,N_120);
or U780 (N_780,N_199,N_98);
and U781 (N_781,N_298,N_544);
or U782 (N_782,N_335,N_582);
nand U783 (N_783,N_22,N_255);
nand U784 (N_784,N_149,N_488);
or U785 (N_785,N_238,N_432);
and U786 (N_786,N_186,N_496);
or U787 (N_787,N_41,N_491);
nor U788 (N_788,N_243,N_303);
nand U789 (N_789,N_31,N_138);
nand U790 (N_790,N_157,N_406);
nor U791 (N_791,N_70,N_137);
nor U792 (N_792,N_134,N_367);
or U793 (N_793,N_320,N_182);
nand U794 (N_794,N_315,N_220);
and U795 (N_795,N_361,N_194);
or U796 (N_796,N_470,N_377);
nand U797 (N_797,N_235,N_437);
nand U798 (N_798,N_54,N_259);
nand U799 (N_799,N_101,N_430);
nand U800 (N_800,N_501,N_42);
or U801 (N_801,N_528,N_104);
nand U802 (N_802,N_76,N_561);
nor U803 (N_803,N_506,N_507);
nor U804 (N_804,N_169,N_215);
and U805 (N_805,N_322,N_125);
nand U806 (N_806,N_158,N_547);
or U807 (N_807,N_427,N_163);
nor U808 (N_808,N_293,N_291);
nor U809 (N_809,N_250,N_99);
nand U810 (N_810,N_311,N_277);
nor U811 (N_811,N_71,N_512);
and U812 (N_812,N_580,N_185);
nand U813 (N_813,N_596,N_211);
nor U814 (N_814,N_476,N_453);
and U815 (N_815,N_193,N_21);
nor U816 (N_816,N_360,N_102);
nand U817 (N_817,N_278,N_336);
and U818 (N_818,N_314,N_331);
or U819 (N_819,N_274,N_329);
nor U820 (N_820,N_38,N_228);
or U821 (N_821,N_570,N_403);
nor U822 (N_822,N_13,N_433);
nand U823 (N_823,N_358,N_150);
nand U824 (N_824,N_521,N_583);
nand U825 (N_825,N_300,N_364);
nand U826 (N_826,N_183,N_178);
or U827 (N_827,N_497,N_562);
or U828 (N_828,N_103,N_2);
nand U829 (N_829,N_151,N_299);
nand U830 (N_830,N_417,N_281);
nor U831 (N_831,N_187,N_223);
nor U832 (N_832,N_565,N_58);
or U833 (N_833,N_584,N_513);
or U834 (N_834,N_266,N_145);
nor U835 (N_835,N_522,N_410);
nand U836 (N_836,N_564,N_273);
and U837 (N_837,N_209,N_567);
or U838 (N_838,N_6,N_109);
or U839 (N_839,N_57,N_362);
or U840 (N_840,N_481,N_129);
nor U841 (N_841,N_308,N_10);
nand U842 (N_842,N_269,N_424);
and U843 (N_843,N_333,N_121);
nor U844 (N_844,N_271,N_305);
nor U845 (N_845,N_556,N_366);
or U846 (N_846,N_45,N_275);
and U847 (N_847,N_12,N_418);
xnor U848 (N_848,N_100,N_502);
and U849 (N_849,N_165,N_43);
nand U850 (N_850,N_585,N_525);
and U851 (N_851,N_508,N_376);
or U852 (N_852,N_63,N_434);
and U853 (N_853,N_166,N_394);
and U854 (N_854,N_55,N_29);
nand U855 (N_855,N_139,N_117);
and U856 (N_856,N_534,N_195);
or U857 (N_857,N_177,N_505);
and U858 (N_858,N_268,N_390);
nand U859 (N_859,N_415,N_52);
or U860 (N_860,N_267,N_389);
nand U861 (N_861,N_342,N_47);
nand U862 (N_862,N_514,N_368);
or U863 (N_863,N_62,N_545);
nor U864 (N_864,N_297,N_372);
or U865 (N_865,N_529,N_578);
nand U866 (N_866,N_555,N_39);
nor U867 (N_867,N_348,N_252);
nor U868 (N_868,N_181,N_118);
and U869 (N_869,N_201,N_61);
nor U870 (N_870,N_153,N_558);
and U871 (N_871,N_0,N_20);
nor U872 (N_872,N_509,N_425);
or U873 (N_873,N_345,N_17);
and U874 (N_874,N_146,N_156);
and U875 (N_875,N_542,N_381);
nor U876 (N_876,N_251,N_378);
or U877 (N_877,N_16,N_188);
or U878 (N_878,N_451,N_212);
and U879 (N_879,N_191,N_568);
or U880 (N_880,N_343,N_30);
or U881 (N_881,N_128,N_591);
and U882 (N_882,N_221,N_460);
nor U883 (N_883,N_115,N_592);
or U884 (N_884,N_436,N_548);
or U885 (N_885,N_500,N_312);
and U886 (N_886,N_469,N_518);
or U887 (N_887,N_40,N_530);
nand U888 (N_888,N_452,N_210);
nand U889 (N_889,N_557,N_148);
or U890 (N_890,N_68,N_351);
and U891 (N_891,N_550,N_370);
nand U892 (N_892,N_141,N_184);
xnor U893 (N_893,N_213,N_132);
and U894 (N_894,N_357,N_168);
or U895 (N_895,N_332,N_349);
nor U896 (N_896,N_408,N_242);
nor U897 (N_897,N_493,N_594);
and U898 (N_898,N_398,N_200);
or U899 (N_899,N_459,N_423);
nand U900 (N_900,N_379,N_197);
nand U901 (N_901,N_112,N_3);
and U902 (N_902,N_492,N_579);
and U903 (N_903,N_168,N_232);
or U904 (N_904,N_293,N_42);
and U905 (N_905,N_500,N_238);
and U906 (N_906,N_268,N_224);
nor U907 (N_907,N_594,N_205);
and U908 (N_908,N_211,N_96);
and U909 (N_909,N_39,N_236);
nor U910 (N_910,N_198,N_15);
nor U911 (N_911,N_570,N_567);
nor U912 (N_912,N_495,N_383);
nand U913 (N_913,N_491,N_413);
nand U914 (N_914,N_369,N_130);
nor U915 (N_915,N_5,N_273);
and U916 (N_916,N_553,N_376);
nor U917 (N_917,N_7,N_515);
and U918 (N_918,N_224,N_287);
nor U919 (N_919,N_442,N_428);
nand U920 (N_920,N_448,N_387);
and U921 (N_921,N_410,N_122);
and U922 (N_922,N_166,N_490);
nor U923 (N_923,N_365,N_312);
nor U924 (N_924,N_555,N_479);
nor U925 (N_925,N_476,N_76);
or U926 (N_926,N_178,N_446);
and U927 (N_927,N_265,N_275);
nand U928 (N_928,N_527,N_510);
or U929 (N_929,N_60,N_56);
nor U930 (N_930,N_60,N_397);
nand U931 (N_931,N_271,N_274);
nand U932 (N_932,N_3,N_282);
or U933 (N_933,N_586,N_346);
or U934 (N_934,N_244,N_239);
nor U935 (N_935,N_500,N_308);
and U936 (N_936,N_193,N_114);
and U937 (N_937,N_383,N_69);
nor U938 (N_938,N_300,N_256);
nand U939 (N_939,N_223,N_394);
or U940 (N_940,N_573,N_231);
nor U941 (N_941,N_148,N_149);
nor U942 (N_942,N_536,N_404);
nand U943 (N_943,N_183,N_333);
nand U944 (N_944,N_47,N_336);
nand U945 (N_945,N_12,N_484);
or U946 (N_946,N_111,N_506);
or U947 (N_947,N_13,N_492);
or U948 (N_948,N_403,N_193);
nor U949 (N_949,N_524,N_274);
and U950 (N_950,N_147,N_508);
and U951 (N_951,N_309,N_103);
or U952 (N_952,N_433,N_170);
or U953 (N_953,N_70,N_60);
or U954 (N_954,N_592,N_315);
and U955 (N_955,N_370,N_328);
nor U956 (N_956,N_211,N_267);
and U957 (N_957,N_352,N_307);
or U958 (N_958,N_66,N_117);
and U959 (N_959,N_17,N_330);
nand U960 (N_960,N_35,N_229);
nor U961 (N_961,N_177,N_84);
nand U962 (N_962,N_33,N_181);
xor U963 (N_963,N_494,N_208);
nand U964 (N_964,N_184,N_372);
and U965 (N_965,N_555,N_119);
nor U966 (N_966,N_105,N_141);
nor U967 (N_967,N_211,N_174);
and U968 (N_968,N_456,N_368);
or U969 (N_969,N_368,N_548);
nand U970 (N_970,N_473,N_374);
and U971 (N_971,N_444,N_142);
and U972 (N_972,N_168,N_41);
or U973 (N_973,N_55,N_267);
and U974 (N_974,N_447,N_129);
or U975 (N_975,N_416,N_518);
or U976 (N_976,N_173,N_298);
nand U977 (N_977,N_2,N_543);
nand U978 (N_978,N_140,N_453);
xnor U979 (N_979,N_502,N_3);
nand U980 (N_980,N_339,N_278);
nand U981 (N_981,N_579,N_393);
and U982 (N_982,N_388,N_327);
and U983 (N_983,N_385,N_146);
or U984 (N_984,N_274,N_341);
and U985 (N_985,N_135,N_566);
or U986 (N_986,N_456,N_382);
and U987 (N_987,N_576,N_69);
or U988 (N_988,N_10,N_53);
and U989 (N_989,N_173,N_14);
nor U990 (N_990,N_590,N_4);
nor U991 (N_991,N_252,N_420);
nor U992 (N_992,N_130,N_565);
and U993 (N_993,N_41,N_113);
nand U994 (N_994,N_281,N_165);
nand U995 (N_995,N_313,N_263);
nand U996 (N_996,N_192,N_189);
nand U997 (N_997,N_26,N_189);
or U998 (N_998,N_216,N_38);
or U999 (N_999,N_494,N_89);
or U1000 (N_1000,N_433,N_91);
nand U1001 (N_1001,N_401,N_50);
nor U1002 (N_1002,N_556,N_495);
nand U1003 (N_1003,N_449,N_69);
or U1004 (N_1004,N_464,N_337);
nor U1005 (N_1005,N_506,N_340);
or U1006 (N_1006,N_346,N_521);
nor U1007 (N_1007,N_468,N_4);
nor U1008 (N_1008,N_314,N_470);
and U1009 (N_1009,N_111,N_109);
and U1010 (N_1010,N_437,N_102);
nor U1011 (N_1011,N_300,N_83);
or U1012 (N_1012,N_157,N_559);
or U1013 (N_1013,N_110,N_102);
or U1014 (N_1014,N_430,N_486);
nor U1015 (N_1015,N_421,N_273);
or U1016 (N_1016,N_424,N_200);
or U1017 (N_1017,N_425,N_128);
and U1018 (N_1018,N_12,N_386);
or U1019 (N_1019,N_276,N_154);
and U1020 (N_1020,N_58,N_130);
or U1021 (N_1021,N_187,N_525);
and U1022 (N_1022,N_113,N_272);
nor U1023 (N_1023,N_227,N_127);
nand U1024 (N_1024,N_80,N_179);
nand U1025 (N_1025,N_203,N_77);
or U1026 (N_1026,N_305,N_157);
and U1027 (N_1027,N_410,N_232);
nor U1028 (N_1028,N_435,N_14);
nor U1029 (N_1029,N_331,N_362);
and U1030 (N_1030,N_104,N_458);
nor U1031 (N_1031,N_322,N_559);
nor U1032 (N_1032,N_447,N_256);
nand U1033 (N_1033,N_121,N_241);
and U1034 (N_1034,N_509,N_350);
or U1035 (N_1035,N_300,N_505);
and U1036 (N_1036,N_394,N_280);
or U1037 (N_1037,N_173,N_432);
nor U1038 (N_1038,N_215,N_159);
or U1039 (N_1039,N_31,N_336);
and U1040 (N_1040,N_90,N_443);
or U1041 (N_1041,N_425,N_244);
and U1042 (N_1042,N_457,N_42);
or U1043 (N_1043,N_98,N_379);
or U1044 (N_1044,N_34,N_140);
nand U1045 (N_1045,N_476,N_95);
nor U1046 (N_1046,N_206,N_49);
nor U1047 (N_1047,N_219,N_65);
nand U1048 (N_1048,N_207,N_366);
nor U1049 (N_1049,N_529,N_346);
nand U1050 (N_1050,N_287,N_186);
or U1051 (N_1051,N_119,N_291);
nor U1052 (N_1052,N_45,N_506);
and U1053 (N_1053,N_394,N_526);
nor U1054 (N_1054,N_377,N_545);
and U1055 (N_1055,N_191,N_325);
nor U1056 (N_1056,N_498,N_105);
nor U1057 (N_1057,N_157,N_129);
or U1058 (N_1058,N_363,N_135);
or U1059 (N_1059,N_570,N_353);
and U1060 (N_1060,N_491,N_386);
nor U1061 (N_1061,N_208,N_101);
nor U1062 (N_1062,N_530,N_87);
or U1063 (N_1063,N_452,N_113);
and U1064 (N_1064,N_160,N_25);
or U1065 (N_1065,N_103,N_427);
nand U1066 (N_1066,N_319,N_393);
and U1067 (N_1067,N_13,N_544);
nand U1068 (N_1068,N_539,N_220);
and U1069 (N_1069,N_62,N_298);
nand U1070 (N_1070,N_273,N_538);
nor U1071 (N_1071,N_461,N_92);
or U1072 (N_1072,N_181,N_43);
nor U1073 (N_1073,N_308,N_129);
nor U1074 (N_1074,N_383,N_385);
nand U1075 (N_1075,N_216,N_343);
or U1076 (N_1076,N_214,N_25);
nor U1077 (N_1077,N_527,N_28);
nand U1078 (N_1078,N_222,N_493);
nor U1079 (N_1079,N_107,N_116);
and U1080 (N_1080,N_411,N_98);
or U1081 (N_1081,N_42,N_452);
and U1082 (N_1082,N_37,N_488);
nand U1083 (N_1083,N_109,N_330);
and U1084 (N_1084,N_281,N_587);
nand U1085 (N_1085,N_445,N_194);
or U1086 (N_1086,N_229,N_531);
or U1087 (N_1087,N_234,N_10);
nor U1088 (N_1088,N_480,N_351);
and U1089 (N_1089,N_145,N_60);
nor U1090 (N_1090,N_88,N_443);
nor U1091 (N_1091,N_506,N_390);
nand U1092 (N_1092,N_343,N_345);
nand U1093 (N_1093,N_340,N_198);
or U1094 (N_1094,N_217,N_407);
and U1095 (N_1095,N_591,N_595);
nor U1096 (N_1096,N_589,N_412);
nand U1097 (N_1097,N_307,N_219);
and U1098 (N_1098,N_46,N_82);
or U1099 (N_1099,N_564,N_70);
nor U1100 (N_1100,N_417,N_457);
nand U1101 (N_1101,N_192,N_87);
or U1102 (N_1102,N_471,N_259);
or U1103 (N_1103,N_225,N_511);
or U1104 (N_1104,N_330,N_67);
nor U1105 (N_1105,N_517,N_161);
nor U1106 (N_1106,N_124,N_270);
nand U1107 (N_1107,N_296,N_220);
or U1108 (N_1108,N_414,N_37);
and U1109 (N_1109,N_449,N_30);
and U1110 (N_1110,N_531,N_86);
or U1111 (N_1111,N_547,N_129);
nor U1112 (N_1112,N_159,N_580);
nand U1113 (N_1113,N_111,N_120);
nor U1114 (N_1114,N_48,N_404);
nand U1115 (N_1115,N_78,N_567);
or U1116 (N_1116,N_373,N_21);
or U1117 (N_1117,N_354,N_1);
or U1118 (N_1118,N_212,N_449);
nand U1119 (N_1119,N_340,N_508);
or U1120 (N_1120,N_88,N_435);
nand U1121 (N_1121,N_79,N_542);
nor U1122 (N_1122,N_303,N_412);
nor U1123 (N_1123,N_452,N_50);
and U1124 (N_1124,N_208,N_268);
nor U1125 (N_1125,N_440,N_432);
nor U1126 (N_1126,N_252,N_506);
nand U1127 (N_1127,N_493,N_236);
nor U1128 (N_1128,N_74,N_423);
nor U1129 (N_1129,N_571,N_166);
nor U1130 (N_1130,N_340,N_273);
nor U1131 (N_1131,N_19,N_130);
nand U1132 (N_1132,N_349,N_574);
or U1133 (N_1133,N_327,N_572);
and U1134 (N_1134,N_153,N_237);
nor U1135 (N_1135,N_573,N_429);
and U1136 (N_1136,N_255,N_297);
or U1137 (N_1137,N_470,N_110);
nor U1138 (N_1138,N_96,N_592);
or U1139 (N_1139,N_513,N_562);
nor U1140 (N_1140,N_67,N_336);
nor U1141 (N_1141,N_203,N_441);
nor U1142 (N_1142,N_36,N_461);
and U1143 (N_1143,N_32,N_529);
or U1144 (N_1144,N_157,N_432);
and U1145 (N_1145,N_160,N_500);
or U1146 (N_1146,N_207,N_127);
nand U1147 (N_1147,N_224,N_56);
nor U1148 (N_1148,N_502,N_414);
nand U1149 (N_1149,N_594,N_89);
nand U1150 (N_1150,N_1,N_326);
nor U1151 (N_1151,N_537,N_75);
nand U1152 (N_1152,N_475,N_279);
nor U1153 (N_1153,N_47,N_430);
or U1154 (N_1154,N_275,N_542);
or U1155 (N_1155,N_313,N_233);
nand U1156 (N_1156,N_314,N_377);
nand U1157 (N_1157,N_583,N_273);
nor U1158 (N_1158,N_127,N_137);
nor U1159 (N_1159,N_586,N_460);
nor U1160 (N_1160,N_578,N_429);
and U1161 (N_1161,N_364,N_381);
and U1162 (N_1162,N_137,N_390);
and U1163 (N_1163,N_480,N_409);
or U1164 (N_1164,N_550,N_326);
nand U1165 (N_1165,N_598,N_521);
and U1166 (N_1166,N_64,N_565);
or U1167 (N_1167,N_267,N_471);
and U1168 (N_1168,N_462,N_1);
nor U1169 (N_1169,N_236,N_232);
and U1170 (N_1170,N_516,N_21);
nand U1171 (N_1171,N_108,N_532);
nand U1172 (N_1172,N_323,N_599);
and U1173 (N_1173,N_3,N_584);
nor U1174 (N_1174,N_542,N_447);
and U1175 (N_1175,N_116,N_271);
and U1176 (N_1176,N_503,N_281);
or U1177 (N_1177,N_69,N_564);
and U1178 (N_1178,N_42,N_437);
and U1179 (N_1179,N_584,N_467);
and U1180 (N_1180,N_499,N_227);
or U1181 (N_1181,N_387,N_518);
nor U1182 (N_1182,N_499,N_472);
nor U1183 (N_1183,N_71,N_394);
or U1184 (N_1184,N_511,N_589);
or U1185 (N_1185,N_534,N_276);
and U1186 (N_1186,N_37,N_516);
nor U1187 (N_1187,N_86,N_518);
nand U1188 (N_1188,N_529,N_509);
and U1189 (N_1189,N_226,N_178);
and U1190 (N_1190,N_150,N_540);
nand U1191 (N_1191,N_423,N_312);
nor U1192 (N_1192,N_264,N_226);
nand U1193 (N_1193,N_555,N_348);
nand U1194 (N_1194,N_342,N_159);
nand U1195 (N_1195,N_289,N_518);
nor U1196 (N_1196,N_431,N_12);
nand U1197 (N_1197,N_271,N_408);
nand U1198 (N_1198,N_314,N_492);
nor U1199 (N_1199,N_69,N_130);
and U1200 (N_1200,N_931,N_1172);
and U1201 (N_1201,N_757,N_627);
nand U1202 (N_1202,N_750,N_958);
nor U1203 (N_1203,N_809,N_1007);
and U1204 (N_1204,N_670,N_992);
and U1205 (N_1205,N_1063,N_1197);
and U1206 (N_1206,N_957,N_788);
nor U1207 (N_1207,N_791,N_1159);
or U1208 (N_1208,N_1150,N_999);
and U1209 (N_1209,N_1141,N_853);
and U1210 (N_1210,N_681,N_1066);
and U1211 (N_1211,N_756,N_994);
nor U1212 (N_1212,N_644,N_888);
or U1213 (N_1213,N_1006,N_1005);
or U1214 (N_1214,N_612,N_688);
nor U1215 (N_1215,N_1021,N_1056);
or U1216 (N_1216,N_658,N_872);
nor U1217 (N_1217,N_876,N_921);
or U1218 (N_1218,N_881,N_641);
and U1219 (N_1219,N_1118,N_600);
nor U1220 (N_1220,N_1017,N_1038);
nor U1221 (N_1221,N_653,N_1097);
nand U1222 (N_1222,N_747,N_655);
nor U1223 (N_1223,N_669,N_1047);
nand U1224 (N_1224,N_822,N_649);
or U1225 (N_1225,N_1127,N_717);
and U1226 (N_1226,N_1036,N_713);
nand U1227 (N_1227,N_1057,N_942);
or U1228 (N_1228,N_1155,N_810);
nor U1229 (N_1229,N_870,N_1042);
nand U1230 (N_1230,N_639,N_718);
and U1231 (N_1231,N_1078,N_904);
nor U1232 (N_1232,N_1163,N_1059);
nor U1233 (N_1233,N_730,N_825);
and U1234 (N_1234,N_826,N_640);
or U1235 (N_1235,N_1094,N_613);
and U1236 (N_1236,N_898,N_603);
and U1237 (N_1237,N_1187,N_961);
or U1238 (N_1238,N_1028,N_917);
and U1239 (N_1239,N_1000,N_980);
and U1240 (N_1240,N_787,N_871);
or U1241 (N_1241,N_1031,N_831);
xor U1242 (N_1242,N_650,N_857);
or U1243 (N_1243,N_624,N_910);
and U1244 (N_1244,N_947,N_836);
and U1245 (N_1245,N_847,N_1024);
nand U1246 (N_1246,N_1122,N_715);
nor U1247 (N_1247,N_1195,N_767);
and U1248 (N_1248,N_708,N_1162);
nor U1249 (N_1249,N_667,N_753);
and U1250 (N_1250,N_657,N_1130);
nand U1251 (N_1251,N_1107,N_834);
nand U1252 (N_1252,N_944,N_893);
and U1253 (N_1253,N_979,N_937);
nand U1254 (N_1254,N_1064,N_1022);
nor U1255 (N_1255,N_1085,N_1117);
nand U1256 (N_1256,N_816,N_647);
or U1257 (N_1257,N_1039,N_666);
or U1258 (N_1258,N_1009,N_1161);
nor U1259 (N_1259,N_812,N_776);
and U1260 (N_1260,N_1061,N_1087);
nor U1261 (N_1261,N_1138,N_1091);
nor U1262 (N_1262,N_780,N_1167);
nand U1263 (N_1263,N_790,N_785);
and U1264 (N_1264,N_1067,N_965);
nand U1265 (N_1265,N_697,N_779);
nor U1266 (N_1266,N_1192,N_799);
or U1267 (N_1267,N_751,N_850);
or U1268 (N_1268,N_900,N_820);
or U1269 (N_1269,N_854,N_1133);
or U1270 (N_1270,N_977,N_913);
or U1271 (N_1271,N_861,N_967);
nand U1272 (N_1272,N_1121,N_929);
nor U1273 (N_1273,N_1025,N_629);
and U1274 (N_1274,N_997,N_731);
nor U1275 (N_1275,N_795,N_839);
nand U1276 (N_1276,N_694,N_687);
nor U1277 (N_1277,N_941,N_927);
nor U1278 (N_1278,N_1041,N_1132);
nand U1279 (N_1279,N_919,N_887);
or U1280 (N_1280,N_1196,N_1105);
and U1281 (N_1281,N_766,N_1108);
nor U1282 (N_1282,N_995,N_1136);
nand U1283 (N_1283,N_609,N_1016);
nor U1284 (N_1284,N_891,N_877);
or U1285 (N_1285,N_763,N_869);
or U1286 (N_1286,N_698,N_863);
nand U1287 (N_1287,N_956,N_1128);
or U1288 (N_1288,N_680,N_843);
and U1289 (N_1289,N_824,N_1158);
nand U1290 (N_1290,N_914,N_659);
nor U1291 (N_1291,N_915,N_761);
nor U1292 (N_1292,N_1112,N_936);
nor U1293 (N_1293,N_846,N_923);
nand U1294 (N_1294,N_679,N_840);
nor U1295 (N_1295,N_890,N_668);
or U1296 (N_1296,N_725,N_1154);
or U1297 (N_1297,N_844,N_823);
and U1298 (N_1298,N_983,N_671);
and U1299 (N_1299,N_648,N_622);
nand U1300 (N_1300,N_616,N_752);
and U1301 (N_1301,N_912,N_1075);
and U1302 (N_1302,N_608,N_741);
nand U1303 (N_1303,N_651,N_1173);
nor U1304 (N_1304,N_1052,N_883);
nor U1305 (N_1305,N_726,N_768);
nor U1306 (N_1306,N_625,N_973);
or U1307 (N_1307,N_852,N_1008);
nor U1308 (N_1308,N_1184,N_692);
and U1309 (N_1309,N_925,N_971);
nand U1310 (N_1310,N_703,N_990);
or U1311 (N_1311,N_646,N_827);
or U1312 (N_1312,N_833,N_974);
and U1313 (N_1313,N_714,N_631);
nand U1314 (N_1314,N_738,N_989);
nor U1315 (N_1315,N_691,N_1058);
nor U1316 (N_1316,N_885,N_1046);
nor U1317 (N_1317,N_1106,N_1190);
and U1318 (N_1318,N_946,N_772);
or U1319 (N_1319,N_792,N_902);
nor U1320 (N_1320,N_832,N_894);
nor U1321 (N_1321,N_606,N_793);
and U1322 (N_1322,N_742,N_1160);
nand U1323 (N_1323,N_699,N_722);
nand U1324 (N_1324,N_709,N_797);
nor U1325 (N_1325,N_1142,N_1020);
and U1326 (N_1326,N_734,N_801);
and U1327 (N_1327,N_1169,N_862);
nor U1328 (N_1328,N_950,N_1065);
nand U1329 (N_1329,N_719,N_908);
or U1330 (N_1330,N_728,N_1177);
or U1331 (N_1331,N_1082,N_1072);
nand U1332 (N_1332,N_638,N_1183);
and U1333 (N_1333,N_1090,N_866);
and U1334 (N_1334,N_1111,N_656);
nand U1335 (N_1335,N_951,N_633);
nor U1336 (N_1336,N_1018,N_849);
and U1337 (N_1337,N_777,N_918);
nor U1338 (N_1338,N_1026,N_909);
nor U1339 (N_1339,N_1001,N_1043);
nor U1340 (N_1340,N_1149,N_1140);
nand U1341 (N_1341,N_884,N_978);
and U1342 (N_1342,N_986,N_838);
nand U1343 (N_1343,N_837,N_1174);
nor U1344 (N_1344,N_1030,N_1102);
xnor U1345 (N_1345,N_605,N_601);
and U1346 (N_1346,N_701,N_604);
or U1347 (N_1347,N_618,N_855);
or U1348 (N_1348,N_781,N_773);
nor U1349 (N_1349,N_1083,N_1080);
nor U1350 (N_1350,N_1034,N_611);
or U1351 (N_1351,N_1114,N_945);
nor U1352 (N_1352,N_1126,N_702);
nand U1353 (N_1353,N_1179,N_959);
nor U1354 (N_1354,N_1151,N_819);
xor U1355 (N_1355,N_1168,N_1048);
and U1356 (N_1356,N_758,N_1170);
nand U1357 (N_1357,N_930,N_1033);
and U1358 (N_1358,N_1123,N_1113);
nor U1359 (N_1359,N_802,N_993);
or U1360 (N_1360,N_953,N_664);
and U1361 (N_1361,N_1079,N_673);
xnor U1362 (N_1362,N_859,N_952);
nand U1363 (N_1363,N_814,N_848);
nor U1364 (N_1364,N_879,N_1050);
nor U1365 (N_1365,N_628,N_686);
and U1366 (N_1366,N_1076,N_743);
or U1367 (N_1367,N_732,N_693);
nor U1368 (N_1368,N_774,N_1040);
and U1369 (N_1369,N_830,N_1089);
nor U1370 (N_1370,N_1077,N_783);
nand U1371 (N_1371,N_602,N_733);
nand U1372 (N_1372,N_782,N_706);
nand U1373 (N_1373,N_1131,N_1186);
nand U1374 (N_1374,N_1032,N_1099);
nand U1375 (N_1375,N_710,N_1011);
or U1376 (N_1376,N_932,N_1101);
or U1377 (N_1377,N_928,N_991);
nor U1378 (N_1378,N_896,N_1068);
nand U1379 (N_1379,N_1182,N_610);
nor U1380 (N_1380,N_829,N_1088);
or U1381 (N_1381,N_845,N_1002);
and U1382 (N_1382,N_665,N_939);
and U1383 (N_1383,N_765,N_723);
or U1384 (N_1384,N_720,N_1104);
nor U1385 (N_1385,N_1027,N_642);
nand U1386 (N_1386,N_740,N_778);
nand U1387 (N_1387,N_806,N_1037);
nand U1388 (N_1388,N_821,N_1055);
nand U1389 (N_1389,N_878,N_684);
nor U1390 (N_1390,N_672,N_721);
or U1391 (N_1391,N_736,N_1093);
or U1392 (N_1392,N_1164,N_1125);
nand U1393 (N_1393,N_796,N_815);
nand U1394 (N_1394,N_865,N_700);
nand U1395 (N_1395,N_615,N_1178);
nand U1396 (N_1396,N_935,N_1191);
and U1397 (N_1397,N_784,N_800);
and U1398 (N_1398,N_770,N_916);
nor U1399 (N_1399,N_828,N_972);
or U1400 (N_1400,N_963,N_798);
nand U1401 (N_1401,N_704,N_1147);
or U1402 (N_1402,N_1148,N_911);
and U1403 (N_1403,N_1069,N_1073);
nand U1404 (N_1404,N_841,N_634);
nand U1405 (N_1405,N_716,N_907);
and U1406 (N_1406,N_851,N_1139);
nand U1407 (N_1407,N_689,N_696);
nand U1408 (N_1408,N_744,N_678);
nor U1409 (N_1409,N_985,N_988);
nor U1410 (N_1410,N_674,N_660);
nand U1411 (N_1411,N_1062,N_676);
nand U1412 (N_1412,N_835,N_1003);
and U1413 (N_1413,N_1054,N_707);
and U1414 (N_1414,N_1096,N_663);
and U1415 (N_1415,N_636,N_964);
xor U1416 (N_1416,N_955,N_1189);
or U1417 (N_1417,N_760,N_1060);
nor U1418 (N_1418,N_899,N_755);
nand U1419 (N_1419,N_1100,N_1012);
nand U1420 (N_1420,N_922,N_635);
or U1421 (N_1421,N_818,N_735);
nand U1422 (N_1422,N_984,N_817);
nand U1423 (N_1423,N_969,N_739);
or U1424 (N_1424,N_1044,N_938);
or U1425 (N_1425,N_654,N_764);
nor U1426 (N_1426,N_1188,N_1181);
nand U1427 (N_1427,N_632,N_1152);
nand U1428 (N_1428,N_1157,N_1103);
or U1429 (N_1429,N_1180,N_1144);
and U1430 (N_1430,N_1081,N_1166);
and U1431 (N_1431,N_1175,N_968);
and U1432 (N_1432,N_1023,N_607);
nand U1433 (N_1433,N_1145,N_874);
nor U1434 (N_1434,N_749,N_794);
or U1435 (N_1435,N_620,N_1193);
and U1436 (N_1436,N_1176,N_1092);
and U1437 (N_1437,N_868,N_905);
nor U1438 (N_1438,N_1035,N_976);
nor U1439 (N_1439,N_711,N_1071);
and U1440 (N_1440,N_903,N_1115);
or U1441 (N_1441,N_645,N_1134);
nand U1442 (N_1442,N_1165,N_954);
or U1443 (N_1443,N_1110,N_970);
nor U1444 (N_1444,N_1124,N_1010);
nor U1445 (N_1445,N_1070,N_1095);
and U1446 (N_1446,N_748,N_1015);
nand U1447 (N_1447,N_1153,N_775);
or U1448 (N_1448,N_1051,N_727);
nand U1449 (N_1449,N_705,N_729);
and U1450 (N_1450,N_808,N_737);
or U1451 (N_1451,N_695,N_682);
nor U1452 (N_1452,N_643,N_1185);
and U1453 (N_1453,N_626,N_762);
nor U1454 (N_1454,N_811,N_614);
and U1455 (N_1455,N_637,N_803);
nor U1456 (N_1456,N_1198,N_1137);
nor U1457 (N_1457,N_867,N_1143);
and U1458 (N_1458,N_1086,N_886);
and U1459 (N_1459,N_1199,N_880);
and U1460 (N_1460,N_1120,N_949);
and U1461 (N_1461,N_975,N_875);
nand U1462 (N_1462,N_1119,N_882);
nor U1463 (N_1463,N_1109,N_786);
xnor U1464 (N_1464,N_617,N_860);
nor U1465 (N_1465,N_1129,N_858);
and U1466 (N_1466,N_789,N_920);
xnor U1467 (N_1467,N_926,N_873);
or U1468 (N_1468,N_805,N_677);
and U1469 (N_1469,N_662,N_1045);
and U1470 (N_1470,N_864,N_960);
nor U1471 (N_1471,N_892,N_998);
and U1472 (N_1472,N_712,N_661);
and U1473 (N_1473,N_675,N_1156);
nor U1474 (N_1474,N_813,N_771);
nor U1475 (N_1475,N_746,N_895);
or U1476 (N_1476,N_1004,N_982);
or U1477 (N_1477,N_943,N_934);
nand U1478 (N_1478,N_1135,N_683);
or U1479 (N_1479,N_1049,N_1019);
or U1480 (N_1480,N_981,N_621);
and U1481 (N_1481,N_690,N_685);
or U1482 (N_1482,N_1084,N_901);
and U1483 (N_1483,N_807,N_652);
nand U1484 (N_1484,N_924,N_724);
nand U1485 (N_1485,N_966,N_1116);
or U1486 (N_1486,N_1146,N_948);
and U1487 (N_1487,N_842,N_962);
or U1488 (N_1488,N_1053,N_1098);
nor U1489 (N_1489,N_623,N_1029);
and U1490 (N_1490,N_630,N_889);
nand U1491 (N_1491,N_1014,N_619);
nand U1492 (N_1492,N_1013,N_754);
and U1493 (N_1493,N_856,N_940);
nor U1494 (N_1494,N_1074,N_987);
or U1495 (N_1495,N_759,N_1171);
and U1496 (N_1496,N_906,N_804);
nor U1497 (N_1497,N_1194,N_897);
or U1498 (N_1498,N_996,N_745);
nand U1499 (N_1499,N_933,N_769);
and U1500 (N_1500,N_838,N_894);
nor U1501 (N_1501,N_717,N_624);
or U1502 (N_1502,N_818,N_1003);
and U1503 (N_1503,N_960,N_816);
nor U1504 (N_1504,N_973,N_896);
or U1505 (N_1505,N_640,N_627);
or U1506 (N_1506,N_754,N_694);
and U1507 (N_1507,N_606,N_1033);
nor U1508 (N_1508,N_727,N_770);
nor U1509 (N_1509,N_811,N_1045);
nand U1510 (N_1510,N_1051,N_866);
nand U1511 (N_1511,N_828,N_830);
nor U1512 (N_1512,N_629,N_920);
nand U1513 (N_1513,N_1153,N_716);
and U1514 (N_1514,N_1144,N_1022);
or U1515 (N_1515,N_1186,N_903);
and U1516 (N_1516,N_892,N_758);
nand U1517 (N_1517,N_747,N_829);
and U1518 (N_1518,N_624,N_785);
and U1519 (N_1519,N_786,N_1088);
and U1520 (N_1520,N_601,N_756);
and U1521 (N_1521,N_721,N_756);
nor U1522 (N_1522,N_706,N_1161);
nand U1523 (N_1523,N_831,N_985);
nand U1524 (N_1524,N_858,N_1110);
and U1525 (N_1525,N_1151,N_1168);
nand U1526 (N_1526,N_803,N_765);
nand U1527 (N_1527,N_991,N_1129);
or U1528 (N_1528,N_1171,N_981);
and U1529 (N_1529,N_873,N_776);
nor U1530 (N_1530,N_970,N_716);
and U1531 (N_1531,N_1120,N_743);
or U1532 (N_1532,N_946,N_622);
or U1533 (N_1533,N_1133,N_848);
nand U1534 (N_1534,N_1099,N_967);
and U1535 (N_1535,N_601,N_939);
nand U1536 (N_1536,N_764,N_945);
and U1537 (N_1537,N_872,N_959);
nand U1538 (N_1538,N_646,N_791);
nor U1539 (N_1539,N_621,N_777);
nor U1540 (N_1540,N_983,N_820);
nor U1541 (N_1541,N_1122,N_938);
nor U1542 (N_1542,N_1063,N_951);
or U1543 (N_1543,N_893,N_897);
nor U1544 (N_1544,N_779,N_935);
nand U1545 (N_1545,N_1159,N_939);
or U1546 (N_1546,N_721,N_877);
nor U1547 (N_1547,N_1005,N_805);
or U1548 (N_1548,N_875,N_819);
or U1549 (N_1549,N_1017,N_861);
or U1550 (N_1550,N_610,N_891);
nor U1551 (N_1551,N_692,N_1130);
nor U1552 (N_1552,N_916,N_1000);
or U1553 (N_1553,N_743,N_744);
nor U1554 (N_1554,N_696,N_1059);
and U1555 (N_1555,N_775,N_887);
nand U1556 (N_1556,N_719,N_767);
and U1557 (N_1557,N_872,N_886);
nand U1558 (N_1558,N_951,N_617);
nand U1559 (N_1559,N_948,N_1116);
nand U1560 (N_1560,N_1059,N_1054);
nor U1561 (N_1561,N_1089,N_615);
nand U1562 (N_1562,N_903,N_972);
or U1563 (N_1563,N_901,N_853);
nand U1564 (N_1564,N_749,N_914);
and U1565 (N_1565,N_993,N_790);
or U1566 (N_1566,N_1079,N_814);
or U1567 (N_1567,N_743,N_1015);
and U1568 (N_1568,N_983,N_1053);
nand U1569 (N_1569,N_1162,N_1115);
nand U1570 (N_1570,N_633,N_974);
nor U1571 (N_1571,N_624,N_856);
or U1572 (N_1572,N_661,N_1049);
and U1573 (N_1573,N_677,N_602);
and U1574 (N_1574,N_1149,N_762);
nand U1575 (N_1575,N_801,N_1132);
or U1576 (N_1576,N_1112,N_1095);
nand U1577 (N_1577,N_644,N_1025);
or U1578 (N_1578,N_1193,N_1019);
nand U1579 (N_1579,N_865,N_1103);
and U1580 (N_1580,N_710,N_628);
or U1581 (N_1581,N_632,N_770);
nand U1582 (N_1582,N_870,N_793);
and U1583 (N_1583,N_905,N_1057);
and U1584 (N_1584,N_1173,N_604);
and U1585 (N_1585,N_679,N_1105);
nand U1586 (N_1586,N_688,N_606);
or U1587 (N_1587,N_921,N_1188);
or U1588 (N_1588,N_777,N_765);
nand U1589 (N_1589,N_1115,N_1075);
nand U1590 (N_1590,N_800,N_692);
or U1591 (N_1591,N_705,N_1017);
or U1592 (N_1592,N_787,N_741);
nand U1593 (N_1593,N_725,N_908);
or U1594 (N_1594,N_844,N_915);
nand U1595 (N_1595,N_664,N_915);
nand U1596 (N_1596,N_931,N_716);
nor U1597 (N_1597,N_1124,N_674);
or U1598 (N_1598,N_815,N_707);
nand U1599 (N_1599,N_715,N_750);
and U1600 (N_1600,N_948,N_1053);
nor U1601 (N_1601,N_1092,N_700);
nand U1602 (N_1602,N_633,N_693);
or U1603 (N_1603,N_1085,N_759);
and U1604 (N_1604,N_608,N_1093);
nand U1605 (N_1605,N_826,N_720);
or U1606 (N_1606,N_968,N_1199);
nor U1607 (N_1607,N_777,N_637);
and U1608 (N_1608,N_1047,N_683);
nor U1609 (N_1609,N_749,N_951);
and U1610 (N_1610,N_1192,N_683);
and U1611 (N_1611,N_935,N_902);
nand U1612 (N_1612,N_903,N_692);
and U1613 (N_1613,N_631,N_925);
nor U1614 (N_1614,N_845,N_1117);
and U1615 (N_1615,N_802,N_1030);
and U1616 (N_1616,N_732,N_866);
or U1617 (N_1617,N_893,N_823);
nor U1618 (N_1618,N_1188,N_1127);
nand U1619 (N_1619,N_732,N_1077);
and U1620 (N_1620,N_625,N_861);
nand U1621 (N_1621,N_956,N_812);
nor U1622 (N_1622,N_652,N_1115);
and U1623 (N_1623,N_1189,N_1117);
and U1624 (N_1624,N_765,N_864);
nor U1625 (N_1625,N_1148,N_818);
nor U1626 (N_1626,N_787,N_863);
nand U1627 (N_1627,N_690,N_847);
nand U1628 (N_1628,N_753,N_937);
nand U1629 (N_1629,N_647,N_874);
nor U1630 (N_1630,N_823,N_620);
nor U1631 (N_1631,N_1142,N_797);
nand U1632 (N_1632,N_1129,N_708);
nor U1633 (N_1633,N_767,N_604);
nor U1634 (N_1634,N_680,N_960);
and U1635 (N_1635,N_848,N_807);
and U1636 (N_1636,N_753,N_1052);
or U1637 (N_1637,N_1171,N_675);
nor U1638 (N_1638,N_801,N_900);
nand U1639 (N_1639,N_1067,N_1177);
nor U1640 (N_1640,N_774,N_807);
and U1641 (N_1641,N_1132,N_940);
nor U1642 (N_1642,N_799,N_1101);
and U1643 (N_1643,N_935,N_987);
nand U1644 (N_1644,N_1126,N_1061);
and U1645 (N_1645,N_1131,N_947);
nor U1646 (N_1646,N_986,N_869);
or U1647 (N_1647,N_959,N_971);
nand U1648 (N_1648,N_785,N_866);
nand U1649 (N_1649,N_707,N_1108);
and U1650 (N_1650,N_824,N_612);
nand U1651 (N_1651,N_1103,N_1012);
nor U1652 (N_1652,N_936,N_895);
nor U1653 (N_1653,N_1101,N_716);
and U1654 (N_1654,N_991,N_1168);
or U1655 (N_1655,N_767,N_786);
or U1656 (N_1656,N_608,N_1001);
nor U1657 (N_1657,N_765,N_860);
or U1658 (N_1658,N_1142,N_848);
or U1659 (N_1659,N_812,N_948);
nand U1660 (N_1660,N_607,N_1039);
xor U1661 (N_1661,N_948,N_877);
nand U1662 (N_1662,N_670,N_703);
or U1663 (N_1663,N_852,N_693);
nand U1664 (N_1664,N_789,N_865);
and U1665 (N_1665,N_612,N_822);
nor U1666 (N_1666,N_735,N_611);
nor U1667 (N_1667,N_639,N_1008);
nand U1668 (N_1668,N_896,N_859);
nor U1669 (N_1669,N_1198,N_1129);
or U1670 (N_1670,N_1097,N_621);
or U1671 (N_1671,N_635,N_1190);
or U1672 (N_1672,N_633,N_1122);
or U1673 (N_1673,N_974,N_729);
nand U1674 (N_1674,N_1063,N_689);
nand U1675 (N_1675,N_1129,N_958);
nor U1676 (N_1676,N_1088,N_696);
nor U1677 (N_1677,N_1040,N_978);
nor U1678 (N_1678,N_801,N_1123);
or U1679 (N_1679,N_880,N_1164);
or U1680 (N_1680,N_672,N_674);
nand U1681 (N_1681,N_959,N_1083);
and U1682 (N_1682,N_667,N_1165);
nor U1683 (N_1683,N_893,N_983);
nand U1684 (N_1684,N_695,N_660);
or U1685 (N_1685,N_840,N_954);
nand U1686 (N_1686,N_624,N_687);
nor U1687 (N_1687,N_1136,N_1199);
and U1688 (N_1688,N_1059,N_1148);
nor U1689 (N_1689,N_715,N_963);
and U1690 (N_1690,N_1079,N_1157);
nor U1691 (N_1691,N_1083,N_1148);
or U1692 (N_1692,N_813,N_912);
or U1693 (N_1693,N_1078,N_931);
nor U1694 (N_1694,N_1193,N_645);
and U1695 (N_1695,N_827,N_732);
nand U1696 (N_1696,N_1156,N_908);
or U1697 (N_1697,N_641,N_682);
nor U1698 (N_1698,N_1180,N_619);
or U1699 (N_1699,N_829,N_1136);
and U1700 (N_1700,N_664,N_1153);
and U1701 (N_1701,N_898,N_715);
and U1702 (N_1702,N_830,N_1097);
nor U1703 (N_1703,N_931,N_1016);
nor U1704 (N_1704,N_917,N_619);
and U1705 (N_1705,N_713,N_610);
nor U1706 (N_1706,N_706,N_849);
and U1707 (N_1707,N_1017,N_1123);
nor U1708 (N_1708,N_901,N_601);
nor U1709 (N_1709,N_1046,N_892);
nand U1710 (N_1710,N_905,N_699);
or U1711 (N_1711,N_650,N_725);
nor U1712 (N_1712,N_807,N_757);
or U1713 (N_1713,N_1110,N_854);
and U1714 (N_1714,N_653,N_658);
or U1715 (N_1715,N_697,N_701);
and U1716 (N_1716,N_1047,N_624);
or U1717 (N_1717,N_791,N_634);
and U1718 (N_1718,N_788,N_795);
or U1719 (N_1719,N_960,N_965);
nand U1720 (N_1720,N_954,N_1181);
nor U1721 (N_1721,N_607,N_833);
or U1722 (N_1722,N_1025,N_894);
nor U1723 (N_1723,N_953,N_940);
and U1724 (N_1724,N_915,N_624);
xor U1725 (N_1725,N_958,N_886);
nor U1726 (N_1726,N_774,N_1010);
nand U1727 (N_1727,N_682,N_971);
nand U1728 (N_1728,N_1167,N_995);
and U1729 (N_1729,N_678,N_916);
nand U1730 (N_1730,N_1014,N_1052);
and U1731 (N_1731,N_1174,N_813);
nand U1732 (N_1732,N_1079,N_956);
or U1733 (N_1733,N_944,N_701);
nand U1734 (N_1734,N_1101,N_1177);
and U1735 (N_1735,N_808,N_778);
or U1736 (N_1736,N_655,N_918);
xnor U1737 (N_1737,N_828,N_600);
and U1738 (N_1738,N_691,N_901);
or U1739 (N_1739,N_613,N_1086);
nand U1740 (N_1740,N_914,N_1190);
or U1741 (N_1741,N_685,N_1088);
or U1742 (N_1742,N_883,N_894);
or U1743 (N_1743,N_1137,N_956);
or U1744 (N_1744,N_1166,N_738);
or U1745 (N_1745,N_955,N_608);
nor U1746 (N_1746,N_947,N_859);
nand U1747 (N_1747,N_899,N_895);
or U1748 (N_1748,N_910,N_869);
nand U1749 (N_1749,N_1113,N_905);
nand U1750 (N_1750,N_1064,N_870);
nand U1751 (N_1751,N_1131,N_648);
or U1752 (N_1752,N_969,N_1084);
and U1753 (N_1753,N_680,N_922);
nand U1754 (N_1754,N_786,N_918);
and U1755 (N_1755,N_727,N_829);
or U1756 (N_1756,N_1026,N_671);
nor U1757 (N_1757,N_1055,N_682);
or U1758 (N_1758,N_1012,N_1065);
nor U1759 (N_1759,N_802,N_909);
nand U1760 (N_1760,N_958,N_676);
nor U1761 (N_1761,N_820,N_654);
and U1762 (N_1762,N_1167,N_1172);
nand U1763 (N_1763,N_1093,N_824);
nor U1764 (N_1764,N_662,N_1165);
and U1765 (N_1765,N_662,N_1101);
nand U1766 (N_1766,N_740,N_1060);
or U1767 (N_1767,N_690,N_1117);
nor U1768 (N_1768,N_695,N_1160);
and U1769 (N_1769,N_711,N_774);
or U1770 (N_1770,N_1173,N_869);
and U1771 (N_1771,N_905,N_1016);
and U1772 (N_1772,N_765,N_781);
nor U1773 (N_1773,N_1130,N_959);
or U1774 (N_1774,N_744,N_697);
and U1775 (N_1775,N_766,N_981);
nand U1776 (N_1776,N_1078,N_1088);
or U1777 (N_1777,N_856,N_1178);
and U1778 (N_1778,N_641,N_1010);
nand U1779 (N_1779,N_996,N_860);
and U1780 (N_1780,N_1118,N_810);
or U1781 (N_1781,N_950,N_737);
nand U1782 (N_1782,N_656,N_1175);
and U1783 (N_1783,N_962,N_608);
or U1784 (N_1784,N_1040,N_1000);
nand U1785 (N_1785,N_1026,N_1137);
or U1786 (N_1786,N_845,N_776);
nor U1787 (N_1787,N_1188,N_652);
xor U1788 (N_1788,N_848,N_1190);
or U1789 (N_1789,N_1035,N_632);
or U1790 (N_1790,N_712,N_776);
nand U1791 (N_1791,N_1196,N_739);
nor U1792 (N_1792,N_757,N_862);
nand U1793 (N_1793,N_881,N_1049);
nand U1794 (N_1794,N_614,N_927);
and U1795 (N_1795,N_736,N_867);
nand U1796 (N_1796,N_1134,N_919);
nor U1797 (N_1797,N_629,N_853);
nand U1798 (N_1798,N_1178,N_1099);
nand U1799 (N_1799,N_1017,N_1110);
and U1800 (N_1800,N_1473,N_1761);
and U1801 (N_1801,N_1360,N_1249);
or U1802 (N_1802,N_1621,N_1612);
and U1803 (N_1803,N_1518,N_1247);
nand U1804 (N_1804,N_1710,N_1379);
or U1805 (N_1805,N_1436,N_1289);
and U1806 (N_1806,N_1718,N_1276);
or U1807 (N_1807,N_1425,N_1726);
or U1808 (N_1808,N_1377,N_1534);
or U1809 (N_1809,N_1799,N_1245);
nor U1810 (N_1810,N_1508,N_1331);
nor U1811 (N_1811,N_1202,N_1638);
nand U1812 (N_1812,N_1560,N_1465);
nand U1813 (N_1813,N_1648,N_1305);
nand U1814 (N_1814,N_1227,N_1218);
or U1815 (N_1815,N_1502,N_1784);
or U1816 (N_1816,N_1579,N_1758);
and U1817 (N_1817,N_1330,N_1431);
and U1818 (N_1818,N_1443,N_1746);
or U1819 (N_1819,N_1216,N_1631);
nor U1820 (N_1820,N_1322,N_1386);
nand U1821 (N_1821,N_1597,N_1456);
or U1822 (N_1822,N_1676,N_1529);
nor U1823 (N_1823,N_1312,N_1258);
and U1824 (N_1824,N_1756,N_1513);
nor U1825 (N_1825,N_1624,N_1486);
or U1826 (N_1826,N_1757,N_1441);
and U1827 (N_1827,N_1266,N_1690);
and U1828 (N_1828,N_1482,N_1461);
and U1829 (N_1829,N_1393,N_1248);
and U1830 (N_1830,N_1319,N_1556);
nand U1831 (N_1831,N_1527,N_1469);
or U1832 (N_1832,N_1285,N_1582);
and U1833 (N_1833,N_1584,N_1222);
and U1834 (N_1834,N_1279,N_1596);
and U1835 (N_1835,N_1476,N_1740);
or U1836 (N_1836,N_1432,N_1449);
or U1837 (N_1837,N_1491,N_1576);
or U1838 (N_1838,N_1563,N_1338);
nor U1839 (N_1839,N_1774,N_1762);
or U1840 (N_1840,N_1419,N_1640);
nand U1841 (N_1841,N_1736,N_1547);
nor U1842 (N_1842,N_1472,N_1633);
or U1843 (N_1843,N_1646,N_1341);
or U1844 (N_1844,N_1274,N_1651);
nor U1845 (N_1845,N_1327,N_1385);
nor U1846 (N_1846,N_1735,N_1686);
and U1847 (N_1847,N_1376,N_1585);
nor U1848 (N_1848,N_1553,N_1670);
nand U1849 (N_1849,N_1378,N_1531);
or U1850 (N_1850,N_1308,N_1260);
or U1851 (N_1851,N_1742,N_1641);
nand U1852 (N_1852,N_1470,N_1437);
or U1853 (N_1853,N_1255,N_1243);
nand U1854 (N_1854,N_1201,N_1204);
nand U1855 (N_1855,N_1323,N_1694);
nand U1856 (N_1856,N_1734,N_1684);
nand U1857 (N_1857,N_1251,N_1480);
nor U1858 (N_1858,N_1667,N_1453);
or U1859 (N_1859,N_1280,N_1388);
xor U1860 (N_1860,N_1446,N_1399);
nor U1861 (N_1861,N_1656,N_1775);
and U1862 (N_1862,N_1776,N_1550);
nand U1863 (N_1863,N_1728,N_1615);
nor U1864 (N_1864,N_1233,N_1355);
and U1865 (N_1865,N_1221,N_1254);
and U1866 (N_1866,N_1496,N_1717);
or U1867 (N_1867,N_1600,N_1727);
or U1868 (N_1868,N_1619,N_1543);
or U1869 (N_1869,N_1760,N_1206);
nor U1870 (N_1870,N_1632,N_1752);
nor U1871 (N_1871,N_1366,N_1219);
nor U1872 (N_1872,N_1445,N_1643);
nor U1873 (N_1873,N_1235,N_1724);
nand U1874 (N_1874,N_1241,N_1603);
or U1875 (N_1875,N_1252,N_1711);
or U1876 (N_1876,N_1702,N_1297);
or U1877 (N_1877,N_1283,N_1662);
or U1878 (N_1878,N_1272,N_1680);
or U1879 (N_1879,N_1374,N_1382);
nor U1880 (N_1880,N_1215,N_1623);
and U1881 (N_1881,N_1304,N_1627);
or U1882 (N_1882,N_1709,N_1611);
nor U1883 (N_1883,N_1575,N_1787);
nand U1884 (N_1884,N_1701,N_1411);
and U1885 (N_1885,N_1413,N_1505);
nand U1886 (N_1886,N_1715,N_1238);
nand U1887 (N_1887,N_1592,N_1363);
xor U1888 (N_1888,N_1609,N_1636);
nand U1889 (N_1889,N_1677,N_1339);
nand U1890 (N_1890,N_1301,N_1739);
nand U1891 (N_1891,N_1687,N_1681);
or U1892 (N_1892,N_1217,N_1792);
nand U1893 (N_1893,N_1314,N_1264);
nor U1894 (N_1894,N_1708,N_1796);
nand U1895 (N_1895,N_1653,N_1299);
or U1896 (N_1896,N_1691,N_1412);
nor U1897 (N_1897,N_1454,N_1771);
or U1898 (N_1898,N_1464,N_1337);
nor U1899 (N_1899,N_1240,N_1346);
nor U1900 (N_1900,N_1253,N_1294);
or U1901 (N_1901,N_1610,N_1566);
nor U1902 (N_1902,N_1523,N_1741);
and U1903 (N_1903,N_1683,N_1259);
or U1904 (N_1904,N_1537,N_1540);
nor U1905 (N_1905,N_1481,N_1703);
or U1906 (N_1906,N_1407,N_1270);
nor U1907 (N_1907,N_1554,N_1356);
and U1908 (N_1908,N_1414,N_1406);
nand U1909 (N_1909,N_1391,N_1786);
and U1910 (N_1910,N_1390,N_1451);
nand U1911 (N_1911,N_1364,N_1521);
or U1912 (N_1912,N_1422,N_1466);
nand U1913 (N_1913,N_1781,N_1581);
and U1914 (N_1914,N_1350,N_1665);
nor U1915 (N_1915,N_1755,N_1688);
or U1916 (N_1916,N_1321,N_1606);
nor U1917 (N_1917,N_1557,N_1444);
nor U1918 (N_1918,N_1599,N_1284);
nor U1919 (N_1919,N_1616,N_1777);
and U1920 (N_1920,N_1532,N_1309);
and U1921 (N_1921,N_1380,N_1569);
and U1922 (N_1922,N_1660,N_1595);
or U1923 (N_1923,N_1555,N_1438);
or U1924 (N_1924,N_1524,N_1403);
or U1925 (N_1925,N_1797,N_1239);
or U1926 (N_1926,N_1509,N_1507);
nand U1927 (N_1927,N_1737,N_1489);
nor U1928 (N_1928,N_1424,N_1261);
nand U1929 (N_1929,N_1561,N_1571);
or U1930 (N_1930,N_1562,N_1589);
or U1931 (N_1931,N_1712,N_1673);
or U1932 (N_1932,N_1598,N_1544);
nand U1933 (N_1933,N_1429,N_1310);
nand U1934 (N_1934,N_1345,N_1488);
nor U1935 (N_1935,N_1499,N_1504);
nor U1936 (N_1936,N_1546,N_1542);
nor U1937 (N_1937,N_1516,N_1352);
nand U1938 (N_1938,N_1371,N_1315);
nor U1939 (N_1939,N_1211,N_1333);
nor U1940 (N_1940,N_1675,N_1765);
nand U1941 (N_1941,N_1789,N_1394);
or U1942 (N_1942,N_1794,N_1793);
nand U1943 (N_1943,N_1520,N_1591);
nand U1944 (N_1944,N_1763,N_1649);
and U1945 (N_1945,N_1250,N_1244);
nand U1946 (N_1946,N_1617,N_1626);
or U1947 (N_1947,N_1428,N_1590);
nand U1948 (N_1948,N_1398,N_1286);
nor U1949 (N_1949,N_1427,N_1652);
or U1950 (N_1950,N_1313,N_1334);
or U1951 (N_1951,N_1408,N_1410);
and U1952 (N_1952,N_1630,N_1203);
xnor U1953 (N_1953,N_1722,N_1256);
and U1954 (N_1954,N_1290,N_1664);
and U1955 (N_1955,N_1316,N_1318);
or U1956 (N_1956,N_1493,N_1423);
or U1957 (N_1957,N_1522,N_1440);
nand U1958 (N_1958,N_1629,N_1383);
nor U1959 (N_1959,N_1705,N_1359);
nand U1960 (N_1960,N_1369,N_1528);
nand U1961 (N_1961,N_1679,N_1692);
nand U1962 (N_1962,N_1232,N_1200);
nor U1963 (N_1963,N_1373,N_1311);
or U1964 (N_1964,N_1209,N_1788);
nor U1965 (N_1965,N_1700,N_1699);
nor U1966 (N_1966,N_1666,N_1501);
and U1967 (N_1967,N_1568,N_1336);
or U1968 (N_1968,N_1298,N_1678);
nand U1969 (N_1969,N_1668,N_1753);
nand U1970 (N_1970,N_1577,N_1574);
and U1971 (N_1971,N_1320,N_1275);
nand U1972 (N_1972,N_1426,N_1292);
nor U1973 (N_1973,N_1401,N_1271);
nand U1974 (N_1974,N_1262,N_1778);
and U1975 (N_1975,N_1220,N_1353);
and U1976 (N_1976,N_1479,N_1452);
or U1977 (N_1977,N_1706,N_1430);
nand U1978 (N_1978,N_1358,N_1485);
or U1979 (N_1979,N_1541,N_1759);
nand U1980 (N_1980,N_1417,N_1693);
and U1981 (N_1981,N_1392,N_1580);
nor U1982 (N_1982,N_1354,N_1768);
xnor U1983 (N_1983,N_1368,N_1697);
or U1984 (N_1984,N_1303,N_1395);
and U1985 (N_1985,N_1512,N_1224);
and U1986 (N_1986,N_1267,N_1492);
or U1987 (N_1987,N_1347,N_1389);
nor U1988 (N_1988,N_1287,N_1572);
nor U1989 (N_1989,N_1340,N_1498);
nand U1990 (N_1990,N_1367,N_1223);
or U1991 (N_1991,N_1608,N_1536);
xor U1992 (N_1992,N_1418,N_1764);
and U1993 (N_1993,N_1291,N_1559);
and U1994 (N_1994,N_1548,N_1647);
nand U1995 (N_1995,N_1663,N_1442);
nand U1996 (N_1996,N_1510,N_1295);
nand U1997 (N_1997,N_1332,N_1745);
and U1998 (N_1998,N_1767,N_1689);
and U1999 (N_1999,N_1421,N_1685);
and U2000 (N_2000,N_1387,N_1361);
nor U2001 (N_2001,N_1733,N_1351);
nand U2002 (N_2002,N_1458,N_1342);
and U2003 (N_2003,N_1234,N_1533);
or U2004 (N_2004,N_1655,N_1783);
or U2005 (N_2005,N_1230,N_1375);
nor U2006 (N_2006,N_1748,N_1578);
nor U2007 (N_2007,N_1798,N_1357);
or U2008 (N_2008,N_1785,N_1511);
nor U2009 (N_2009,N_1729,N_1293);
or U2010 (N_2010,N_1503,N_1669);
nor U2011 (N_2011,N_1645,N_1618);
nor U2012 (N_2012,N_1642,N_1564);
and U2013 (N_2013,N_1459,N_1657);
nand U2014 (N_2014,N_1790,N_1658);
nand U2015 (N_2015,N_1519,N_1497);
and U2016 (N_2016,N_1720,N_1695);
nand U2017 (N_2017,N_1474,N_1780);
nand U2018 (N_2018,N_1738,N_1236);
or U2019 (N_2019,N_1749,N_1242);
nor U2020 (N_2020,N_1302,N_1732);
or U2021 (N_2021,N_1281,N_1719);
or U2022 (N_2022,N_1674,N_1634);
or U2023 (N_2023,N_1614,N_1343);
and U2024 (N_2024,N_1730,N_1770);
nor U2025 (N_2025,N_1751,N_1463);
nand U2026 (N_2026,N_1384,N_1484);
or U2027 (N_2027,N_1558,N_1593);
and U2028 (N_2028,N_1713,N_1226);
nand U2029 (N_2029,N_1644,N_1682);
nor U2030 (N_2030,N_1620,N_1362);
and U2031 (N_2031,N_1744,N_1604);
and U2032 (N_2032,N_1483,N_1628);
or U2033 (N_2033,N_1208,N_1471);
nor U2034 (N_2034,N_1766,N_1535);
nand U2035 (N_2035,N_1795,N_1525);
and U2036 (N_2036,N_1439,N_1317);
or U2037 (N_2037,N_1494,N_1213);
or U2038 (N_2038,N_1273,N_1716);
and U2039 (N_2039,N_1263,N_1434);
and U2040 (N_2040,N_1268,N_1467);
nand U2041 (N_2041,N_1468,N_1588);
or U2042 (N_2042,N_1607,N_1514);
nand U2043 (N_2043,N_1517,N_1601);
nand U2044 (N_2044,N_1420,N_1225);
or U2045 (N_2045,N_1307,N_1402);
or U2046 (N_2046,N_1475,N_1448);
and U2047 (N_2047,N_1754,N_1567);
and U2048 (N_2048,N_1613,N_1515);
nor U2049 (N_2049,N_1477,N_1573);
or U2050 (N_2050,N_1622,N_1278);
nand U2051 (N_2051,N_1328,N_1506);
nand U2052 (N_2052,N_1265,N_1725);
or U2053 (N_2053,N_1602,N_1282);
nand U2054 (N_2054,N_1329,N_1397);
or U2055 (N_2055,N_1791,N_1731);
nor U2056 (N_2056,N_1457,N_1450);
or U2057 (N_2057,N_1257,N_1625);
nand U2058 (N_2058,N_1381,N_1415);
nand U2059 (N_2059,N_1455,N_1594);
nand U2060 (N_2060,N_1661,N_1296);
or U2061 (N_2061,N_1269,N_1539);
nor U2062 (N_2062,N_1433,N_1409);
and U2063 (N_2063,N_1570,N_1698);
or U2064 (N_2064,N_1586,N_1587);
nand U2065 (N_2065,N_1372,N_1344);
nor U2066 (N_2066,N_1228,N_1779);
nand U2067 (N_2067,N_1635,N_1704);
or U2068 (N_2068,N_1743,N_1400);
nor U2069 (N_2069,N_1782,N_1335);
nor U2070 (N_2070,N_1769,N_1500);
or U2071 (N_2071,N_1723,N_1552);
or U2072 (N_2072,N_1495,N_1530);
or U2073 (N_2073,N_1288,N_1637);
nand U2074 (N_2074,N_1325,N_1549);
nor U2075 (N_2075,N_1306,N_1348);
and U2076 (N_2076,N_1229,N_1605);
nor U2077 (N_2077,N_1396,N_1707);
or U2078 (N_2078,N_1214,N_1696);
and U2079 (N_2079,N_1277,N_1639);
or U2080 (N_2080,N_1672,N_1654);
nand U2081 (N_2081,N_1551,N_1205);
nand U2082 (N_2082,N_1404,N_1671);
and U2083 (N_2083,N_1650,N_1207);
nand U2084 (N_2084,N_1462,N_1750);
nor U2085 (N_2085,N_1231,N_1460);
or U2086 (N_2086,N_1212,N_1773);
and U2087 (N_2087,N_1324,N_1714);
and U2088 (N_2088,N_1447,N_1300);
or U2089 (N_2089,N_1435,N_1747);
or U2090 (N_2090,N_1538,N_1405);
and U2091 (N_2091,N_1526,N_1583);
or U2092 (N_2092,N_1772,N_1326);
or U2093 (N_2093,N_1210,N_1365);
and U2094 (N_2094,N_1490,N_1545);
nor U2095 (N_2095,N_1478,N_1349);
and U2096 (N_2096,N_1721,N_1565);
nor U2097 (N_2097,N_1416,N_1370);
nand U2098 (N_2098,N_1246,N_1237);
nand U2099 (N_2099,N_1659,N_1487);
or U2100 (N_2100,N_1583,N_1263);
nand U2101 (N_2101,N_1637,N_1238);
nor U2102 (N_2102,N_1574,N_1582);
and U2103 (N_2103,N_1703,N_1327);
nor U2104 (N_2104,N_1205,N_1358);
nor U2105 (N_2105,N_1552,N_1331);
nor U2106 (N_2106,N_1272,N_1775);
or U2107 (N_2107,N_1580,N_1583);
nor U2108 (N_2108,N_1788,N_1794);
or U2109 (N_2109,N_1664,N_1570);
nor U2110 (N_2110,N_1675,N_1334);
or U2111 (N_2111,N_1655,N_1528);
or U2112 (N_2112,N_1607,N_1393);
or U2113 (N_2113,N_1323,N_1796);
nor U2114 (N_2114,N_1298,N_1325);
nand U2115 (N_2115,N_1519,N_1779);
nand U2116 (N_2116,N_1465,N_1237);
or U2117 (N_2117,N_1622,N_1220);
and U2118 (N_2118,N_1455,N_1457);
or U2119 (N_2119,N_1448,N_1616);
nand U2120 (N_2120,N_1475,N_1599);
nand U2121 (N_2121,N_1383,N_1418);
or U2122 (N_2122,N_1292,N_1433);
nor U2123 (N_2123,N_1305,N_1510);
xnor U2124 (N_2124,N_1411,N_1372);
nand U2125 (N_2125,N_1238,N_1770);
or U2126 (N_2126,N_1629,N_1422);
or U2127 (N_2127,N_1636,N_1611);
nand U2128 (N_2128,N_1459,N_1317);
nand U2129 (N_2129,N_1712,N_1440);
nand U2130 (N_2130,N_1530,N_1437);
or U2131 (N_2131,N_1750,N_1517);
or U2132 (N_2132,N_1638,N_1354);
nand U2133 (N_2133,N_1790,N_1650);
nor U2134 (N_2134,N_1553,N_1596);
nor U2135 (N_2135,N_1575,N_1274);
or U2136 (N_2136,N_1491,N_1684);
nand U2137 (N_2137,N_1550,N_1636);
nor U2138 (N_2138,N_1460,N_1238);
and U2139 (N_2139,N_1559,N_1728);
nor U2140 (N_2140,N_1417,N_1776);
nand U2141 (N_2141,N_1364,N_1516);
nand U2142 (N_2142,N_1215,N_1784);
nor U2143 (N_2143,N_1250,N_1653);
or U2144 (N_2144,N_1647,N_1499);
and U2145 (N_2145,N_1535,N_1557);
nand U2146 (N_2146,N_1635,N_1615);
or U2147 (N_2147,N_1515,N_1285);
nor U2148 (N_2148,N_1724,N_1638);
nor U2149 (N_2149,N_1510,N_1738);
or U2150 (N_2150,N_1411,N_1447);
and U2151 (N_2151,N_1715,N_1408);
nor U2152 (N_2152,N_1532,N_1764);
or U2153 (N_2153,N_1720,N_1334);
nand U2154 (N_2154,N_1794,N_1543);
nand U2155 (N_2155,N_1749,N_1446);
nand U2156 (N_2156,N_1342,N_1542);
or U2157 (N_2157,N_1676,N_1476);
and U2158 (N_2158,N_1400,N_1413);
and U2159 (N_2159,N_1736,N_1520);
nor U2160 (N_2160,N_1622,N_1459);
nand U2161 (N_2161,N_1569,N_1611);
nand U2162 (N_2162,N_1250,N_1511);
and U2163 (N_2163,N_1746,N_1423);
and U2164 (N_2164,N_1723,N_1414);
nand U2165 (N_2165,N_1306,N_1432);
and U2166 (N_2166,N_1719,N_1775);
and U2167 (N_2167,N_1402,N_1628);
nand U2168 (N_2168,N_1668,N_1796);
or U2169 (N_2169,N_1711,N_1427);
or U2170 (N_2170,N_1384,N_1628);
nand U2171 (N_2171,N_1291,N_1512);
and U2172 (N_2172,N_1659,N_1517);
and U2173 (N_2173,N_1600,N_1288);
and U2174 (N_2174,N_1280,N_1714);
nand U2175 (N_2175,N_1233,N_1648);
and U2176 (N_2176,N_1702,N_1442);
and U2177 (N_2177,N_1725,N_1665);
and U2178 (N_2178,N_1568,N_1766);
and U2179 (N_2179,N_1352,N_1296);
nand U2180 (N_2180,N_1347,N_1267);
nand U2181 (N_2181,N_1276,N_1677);
or U2182 (N_2182,N_1701,N_1755);
and U2183 (N_2183,N_1419,N_1527);
nor U2184 (N_2184,N_1749,N_1532);
nor U2185 (N_2185,N_1255,N_1679);
nor U2186 (N_2186,N_1251,N_1685);
and U2187 (N_2187,N_1546,N_1627);
nor U2188 (N_2188,N_1402,N_1361);
and U2189 (N_2189,N_1387,N_1663);
or U2190 (N_2190,N_1469,N_1258);
and U2191 (N_2191,N_1490,N_1281);
and U2192 (N_2192,N_1635,N_1478);
nor U2193 (N_2193,N_1538,N_1441);
nand U2194 (N_2194,N_1283,N_1333);
or U2195 (N_2195,N_1277,N_1629);
and U2196 (N_2196,N_1428,N_1703);
or U2197 (N_2197,N_1560,N_1352);
and U2198 (N_2198,N_1318,N_1627);
nor U2199 (N_2199,N_1422,N_1500);
or U2200 (N_2200,N_1273,N_1676);
nor U2201 (N_2201,N_1541,N_1767);
or U2202 (N_2202,N_1429,N_1794);
or U2203 (N_2203,N_1557,N_1378);
and U2204 (N_2204,N_1793,N_1752);
nand U2205 (N_2205,N_1656,N_1447);
nor U2206 (N_2206,N_1316,N_1705);
or U2207 (N_2207,N_1698,N_1507);
and U2208 (N_2208,N_1224,N_1230);
and U2209 (N_2209,N_1291,N_1642);
or U2210 (N_2210,N_1357,N_1743);
nand U2211 (N_2211,N_1588,N_1704);
and U2212 (N_2212,N_1419,N_1261);
nor U2213 (N_2213,N_1388,N_1677);
nor U2214 (N_2214,N_1421,N_1447);
or U2215 (N_2215,N_1593,N_1680);
nor U2216 (N_2216,N_1262,N_1728);
or U2217 (N_2217,N_1387,N_1776);
and U2218 (N_2218,N_1736,N_1581);
and U2219 (N_2219,N_1504,N_1267);
nand U2220 (N_2220,N_1690,N_1660);
and U2221 (N_2221,N_1632,N_1559);
or U2222 (N_2222,N_1706,N_1654);
and U2223 (N_2223,N_1516,N_1224);
nor U2224 (N_2224,N_1553,N_1202);
or U2225 (N_2225,N_1726,N_1713);
or U2226 (N_2226,N_1589,N_1645);
or U2227 (N_2227,N_1533,N_1318);
nand U2228 (N_2228,N_1619,N_1644);
nor U2229 (N_2229,N_1582,N_1532);
nor U2230 (N_2230,N_1435,N_1336);
xnor U2231 (N_2231,N_1614,N_1676);
and U2232 (N_2232,N_1346,N_1693);
nand U2233 (N_2233,N_1566,N_1283);
or U2234 (N_2234,N_1652,N_1417);
nor U2235 (N_2235,N_1246,N_1278);
and U2236 (N_2236,N_1362,N_1257);
or U2237 (N_2237,N_1763,N_1603);
nand U2238 (N_2238,N_1477,N_1405);
and U2239 (N_2239,N_1648,N_1755);
nand U2240 (N_2240,N_1650,N_1590);
or U2241 (N_2241,N_1520,N_1387);
or U2242 (N_2242,N_1580,N_1712);
and U2243 (N_2243,N_1657,N_1736);
nand U2244 (N_2244,N_1316,N_1520);
or U2245 (N_2245,N_1456,N_1487);
nand U2246 (N_2246,N_1239,N_1688);
nand U2247 (N_2247,N_1356,N_1694);
nand U2248 (N_2248,N_1508,N_1212);
nor U2249 (N_2249,N_1603,N_1498);
nand U2250 (N_2250,N_1729,N_1460);
or U2251 (N_2251,N_1309,N_1543);
nand U2252 (N_2252,N_1396,N_1655);
and U2253 (N_2253,N_1390,N_1376);
nand U2254 (N_2254,N_1387,N_1381);
xnor U2255 (N_2255,N_1381,N_1762);
or U2256 (N_2256,N_1796,N_1494);
and U2257 (N_2257,N_1568,N_1246);
and U2258 (N_2258,N_1757,N_1655);
nor U2259 (N_2259,N_1787,N_1784);
and U2260 (N_2260,N_1729,N_1581);
or U2261 (N_2261,N_1353,N_1341);
nand U2262 (N_2262,N_1200,N_1576);
nor U2263 (N_2263,N_1358,N_1263);
nand U2264 (N_2264,N_1228,N_1203);
and U2265 (N_2265,N_1575,N_1606);
nand U2266 (N_2266,N_1275,N_1460);
or U2267 (N_2267,N_1718,N_1302);
nor U2268 (N_2268,N_1404,N_1702);
nor U2269 (N_2269,N_1770,N_1353);
and U2270 (N_2270,N_1466,N_1583);
and U2271 (N_2271,N_1673,N_1660);
nor U2272 (N_2272,N_1281,N_1220);
nor U2273 (N_2273,N_1230,N_1500);
nand U2274 (N_2274,N_1462,N_1788);
nor U2275 (N_2275,N_1449,N_1207);
or U2276 (N_2276,N_1488,N_1238);
nand U2277 (N_2277,N_1565,N_1728);
nor U2278 (N_2278,N_1212,N_1618);
or U2279 (N_2279,N_1521,N_1514);
nor U2280 (N_2280,N_1660,N_1496);
or U2281 (N_2281,N_1344,N_1205);
nand U2282 (N_2282,N_1221,N_1750);
and U2283 (N_2283,N_1565,N_1791);
or U2284 (N_2284,N_1588,N_1732);
and U2285 (N_2285,N_1743,N_1279);
nor U2286 (N_2286,N_1750,N_1412);
nand U2287 (N_2287,N_1353,N_1284);
xnor U2288 (N_2288,N_1354,N_1750);
or U2289 (N_2289,N_1384,N_1673);
nand U2290 (N_2290,N_1247,N_1595);
nor U2291 (N_2291,N_1233,N_1568);
nor U2292 (N_2292,N_1624,N_1211);
nand U2293 (N_2293,N_1402,N_1632);
nor U2294 (N_2294,N_1253,N_1218);
and U2295 (N_2295,N_1737,N_1788);
nand U2296 (N_2296,N_1598,N_1488);
or U2297 (N_2297,N_1308,N_1330);
nor U2298 (N_2298,N_1295,N_1670);
nand U2299 (N_2299,N_1291,N_1292);
nand U2300 (N_2300,N_1718,N_1298);
and U2301 (N_2301,N_1573,N_1225);
nand U2302 (N_2302,N_1521,N_1519);
nand U2303 (N_2303,N_1610,N_1379);
nor U2304 (N_2304,N_1534,N_1743);
nand U2305 (N_2305,N_1707,N_1323);
and U2306 (N_2306,N_1513,N_1414);
or U2307 (N_2307,N_1738,N_1200);
nor U2308 (N_2308,N_1417,N_1339);
or U2309 (N_2309,N_1655,N_1479);
or U2310 (N_2310,N_1205,N_1585);
nand U2311 (N_2311,N_1739,N_1519);
nand U2312 (N_2312,N_1703,N_1475);
and U2313 (N_2313,N_1797,N_1719);
or U2314 (N_2314,N_1449,N_1297);
nor U2315 (N_2315,N_1753,N_1422);
and U2316 (N_2316,N_1699,N_1313);
and U2317 (N_2317,N_1445,N_1319);
nand U2318 (N_2318,N_1591,N_1408);
nand U2319 (N_2319,N_1337,N_1768);
or U2320 (N_2320,N_1531,N_1399);
nor U2321 (N_2321,N_1567,N_1650);
and U2322 (N_2322,N_1274,N_1582);
or U2323 (N_2323,N_1317,N_1268);
nor U2324 (N_2324,N_1274,N_1414);
and U2325 (N_2325,N_1717,N_1642);
nor U2326 (N_2326,N_1527,N_1355);
or U2327 (N_2327,N_1381,N_1202);
nor U2328 (N_2328,N_1740,N_1372);
or U2329 (N_2329,N_1485,N_1296);
nand U2330 (N_2330,N_1531,N_1551);
nor U2331 (N_2331,N_1446,N_1553);
nor U2332 (N_2332,N_1380,N_1551);
nand U2333 (N_2333,N_1543,N_1496);
nand U2334 (N_2334,N_1212,N_1208);
and U2335 (N_2335,N_1486,N_1269);
and U2336 (N_2336,N_1545,N_1783);
nand U2337 (N_2337,N_1663,N_1441);
nor U2338 (N_2338,N_1781,N_1330);
nand U2339 (N_2339,N_1646,N_1308);
or U2340 (N_2340,N_1444,N_1689);
nand U2341 (N_2341,N_1367,N_1570);
nor U2342 (N_2342,N_1658,N_1510);
nor U2343 (N_2343,N_1657,N_1500);
nor U2344 (N_2344,N_1665,N_1289);
nor U2345 (N_2345,N_1599,N_1254);
nand U2346 (N_2346,N_1463,N_1312);
nor U2347 (N_2347,N_1578,N_1502);
nor U2348 (N_2348,N_1608,N_1386);
nand U2349 (N_2349,N_1399,N_1655);
nor U2350 (N_2350,N_1373,N_1680);
and U2351 (N_2351,N_1482,N_1542);
and U2352 (N_2352,N_1342,N_1548);
nor U2353 (N_2353,N_1650,N_1315);
and U2354 (N_2354,N_1590,N_1673);
nor U2355 (N_2355,N_1291,N_1306);
or U2356 (N_2356,N_1799,N_1791);
nor U2357 (N_2357,N_1521,N_1376);
and U2358 (N_2358,N_1716,N_1771);
nand U2359 (N_2359,N_1699,N_1354);
nor U2360 (N_2360,N_1538,N_1768);
or U2361 (N_2361,N_1741,N_1724);
nor U2362 (N_2362,N_1349,N_1714);
and U2363 (N_2363,N_1278,N_1289);
and U2364 (N_2364,N_1544,N_1580);
or U2365 (N_2365,N_1505,N_1699);
or U2366 (N_2366,N_1325,N_1247);
nand U2367 (N_2367,N_1557,N_1511);
or U2368 (N_2368,N_1333,N_1747);
or U2369 (N_2369,N_1585,N_1538);
nor U2370 (N_2370,N_1272,N_1704);
nand U2371 (N_2371,N_1397,N_1316);
nand U2372 (N_2372,N_1267,N_1200);
and U2373 (N_2373,N_1320,N_1220);
and U2374 (N_2374,N_1407,N_1244);
and U2375 (N_2375,N_1206,N_1268);
nand U2376 (N_2376,N_1653,N_1607);
nand U2377 (N_2377,N_1314,N_1382);
nor U2378 (N_2378,N_1274,N_1772);
nand U2379 (N_2379,N_1588,N_1496);
and U2380 (N_2380,N_1595,N_1222);
nand U2381 (N_2381,N_1465,N_1407);
or U2382 (N_2382,N_1569,N_1680);
nor U2383 (N_2383,N_1666,N_1675);
or U2384 (N_2384,N_1622,N_1766);
or U2385 (N_2385,N_1429,N_1280);
and U2386 (N_2386,N_1753,N_1363);
or U2387 (N_2387,N_1494,N_1498);
nor U2388 (N_2388,N_1293,N_1610);
or U2389 (N_2389,N_1364,N_1248);
or U2390 (N_2390,N_1300,N_1594);
and U2391 (N_2391,N_1313,N_1246);
nor U2392 (N_2392,N_1204,N_1629);
or U2393 (N_2393,N_1492,N_1408);
nand U2394 (N_2394,N_1266,N_1646);
and U2395 (N_2395,N_1659,N_1316);
nand U2396 (N_2396,N_1787,N_1202);
nor U2397 (N_2397,N_1374,N_1682);
or U2398 (N_2398,N_1660,N_1333);
and U2399 (N_2399,N_1551,N_1235);
or U2400 (N_2400,N_2088,N_2111);
nand U2401 (N_2401,N_1921,N_2086);
nand U2402 (N_2402,N_2181,N_2003);
nand U2403 (N_2403,N_2265,N_1899);
and U2404 (N_2404,N_2136,N_2192);
nand U2405 (N_2405,N_2205,N_1855);
nand U2406 (N_2406,N_2150,N_1963);
nand U2407 (N_2407,N_1902,N_1852);
and U2408 (N_2408,N_2305,N_2124);
nor U2409 (N_2409,N_2399,N_2174);
and U2410 (N_2410,N_1823,N_2023);
nor U2411 (N_2411,N_2197,N_2266);
and U2412 (N_2412,N_2047,N_1976);
or U2413 (N_2413,N_1888,N_2084);
nor U2414 (N_2414,N_2015,N_2147);
nor U2415 (N_2415,N_1811,N_1965);
nor U2416 (N_2416,N_2291,N_1885);
and U2417 (N_2417,N_2384,N_1996);
nand U2418 (N_2418,N_1840,N_2229);
nand U2419 (N_2419,N_2210,N_2326);
nand U2420 (N_2420,N_2089,N_1817);
nor U2421 (N_2421,N_2158,N_2020);
nand U2422 (N_2422,N_1898,N_2043);
nand U2423 (N_2423,N_1914,N_2321);
nor U2424 (N_2424,N_1828,N_2100);
and U2425 (N_2425,N_1826,N_2264);
or U2426 (N_2426,N_2354,N_2040);
nor U2427 (N_2427,N_1931,N_2137);
nand U2428 (N_2428,N_2090,N_1911);
and U2429 (N_2429,N_2002,N_1954);
nand U2430 (N_2430,N_2268,N_1889);
nor U2431 (N_2431,N_2159,N_2302);
nor U2432 (N_2432,N_2343,N_2118);
nand U2433 (N_2433,N_2218,N_2144);
and U2434 (N_2434,N_2281,N_1867);
or U2435 (N_2435,N_2350,N_1932);
nand U2436 (N_2436,N_2065,N_2240);
and U2437 (N_2437,N_2132,N_2295);
and U2438 (N_2438,N_2012,N_2358);
and U2439 (N_2439,N_2226,N_1829);
or U2440 (N_2440,N_1930,N_2119);
nor U2441 (N_2441,N_2194,N_2336);
xnor U2442 (N_2442,N_2180,N_1944);
nand U2443 (N_2443,N_2106,N_2287);
nor U2444 (N_2444,N_2101,N_2289);
nor U2445 (N_2445,N_2203,N_2075);
or U2446 (N_2446,N_2293,N_2365);
xor U2447 (N_2447,N_2056,N_2338);
nand U2448 (N_2448,N_2004,N_1915);
or U2449 (N_2449,N_2055,N_2367);
nand U2450 (N_2450,N_1979,N_2374);
or U2451 (N_2451,N_2379,N_2083);
nand U2452 (N_2452,N_2102,N_2298);
nand U2453 (N_2453,N_2247,N_1992);
nand U2454 (N_2454,N_2269,N_1919);
or U2455 (N_2455,N_1928,N_2335);
nand U2456 (N_2456,N_2370,N_2064);
nand U2457 (N_2457,N_1864,N_2311);
or U2458 (N_2458,N_2233,N_2307);
nor U2459 (N_2459,N_2183,N_1977);
or U2460 (N_2460,N_2388,N_2241);
or U2461 (N_2461,N_2087,N_2373);
and U2462 (N_2462,N_1830,N_2392);
and U2463 (N_2463,N_2317,N_2188);
nand U2464 (N_2464,N_2208,N_2245);
nand U2465 (N_2465,N_2278,N_2034);
or U2466 (N_2466,N_2185,N_2273);
nor U2467 (N_2467,N_1981,N_2117);
and U2468 (N_2468,N_2364,N_1883);
or U2469 (N_2469,N_2267,N_2073);
nor U2470 (N_2470,N_1809,N_2103);
nand U2471 (N_2471,N_1842,N_2257);
or U2472 (N_2472,N_2025,N_2391);
nor U2473 (N_2473,N_1958,N_2169);
and U2474 (N_2474,N_2098,N_2186);
and U2475 (N_2475,N_2272,N_2067);
or U2476 (N_2476,N_2104,N_1832);
or U2477 (N_2477,N_2189,N_2363);
nand U2478 (N_2478,N_2076,N_2062);
and U2479 (N_2479,N_1938,N_2096);
nor U2480 (N_2480,N_2386,N_2351);
or U2481 (N_2481,N_2313,N_1892);
or U2482 (N_2482,N_2014,N_2161);
and U2483 (N_2483,N_2061,N_2206);
nand U2484 (N_2484,N_1815,N_1967);
nand U2485 (N_2485,N_2275,N_2110);
nor U2486 (N_2486,N_1939,N_2165);
nor U2487 (N_2487,N_1808,N_2377);
nor U2488 (N_2488,N_2258,N_2286);
and U2489 (N_2489,N_2044,N_1982);
nor U2490 (N_2490,N_2116,N_2079);
nand U2491 (N_2491,N_2195,N_1917);
and U2492 (N_2492,N_2091,N_2152);
or U2493 (N_2493,N_2122,N_2228);
or U2494 (N_2494,N_1973,N_1875);
or U2495 (N_2495,N_2348,N_2344);
or U2496 (N_2496,N_1833,N_2382);
or U2497 (N_2497,N_2304,N_2243);
nand U2498 (N_2498,N_1847,N_2239);
nand U2499 (N_2499,N_2332,N_1908);
or U2500 (N_2500,N_1945,N_1886);
nand U2501 (N_2501,N_2109,N_1904);
or U2502 (N_2502,N_2177,N_2138);
nor U2503 (N_2503,N_2139,N_1821);
nand U2504 (N_2504,N_2296,N_2080);
nand U2505 (N_2505,N_1856,N_1959);
and U2506 (N_2506,N_2389,N_2204);
nand U2507 (N_2507,N_2325,N_1952);
nand U2508 (N_2508,N_2074,N_2066);
and U2509 (N_2509,N_1844,N_1937);
or U2510 (N_2510,N_1946,N_2309);
nor U2511 (N_2511,N_2097,N_2166);
and U2512 (N_2512,N_1819,N_2261);
nor U2513 (N_2513,N_1870,N_2316);
and U2514 (N_2514,N_2054,N_1858);
or U2515 (N_2515,N_2320,N_2360);
or U2516 (N_2516,N_2323,N_2176);
nand U2517 (N_2517,N_2340,N_2346);
and U2518 (N_2518,N_2143,N_2246);
and U2519 (N_2519,N_2153,N_2366);
or U2520 (N_2520,N_2170,N_2256);
and U2521 (N_2521,N_2394,N_2230);
and U2522 (N_2522,N_2253,N_1906);
or U2523 (N_2523,N_1956,N_1934);
nand U2524 (N_2524,N_1922,N_2000);
or U2525 (N_2525,N_2115,N_1860);
and U2526 (N_2526,N_1834,N_1803);
and U2527 (N_2527,N_2198,N_2049);
nand U2528 (N_2528,N_2237,N_1940);
or U2529 (N_2529,N_2085,N_1800);
or U2530 (N_2530,N_2050,N_2045);
or U2531 (N_2531,N_1929,N_2251);
nor U2532 (N_2532,N_2133,N_1814);
nand U2533 (N_2533,N_2028,N_1975);
or U2534 (N_2534,N_2127,N_2215);
nor U2535 (N_2535,N_2331,N_2398);
nand U2536 (N_2536,N_2276,N_2008);
nor U2537 (N_2537,N_2190,N_2337);
and U2538 (N_2538,N_2285,N_2038);
or U2539 (N_2539,N_2068,N_2128);
or U2540 (N_2540,N_2007,N_1845);
nor U2541 (N_2541,N_2371,N_2224);
and U2542 (N_2542,N_2292,N_2125);
or U2543 (N_2543,N_2027,N_1894);
nand U2544 (N_2544,N_1960,N_2018);
and U2545 (N_2545,N_1943,N_1891);
and U2546 (N_2546,N_2310,N_2123);
or U2547 (N_2547,N_2312,N_2162);
nor U2548 (N_2548,N_1927,N_1801);
nor U2549 (N_2549,N_2319,N_2328);
or U2550 (N_2550,N_1951,N_1802);
or U2551 (N_2551,N_2383,N_2154);
nor U2552 (N_2552,N_1881,N_2283);
or U2553 (N_2553,N_2172,N_2010);
nand U2554 (N_2554,N_2157,N_2306);
or U2555 (N_2555,N_1972,N_2178);
nor U2556 (N_2556,N_2077,N_2236);
nor U2557 (N_2557,N_2220,N_2259);
and U2558 (N_2558,N_2013,N_1961);
nor U2559 (N_2559,N_1812,N_2042);
nand U2560 (N_2560,N_2284,N_1876);
and U2561 (N_2561,N_2372,N_2378);
nand U2562 (N_2562,N_2255,N_1920);
and U2563 (N_2563,N_1985,N_1918);
or U2564 (N_2564,N_2260,N_1869);
nand U2565 (N_2565,N_1807,N_2290);
and U2566 (N_2566,N_2209,N_1990);
or U2567 (N_2567,N_2072,N_1804);
or U2568 (N_2568,N_1962,N_2029);
and U2569 (N_2569,N_2242,N_2134);
nor U2570 (N_2570,N_1912,N_2095);
or U2571 (N_2571,N_2082,N_1936);
nand U2572 (N_2572,N_2271,N_1818);
nor U2573 (N_2573,N_2011,N_2222);
nor U2574 (N_2574,N_2288,N_1947);
and U2575 (N_2575,N_2359,N_2381);
nand U2576 (N_2576,N_2071,N_1993);
xnor U2577 (N_2577,N_1933,N_2022);
nand U2578 (N_2578,N_2216,N_2387);
nor U2579 (N_2579,N_1824,N_1838);
or U2580 (N_2580,N_2207,N_1942);
and U2581 (N_2581,N_2006,N_2175);
nor U2582 (N_2582,N_1949,N_1890);
nor U2583 (N_2583,N_2121,N_2249);
nor U2584 (N_2584,N_1953,N_2324);
nand U2585 (N_2585,N_1941,N_2353);
and U2586 (N_2586,N_2094,N_2130);
and U2587 (N_2587,N_2167,N_1836);
nand U2588 (N_2588,N_2303,N_2248);
or U2589 (N_2589,N_2390,N_2114);
nand U2590 (N_2590,N_1948,N_1879);
and U2591 (N_2591,N_2199,N_2164);
or U2592 (N_2592,N_1987,N_2395);
nor U2593 (N_2593,N_1997,N_1970);
nor U2594 (N_2594,N_2212,N_2300);
nor U2595 (N_2595,N_1900,N_1866);
and U2596 (N_2596,N_1896,N_2155);
nor U2597 (N_2597,N_1989,N_2282);
nor U2598 (N_2598,N_2252,N_1994);
nor U2599 (N_2599,N_2173,N_2182);
or U2600 (N_2600,N_1839,N_2030);
or U2601 (N_2601,N_1974,N_2297);
nor U2602 (N_2602,N_2019,N_2107);
and U2603 (N_2603,N_2235,N_2026);
or U2604 (N_2604,N_1983,N_1895);
nor U2605 (N_2605,N_1964,N_2238);
nand U2606 (N_2606,N_1810,N_1877);
nor U2607 (N_2607,N_2046,N_1913);
and U2608 (N_2608,N_1846,N_2279);
and U2609 (N_2609,N_2345,N_2223);
and U2610 (N_2610,N_2037,N_2201);
nand U2611 (N_2611,N_2039,N_1969);
nand U2612 (N_2612,N_2131,N_1859);
or U2613 (N_2613,N_1924,N_1978);
and U2614 (N_2614,N_2151,N_1980);
and U2615 (N_2615,N_1926,N_1995);
and U2616 (N_2616,N_2009,N_1887);
nor U2617 (N_2617,N_1882,N_2231);
nor U2618 (N_2618,N_1907,N_2070);
or U2619 (N_2619,N_1955,N_2191);
nor U2620 (N_2620,N_2254,N_2032);
nor U2621 (N_2621,N_2021,N_2168);
and U2622 (N_2622,N_2219,N_1835);
and U2623 (N_2623,N_1820,N_1903);
nor U2624 (N_2624,N_2179,N_1998);
or U2625 (N_2625,N_2017,N_1878);
or U2626 (N_2626,N_1909,N_1923);
nor U2627 (N_2627,N_2160,N_1905);
or U2628 (N_2628,N_2385,N_1853);
and U2629 (N_2629,N_2299,N_2202);
or U2630 (N_2630,N_2211,N_1849);
or U2631 (N_2631,N_1966,N_2035);
nand U2632 (N_2632,N_2016,N_2361);
nand U2633 (N_2633,N_1851,N_1897);
nor U2634 (N_2634,N_1857,N_2057);
or U2635 (N_2635,N_2156,N_1813);
nand U2636 (N_2636,N_2263,N_2187);
nor U2637 (N_2637,N_2052,N_2397);
and U2638 (N_2638,N_2051,N_2196);
and U2639 (N_2639,N_2357,N_1806);
or U2640 (N_2640,N_2396,N_2314);
and U2641 (N_2641,N_2274,N_2141);
nor U2642 (N_2642,N_2327,N_2033);
and U2643 (N_2643,N_2301,N_2200);
and U2644 (N_2644,N_1862,N_2149);
and U2645 (N_2645,N_2308,N_1925);
nor U2646 (N_2646,N_2333,N_1893);
nand U2647 (N_2647,N_2081,N_2380);
nor U2648 (N_2648,N_2213,N_1901);
or U2649 (N_2649,N_2214,N_2092);
nor U2650 (N_2650,N_1827,N_1863);
nand U2651 (N_2651,N_2112,N_1999);
or U2652 (N_2652,N_2330,N_2135);
and U2653 (N_2653,N_2146,N_2318);
or U2654 (N_2654,N_1872,N_1873);
and U2655 (N_2655,N_2093,N_2145);
or U2656 (N_2656,N_2355,N_2069);
and U2657 (N_2657,N_1971,N_1854);
or U2658 (N_2658,N_2234,N_2329);
nor U2659 (N_2659,N_1837,N_2041);
nand U2660 (N_2660,N_2232,N_1822);
nand U2661 (N_2661,N_1916,N_2105);
and U2662 (N_2662,N_2250,N_1871);
and U2663 (N_2663,N_2048,N_2053);
or U2664 (N_2664,N_2334,N_2060);
nand U2665 (N_2665,N_2163,N_2113);
and U2666 (N_2666,N_2368,N_2078);
and U2667 (N_2667,N_1988,N_1841);
xor U2668 (N_2668,N_1861,N_2315);
nand U2669 (N_2669,N_2217,N_1910);
or U2670 (N_2670,N_2005,N_2294);
nand U2671 (N_2671,N_2129,N_2262);
and U2672 (N_2672,N_2036,N_2184);
nor U2673 (N_2673,N_2342,N_1968);
and U2674 (N_2674,N_1935,N_2225);
nand U2675 (N_2675,N_1957,N_2352);
xnor U2676 (N_2676,N_1831,N_1816);
or U2677 (N_2677,N_2322,N_2063);
and U2678 (N_2678,N_2059,N_2280);
nand U2679 (N_2679,N_1986,N_2171);
or U2680 (N_2680,N_1848,N_1874);
and U2681 (N_2681,N_2277,N_2120);
or U2682 (N_2682,N_2339,N_2193);
or U2683 (N_2683,N_2108,N_2142);
nand U2684 (N_2684,N_2001,N_1805);
or U2685 (N_2685,N_1880,N_2140);
nand U2686 (N_2686,N_2347,N_2393);
nand U2687 (N_2687,N_1950,N_1865);
or U2688 (N_2688,N_1843,N_1868);
and U2689 (N_2689,N_2227,N_2024);
nor U2690 (N_2690,N_2356,N_1884);
or U2691 (N_2691,N_2369,N_2221);
and U2692 (N_2692,N_2244,N_2148);
nor U2693 (N_2693,N_2126,N_2341);
nor U2694 (N_2694,N_2376,N_1991);
and U2695 (N_2695,N_1825,N_2349);
or U2696 (N_2696,N_1984,N_2031);
and U2697 (N_2697,N_1850,N_2058);
and U2698 (N_2698,N_2099,N_2375);
and U2699 (N_2699,N_2362,N_2270);
nand U2700 (N_2700,N_1990,N_2045);
and U2701 (N_2701,N_2152,N_2146);
or U2702 (N_2702,N_1850,N_2332);
nand U2703 (N_2703,N_2283,N_2086);
nand U2704 (N_2704,N_2263,N_2316);
nor U2705 (N_2705,N_1815,N_1937);
and U2706 (N_2706,N_2007,N_2272);
or U2707 (N_2707,N_2143,N_2316);
nand U2708 (N_2708,N_1815,N_2155);
and U2709 (N_2709,N_2189,N_2179);
nand U2710 (N_2710,N_2171,N_1901);
and U2711 (N_2711,N_2370,N_1872);
or U2712 (N_2712,N_2291,N_2281);
xnor U2713 (N_2713,N_2031,N_2157);
nand U2714 (N_2714,N_2399,N_2273);
and U2715 (N_2715,N_2285,N_2295);
or U2716 (N_2716,N_2066,N_1932);
nor U2717 (N_2717,N_2275,N_2388);
nor U2718 (N_2718,N_1965,N_1941);
or U2719 (N_2719,N_2229,N_1913);
nand U2720 (N_2720,N_2287,N_2000);
nand U2721 (N_2721,N_2044,N_1808);
nand U2722 (N_2722,N_1886,N_2094);
or U2723 (N_2723,N_1901,N_2147);
or U2724 (N_2724,N_2016,N_2328);
nand U2725 (N_2725,N_1937,N_2385);
nand U2726 (N_2726,N_2377,N_2237);
or U2727 (N_2727,N_2285,N_1987);
or U2728 (N_2728,N_2139,N_1939);
or U2729 (N_2729,N_2016,N_2358);
nor U2730 (N_2730,N_2188,N_2381);
nor U2731 (N_2731,N_2237,N_2356);
nor U2732 (N_2732,N_2183,N_2189);
and U2733 (N_2733,N_1938,N_2276);
nor U2734 (N_2734,N_2239,N_1905);
nor U2735 (N_2735,N_2198,N_2256);
nand U2736 (N_2736,N_1975,N_2222);
or U2737 (N_2737,N_2372,N_2310);
or U2738 (N_2738,N_1819,N_2170);
nor U2739 (N_2739,N_1903,N_1973);
and U2740 (N_2740,N_2265,N_1833);
or U2741 (N_2741,N_2034,N_1861);
nor U2742 (N_2742,N_2276,N_2038);
and U2743 (N_2743,N_2117,N_1963);
and U2744 (N_2744,N_2011,N_1835);
and U2745 (N_2745,N_2375,N_1800);
xor U2746 (N_2746,N_2053,N_1802);
and U2747 (N_2747,N_2230,N_2341);
or U2748 (N_2748,N_2275,N_2040);
or U2749 (N_2749,N_2361,N_1977);
nand U2750 (N_2750,N_2196,N_2344);
or U2751 (N_2751,N_2074,N_1826);
nand U2752 (N_2752,N_2227,N_2240);
and U2753 (N_2753,N_1912,N_2061);
and U2754 (N_2754,N_2113,N_2062);
nor U2755 (N_2755,N_2025,N_2229);
nand U2756 (N_2756,N_1919,N_1962);
and U2757 (N_2757,N_1936,N_2137);
and U2758 (N_2758,N_2294,N_1879);
and U2759 (N_2759,N_2204,N_1896);
and U2760 (N_2760,N_2352,N_2275);
or U2761 (N_2761,N_2040,N_1974);
xor U2762 (N_2762,N_2260,N_1973);
nor U2763 (N_2763,N_2245,N_2101);
or U2764 (N_2764,N_2353,N_2278);
nor U2765 (N_2765,N_1839,N_2170);
nand U2766 (N_2766,N_2136,N_2031);
or U2767 (N_2767,N_2040,N_2095);
or U2768 (N_2768,N_2371,N_2200);
and U2769 (N_2769,N_1979,N_2109);
or U2770 (N_2770,N_2197,N_2045);
nand U2771 (N_2771,N_2099,N_2145);
nand U2772 (N_2772,N_1805,N_1828);
and U2773 (N_2773,N_2290,N_2149);
and U2774 (N_2774,N_2005,N_2204);
or U2775 (N_2775,N_2277,N_1821);
nand U2776 (N_2776,N_2393,N_1918);
and U2777 (N_2777,N_2207,N_1827);
nand U2778 (N_2778,N_1811,N_2143);
and U2779 (N_2779,N_1921,N_2060);
and U2780 (N_2780,N_2131,N_2172);
nor U2781 (N_2781,N_2359,N_2014);
nand U2782 (N_2782,N_2342,N_1825);
nor U2783 (N_2783,N_1829,N_2103);
or U2784 (N_2784,N_2285,N_2147);
nor U2785 (N_2785,N_1828,N_2365);
nand U2786 (N_2786,N_1860,N_2062);
nor U2787 (N_2787,N_2029,N_2302);
nand U2788 (N_2788,N_1840,N_2205);
or U2789 (N_2789,N_1909,N_2315);
nand U2790 (N_2790,N_2003,N_2276);
nand U2791 (N_2791,N_1905,N_1960);
or U2792 (N_2792,N_2087,N_1999);
and U2793 (N_2793,N_2182,N_2066);
xnor U2794 (N_2794,N_1858,N_2271);
nand U2795 (N_2795,N_1816,N_1813);
nand U2796 (N_2796,N_1845,N_2105);
nor U2797 (N_2797,N_2116,N_2206);
or U2798 (N_2798,N_2375,N_1916);
and U2799 (N_2799,N_1859,N_2098);
nand U2800 (N_2800,N_2055,N_2098);
nand U2801 (N_2801,N_1958,N_2038);
nand U2802 (N_2802,N_2197,N_1830);
nor U2803 (N_2803,N_2274,N_2053);
nor U2804 (N_2804,N_1904,N_1945);
and U2805 (N_2805,N_1938,N_2216);
nand U2806 (N_2806,N_1856,N_2159);
nand U2807 (N_2807,N_2197,N_2333);
nand U2808 (N_2808,N_2095,N_2338);
nor U2809 (N_2809,N_2116,N_2140);
nand U2810 (N_2810,N_2310,N_2279);
or U2811 (N_2811,N_1943,N_2260);
or U2812 (N_2812,N_2374,N_2105);
nor U2813 (N_2813,N_1983,N_1918);
and U2814 (N_2814,N_1955,N_1848);
or U2815 (N_2815,N_2073,N_1863);
nand U2816 (N_2816,N_2181,N_2048);
nor U2817 (N_2817,N_1810,N_2377);
nand U2818 (N_2818,N_1875,N_2224);
and U2819 (N_2819,N_2074,N_1844);
nor U2820 (N_2820,N_1953,N_2316);
nand U2821 (N_2821,N_2299,N_2099);
nand U2822 (N_2822,N_2153,N_2195);
nand U2823 (N_2823,N_2291,N_2374);
or U2824 (N_2824,N_2286,N_1817);
or U2825 (N_2825,N_1980,N_1903);
or U2826 (N_2826,N_2368,N_2315);
or U2827 (N_2827,N_2026,N_2121);
nor U2828 (N_2828,N_1841,N_2325);
or U2829 (N_2829,N_2013,N_1953);
nand U2830 (N_2830,N_2009,N_2397);
nand U2831 (N_2831,N_2108,N_2168);
and U2832 (N_2832,N_1871,N_2071);
and U2833 (N_2833,N_1958,N_2226);
nand U2834 (N_2834,N_2086,N_2186);
nor U2835 (N_2835,N_2232,N_2382);
nand U2836 (N_2836,N_2394,N_2050);
or U2837 (N_2837,N_2015,N_2021);
nor U2838 (N_2838,N_2195,N_2050);
xnor U2839 (N_2839,N_1926,N_2100);
and U2840 (N_2840,N_1916,N_1918);
or U2841 (N_2841,N_1833,N_2255);
nand U2842 (N_2842,N_2367,N_2125);
or U2843 (N_2843,N_2011,N_2314);
nor U2844 (N_2844,N_2035,N_2168);
nand U2845 (N_2845,N_1941,N_2019);
or U2846 (N_2846,N_2291,N_1919);
and U2847 (N_2847,N_2151,N_2387);
nand U2848 (N_2848,N_2062,N_2145);
nor U2849 (N_2849,N_2231,N_2105);
nand U2850 (N_2850,N_2244,N_2338);
and U2851 (N_2851,N_2360,N_1957);
and U2852 (N_2852,N_1814,N_1950);
or U2853 (N_2853,N_1961,N_2075);
and U2854 (N_2854,N_2291,N_2223);
and U2855 (N_2855,N_1872,N_2191);
nor U2856 (N_2856,N_1895,N_2294);
nand U2857 (N_2857,N_2154,N_1904);
nor U2858 (N_2858,N_2151,N_1928);
nand U2859 (N_2859,N_2023,N_1944);
nand U2860 (N_2860,N_2088,N_2349);
nand U2861 (N_2861,N_2377,N_2225);
nor U2862 (N_2862,N_2033,N_2268);
nand U2863 (N_2863,N_2089,N_2028);
nand U2864 (N_2864,N_2382,N_2074);
or U2865 (N_2865,N_2357,N_2156);
and U2866 (N_2866,N_2278,N_2247);
or U2867 (N_2867,N_2096,N_2030);
nor U2868 (N_2868,N_1916,N_1821);
nor U2869 (N_2869,N_1984,N_2099);
and U2870 (N_2870,N_1998,N_2364);
nand U2871 (N_2871,N_2003,N_2126);
nor U2872 (N_2872,N_2165,N_2200);
and U2873 (N_2873,N_2261,N_2210);
or U2874 (N_2874,N_2318,N_1966);
nor U2875 (N_2875,N_1838,N_1998);
and U2876 (N_2876,N_2228,N_1993);
nand U2877 (N_2877,N_1882,N_2092);
and U2878 (N_2878,N_2090,N_2179);
and U2879 (N_2879,N_2189,N_2219);
or U2880 (N_2880,N_1935,N_2052);
and U2881 (N_2881,N_2115,N_2185);
and U2882 (N_2882,N_2285,N_2306);
nand U2883 (N_2883,N_1821,N_2150);
and U2884 (N_2884,N_1841,N_1839);
or U2885 (N_2885,N_1898,N_1949);
and U2886 (N_2886,N_1960,N_1944);
and U2887 (N_2887,N_1975,N_2322);
and U2888 (N_2888,N_1926,N_1871);
or U2889 (N_2889,N_1946,N_2180);
and U2890 (N_2890,N_1970,N_2096);
nand U2891 (N_2891,N_2110,N_2240);
or U2892 (N_2892,N_2375,N_1882);
or U2893 (N_2893,N_2057,N_1875);
nand U2894 (N_2894,N_2010,N_2393);
or U2895 (N_2895,N_2166,N_1879);
or U2896 (N_2896,N_1859,N_2219);
or U2897 (N_2897,N_1950,N_2220);
nor U2898 (N_2898,N_2066,N_2174);
nor U2899 (N_2899,N_1888,N_1816);
or U2900 (N_2900,N_1894,N_1820);
nor U2901 (N_2901,N_1816,N_1814);
or U2902 (N_2902,N_2350,N_1976);
and U2903 (N_2903,N_2308,N_1986);
and U2904 (N_2904,N_2187,N_1805);
and U2905 (N_2905,N_2387,N_2384);
or U2906 (N_2906,N_2270,N_2006);
nor U2907 (N_2907,N_2358,N_2025);
and U2908 (N_2908,N_2321,N_2163);
nor U2909 (N_2909,N_2294,N_2115);
or U2910 (N_2910,N_2035,N_1975);
or U2911 (N_2911,N_1817,N_1964);
or U2912 (N_2912,N_2337,N_1899);
nand U2913 (N_2913,N_2234,N_2332);
nor U2914 (N_2914,N_2388,N_2068);
or U2915 (N_2915,N_2104,N_2041);
and U2916 (N_2916,N_2034,N_2059);
and U2917 (N_2917,N_2208,N_2275);
or U2918 (N_2918,N_2382,N_2096);
and U2919 (N_2919,N_2055,N_2189);
nand U2920 (N_2920,N_1806,N_1927);
nor U2921 (N_2921,N_1916,N_2059);
or U2922 (N_2922,N_2015,N_1889);
or U2923 (N_2923,N_2045,N_2329);
or U2924 (N_2924,N_2379,N_2299);
or U2925 (N_2925,N_2124,N_2190);
and U2926 (N_2926,N_2108,N_1881);
and U2927 (N_2927,N_2032,N_2385);
nand U2928 (N_2928,N_1871,N_2387);
or U2929 (N_2929,N_1928,N_2340);
nor U2930 (N_2930,N_1898,N_1948);
or U2931 (N_2931,N_1813,N_2339);
nor U2932 (N_2932,N_2060,N_1928);
nand U2933 (N_2933,N_1964,N_2112);
nor U2934 (N_2934,N_1866,N_2090);
and U2935 (N_2935,N_2093,N_2369);
and U2936 (N_2936,N_2220,N_1877);
or U2937 (N_2937,N_2384,N_1927);
nor U2938 (N_2938,N_1967,N_2057);
nor U2939 (N_2939,N_1887,N_1851);
or U2940 (N_2940,N_2040,N_2140);
or U2941 (N_2941,N_2386,N_1842);
nor U2942 (N_2942,N_2165,N_2149);
and U2943 (N_2943,N_2341,N_2064);
or U2944 (N_2944,N_2284,N_2052);
or U2945 (N_2945,N_2268,N_1826);
nor U2946 (N_2946,N_2172,N_1816);
nand U2947 (N_2947,N_1998,N_2069);
nand U2948 (N_2948,N_2134,N_2190);
nand U2949 (N_2949,N_2161,N_2373);
and U2950 (N_2950,N_2295,N_2215);
and U2951 (N_2951,N_2008,N_2099);
nand U2952 (N_2952,N_1919,N_2225);
nand U2953 (N_2953,N_1973,N_2167);
nor U2954 (N_2954,N_2394,N_2112);
or U2955 (N_2955,N_2115,N_2110);
or U2956 (N_2956,N_1970,N_2280);
and U2957 (N_2957,N_1985,N_2293);
nor U2958 (N_2958,N_2047,N_2298);
nand U2959 (N_2959,N_2351,N_2022);
nand U2960 (N_2960,N_2180,N_2159);
nand U2961 (N_2961,N_2074,N_2359);
and U2962 (N_2962,N_2314,N_2255);
nor U2963 (N_2963,N_2210,N_2310);
or U2964 (N_2964,N_2104,N_2058);
nand U2965 (N_2965,N_2218,N_1878);
or U2966 (N_2966,N_1922,N_1935);
or U2967 (N_2967,N_1831,N_1882);
nor U2968 (N_2968,N_2163,N_2395);
nor U2969 (N_2969,N_2123,N_2258);
or U2970 (N_2970,N_1888,N_2224);
and U2971 (N_2971,N_2034,N_2123);
nand U2972 (N_2972,N_2009,N_2116);
nor U2973 (N_2973,N_1886,N_2375);
and U2974 (N_2974,N_2393,N_2211);
and U2975 (N_2975,N_2293,N_2336);
nor U2976 (N_2976,N_2243,N_2341);
or U2977 (N_2977,N_1848,N_2108);
nor U2978 (N_2978,N_2009,N_2206);
nand U2979 (N_2979,N_1802,N_1941);
nor U2980 (N_2980,N_2359,N_2097);
or U2981 (N_2981,N_2183,N_2179);
nor U2982 (N_2982,N_2196,N_2215);
nor U2983 (N_2983,N_1837,N_2321);
nor U2984 (N_2984,N_2237,N_1826);
nor U2985 (N_2985,N_2213,N_2327);
nand U2986 (N_2986,N_2091,N_2357);
or U2987 (N_2987,N_2176,N_2137);
nand U2988 (N_2988,N_2090,N_2027);
nand U2989 (N_2989,N_2038,N_1824);
nor U2990 (N_2990,N_2247,N_2169);
and U2991 (N_2991,N_2347,N_1801);
or U2992 (N_2992,N_1899,N_1947);
or U2993 (N_2993,N_2079,N_2120);
nand U2994 (N_2994,N_1808,N_1980);
or U2995 (N_2995,N_2131,N_1903);
nor U2996 (N_2996,N_2215,N_2015);
nand U2997 (N_2997,N_2039,N_2377);
or U2998 (N_2998,N_1819,N_1958);
or U2999 (N_2999,N_2314,N_2203);
or UO_0 (O_0,N_2449,N_2652);
nor UO_1 (O_1,N_2974,N_2406);
or UO_2 (O_2,N_2711,N_2849);
nand UO_3 (O_3,N_2760,N_2848);
and UO_4 (O_4,N_2740,N_2705);
nand UO_5 (O_5,N_2425,N_2748);
and UO_6 (O_6,N_2498,N_2957);
and UO_7 (O_7,N_2643,N_2684);
or UO_8 (O_8,N_2818,N_2501);
nand UO_9 (O_9,N_2738,N_2701);
and UO_10 (O_10,N_2671,N_2942);
and UO_11 (O_11,N_2904,N_2610);
nand UO_12 (O_12,N_2598,N_2800);
nand UO_13 (O_13,N_2785,N_2676);
nand UO_14 (O_14,N_2489,N_2654);
or UO_15 (O_15,N_2504,N_2969);
nor UO_16 (O_16,N_2958,N_2524);
nor UO_17 (O_17,N_2685,N_2772);
nand UO_18 (O_18,N_2719,N_2499);
and UO_19 (O_19,N_2949,N_2619);
and UO_20 (O_20,N_2722,N_2548);
and UO_21 (O_21,N_2846,N_2412);
and UO_22 (O_22,N_2894,N_2820);
and UO_23 (O_23,N_2952,N_2693);
and UO_24 (O_24,N_2937,N_2821);
xor UO_25 (O_25,N_2703,N_2727);
and UO_26 (O_26,N_2717,N_2563);
nor UO_27 (O_27,N_2561,N_2745);
nor UO_28 (O_28,N_2567,N_2679);
and UO_29 (O_29,N_2825,N_2658);
and UO_30 (O_30,N_2782,N_2812);
nand UO_31 (O_31,N_2605,N_2726);
nand UO_32 (O_32,N_2988,N_2669);
or UO_33 (O_33,N_2990,N_2966);
nor UO_34 (O_34,N_2634,N_2427);
and UO_35 (O_35,N_2411,N_2421);
and UO_36 (O_36,N_2809,N_2989);
nor UO_37 (O_37,N_2930,N_2725);
nor UO_38 (O_38,N_2569,N_2761);
nor UO_39 (O_39,N_2571,N_2845);
and UO_40 (O_40,N_2746,N_2729);
nand UO_41 (O_41,N_2650,N_2852);
nand UO_42 (O_42,N_2649,N_2987);
nor UO_43 (O_43,N_2624,N_2826);
and UO_44 (O_44,N_2662,N_2886);
or UO_45 (O_45,N_2781,N_2739);
and UO_46 (O_46,N_2713,N_2919);
or UO_47 (O_47,N_2622,N_2796);
and UO_48 (O_48,N_2514,N_2776);
or UO_49 (O_49,N_2842,N_2774);
nor UO_50 (O_50,N_2881,N_2480);
nand UO_51 (O_51,N_2893,N_2420);
nor UO_52 (O_52,N_2418,N_2996);
and UO_53 (O_53,N_2759,N_2707);
and UO_54 (O_54,N_2861,N_2606);
nor UO_55 (O_55,N_2699,N_2939);
nor UO_56 (O_56,N_2494,N_2803);
nand UO_57 (O_57,N_2674,N_2791);
nor UO_58 (O_58,N_2793,N_2595);
or UO_59 (O_59,N_2899,N_2863);
nor UO_60 (O_60,N_2922,N_2664);
and UO_61 (O_61,N_2604,N_2520);
nand UO_62 (O_62,N_2445,N_2545);
nand UO_63 (O_63,N_2710,N_2709);
nand UO_64 (O_64,N_2733,N_2630);
or UO_65 (O_65,N_2638,N_2801);
nor UO_66 (O_66,N_2694,N_2751);
and UO_67 (O_67,N_2461,N_2565);
nand UO_68 (O_68,N_2933,N_2683);
nor UO_69 (O_69,N_2542,N_2534);
nor UO_70 (O_70,N_2889,N_2620);
nand UO_71 (O_71,N_2491,N_2764);
or UO_72 (O_72,N_2730,N_2997);
or UO_73 (O_73,N_2452,N_2768);
nor UO_74 (O_74,N_2525,N_2581);
and UO_75 (O_75,N_2758,N_2515);
nor UO_76 (O_76,N_2871,N_2962);
or UO_77 (O_77,N_2789,N_2872);
nor UO_78 (O_78,N_2923,N_2435);
nor UO_79 (O_79,N_2478,N_2940);
and UO_80 (O_80,N_2559,N_2436);
nand UO_81 (O_81,N_2568,N_2955);
nand UO_82 (O_82,N_2858,N_2762);
and UO_83 (O_83,N_2792,N_2991);
nor UO_84 (O_84,N_2680,N_2844);
and UO_85 (O_85,N_2602,N_2765);
nor UO_86 (O_86,N_2831,N_2413);
and UO_87 (O_87,N_2843,N_2552);
and UO_88 (O_88,N_2407,N_2967);
and UO_89 (O_89,N_2742,N_2888);
or UO_90 (O_90,N_2932,N_2579);
and UO_91 (O_91,N_2496,N_2948);
nor UO_92 (O_92,N_2814,N_2516);
nor UO_93 (O_93,N_2799,N_2455);
nand UO_94 (O_94,N_2657,N_2954);
or UO_95 (O_95,N_2651,N_2484);
or UO_96 (O_96,N_2783,N_2440);
nand UO_97 (O_97,N_2497,N_2655);
nand UO_98 (O_98,N_2806,N_2934);
or UO_99 (O_99,N_2599,N_2750);
and UO_100 (O_100,N_2891,N_2464);
nand UO_101 (O_101,N_2840,N_2867);
nand UO_102 (O_102,N_2741,N_2572);
and UO_103 (O_103,N_2626,N_2453);
or UO_104 (O_104,N_2928,N_2656);
nor UO_105 (O_105,N_2535,N_2859);
nand UO_106 (O_106,N_2860,N_2482);
xnor UO_107 (O_107,N_2476,N_2580);
nand UO_108 (O_108,N_2855,N_2551);
and UO_109 (O_109,N_2704,N_2743);
or UO_110 (O_110,N_2659,N_2526);
or UO_111 (O_111,N_2841,N_2414);
nand UO_112 (O_112,N_2540,N_2999);
or UO_113 (O_113,N_2698,N_2457);
or UO_114 (O_114,N_2570,N_2640);
nand UO_115 (O_115,N_2965,N_2635);
nand UO_116 (O_116,N_2943,N_2441);
or UO_117 (O_117,N_2603,N_2788);
or UO_118 (O_118,N_2981,N_2797);
or UO_119 (O_119,N_2992,N_2837);
nor UO_120 (O_120,N_2682,N_2500);
nor UO_121 (O_121,N_2884,N_2824);
or UO_122 (O_122,N_2926,N_2642);
or UO_123 (O_123,N_2446,N_2465);
or UO_124 (O_124,N_2834,N_2578);
nor UO_125 (O_125,N_2877,N_2616);
and UO_126 (O_126,N_2876,N_2617);
or UO_127 (O_127,N_2665,N_2503);
nand UO_128 (O_128,N_2442,N_2668);
and UO_129 (O_129,N_2778,N_2550);
or UO_130 (O_130,N_2632,N_2790);
or UO_131 (O_131,N_2596,N_2558);
nor UO_132 (O_132,N_2838,N_2645);
nand UO_133 (O_133,N_2405,N_2973);
nand UO_134 (O_134,N_2646,N_2708);
or UO_135 (O_135,N_2927,N_2663);
or UO_136 (O_136,N_2555,N_2444);
nand UO_137 (O_137,N_2416,N_2808);
nor UO_138 (O_138,N_2623,N_2544);
or UO_139 (O_139,N_2731,N_2985);
nand UO_140 (O_140,N_2979,N_2404);
nor UO_141 (O_141,N_2470,N_2766);
nand UO_142 (O_142,N_2787,N_2994);
and UO_143 (O_143,N_2706,N_2865);
or UO_144 (O_144,N_2467,N_2850);
nand UO_145 (O_145,N_2475,N_2970);
nor UO_146 (O_146,N_2753,N_2718);
nor UO_147 (O_147,N_2784,N_2590);
nor UO_148 (O_148,N_2944,N_2666);
nand UO_149 (O_149,N_2980,N_2828);
nand UO_150 (O_150,N_2870,N_2851);
nand UO_151 (O_151,N_2408,N_2830);
and UO_152 (O_152,N_2529,N_2660);
nor UO_153 (O_153,N_2959,N_2873);
or UO_154 (O_154,N_2816,N_2953);
nor UO_155 (O_155,N_2433,N_2462);
or UO_156 (O_156,N_2409,N_2417);
nand UO_157 (O_157,N_2908,N_2874);
nand UO_158 (O_158,N_2528,N_2530);
nor UO_159 (O_159,N_2786,N_2920);
nor UO_160 (O_160,N_2594,N_2907);
nor UO_161 (O_161,N_2681,N_2986);
xnor UO_162 (O_162,N_2607,N_2913);
nor UO_163 (O_163,N_2724,N_2403);
and UO_164 (O_164,N_2755,N_2511);
nor UO_165 (O_165,N_2575,N_2495);
or UO_166 (O_166,N_2805,N_2431);
and UO_167 (O_167,N_2744,N_2715);
nand UO_168 (O_168,N_2956,N_2687);
or UO_169 (O_169,N_2775,N_2773);
or UO_170 (O_170,N_2631,N_2895);
and UO_171 (O_171,N_2589,N_2438);
nand UO_172 (O_172,N_2911,N_2835);
and UO_173 (O_173,N_2424,N_2880);
nor UO_174 (O_174,N_2609,N_2422);
nand UO_175 (O_175,N_2400,N_2771);
and UO_176 (O_176,N_2519,N_2734);
nor UO_177 (O_177,N_2536,N_2882);
nor UO_178 (O_178,N_2915,N_2938);
and UO_179 (O_179,N_2521,N_2560);
and UO_180 (O_180,N_2833,N_2747);
nand UO_181 (O_181,N_2639,N_2728);
or UO_182 (O_182,N_2419,N_2829);
or UO_183 (O_183,N_2615,N_2901);
nand UO_184 (O_184,N_2592,N_2976);
and UO_185 (O_185,N_2921,N_2960);
or UO_186 (O_186,N_2968,N_2857);
and UO_187 (O_187,N_2532,N_2853);
or UO_188 (O_188,N_2777,N_2716);
nand UO_189 (O_189,N_2736,N_2839);
and UO_190 (O_190,N_2443,N_2430);
and UO_191 (O_191,N_2804,N_2512);
nor UO_192 (O_192,N_2896,N_2754);
and UO_193 (O_193,N_2964,N_2897);
nand UO_194 (O_194,N_2869,N_2584);
nor UO_195 (O_195,N_2410,N_2629);
nor UO_196 (O_196,N_2636,N_2518);
or UO_197 (O_197,N_2672,N_2454);
or UO_198 (O_198,N_2537,N_2677);
or UO_199 (O_199,N_2434,N_2696);
or UO_200 (O_200,N_2914,N_2533);
nand UO_201 (O_201,N_2678,N_2557);
and UO_202 (O_202,N_2608,N_2924);
nor UO_203 (O_203,N_2688,N_2689);
nand UO_204 (O_204,N_2628,N_2813);
nand UO_205 (O_205,N_2582,N_2459);
nor UO_206 (O_206,N_2721,N_2898);
and UO_207 (O_207,N_2735,N_2902);
or UO_208 (O_208,N_2866,N_2505);
nor UO_209 (O_209,N_2692,N_2998);
and UO_210 (O_210,N_2458,N_2490);
or UO_211 (O_211,N_2903,N_2890);
or UO_212 (O_212,N_2673,N_2538);
or UO_213 (O_213,N_2509,N_2426);
and UO_214 (O_214,N_2428,N_2702);
nand UO_215 (O_215,N_2633,N_2507);
or UO_216 (O_216,N_2946,N_2597);
or UO_217 (O_217,N_2593,N_2466);
nor UO_218 (O_218,N_2982,N_2448);
nor UO_219 (O_219,N_2543,N_2947);
nor UO_220 (O_220,N_2802,N_2963);
nor UO_221 (O_221,N_2648,N_2941);
nor UO_222 (O_222,N_2492,N_2527);
or UO_223 (O_223,N_2690,N_2720);
and UO_224 (O_224,N_2574,N_2749);
and UO_225 (O_225,N_2862,N_2637);
or UO_226 (O_226,N_2807,N_2474);
or UO_227 (O_227,N_2686,N_2779);
and UO_228 (O_228,N_2832,N_2487);
nand UO_229 (O_229,N_2780,N_2469);
or UO_230 (O_230,N_2613,N_2883);
or UO_231 (O_231,N_2795,N_2670);
nor UO_232 (O_232,N_2879,N_2547);
or UO_233 (O_233,N_2556,N_2910);
or UO_234 (O_234,N_2611,N_2506);
nand UO_235 (O_235,N_2697,N_2432);
nor UO_236 (O_236,N_2591,N_2522);
nand UO_237 (O_237,N_2588,N_2647);
nand UO_238 (O_238,N_2401,N_2485);
and UO_239 (O_239,N_2577,N_2752);
nor UO_240 (O_240,N_2885,N_2864);
or UO_241 (O_241,N_2463,N_2798);
or UO_242 (O_242,N_2539,N_2479);
and UO_243 (O_243,N_2732,N_2481);
and UO_244 (O_244,N_2827,N_2936);
or UO_245 (O_245,N_2977,N_2460);
nand UO_246 (O_246,N_2868,N_2887);
or UO_247 (O_247,N_2586,N_2916);
or UO_248 (O_248,N_2429,N_2925);
nor UO_249 (O_249,N_2439,N_2486);
nor UO_250 (O_250,N_2437,N_2587);
or UO_251 (O_251,N_2723,N_2553);
or UO_252 (O_252,N_2661,N_2810);
or UO_253 (O_253,N_2614,N_2971);
nand UO_254 (O_254,N_2945,N_2667);
and UO_255 (O_255,N_2714,N_2935);
nor UO_256 (O_256,N_2618,N_2905);
and UO_257 (O_257,N_2585,N_2531);
nand UO_258 (O_258,N_2508,N_2456);
nand UO_259 (O_259,N_2906,N_2601);
nand UO_260 (O_260,N_2566,N_2917);
and UO_261 (O_261,N_2468,N_2415);
nor UO_262 (O_262,N_2929,N_2493);
nand UO_263 (O_263,N_2819,N_2909);
nor UO_264 (O_264,N_2447,N_2875);
nand UO_265 (O_265,N_2811,N_2767);
nor UO_266 (O_266,N_2961,N_2600);
nand UO_267 (O_267,N_2918,N_2576);
or UO_268 (O_268,N_2878,N_2621);
or UO_269 (O_269,N_2978,N_2972);
nand UO_270 (O_270,N_2984,N_2471);
and UO_271 (O_271,N_2712,N_2912);
and UO_272 (O_272,N_2562,N_2477);
and UO_273 (O_273,N_2513,N_2402);
and UO_274 (O_274,N_2757,N_2695);
or UO_275 (O_275,N_2423,N_2854);
nand UO_276 (O_276,N_2541,N_2951);
nand UO_277 (O_277,N_2625,N_2770);
nor UO_278 (O_278,N_2892,N_2737);
nand UO_279 (O_279,N_2564,N_2644);
nor UO_280 (O_280,N_2510,N_2627);
nor UO_281 (O_281,N_2950,N_2488);
and UO_282 (O_282,N_2546,N_2554);
or UO_283 (O_283,N_2856,N_2641);
nand UO_284 (O_284,N_2472,N_2502);
nor UO_285 (O_285,N_2573,N_2815);
and UO_286 (O_286,N_2822,N_2517);
nor UO_287 (O_287,N_2794,N_2700);
nor UO_288 (O_288,N_2675,N_2483);
nand UO_289 (O_289,N_2769,N_2763);
and UO_290 (O_290,N_2823,N_2931);
and UO_291 (O_291,N_2993,N_2817);
nor UO_292 (O_292,N_2523,N_2983);
nand UO_293 (O_293,N_2975,N_2756);
or UO_294 (O_294,N_2473,N_2847);
nor UO_295 (O_295,N_2612,N_2451);
and UO_296 (O_296,N_2836,N_2691);
nand UO_297 (O_297,N_2995,N_2450);
nand UO_298 (O_298,N_2653,N_2900);
nor UO_299 (O_299,N_2549,N_2583);
nor UO_300 (O_300,N_2969,N_2849);
and UO_301 (O_301,N_2865,N_2967);
nor UO_302 (O_302,N_2676,N_2624);
nand UO_303 (O_303,N_2503,N_2425);
nand UO_304 (O_304,N_2820,N_2401);
or UO_305 (O_305,N_2589,N_2833);
and UO_306 (O_306,N_2943,N_2559);
nand UO_307 (O_307,N_2609,N_2660);
and UO_308 (O_308,N_2881,N_2991);
nor UO_309 (O_309,N_2912,N_2562);
and UO_310 (O_310,N_2574,N_2664);
nor UO_311 (O_311,N_2444,N_2469);
or UO_312 (O_312,N_2545,N_2688);
and UO_313 (O_313,N_2985,N_2689);
and UO_314 (O_314,N_2933,N_2623);
and UO_315 (O_315,N_2881,N_2982);
or UO_316 (O_316,N_2571,N_2591);
or UO_317 (O_317,N_2783,N_2576);
nand UO_318 (O_318,N_2872,N_2684);
and UO_319 (O_319,N_2482,N_2746);
nor UO_320 (O_320,N_2856,N_2709);
or UO_321 (O_321,N_2524,N_2916);
or UO_322 (O_322,N_2777,N_2799);
nor UO_323 (O_323,N_2637,N_2953);
nand UO_324 (O_324,N_2883,N_2888);
or UO_325 (O_325,N_2822,N_2585);
and UO_326 (O_326,N_2821,N_2946);
or UO_327 (O_327,N_2476,N_2839);
and UO_328 (O_328,N_2581,N_2845);
nand UO_329 (O_329,N_2911,N_2760);
and UO_330 (O_330,N_2686,N_2980);
or UO_331 (O_331,N_2950,N_2549);
or UO_332 (O_332,N_2976,N_2603);
nor UO_333 (O_333,N_2901,N_2960);
and UO_334 (O_334,N_2784,N_2595);
and UO_335 (O_335,N_2689,N_2461);
nand UO_336 (O_336,N_2526,N_2758);
nand UO_337 (O_337,N_2713,N_2734);
nor UO_338 (O_338,N_2484,N_2903);
or UO_339 (O_339,N_2923,N_2769);
and UO_340 (O_340,N_2422,N_2712);
nand UO_341 (O_341,N_2429,N_2804);
or UO_342 (O_342,N_2775,N_2853);
and UO_343 (O_343,N_2576,N_2930);
nand UO_344 (O_344,N_2982,N_2723);
or UO_345 (O_345,N_2980,N_2748);
nor UO_346 (O_346,N_2923,N_2832);
and UO_347 (O_347,N_2908,N_2734);
or UO_348 (O_348,N_2976,N_2462);
nand UO_349 (O_349,N_2810,N_2538);
and UO_350 (O_350,N_2956,N_2651);
and UO_351 (O_351,N_2800,N_2558);
nand UO_352 (O_352,N_2556,N_2734);
nor UO_353 (O_353,N_2862,N_2590);
nand UO_354 (O_354,N_2973,N_2977);
and UO_355 (O_355,N_2730,N_2787);
nor UO_356 (O_356,N_2628,N_2926);
nand UO_357 (O_357,N_2775,N_2924);
xnor UO_358 (O_358,N_2922,N_2809);
and UO_359 (O_359,N_2892,N_2971);
and UO_360 (O_360,N_2799,N_2986);
nor UO_361 (O_361,N_2629,N_2776);
or UO_362 (O_362,N_2867,N_2431);
and UO_363 (O_363,N_2424,N_2456);
nor UO_364 (O_364,N_2710,N_2994);
and UO_365 (O_365,N_2890,N_2778);
nand UO_366 (O_366,N_2923,N_2427);
and UO_367 (O_367,N_2561,N_2654);
and UO_368 (O_368,N_2549,N_2925);
nor UO_369 (O_369,N_2687,N_2731);
or UO_370 (O_370,N_2887,N_2588);
nor UO_371 (O_371,N_2710,N_2641);
nor UO_372 (O_372,N_2734,N_2816);
nand UO_373 (O_373,N_2949,N_2532);
nor UO_374 (O_374,N_2435,N_2669);
and UO_375 (O_375,N_2627,N_2692);
nand UO_376 (O_376,N_2778,N_2663);
and UO_377 (O_377,N_2758,N_2765);
and UO_378 (O_378,N_2501,N_2640);
and UO_379 (O_379,N_2459,N_2994);
and UO_380 (O_380,N_2685,N_2501);
or UO_381 (O_381,N_2455,N_2704);
or UO_382 (O_382,N_2621,N_2550);
nor UO_383 (O_383,N_2744,N_2828);
and UO_384 (O_384,N_2953,N_2858);
nand UO_385 (O_385,N_2981,N_2637);
and UO_386 (O_386,N_2536,N_2438);
nor UO_387 (O_387,N_2841,N_2977);
or UO_388 (O_388,N_2889,N_2950);
nor UO_389 (O_389,N_2742,N_2462);
or UO_390 (O_390,N_2845,N_2627);
nor UO_391 (O_391,N_2557,N_2969);
nor UO_392 (O_392,N_2970,N_2500);
nand UO_393 (O_393,N_2417,N_2837);
nand UO_394 (O_394,N_2538,N_2628);
nand UO_395 (O_395,N_2557,N_2463);
or UO_396 (O_396,N_2872,N_2548);
nor UO_397 (O_397,N_2413,N_2867);
nor UO_398 (O_398,N_2568,N_2891);
and UO_399 (O_399,N_2962,N_2463);
nor UO_400 (O_400,N_2569,N_2495);
nor UO_401 (O_401,N_2973,N_2462);
xnor UO_402 (O_402,N_2876,N_2822);
nor UO_403 (O_403,N_2983,N_2896);
or UO_404 (O_404,N_2677,N_2999);
or UO_405 (O_405,N_2913,N_2741);
and UO_406 (O_406,N_2573,N_2602);
xor UO_407 (O_407,N_2539,N_2871);
nand UO_408 (O_408,N_2545,N_2917);
nor UO_409 (O_409,N_2522,N_2954);
and UO_410 (O_410,N_2682,N_2782);
nor UO_411 (O_411,N_2596,N_2664);
and UO_412 (O_412,N_2744,N_2953);
or UO_413 (O_413,N_2947,N_2740);
and UO_414 (O_414,N_2814,N_2540);
nor UO_415 (O_415,N_2472,N_2589);
and UO_416 (O_416,N_2783,N_2686);
and UO_417 (O_417,N_2806,N_2461);
or UO_418 (O_418,N_2822,N_2439);
or UO_419 (O_419,N_2549,N_2495);
or UO_420 (O_420,N_2678,N_2793);
and UO_421 (O_421,N_2747,N_2460);
and UO_422 (O_422,N_2492,N_2647);
and UO_423 (O_423,N_2736,N_2742);
or UO_424 (O_424,N_2458,N_2433);
or UO_425 (O_425,N_2594,N_2977);
nor UO_426 (O_426,N_2800,N_2493);
or UO_427 (O_427,N_2610,N_2586);
nor UO_428 (O_428,N_2868,N_2971);
or UO_429 (O_429,N_2604,N_2649);
nand UO_430 (O_430,N_2627,N_2994);
nor UO_431 (O_431,N_2732,N_2400);
nand UO_432 (O_432,N_2720,N_2768);
nor UO_433 (O_433,N_2467,N_2622);
or UO_434 (O_434,N_2943,N_2640);
nand UO_435 (O_435,N_2878,N_2648);
or UO_436 (O_436,N_2458,N_2432);
nor UO_437 (O_437,N_2839,N_2446);
nand UO_438 (O_438,N_2433,N_2982);
nor UO_439 (O_439,N_2828,N_2526);
and UO_440 (O_440,N_2901,N_2823);
or UO_441 (O_441,N_2910,N_2692);
nand UO_442 (O_442,N_2674,N_2953);
and UO_443 (O_443,N_2758,N_2746);
or UO_444 (O_444,N_2448,N_2835);
or UO_445 (O_445,N_2627,N_2847);
and UO_446 (O_446,N_2760,N_2927);
nor UO_447 (O_447,N_2719,N_2534);
nor UO_448 (O_448,N_2687,N_2800);
nand UO_449 (O_449,N_2448,N_2810);
and UO_450 (O_450,N_2516,N_2767);
or UO_451 (O_451,N_2442,N_2555);
nand UO_452 (O_452,N_2662,N_2748);
nor UO_453 (O_453,N_2770,N_2789);
nor UO_454 (O_454,N_2746,N_2559);
or UO_455 (O_455,N_2784,N_2682);
nand UO_456 (O_456,N_2993,N_2496);
nand UO_457 (O_457,N_2988,N_2490);
or UO_458 (O_458,N_2929,N_2670);
nor UO_459 (O_459,N_2895,N_2546);
nor UO_460 (O_460,N_2701,N_2654);
nor UO_461 (O_461,N_2512,N_2746);
nand UO_462 (O_462,N_2877,N_2712);
nand UO_463 (O_463,N_2711,N_2506);
and UO_464 (O_464,N_2686,N_2941);
and UO_465 (O_465,N_2465,N_2618);
and UO_466 (O_466,N_2960,N_2756);
nor UO_467 (O_467,N_2409,N_2880);
nor UO_468 (O_468,N_2799,N_2599);
nor UO_469 (O_469,N_2683,N_2449);
or UO_470 (O_470,N_2400,N_2786);
and UO_471 (O_471,N_2883,N_2489);
or UO_472 (O_472,N_2617,N_2896);
nor UO_473 (O_473,N_2691,N_2759);
nor UO_474 (O_474,N_2527,N_2411);
or UO_475 (O_475,N_2403,N_2665);
or UO_476 (O_476,N_2732,N_2575);
and UO_477 (O_477,N_2439,N_2733);
or UO_478 (O_478,N_2513,N_2531);
nand UO_479 (O_479,N_2960,N_2708);
or UO_480 (O_480,N_2637,N_2912);
and UO_481 (O_481,N_2421,N_2951);
nor UO_482 (O_482,N_2874,N_2788);
or UO_483 (O_483,N_2435,N_2892);
or UO_484 (O_484,N_2562,N_2639);
and UO_485 (O_485,N_2415,N_2646);
and UO_486 (O_486,N_2411,N_2876);
nand UO_487 (O_487,N_2707,N_2661);
or UO_488 (O_488,N_2423,N_2587);
nand UO_489 (O_489,N_2989,N_2865);
xnor UO_490 (O_490,N_2951,N_2708);
nor UO_491 (O_491,N_2822,N_2587);
nand UO_492 (O_492,N_2663,N_2711);
or UO_493 (O_493,N_2475,N_2404);
and UO_494 (O_494,N_2761,N_2907);
and UO_495 (O_495,N_2817,N_2682);
or UO_496 (O_496,N_2708,N_2838);
or UO_497 (O_497,N_2826,N_2432);
or UO_498 (O_498,N_2751,N_2800);
or UO_499 (O_499,N_2596,N_2803);
endmodule