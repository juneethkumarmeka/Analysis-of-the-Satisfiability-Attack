module basic_750_5000_1000_2_levels_5xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2525,N_2527,N_2528,N_2529,N_2530,N_2532,N_2533,N_2534,N_2535,N_2536,N_2538,N_2539,N_2540,N_2543,N_2544,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2566,N_2568,N_2569,N_2570,N_2571,N_2572,N_2574,N_2575,N_2576,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2599,N_2600,N_2601,N_2602,N_2604,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2644,N_2645,N_2646,N_2647,N_2648,N_2650,N_2651,N_2652,N_2654,N_2655,N_2656,N_2658,N_2659,N_2661,N_2663,N_2665,N_2666,N_2669,N_2671,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2714,N_2716,N_2717,N_2720,N_2721,N_2722,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2732,N_2733,N_2734,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2752,N_2753,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2766,N_2767,N_2768,N_2770,N_2771,N_2772,N_2775,N_2776,N_2778,N_2781,N_2782,N_2784,N_2786,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2805,N_2806,N_2808,N_2809,N_2810,N_2812,N_2813,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2824,N_2825,N_2826,N_2827,N_2829,N_2830,N_2831,N_2832,N_2834,N_2836,N_2837,N_2838,N_2839,N_2841,N_2842,N_2844,N_2845,N_2846,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2857,N_2859,N_2860,N_2862,N_2863,N_2864,N_2865,N_2866,N_2868,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2880,N_2881,N_2882,N_2883,N_2884,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2967,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2977,N_2978,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2989,N_2990,N_2991,N_2993,N_2994,N_2995,N_2996,N_2997,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3007,N_3008,N_3012,N_3013,N_3014,N_3016,N_3018,N_3020,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3059,N_3061,N_3062,N_3063,N_3064,N_3065,N_3067,N_3070,N_3072,N_3074,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3097,N_3099,N_3100,N_3101,N_3102,N_3104,N_3106,N_3107,N_3110,N_3111,N_3112,N_3113,N_3114,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3129,N_3130,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3140,N_3141,N_3143,N_3144,N_3145,N_3146,N_3148,N_3150,N_3151,N_3155,N_3157,N_3160,N_3161,N_3162,N_3164,N_3165,N_3166,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3176,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3189,N_3190,N_3191,N_3192,N_3193,N_3195,N_3196,N_3198,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3214,N_3215,N_3216,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3228,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3241,N_3242,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3252,N_3253,N_3254,N_3255,N_3258,N_3259,N_3261,N_3262,N_3264,N_3265,N_3266,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3280,N_3281,N_3283,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3315,N_3316,N_3319,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3340,N_3341,N_3344,N_3346,N_3349,N_3350,N_3355,N_3356,N_3357,N_3358,N_3359,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3391,N_3392,N_3393,N_3394,N_3396,N_3397,N_3398,N_3399,N_3400,N_3402,N_3403,N_3404,N_3405,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3420,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3435,N_3436,N_3438,N_3439,N_3440,N_3441,N_3443,N_3444,N_3447,N_3448,N_3449,N_3450,N_3451,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3477,N_3478,N_3479,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3498,N_3499,N_3500,N_3501,N_3502,N_3504,N_3506,N_3507,N_3508,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3538,N_3539,N_3541,N_3542,N_3543,N_3544,N_3546,N_3547,N_3548,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3558,N_3559,N_3560,N_3561,N_3562,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3585,N_3586,N_3587,N_3589,N_3590,N_3591,N_3592,N_3594,N_3595,N_3596,N_3598,N_3599,N_3602,N_3603,N_3604,N_3606,N_3609,N_3610,N_3611,N_3612,N_3613,N_3615,N_3616,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3632,N_3634,N_3635,N_3636,N_3637,N_3638,N_3640,N_3641,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3653,N_3654,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3682,N_3683,N_3684,N_3685,N_3687,N_3689,N_3692,N_3693,N_3694,N_3695,N_3696,N_3698,N_3699,N_3700,N_3701,N_3702,N_3704,N_3706,N_3707,N_3709,N_3710,N_3712,N_3714,N_3715,N_3716,N_3717,N_3719,N_3720,N_3721,N_3722,N_3723,N_3725,N_3726,N_3727,N_3728,N_3729,N_3731,N_3732,N_3734,N_3736,N_3737,N_3738,N_3739,N_3742,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3751,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3777,N_3778,N_3779,N_3782,N_3783,N_3784,N_3785,N_3787,N_3788,N_3789,N_3790,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3801,N_3802,N_3803,N_3804,N_3806,N_3809,N_3810,N_3811,N_3814,N_3815,N_3816,N_3818,N_3819,N_3821,N_3822,N_3823,N_3824,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3843,N_3845,N_3846,N_3847,N_3848,N_3849,N_3851,N_3852,N_3854,N_3855,N_3856,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3904,N_3905,N_3907,N_3908,N_3909,N_3910,N_3912,N_3913,N_3914,N_3915,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3952,N_3953,N_3954,N_3957,N_3959,N_3961,N_3962,N_3964,N_3965,N_3967,N_3968,N_3969,N_3970,N_3972,N_3973,N_3974,N_3975,N_3976,N_3979,N_3980,N_3983,N_3985,N_3986,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4003,N_4004,N_4005,N_4006,N_4008,N_4010,N_4011,N_4012,N_4013,N_4014,N_4017,N_4018,N_4020,N_4021,N_4022,N_4023,N_4024,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4037,N_4038,N_4040,N_4042,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4055,N_4056,N_4057,N_4060,N_4061,N_4062,N_4063,N_4065,N_4066,N_4067,N_4068,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4079,N_4081,N_4082,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4105,N_4107,N_4109,N_4110,N_4111,N_4112,N_4113,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4126,N_4127,N_4128,N_4130,N_4131,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4152,N_4153,N_4154,N_4156,N_4157,N_4158,N_4159,N_4161,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4170,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4182,N_4183,N_4184,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4215,N_4216,N_4217,N_4218,N_4219,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4228,N_4229,N_4230,N_4231,N_4233,N_4234,N_4235,N_4236,N_4238,N_4239,N_4241,N_4242,N_4245,N_4246,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4262,N_4263,N_4266,N_4267,N_4268,N_4269,N_4270,N_4272,N_4273,N_4275,N_4276,N_4277,N_4278,N_4279,N_4281,N_4282,N_4283,N_4285,N_4286,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4315,N_4316,N_4317,N_4318,N_4319,N_4321,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4344,N_4345,N_4348,N_4349,N_4350,N_4352,N_4353,N_4355,N_4357,N_4358,N_4359,N_4360,N_4361,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4377,N_4379,N_4380,N_4381,N_4382,N_4385,N_4387,N_4388,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4407,N_4408,N_4409,N_4410,N_4411,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4429,N_4431,N_4432,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4442,N_4443,N_4444,N_4445,N_4448,N_4449,N_4450,N_4451,N_4452,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4472,N_4473,N_4474,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4496,N_4497,N_4498,N_4499,N_4501,N_4503,N_4504,N_4505,N_4508,N_4509,N_4510,N_4513,N_4514,N_4515,N_4516,N_4517,N_4519,N_4520,N_4521,N_4523,N_4524,N_4525,N_4526,N_4529,N_4530,N_4531,N_4532,N_4533,N_4535,N_4536,N_4537,N_4538,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4548,N_4549,N_4550,N_4552,N_4554,N_4555,N_4557,N_4558,N_4559,N_4560,N_4561,N_4563,N_4565,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4624,N_4626,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4639,N_4640,N_4642,N_4643,N_4644,N_4645,N_4646,N_4649,N_4650,N_4651,N_4652,N_4653,N_4655,N_4656,N_4657,N_4658,N_4660,N_4662,N_4664,N_4665,N_4666,N_4667,N_4669,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4691,N_4692,N_4693,N_4695,N_4696,N_4697,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4708,N_4709,N_4711,N_4712,N_4714,N_4715,N_4716,N_4717,N_4719,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4752,N_4753,N_4754,N_4755,N_4756,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4773,N_4774,N_4775,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4801,N_4802,N_4803,N_4804,N_4807,N_4808,N_4810,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4824,N_4825,N_4826,N_4828,N_4829,N_4830,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4843,N_4846,N_4847,N_4849,N_4851,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4862,N_4864,N_4865,N_4866,N_4867,N_4868,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4878,N_4880,N_4882,N_4883,N_4884,N_4885,N_4886,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4902,N_4904,N_4906,N_4908,N_4909,N_4910,N_4911,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4923,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4944,N_4946,N_4947,N_4948,N_4949,N_4950,N_4952,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4980,N_4982,N_4983,N_4984,N_4986,N_4987,N_4988,N_4990,N_4991,N_4992,N_4993,N_4995,N_4996,N_4997,N_4998;
nand U0 (N_0,In_134,In_124);
nor U1 (N_1,In_412,In_709);
and U2 (N_2,In_555,In_644);
nand U3 (N_3,In_117,In_546);
and U4 (N_4,In_172,In_460);
or U5 (N_5,In_461,In_59);
nor U6 (N_6,In_469,In_83);
and U7 (N_7,In_636,In_20);
or U8 (N_8,In_231,In_748);
xnor U9 (N_9,In_501,In_122);
or U10 (N_10,In_150,In_384);
nand U11 (N_11,In_549,In_648);
or U12 (N_12,In_380,In_151);
or U13 (N_13,In_545,In_726);
nand U14 (N_14,In_429,In_49);
xor U15 (N_15,In_656,In_670);
and U16 (N_16,In_586,In_686);
xor U17 (N_17,In_200,In_326);
nand U18 (N_18,In_10,In_374);
and U19 (N_19,In_19,In_133);
xor U20 (N_20,In_320,In_746);
nand U21 (N_21,In_189,In_17);
xnor U22 (N_22,In_599,In_243);
nor U23 (N_23,In_417,In_728);
nor U24 (N_24,In_332,In_74);
nor U25 (N_25,In_287,In_46);
or U26 (N_26,In_107,In_705);
and U27 (N_27,In_249,In_732);
nor U28 (N_28,In_93,In_439);
or U29 (N_29,In_588,In_258);
or U30 (N_30,In_94,In_527);
or U31 (N_31,In_508,In_330);
or U32 (N_32,In_671,In_111);
and U33 (N_33,In_254,In_470);
nor U34 (N_34,In_323,In_227);
and U35 (N_35,In_259,In_196);
nor U36 (N_36,In_431,In_281);
and U37 (N_37,In_197,In_472);
and U38 (N_38,In_474,In_95);
nor U39 (N_39,In_698,In_727);
nor U40 (N_40,In_625,In_136);
nor U41 (N_41,In_414,In_687);
nor U42 (N_42,In_2,In_445);
xor U43 (N_43,In_168,In_140);
nand U44 (N_44,In_657,In_264);
and U45 (N_45,In_403,In_525);
nor U46 (N_46,In_145,In_542);
or U47 (N_47,In_738,In_115);
or U48 (N_48,In_580,In_740);
nand U49 (N_49,In_576,In_9);
or U50 (N_50,In_365,In_430);
or U51 (N_51,In_560,In_317);
or U52 (N_52,In_4,In_554);
nand U53 (N_53,In_314,In_118);
and U54 (N_54,In_604,In_250);
or U55 (N_55,In_483,In_295);
nand U56 (N_56,In_719,In_516);
nand U57 (N_57,In_399,In_99);
and U58 (N_58,In_669,In_362);
or U59 (N_59,In_477,In_366);
nand U60 (N_60,In_611,In_342);
nor U61 (N_61,In_98,In_225);
nand U62 (N_62,In_171,In_275);
nor U63 (N_63,In_324,In_574);
and U64 (N_64,In_462,In_106);
and U65 (N_65,In_504,In_480);
nor U66 (N_66,In_497,In_658);
or U67 (N_67,In_663,In_531);
nor U68 (N_68,In_419,In_128);
or U69 (N_69,In_22,In_188);
nand U70 (N_70,In_206,In_379);
or U71 (N_71,In_742,In_708);
and U72 (N_72,In_63,In_421);
nor U73 (N_73,In_293,In_103);
nor U74 (N_74,In_194,In_593);
xnor U75 (N_75,In_487,In_48);
nand U76 (N_76,In_210,In_597);
xnor U77 (N_77,In_603,In_540);
nand U78 (N_78,In_5,In_32);
nand U79 (N_79,In_695,In_340);
nor U80 (N_80,In_596,In_486);
nand U81 (N_81,In_68,In_302);
and U82 (N_82,In_494,In_616);
nor U83 (N_83,In_169,In_442);
or U84 (N_84,In_266,In_343);
and U85 (N_85,In_325,In_334);
nand U86 (N_86,In_488,In_450);
nor U87 (N_87,In_251,In_521);
xor U88 (N_88,In_587,In_52);
or U89 (N_89,In_289,In_58);
nor U90 (N_90,In_24,In_637);
nand U91 (N_91,In_211,In_711);
or U92 (N_92,In_731,In_363);
nand U93 (N_93,In_256,In_524);
nand U94 (N_94,In_143,In_680);
and U95 (N_95,In_561,In_413);
nor U96 (N_96,In_141,In_290);
nand U97 (N_97,In_244,In_237);
or U98 (N_98,In_396,In_18);
and U99 (N_99,In_535,In_675);
nand U100 (N_100,In_185,In_602);
and U101 (N_101,In_204,In_14);
and U102 (N_102,In_224,In_267);
nor U103 (N_103,In_659,In_473);
nor U104 (N_104,In_162,In_255);
nor U105 (N_105,In_406,In_393);
nand U106 (N_106,In_350,In_427);
xnor U107 (N_107,In_515,In_81);
or U108 (N_108,In_548,In_154);
or U109 (N_109,In_617,In_454);
nand U110 (N_110,In_411,In_667);
and U111 (N_111,In_674,In_31);
nor U112 (N_112,In_8,In_282);
nand U113 (N_113,In_329,In_492);
nand U114 (N_114,In_21,In_736);
and U115 (N_115,In_579,In_205);
and U116 (N_116,In_352,In_62);
nor U117 (N_117,In_405,In_730);
and U118 (N_118,In_43,In_433);
nand U119 (N_119,In_386,In_92);
or U120 (N_120,In_533,In_1);
and U121 (N_121,In_436,In_50);
nand U122 (N_122,In_56,In_166);
and U123 (N_123,In_685,In_621);
and U124 (N_124,In_218,In_743);
nand U125 (N_125,In_739,In_184);
nand U126 (N_126,In_131,In_688);
and U127 (N_127,In_212,In_319);
or U128 (N_128,In_90,In_35);
xnor U129 (N_129,In_163,In_191);
nand U130 (N_130,In_679,In_485);
xor U131 (N_131,In_38,In_410);
nor U132 (N_132,In_66,In_353);
or U133 (N_133,In_517,In_110);
nand U134 (N_134,In_394,In_130);
nor U135 (N_135,In_539,In_645);
and U136 (N_136,In_214,In_236);
or U137 (N_137,In_327,In_369);
or U138 (N_138,In_407,In_64);
or U139 (N_139,In_400,In_39);
or U140 (N_140,In_553,In_228);
xnor U141 (N_141,In_82,In_271);
and U142 (N_142,In_344,In_478);
xor U143 (N_143,In_720,In_567);
and U144 (N_144,In_121,In_747);
and U145 (N_145,In_677,In_672);
nor U146 (N_146,In_312,In_335);
nand U147 (N_147,In_502,In_724);
nor U148 (N_148,In_370,In_459);
or U149 (N_149,In_345,In_159);
and U150 (N_150,In_397,In_89);
or U151 (N_151,In_272,In_591);
nand U152 (N_152,In_428,In_543);
nor U153 (N_153,In_479,In_457);
nand U154 (N_154,In_498,In_594);
or U155 (N_155,In_717,In_499);
and U156 (N_156,In_467,In_507);
nand U157 (N_157,In_707,In_618);
nand U158 (N_158,In_661,In_590);
and U159 (N_159,In_676,In_284);
or U160 (N_160,In_125,In_630);
nand U161 (N_161,In_186,In_139);
or U162 (N_162,In_360,In_41);
or U163 (N_163,In_349,In_104);
nand U164 (N_164,In_565,In_437);
nor U165 (N_165,In_181,In_148);
xor U166 (N_166,In_142,In_577);
or U167 (N_167,In_426,In_313);
and U168 (N_168,In_744,In_311);
and U169 (N_169,In_67,In_526);
xor U170 (N_170,In_368,In_699);
nand U171 (N_171,In_605,In_649);
nand U172 (N_172,In_514,In_226);
xnor U173 (N_173,In_322,In_265);
nand U174 (N_174,In_650,In_468);
and U175 (N_175,In_633,In_338);
and U176 (N_176,In_598,In_192);
nor U177 (N_177,In_615,In_532);
and U178 (N_178,In_600,In_547);
nor U179 (N_179,In_190,In_519);
and U180 (N_180,In_372,In_202);
or U181 (N_181,In_511,In_57);
nand U182 (N_182,In_690,In_199);
and U183 (N_183,In_96,In_29);
nor U184 (N_184,In_383,In_627);
and U185 (N_185,In_180,In_456);
nor U186 (N_186,In_47,In_253);
nor U187 (N_187,In_176,In_129);
nor U188 (N_188,In_109,In_174);
or U189 (N_189,In_203,In_215);
or U190 (N_190,In_377,In_376);
nand U191 (N_191,In_438,In_595);
nor U192 (N_192,In_443,In_299);
nand U193 (N_193,In_167,In_309);
nor U194 (N_194,In_713,In_348);
nor U195 (N_195,In_449,In_51);
nor U196 (N_196,In_232,In_308);
and U197 (N_197,In_61,In_120);
and U198 (N_198,In_425,In_239);
nor U199 (N_199,In_357,In_476);
nor U200 (N_200,In_321,In_77);
or U201 (N_201,In_655,In_528);
nand U202 (N_202,In_700,In_513);
xor U203 (N_203,In_359,In_571);
xnor U204 (N_204,In_161,In_222);
or U205 (N_205,In_155,In_355);
or U206 (N_206,In_569,In_512);
or U207 (N_207,In_55,In_337);
and U208 (N_208,In_0,In_704);
and U209 (N_209,In_635,In_356);
or U210 (N_210,In_187,In_714);
xor U211 (N_211,In_570,In_173);
nor U212 (N_212,In_294,In_651);
or U213 (N_213,In_375,In_273);
nand U214 (N_214,In_105,In_398);
or U215 (N_215,In_354,In_100);
or U216 (N_216,In_440,In_16);
nand U217 (N_217,In_71,In_69);
or U218 (N_218,In_13,In_135);
and U219 (N_219,In_296,In_453);
xor U220 (N_220,In_292,In_606);
nand U221 (N_221,In_722,In_36);
nand U222 (N_222,In_706,In_522);
and U223 (N_223,In_248,In_182);
nand U224 (N_224,In_609,In_91);
or U225 (N_225,In_592,In_614);
nor U226 (N_226,In_446,In_691);
and U227 (N_227,In_219,In_529);
nor U228 (N_228,In_114,In_471);
nor U229 (N_229,In_652,In_568);
nor U230 (N_230,In_523,In_33);
nor U231 (N_231,In_475,In_581);
xnor U232 (N_232,In_518,In_156);
nand U233 (N_233,In_392,In_87);
nand U234 (N_234,In_378,In_631);
nor U235 (N_235,In_654,In_364);
nor U236 (N_236,In_583,In_402);
nand U237 (N_237,In_358,In_391);
nor U238 (N_238,In_116,In_164);
and U239 (N_239,In_245,In_307);
xor U240 (N_240,In_252,In_213);
and U241 (N_241,In_298,In_119);
or U242 (N_242,In_703,In_170);
or U243 (N_243,In_573,In_144);
and U244 (N_244,In_268,In_333);
and U245 (N_245,In_640,In_733);
nor U246 (N_246,In_276,In_389);
xor U247 (N_247,In_341,In_367);
nor U248 (N_248,In_158,In_315);
nor U249 (N_249,In_318,In_660);
and U250 (N_250,In_301,In_589);
nand U251 (N_251,In_647,In_278);
or U252 (N_252,In_584,In_261);
and U253 (N_253,In_387,In_336);
nor U254 (N_254,In_666,In_84);
nand U255 (N_255,In_361,In_534);
or U256 (N_256,In_506,In_7);
and U257 (N_257,In_628,In_683);
nor U258 (N_258,In_79,In_132);
nor U259 (N_259,In_493,In_613);
xnor U260 (N_260,In_496,In_220);
or U261 (N_261,In_388,In_612);
nand U262 (N_262,In_316,In_435);
nand U263 (N_263,In_424,In_701);
or U264 (N_264,In_85,In_557);
nand U265 (N_265,In_238,In_601);
and U266 (N_266,In_73,In_716);
and U267 (N_267,In_702,In_490);
nand U268 (N_268,In_37,In_97);
or U269 (N_269,In_664,In_72);
and U270 (N_270,In_734,In_585);
and U271 (N_271,In_65,In_277);
nor U272 (N_272,In_138,In_70);
nor U273 (N_273,In_416,In_44);
xnor U274 (N_274,In_217,In_422);
nand U275 (N_275,In_30,In_195);
and U276 (N_276,In_575,In_102);
nor U277 (N_277,In_694,In_233);
xnor U278 (N_278,In_390,In_432);
and U279 (N_279,In_420,In_668);
nor U280 (N_280,In_622,In_149);
and U281 (N_281,In_452,In_160);
nand U282 (N_282,In_112,In_274);
or U283 (N_283,In_88,In_749);
and U284 (N_284,In_305,In_626);
xor U285 (N_285,In_444,In_34);
or U286 (N_286,In_455,In_381);
nand U287 (N_287,In_608,In_263);
nor U288 (N_288,In_578,In_489);
nand U289 (N_289,In_165,In_418);
or U290 (N_290,In_157,In_193);
nor U291 (N_291,In_234,In_28);
or U292 (N_292,In_551,In_536);
or U293 (N_293,In_491,In_544);
and U294 (N_294,In_441,In_619);
and U295 (N_295,In_715,In_642);
nand U296 (N_296,In_395,In_347);
or U297 (N_297,In_198,In_481);
and U298 (N_298,In_623,In_415);
and U299 (N_299,In_328,In_288);
and U300 (N_300,In_241,In_710);
nor U301 (N_301,In_505,In_297);
nand U302 (N_302,In_404,In_247);
and U303 (N_303,In_175,In_146);
nand U304 (N_304,In_530,In_303);
and U305 (N_305,In_42,In_152);
nor U306 (N_306,In_566,In_673);
or U307 (N_307,In_351,In_270);
xor U308 (N_308,In_286,In_76);
xor U309 (N_309,In_484,In_306);
or U310 (N_310,In_464,In_183);
nand U311 (N_311,In_653,In_283);
nor U312 (N_312,In_6,In_25);
xor U313 (N_313,In_86,In_280);
nand U314 (N_314,In_482,In_27);
and U315 (N_315,In_629,In_563);
nor U316 (N_316,In_279,In_382);
or U317 (N_317,In_610,In_147);
nor U318 (N_318,In_53,In_201);
or U319 (N_319,In_127,In_696);
or U320 (N_320,In_643,In_209);
nand U321 (N_321,In_681,In_221);
and U322 (N_322,In_291,In_54);
nand U323 (N_323,In_538,In_285);
nor U324 (N_324,In_463,In_447);
or U325 (N_325,In_451,In_684);
and U326 (N_326,In_207,In_624);
nor U327 (N_327,In_385,In_556);
nand U328 (N_328,In_723,In_646);
nand U329 (N_329,In_208,In_409);
or U330 (N_330,In_745,In_178);
or U331 (N_331,In_269,In_510);
xnor U332 (N_332,In_26,In_113);
nand U333 (N_333,In_45,In_620);
or U334 (N_334,In_262,In_634);
and U335 (N_335,In_371,In_257);
and U336 (N_336,In_235,In_466);
or U337 (N_337,In_331,In_310);
and U338 (N_338,In_500,In_725);
and U339 (N_339,In_692,In_108);
nand U340 (N_340,In_718,In_559);
nand U341 (N_341,In_177,In_582);
nand U342 (N_342,In_552,In_665);
nor U343 (N_343,In_520,In_80);
or U344 (N_344,In_509,In_300);
and U345 (N_345,In_662,In_423);
nand U346 (N_346,In_179,In_246);
xnor U347 (N_347,In_401,In_737);
and U348 (N_348,In_741,In_458);
and U349 (N_349,In_465,In_101);
nand U350 (N_350,In_712,In_15);
and U351 (N_351,In_223,In_541);
and U352 (N_352,In_641,In_260);
or U353 (N_353,In_12,In_721);
and U354 (N_354,In_448,In_242);
or U355 (N_355,In_729,In_689);
nor U356 (N_356,In_216,In_564);
and U357 (N_357,In_346,In_607);
or U358 (N_358,In_503,In_693);
xnor U359 (N_359,In_339,In_373);
or U360 (N_360,In_229,In_40);
nand U361 (N_361,In_697,In_60);
or U362 (N_362,In_682,In_240);
xnor U363 (N_363,In_558,In_408);
and U364 (N_364,In_126,In_735);
or U365 (N_365,In_562,In_638);
and U366 (N_366,In_632,In_537);
or U367 (N_367,In_550,In_137);
and U368 (N_368,In_123,In_572);
nand U369 (N_369,In_153,In_678);
and U370 (N_370,In_3,In_75);
nor U371 (N_371,In_639,In_230);
nand U372 (N_372,In_304,In_78);
nand U373 (N_373,In_434,In_495);
nand U374 (N_374,In_23,In_11);
nand U375 (N_375,In_497,In_623);
xnor U376 (N_376,In_202,In_242);
or U377 (N_377,In_387,In_90);
nor U378 (N_378,In_584,In_592);
and U379 (N_379,In_725,In_551);
nand U380 (N_380,In_93,In_641);
nand U381 (N_381,In_408,In_705);
or U382 (N_382,In_732,In_222);
xnor U383 (N_383,In_370,In_485);
nand U384 (N_384,In_330,In_506);
or U385 (N_385,In_87,In_150);
nor U386 (N_386,In_582,In_425);
or U387 (N_387,In_237,In_360);
or U388 (N_388,In_604,In_405);
nand U389 (N_389,In_170,In_143);
nand U390 (N_390,In_738,In_654);
xnor U391 (N_391,In_391,In_694);
nand U392 (N_392,In_36,In_426);
nor U393 (N_393,In_646,In_251);
nor U394 (N_394,In_241,In_386);
or U395 (N_395,In_475,In_48);
nand U396 (N_396,In_177,In_246);
or U397 (N_397,In_308,In_209);
nand U398 (N_398,In_112,In_474);
nor U399 (N_399,In_739,In_387);
nor U400 (N_400,In_158,In_711);
nand U401 (N_401,In_660,In_440);
nand U402 (N_402,In_529,In_306);
or U403 (N_403,In_480,In_45);
nand U404 (N_404,In_95,In_283);
or U405 (N_405,In_306,In_734);
or U406 (N_406,In_8,In_609);
nand U407 (N_407,In_650,In_71);
nand U408 (N_408,In_655,In_710);
or U409 (N_409,In_677,In_405);
or U410 (N_410,In_46,In_377);
and U411 (N_411,In_713,In_410);
xor U412 (N_412,In_207,In_5);
and U413 (N_413,In_666,In_561);
and U414 (N_414,In_387,In_569);
nand U415 (N_415,In_340,In_124);
xnor U416 (N_416,In_572,In_437);
nor U417 (N_417,In_124,In_481);
and U418 (N_418,In_307,In_303);
or U419 (N_419,In_479,In_246);
nand U420 (N_420,In_745,In_588);
nor U421 (N_421,In_250,In_152);
nand U422 (N_422,In_370,In_683);
or U423 (N_423,In_550,In_394);
or U424 (N_424,In_74,In_204);
or U425 (N_425,In_333,In_468);
nand U426 (N_426,In_30,In_610);
and U427 (N_427,In_713,In_724);
and U428 (N_428,In_584,In_489);
and U429 (N_429,In_335,In_559);
xnor U430 (N_430,In_385,In_270);
or U431 (N_431,In_469,In_245);
and U432 (N_432,In_56,In_496);
and U433 (N_433,In_476,In_498);
xor U434 (N_434,In_452,In_240);
or U435 (N_435,In_236,In_30);
and U436 (N_436,In_41,In_223);
or U437 (N_437,In_612,In_574);
and U438 (N_438,In_74,In_185);
or U439 (N_439,In_742,In_51);
nor U440 (N_440,In_453,In_709);
xor U441 (N_441,In_23,In_739);
or U442 (N_442,In_640,In_525);
or U443 (N_443,In_522,In_238);
or U444 (N_444,In_196,In_24);
and U445 (N_445,In_258,In_287);
or U446 (N_446,In_320,In_405);
or U447 (N_447,In_64,In_264);
xnor U448 (N_448,In_313,In_287);
nor U449 (N_449,In_730,In_192);
nor U450 (N_450,In_21,In_673);
nand U451 (N_451,In_294,In_81);
nor U452 (N_452,In_349,In_70);
or U453 (N_453,In_43,In_36);
and U454 (N_454,In_536,In_569);
xnor U455 (N_455,In_593,In_481);
xnor U456 (N_456,In_635,In_90);
xor U457 (N_457,In_432,In_538);
and U458 (N_458,In_332,In_449);
xnor U459 (N_459,In_94,In_88);
or U460 (N_460,In_157,In_524);
and U461 (N_461,In_499,In_234);
or U462 (N_462,In_144,In_682);
nor U463 (N_463,In_288,In_14);
or U464 (N_464,In_388,In_420);
nand U465 (N_465,In_467,In_228);
nand U466 (N_466,In_389,In_354);
or U467 (N_467,In_527,In_617);
or U468 (N_468,In_556,In_600);
and U469 (N_469,In_308,In_705);
or U470 (N_470,In_741,In_366);
or U471 (N_471,In_55,In_502);
nor U472 (N_472,In_175,In_483);
and U473 (N_473,In_727,In_401);
xnor U474 (N_474,In_162,In_611);
or U475 (N_475,In_731,In_396);
nand U476 (N_476,In_198,In_628);
xnor U477 (N_477,In_356,In_161);
nor U478 (N_478,In_245,In_340);
nor U479 (N_479,In_343,In_461);
and U480 (N_480,In_5,In_291);
and U481 (N_481,In_687,In_626);
or U482 (N_482,In_676,In_460);
nand U483 (N_483,In_729,In_714);
nand U484 (N_484,In_696,In_29);
or U485 (N_485,In_689,In_67);
or U486 (N_486,In_392,In_247);
nor U487 (N_487,In_662,In_455);
nand U488 (N_488,In_143,In_209);
nor U489 (N_489,In_274,In_464);
and U490 (N_490,In_83,In_247);
or U491 (N_491,In_685,In_130);
nand U492 (N_492,In_315,In_709);
or U493 (N_493,In_310,In_367);
and U494 (N_494,In_156,In_720);
and U495 (N_495,In_250,In_187);
or U496 (N_496,In_463,In_374);
or U497 (N_497,In_736,In_174);
nor U498 (N_498,In_614,In_639);
xnor U499 (N_499,In_145,In_179);
and U500 (N_500,In_322,In_721);
nor U501 (N_501,In_447,In_527);
xor U502 (N_502,In_534,In_442);
and U503 (N_503,In_23,In_467);
or U504 (N_504,In_229,In_459);
and U505 (N_505,In_714,In_479);
and U506 (N_506,In_449,In_280);
and U507 (N_507,In_699,In_134);
nor U508 (N_508,In_247,In_158);
or U509 (N_509,In_692,In_50);
nand U510 (N_510,In_581,In_483);
nor U511 (N_511,In_599,In_272);
or U512 (N_512,In_60,In_64);
xnor U513 (N_513,In_182,In_395);
nor U514 (N_514,In_236,In_176);
and U515 (N_515,In_227,In_628);
and U516 (N_516,In_657,In_664);
or U517 (N_517,In_334,In_104);
and U518 (N_518,In_401,In_652);
nor U519 (N_519,In_193,In_498);
nand U520 (N_520,In_379,In_483);
nor U521 (N_521,In_104,In_673);
or U522 (N_522,In_218,In_326);
and U523 (N_523,In_79,In_173);
nand U524 (N_524,In_469,In_217);
nor U525 (N_525,In_271,In_675);
nor U526 (N_526,In_296,In_153);
and U527 (N_527,In_700,In_746);
nor U528 (N_528,In_619,In_56);
and U529 (N_529,In_279,In_615);
nor U530 (N_530,In_176,In_486);
and U531 (N_531,In_577,In_597);
nor U532 (N_532,In_94,In_22);
or U533 (N_533,In_84,In_364);
and U534 (N_534,In_125,In_691);
or U535 (N_535,In_159,In_733);
and U536 (N_536,In_227,In_660);
xnor U537 (N_537,In_462,In_309);
xnor U538 (N_538,In_513,In_473);
and U539 (N_539,In_105,In_35);
or U540 (N_540,In_686,In_50);
and U541 (N_541,In_247,In_638);
or U542 (N_542,In_580,In_630);
nor U543 (N_543,In_0,In_377);
or U544 (N_544,In_357,In_571);
or U545 (N_545,In_575,In_156);
nand U546 (N_546,In_291,In_129);
xnor U547 (N_547,In_147,In_433);
and U548 (N_548,In_261,In_146);
or U549 (N_549,In_692,In_2);
nand U550 (N_550,In_497,In_196);
or U551 (N_551,In_248,In_654);
and U552 (N_552,In_289,In_441);
and U553 (N_553,In_554,In_21);
nor U554 (N_554,In_392,In_228);
nand U555 (N_555,In_77,In_24);
nand U556 (N_556,In_293,In_687);
nand U557 (N_557,In_749,In_656);
nor U558 (N_558,In_577,In_316);
or U559 (N_559,In_2,In_214);
or U560 (N_560,In_516,In_251);
xor U561 (N_561,In_16,In_749);
xor U562 (N_562,In_274,In_736);
nor U563 (N_563,In_266,In_198);
and U564 (N_564,In_269,In_525);
nand U565 (N_565,In_297,In_628);
nor U566 (N_566,In_744,In_30);
or U567 (N_567,In_381,In_608);
nor U568 (N_568,In_225,In_332);
or U569 (N_569,In_392,In_749);
nand U570 (N_570,In_587,In_73);
nor U571 (N_571,In_454,In_512);
nor U572 (N_572,In_217,In_568);
and U573 (N_573,In_604,In_742);
and U574 (N_574,In_17,In_286);
nand U575 (N_575,In_32,In_589);
nand U576 (N_576,In_572,In_501);
or U577 (N_577,In_36,In_498);
or U578 (N_578,In_279,In_516);
and U579 (N_579,In_222,In_60);
nor U580 (N_580,In_490,In_58);
or U581 (N_581,In_260,In_348);
or U582 (N_582,In_610,In_730);
and U583 (N_583,In_248,In_275);
or U584 (N_584,In_280,In_195);
nor U585 (N_585,In_736,In_546);
or U586 (N_586,In_460,In_429);
and U587 (N_587,In_110,In_508);
and U588 (N_588,In_6,In_522);
or U589 (N_589,In_746,In_12);
or U590 (N_590,In_230,In_384);
or U591 (N_591,In_548,In_590);
nand U592 (N_592,In_292,In_210);
and U593 (N_593,In_410,In_71);
or U594 (N_594,In_454,In_258);
nor U595 (N_595,In_427,In_117);
nor U596 (N_596,In_64,In_179);
and U597 (N_597,In_441,In_429);
nand U598 (N_598,In_307,In_528);
xor U599 (N_599,In_579,In_318);
or U600 (N_600,In_145,In_731);
or U601 (N_601,In_621,In_96);
nand U602 (N_602,In_686,In_409);
and U603 (N_603,In_390,In_186);
nand U604 (N_604,In_221,In_367);
or U605 (N_605,In_656,In_275);
and U606 (N_606,In_664,In_112);
nor U607 (N_607,In_81,In_137);
nand U608 (N_608,In_672,In_716);
xor U609 (N_609,In_203,In_691);
nor U610 (N_610,In_579,In_134);
or U611 (N_611,In_662,In_204);
nand U612 (N_612,In_566,In_552);
nand U613 (N_613,In_688,In_0);
xor U614 (N_614,In_261,In_58);
xor U615 (N_615,In_226,In_270);
or U616 (N_616,In_458,In_544);
and U617 (N_617,In_275,In_426);
nand U618 (N_618,In_318,In_479);
xor U619 (N_619,In_741,In_680);
nor U620 (N_620,In_490,In_602);
nor U621 (N_621,In_63,In_654);
xor U622 (N_622,In_485,In_89);
or U623 (N_623,In_263,In_75);
and U624 (N_624,In_156,In_158);
and U625 (N_625,In_683,In_61);
nand U626 (N_626,In_341,In_75);
and U627 (N_627,In_178,In_30);
nor U628 (N_628,In_239,In_665);
and U629 (N_629,In_245,In_232);
and U630 (N_630,In_316,In_544);
nor U631 (N_631,In_367,In_475);
nand U632 (N_632,In_727,In_719);
nand U633 (N_633,In_638,In_651);
nand U634 (N_634,In_575,In_576);
or U635 (N_635,In_18,In_443);
nor U636 (N_636,In_218,In_553);
nand U637 (N_637,In_542,In_78);
nor U638 (N_638,In_24,In_55);
nand U639 (N_639,In_136,In_590);
nand U640 (N_640,In_47,In_697);
nor U641 (N_641,In_510,In_663);
nand U642 (N_642,In_552,In_572);
nor U643 (N_643,In_304,In_544);
and U644 (N_644,In_233,In_64);
nand U645 (N_645,In_694,In_312);
nor U646 (N_646,In_336,In_685);
or U647 (N_647,In_659,In_353);
nor U648 (N_648,In_638,In_503);
nand U649 (N_649,In_202,In_138);
and U650 (N_650,In_414,In_589);
xor U651 (N_651,In_707,In_546);
nor U652 (N_652,In_672,In_231);
and U653 (N_653,In_387,In_164);
and U654 (N_654,In_482,In_532);
and U655 (N_655,In_610,In_21);
nor U656 (N_656,In_443,In_539);
nor U657 (N_657,In_290,In_435);
nor U658 (N_658,In_532,In_66);
nand U659 (N_659,In_261,In_558);
or U660 (N_660,In_109,In_183);
nor U661 (N_661,In_533,In_608);
nor U662 (N_662,In_468,In_413);
nand U663 (N_663,In_353,In_550);
and U664 (N_664,In_416,In_726);
nor U665 (N_665,In_173,In_529);
xor U666 (N_666,In_498,In_502);
xor U667 (N_667,In_39,In_169);
nor U668 (N_668,In_109,In_590);
xor U669 (N_669,In_280,In_380);
nand U670 (N_670,In_252,In_381);
xor U671 (N_671,In_440,In_350);
nor U672 (N_672,In_361,In_191);
nor U673 (N_673,In_595,In_193);
or U674 (N_674,In_488,In_434);
or U675 (N_675,In_401,In_518);
nor U676 (N_676,In_594,In_244);
nor U677 (N_677,In_54,In_415);
nand U678 (N_678,In_523,In_528);
nor U679 (N_679,In_117,In_534);
and U680 (N_680,In_519,In_545);
or U681 (N_681,In_43,In_473);
or U682 (N_682,In_429,In_589);
nor U683 (N_683,In_725,In_215);
and U684 (N_684,In_384,In_209);
or U685 (N_685,In_482,In_550);
or U686 (N_686,In_7,In_270);
or U687 (N_687,In_186,In_434);
nand U688 (N_688,In_104,In_627);
xor U689 (N_689,In_746,In_134);
nand U690 (N_690,In_124,In_373);
nor U691 (N_691,In_27,In_330);
nor U692 (N_692,In_283,In_184);
or U693 (N_693,In_40,In_367);
nor U694 (N_694,In_114,In_720);
or U695 (N_695,In_662,In_178);
and U696 (N_696,In_682,In_719);
and U697 (N_697,In_529,In_619);
or U698 (N_698,In_131,In_672);
nand U699 (N_699,In_56,In_645);
or U700 (N_700,In_621,In_184);
or U701 (N_701,In_555,In_454);
and U702 (N_702,In_169,In_513);
or U703 (N_703,In_707,In_399);
and U704 (N_704,In_596,In_635);
nor U705 (N_705,In_330,In_266);
xnor U706 (N_706,In_552,In_159);
nand U707 (N_707,In_734,In_346);
nand U708 (N_708,In_480,In_70);
and U709 (N_709,In_673,In_373);
or U710 (N_710,In_553,In_170);
nand U711 (N_711,In_580,In_309);
nand U712 (N_712,In_28,In_7);
nor U713 (N_713,In_234,In_348);
and U714 (N_714,In_269,In_306);
nand U715 (N_715,In_258,In_678);
nor U716 (N_716,In_548,In_243);
nor U717 (N_717,In_408,In_550);
or U718 (N_718,In_688,In_625);
and U719 (N_719,In_75,In_627);
nor U720 (N_720,In_271,In_32);
and U721 (N_721,In_572,In_253);
and U722 (N_722,In_10,In_340);
nor U723 (N_723,In_608,In_30);
or U724 (N_724,In_561,In_509);
nand U725 (N_725,In_644,In_361);
and U726 (N_726,In_160,In_165);
nor U727 (N_727,In_443,In_120);
nand U728 (N_728,In_275,In_450);
nand U729 (N_729,In_657,In_247);
xor U730 (N_730,In_529,In_257);
nand U731 (N_731,In_548,In_50);
nand U732 (N_732,In_236,In_10);
nor U733 (N_733,In_494,In_673);
or U734 (N_734,In_652,In_623);
nor U735 (N_735,In_237,In_579);
xnor U736 (N_736,In_664,In_547);
nand U737 (N_737,In_480,In_197);
nand U738 (N_738,In_356,In_171);
and U739 (N_739,In_85,In_289);
or U740 (N_740,In_642,In_381);
nor U741 (N_741,In_686,In_208);
nor U742 (N_742,In_657,In_432);
nor U743 (N_743,In_690,In_378);
nand U744 (N_744,In_405,In_433);
or U745 (N_745,In_157,In_547);
nor U746 (N_746,In_622,In_560);
and U747 (N_747,In_536,In_64);
or U748 (N_748,In_403,In_740);
or U749 (N_749,In_257,In_645);
and U750 (N_750,In_648,In_485);
nand U751 (N_751,In_130,In_68);
nand U752 (N_752,In_449,In_714);
nand U753 (N_753,In_239,In_476);
and U754 (N_754,In_110,In_547);
xor U755 (N_755,In_677,In_697);
nand U756 (N_756,In_242,In_98);
or U757 (N_757,In_518,In_116);
and U758 (N_758,In_450,In_318);
and U759 (N_759,In_280,In_641);
and U760 (N_760,In_381,In_177);
and U761 (N_761,In_1,In_625);
or U762 (N_762,In_408,In_269);
nor U763 (N_763,In_695,In_60);
nand U764 (N_764,In_32,In_204);
and U765 (N_765,In_227,In_368);
nand U766 (N_766,In_61,In_665);
or U767 (N_767,In_548,In_734);
nor U768 (N_768,In_381,In_509);
nor U769 (N_769,In_673,In_700);
or U770 (N_770,In_303,In_317);
and U771 (N_771,In_562,In_360);
nor U772 (N_772,In_306,In_335);
xnor U773 (N_773,In_177,In_368);
nand U774 (N_774,In_235,In_5);
xor U775 (N_775,In_6,In_162);
nand U776 (N_776,In_628,In_130);
or U777 (N_777,In_349,In_451);
and U778 (N_778,In_40,In_636);
or U779 (N_779,In_414,In_290);
and U780 (N_780,In_655,In_562);
nand U781 (N_781,In_269,In_20);
nor U782 (N_782,In_664,In_353);
or U783 (N_783,In_242,In_119);
nor U784 (N_784,In_134,In_518);
or U785 (N_785,In_87,In_229);
or U786 (N_786,In_161,In_56);
or U787 (N_787,In_88,In_129);
and U788 (N_788,In_288,In_377);
or U789 (N_789,In_223,In_476);
xnor U790 (N_790,In_354,In_660);
or U791 (N_791,In_402,In_0);
or U792 (N_792,In_27,In_653);
xor U793 (N_793,In_28,In_626);
nor U794 (N_794,In_351,In_136);
nor U795 (N_795,In_347,In_584);
nor U796 (N_796,In_221,In_601);
and U797 (N_797,In_473,In_279);
or U798 (N_798,In_687,In_404);
or U799 (N_799,In_100,In_26);
nand U800 (N_800,In_16,In_742);
nor U801 (N_801,In_559,In_343);
nor U802 (N_802,In_657,In_116);
nor U803 (N_803,In_24,In_668);
nor U804 (N_804,In_430,In_725);
nand U805 (N_805,In_7,In_749);
or U806 (N_806,In_493,In_593);
and U807 (N_807,In_135,In_275);
nand U808 (N_808,In_591,In_734);
xor U809 (N_809,In_573,In_626);
or U810 (N_810,In_254,In_125);
or U811 (N_811,In_729,In_610);
or U812 (N_812,In_215,In_76);
nor U813 (N_813,In_50,In_536);
nor U814 (N_814,In_609,In_168);
or U815 (N_815,In_57,In_22);
or U816 (N_816,In_641,In_590);
xor U817 (N_817,In_637,In_429);
nor U818 (N_818,In_645,In_605);
nand U819 (N_819,In_441,In_408);
nand U820 (N_820,In_711,In_641);
nor U821 (N_821,In_487,In_522);
or U822 (N_822,In_228,In_50);
or U823 (N_823,In_221,In_521);
or U824 (N_824,In_17,In_282);
nor U825 (N_825,In_56,In_9);
or U826 (N_826,In_523,In_368);
nor U827 (N_827,In_345,In_577);
nor U828 (N_828,In_481,In_487);
and U829 (N_829,In_541,In_179);
or U830 (N_830,In_231,In_141);
nor U831 (N_831,In_247,In_132);
or U832 (N_832,In_280,In_678);
and U833 (N_833,In_335,In_284);
xor U834 (N_834,In_83,In_196);
nand U835 (N_835,In_556,In_311);
nand U836 (N_836,In_53,In_557);
xor U837 (N_837,In_157,In_719);
nand U838 (N_838,In_536,In_126);
nand U839 (N_839,In_362,In_606);
nand U840 (N_840,In_363,In_568);
xor U841 (N_841,In_550,In_63);
nor U842 (N_842,In_445,In_105);
and U843 (N_843,In_723,In_522);
or U844 (N_844,In_697,In_14);
nand U845 (N_845,In_688,In_510);
or U846 (N_846,In_610,In_346);
and U847 (N_847,In_425,In_519);
nand U848 (N_848,In_475,In_683);
nand U849 (N_849,In_186,In_366);
nor U850 (N_850,In_449,In_17);
nor U851 (N_851,In_543,In_104);
nor U852 (N_852,In_114,In_523);
and U853 (N_853,In_336,In_382);
nand U854 (N_854,In_278,In_631);
and U855 (N_855,In_569,In_100);
nand U856 (N_856,In_104,In_233);
and U857 (N_857,In_353,In_466);
nor U858 (N_858,In_478,In_362);
nand U859 (N_859,In_250,In_32);
and U860 (N_860,In_92,In_168);
xnor U861 (N_861,In_441,In_435);
nor U862 (N_862,In_537,In_727);
nand U863 (N_863,In_618,In_138);
xor U864 (N_864,In_32,In_728);
xnor U865 (N_865,In_544,In_114);
or U866 (N_866,In_250,In_261);
and U867 (N_867,In_490,In_68);
or U868 (N_868,In_530,In_627);
nor U869 (N_869,In_397,In_169);
nor U870 (N_870,In_703,In_264);
nor U871 (N_871,In_664,In_536);
nor U872 (N_872,In_66,In_506);
xor U873 (N_873,In_77,In_92);
nor U874 (N_874,In_734,In_437);
and U875 (N_875,In_195,In_162);
nand U876 (N_876,In_682,In_343);
or U877 (N_877,In_317,In_398);
xnor U878 (N_878,In_277,In_538);
and U879 (N_879,In_377,In_172);
nor U880 (N_880,In_309,In_450);
nand U881 (N_881,In_469,In_386);
or U882 (N_882,In_704,In_741);
nor U883 (N_883,In_515,In_44);
nor U884 (N_884,In_390,In_597);
nand U885 (N_885,In_8,In_171);
xor U886 (N_886,In_164,In_302);
nor U887 (N_887,In_537,In_1);
nor U888 (N_888,In_584,In_22);
nand U889 (N_889,In_670,In_618);
or U890 (N_890,In_595,In_357);
nand U891 (N_891,In_501,In_261);
nand U892 (N_892,In_2,In_634);
nor U893 (N_893,In_498,In_679);
nand U894 (N_894,In_649,In_620);
nand U895 (N_895,In_499,In_507);
and U896 (N_896,In_61,In_239);
and U897 (N_897,In_343,In_210);
nand U898 (N_898,In_491,In_661);
nor U899 (N_899,In_397,In_188);
or U900 (N_900,In_60,In_412);
or U901 (N_901,In_587,In_664);
and U902 (N_902,In_623,In_413);
or U903 (N_903,In_299,In_596);
nor U904 (N_904,In_459,In_274);
nand U905 (N_905,In_311,In_362);
or U906 (N_906,In_510,In_687);
nand U907 (N_907,In_10,In_567);
xor U908 (N_908,In_149,In_287);
or U909 (N_909,In_472,In_727);
nand U910 (N_910,In_358,In_668);
or U911 (N_911,In_480,In_438);
nor U912 (N_912,In_522,In_265);
xor U913 (N_913,In_667,In_624);
and U914 (N_914,In_490,In_197);
nand U915 (N_915,In_254,In_333);
nand U916 (N_916,In_419,In_342);
nor U917 (N_917,In_252,In_84);
and U918 (N_918,In_576,In_446);
nor U919 (N_919,In_378,In_581);
xnor U920 (N_920,In_618,In_716);
and U921 (N_921,In_198,In_120);
nor U922 (N_922,In_195,In_362);
xnor U923 (N_923,In_585,In_85);
nor U924 (N_924,In_151,In_655);
nand U925 (N_925,In_558,In_200);
xor U926 (N_926,In_210,In_677);
and U927 (N_927,In_658,In_110);
or U928 (N_928,In_123,In_433);
nor U929 (N_929,In_488,In_456);
nor U930 (N_930,In_101,In_36);
and U931 (N_931,In_484,In_587);
nand U932 (N_932,In_386,In_707);
nand U933 (N_933,In_423,In_208);
nor U934 (N_934,In_734,In_54);
or U935 (N_935,In_16,In_185);
or U936 (N_936,In_572,In_414);
or U937 (N_937,In_76,In_343);
or U938 (N_938,In_295,In_692);
or U939 (N_939,In_539,In_260);
nor U940 (N_940,In_252,In_495);
nor U941 (N_941,In_485,In_563);
and U942 (N_942,In_375,In_479);
and U943 (N_943,In_694,In_266);
or U944 (N_944,In_526,In_649);
nand U945 (N_945,In_675,In_11);
xor U946 (N_946,In_615,In_481);
and U947 (N_947,In_342,In_142);
xnor U948 (N_948,In_702,In_270);
nand U949 (N_949,In_386,In_539);
nand U950 (N_950,In_384,In_79);
xnor U951 (N_951,In_749,In_529);
and U952 (N_952,In_32,In_472);
nor U953 (N_953,In_351,In_91);
nand U954 (N_954,In_170,In_594);
nand U955 (N_955,In_116,In_267);
xor U956 (N_956,In_228,In_549);
nand U957 (N_957,In_463,In_310);
or U958 (N_958,In_616,In_474);
nor U959 (N_959,In_443,In_652);
or U960 (N_960,In_393,In_467);
nor U961 (N_961,In_85,In_27);
nor U962 (N_962,In_681,In_242);
and U963 (N_963,In_686,In_638);
or U964 (N_964,In_255,In_301);
nand U965 (N_965,In_614,In_538);
and U966 (N_966,In_568,In_731);
and U967 (N_967,In_194,In_288);
or U968 (N_968,In_417,In_20);
and U969 (N_969,In_57,In_353);
nand U970 (N_970,In_80,In_509);
nor U971 (N_971,In_537,In_422);
and U972 (N_972,In_309,In_625);
or U973 (N_973,In_273,In_359);
nand U974 (N_974,In_366,In_634);
nor U975 (N_975,In_422,In_625);
or U976 (N_976,In_444,In_331);
nand U977 (N_977,In_213,In_231);
nor U978 (N_978,In_289,In_630);
and U979 (N_979,In_422,In_629);
nor U980 (N_980,In_207,In_44);
nor U981 (N_981,In_650,In_311);
nor U982 (N_982,In_258,In_691);
xnor U983 (N_983,In_728,In_74);
nor U984 (N_984,In_577,In_568);
and U985 (N_985,In_235,In_747);
and U986 (N_986,In_591,In_188);
and U987 (N_987,In_611,In_383);
or U988 (N_988,In_183,In_177);
nor U989 (N_989,In_685,In_274);
and U990 (N_990,In_406,In_476);
and U991 (N_991,In_73,In_124);
or U992 (N_992,In_696,In_54);
nor U993 (N_993,In_157,In_206);
or U994 (N_994,In_95,In_290);
and U995 (N_995,In_215,In_560);
and U996 (N_996,In_218,In_37);
and U997 (N_997,In_26,In_224);
or U998 (N_998,In_470,In_656);
nor U999 (N_999,In_632,In_286);
nor U1000 (N_1000,In_236,In_729);
nor U1001 (N_1001,In_40,In_729);
and U1002 (N_1002,In_268,In_148);
and U1003 (N_1003,In_525,In_593);
and U1004 (N_1004,In_534,In_499);
and U1005 (N_1005,In_109,In_85);
xnor U1006 (N_1006,In_353,In_102);
nor U1007 (N_1007,In_147,In_646);
nor U1008 (N_1008,In_630,In_233);
or U1009 (N_1009,In_427,In_635);
xor U1010 (N_1010,In_628,In_373);
and U1011 (N_1011,In_271,In_258);
nor U1012 (N_1012,In_504,In_68);
nand U1013 (N_1013,In_58,In_408);
or U1014 (N_1014,In_333,In_392);
xor U1015 (N_1015,In_121,In_709);
or U1016 (N_1016,In_310,In_589);
nand U1017 (N_1017,In_492,In_555);
nor U1018 (N_1018,In_133,In_39);
nand U1019 (N_1019,In_55,In_68);
nor U1020 (N_1020,In_94,In_353);
nand U1021 (N_1021,In_491,In_273);
and U1022 (N_1022,In_431,In_494);
and U1023 (N_1023,In_329,In_237);
nand U1024 (N_1024,In_692,In_187);
and U1025 (N_1025,In_370,In_234);
nand U1026 (N_1026,In_396,In_357);
nor U1027 (N_1027,In_680,In_9);
nor U1028 (N_1028,In_440,In_642);
and U1029 (N_1029,In_417,In_632);
and U1030 (N_1030,In_278,In_163);
and U1031 (N_1031,In_587,In_134);
and U1032 (N_1032,In_62,In_518);
and U1033 (N_1033,In_187,In_70);
nand U1034 (N_1034,In_544,In_680);
or U1035 (N_1035,In_26,In_580);
nor U1036 (N_1036,In_87,In_368);
nand U1037 (N_1037,In_540,In_684);
and U1038 (N_1038,In_624,In_260);
nand U1039 (N_1039,In_424,In_234);
nand U1040 (N_1040,In_685,In_332);
or U1041 (N_1041,In_17,In_257);
nor U1042 (N_1042,In_673,In_625);
nand U1043 (N_1043,In_473,In_466);
nor U1044 (N_1044,In_360,In_392);
nand U1045 (N_1045,In_94,In_56);
and U1046 (N_1046,In_0,In_122);
nand U1047 (N_1047,In_137,In_320);
xnor U1048 (N_1048,In_271,In_74);
nor U1049 (N_1049,In_465,In_347);
nor U1050 (N_1050,In_336,In_99);
nand U1051 (N_1051,In_273,In_218);
and U1052 (N_1052,In_164,In_694);
nand U1053 (N_1053,In_579,In_598);
and U1054 (N_1054,In_524,In_382);
nand U1055 (N_1055,In_678,In_683);
nand U1056 (N_1056,In_37,In_735);
nand U1057 (N_1057,In_7,In_234);
xor U1058 (N_1058,In_231,In_691);
and U1059 (N_1059,In_359,In_633);
nor U1060 (N_1060,In_315,In_259);
and U1061 (N_1061,In_602,In_353);
xor U1062 (N_1062,In_666,In_267);
and U1063 (N_1063,In_274,In_260);
nor U1064 (N_1064,In_467,In_594);
xnor U1065 (N_1065,In_639,In_424);
nor U1066 (N_1066,In_289,In_597);
and U1067 (N_1067,In_216,In_609);
xor U1068 (N_1068,In_362,In_308);
nand U1069 (N_1069,In_219,In_554);
and U1070 (N_1070,In_458,In_45);
or U1071 (N_1071,In_168,In_741);
or U1072 (N_1072,In_429,In_76);
xor U1073 (N_1073,In_704,In_480);
nand U1074 (N_1074,In_496,In_145);
or U1075 (N_1075,In_76,In_530);
nor U1076 (N_1076,In_522,In_365);
nand U1077 (N_1077,In_313,In_141);
nand U1078 (N_1078,In_612,In_102);
nand U1079 (N_1079,In_193,In_407);
or U1080 (N_1080,In_332,In_522);
nand U1081 (N_1081,In_27,In_423);
nand U1082 (N_1082,In_200,In_579);
or U1083 (N_1083,In_43,In_247);
and U1084 (N_1084,In_304,In_718);
or U1085 (N_1085,In_580,In_403);
xor U1086 (N_1086,In_622,In_258);
and U1087 (N_1087,In_1,In_547);
nor U1088 (N_1088,In_709,In_147);
and U1089 (N_1089,In_198,In_505);
nand U1090 (N_1090,In_161,In_83);
nor U1091 (N_1091,In_119,In_490);
and U1092 (N_1092,In_199,In_119);
or U1093 (N_1093,In_263,In_501);
nor U1094 (N_1094,In_454,In_631);
nand U1095 (N_1095,In_401,In_706);
or U1096 (N_1096,In_588,In_180);
nor U1097 (N_1097,In_598,In_40);
nor U1098 (N_1098,In_466,In_330);
or U1099 (N_1099,In_289,In_273);
and U1100 (N_1100,In_84,In_469);
nand U1101 (N_1101,In_30,In_228);
or U1102 (N_1102,In_24,In_408);
or U1103 (N_1103,In_547,In_70);
nor U1104 (N_1104,In_70,In_92);
nor U1105 (N_1105,In_315,In_613);
nor U1106 (N_1106,In_600,In_699);
or U1107 (N_1107,In_165,In_141);
or U1108 (N_1108,In_43,In_624);
nand U1109 (N_1109,In_174,In_550);
and U1110 (N_1110,In_701,In_17);
or U1111 (N_1111,In_344,In_251);
or U1112 (N_1112,In_231,In_325);
and U1113 (N_1113,In_180,In_655);
nand U1114 (N_1114,In_256,In_306);
and U1115 (N_1115,In_279,In_154);
or U1116 (N_1116,In_581,In_695);
nor U1117 (N_1117,In_396,In_199);
nand U1118 (N_1118,In_31,In_358);
nand U1119 (N_1119,In_321,In_573);
nand U1120 (N_1120,In_670,In_443);
or U1121 (N_1121,In_119,In_196);
and U1122 (N_1122,In_745,In_371);
and U1123 (N_1123,In_711,In_125);
nor U1124 (N_1124,In_173,In_493);
nand U1125 (N_1125,In_432,In_349);
or U1126 (N_1126,In_662,In_192);
or U1127 (N_1127,In_569,In_708);
or U1128 (N_1128,In_542,In_743);
nand U1129 (N_1129,In_450,In_325);
nor U1130 (N_1130,In_32,In_705);
or U1131 (N_1131,In_529,In_246);
xor U1132 (N_1132,In_231,In_81);
and U1133 (N_1133,In_679,In_569);
and U1134 (N_1134,In_435,In_155);
or U1135 (N_1135,In_563,In_33);
nor U1136 (N_1136,In_231,In_569);
and U1137 (N_1137,In_71,In_440);
nand U1138 (N_1138,In_206,In_630);
and U1139 (N_1139,In_625,In_39);
and U1140 (N_1140,In_335,In_378);
nand U1141 (N_1141,In_552,In_521);
nor U1142 (N_1142,In_141,In_716);
or U1143 (N_1143,In_254,In_690);
nor U1144 (N_1144,In_228,In_627);
or U1145 (N_1145,In_519,In_395);
xnor U1146 (N_1146,In_240,In_76);
nand U1147 (N_1147,In_677,In_500);
nor U1148 (N_1148,In_418,In_182);
or U1149 (N_1149,In_732,In_261);
or U1150 (N_1150,In_99,In_582);
or U1151 (N_1151,In_298,In_602);
and U1152 (N_1152,In_30,In_419);
or U1153 (N_1153,In_605,In_679);
and U1154 (N_1154,In_41,In_37);
xnor U1155 (N_1155,In_175,In_499);
nand U1156 (N_1156,In_466,In_305);
nor U1157 (N_1157,In_647,In_522);
and U1158 (N_1158,In_23,In_271);
nor U1159 (N_1159,In_328,In_88);
nand U1160 (N_1160,In_61,In_431);
xor U1161 (N_1161,In_345,In_290);
or U1162 (N_1162,In_84,In_17);
and U1163 (N_1163,In_24,In_736);
and U1164 (N_1164,In_362,In_278);
xor U1165 (N_1165,In_290,In_102);
nor U1166 (N_1166,In_237,In_721);
nor U1167 (N_1167,In_571,In_94);
or U1168 (N_1168,In_397,In_97);
nand U1169 (N_1169,In_75,In_583);
nand U1170 (N_1170,In_311,In_32);
and U1171 (N_1171,In_38,In_559);
or U1172 (N_1172,In_176,In_215);
nor U1173 (N_1173,In_421,In_350);
or U1174 (N_1174,In_256,In_312);
xor U1175 (N_1175,In_556,In_659);
and U1176 (N_1176,In_174,In_235);
xor U1177 (N_1177,In_749,In_569);
or U1178 (N_1178,In_626,In_631);
and U1179 (N_1179,In_116,In_566);
or U1180 (N_1180,In_516,In_623);
and U1181 (N_1181,In_118,In_156);
nand U1182 (N_1182,In_313,In_620);
and U1183 (N_1183,In_737,In_607);
nor U1184 (N_1184,In_549,In_724);
and U1185 (N_1185,In_453,In_148);
or U1186 (N_1186,In_69,In_194);
or U1187 (N_1187,In_50,In_363);
and U1188 (N_1188,In_708,In_472);
xor U1189 (N_1189,In_141,In_530);
nor U1190 (N_1190,In_695,In_624);
or U1191 (N_1191,In_392,In_543);
nand U1192 (N_1192,In_372,In_652);
and U1193 (N_1193,In_30,In_690);
nor U1194 (N_1194,In_27,In_348);
xor U1195 (N_1195,In_709,In_402);
nor U1196 (N_1196,In_51,In_16);
nand U1197 (N_1197,In_200,In_636);
nand U1198 (N_1198,In_511,In_692);
xnor U1199 (N_1199,In_721,In_431);
nand U1200 (N_1200,In_718,In_438);
nor U1201 (N_1201,In_230,In_409);
nor U1202 (N_1202,In_737,In_446);
nand U1203 (N_1203,In_482,In_324);
and U1204 (N_1204,In_291,In_13);
and U1205 (N_1205,In_521,In_253);
or U1206 (N_1206,In_436,In_38);
and U1207 (N_1207,In_411,In_711);
nor U1208 (N_1208,In_215,In_506);
nor U1209 (N_1209,In_310,In_701);
nor U1210 (N_1210,In_713,In_137);
or U1211 (N_1211,In_41,In_272);
or U1212 (N_1212,In_39,In_511);
nand U1213 (N_1213,In_303,In_363);
and U1214 (N_1214,In_245,In_101);
nor U1215 (N_1215,In_383,In_583);
xor U1216 (N_1216,In_678,In_629);
nor U1217 (N_1217,In_272,In_27);
or U1218 (N_1218,In_504,In_643);
nor U1219 (N_1219,In_500,In_23);
and U1220 (N_1220,In_474,In_334);
nand U1221 (N_1221,In_26,In_677);
xor U1222 (N_1222,In_747,In_449);
nand U1223 (N_1223,In_52,In_93);
or U1224 (N_1224,In_584,In_12);
nor U1225 (N_1225,In_166,In_635);
and U1226 (N_1226,In_205,In_68);
and U1227 (N_1227,In_13,In_439);
or U1228 (N_1228,In_473,In_611);
or U1229 (N_1229,In_13,In_247);
xor U1230 (N_1230,In_223,In_629);
xor U1231 (N_1231,In_602,In_158);
and U1232 (N_1232,In_369,In_242);
nand U1233 (N_1233,In_2,In_547);
nand U1234 (N_1234,In_26,In_255);
nand U1235 (N_1235,In_718,In_5);
nand U1236 (N_1236,In_711,In_208);
or U1237 (N_1237,In_709,In_639);
nor U1238 (N_1238,In_594,In_609);
or U1239 (N_1239,In_643,In_748);
nand U1240 (N_1240,In_347,In_170);
or U1241 (N_1241,In_549,In_161);
and U1242 (N_1242,In_350,In_337);
nor U1243 (N_1243,In_144,In_552);
nor U1244 (N_1244,In_493,In_154);
nand U1245 (N_1245,In_692,In_630);
xor U1246 (N_1246,In_105,In_204);
nor U1247 (N_1247,In_498,In_63);
and U1248 (N_1248,In_326,In_164);
or U1249 (N_1249,In_245,In_502);
or U1250 (N_1250,In_142,In_241);
nor U1251 (N_1251,In_705,In_110);
and U1252 (N_1252,In_463,In_58);
or U1253 (N_1253,In_564,In_531);
xnor U1254 (N_1254,In_724,In_181);
and U1255 (N_1255,In_20,In_711);
nor U1256 (N_1256,In_743,In_444);
xor U1257 (N_1257,In_520,In_744);
nor U1258 (N_1258,In_7,In_42);
and U1259 (N_1259,In_67,In_663);
and U1260 (N_1260,In_698,In_18);
and U1261 (N_1261,In_632,In_363);
or U1262 (N_1262,In_378,In_529);
nor U1263 (N_1263,In_18,In_497);
nor U1264 (N_1264,In_23,In_47);
nor U1265 (N_1265,In_147,In_92);
or U1266 (N_1266,In_427,In_376);
or U1267 (N_1267,In_623,In_157);
xnor U1268 (N_1268,In_87,In_343);
and U1269 (N_1269,In_147,In_399);
and U1270 (N_1270,In_498,In_431);
and U1271 (N_1271,In_321,In_651);
xor U1272 (N_1272,In_161,In_178);
and U1273 (N_1273,In_383,In_121);
or U1274 (N_1274,In_184,In_493);
or U1275 (N_1275,In_55,In_714);
or U1276 (N_1276,In_726,In_61);
nand U1277 (N_1277,In_730,In_320);
xnor U1278 (N_1278,In_337,In_616);
or U1279 (N_1279,In_6,In_114);
and U1280 (N_1280,In_599,In_277);
or U1281 (N_1281,In_89,In_499);
xor U1282 (N_1282,In_385,In_709);
nor U1283 (N_1283,In_749,In_424);
nand U1284 (N_1284,In_471,In_239);
or U1285 (N_1285,In_312,In_82);
and U1286 (N_1286,In_134,In_515);
nand U1287 (N_1287,In_106,In_51);
or U1288 (N_1288,In_737,In_386);
nor U1289 (N_1289,In_227,In_486);
or U1290 (N_1290,In_418,In_309);
and U1291 (N_1291,In_527,In_265);
nor U1292 (N_1292,In_68,In_188);
and U1293 (N_1293,In_532,In_104);
and U1294 (N_1294,In_136,In_708);
or U1295 (N_1295,In_311,In_133);
nor U1296 (N_1296,In_43,In_282);
nand U1297 (N_1297,In_675,In_609);
or U1298 (N_1298,In_70,In_696);
and U1299 (N_1299,In_260,In_533);
or U1300 (N_1300,In_186,In_250);
or U1301 (N_1301,In_434,In_728);
nand U1302 (N_1302,In_362,In_243);
nor U1303 (N_1303,In_376,In_259);
nor U1304 (N_1304,In_121,In_685);
xor U1305 (N_1305,In_571,In_295);
nand U1306 (N_1306,In_491,In_637);
nand U1307 (N_1307,In_261,In_214);
and U1308 (N_1308,In_292,In_28);
nand U1309 (N_1309,In_651,In_54);
nand U1310 (N_1310,In_6,In_136);
xor U1311 (N_1311,In_596,In_393);
nand U1312 (N_1312,In_98,In_158);
or U1313 (N_1313,In_259,In_137);
or U1314 (N_1314,In_225,In_391);
nand U1315 (N_1315,In_716,In_625);
nor U1316 (N_1316,In_561,In_406);
xor U1317 (N_1317,In_419,In_60);
nor U1318 (N_1318,In_110,In_385);
nor U1319 (N_1319,In_342,In_59);
or U1320 (N_1320,In_108,In_437);
nor U1321 (N_1321,In_175,In_419);
and U1322 (N_1322,In_403,In_354);
nand U1323 (N_1323,In_277,In_226);
nand U1324 (N_1324,In_145,In_253);
nor U1325 (N_1325,In_637,In_617);
xor U1326 (N_1326,In_458,In_555);
nor U1327 (N_1327,In_157,In_75);
and U1328 (N_1328,In_138,In_190);
or U1329 (N_1329,In_168,In_224);
nand U1330 (N_1330,In_414,In_16);
nor U1331 (N_1331,In_253,In_79);
and U1332 (N_1332,In_716,In_452);
nand U1333 (N_1333,In_563,In_525);
xor U1334 (N_1334,In_371,In_285);
nand U1335 (N_1335,In_517,In_232);
nand U1336 (N_1336,In_649,In_717);
and U1337 (N_1337,In_200,In_497);
nand U1338 (N_1338,In_93,In_479);
and U1339 (N_1339,In_588,In_678);
nor U1340 (N_1340,In_748,In_702);
nand U1341 (N_1341,In_408,In_549);
nand U1342 (N_1342,In_507,In_331);
xor U1343 (N_1343,In_79,In_197);
nand U1344 (N_1344,In_688,In_201);
and U1345 (N_1345,In_644,In_707);
nor U1346 (N_1346,In_613,In_273);
nor U1347 (N_1347,In_214,In_33);
nor U1348 (N_1348,In_646,In_538);
nand U1349 (N_1349,In_427,In_625);
nand U1350 (N_1350,In_91,In_268);
nand U1351 (N_1351,In_615,In_575);
nor U1352 (N_1352,In_672,In_177);
or U1353 (N_1353,In_158,In_599);
nor U1354 (N_1354,In_6,In_117);
or U1355 (N_1355,In_240,In_626);
or U1356 (N_1356,In_266,In_202);
or U1357 (N_1357,In_233,In_178);
nand U1358 (N_1358,In_416,In_600);
nand U1359 (N_1359,In_643,In_192);
nor U1360 (N_1360,In_581,In_467);
or U1361 (N_1361,In_324,In_446);
or U1362 (N_1362,In_740,In_285);
nor U1363 (N_1363,In_204,In_315);
nor U1364 (N_1364,In_200,In_540);
or U1365 (N_1365,In_70,In_199);
xor U1366 (N_1366,In_622,In_232);
and U1367 (N_1367,In_488,In_274);
or U1368 (N_1368,In_526,In_573);
nand U1369 (N_1369,In_10,In_271);
nor U1370 (N_1370,In_566,In_626);
nand U1371 (N_1371,In_676,In_293);
and U1372 (N_1372,In_630,In_127);
nand U1373 (N_1373,In_675,In_130);
nor U1374 (N_1374,In_599,In_27);
nand U1375 (N_1375,In_513,In_424);
or U1376 (N_1376,In_561,In_148);
xnor U1377 (N_1377,In_440,In_717);
nand U1378 (N_1378,In_458,In_495);
nor U1379 (N_1379,In_664,In_574);
nand U1380 (N_1380,In_534,In_151);
nor U1381 (N_1381,In_283,In_240);
or U1382 (N_1382,In_348,In_516);
nand U1383 (N_1383,In_67,In_64);
xnor U1384 (N_1384,In_643,In_237);
nand U1385 (N_1385,In_554,In_78);
xor U1386 (N_1386,In_190,In_627);
nand U1387 (N_1387,In_598,In_227);
nor U1388 (N_1388,In_365,In_658);
nand U1389 (N_1389,In_21,In_540);
or U1390 (N_1390,In_230,In_478);
and U1391 (N_1391,In_225,In_92);
nor U1392 (N_1392,In_601,In_85);
and U1393 (N_1393,In_548,In_710);
nand U1394 (N_1394,In_347,In_531);
nor U1395 (N_1395,In_537,In_354);
or U1396 (N_1396,In_534,In_295);
xor U1397 (N_1397,In_327,In_533);
nor U1398 (N_1398,In_591,In_449);
and U1399 (N_1399,In_575,In_608);
and U1400 (N_1400,In_201,In_641);
or U1401 (N_1401,In_315,In_612);
and U1402 (N_1402,In_25,In_459);
or U1403 (N_1403,In_220,In_401);
nand U1404 (N_1404,In_125,In_266);
xor U1405 (N_1405,In_575,In_408);
nand U1406 (N_1406,In_469,In_413);
and U1407 (N_1407,In_101,In_532);
nor U1408 (N_1408,In_29,In_570);
xnor U1409 (N_1409,In_516,In_665);
nor U1410 (N_1410,In_119,In_66);
nor U1411 (N_1411,In_289,In_178);
nand U1412 (N_1412,In_154,In_42);
or U1413 (N_1413,In_644,In_678);
and U1414 (N_1414,In_611,In_51);
xor U1415 (N_1415,In_54,In_430);
or U1416 (N_1416,In_720,In_550);
nor U1417 (N_1417,In_401,In_28);
nor U1418 (N_1418,In_535,In_472);
nor U1419 (N_1419,In_433,In_187);
and U1420 (N_1420,In_295,In_266);
xnor U1421 (N_1421,In_639,In_433);
and U1422 (N_1422,In_91,In_525);
nor U1423 (N_1423,In_517,In_324);
xnor U1424 (N_1424,In_616,In_373);
nor U1425 (N_1425,In_612,In_657);
or U1426 (N_1426,In_141,In_292);
or U1427 (N_1427,In_154,In_629);
or U1428 (N_1428,In_121,In_79);
and U1429 (N_1429,In_564,In_164);
xnor U1430 (N_1430,In_435,In_468);
and U1431 (N_1431,In_634,In_213);
or U1432 (N_1432,In_198,In_418);
nor U1433 (N_1433,In_662,In_183);
nand U1434 (N_1434,In_553,In_401);
and U1435 (N_1435,In_487,In_46);
nand U1436 (N_1436,In_62,In_501);
and U1437 (N_1437,In_735,In_357);
or U1438 (N_1438,In_95,In_226);
xnor U1439 (N_1439,In_736,In_399);
nand U1440 (N_1440,In_570,In_534);
and U1441 (N_1441,In_137,In_343);
and U1442 (N_1442,In_488,In_685);
or U1443 (N_1443,In_339,In_398);
or U1444 (N_1444,In_123,In_168);
nor U1445 (N_1445,In_84,In_465);
and U1446 (N_1446,In_144,In_317);
nand U1447 (N_1447,In_743,In_3);
nand U1448 (N_1448,In_146,In_687);
and U1449 (N_1449,In_354,In_153);
or U1450 (N_1450,In_400,In_258);
nor U1451 (N_1451,In_315,In_699);
and U1452 (N_1452,In_417,In_525);
and U1453 (N_1453,In_291,In_353);
and U1454 (N_1454,In_487,In_625);
and U1455 (N_1455,In_2,In_644);
or U1456 (N_1456,In_113,In_654);
xor U1457 (N_1457,In_662,In_720);
nor U1458 (N_1458,In_24,In_203);
and U1459 (N_1459,In_615,In_365);
or U1460 (N_1460,In_53,In_133);
xnor U1461 (N_1461,In_404,In_16);
nor U1462 (N_1462,In_247,In_592);
nand U1463 (N_1463,In_585,In_285);
and U1464 (N_1464,In_115,In_638);
nand U1465 (N_1465,In_165,In_183);
or U1466 (N_1466,In_401,In_385);
nand U1467 (N_1467,In_349,In_561);
nand U1468 (N_1468,In_160,In_401);
nor U1469 (N_1469,In_521,In_386);
and U1470 (N_1470,In_17,In_393);
xnor U1471 (N_1471,In_443,In_344);
nand U1472 (N_1472,In_422,In_314);
and U1473 (N_1473,In_98,In_635);
nand U1474 (N_1474,In_2,In_325);
or U1475 (N_1475,In_167,In_357);
nor U1476 (N_1476,In_618,In_48);
nand U1477 (N_1477,In_645,In_75);
nand U1478 (N_1478,In_281,In_42);
nand U1479 (N_1479,In_51,In_438);
xnor U1480 (N_1480,In_527,In_456);
or U1481 (N_1481,In_336,In_676);
nand U1482 (N_1482,In_497,In_190);
and U1483 (N_1483,In_435,In_9);
and U1484 (N_1484,In_68,In_531);
xor U1485 (N_1485,In_374,In_574);
and U1486 (N_1486,In_13,In_444);
or U1487 (N_1487,In_342,In_328);
xnor U1488 (N_1488,In_681,In_745);
and U1489 (N_1489,In_187,In_223);
or U1490 (N_1490,In_201,In_406);
nor U1491 (N_1491,In_676,In_346);
nor U1492 (N_1492,In_550,In_164);
xor U1493 (N_1493,In_602,In_223);
nand U1494 (N_1494,In_190,In_304);
or U1495 (N_1495,In_425,In_517);
nor U1496 (N_1496,In_716,In_50);
nand U1497 (N_1497,In_550,In_395);
nor U1498 (N_1498,In_602,In_236);
nor U1499 (N_1499,In_187,In_263);
and U1500 (N_1500,In_29,In_644);
nor U1501 (N_1501,In_649,In_6);
and U1502 (N_1502,In_298,In_406);
xnor U1503 (N_1503,In_320,In_80);
xor U1504 (N_1504,In_551,In_368);
nand U1505 (N_1505,In_316,In_423);
nor U1506 (N_1506,In_449,In_63);
and U1507 (N_1507,In_220,In_272);
or U1508 (N_1508,In_536,In_132);
xor U1509 (N_1509,In_181,In_407);
nand U1510 (N_1510,In_518,In_20);
or U1511 (N_1511,In_210,In_114);
and U1512 (N_1512,In_160,In_100);
nand U1513 (N_1513,In_231,In_433);
nor U1514 (N_1514,In_657,In_9);
and U1515 (N_1515,In_730,In_473);
and U1516 (N_1516,In_272,In_723);
nand U1517 (N_1517,In_629,In_742);
xnor U1518 (N_1518,In_11,In_684);
nand U1519 (N_1519,In_560,In_550);
nand U1520 (N_1520,In_652,In_49);
nand U1521 (N_1521,In_727,In_251);
xnor U1522 (N_1522,In_486,In_92);
and U1523 (N_1523,In_352,In_205);
nor U1524 (N_1524,In_83,In_657);
or U1525 (N_1525,In_670,In_123);
or U1526 (N_1526,In_642,In_444);
or U1527 (N_1527,In_197,In_140);
nand U1528 (N_1528,In_608,In_68);
xnor U1529 (N_1529,In_376,In_485);
or U1530 (N_1530,In_98,In_294);
and U1531 (N_1531,In_418,In_616);
nand U1532 (N_1532,In_741,In_608);
nand U1533 (N_1533,In_173,In_146);
nor U1534 (N_1534,In_443,In_550);
and U1535 (N_1535,In_156,In_228);
or U1536 (N_1536,In_598,In_459);
nand U1537 (N_1537,In_169,In_201);
or U1538 (N_1538,In_356,In_234);
and U1539 (N_1539,In_403,In_532);
xnor U1540 (N_1540,In_35,In_446);
and U1541 (N_1541,In_633,In_420);
nand U1542 (N_1542,In_46,In_349);
and U1543 (N_1543,In_628,In_149);
xnor U1544 (N_1544,In_153,In_367);
or U1545 (N_1545,In_586,In_434);
or U1546 (N_1546,In_739,In_236);
nand U1547 (N_1547,In_203,In_615);
nor U1548 (N_1548,In_232,In_606);
or U1549 (N_1549,In_46,In_382);
xnor U1550 (N_1550,In_555,In_548);
or U1551 (N_1551,In_433,In_656);
nand U1552 (N_1552,In_459,In_566);
and U1553 (N_1553,In_149,In_547);
nand U1554 (N_1554,In_451,In_597);
xor U1555 (N_1555,In_711,In_563);
xor U1556 (N_1556,In_124,In_676);
xnor U1557 (N_1557,In_639,In_559);
or U1558 (N_1558,In_274,In_215);
nand U1559 (N_1559,In_480,In_577);
nor U1560 (N_1560,In_266,In_385);
nor U1561 (N_1561,In_219,In_437);
or U1562 (N_1562,In_547,In_119);
nor U1563 (N_1563,In_200,In_682);
nand U1564 (N_1564,In_549,In_354);
or U1565 (N_1565,In_266,In_26);
nand U1566 (N_1566,In_450,In_467);
nand U1567 (N_1567,In_238,In_245);
and U1568 (N_1568,In_199,In_331);
or U1569 (N_1569,In_245,In_556);
nand U1570 (N_1570,In_305,In_404);
and U1571 (N_1571,In_426,In_723);
nand U1572 (N_1572,In_29,In_282);
nor U1573 (N_1573,In_471,In_450);
nand U1574 (N_1574,In_300,In_340);
and U1575 (N_1575,In_99,In_696);
or U1576 (N_1576,In_58,In_337);
and U1577 (N_1577,In_598,In_345);
and U1578 (N_1578,In_163,In_619);
xnor U1579 (N_1579,In_696,In_675);
nor U1580 (N_1580,In_625,In_316);
and U1581 (N_1581,In_36,In_2);
nor U1582 (N_1582,In_99,In_145);
or U1583 (N_1583,In_51,In_78);
or U1584 (N_1584,In_386,In_394);
nand U1585 (N_1585,In_19,In_571);
or U1586 (N_1586,In_708,In_126);
and U1587 (N_1587,In_681,In_298);
nor U1588 (N_1588,In_103,In_335);
nor U1589 (N_1589,In_473,In_640);
and U1590 (N_1590,In_598,In_667);
nor U1591 (N_1591,In_568,In_338);
and U1592 (N_1592,In_189,In_362);
nand U1593 (N_1593,In_539,In_545);
nand U1594 (N_1594,In_522,In_19);
and U1595 (N_1595,In_665,In_4);
and U1596 (N_1596,In_685,In_745);
nor U1597 (N_1597,In_517,In_471);
and U1598 (N_1598,In_478,In_301);
nor U1599 (N_1599,In_98,In_84);
or U1600 (N_1600,In_390,In_669);
nor U1601 (N_1601,In_376,In_608);
nand U1602 (N_1602,In_628,In_100);
or U1603 (N_1603,In_135,In_681);
nand U1604 (N_1604,In_21,In_238);
or U1605 (N_1605,In_541,In_742);
nor U1606 (N_1606,In_452,In_696);
and U1607 (N_1607,In_25,In_397);
nor U1608 (N_1608,In_455,In_50);
and U1609 (N_1609,In_279,In_634);
nand U1610 (N_1610,In_105,In_304);
nand U1611 (N_1611,In_364,In_675);
nand U1612 (N_1612,In_655,In_463);
or U1613 (N_1613,In_73,In_103);
and U1614 (N_1614,In_394,In_280);
xnor U1615 (N_1615,In_485,In_504);
nor U1616 (N_1616,In_235,In_463);
nand U1617 (N_1617,In_308,In_23);
nor U1618 (N_1618,In_647,In_90);
nor U1619 (N_1619,In_194,In_90);
nor U1620 (N_1620,In_722,In_13);
nor U1621 (N_1621,In_160,In_553);
nand U1622 (N_1622,In_452,In_470);
xor U1623 (N_1623,In_673,In_178);
or U1624 (N_1624,In_417,In_634);
nor U1625 (N_1625,In_89,In_205);
nor U1626 (N_1626,In_466,In_449);
nand U1627 (N_1627,In_638,In_8);
nand U1628 (N_1628,In_179,In_591);
or U1629 (N_1629,In_172,In_399);
and U1630 (N_1630,In_728,In_621);
nand U1631 (N_1631,In_604,In_320);
or U1632 (N_1632,In_234,In_300);
nor U1633 (N_1633,In_214,In_123);
nand U1634 (N_1634,In_201,In_392);
nor U1635 (N_1635,In_694,In_17);
nand U1636 (N_1636,In_156,In_329);
and U1637 (N_1637,In_543,In_290);
and U1638 (N_1638,In_667,In_542);
xor U1639 (N_1639,In_240,In_47);
xnor U1640 (N_1640,In_230,In_669);
nor U1641 (N_1641,In_260,In_68);
nand U1642 (N_1642,In_277,In_194);
and U1643 (N_1643,In_620,In_219);
nor U1644 (N_1644,In_103,In_170);
and U1645 (N_1645,In_443,In_609);
xor U1646 (N_1646,In_258,In_189);
nand U1647 (N_1647,In_427,In_458);
xor U1648 (N_1648,In_738,In_196);
nand U1649 (N_1649,In_373,In_80);
nor U1650 (N_1650,In_56,In_749);
nor U1651 (N_1651,In_376,In_0);
or U1652 (N_1652,In_168,In_349);
or U1653 (N_1653,In_722,In_742);
or U1654 (N_1654,In_90,In_743);
xor U1655 (N_1655,In_385,In_475);
xor U1656 (N_1656,In_744,In_587);
or U1657 (N_1657,In_521,In_430);
nand U1658 (N_1658,In_443,In_347);
nor U1659 (N_1659,In_317,In_12);
or U1660 (N_1660,In_683,In_211);
and U1661 (N_1661,In_741,In_604);
and U1662 (N_1662,In_723,In_209);
nor U1663 (N_1663,In_298,In_726);
or U1664 (N_1664,In_679,In_24);
or U1665 (N_1665,In_87,In_575);
or U1666 (N_1666,In_557,In_715);
nor U1667 (N_1667,In_226,In_114);
xor U1668 (N_1668,In_698,In_15);
xor U1669 (N_1669,In_707,In_241);
or U1670 (N_1670,In_194,In_286);
or U1671 (N_1671,In_544,In_542);
or U1672 (N_1672,In_306,In_546);
nor U1673 (N_1673,In_345,In_104);
or U1674 (N_1674,In_549,In_426);
and U1675 (N_1675,In_526,In_404);
xor U1676 (N_1676,In_301,In_225);
or U1677 (N_1677,In_722,In_71);
and U1678 (N_1678,In_195,In_589);
and U1679 (N_1679,In_509,In_101);
or U1680 (N_1680,In_615,In_595);
nor U1681 (N_1681,In_136,In_180);
or U1682 (N_1682,In_522,In_687);
or U1683 (N_1683,In_352,In_241);
nor U1684 (N_1684,In_84,In_23);
xor U1685 (N_1685,In_225,In_532);
nor U1686 (N_1686,In_390,In_385);
nand U1687 (N_1687,In_594,In_253);
or U1688 (N_1688,In_717,In_225);
nor U1689 (N_1689,In_671,In_560);
and U1690 (N_1690,In_624,In_175);
nand U1691 (N_1691,In_336,In_532);
and U1692 (N_1692,In_354,In_650);
nand U1693 (N_1693,In_310,In_537);
nand U1694 (N_1694,In_370,In_628);
nand U1695 (N_1695,In_341,In_346);
and U1696 (N_1696,In_309,In_312);
xnor U1697 (N_1697,In_702,In_707);
nand U1698 (N_1698,In_569,In_281);
or U1699 (N_1699,In_42,In_11);
and U1700 (N_1700,In_393,In_6);
or U1701 (N_1701,In_381,In_303);
nor U1702 (N_1702,In_593,In_126);
and U1703 (N_1703,In_401,In_659);
nor U1704 (N_1704,In_175,In_9);
xor U1705 (N_1705,In_496,In_57);
or U1706 (N_1706,In_447,In_322);
nand U1707 (N_1707,In_61,In_220);
nand U1708 (N_1708,In_521,In_179);
xor U1709 (N_1709,In_505,In_654);
xnor U1710 (N_1710,In_407,In_161);
and U1711 (N_1711,In_545,In_578);
and U1712 (N_1712,In_293,In_320);
and U1713 (N_1713,In_316,In_587);
nor U1714 (N_1714,In_644,In_479);
or U1715 (N_1715,In_214,In_487);
nand U1716 (N_1716,In_576,In_619);
nor U1717 (N_1717,In_411,In_244);
and U1718 (N_1718,In_357,In_26);
nor U1719 (N_1719,In_492,In_489);
xor U1720 (N_1720,In_503,In_343);
nand U1721 (N_1721,In_548,In_623);
and U1722 (N_1722,In_307,In_559);
nor U1723 (N_1723,In_234,In_495);
or U1724 (N_1724,In_727,In_55);
and U1725 (N_1725,In_215,In_748);
and U1726 (N_1726,In_125,In_738);
nor U1727 (N_1727,In_370,In_427);
xnor U1728 (N_1728,In_499,In_396);
xnor U1729 (N_1729,In_385,In_693);
nor U1730 (N_1730,In_730,In_526);
and U1731 (N_1731,In_732,In_64);
xnor U1732 (N_1732,In_376,In_670);
and U1733 (N_1733,In_450,In_257);
nor U1734 (N_1734,In_444,In_209);
or U1735 (N_1735,In_733,In_43);
nand U1736 (N_1736,In_455,In_134);
and U1737 (N_1737,In_271,In_716);
nand U1738 (N_1738,In_702,In_521);
and U1739 (N_1739,In_16,In_680);
and U1740 (N_1740,In_186,In_21);
xor U1741 (N_1741,In_207,In_406);
or U1742 (N_1742,In_493,In_207);
or U1743 (N_1743,In_183,In_67);
or U1744 (N_1744,In_136,In_84);
xnor U1745 (N_1745,In_701,In_351);
xor U1746 (N_1746,In_542,In_728);
and U1747 (N_1747,In_618,In_244);
or U1748 (N_1748,In_453,In_377);
nor U1749 (N_1749,In_600,In_425);
nor U1750 (N_1750,In_122,In_271);
or U1751 (N_1751,In_162,In_106);
xor U1752 (N_1752,In_374,In_720);
or U1753 (N_1753,In_523,In_705);
xnor U1754 (N_1754,In_29,In_99);
nor U1755 (N_1755,In_584,In_131);
or U1756 (N_1756,In_97,In_746);
or U1757 (N_1757,In_513,In_673);
xor U1758 (N_1758,In_60,In_330);
nand U1759 (N_1759,In_179,In_216);
and U1760 (N_1760,In_537,In_665);
nand U1761 (N_1761,In_362,In_406);
or U1762 (N_1762,In_333,In_666);
nand U1763 (N_1763,In_740,In_733);
or U1764 (N_1764,In_264,In_643);
and U1765 (N_1765,In_568,In_494);
and U1766 (N_1766,In_95,In_212);
and U1767 (N_1767,In_632,In_330);
nor U1768 (N_1768,In_172,In_359);
xor U1769 (N_1769,In_448,In_220);
nor U1770 (N_1770,In_622,In_42);
or U1771 (N_1771,In_186,In_412);
nor U1772 (N_1772,In_4,In_612);
nand U1773 (N_1773,In_677,In_582);
nor U1774 (N_1774,In_336,In_677);
or U1775 (N_1775,In_41,In_48);
xor U1776 (N_1776,In_190,In_533);
nor U1777 (N_1777,In_404,In_531);
and U1778 (N_1778,In_705,In_508);
nor U1779 (N_1779,In_647,In_575);
nand U1780 (N_1780,In_151,In_257);
nand U1781 (N_1781,In_48,In_349);
and U1782 (N_1782,In_201,In_415);
xor U1783 (N_1783,In_710,In_290);
and U1784 (N_1784,In_29,In_546);
nor U1785 (N_1785,In_238,In_525);
nand U1786 (N_1786,In_75,In_23);
or U1787 (N_1787,In_254,In_308);
nand U1788 (N_1788,In_187,In_106);
nor U1789 (N_1789,In_148,In_108);
xor U1790 (N_1790,In_92,In_678);
and U1791 (N_1791,In_280,In_108);
nor U1792 (N_1792,In_613,In_333);
nor U1793 (N_1793,In_277,In_19);
nand U1794 (N_1794,In_550,In_581);
nor U1795 (N_1795,In_64,In_477);
nor U1796 (N_1796,In_512,In_420);
and U1797 (N_1797,In_537,In_292);
nand U1798 (N_1798,In_247,In_1);
or U1799 (N_1799,In_11,In_49);
and U1800 (N_1800,In_614,In_198);
or U1801 (N_1801,In_695,In_63);
nand U1802 (N_1802,In_170,In_91);
or U1803 (N_1803,In_247,In_706);
nor U1804 (N_1804,In_509,In_683);
nor U1805 (N_1805,In_51,In_693);
nor U1806 (N_1806,In_328,In_442);
or U1807 (N_1807,In_258,In_427);
nor U1808 (N_1808,In_113,In_112);
or U1809 (N_1809,In_397,In_129);
or U1810 (N_1810,In_96,In_102);
nor U1811 (N_1811,In_562,In_726);
nor U1812 (N_1812,In_589,In_212);
nand U1813 (N_1813,In_524,In_63);
or U1814 (N_1814,In_498,In_743);
or U1815 (N_1815,In_213,In_484);
xor U1816 (N_1816,In_306,In_495);
nor U1817 (N_1817,In_347,In_714);
or U1818 (N_1818,In_86,In_729);
nor U1819 (N_1819,In_509,In_578);
nand U1820 (N_1820,In_129,In_655);
or U1821 (N_1821,In_519,In_88);
and U1822 (N_1822,In_74,In_445);
or U1823 (N_1823,In_60,In_72);
nand U1824 (N_1824,In_544,In_330);
nand U1825 (N_1825,In_355,In_499);
xnor U1826 (N_1826,In_149,In_81);
and U1827 (N_1827,In_576,In_117);
nand U1828 (N_1828,In_311,In_298);
or U1829 (N_1829,In_512,In_539);
nor U1830 (N_1830,In_70,In_463);
or U1831 (N_1831,In_176,In_533);
nand U1832 (N_1832,In_380,In_225);
nand U1833 (N_1833,In_660,In_437);
nor U1834 (N_1834,In_473,In_487);
nor U1835 (N_1835,In_492,In_695);
or U1836 (N_1836,In_582,In_199);
or U1837 (N_1837,In_726,In_700);
and U1838 (N_1838,In_81,In_264);
and U1839 (N_1839,In_625,In_42);
and U1840 (N_1840,In_321,In_660);
nand U1841 (N_1841,In_159,In_13);
or U1842 (N_1842,In_4,In_40);
or U1843 (N_1843,In_363,In_631);
nand U1844 (N_1844,In_678,In_54);
nor U1845 (N_1845,In_723,In_555);
and U1846 (N_1846,In_407,In_134);
and U1847 (N_1847,In_265,In_413);
nor U1848 (N_1848,In_31,In_226);
nand U1849 (N_1849,In_331,In_463);
nand U1850 (N_1850,In_90,In_114);
or U1851 (N_1851,In_460,In_445);
nor U1852 (N_1852,In_475,In_312);
or U1853 (N_1853,In_116,In_562);
or U1854 (N_1854,In_570,In_553);
or U1855 (N_1855,In_646,In_667);
or U1856 (N_1856,In_710,In_520);
xnor U1857 (N_1857,In_426,In_524);
or U1858 (N_1858,In_712,In_719);
and U1859 (N_1859,In_368,In_240);
nor U1860 (N_1860,In_54,In_566);
nor U1861 (N_1861,In_603,In_605);
and U1862 (N_1862,In_557,In_423);
nor U1863 (N_1863,In_506,In_44);
xnor U1864 (N_1864,In_26,In_572);
nand U1865 (N_1865,In_72,In_278);
xor U1866 (N_1866,In_333,In_224);
or U1867 (N_1867,In_615,In_280);
nor U1868 (N_1868,In_681,In_59);
nor U1869 (N_1869,In_219,In_673);
or U1870 (N_1870,In_548,In_178);
and U1871 (N_1871,In_567,In_26);
and U1872 (N_1872,In_442,In_436);
xnor U1873 (N_1873,In_326,In_337);
and U1874 (N_1874,In_214,In_740);
or U1875 (N_1875,In_518,In_430);
or U1876 (N_1876,In_178,In_112);
and U1877 (N_1877,In_707,In_289);
nor U1878 (N_1878,In_618,In_516);
xnor U1879 (N_1879,In_379,In_16);
and U1880 (N_1880,In_14,In_162);
or U1881 (N_1881,In_667,In_402);
xor U1882 (N_1882,In_128,In_439);
xnor U1883 (N_1883,In_116,In_715);
nor U1884 (N_1884,In_156,In_312);
and U1885 (N_1885,In_515,In_196);
and U1886 (N_1886,In_680,In_519);
nor U1887 (N_1887,In_499,In_746);
or U1888 (N_1888,In_620,In_731);
and U1889 (N_1889,In_81,In_711);
or U1890 (N_1890,In_59,In_172);
nand U1891 (N_1891,In_297,In_448);
and U1892 (N_1892,In_572,In_595);
nand U1893 (N_1893,In_161,In_456);
nor U1894 (N_1894,In_640,In_534);
nand U1895 (N_1895,In_267,In_93);
xnor U1896 (N_1896,In_49,In_0);
nor U1897 (N_1897,In_86,In_333);
or U1898 (N_1898,In_692,In_647);
and U1899 (N_1899,In_657,In_70);
nor U1900 (N_1900,In_93,In_688);
and U1901 (N_1901,In_497,In_377);
xnor U1902 (N_1902,In_571,In_543);
and U1903 (N_1903,In_15,In_377);
or U1904 (N_1904,In_603,In_152);
or U1905 (N_1905,In_379,In_13);
or U1906 (N_1906,In_681,In_115);
or U1907 (N_1907,In_635,In_568);
and U1908 (N_1908,In_742,In_2);
or U1909 (N_1909,In_189,In_435);
nor U1910 (N_1910,In_649,In_325);
nand U1911 (N_1911,In_375,In_208);
and U1912 (N_1912,In_486,In_695);
or U1913 (N_1913,In_728,In_517);
and U1914 (N_1914,In_63,In_470);
or U1915 (N_1915,In_196,In_483);
xnor U1916 (N_1916,In_8,In_81);
or U1917 (N_1917,In_159,In_429);
nor U1918 (N_1918,In_253,In_739);
nand U1919 (N_1919,In_690,In_27);
nor U1920 (N_1920,In_578,In_490);
nand U1921 (N_1921,In_44,In_502);
nand U1922 (N_1922,In_559,In_365);
nand U1923 (N_1923,In_250,In_238);
and U1924 (N_1924,In_405,In_651);
or U1925 (N_1925,In_395,In_313);
nand U1926 (N_1926,In_660,In_435);
or U1927 (N_1927,In_402,In_92);
and U1928 (N_1928,In_464,In_592);
xor U1929 (N_1929,In_446,In_610);
nor U1930 (N_1930,In_35,In_648);
nand U1931 (N_1931,In_725,In_157);
nor U1932 (N_1932,In_732,In_38);
nor U1933 (N_1933,In_389,In_662);
and U1934 (N_1934,In_61,In_286);
and U1935 (N_1935,In_122,In_375);
nor U1936 (N_1936,In_430,In_174);
or U1937 (N_1937,In_535,In_199);
nor U1938 (N_1938,In_595,In_473);
and U1939 (N_1939,In_24,In_535);
nand U1940 (N_1940,In_438,In_332);
nor U1941 (N_1941,In_17,In_474);
nand U1942 (N_1942,In_695,In_168);
nor U1943 (N_1943,In_732,In_395);
nor U1944 (N_1944,In_496,In_651);
and U1945 (N_1945,In_231,In_625);
nand U1946 (N_1946,In_347,In_529);
nand U1947 (N_1947,In_497,In_428);
xnor U1948 (N_1948,In_181,In_706);
or U1949 (N_1949,In_266,In_639);
nor U1950 (N_1950,In_154,In_369);
and U1951 (N_1951,In_16,In_407);
and U1952 (N_1952,In_61,In_69);
and U1953 (N_1953,In_665,In_673);
nand U1954 (N_1954,In_298,In_107);
or U1955 (N_1955,In_682,In_71);
nand U1956 (N_1956,In_51,In_656);
nor U1957 (N_1957,In_589,In_560);
and U1958 (N_1958,In_721,In_69);
or U1959 (N_1959,In_225,In_620);
and U1960 (N_1960,In_654,In_328);
and U1961 (N_1961,In_459,In_35);
nand U1962 (N_1962,In_408,In_613);
and U1963 (N_1963,In_342,In_715);
and U1964 (N_1964,In_233,In_271);
nand U1965 (N_1965,In_97,In_66);
xor U1966 (N_1966,In_62,In_132);
or U1967 (N_1967,In_142,In_655);
nand U1968 (N_1968,In_722,In_427);
or U1969 (N_1969,In_676,In_644);
nor U1970 (N_1970,In_730,In_208);
and U1971 (N_1971,In_437,In_275);
nand U1972 (N_1972,In_104,In_39);
nand U1973 (N_1973,In_582,In_83);
and U1974 (N_1974,In_274,In_466);
or U1975 (N_1975,In_135,In_309);
or U1976 (N_1976,In_697,In_285);
and U1977 (N_1977,In_297,In_385);
and U1978 (N_1978,In_209,In_689);
or U1979 (N_1979,In_171,In_542);
and U1980 (N_1980,In_341,In_3);
and U1981 (N_1981,In_689,In_151);
and U1982 (N_1982,In_317,In_305);
nand U1983 (N_1983,In_625,In_229);
and U1984 (N_1984,In_300,In_410);
or U1985 (N_1985,In_340,In_418);
nand U1986 (N_1986,In_683,In_742);
and U1987 (N_1987,In_70,In_699);
xnor U1988 (N_1988,In_442,In_668);
nand U1989 (N_1989,In_538,In_339);
nor U1990 (N_1990,In_255,In_29);
nor U1991 (N_1991,In_732,In_246);
or U1992 (N_1992,In_226,In_123);
nand U1993 (N_1993,In_538,In_642);
nand U1994 (N_1994,In_157,In_695);
and U1995 (N_1995,In_643,In_370);
nand U1996 (N_1996,In_232,In_324);
or U1997 (N_1997,In_491,In_479);
nor U1998 (N_1998,In_417,In_269);
or U1999 (N_1999,In_504,In_283);
and U2000 (N_2000,In_496,In_650);
and U2001 (N_2001,In_544,In_487);
nor U2002 (N_2002,In_653,In_228);
nor U2003 (N_2003,In_300,In_614);
or U2004 (N_2004,In_674,In_715);
and U2005 (N_2005,In_428,In_430);
and U2006 (N_2006,In_612,In_461);
and U2007 (N_2007,In_719,In_380);
and U2008 (N_2008,In_34,In_89);
nor U2009 (N_2009,In_307,In_416);
xnor U2010 (N_2010,In_558,In_522);
or U2011 (N_2011,In_580,In_350);
and U2012 (N_2012,In_725,In_315);
nor U2013 (N_2013,In_367,In_155);
and U2014 (N_2014,In_480,In_72);
and U2015 (N_2015,In_51,In_226);
and U2016 (N_2016,In_296,In_326);
nand U2017 (N_2017,In_58,In_308);
and U2018 (N_2018,In_257,In_636);
nor U2019 (N_2019,In_318,In_706);
and U2020 (N_2020,In_603,In_94);
nand U2021 (N_2021,In_17,In_657);
xnor U2022 (N_2022,In_113,In_263);
or U2023 (N_2023,In_653,In_64);
nor U2024 (N_2024,In_15,In_603);
nor U2025 (N_2025,In_310,In_55);
and U2026 (N_2026,In_58,In_249);
nor U2027 (N_2027,In_570,In_671);
nor U2028 (N_2028,In_414,In_210);
and U2029 (N_2029,In_570,In_363);
nand U2030 (N_2030,In_39,In_194);
nor U2031 (N_2031,In_578,In_199);
nor U2032 (N_2032,In_508,In_746);
nand U2033 (N_2033,In_544,In_207);
or U2034 (N_2034,In_580,In_48);
and U2035 (N_2035,In_279,In_354);
nor U2036 (N_2036,In_345,In_314);
nor U2037 (N_2037,In_350,In_480);
xnor U2038 (N_2038,In_480,In_373);
nor U2039 (N_2039,In_272,In_72);
nand U2040 (N_2040,In_584,In_214);
and U2041 (N_2041,In_382,In_668);
nor U2042 (N_2042,In_724,In_386);
nor U2043 (N_2043,In_521,In_559);
and U2044 (N_2044,In_327,In_539);
or U2045 (N_2045,In_716,In_534);
xor U2046 (N_2046,In_375,In_243);
or U2047 (N_2047,In_636,In_84);
nor U2048 (N_2048,In_655,In_591);
nand U2049 (N_2049,In_612,In_205);
and U2050 (N_2050,In_351,In_347);
xor U2051 (N_2051,In_333,In_185);
nand U2052 (N_2052,In_412,In_742);
or U2053 (N_2053,In_625,In_700);
or U2054 (N_2054,In_239,In_39);
nand U2055 (N_2055,In_333,In_568);
nand U2056 (N_2056,In_228,In_529);
nand U2057 (N_2057,In_330,In_588);
or U2058 (N_2058,In_600,In_418);
or U2059 (N_2059,In_390,In_488);
and U2060 (N_2060,In_144,In_401);
or U2061 (N_2061,In_675,In_476);
nand U2062 (N_2062,In_688,In_374);
or U2063 (N_2063,In_46,In_372);
or U2064 (N_2064,In_690,In_21);
xor U2065 (N_2065,In_154,In_335);
or U2066 (N_2066,In_709,In_187);
nor U2067 (N_2067,In_168,In_330);
or U2068 (N_2068,In_50,In_183);
xnor U2069 (N_2069,In_183,In_714);
xor U2070 (N_2070,In_546,In_383);
nor U2071 (N_2071,In_402,In_571);
nand U2072 (N_2072,In_698,In_215);
or U2073 (N_2073,In_702,In_625);
nand U2074 (N_2074,In_425,In_61);
and U2075 (N_2075,In_538,In_45);
or U2076 (N_2076,In_287,In_540);
or U2077 (N_2077,In_367,In_253);
nor U2078 (N_2078,In_655,In_194);
nand U2079 (N_2079,In_222,In_154);
or U2080 (N_2080,In_386,In_626);
nand U2081 (N_2081,In_53,In_219);
nand U2082 (N_2082,In_748,In_398);
and U2083 (N_2083,In_164,In_373);
nor U2084 (N_2084,In_420,In_396);
nor U2085 (N_2085,In_36,In_287);
nor U2086 (N_2086,In_562,In_382);
nor U2087 (N_2087,In_703,In_320);
and U2088 (N_2088,In_141,In_635);
or U2089 (N_2089,In_475,In_433);
and U2090 (N_2090,In_265,In_219);
nand U2091 (N_2091,In_299,In_118);
nor U2092 (N_2092,In_335,In_723);
xnor U2093 (N_2093,In_279,In_221);
nand U2094 (N_2094,In_53,In_723);
nand U2095 (N_2095,In_485,In_428);
nand U2096 (N_2096,In_48,In_204);
and U2097 (N_2097,In_103,In_531);
xor U2098 (N_2098,In_388,In_225);
and U2099 (N_2099,In_321,In_36);
or U2100 (N_2100,In_484,In_718);
nor U2101 (N_2101,In_210,In_365);
or U2102 (N_2102,In_292,In_458);
and U2103 (N_2103,In_425,In_242);
nor U2104 (N_2104,In_155,In_673);
or U2105 (N_2105,In_100,In_582);
or U2106 (N_2106,In_29,In_727);
or U2107 (N_2107,In_720,In_200);
or U2108 (N_2108,In_408,In_522);
or U2109 (N_2109,In_269,In_56);
and U2110 (N_2110,In_539,In_358);
nand U2111 (N_2111,In_362,In_345);
or U2112 (N_2112,In_504,In_423);
nand U2113 (N_2113,In_480,In_421);
nand U2114 (N_2114,In_714,In_117);
nor U2115 (N_2115,In_40,In_228);
nand U2116 (N_2116,In_156,In_661);
or U2117 (N_2117,In_243,In_456);
nor U2118 (N_2118,In_593,In_548);
nor U2119 (N_2119,In_571,In_301);
xor U2120 (N_2120,In_491,In_327);
nand U2121 (N_2121,In_318,In_156);
nor U2122 (N_2122,In_120,In_240);
and U2123 (N_2123,In_315,In_232);
and U2124 (N_2124,In_564,In_78);
nand U2125 (N_2125,In_526,In_348);
xnor U2126 (N_2126,In_679,In_15);
nor U2127 (N_2127,In_191,In_690);
and U2128 (N_2128,In_55,In_340);
or U2129 (N_2129,In_266,In_664);
nand U2130 (N_2130,In_401,In_520);
or U2131 (N_2131,In_172,In_132);
nand U2132 (N_2132,In_340,In_284);
and U2133 (N_2133,In_206,In_586);
and U2134 (N_2134,In_394,In_620);
nor U2135 (N_2135,In_42,In_129);
nor U2136 (N_2136,In_456,In_625);
and U2137 (N_2137,In_732,In_592);
nor U2138 (N_2138,In_547,In_571);
or U2139 (N_2139,In_78,In_615);
xnor U2140 (N_2140,In_611,In_528);
xor U2141 (N_2141,In_695,In_471);
nand U2142 (N_2142,In_690,In_587);
and U2143 (N_2143,In_662,In_169);
nor U2144 (N_2144,In_49,In_484);
and U2145 (N_2145,In_162,In_698);
and U2146 (N_2146,In_563,In_315);
nor U2147 (N_2147,In_443,In_122);
nor U2148 (N_2148,In_508,In_355);
or U2149 (N_2149,In_128,In_653);
or U2150 (N_2150,In_364,In_149);
nor U2151 (N_2151,In_561,In_234);
nand U2152 (N_2152,In_41,In_222);
nor U2153 (N_2153,In_467,In_555);
nand U2154 (N_2154,In_219,In_613);
or U2155 (N_2155,In_286,In_710);
or U2156 (N_2156,In_547,In_363);
and U2157 (N_2157,In_187,In_120);
or U2158 (N_2158,In_238,In_65);
or U2159 (N_2159,In_531,In_441);
and U2160 (N_2160,In_500,In_113);
or U2161 (N_2161,In_226,In_372);
or U2162 (N_2162,In_431,In_557);
nor U2163 (N_2163,In_160,In_273);
xor U2164 (N_2164,In_133,In_479);
and U2165 (N_2165,In_195,In_550);
xnor U2166 (N_2166,In_426,In_49);
nand U2167 (N_2167,In_417,In_326);
nand U2168 (N_2168,In_61,In_692);
or U2169 (N_2169,In_665,In_515);
nor U2170 (N_2170,In_347,In_314);
and U2171 (N_2171,In_340,In_211);
xnor U2172 (N_2172,In_516,In_732);
nor U2173 (N_2173,In_670,In_420);
nand U2174 (N_2174,In_572,In_596);
nand U2175 (N_2175,In_691,In_670);
xor U2176 (N_2176,In_651,In_577);
and U2177 (N_2177,In_269,In_452);
or U2178 (N_2178,In_544,In_26);
nand U2179 (N_2179,In_471,In_253);
or U2180 (N_2180,In_570,In_501);
and U2181 (N_2181,In_174,In_245);
nand U2182 (N_2182,In_338,In_629);
or U2183 (N_2183,In_99,In_189);
and U2184 (N_2184,In_167,In_1);
or U2185 (N_2185,In_461,In_68);
nand U2186 (N_2186,In_269,In_706);
or U2187 (N_2187,In_569,In_128);
or U2188 (N_2188,In_687,In_607);
or U2189 (N_2189,In_586,In_374);
nor U2190 (N_2190,In_683,In_172);
and U2191 (N_2191,In_312,In_349);
nand U2192 (N_2192,In_241,In_556);
nand U2193 (N_2193,In_635,In_388);
xnor U2194 (N_2194,In_260,In_172);
and U2195 (N_2195,In_454,In_746);
nand U2196 (N_2196,In_661,In_680);
and U2197 (N_2197,In_287,In_749);
and U2198 (N_2198,In_748,In_35);
and U2199 (N_2199,In_637,In_375);
nor U2200 (N_2200,In_703,In_578);
and U2201 (N_2201,In_477,In_525);
and U2202 (N_2202,In_248,In_348);
nor U2203 (N_2203,In_490,In_203);
or U2204 (N_2204,In_289,In_419);
xnor U2205 (N_2205,In_230,In_635);
nor U2206 (N_2206,In_241,In_446);
nor U2207 (N_2207,In_544,In_617);
nor U2208 (N_2208,In_296,In_306);
nand U2209 (N_2209,In_645,In_91);
nor U2210 (N_2210,In_15,In_567);
xor U2211 (N_2211,In_691,In_520);
nand U2212 (N_2212,In_634,In_452);
nor U2213 (N_2213,In_599,In_370);
xnor U2214 (N_2214,In_625,In_276);
nor U2215 (N_2215,In_635,In_220);
nand U2216 (N_2216,In_548,In_284);
or U2217 (N_2217,In_480,In_605);
xnor U2218 (N_2218,In_426,In_525);
nand U2219 (N_2219,In_255,In_278);
nor U2220 (N_2220,In_97,In_542);
or U2221 (N_2221,In_156,In_538);
or U2222 (N_2222,In_653,In_442);
nand U2223 (N_2223,In_556,In_20);
xor U2224 (N_2224,In_582,In_254);
or U2225 (N_2225,In_1,In_457);
nor U2226 (N_2226,In_408,In_487);
or U2227 (N_2227,In_221,In_211);
nand U2228 (N_2228,In_443,In_169);
or U2229 (N_2229,In_709,In_283);
xnor U2230 (N_2230,In_586,In_556);
nand U2231 (N_2231,In_264,In_209);
and U2232 (N_2232,In_454,In_248);
or U2233 (N_2233,In_152,In_112);
nor U2234 (N_2234,In_64,In_474);
and U2235 (N_2235,In_590,In_372);
nor U2236 (N_2236,In_375,In_89);
nand U2237 (N_2237,In_283,In_21);
and U2238 (N_2238,In_741,In_267);
nor U2239 (N_2239,In_401,In_665);
nor U2240 (N_2240,In_187,In_319);
nor U2241 (N_2241,In_702,In_197);
and U2242 (N_2242,In_248,In_57);
nand U2243 (N_2243,In_382,In_0);
and U2244 (N_2244,In_132,In_44);
or U2245 (N_2245,In_478,In_496);
nor U2246 (N_2246,In_288,In_306);
and U2247 (N_2247,In_528,In_509);
nand U2248 (N_2248,In_736,In_395);
nand U2249 (N_2249,In_105,In_95);
xor U2250 (N_2250,In_588,In_136);
and U2251 (N_2251,In_20,In_507);
xnor U2252 (N_2252,In_338,In_649);
nand U2253 (N_2253,In_376,In_112);
and U2254 (N_2254,In_546,In_540);
or U2255 (N_2255,In_116,In_579);
or U2256 (N_2256,In_542,In_268);
xor U2257 (N_2257,In_539,In_692);
or U2258 (N_2258,In_469,In_618);
or U2259 (N_2259,In_224,In_738);
and U2260 (N_2260,In_7,In_237);
and U2261 (N_2261,In_122,In_308);
nor U2262 (N_2262,In_103,In_609);
xor U2263 (N_2263,In_377,In_234);
or U2264 (N_2264,In_595,In_328);
or U2265 (N_2265,In_485,In_153);
and U2266 (N_2266,In_340,In_540);
or U2267 (N_2267,In_177,In_564);
or U2268 (N_2268,In_112,In_708);
nor U2269 (N_2269,In_674,In_381);
and U2270 (N_2270,In_703,In_695);
or U2271 (N_2271,In_406,In_531);
nor U2272 (N_2272,In_645,In_35);
and U2273 (N_2273,In_742,In_109);
or U2274 (N_2274,In_538,In_167);
and U2275 (N_2275,In_659,In_621);
or U2276 (N_2276,In_75,In_6);
nand U2277 (N_2277,In_661,In_438);
or U2278 (N_2278,In_257,In_679);
nor U2279 (N_2279,In_502,In_661);
nor U2280 (N_2280,In_135,In_208);
and U2281 (N_2281,In_431,In_213);
nor U2282 (N_2282,In_3,In_590);
nor U2283 (N_2283,In_208,In_226);
xor U2284 (N_2284,In_573,In_119);
nor U2285 (N_2285,In_239,In_538);
nor U2286 (N_2286,In_4,In_204);
nor U2287 (N_2287,In_103,In_657);
and U2288 (N_2288,In_530,In_293);
nand U2289 (N_2289,In_544,In_492);
xnor U2290 (N_2290,In_526,In_42);
xnor U2291 (N_2291,In_279,In_149);
and U2292 (N_2292,In_711,In_649);
xnor U2293 (N_2293,In_554,In_483);
nand U2294 (N_2294,In_550,In_362);
or U2295 (N_2295,In_570,In_511);
or U2296 (N_2296,In_281,In_303);
nor U2297 (N_2297,In_110,In_286);
nand U2298 (N_2298,In_651,In_355);
and U2299 (N_2299,In_668,In_408);
and U2300 (N_2300,In_735,In_456);
nor U2301 (N_2301,In_26,In_253);
xnor U2302 (N_2302,In_112,In_91);
xor U2303 (N_2303,In_127,In_670);
and U2304 (N_2304,In_351,In_745);
or U2305 (N_2305,In_92,In_512);
nand U2306 (N_2306,In_377,In_23);
or U2307 (N_2307,In_434,In_610);
and U2308 (N_2308,In_585,In_314);
or U2309 (N_2309,In_547,In_384);
or U2310 (N_2310,In_281,In_623);
nand U2311 (N_2311,In_736,In_573);
xnor U2312 (N_2312,In_96,In_228);
and U2313 (N_2313,In_626,In_332);
nand U2314 (N_2314,In_585,In_615);
or U2315 (N_2315,In_724,In_528);
nand U2316 (N_2316,In_506,In_648);
xor U2317 (N_2317,In_326,In_627);
and U2318 (N_2318,In_597,In_686);
nor U2319 (N_2319,In_700,In_563);
nand U2320 (N_2320,In_684,In_165);
nand U2321 (N_2321,In_243,In_348);
and U2322 (N_2322,In_160,In_320);
and U2323 (N_2323,In_340,In_148);
or U2324 (N_2324,In_514,In_493);
xnor U2325 (N_2325,In_574,In_406);
nor U2326 (N_2326,In_427,In_323);
or U2327 (N_2327,In_697,In_165);
nor U2328 (N_2328,In_165,In_601);
or U2329 (N_2329,In_291,In_98);
nor U2330 (N_2330,In_245,In_676);
nand U2331 (N_2331,In_244,In_465);
and U2332 (N_2332,In_295,In_372);
nand U2333 (N_2333,In_589,In_511);
or U2334 (N_2334,In_211,In_582);
or U2335 (N_2335,In_236,In_249);
and U2336 (N_2336,In_729,In_533);
nand U2337 (N_2337,In_527,In_158);
nand U2338 (N_2338,In_82,In_130);
nand U2339 (N_2339,In_660,In_254);
and U2340 (N_2340,In_588,In_410);
and U2341 (N_2341,In_549,In_210);
and U2342 (N_2342,In_638,In_632);
or U2343 (N_2343,In_500,In_699);
nor U2344 (N_2344,In_532,In_430);
and U2345 (N_2345,In_577,In_132);
and U2346 (N_2346,In_95,In_598);
or U2347 (N_2347,In_672,In_345);
and U2348 (N_2348,In_105,In_585);
or U2349 (N_2349,In_148,In_334);
nor U2350 (N_2350,In_499,In_190);
nand U2351 (N_2351,In_714,In_99);
nor U2352 (N_2352,In_718,In_384);
nand U2353 (N_2353,In_383,In_607);
xnor U2354 (N_2354,In_449,In_744);
and U2355 (N_2355,In_183,In_102);
nor U2356 (N_2356,In_245,In_253);
and U2357 (N_2357,In_612,In_480);
xor U2358 (N_2358,In_285,In_182);
nand U2359 (N_2359,In_606,In_560);
nor U2360 (N_2360,In_656,In_284);
and U2361 (N_2361,In_203,In_498);
nand U2362 (N_2362,In_168,In_542);
nor U2363 (N_2363,In_406,In_397);
nor U2364 (N_2364,In_617,In_32);
and U2365 (N_2365,In_222,In_503);
or U2366 (N_2366,In_313,In_626);
nor U2367 (N_2367,In_435,In_222);
nor U2368 (N_2368,In_29,In_15);
nand U2369 (N_2369,In_65,In_400);
and U2370 (N_2370,In_217,In_280);
and U2371 (N_2371,In_87,In_472);
or U2372 (N_2372,In_283,In_23);
or U2373 (N_2373,In_346,In_609);
nand U2374 (N_2374,In_122,In_662);
xor U2375 (N_2375,In_105,In_719);
nand U2376 (N_2376,In_677,In_429);
and U2377 (N_2377,In_505,In_744);
nand U2378 (N_2378,In_557,In_700);
nor U2379 (N_2379,In_490,In_493);
or U2380 (N_2380,In_81,In_746);
and U2381 (N_2381,In_308,In_539);
and U2382 (N_2382,In_535,In_402);
nor U2383 (N_2383,In_403,In_736);
or U2384 (N_2384,In_100,In_515);
nand U2385 (N_2385,In_167,In_430);
nor U2386 (N_2386,In_681,In_664);
xnor U2387 (N_2387,In_426,In_324);
nor U2388 (N_2388,In_581,In_310);
nor U2389 (N_2389,In_248,In_739);
and U2390 (N_2390,In_268,In_252);
xnor U2391 (N_2391,In_214,In_508);
or U2392 (N_2392,In_723,In_731);
or U2393 (N_2393,In_373,In_555);
nand U2394 (N_2394,In_388,In_737);
nor U2395 (N_2395,In_115,In_704);
xnor U2396 (N_2396,In_463,In_69);
and U2397 (N_2397,In_685,In_687);
nand U2398 (N_2398,In_602,In_632);
and U2399 (N_2399,In_484,In_96);
and U2400 (N_2400,In_257,In_675);
or U2401 (N_2401,In_619,In_310);
nor U2402 (N_2402,In_324,In_607);
nand U2403 (N_2403,In_187,In_689);
and U2404 (N_2404,In_375,In_282);
or U2405 (N_2405,In_664,In_678);
or U2406 (N_2406,In_250,In_516);
or U2407 (N_2407,In_123,In_563);
and U2408 (N_2408,In_77,In_626);
nor U2409 (N_2409,In_565,In_396);
nand U2410 (N_2410,In_111,In_23);
nand U2411 (N_2411,In_93,In_15);
and U2412 (N_2412,In_296,In_694);
or U2413 (N_2413,In_661,In_545);
or U2414 (N_2414,In_492,In_45);
or U2415 (N_2415,In_242,In_730);
or U2416 (N_2416,In_401,In_55);
nor U2417 (N_2417,In_107,In_246);
nand U2418 (N_2418,In_744,In_355);
xnor U2419 (N_2419,In_719,In_554);
and U2420 (N_2420,In_213,In_671);
xor U2421 (N_2421,In_107,In_354);
nor U2422 (N_2422,In_128,In_221);
nand U2423 (N_2423,In_128,In_1);
and U2424 (N_2424,In_45,In_194);
or U2425 (N_2425,In_603,In_595);
or U2426 (N_2426,In_606,In_113);
or U2427 (N_2427,In_533,In_297);
and U2428 (N_2428,In_493,In_74);
or U2429 (N_2429,In_469,In_103);
nor U2430 (N_2430,In_4,In_108);
nand U2431 (N_2431,In_42,In_274);
and U2432 (N_2432,In_72,In_158);
or U2433 (N_2433,In_288,In_23);
xor U2434 (N_2434,In_344,In_361);
nand U2435 (N_2435,In_298,In_376);
nand U2436 (N_2436,In_188,In_723);
and U2437 (N_2437,In_455,In_357);
nor U2438 (N_2438,In_32,In_438);
and U2439 (N_2439,In_432,In_9);
nand U2440 (N_2440,In_83,In_521);
or U2441 (N_2441,In_397,In_487);
or U2442 (N_2442,In_216,In_591);
and U2443 (N_2443,In_52,In_296);
or U2444 (N_2444,In_652,In_370);
nor U2445 (N_2445,In_23,In_549);
nor U2446 (N_2446,In_161,In_191);
or U2447 (N_2447,In_401,In_691);
nor U2448 (N_2448,In_452,In_134);
nor U2449 (N_2449,In_377,In_610);
or U2450 (N_2450,In_483,In_572);
nor U2451 (N_2451,In_258,In_618);
xor U2452 (N_2452,In_309,In_542);
xnor U2453 (N_2453,In_428,In_227);
nor U2454 (N_2454,In_460,In_727);
nor U2455 (N_2455,In_108,In_2);
and U2456 (N_2456,In_301,In_362);
nor U2457 (N_2457,In_84,In_421);
or U2458 (N_2458,In_257,In_709);
nor U2459 (N_2459,In_325,In_635);
or U2460 (N_2460,In_423,In_480);
and U2461 (N_2461,In_699,In_413);
or U2462 (N_2462,In_477,In_489);
xnor U2463 (N_2463,In_57,In_399);
or U2464 (N_2464,In_457,In_397);
and U2465 (N_2465,In_734,In_634);
nor U2466 (N_2466,In_187,In_521);
nor U2467 (N_2467,In_150,In_83);
nor U2468 (N_2468,In_497,In_544);
nand U2469 (N_2469,In_222,In_316);
xor U2470 (N_2470,In_489,In_716);
or U2471 (N_2471,In_596,In_179);
nand U2472 (N_2472,In_288,In_214);
nand U2473 (N_2473,In_359,In_196);
or U2474 (N_2474,In_431,In_76);
nor U2475 (N_2475,In_192,In_704);
or U2476 (N_2476,In_36,In_593);
and U2477 (N_2477,In_171,In_423);
and U2478 (N_2478,In_551,In_708);
and U2479 (N_2479,In_292,In_455);
nor U2480 (N_2480,In_636,In_375);
nor U2481 (N_2481,In_116,In_8);
nand U2482 (N_2482,In_516,In_709);
and U2483 (N_2483,In_158,In_703);
nand U2484 (N_2484,In_61,In_487);
nand U2485 (N_2485,In_670,In_688);
and U2486 (N_2486,In_645,In_687);
and U2487 (N_2487,In_431,In_8);
xor U2488 (N_2488,In_121,In_432);
or U2489 (N_2489,In_510,In_202);
nor U2490 (N_2490,In_523,In_680);
or U2491 (N_2491,In_717,In_168);
nor U2492 (N_2492,In_488,In_334);
nand U2493 (N_2493,In_368,In_692);
nand U2494 (N_2494,In_729,In_71);
and U2495 (N_2495,In_383,In_163);
nand U2496 (N_2496,In_485,In_39);
nor U2497 (N_2497,In_617,In_49);
or U2498 (N_2498,In_723,In_631);
nor U2499 (N_2499,In_722,In_689);
or U2500 (N_2500,N_1745,N_1336);
or U2501 (N_2501,N_2103,N_160);
nor U2502 (N_2502,N_1510,N_2377);
and U2503 (N_2503,N_2401,N_1008);
nor U2504 (N_2504,N_957,N_1825);
or U2505 (N_2505,N_582,N_2381);
and U2506 (N_2506,N_2244,N_2288);
nor U2507 (N_2507,N_301,N_555);
nand U2508 (N_2508,N_657,N_1175);
nor U2509 (N_2509,N_950,N_2264);
and U2510 (N_2510,N_2398,N_238);
nand U2511 (N_2511,N_2125,N_574);
or U2512 (N_2512,N_723,N_2310);
xnor U2513 (N_2513,N_1562,N_115);
and U2514 (N_2514,N_1579,N_862);
nand U2515 (N_2515,N_2253,N_2388);
nor U2516 (N_2516,N_2009,N_1381);
nand U2517 (N_2517,N_2224,N_2087);
and U2518 (N_2518,N_1376,N_528);
nand U2519 (N_2519,N_350,N_763);
nor U2520 (N_2520,N_1004,N_2221);
nor U2521 (N_2521,N_1833,N_822);
nand U2522 (N_2522,N_2022,N_2013);
xnor U2523 (N_2523,N_2171,N_821);
nand U2524 (N_2524,N_1598,N_664);
or U2525 (N_2525,N_1076,N_1091);
nand U2526 (N_2526,N_1209,N_534);
nand U2527 (N_2527,N_721,N_403);
or U2528 (N_2528,N_2240,N_522);
nor U2529 (N_2529,N_316,N_1742);
and U2530 (N_2530,N_1037,N_2234);
nor U2531 (N_2531,N_1962,N_2219);
nor U2532 (N_2532,N_1026,N_652);
nand U2533 (N_2533,N_111,N_1186);
or U2534 (N_2534,N_711,N_1880);
nor U2535 (N_2535,N_1587,N_2043);
nand U2536 (N_2536,N_1838,N_938);
and U2537 (N_2537,N_1608,N_632);
xor U2538 (N_2538,N_1786,N_1721);
xor U2539 (N_2539,N_145,N_1372);
and U2540 (N_2540,N_333,N_490);
nor U2541 (N_2541,N_1214,N_1911);
nor U2542 (N_2542,N_865,N_891);
and U2543 (N_2543,N_1730,N_2044);
nor U2544 (N_2544,N_1736,N_2050);
and U2545 (N_2545,N_2478,N_2471);
and U2546 (N_2546,N_2448,N_2169);
or U2547 (N_2547,N_1047,N_643);
and U2548 (N_2548,N_1610,N_52);
or U2549 (N_2549,N_36,N_182);
and U2550 (N_2550,N_1364,N_1671);
xnor U2551 (N_2551,N_1177,N_1319);
nor U2552 (N_2552,N_1399,N_1571);
or U2553 (N_2553,N_1380,N_152);
nor U2554 (N_2554,N_1808,N_880);
xnor U2555 (N_2555,N_307,N_2024);
xor U2556 (N_2556,N_712,N_927);
and U2557 (N_2557,N_2294,N_1289);
xnor U2558 (N_2558,N_2152,N_2198);
nor U2559 (N_2559,N_1614,N_16);
nand U2560 (N_2560,N_2162,N_746);
nor U2561 (N_2561,N_1609,N_287);
xor U2562 (N_2562,N_1233,N_461);
or U2563 (N_2563,N_493,N_349);
nand U2564 (N_2564,N_1797,N_737);
nor U2565 (N_2565,N_743,N_1052);
nand U2566 (N_2566,N_1750,N_964);
and U2567 (N_2567,N_1088,N_903);
or U2568 (N_2568,N_179,N_1207);
nor U2569 (N_2569,N_703,N_1492);
nor U2570 (N_2570,N_398,N_788);
nand U2571 (N_2571,N_1035,N_1639);
xnor U2572 (N_2572,N_2480,N_270);
and U2573 (N_2573,N_2469,N_852);
nand U2574 (N_2574,N_1877,N_654);
nor U2575 (N_2575,N_1149,N_1862);
or U2576 (N_2576,N_1988,N_2106);
nand U2577 (N_2577,N_1627,N_1200);
xor U2578 (N_2578,N_91,N_2371);
nor U2579 (N_2579,N_2322,N_1078);
nor U2580 (N_2580,N_2316,N_66);
and U2581 (N_2581,N_2444,N_1161);
and U2582 (N_2582,N_1813,N_1092);
nand U2583 (N_2583,N_1955,N_2339);
nor U2584 (N_2584,N_363,N_277);
or U2585 (N_2585,N_974,N_1171);
xor U2586 (N_2586,N_1728,N_1107);
and U2587 (N_2587,N_2456,N_736);
or U2588 (N_2588,N_1507,N_1864);
xnor U2589 (N_2589,N_760,N_45);
nand U2590 (N_2590,N_835,N_190);
and U2591 (N_2591,N_2001,N_1892);
nand U2592 (N_2592,N_2386,N_607);
nand U2593 (N_2593,N_569,N_2428);
nor U2594 (N_2594,N_221,N_186);
or U2595 (N_2595,N_629,N_876);
nand U2596 (N_2596,N_444,N_188);
nor U2597 (N_2597,N_2158,N_2399);
nor U2598 (N_2598,N_617,N_177);
nand U2599 (N_2599,N_1406,N_1592);
or U2600 (N_2600,N_494,N_1909);
nor U2601 (N_2601,N_1857,N_2031);
nor U2602 (N_2602,N_1606,N_706);
xnor U2603 (N_2603,N_244,N_1675);
or U2604 (N_2604,N_1112,N_2166);
and U2605 (N_2605,N_22,N_2220);
and U2606 (N_2606,N_1603,N_26);
nor U2607 (N_2607,N_1656,N_1338);
and U2608 (N_2608,N_1873,N_1240);
and U2609 (N_2609,N_2475,N_2281);
or U2610 (N_2610,N_1600,N_41);
or U2611 (N_2611,N_304,N_396);
or U2612 (N_2612,N_1663,N_914);
nor U2613 (N_2613,N_2330,N_1064);
nand U2614 (N_2614,N_1535,N_2095);
nor U2615 (N_2615,N_1071,N_8);
nor U2616 (N_2616,N_1520,N_1999);
and U2617 (N_2617,N_1926,N_1767);
nand U2618 (N_2618,N_457,N_1717);
nand U2619 (N_2619,N_738,N_949);
nand U2620 (N_2620,N_1053,N_1096);
xnor U2621 (N_2621,N_2473,N_410);
or U2622 (N_2622,N_2053,N_806);
and U2623 (N_2623,N_171,N_1538);
and U2624 (N_2624,N_1811,N_1463);
or U2625 (N_2625,N_2216,N_1426);
nand U2626 (N_2626,N_1132,N_1036);
and U2627 (N_2627,N_1824,N_463);
nand U2628 (N_2628,N_40,N_2062);
nand U2629 (N_2629,N_2236,N_527);
or U2630 (N_2630,N_1396,N_1324);
and U2631 (N_2631,N_904,N_2445);
nand U2632 (N_2632,N_668,N_1849);
nor U2633 (N_2633,N_861,N_925);
xnor U2634 (N_2634,N_1701,N_1589);
nor U2635 (N_2635,N_133,N_722);
nand U2636 (N_2636,N_83,N_2078);
or U2637 (N_2637,N_1753,N_2483);
xor U2638 (N_2638,N_2183,N_2276);
xnor U2639 (N_2639,N_2429,N_198);
and U2640 (N_2640,N_1853,N_1693);
xnor U2641 (N_2641,N_954,N_1633);
nor U2642 (N_2642,N_1323,N_1586);
nor U2643 (N_2643,N_1859,N_2085);
nor U2644 (N_2644,N_2482,N_536);
xnor U2645 (N_2645,N_948,N_230);
nor U2646 (N_2646,N_757,N_1073);
nor U2647 (N_2647,N_1201,N_2061);
and U2648 (N_2648,N_2477,N_597);
or U2649 (N_2649,N_1144,N_2476);
or U2650 (N_2650,N_2467,N_749);
and U2651 (N_2651,N_1795,N_1006);
nand U2652 (N_2652,N_1789,N_69);
and U2653 (N_2653,N_877,N_2360);
or U2654 (N_2654,N_1652,N_1502);
nand U2655 (N_2655,N_2091,N_35);
nor U2656 (N_2656,N_2203,N_1725);
and U2657 (N_2657,N_2327,N_1832);
and U2658 (N_2658,N_2283,N_2359);
nor U2659 (N_2659,N_933,N_1147);
nand U2660 (N_2660,N_2334,N_1653);
nand U2661 (N_2661,N_2286,N_1162);
and U2662 (N_2662,N_1125,N_2116);
nand U2663 (N_2663,N_1526,N_1418);
nand U2664 (N_2664,N_2020,N_1852);
nand U2665 (N_2665,N_1109,N_773);
or U2666 (N_2666,N_382,N_1749);
nand U2667 (N_2667,N_1844,N_1398);
nand U2668 (N_2668,N_1952,N_838);
and U2669 (N_2669,N_2356,N_1294);
xor U2670 (N_2670,N_358,N_2173);
and U2671 (N_2671,N_584,N_2262);
nor U2672 (N_2672,N_850,N_1706);
nor U2673 (N_2673,N_264,N_1575);
or U2674 (N_2674,N_843,N_430);
nor U2675 (N_2675,N_1413,N_480);
or U2676 (N_2676,N_618,N_1970);
xnor U2677 (N_2677,N_2256,N_1645);
and U2678 (N_2678,N_2493,N_1243);
xor U2679 (N_2679,N_2351,N_2230);
and U2680 (N_2680,N_405,N_951);
and U2681 (N_2681,N_2113,N_899);
or U2682 (N_2682,N_745,N_248);
nor U2683 (N_2683,N_104,N_110);
and U2684 (N_2684,N_1508,N_1607);
and U2685 (N_2685,N_1868,N_353);
or U2686 (N_2686,N_1395,N_1595);
nor U2687 (N_2687,N_2122,N_1889);
and U2688 (N_2688,N_946,N_550);
nor U2689 (N_2689,N_941,N_795);
nand U2690 (N_2690,N_1130,N_408);
nor U2691 (N_2691,N_693,N_49);
or U2692 (N_2692,N_691,N_2098);
nor U2693 (N_2693,N_11,N_1194);
and U2694 (N_2694,N_646,N_1156);
xor U2695 (N_2695,N_174,N_1099);
nor U2696 (N_2696,N_2079,N_2425);
nor U2697 (N_2697,N_1192,N_2238);
nand U2698 (N_2698,N_300,N_639);
nor U2699 (N_2699,N_1814,N_709);
or U2700 (N_2700,N_1541,N_1963);
and U2701 (N_2701,N_165,N_2023);
or U2702 (N_2702,N_208,N_671);
and U2703 (N_2703,N_21,N_537);
nor U2704 (N_2704,N_1257,N_934);
nor U2705 (N_2705,N_59,N_1943);
or U2706 (N_2706,N_1895,N_2352);
nor U2707 (N_2707,N_1225,N_2128);
and U2708 (N_2708,N_1993,N_585);
nor U2709 (N_2709,N_355,N_1268);
and U2710 (N_2710,N_1618,N_168);
nand U2711 (N_2711,N_1643,N_261);
and U2712 (N_2712,N_1779,N_2350);
nor U2713 (N_2713,N_972,N_1140);
nand U2714 (N_2714,N_678,N_624);
nand U2715 (N_2715,N_1906,N_46);
xnor U2716 (N_2716,N_1439,N_1114);
and U2717 (N_2717,N_1856,N_2227);
nand U2718 (N_2718,N_181,N_793);
nor U2719 (N_2719,N_1776,N_1945);
or U2720 (N_2720,N_2075,N_784);
and U2721 (N_2721,N_718,N_1145);
and U2722 (N_2722,N_1001,N_1165);
nand U2723 (N_2723,N_660,N_1641);
xor U2724 (N_2724,N_2189,N_2083);
nand U2725 (N_2725,N_2251,N_1922);
nand U2726 (N_2726,N_1404,N_692);
nand U2727 (N_2727,N_622,N_1069);
and U2728 (N_2728,N_2414,N_176);
nor U2729 (N_2729,N_1573,N_2474);
and U2730 (N_2730,N_2285,N_2046);
and U2731 (N_2731,N_251,N_1479);
nand U2732 (N_2732,N_78,N_1707);
or U2733 (N_2733,N_467,N_869);
xor U2734 (N_2734,N_565,N_859);
xor U2735 (N_2735,N_1084,N_1456);
nand U2736 (N_2736,N_1460,N_1664);
and U2737 (N_2737,N_71,N_762);
nand U2738 (N_2738,N_436,N_583);
or U2739 (N_2739,N_328,N_282);
nand U2740 (N_2740,N_364,N_2051);
nor U2741 (N_2741,N_337,N_223);
and U2742 (N_2742,N_438,N_2287);
nand U2743 (N_2743,N_1138,N_1483);
nor U2744 (N_2744,N_2435,N_1155);
nor U2745 (N_2745,N_779,N_1847);
or U2746 (N_2746,N_605,N_1139);
or U2747 (N_2747,N_663,N_1836);
and U2748 (N_2748,N_2226,N_1699);
and U2749 (N_2749,N_295,N_2324);
nor U2750 (N_2750,N_978,N_1260);
nand U2751 (N_2751,N_983,N_923);
or U2752 (N_2752,N_1710,N_1254);
nand U2753 (N_2753,N_2459,N_94);
or U2754 (N_2754,N_2084,N_1668);
nor U2755 (N_2755,N_2120,N_1489);
nor U2756 (N_2756,N_404,N_23);
or U2757 (N_2757,N_1111,N_1017);
or U2758 (N_2758,N_766,N_219);
nand U2759 (N_2759,N_125,N_807);
nand U2760 (N_2760,N_1075,N_1764);
or U2761 (N_2761,N_412,N_1477);
xor U2762 (N_2762,N_1676,N_2003);
nor U2763 (N_2763,N_871,N_95);
xnor U2764 (N_2764,N_2011,N_330);
or U2765 (N_2765,N_2194,N_714);
nor U2766 (N_2766,N_370,N_1119);
nor U2767 (N_2767,N_982,N_518);
and U2768 (N_2768,N_1235,N_921);
or U2769 (N_2769,N_1224,N_540);
nand U2770 (N_2770,N_342,N_1085);
nand U2771 (N_2771,N_2118,N_554);
and U2772 (N_2772,N_478,N_1842);
nor U2773 (N_2773,N_1431,N_28);
xnor U2774 (N_2774,N_1291,N_39);
and U2775 (N_2775,N_68,N_1079);
and U2776 (N_2776,N_427,N_1444);
nor U2777 (N_2777,N_361,N_2358);
nor U2778 (N_2778,N_2153,N_936);
xor U2779 (N_2779,N_2277,N_2060);
nor U2780 (N_2780,N_484,N_1995);
xor U2781 (N_2781,N_228,N_1785);
nand U2782 (N_2782,N_523,N_2252);
and U2783 (N_2783,N_2298,N_486);
or U2784 (N_2784,N_1584,N_2301);
nor U2785 (N_2785,N_1060,N_1488);
nor U2786 (N_2786,N_827,N_1296);
nand U2787 (N_2787,N_2034,N_1553);
nor U2788 (N_2788,N_620,N_836);
or U2789 (N_2789,N_415,N_546);
nor U2790 (N_2790,N_1160,N_1232);
or U2791 (N_2791,N_2415,N_775);
or U2792 (N_2792,N_18,N_1977);
nand U2793 (N_2793,N_659,N_2434);
and U2794 (N_2794,N_10,N_1360);
nor U2795 (N_2795,N_258,N_602);
nor U2796 (N_2796,N_1694,N_1992);
and U2797 (N_2797,N_2133,N_1283);
nor U2798 (N_2798,N_92,N_1419);
and U2799 (N_2799,N_846,N_102);
nor U2800 (N_2800,N_82,N_858);
nand U2801 (N_2801,N_1027,N_1332);
and U2802 (N_2802,N_2259,N_1950);
nand U2803 (N_2803,N_1490,N_2320);
xor U2804 (N_2804,N_2232,N_2270);
nand U2805 (N_2805,N_625,N_1495);
and U2806 (N_2806,N_2427,N_2041);
nand U2807 (N_2807,N_1890,N_591);
nor U2808 (N_2808,N_227,N_720);
nand U2809 (N_2809,N_1054,N_1465);
or U2810 (N_2810,N_1588,N_1978);
and U2811 (N_2811,N_2154,N_2010);
and U2812 (N_2812,N_1215,N_1000);
or U2813 (N_2813,N_1961,N_854);
or U2814 (N_2814,N_1702,N_2181);
or U2815 (N_2815,N_1255,N_2250);
and U2816 (N_2816,N_1131,N_1407);
nor U2817 (N_2817,N_1397,N_2172);
nor U2818 (N_2818,N_42,N_1496);
and U2819 (N_2819,N_1025,N_2484);
xnor U2820 (N_2820,N_1931,N_553);
and U2821 (N_2821,N_2443,N_906);
nand U2822 (N_2822,N_1441,N_2109);
nor U2823 (N_2823,N_1427,N_1270);
nand U2824 (N_2824,N_814,N_1744);
nand U2825 (N_2825,N_772,N_1732);
nand U2826 (N_2826,N_767,N_20);
or U2827 (N_2827,N_1285,N_699);
and U2828 (N_2828,N_105,N_2247);
nand U2829 (N_2829,N_2197,N_2059);
or U2830 (N_2830,N_2054,N_1547);
and U2831 (N_2831,N_1980,N_1433);
or U2832 (N_2832,N_1470,N_2384);
nor U2833 (N_2833,N_2317,N_1485);
xnor U2834 (N_2834,N_675,N_810);
nand U2835 (N_2835,N_634,N_1846);
or U2836 (N_2836,N_1946,N_1590);
or U2837 (N_2837,N_1392,N_524);
nand U2838 (N_2838,N_2290,N_103);
or U2839 (N_2839,N_1282,N_1902);
nor U2840 (N_2840,N_291,N_1964);
nor U2841 (N_2841,N_774,N_2184);
or U2842 (N_2842,N_2159,N_1660);
nor U2843 (N_2843,N_1518,N_2305);
or U2844 (N_2844,N_323,N_588);
and U2845 (N_2845,N_447,N_1297);
and U2846 (N_2846,N_544,N_2392);
xnor U2847 (N_2847,N_1793,N_1379);
nor U2848 (N_2848,N_2265,N_2295);
or U2849 (N_2849,N_2257,N_2405);
nor U2850 (N_2850,N_1712,N_794);
nor U2851 (N_2851,N_1637,N_193);
nand U2852 (N_2852,N_320,N_191);
or U2853 (N_2853,N_621,N_579);
and U2854 (N_2854,N_2457,N_1913);
or U2855 (N_2855,N_1059,N_1686);
or U2856 (N_2856,N_2312,N_2329);
or U2857 (N_2857,N_1472,N_2037);
nand U2858 (N_2858,N_321,N_2182);
or U2859 (N_2859,N_991,N_1788);
nand U2860 (N_2860,N_820,N_1030);
nand U2861 (N_2861,N_677,N_389);
nand U2862 (N_2862,N_2389,N_481);
and U2863 (N_2863,N_1436,N_860);
or U2864 (N_2864,N_2096,N_2307);
and U2865 (N_2865,N_2354,N_817);
or U2866 (N_2866,N_944,N_1416);
or U2867 (N_2867,N_85,N_1141);
or U2868 (N_2868,N_2292,N_1122);
and U2869 (N_2869,N_2180,N_1661);
nand U2870 (N_2870,N_2325,N_2077);
xnor U2871 (N_2871,N_1312,N_1947);
nor U2872 (N_2872,N_1056,N_2357);
and U2873 (N_2873,N_1208,N_1594);
xor U2874 (N_2874,N_2452,N_804);
or U2875 (N_2875,N_1576,N_882);
and U2876 (N_2876,N_1128,N_360);
nor U2877 (N_2877,N_1623,N_1135);
nor U2878 (N_2878,N_556,N_799);
nor U2879 (N_2879,N_833,N_246);
and U2880 (N_2880,N_159,N_729);
nor U2881 (N_2881,N_898,N_1183);
nand U2882 (N_2882,N_651,N_1043);
nand U2883 (N_2883,N_255,N_765);
nand U2884 (N_2884,N_637,N_612);
xor U2885 (N_2885,N_2461,N_2313);
and U2886 (N_2886,N_2174,N_756);
or U2887 (N_2887,N_1309,N_1932);
nor U2888 (N_2888,N_1173,N_302);
or U2889 (N_2889,N_521,N_2396);
nand U2890 (N_2890,N_840,N_520);
nand U2891 (N_2891,N_263,N_672);
xnor U2892 (N_2892,N_900,N_2291);
or U2893 (N_2893,N_768,N_1040);
or U2894 (N_2894,N_202,N_30);
nor U2895 (N_2895,N_1998,N_2261);
or U2896 (N_2896,N_1835,N_2245);
and U2897 (N_2897,N_1956,N_506);
or U2898 (N_2898,N_1718,N_1377);
nor U2899 (N_2899,N_1415,N_236);
or U2900 (N_2900,N_378,N_1041);
nand U2901 (N_2901,N_894,N_1601);
nand U2902 (N_2902,N_281,N_1790);
xnor U2903 (N_2903,N_2165,N_939);
xor U2904 (N_2904,N_770,N_510);
nand U2905 (N_2905,N_2460,N_252);
nand U2906 (N_2906,N_2047,N_1654);
nor U2907 (N_2907,N_1839,N_1615);
nand U2908 (N_2908,N_464,N_2092);
xnor U2909 (N_2909,N_2488,N_568);
nand U2910 (N_2910,N_2055,N_1672);
nand U2911 (N_2911,N_379,N_593);
and U2912 (N_2912,N_99,N_2404);
or U2913 (N_2913,N_93,N_1024);
or U2914 (N_2914,N_1727,N_1443);
xor U2915 (N_2915,N_1755,N_2453);
or U2916 (N_2916,N_1534,N_2437);
and U2917 (N_2917,N_213,N_2136);
nor U2918 (N_2918,N_1972,N_2306);
nand U2919 (N_2919,N_2433,N_1734);
nor U2920 (N_2920,N_598,N_1003);
or U2921 (N_2921,N_178,N_217);
and U2922 (N_2922,N_1002,N_2487);
nand U2923 (N_2923,N_895,N_1166);
xnor U2924 (N_2924,N_2279,N_351);
and U2925 (N_2925,N_34,N_1348);
nand U2926 (N_2926,N_1363,N_1910);
and U2927 (N_2927,N_279,N_1735);
nand U2928 (N_2928,N_2099,N_313);
xor U2929 (N_2929,N_1371,N_2243);
nand U2930 (N_2930,N_1723,N_390);
nand U2931 (N_2931,N_1687,N_790);
and U2932 (N_2932,N_750,N_1638);
and U2933 (N_2933,N_1359,N_1320);
nand U2934 (N_2934,N_940,N_1751);
and U2935 (N_2935,N_1559,N_1934);
nor U2936 (N_2936,N_108,N_454);
or U2937 (N_2937,N_1498,N_1787);
or U2938 (N_2938,N_1630,N_2093);
nand U2939 (N_2939,N_1012,N_823);
or U2940 (N_2940,N_1265,N_1599);
or U2941 (N_2941,N_2101,N_2150);
or U2942 (N_2942,N_142,N_803);
xnor U2943 (N_2943,N_2366,N_2208);
xor U2944 (N_2944,N_931,N_1546);
or U2945 (N_2945,N_1860,N_753);
nand U2946 (N_2946,N_437,N_292);
nand U2947 (N_2947,N_462,N_685);
or U2948 (N_2948,N_1301,N_1848);
xnor U2949 (N_2949,N_1110,N_1869);
or U2950 (N_2950,N_326,N_1072);
nor U2951 (N_2951,N_1150,N_1368);
or U2952 (N_2952,N_240,N_2089);
or U2953 (N_2953,N_2088,N_1794);
and U2954 (N_2954,N_2048,N_1516);
and U2955 (N_2955,N_673,N_451);
nand U2956 (N_2956,N_815,N_241);
xnor U2957 (N_2957,N_674,N_1533);
or U2958 (N_2958,N_764,N_2248);
nor U2959 (N_2959,N_2289,N_1605);
nor U2960 (N_2960,N_1420,N_679);
nand U2961 (N_2961,N_2056,N_497);
nand U2962 (N_2962,N_294,N_1976);
xnor U2963 (N_2963,N_780,N_590);
nor U2964 (N_2964,N_2438,N_485);
or U2965 (N_2965,N_2032,N_2027);
and U2966 (N_2966,N_1773,N_531);
nand U2967 (N_2967,N_1213,N_1275);
nor U2968 (N_2968,N_1828,N_124);
or U2969 (N_2969,N_368,N_1816);
or U2970 (N_2970,N_127,N_530);
xnor U2971 (N_2971,N_1386,N_1731);
and U2972 (N_2972,N_2464,N_334);
nand U2973 (N_2973,N_1929,N_2319);
xor U2974 (N_2974,N_1557,N_340);
nand U2975 (N_2975,N_2374,N_832);
nand U2976 (N_2976,N_477,N_2353);
nor U2977 (N_2977,N_797,N_1369);
nand U2978 (N_2978,N_2315,N_220);
or U2979 (N_2979,N_489,N_2297);
and U2980 (N_2980,N_1180,N_312);
or U2981 (N_2981,N_29,N_813);
or U2982 (N_2982,N_1228,N_798);
nand U2983 (N_2983,N_232,N_1887);
nand U2984 (N_2984,N_495,N_689);
or U2985 (N_2985,N_233,N_455);
nand U2986 (N_2986,N_1113,N_377);
nand U2987 (N_2987,N_2217,N_1087);
nor U2988 (N_2988,N_2402,N_365);
or U2989 (N_2989,N_1062,N_1246);
and U2990 (N_2990,N_369,N_1329);
xor U2991 (N_2991,N_2465,N_1237);
or U2992 (N_2992,N_834,N_7);
nor U2993 (N_2993,N_1827,N_440);
nand U2994 (N_2994,N_700,N_1021);
and U2995 (N_2995,N_919,N_658);
nand U2996 (N_2996,N_421,N_96);
or U2997 (N_2997,N_1897,N_331);
or U2998 (N_2998,N_696,N_1525);
or U2999 (N_2999,N_2213,N_1804);
and U3000 (N_3000,N_2364,N_2454);
or U3001 (N_3001,N_2123,N_1861);
nand U3002 (N_3002,N_1184,N_206);
nor U3003 (N_3003,N_2400,N_879);
nor U3004 (N_3004,N_1975,N_2407);
and U3005 (N_3005,N_1366,N_908);
or U3006 (N_3006,N_1311,N_419);
and U3007 (N_3007,N_1883,N_1777);
or U3008 (N_3008,N_2223,N_640);
or U3009 (N_3009,N_1137,N_187);
nor U3010 (N_3010,N_2496,N_1322);
xor U3011 (N_3011,N_1045,N_1919);
and U3012 (N_3012,N_647,N_1709);
or U3013 (N_3013,N_380,N_2112);
nand U3014 (N_3014,N_2202,N_1494);
or U3015 (N_3015,N_1662,N_1127);
nor U3016 (N_3016,N_911,N_2030);
or U3017 (N_3017,N_1680,N_2071);
nor U3018 (N_3018,N_2212,N_1146);
nor U3019 (N_3019,N_1537,N_189);
nor U3020 (N_3020,N_308,N_1841);
xor U3021 (N_3021,N_2342,N_2378);
nand U3022 (N_3022,N_2470,N_603);
nor U3023 (N_3023,N_2309,N_937);
xnor U3024 (N_3024,N_1983,N_1010);
nor U3025 (N_3025,N_564,N_247);
or U3026 (N_3026,N_1651,N_805);
xnor U3027 (N_3027,N_286,N_2332);
nor U3028 (N_3028,N_2390,N_2318);
and U3029 (N_3029,N_2127,N_1429);
nand U3030 (N_3030,N_214,N_848);
nand U3031 (N_3031,N_395,N_1837);
nor U3032 (N_3032,N_761,N_1249);
nand U3033 (N_3033,N_1252,N_655);
and U3034 (N_3034,N_2178,N_730);
nand U3035 (N_3035,N_155,N_1038);
nor U3036 (N_3036,N_708,N_1310);
and U3037 (N_3037,N_141,N_563);
nand U3038 (N_3038,N_2458,N_1046);
nor U3039 (N_3039,N_293,N_53);
nand U3040 (N_3040,N_429,N_1343);
nor U3041 (N_3041,N_303,N_1362);
nand U3042 (N_3042,N_686,N_1352);
nor U3043 (N_3043,N_1245,N_1400);
or U3044 (N_3044,N_1741,N_844);
nand U3045 (N_3045,N_1628,N_257);
nor U3046 (N_3046,N_271,N_1039);
nor U3047 (N_3047,N_1152,N_1905);
xor U3048 (N_3048,N_1871,N_366);
or U3049 (N_3049,N_1048,N_2239);
and U3050 (N_3050,N_733,N_106);
nand U3051 (N_3051,N_1446,N_649);
nor U3052 (N_3052,N_1197,N_596);
and U3053 (N_3053,N_1100,N_1951);
and U3054 (N_3054,N_1115,N_650);
or U3055 (N_3055,N_636,N_1430);
nand U3056 (N_3056,N_2126,N_1994);
or U3057 (N_3057,N_831,N_2468);
nand U3058 (N_3058,N_1780,N_1551);
nand U3059 (N_3059,N_502,N_2214);
or U3060 (N_3060,N_310,N_90);
nand U3061 (N_3061,N_960,N_819);
nand U3062 (N_3062,N_1210,N_782);
nand U3063 (N_3063,N_148,N_509);
or U3064 (N_3064,N_829,N_1341);
nor U3065 (N_3065,N_837,N_1222);
or U3066 (N_3066,N_2385,N_2200);
and U3067 (N_3067,N_1545,N_1840);
nand U3068 (N_3068,N_645,N_1700);
and U3069 (N_3069,N_54,N_595);
and U3070 (N_3070,N_210,N_84);
and U3071 (N_3071,N_2393,N_1271);
nand U3072 (N_3072,N_1891,N_4);
and U3073 (N_3073,N_1304,N_1527);
and U3074 (N_3074,N_1258,N_503);
xor U3075 (N_3075,N_2431,N_1539);
and U3076 (N_3076,N_2254,N_1066);
xor U3077 (N_3077,N_386,N_913);
xnor U3078 (N_3078,N_2311,N_732);
or U3079 (N_3079,N_529,N_2090);
and U3080 (N_3080,N_2105,N_107);
or U3081 (N_3081,N_1681,N_1879);
or U3082 (N_3082,N_117,N_1300);
and U3083 (N_3083,N_548,N_348);
xnor U3084 (N_3084,N_1558,N_2025);
or U3085 (N_3085,N_969,N_383);
nand U3086 (N_3086,N_2215,N_2142);
nor U3087 (N_3087,N_1358,N_1335);
and U3088 (N_3088,N_816,N_216);
xnor U3089 (N_3089,N_2394,N_443);
nand U3090 (N_3090,N_2175,N_98);
xor U3091 (N_3091,N_1874,N_2066);
or U3092 (N_3092,N_1308,N_1050);
and U3093 (N_3093,N_2004,N_1893);
nand U3094 (N_3094,N_1515,N_2280);
xnor U3095 (N_3095,N_1529,N_1888);
or U3096 (N_3096,N_1298,N_184);
nand U3097 (N_3097,N_715,N_1552);
and U3098 (N_3098,N_1782,N_2347);
nor U3099 (N_3099,N_1617,N_414);
or U3100 (N_3100,N_698,N_586);
and U3101 (N_3101,N_839,N_381);
xnor U3102 (N_3102,N_992,N_1355);
nand U3103 (N_3103,N_254,N_356);
or U3104 (N_3104,N_955,N_2333);
nor U3105 (N_3105,N_1034,N_55);
and U3106 (N_3106,N_1758,N_48);
and U3107 (N_3107,N_439,N_1991);
xnor U3108 (N_3108,N_2284,N_1522);
nor U3109 (N_3109,N_734,N_2049);
nand U3110 (N_3110,N_362,N_2492);
or U3111 (N_3111,N_2145,N_47);
nor U3112 (N_3112,N_1373,N_499);
nand U3113 (N_3113,N_161,N_357);
nand U3114 (N_3114,N_2370,N_2177);
and U3115 (N_3115,N_2100,N_1080);
nor U3116 (N_3116,N_147,N_2372);
nor U3117 (N_3117,N_327,N_559);
xor U3118 (N_3118,N_1277,N_151);
nor U3119 (N_3119,N_2341,N_64);
or U3120 (N_3120,N_1611,N_947);
nand U3121 (N_3121,N_1747,N_1044);
nand U3122 (N_3122,N_1854,N_997);
and U3123 (N_3123,N_2029,N_1164);
and U3124 (N_3124,N_920,N_1765);
nand U3125 (N_3125,N_1061,N_1195);
or U3126 (N_3126,N_628,N_470);
nand U3127 (N_3127,N_1969,N_1982);
and U3128 (N_3128,N_1568,N_450);
or U3129 (N_3129,N_1221,N_2255);
or U3130 (N_3130,N_1944,N_1410);
nand U3131 (N_3131,N_2074,N_154);
or U3132 (N_3132,N_1981,N_1163);
or U3133 (N_3133,N_2368,N_1915);
nand U3134 (N_3134,N_2225,N_1691);
or U3135 (N_3135,N_508,N_2131);
nand U3136 (N_3136,N_1333,N_1448);
nor U3137 (N_3137,N_2472,N_2107);
nor U3138 (N_3138,N_2422,N_1960);
or U3139 (N_3139,N_1582,N_31);
or U3140 (N_3140,N_606,N_1388);
xnor U3141 (N_3141,N_1281,N_128);
xnor U3142 (N_3142,N_1885,N_885);
nand U3143 (N_3143,N_1914,N_2361);
nand U3144 (N_3144,N_423,N_322);
or U3145 (N_3145,N_329,N_1548);
or U3146 (N_3146,N_2380,N_881);
and U3147 (N_3147,N_1015,N_1331);
and U3148 (N_3148,N_1279,N_290);
or U3149 (N_3149,N_1218,N_2209);
nand U3150 (N_3150,N_2017,N_2211);
and U3151 (N_3151,N_118,N_1449);
nand U3152 (N_3152,N_173,N_1345);
nand U3153 (N_3153,N_2419,N_269);
and U3154 (N_3154,N_1826,N_1154);
nor U3155 (N_3155,N_88,N_751);
and U3156 (N_3156,N_2387,N_619);
nand U3157 (N_3157,N_578,N_735);
nor U3158 (N_3158,N_1011,N_2263);
and U3159 (N_3159,N_901,N_371);
nand U3160 (N_3160,N_1350,N_1462);
or U3161 (N_3161,N_995,N_2146);
xnor U3162 (N_3162,N_459,N_1626);
or U3163 (N_3163,N_1158,N_433);
nor U3164 (N_3164,N_610,N_50);
or U3165 (N_3165,N_1239,N_393);
nor U3166 (N_3166,N_1196,N_1126);
or U3167 (N_3167,N_1306,N_149);
nand U3168 (N_3168,N_1695,N_1583);
and U3169 (N_3169,N_1666,N_1435);
nor U3170 (N_3170,N_460,N_339);
and U3171 (N_3171,N_1683,N_1005);
or U3172 (N_3172,N_122,N_2160);
nor U3173 (N_3173,N_1667,N_1917);
nand U3174 (N_3174,N_627,N_2163);
or U3175 (N_3175,N_1159,N_1968);
nor U3176 (N_3176,N_1678,N_961);
nor U3177 (N_3177,N_1855,N_1646);
and U3178 (N_3178,N_1190,N_987);
and U3179 (N_3179,N_1028,N_539);
nand U3180 (N_3180,N_315,N_1471);
or U3181 (N_3181,N_662,N_630);
nand U3182 (N_3182,N_62,N_1930);
and U3183 (N_3183,N_2272,N_1512);
and U3184 (N_3184,N_2489,N_971);
nand U3185 (N_3185,N_483,N_175);
or U3186 (N_3186,N_1941,N_2348);
or U3187 (N_3187,N_1886,N_1295);
and U3188 (N_3188,N_131,N_1230);
xnor U3189 (N_3189,N_2115,N_2148);
nand U3190 (N_3190,N_1440,N_1467);
nor U3191 (N_3191,N_2343,N_1182);
xnor U3192 (N_3192,N_472,N_778);
or U3193 (N_3193,N_545,N_1649);
and U3194 (N_3194,N_1468,N_2072);
or U3195 (N_3195,N_849,N_1104);
nor U3196 (N_3196,N_996,N_1942);
or U3197 (N_3197,N_2063,N_916);
and U3198 (N_3198,N_132,N_1058);
nand U3199 (N_3199,N_571,N_1697);
nand U3200 (N_3200,N_129,N_1719);
nand U3201 (N_3201,N_2455,N_140);
or U3202 (N_3202,N_867,N_237);
or U3203 (N_3203,N_401,N_697);
nor U3204 (N_3204,N_139,N_1670);
nor U3205 (N_3205,N_1083,N_14);
nand U3206 (N_3206,N_1784,N_1455);
and U3207 (N_3207,N_1242,N_926);
or U3208 (N_3208,N_249,N_710);
nand U3209 (N_3209,N_2218,N_1437);
and U3210 (N_3210,N_2052,N_1031);
or U3211 (N_3211,N_2137,N_1997);
and U3212 (N_3212,N_1097,N_2331);
and U3213 (N_3213,N_1798,N_409);
nand U3214 (N_3214,N_1901,N_1899);
or U3215 (N_3215,N_896,N_2);
nand U3216 (N_3216,N_212,N_260);
or U3217 (N_3217,N_776,N_163);
nor U3218 (N_3218,N_1572,N_726);
nor U3219 (N_3219,N_1227,N_1267);
xnor U3220 (N_3220,N_1434,N_1933);
or U3221 (N_3221,N_1935,N_2426);
nand U3222 (N_3222,N_1123,N_694);
or U3223 (N_3223,N_1148,N_1370);
nor U3224 (N_3224,N_426,N_2447);
nor U3225 (N_3225,N_1428,N_1401);
nand U3226 (N_3226,N_2375,N_374);
or U3227 (N_3227,N_1684,N_1685);
nand U3228 (N_3228,N_121,N_1894);
or U3229 (N_3229,N_1866,N_547);
xor U3230 (N_3230,N_250,N_552);
nor U3231 (N_3231,N_1738,N_442);
nand U3232 (N_3232,N_343,N_32);
or U3233 (N_3233,N_1303,N_1269);
or U3234 (N_3234,N_1851,N_1106);
nand U3235 (N_3235,N_1715,N_1830);
and U3236 (N_3236,N_884,N_33);
nor U3237 (N_3237,N_2104,N_592);
xnor U3238 (N_3238,N_2450,N_2403);
and U3239 (N_3239,N_296,N_2039);
and U3240 (N_3240,N_97,N_2308);
or U3241 (N_3241,N_134,N_1484);
nand U3242 (N_3242,N_2269,N_2018);
and U3243 (N_3243,N_1602,N_311);
or U3244 (N_3244,N_2143,N_1530);
and U3245 (N_3245,N_812,N_935);
nand U3246 (N_3246,N_456,N_259);
nand U3247 (N_3247,N_1,N_1390);
nand U3248 (N_3248,N_243,N_2373);
nand U3249 (N_3249,N_2204,N_988);
nor U3250 (N_3250,N_809,N_2242);
and U3251 (N_3251,N_1247,N_1105);
nor U3252 (N_3252,N_13,N_1740);
and U3253 (N_3253,N_2206,N_2210);
or U3254 (N_3254,N_397,N_72);
nand U3255 (N_3255,N_2418,N_2124);
xor U3256 (N_3256,N_1014,N_1803);
xnor U3257 (N_3257,N_1274,N_1262);
nor U3258 (N_3258,N_786,N_1328);
nor U3259 (N_3259,N_1705,N_648);
and U3260 (N_3260,N_2019,N_532);
or U3261 (N_3261,N_2021,N_158);
nor U3262 (N_3262,N_1339,N_985);
or U3263 (N_3263,N_435,N_56);
nand U3264 (N_3264,N_458,N_1616);
nand U3265 (N_3265,N_1278,N_2149);
nand U3266 (N_3266,N_1187,N_319);
and U3267 (N_3267,N_2328,N_1923);
and U3268 (N_3268,N_2367,N_2369);
nand U3269 (N_3269,N_2462,N_1973);
nand U3270 (N_3270,N_2005,N_2258);
nand U3271 (N_3271,N_977,N_504);
nor U3272 (N_3272,N_1198,N_870);
nor U3273 (N_3273,N_1577,N_2498);
nand U3274 (N_3274,N_309,N_1256);
nor U3275 (N_3275,N_847,N_1229);
nor U3276 (N_3276,N_962,N_1536);
or U3277 (N_3277,N_2451,N_204);
and U3278 (N_3278,N_2231,N_2246);
nor U3279 (N_3279,N_1018,N_2274);
or U3280 (N_3280,N_2300,N_2119);
nor U3281 (N_3281,N_1387,N_482);
nand U3282 (N_3282,N_981,N_1812);
nand U3283 (N_3283,N_1565,N_1095);
or U3284 (N_3284,N_1938,N_2303);
nand U3285 (N_3285,N_785,N_994);
or U3286 (N_3286,N_2266,N_1665);
nor U3287 (N_3287,N_60,N_1959);
nand U3288 (N_3288,N_43,N_1503);
or U3289 (N_3289,N_1903,N_754);
nor U3290 (N_3290,N_1389,N_1724);
xnor U3291 (N_3291,N_172,N_1464);
or U3292 (N_3292,N_1996,N_864);
nor U3293 (N_3293,N_1409,N_324);
or U3294 (N_3294,N_993,N_1550);
and U3295 (N_3295,N_1402,N_1261);
nor U3296 (N_3296,N_1850,N_2497);
or U3297 (N_3297,N_1349,N_1481);
and U3298 (N_3298,N_1199,N_755);
and U3299 (N_3299,N_1334,N_2144);
nor U3300 (N_3300,N_2070,N_1801);
nand U3301 (N_3301,N_641,N_1457);
nand U3302 (N_3302,N_1733,N_1346);
nand U3303 (N_3303,N_615,N_387);
nor U3304 (N_3304,N_2441,N_1624);
xnor U3305 (N_3305,N_1948,N_1762);
nand U3306 (N_3306,N_2409,N_683);
nand U3307 (N_3307,N_1055,N_2026);
nor U3308 (N_3308,N_771,N_1293);
and U3309 (N_3309,N_1771,N_1193);
nand U3310 (N_3310,N_413,N_345);
nor U3311 (N_3311,N_2228,N_1501);
xor U3312 (N_3312,N_1613,N_2196);
xor U3313 (N_3313,N_769,N_1574);
and U3314 (N_3314,N_80,N_2485);
nor U3315 (N_3315,N_886,N_1807);
nand U3316 (N_3316,N_1523,N_1768);
or U3317 (N_3317,N_990,N_1677);
nor U3318 (N_3318,N_278,N_945);
or U3319 (N_3319,N_1425,N_1327);
or U3320 (N_3320,N_1756,N_1353);
or U3321 (N_3321,N_681,N_740);
and U3322 (N_3322,N_17,N_1958);
and U3323 (N_3323,N_1737,N_1318);
xor U3324 (N_3324,N_157,N_915);
or U3325 (N_3325,N_2129,N_1019);
or U3326 (N_3326,N_1631,N_1965);
nor U3327 (N_3327,N_1241,N_1375);
nand U3328 (N_3328,N_1746,N_2028);
and U3329 (N_3329,N_1564,N_512);
or U3330 (N_3330,N_2033,N_2036);
and U3331 (N_3331,N_1987,N_2436);
and U3332 (N_3332,N_2499,N_245);
nand U3333 (N_3333,N_2007,N_665);
and U3334 (N_3334,N_1136,N_1081);
and U3335 (N_3335,N_1882,N_2132);
or U3336 (N_3336,N_1212,N_2421);
and U3337 (N_3337,N_1405,N_268);
or U3338 (N_3338,N_1819,N_2249);
or U3339 (N_3339,N_1226,N_1834);
or U3340 (N_3340,N_594,N_2408);
or U3341 (N_3341,N_479,N_866);
or U3342 (N_3342,N_1423,N_2410);
or U3343 (N_3343,N_253,N_2335);
nor U3344 (N_3344,N_2164,N_2432);
xnor U3345 (N_3345,N_1936,N_167);
nand U3346 (N_3346,N_2344,N_1473);
and U3347 (N_3347,N_589,N_519);
nor U3348 (N_3348,N_2134,N_2065);
or U3349 (N_3349,N_1089,N_2323);
nand U3350 (N_3350,N_1313,N_958);
nor U3351 (N_3351,N_1822,N_1299);
and U3352 (N_3352,N_1033,N_1635);
nor U3353 (N_3353,N_2086,N_226);
nand U3354 (N_3354,N_2141,N_1453);
nor U3355 (N_3355,N_89,N_61);
nand U3356 (N_3356,N_1703,N_1513);
and U3357 (N_3357,N_420,N_1118);
nor U3358 (N_3358,N_1070,N_558);
and U3359 (N_3359,N_136,N_86);
or U3360 (N_3360,N_1820,N_2201);
nor U3361 (N_3361,N_713,N_1181);
or U3362 (N_3362,N_2486,N_868);
or U3363 (N_3363,N_335,N_1475);
nor U3364 (N_3364,N_1049,N_289);
nand U3365 (N_3365,N_2345,N_1361);
nand U3366 (N_3366,N_1585,N_150);
nand U3367 (N_3367,N_973,N_192);
and U3368 (N_3368,N_731,N_2449);
or U3369 (N_3369,N_626,N_367);
and U3370 (N_3370,N_924,N_476);
nor U3371 (N_3371,N_1876,N_126);
nor U3372 (N_3372,N_239,N_1216);
nand U3373 (N_3373,N_566,N_1103);
xor U3374 (N_3374,N_27,N_1129);
nand U3375 (N_3375,N_2094,N_2417);
or U3376 (N_3376,N_2045,N_873);
nand U3377 (N_3377,N_1517,N_1658);
and U3378 (N_3378,N_446,N_1774);
and U3379 (N_3379,N_1082,N_1458);
nand U3380 (N_3380,N_73,N_38);
and U3381 (N_3381,N_288,N_2157);
nand U3382 (N_3382,N_424,N_2135);
or U3383 (N_3383,N_2195,N_1722);
xor U3384 (N_3384,N_2188,N_372);
or U3385 (N_3385,N_1176,N_828);
nand U3386 (N_3386,N_1486,N_1924);
or U3387 (N_3387,N_2110,N_468);
nor U3388 (N_3388,N_538,N_928);
or U3389 (N_3389,N_1167,N_1286);
nor U3390 (N_3390,N_1452,N_1007);
or U3391 (N_3391,N_274,N_1524);
nor U3392 (N_3392,N_501,N_2491);
and U3393 (N_3393,N_1799,N_1989);
nand U3394 (N_3394,N_1188,N_541);
and U3395 (N_3395,N_1612,N_2014);
nor U3396 (N_3396,N_1912,N_967);
nor U3397 (N_3397,N_1191,N_1634);
and U3398 (N_3398,N_2102,N_1984);
nor U3399 (N_3399,N_1569,N_1791);
and U3400 (N_3400,N_74,N_1493);
or U3401 (N_3401,N_1580,N_488);
nand U3402 (N_3402,N_1365,N_138);
and U3403 (N_3403,N_1650,N_1928);
nand U3404 (N_3404,N_929,N_1204);
or U3405 (N_3405,N_411,N_1287);
xnor U3406 (N_3406,N_1570,N_918);
or U3407 (N_3407,N_853,N_1629);
nor U3408 (N_3408,N_863,N_2040);
and U3409 (N_3409,N_851,N_487);
nand U3410 (N_3410,N_1391,N_701);
xnor U3411 (N_3411,N_1179,N_2191);
nor U3412 (N_3412,N_1307,N_1253);
and U3413 (N_3413,N_2114,N_2155);
or U3414 (N_3414,N_2304,N_199);
nor U3415 (N_3415,N_471,N_2006);
xnor U3416 (N_3416,N_2395,N_146);
nand U3417 (N_3417,N_1250,N_1032);
nor U3418 (N_3418,N_560,N_235);
nor U3419 (N_3419,N_1057,N_1117);
nor U3420 (N_3420,N_2130,N_1648);
nor U3421 (N_3421,N_2439,N_224);
xnor U3422 (N_3422,N_1273,N_1063);
and U3423 (N_3423,N_417,N_441);
and U3424 (N_3424,N_1971,N_1316);
and U3425 (N_3425,N_1625,N_744);
and U3426 (N_3426,N_511,N_9);
nor U3427 (N_3427,N_1022,N_143);
nand U3428 (N_3428,N_1478,N_70);
nand U3429 (N_3429,N_234,N_966);
or U3430 (N_3430,N_2235,N_384);
xnor U3431 (N_3431,N_922,N_917);
and U3432 (N_3432,N_516,N_1519);
nor U3433 (N_3433,N_842,N_169);
and U3434 (N_3434,N_1290,N_2466);
nor U3435 (N_3435,N_2187,N_1679);
nand U3436 (N_3436,N_909,N_561);
nor U3437 (N_3437,N_1337,N_1907);
nand U3438 (N_3438,N_2076,N_196);
nor U3439 (N_3439,N_203,N_114);
nand U3440 (N_3440,N_1474,N_215);
or U3441 (N_3441,N_1778,N_266);
nand U3442 (N_3442,N_1770,N_352);
xnor U3443 (N_3443,N_514,N_1009);
nand U3444 (N_3444,N_728,N_1203);
xnor U3445 (N_3445,N_2111,N_392);
or U3446 (N_3446,N_777,N_613);
nand U3447 (N_3447,N_2383,N_1925);
nor U3448 (N_3448,N_166,N_1563);
nand U3449 (N_3449,N_1757,N_469);
or U3450 (N_3450,N_2282,N_889);
or U3451 (N_3451,N_1094,N_1865);
nand U3452 (N_3452,N_1532,N_1424);
and U3453 (N_3453,N_1986,N_1051);
nor U3454 (N_3454,N_507,N_1920);
nand U3455 (N_3455,N_2185,N_2190);
or U3456 (N_3456,N_739,N_1766);
or U3457 (N_3457,N_1121,N_1326);
and U3458 (N_3458,N_418,N_1823);
and U3459 (N_3459,N_183,N_963);
and U3460 (N_3460,N_2042,N_1640);
and U3461 (N_3461,N_2412,N_2229);
nand U3462 (N_3462,N_407,N_1896);
or U3463 (N_3463,N_1321,N_1168);
nand U3464 (N_3464,N_1597,N_162);
nor U3465 (N_3465,N_608,N_727);
nand U3466 (N_3466,N_385,N_1953);
nor U3467 (N_3467,N_2002,N_856);
xor U3468 (N_3468,N_1174,N_874);
nand U3469 (N_3469,N_1134,N_197);
xnor U3470 (N_3470,N_1916,N_1482);
nand U3471 (N_3471,N_1540,N_580);
xnor U3472 (N_3472,N_284,N_1805);
nor U3473 (N_3473,N_826,N_272);
or U3474 (N_3474,N_1454,N_2326);
nand U3475 (N_3475,N_801,N_44);
nor U3476 (N_3476,N_1711,N_1020);
nor U3477 (N_3477,N_1690,N_1219);
and U3478 (N_3478,N_1591,N_1990);
nand U3479 (N_3479,N_513,N_473);
or U3480 (N_3480,N_1169,N_892);
nand U3481 (N_3481,N_1818,N_1347);
nand U3482 (N_3482,N_57,N_535);
nor U3483 (N_3483,N_1940,N_276);
or U3484 (N_3484,N_1065,N_614);
xor U3485 (N_3485,N_1421,N_716);
or U3486 (N_3486,N_2035,N_500);
nor U3487 (N_3487,N_1432,N_932);
nor U3488 (N_3488,N_1647,N_653);
and U3489 (N_3489,N_332,N_1560);
and U3490 (N_3490,N_1621,N_2302);
nor U3491 (N_3491,N_759,N_705);
nor U3492 (N_3492,N_796,N_116);
nor U3493 (N_3493,N_1090,N_2490);
and U3494 (N_3494,N_1450,N_1497);
or U3495 (N_3495,N_1714,N_1185);
or U3496 (N_3496,N_576,N_789);
nor U3497 (N_3497,N_170,N_1954);
nor U3498 (N_3498,N_855,N_2193);
nor U3499 (N_3499,N_1077,N_741);
nor U3500 (N_3500,N_1817,N_1500);
or U3501 (N_3501,N_2278,N_1674);
xnor U3502 (N_3502,N_1561,N_818);
nand U3503 (N_3503,N_283,N_965);
nand U3504 (N_3504,N_305,N_1330);
and U3505 (N_3505,N_1211,N_2117);
xor U3506 (N_3506,N_830,N_1451);
or U3507 (N_3507,N_2179,N_1422);
xor U3508 (N_3508,N_1783,N_1340);
nand U3509 (N_3509,N_37,N_1673);
nand U3510 (N_3510,N_1775,N_690);
and U3511 (N_3511,N_1949,N_1554);
and U3512 (N_3512,N_1403,N_200);
nand U3513 (N_3513,N_2363,N_897);
nand U3514 (N_3514,N_5,N_207);
nor U3515 (N_3515,N_857,N_2068);
nand U3516 (N_3516,N_262,N_1739);
nor U3517 (N_3517,N_153,N_1029);
nand U3518 (N_3518,N_902,N_1657);
nand U3519 (N_3519,N_1521,N_1476);
or U3520 (N_3520,N_1272,N_218);
nand U3521 (N_3521,N_1531,N_752);
nor U3522 (N_3522,N_341,N_1354);
xor U3523 (N_3523,N_526,N_1881);
or U3524 (N_3524,N_2222,N_63);
nor U3525 (N_3525,N_156,N_1729);
or U3526 (N_3526,N_15,N_2442);
and U3527 (N_3527,N_1511,N_1151);
and U3528 (N_3528,N_1382,N_394);
nor U3529 (N_3529,N_888,N_638);
or U3530 (N_3530,N_1220,N_79);
and U3531 (N_3531,N_298,N_2176);
or U3532 (N_3532,N_1567,N_1178);
nand U3533 (N_3533,N_2271,N_314);
nand U3534 (N_3534,N_275,N_1908);
and U3535 (N_3535,N_256,N_0);
or U3536 (N_3536,N_719,N_2346);
nand U3537 (N_3537,N_2008,N_1244);
or U3538 (N_3538,N_81,N_1264);
and U3539 (N_3539,N_1325,N_1900);
nand U3540 (N_3540,N_687,N_573);
or U3541 (N_3541,N_1317,N_2073);
nor U3542 (N_3542,N_1726,N_318);
and U3543 (N_3543,N_1124,N_781);
or U3544 (N_3544,N_1305,N_562);
nand U3545 (N_3545,N_549,N_1442);
nand U3546 (N_3546,N_496,N_2495);
or U3547 (N_3547,N_2207,N_1985);
or U3548 (N_3548,N_2260,N_1845);
or U3549 (N_3549,N_1172,N_432);
nor U3550 (N_3550,N_1217,N_12);
and U3551 (N_3551,N_2000,N_1596);
and U3552 (N_3552,N_1918,N_2082);
and U3553 (N_3553,N_194,N_2081);
nand U3554 (N_3554,N_428,N_875);
and U3555 (N_3555,N_570,N_346);
or U3556 (N_3556,N_599,N_684);
nand U3557 (N_3557,N_2299,N_2440);
and U3558 (N_3558,N_1542,N_2192);
and U3559 (N_3559,N_811,N_633);
and U3560 (N_3560,N_707,N_1632);
xor U3561 (N_3561,N_575,N_1752);
nor U3562 (N_3562,N_1713,N_6);
xnor U3563 (N_3563,N_135,N_1555);
and U3564 (N_3564,N_1642,N_2233);
or U3565 (N_3565,N_1831,N_1815);
and U3566 (N_3566,N_130,N_1809);
nor U3567 (N_3567,N_1074,N_970);
nor U3568 (N_3568,N_748,N_2397);
xnor U3569 (N_3569,N_669,N_491);
or U3570 (N_3570,N_666,N_1966);
and U3571 (N_3571,N_75,N_445);
or U3572 (N_3572,N_800,N_1967);
or U3573 (N_3573,N_792,N_724);
or U3574 (N_3574,N_572,N_1367);
nor U3575 (N_3575,N_1506,N_2015);
nand U3576 (N_3576,N_2481,N_1102);
nand U3577 (N_3577,N_1202,N_119);
nand U3578 (N_3578,N_58,N_517);
nor U3579 (N_3579,N_297,N_2275);
or U3580 (N_3580,N_2168,N_2267);
nor U3581 (N_3581,N_890,N_285);
nand U3582 (N_3582,N_587,N_2479);
and U3583 (N_3583,N_542,N_1445);
nor U3584 (N_3584,N_910,N_808);
nand U3585 (N_3585,N_2156,N_112);
nor U3586 (N_3586,N_3,N_1098);
xor U3587 (N_3587,N_1509,N_2138);
or U3588 (N_3588,N_1120,N_704);
or U3589 (N_3589,N_1763,N_452);
nand U3590 (N_3590,N_670,N_1636);
or U3591 (N_3591,N_824,N_1806);
xor U3592 (N_3592,N_1266,N_1408);
and U3593 (N_3593,N_51,N_1459);
or U3594 (N_3594,N_1143,N_1013);
or U3595 (N_3595,N_273,N_1491);
or U3596 (N_3596,N_695,N_758);
nand U3597 (N_3597,N_1108,N_1863);
xor U3598 (N_3598,N_1754,N_635);
xnor U3599 (N_3599,N_1315,N_1356);
and U3600 (N_3600,N_2038,N_1236);
and U3601 (N_3601,N_1867,N_1528);
or U3602 (N_3602,N_2423,N_2340);
nor U3603 (N_3603,N_1157,N_611);
nand U3604 (N_3604,N_661,N_209);
nand U3605 (N_3605,N_1383,N_317);
nand U3606 (N_3606,N_434,N_1604);
or U3607 (N_3607,N_1761,N_2336);
or U3608 (N_3608,N_2296,N_1280);
nor U3609 (N_3609,N_642,N_1393);
nand U3610 (N_3610,N_1689,N_1543);
and U3611 (N_3611,N_887,N_1205);
or U3612 (N_3612,N_1870,N_1760);
nand U3613 (N_3613,N_1288,N_1556);
and U3614 (N_3614,N_912,N_2097);
nand U3615 (N_3615,N_1170,N_1802);
and U3616 (N_3616,N_1263,N_953);
nand U3617 (N_3617,N_999,N_1921);
nor U3618 (N_3618,N_968,N_2337);
xor U3619 (N_3619,N_1438,N_1696);
nor U3620 (N_3620,N_2355,N_1769);
nand U3621 (N_3621,N_1655,N_1708);
xor U3622 (N_3622,N_1116,N_1622);
nand U3623 (N_3623,N_1692,N_2186);
nand U3624 (N_3624,N_680,N_1414);
and U3625 (N_3625,N_448,N_498);
nand U3626 (N_3626,N_2057,N_65);
nand U3627 (N_3627,N_1023,N_682);
nor U3628 (N_3628,N_225,N_2413);
or U3629 (N_3629,N_1466,N_980);
or U3630 (N_3630,N_505,N_267);
or U3631 (N_3631,N_525,N_2151);
nor U3632 (N_3632,N_2016,N_2140);
and U3633 (N_3633,N_1759,N_984);
nor U3634 (N_3634,N_120,N_242);
or U3635 (N_3635,N_1974,N_2069);
nand U3636 (N_3636,N_1800,N_1772);
and U3637 (N_3637,N_1875,N_25);
xor U3638 (N_3638,N_791,N_943);
and U3639 (N_3639,N_1101,N_359);
nand U3640 (N_3640,N_959,N_211);
xnor U3641 (N_3641,N_1644,N_557);
or U3642 (N_3642,N_551,N_416);
nand U3643 (N_3643,N_2391,N_2108);
and U3644 (N_3644,N_1068,N_306);
and U3645 (N_3645,N_631,N_2321);
nand U3646 (N_3646,N_2170,N_2430);
and U3647 (N_3647,N_1904,N_2058);
nor U3648 (N_3648,N_1206,N_1342);
nor U3649 (N_3649,N_338,N_1234);
or U3650 (N_3650,N_952,N_137);
and U3651 (N_3651,N_2147,N_1720);
or U3652 (N_3652,N_1276,N_1927);
nand U3653 (N_3653,N_2199,N_2463);
nand U3654 (N_3654,N_976,N_1292);
nand U3655 (N_3655,N_391,N_388);
or U3656 (N_3656,N_299,N_975);
or U3657 (N_3657,N_1480,N_1142);
nand U3658 (N_3658,N_2362,N_1884);
and U3659 (N_3659,N_577,N_702);
nor U3660 (N_3660,N_989,N_1578);
or U3661 (N_3661,N_783,N_1417);
or U3662 (N_3662,N_2268,N_474);
nor U3663 (N_3663,N_1086,N_1374);
or U3664 (N_3664,N_1461,N_1748);
nand U3665 (N_3665,N_325,N_144);
nand U3666 (N_3666,N_1487,N_1469);
or U3667 (N_3667,N_2379,N_344);
nand U3668 (N_3668,N_1238,N_1259);
and U3669 (N_3669,N_87,N_1504);
and U3670 (N_3670,N_742,N_2365);
or U3671 (N_3671,N_515,N_1384);
nor U3672 (N_3672,N_431,N_2494);
or U3673 (N_3673,N_222,N_1412);
nor U3674 (N_3674,N_1314,N_581);
nand U3675 (N_3675,N_1447,N_1620);
or U3676 (N_3676,N_2241,N_449);
and U3677 (N_3677,N_2411,N_354);
and U3678 (N_3678,N_2237,N_229);
nand U3679 (N_3679,N_609,N_533);
or U3680 (N_3680,N_907,N_453);
nand U3681 (N_3681,N_76,N_1619);
or U3682 (N_3682,N_2080,N_747);
nor U3683 (N_3683,N_979,N_2121);
xnor U3684 (N_3684,N_1394,N_1016);
and U3685 (N_3685,N_2205,N_1042);
nor U3686 (N_3686,N_1378,N_425);
or U3687 (N_3687,N_2012,N_1979);
or U3688 (N_3688,N_644,N_1411);
and U3689 (N_3689,N_667,N_400);
nand U3690 (N_3690,N_825,N_100);
or U3691 (N_3691,N_180,N_280);
nor U3692 (N_3692,N_1792,N_872);
nand U3693 (N_3693,N_1829,N_113);
or U3694 (N_3694,N_2067,N_1251);
nor U3695 (N_3695,N_600,N_2382);
or U3696 (N_3696,N_77,N_195);
xnor U3697 (N_3697,N_2416,N_2293);
nor U3698 (N_3698,N_1133,N_1189);
and U3699 (N_3699,N_1357,N_492);
nand U3700 (N_3700,N_1957,N_1344);
or U3701 (N_3701,N_656,N_465);
nand U3702 (N_3702,N_986,N_717);
or U3703 (N_3703,N_1704,N_2446);
nand U3704 (N_3704,N_1351,N_2161);
xor U3705 (N_3705,N_1385,N_1659);
nor U3706 (N_3706,N_1937,N_604);
xor U3707 (N_3707,N_942,N_841);
and U3708 (N_3708,N_231,N_802);
nor U3709 (N_3709,N_375,N_109);
or U3710 (N_3710,N_998,N_1593);
nand U3711 (N_3711,N_905,N_1223);
nand U3712 (N_3712,N_1093,N_185);
and U3713 (N_3713,N_1544,N_930);
xnor U3714 (N_3714,N_1698,N_1939);
and U3715 (N_3715,N_725,N_1248);
xnor U3716 (N_3716,N_787,N_1743);
and U3717 (N_3717,N_19,N_2314);
and U3718 (N_3718,N_543,N_1549);
or U3719 (N_3719,N_1231,N_883);
xor U3720 (N_3720,N_101,N_2424);
nor U3721 (N_3721,N_2338,N_2273);
xnor U3722 (N_3722,N_1716,N_845);
nor U3723 (N_3723,N_1505,N_1898);
nand U3724 (N_3724,N_1153,N_1566);
and U3725 (N_3725,N_205,N_1284);
or U3726 (N_3726,N_676,N_1581);
or U3727 (N_3727,N_2167,N_956);
and U3728 (N_3728,N_1843,N_402);
or U3729 (N_3729,N_373,N_24);
nand U3730 (N_3730,N_1682,N_1878);
nor U3731 (N_3731,N_399,N_347);
xor U3732 (N_3732,N_688,N_2420);
nor U3733 (N_3733,N_623,N_376);
xor U3734 (N_3734,N_2064,N_1067);
or U3735 (N_3735,N_265,N_2139);
nand U3736 (N_3736,N_336,N_878);
nand U3737 (N_3737,N_1810,N_1514);
nand U3738 (N_3738,N_2406,N_1796);
or U3739 (N_3739,N_67,N_2376);
nor U3740 (N_3740,N_1302,N_1872);
nand U3741 (N_3741,N_1858,N_123);
nand U3742 (N_3742,N_1688,N_1499);
and U3743 (N_3743,N_164,N_893);
nand U3744 (N_3744,N_567,N_1821);
nand U3745 (N_3745,N_475,N_601);
or U3746 (N_3746,N_201,N_1669);
or U3747 (N_3747,N_422,N_1781);
xor U3748 (N_3748,N_2349,N_616);
or U3749 (N_3749,N_466,N_406);
nor U3750 (N_3750,N_2102,N_114);
nor U3751 (N_3751,N_1212,N_1221);
nor U3752 (N_3752,N_971,N_467);
nand U3753 (N_3753,N_1910,N_1588);
nand U3754 (N_3754,N_892,N_1789);
nand U3755 (N_3755,N_1483,N_289);
or U3756 (N_3756,N_2166,N_482);
nor U3757 (N_3757,N_2027,N_513);
nand U3758 (N_3758,N_734,N_786);
nand U3759 (N_3759,N_853,N_613);
or U3760 (N_3760,N_53,N_1216);
nor U3761 (N_3761,N_1681,N_2002);
and U3762 (N_3762,N_1401,N_2370);
and U3763 (N_3763,N_16,N_1478);
and U3764 (N_3764,N_1632,N_1711);
or U3765 (N_3765,N_2235,N_2131);
and U3766 (N_3766,N_973,N_2410);
nand U3767 (N_3767,N_421,N_173);
nand U3768 (N_3768,N_763,N_1615);
nand U3769 (N_3769,N_1062,N_764);
nor U3770 (N_3770,N_2067,N_1103);
and U3771 (N_3771,N_123,N_222);
nand U3772 (N_3772,N_271,N_1559);
nor U3773 (N_3773,N_839,N_361);
xnor U3774 (N_3774,N_686,N_2187);
or U3775 (N_3775,N_1532,N_1855);
nor U3776 (N_3776,N_2115,N_1946);
nor U3777 (N_3777,N_2232,N_1892);
and U3778 (N_3778,N_1989,N_1343);
or U3779 (N_3779,N_904,N_1964);
or U3780 (N_3780,N_2423,N_141);
and U3781 (N_3781,N_971,N_1111);
nand U3782 (N_3782,N_268,N_2087);
nand U3783 (N_3783,N_307,N_1223);
or U3784 (N_3784,N_1723,N_526);
nand U3785 (N_3785,N_1469,N_544);
and U3786 (N_3786,N_280,N_2196);
nand U3787 (N_3787,N_1961,N_1377);
nor U3788 (N_3788,N_1284,N_1712);
nand U3789 (N_3789,N_1313,N_2077);
nand U3790 (N_3790,N_2492,N_2257);
or U3791 (N_3791,N_2378,N_2050);
and U3792 (N_3792,N_2137,N_983);
and U3793 (N_3793,N_1637,N_1111);
nor U3794 (N_3794,N_2134,N_1454);
and U3795 (N_3795,N_1203,N_2010);
and U3796 (N_3796,N_1894,N_1273);
and U3797 (N_3797,N_2271,N_1135);
nand U3798 (N_3798,N_1103,N_266);
and U3799 (N_3799,N_1926,N_1181);
or U3800 (N_3800,N_576,N_2085);
nand U3801 (N_3801,N_764,N_884);
xor U3802 (N_3802,N_1000,N_1988);
and U3803 (N_3803,N_788,N_2111);
or U3804 (N_3804,N_1676,N_1925);
nor U3805 (N_3805,N_890,N_307);
nand U3806 (N_3806,N_332,N_1131);
nand U3807 (N_3807,N_584,N_2203);
and U3808 (N_3808,N_1293,N_788);
or U3809 (N_3809,N_1937,N_565);
or U3810 (N_3810,N_124,N_185);
nand U3811 (N_3811,N_560,N_970);
nor U3812 (N_3812,N_797,N_42);
xnor U3813 (N_3813,N_845,N_139);
or U3814 (N_3814,N_2486,N_1270);
nor U3815 (N_3815,N_2196,N_2342);
and U3816 (N_3816,N_643,N_1150);
and U3817 (N_3817,N_305,N_1946);
nor U3818 (N_3818,N_823,N_1625);
nor U3819 (N_3819,N_1117,N_1915);
or U3820 (N_3820,N_1677,N_858);
or U3821 (N_3821,N_1550,N_541);
nor U3822 (N_3822,N_2039,N_1718);
and U3823 (N_3823,N_489,N_530);
and U3824 (N_3824,N_546,N_2105);
xnor U3825 (N_3825,N_2407,N_1839);
nand U3826 (N_3826,N_80,N_789);
nor U3827 (N_3827,N_872,N_2201);
or U3828 (N_3828,N_1761,N_2299);
or U3829 (N_3829,N_1545,N_1029);
nor U3830 (N_3830,N_2147,N_2290);
xor U3831 (N_3831,N_1313,N_142);
nand U3832 (N_3832,N_109,N_1570);
nor U3833 (N_3833,N_2247,N_1731);
or U3834 (N_3834,N_2465,N_1447);
and U3835 (N_3835,N_2410,N_1447);
nor U3836 (N_3836,N_921,N_266);
nand U3837 (N_3837,N_1433,N_314);
and U3838 (N_3838,N_1516,N_361);
or U3839 (N_3839,N_1182,N_1447);
and U3840 (N_3840,N_2257,N_1039);
nor U3841 (N_3841,N_2154,N_2460);
xor U3842 (N_3842,N_1505,N_927);
and U3843 (N_3843,N_1557,N_1858);
nand U3844 (N_3844,N_1156,N_598);
nand U3845 (N_3845,N_1842,N_1278);
xor U3846 (N_3846,N_2374,N_1829);
nand U3847 (N_3847,N_1068,N_1004);
nand U3848 (N_3848,N_393,N_2029);
nand U3849 (N_3849,N_144,N_861);
and U3850 (N_3850,N_268,N_1023);
or U3851 (N_3851,N_2327,N_722);
and U3852 (N_3852,N_1626,N_1277);
nand U3853 (N_3853,N_879,N_1920);
nor U3854 (N_3854,N_1361,N_1889);
or U3855 (N_3855,N_1942,N_1472);
nor U3856 (N_3856,N_679,N_1624);
or U3857 (N_3857,N_1485,N_940);
or U3858 (N_3858,N_192,N_215);
or U3859 (N_3859,N_1185,N_669);
and U3860 (N_3860,N_2279,N_288);
and U3861 (N_3861,N_2106,N_781);
or U3862 (N_3862,N_1689,N_1615);
nor U3863 (N_3863,N_319,N_1150);
nor U3864 (N_3864,N_249,N_1592);
nor U3865 (N_3865,N_507,N_1110);
and U3866 (N_3866,N_998,N_206);
nor U3867 (N_3867,N_418,N_725);
xor U3868 (N_3868,N_1639,N_387);
nor U3869 (N_3869,N_578,N_954);
nand U3870 (N_3870,N_1928,N_1276);
nand U3871 (N_3871,N_427,N_1590);
nand U3872 (N_3872,N_866,N_233);
and U3873 (N_3873,N_1849,N_328);
nand U3874 (N_3874,N_1712,N_1896);
or U3875 (N_3875,N_1714,N_992);
xnor U3876 (N_3876,N_214,N_2082);
nand U3877 (N_3877,N_1494,N_1323);
nand U3878 (N_3878,N_621,N_1769);
or U3879 (N_3879,N_882,N_367);
nand U3880 (N_3880,N_588,N_1429);
or U3881 (N_3881,N_713,N_2054);
nand U3882 (N_3882,N_275,N_554);
and U3883 (N_3883,N_797,N_101);
or U3884 (N_3884,N_153,N_452);
nor U3885 (N_3885,N_2064,N_205);
nor U3886 (N_3886,N_2046,N_1808);
nor U3887 (N_3887,N_2155,N_2109);
and U3888 (N_3888,N_2096,N_32);
xnor U3889 (N_3889,N_1189,N_968);
nor U3890 (N_3890,N_18,N_411);
or U3891 (N_3891,N_274,N_1358);
nor U3892 (N_3892,N_2257,N_1357);
nor U3893 (N_3893,N_1036,N_1191);
nand U3894 (N_3894,N_1236,N_1655);
nor U3895 (N_3895,N_2220,N_1410);
or U3896 (N_3896,N_990,N_1144);
nor U3897 (N_3897,N_1911,N_1129);
nor U3898 (N_3898,N_63,N_273);
nand U3899 (N_3899,N_2158,N_915);
and U3900 (N_3900,N_1754,N_627);
nand U3901 (N_3901,N_785,N_1237);
nand U3902 (N_3902,N_822,N_991);
nand U3903 (N_3903,N_469,N_1889);
nor U3904 (N_3904,N_963,N_2493);
nand U3905 (N_3905,N_1091,N_1305);
nor U3906 (N_3906,N_1095,N_1133);
and U3907 (N_3907,N_764,N_1499);
nand U3908 (N_3908,N_2298,N_2126);
nor U3909 (N_3909,N_388,N_487);
nor U3910 (N_3910,N_225,N_2372);
and U3911 (N_3911,N_1052,N_370);
nand U3912 (N_3912,N_1715,N_2498);
nor U3913 (N_3913,N_1285,N_1284);
nor U3914 (N_3914,N_1233,N_432);
nand U3915 (N_3915,N_944,N_1154);
nor U3916 (N_3916,N_1710,N_1452);
nor U3917 (N_3917,N_656,N_297);
and U3918 (N_3918,N_1610,N_983);
nor U3919 (N_3919,N_449,N_711);
nor U3920 (N_3920,N_160,N_1167);
or U3921 (N_3921,N_1916,N_1066);
or U3922 (N_3922,N_964,N_1634);
xor U3923 (N_3923,N_900,N_549);
nor U3924 (N_3924,N_439,N_837);
and U3925 (N_3925,N_851,N_1397);
nor U3926 (N_3926,N_1086,N_754);
nor U3927 (N_3927,N_459,N_847);
nor U3928 (N_3928,N_199,N_1870);
or U3929 (N_3929,N_1002,N_1468);
xor U3930 (N_3930,N_730,N_462);
and U3931 (N_3931,N_1153,N_2107);
nor U3932 (N_3932,N_1213,N_1658);
xor U3933 (N_3933,N_1974,N_1123);
nand U3934 (N_3934,N_1237,N_1424);
and U3935 (N_3935,N_2491,N_898);
xnor U3936 (N_3936,N_2067,N_1512);
nor U3937 (N_3937,N_822,N_405);
and U3938 (N_3938,N_1953,N_1161);
xor U3939 (N_3939,N_1433,N_824);
nor U3940 (N_3940,N_1050,N_1355);
nor U3941 (N_3941,N_2242,N_1490);
nor U3942 (N_3942,N_32,N_176);
and U3943 (N_3943,N_1136,N_887);
nand U3944 (N_3944,N_265,N_1267);
or U3945 (N_3945,N_2147,N_2021);
and U3946 (N_3946,N_1763,N_2285);
nand U3947 (N_3947,N_1404,N_698);
nor U3948 (N_3948,N_2238,N_323);
nor U3949 (N_3949,N_382,N_498);
nand U3950 (N_3950,N_1066,N_589);
and U3951 (N_3951,N_1280,N_432);
nand U3952 (N_3952,N_191,N_261);
and U3953 (N_3953,N_1724,N_1067);
nor U3954 (N_3954,N_1547,N_2348);
nand U3955 (N_3955,N_1032,N_2402);
nor U3956 (N_3956,N_957,N_2364);
nor U3957 (N_3957,N_1007,N_1489);
nand U3958 (N_3958,N_2292,N_1207);
and U3959 (N_3959,N_1345,N_1005);
nand U3960 (N_3960,N_315,N_750);
or U3961 (N_3961,N_2138,N_747);
nor U3962 (N_3962,N_2170,N_89);
nand U3963 (N_3963,N_488,N_1651);
and U3964 (N_3964,N_2100,N_824);
and U3965 (N_3965,N_1723,N_1325);
nor U3966 (N_3966,N_494,N_1591);
xnor U3967 (N_3967,N_1442,N_2146);
and U3968 (N_3968,N_2212,N_596);
nand U3969 (N_3969,N_280,N_930);
and U3970 (N_3970,N_188,N_1455);
nor U3971 (N_3971,N_1120,N_1957);
or U3972 (N_3972,N_2122,N_1554);
xor U3973 (N_3973,N_289,N_2238);
nand U3974 (N_3974,N_946,N_227);
or U3975 (N_3975,N_1403,N_506);
and U3976 (N_3976,N_230,N_22);
or U3977 (N_3977,N_2384,N_561);
and U3978 (N_3978,N_1133,N_71);
nand U3979 (N_3979,N_427,N_1269);
or U3980 (N_3980,N_1288,N_1265);
or U3981 (N_3981,N_649,N_2065);
xor U3982 (N_3982,N_1516,N_2267);
nand U3983 (N_3983,N_906,N_713);
or U3984 (N_3984,N_1727,N_1923);
or U3985 (N_3985,N_1627,N_2288);
nand U3986 (N_3986,N_1303,N_1036);
nor U3987 (N_3987,N_851,N_1798);
nand U3988 (N_3988,N_801,N_1345);
and U3989 (N_3989,N_1676,N_1136);
nand U3990 (N_3990,N_1294,N_459);
nor U3991 (N_3991,N_2365,N_654);
or U3992 (N_3992,N_1620,N_1309);
or U3993 (N_3993,N_607,N_1915);
nor U3994 (N_3994,N_1284,N_584);
nor U3995 (N_3995,N_2204,N_1396);
nand U3996 (N_3996,N_958,N_2386);
nand U3997 (N_3997,N_1304,N_1674);
and U3998 (N_3998,N_2185,N_597);
xor U3999 (N_3999,N_1751,N_578);
nand U4000 (N_4000,N_1970,N_1499);
nor U4001 (N_4001,N_1042,N_2255);
or U4002 (N_4002,N_525,N_379);
nor U4003 (N_4003,N_1648,N_1977);
nor U4004 (N_4004,N_1152,N_509);
nor U4005 (N_4005,N_1260,N_1651);
nor U4006 (N_4006,N_2189,N_504);
nand U4007 (N_4007,N_258,N_197);
nand U4008 (N_4008,N_37,N_2085);
and U4009 (N_4009,N_1211,N_1282);
or U4010 (N_4010,N_1390,N_1819);
or U4011 (N_4011,N_2383,N_2036);
nor U4012 (N_4012,N_1678,N_1751);
nor U4013 (N_4013,N_1844,N_1748);
and U4014 (N_4014,N_56,N_355);
nand U4015 (N_4015,N_464,N_1389);
or U4016 (N_4016,N_560,N_815);
nor U4017 (N_4017,N_559,N_683);
nor U4018 (N_4018,N_2130,N_1660);
or U4019 (N_4019,N_2341,N_1625);
or U4020 (N_4020,N_1547,N_1832);
or U4021 (N_4021,N_1845,N_2303);
nand U4022 (N_4022,N_817,N_2398);
nand U4023 (N_4023,N_194,N_1238);
and U4024 (N_4024,N_1652,N_1453);
or U4025 (N_4025,N_2044,N_1908);
and U4026 (N_4026,N_873,N_665);
nand U4027 (N_4027,N_730,N_1995);
xor U4028 (N_4028,N_746,N_2191);
and U4029 (N_4029,N_1753,N_1104);
or U4030 (N_4030,N_517,N_2056);
and U4031 (N_4031,N_1453,N_1218);
nor U4032 (N_4032,N_603,N_1739);
and U4033 (N_4033,N_2311,N_1909);
nor U4034 (N_4034,N_165,N_2276);
and U4035 (N_4035,N_2228,N_1658);
and U4036 (N_4036,N_1687,N_1174);
xnor U4037 (N_4037,N_843,N_1619);
or U4038 (N_4038,N_958,N_1835);
or U4039 (N_4039,N_922,N_983);
nor U4040 (N_4040,N_22,N_854);
xnor U4041 (N_4041,N_1783,N_526);
and U4042 (N_4042,N_1977,N_1715);
nor U4043 (N_4043,N_1031,N_1266);
and U4044 (N_4044,N_2314,N_1803);
nor U4045 (N_4045,N_541,N_2000);
nand U4046 (N_4046,N_1423,N_730);
and U4047 (N_4047,N_486,N_710);
nand U4048 (N_4048,N_1216,N_2360);
and U4049 (N_4049,N_918,N_2474);
nand U4050 (N_4050,N_1744,N_517);
nor U4051 (N_4051,N_680,N_2230);
xnor U4052 (N_4052,N_1949,N_174);
nor U4053 (N_4053,N_326,N_2060);
nor U4054 (N_4054,N_76,N_1333);
nand U4055 (N_4055,N_2490,N_2019);
nand U4056 (N_4056,N_190,N_2158);
nand U4057 (N_4057,N_2022,N_944);
or U4058 (N_4058,N_1244,N_2494);
or U4059 (N_4059,N_2085,N_1573);
and U4060 (N_4060,N_94,N_2254);
nor U4061 (N_4061,N_926,N_793);
nor U4062 (N_4062,N_699,N_1889);
or U4063 (N_4063,N_377,N_1931);
nand U4064 (N_4064,N_293,N_345);
or U4065 (N_4065,N_1717,N_2302);
and U4066 (N_4066,N_599,N_1273);
nand U4067 (N_4067,N_798,N_2173);
xor U4068 (N_4068,N_1405,N_88);
nor U4069 (N_4069,N_161,N_1579);
nor U4070 (N_4070,N_1971,N_490);
and U4071 (N_4071,N_210,N_357);
nand U4072 (N_4072,N_2138,N_690);
xnor U4073 (N_4073,N_1194,N_404);
and U4074 (N_4074,N_1758,N_622);
or U4075 (N_4075,N_981,N_1182);
nor U4076 (N_4076,N_1652,N_2256);
or U4077 (N_4077,N_90,N_1742);
or U4078 (N_4078,N_1169,N_2171);
or U4079 (N_4079,N_2347,N_1772);
and U4080 (N_4080,N_2102,N_912);
nor U4081 (N_4081,N_624,N_2344);
or U4082 (N_4082,N_2254,N_2263);
nor U4083 (N_4083,N_712,N_1461);
or U4084 (N_4084,N_255,N_1240);
or U4085 (N_4085,N_66,N_1634);
nor U4086 (N_4086,N_950,N_1500);
and U4087 (N_4087,N_1226,N_826);
and U4088 (N_4088,N_1571,N_2458);
or U4089 (N_4089,N_2018,N_1901);
nand U4090 (N_4090,N_2085,N_810);
and U4091 (N_4091,N_1342,N_2256);
nor U4092 (N_4092,N_1028,N_917);
or U4093 (N_4093,N_1,N_905);
or U4094 (N_4094,N_1109,N_813);
and U4095 (N_4095,N_2206,N_1175);
and U4096 (N_4096,N_223,N_321);
or U4097 (N_4097,N_2462,N_1876);
nand U4098 (N_4098,N_1134,N_1466);
nor U4099 (N_4099,N_1621,N_2030);
xor U4100 (N_4100,N_1039,N_336);
or U4101 (N_4101,N_1035,N_2085);
or U4102 (N_4102,N_1978,N_41);
or U4103 (N_4103,N_2386,N_1861);
nor U4104 (N_4104,N_1011,N_75);
xor U4105 (N_4105,N_2135,N_1335);
and U4106 (N_4106,N_1540,N_1488);
xor U4107 (N_4107,N_1408,N_763);
nand U4108 (N_4108,N_1917,N_1205);
or U4109 (N_4109,N_352,N_2273);
nor U4110 (N_4110,N_298,N_2090);
nor U4111 (N_4111,N_1405,N_1920);
and U4112 (N_4112,N_566,N_1834);
nand U4113 (N_4113,N_1489,N_2205);
or U4114 (N_4114,N_1838,N_1861);
or U4115 (N_4115,N_74,N_1152);
nand U4116 (N_4116,N_1135,N_2427);
and U4117 (N_4117,N_15,N_2156);
nor U4118 (N_4118,N_154,N_621);
xor U4119 (N_4119,N_558,N_13);
or U4120 (N_4120,N_1598,N_2045);
xnor U4121 (N_4121,N_178,N_244);
and U4122 (N_4122,N_225,N_893);
nor U4123 (N_4123,N_43,N_436);
nor U4124 (N_4124,N_946,N_1058);
or U4125 (N_4125,N_1840,N_1142);
and U4126 (N_4126,N_514,N_1915);
nor U4127 (N_4127,N_405,N_105);
and U4128 (N_4128,N_2118,N_869);
and U4129 (N_4129,N_2286,N_2089);
nand U4130 (N_4130,N_2432,N_2090);
nor U4131 (N_4131,N_1718,N_214);
nor U4132 (N_4132,N_1099,N_608);
or U4133 (N_4133,N_2252,N_1622);
or U4134 (N_4134,N_1791,N_2141);
nor U4135 (N_4135,N_932,N_1983);
nor U4136 (N_4136,N_661,N_456);
or U4137 (N_4137,N_1375,N_202);
nor U4138 (N_4138,N_364,N_2484);
nand U4139 (N_4139,N_2111,N_2187);
or U4140 (N_4140,N_1797,N_892);
nor U4141 (N_4141,N_2125,N_1233);
nand U4142 (N_4142,N_919,N_514);
nor U4143 (N_4143,N_1611,N_1);
and U4144 (N_4144,N_1365,N_1463);
nand U4145 (N_4145,N_1022,N_628);
and U4146 (N_4146,N_2036,N_1609);
and U4147 (N_4147,N_2496,N_671);
nor U4148 (N_4148,N_280,N_281);
nand U4149 (N_4149,N_1392,N_1445);
and U4150 (N_4150,N_1100,N_32);
or U4151 (N_4151,N_649,N_412);
nand U4152 (N_4152,N_367,N_2003);
or U4153 (N_4153,N_1732,N_1373);
nor U4154 (N_4154,N_1409,N_883);
nor U4155 (N_4155,N_786,N_1635);
nor U4156 (N_4156,N_2193,N_1662);
nand U4157 (N_4157,N_2141,N_2269);
or U4158 (N_4158,N_1064,N_721);
and U4159 (N_4159,N_2038,N_1462);
and U4160 (N_4160,N_2286,N_72);
nand U4161 (N_4161,N_1845,N_167);
nand U4162 (N_4162,N_2098,N_8);
or U4163 (N_4163,N_376,N_1589);
and U4164 (N_4164,N_1361,N_707);
and U4165 (N_4165,N_1847,N_287);
or U4166 (N_4166,N_2323,N_2007);
or U4167 (N_4167,N_2056,N_1976);
nor U4168 (N_4168,N_604,N_2335);
nor U4169 (N_4169,N_2480,N_1108);
and U4170 (N_4170,N_734,N_383);
xnor U4171 (N_4171,N_840,N_2261);
xnor U4172 (N_4172,N_2071,N_1198);
or U4173 (N_4173,N_2466,N_1786);
xor U4174 (N_4174,N_1017,N_802);
and U4175 (N_4175,N_922,N_786);
nand U4176 (N_4176,N_1766,N_2443);
and U4177 (N_4177,N_380,N_25);
nor U4178 (N_4178,N_570,N_2008);
or U4179 (N_4179,N_542,N_1492);
nand U4180 (N_4180,N_62,N_2416);
nand U4181 (N_4181,N_483,N_471);
nor U4182 (N_4182,N_93,N_1218);
or U4183 (N_4183,N_1984,N_1302);
nand U4184 (N_4184,N_235,N_1542);
nand U4185 (N_4185,N_1435,N_1473);
nor U4186 (N_4186,N_1370,N_743);
and U4187 (N_4187,N_925,N_2361);
and U4188 (N_4188,N_710,N_1219);
and U4189 (N_4189,N_708,N_196);
or U4190 (N_4190,N_511,N_550);
or U4191 (N_4191,N_669,N_979);
nor U4192 (N_4192,N_2063,N_2206);
nor U4193 (N_4193,N_834,N_919);
xor U4194 (N_4194,N_950,N_388);
and U4195 (N_4195,N_970,N_278);
and U4196 (N_4196,N_741,N_2222);
nand U4197 (N_4197,N_668,N_1307);
xor U4198 (N_4198,N_1049,N_2443);
and U4199 (N_4199,N_2050,N_837);
nor U4200 (N_4200,N_1060,N_2162);
and U4201 (N_4201,N_1152,N_2011);
nand U4202 (N_4202,N_187,N_803);
nand U4203 (N_4203,N_96,N_316);
nor U4204 (N_4204,N_1372,N_1318);
and U4205 (N_4205,N_617,N_785);
xor U4206 (N_4206,N_2109,N_2185);
nor U4207 (N_4207,N_1675,N_161);
and U4208 (N_4208,N_1146,N_1738);
and U4209 (N_4209,N_2066,N_1758);
or U4210 (N_4210,N_58,N_2045);
or U4211 (N_4211,N_1117,N_865);
and U4212 (N_4212,N_1267,N_2132);
nand U4213 (N_4213,N_720,N_2147);
nand U4214 (N_4214,N_1199,N_2473);
nor U4215 (N_4215,N_877,N_891);
nand U4216 (N_4216,N_235,N_379);
or U4217 (N_4217,N_2048,N_1278);
nand U4218 (N_4218,N_1009,N_1572);
xor U4219 (N_4219,N_1144,N_569);
nand U4220 (N_4220,N_997,N_590);
nand U4221 (N_4221,N_2438,N_378);
nand U4222 (N_4222,N_2304,N_462);
and U4223 (N_4223,N_711,N_1491);
nor U4224 (N_4224,N_1877,N_1659);
xnor U4225 (N_4225,N_813,N_1595);
nand U4226 (N_4226,N_2043,N_646);
nand U4227 (N_4227,N_268,N_1850);
and U4228 (N_4228,N_1477,N_21);
nand U4229 (N_4229,N_2310,N_570);
or U4230 (N_4230,N_1805,N_943);
nor U4231 (N_4231,N_604,N_1512);
and U4232 (N_4232,N_2289,N_708);
nand U4233 (N_4233,N_19,N_1);
nor U4234 (N_4234,N_2394,N_472);
nand U4235 (N_4235,N_114,N_1335);
nand U4236 (N_4236,N_150,N_323);
nand U4237 (N_4237,N_1346,N_1066);
nor U4238 (N_4238,N_1357,N_2436);
or U4239 (N_4239,N_343,N_1850);
and U4240 (N_4240,N_1045,N_1631);
nor U4241 (N_4241,N_2401,N_1621);
or U4242 (N_4242,N_887,N_531);
nand U4243 (N_4243,N_2228,N_819);
and U4244 (N_4244,N_1776,N_707);
nand U4245 (N_4245,N_2092,N_1656);
and U4246 (N_4246,N_2347,N_2014);
and U4247 (N_4247,N_1606,N_302);
nand U4248 (N_4248,N_2061,N_1515);
xor U4249 (N_4249,N_1875,N_580);
nand U4250 (N_4250,N_1682,N_976);
nand U4251 (N_4251,N_576,N_1528);
and U4252 (N_4252,N_2349,N_85);
and U4253 (N_4253,N_444,N_461);
and U4254 (N_4254,N_1540,N_1829);
nor U4255 (N_4255,N_922,N_734);
or U4256 (N_4256,N_2002,N_1275);
and U4257 (N_4257,N_1321,N_1521);
and U4258 (N_4258,N_616,N_1630);
nor U4259 (N_4259,N_1147,N_422);
and U4260 (N_4260,N_675,N_2345);
or U4261 (N_4261,N_133,N_1873);
nor U4262 (N_4262,N_128,N_1989);
nand U4263 (N_4263,N_529,N_1194);
nor U4264 (N_4264,N_2481,N_2487);
and U4265 (N_4265,N_2110,N_1821);
nand U4266 (N_4266,N_753,N_1907);
nand U4267 (N_4267,N_2050,N_2103);
and U4268 (N_4268,N_1821,N_1629);
and U4269 (N_4269,N_1925,N_199);
nand U4270 (N_4270,N_208,N_895);
nor U4271 (N_4271,N_2353,N_11);
or U4272 (N_4272,N_758,N_1490);
and U4273 (N_4273,N_680,N_1776);
or U4274 (N_4274,N_877,N_1222);
xor U4275 (N_4275,N_904,N_1838);
xor U4276 (N_4276,N_506,N_19);
nand U4277 (N_4277,N_47,N_1235);
xnor U4278 (N_4278,N_1505,N_165);
nor U4279 (N_4279,N_2310,N_325);
or U4280 (N_4280,N_2395,N_2214);
or U4281 (N_4281,N_620,N_2449);
xnor U4282 (N_4282,N_1573,N_600);
or U4283 (N_4283,N_10,N_739);
and U4284 (N_4284,N_1941,N_510);
or U4285 (N_4285,N_8,N_2012);
and U4286 (N_4286,N_1149,N_1200);
nand U4287 (N_4287,N_1931,N_121);
and U4288 (N_4288,N_1691,N_173);
and U4289 (N_4289,N_2400,N_2014);
or U4290 (N_4290,N_2143,N_1622);
and U4291 (N_4291,N_951,N_935);
xnor U4292 (N_4292,N_1352,N_646);
and U4293 (N_4293,N_1236,N_1735);
or U4294 (N_4294,N_540,N_977);
nand U4295 (N_4295,N_684,N_795);
and U4296 (N_4296,N_1409,N_2311);
nand U4297 (N_4297,N_2091,N_902);
nand U4298 (N_4298,N_1001,N_862);
and U4299 (N_4299,N_2241,N_311);
and U4300 (N_4300,N_1103,N_1691);
or U4301 (N_4301,N_374,N_41);
or U4302 (N_4302,N_2435,N_2125);
nor U4303 (N_4303,N_1015,N_1830);
or U4304 (N_4304,N_915,N_378);
nand U4305 (N_4305,N_1609,N_542);
or U4306 (N_4306,N_1990,N_526);
or U4307 (N_4307,N_936,N_1944);
and U4308 (N_4308,N_2387,N_454);
nor U4309 (N_4309,N_196,N_2234);
nor U4310 (N_4310,N_464,N_1703);
and U4311 (N_4311,N_1775,N_2311);
and U4312 (N_4312,N_2137,N_1425);
nor U4313 (N_4313,N_1638,N_80);
nand U4314 (N_4314,N_2393,N_1503);
nor U4315 (N_4315,N_2171,N_1707);
or U4316 (N_4316,N_1695,N_1302);
nor U4317 (N_4317,N_1343,N_1591);
nand U4318 (N_4318,N_2365,N_2233);
nand U4319 (N_4319,N_88,N_2162);
or U4320 (N_4320,N_1467,N_1511);
nor U4321 (N_4321,N_812,N_1447);
nor U4322 (N_4322,N_1628,N_2474);
and U4323 (N_4323,N_64,N_1170);
nand U4324 (N_4324,N_43,N_2320);
or U4325 (N_4325,N_2231,N_407);
and U4326 (N_4326,N_2311,N_1282);
nand U4327 (N_4327,N_1941,N_1640);
xnor U4328 (N_4328,N_1703,N_632);
nand U4329 (N_4329,N_867,N_600);
or U4330 (N_4330,N_1798,N_1375);
and U4331 (N_4331,N_1615,N_432);
nand U4332 (N_4332,N_1858,N_598);
nand U4333 (N_4333,N_489,N_1995);
and U4334 (N_4334,N_2404,N_1281);
nor U4335 (N_4335,N_1288,N_1231);
nor U4336 (N_4336,N_1046,N_620);
or U4337 (N_4337,N_314,N_557);
nor U4338 (N_4338,N_701,N_1080);
nand U4339 (N_4339,N_265,N_1809);
or U4340 (N_4340,N_825,N_77);
nand U4341 (N_4341,N_1986,N_2439);
nand U4342 (N_4342,N_1201,N_294);
nor U4343 (N_4343,N_1236,N_694);
or U4344 (N_4344,N_2019,N_775);
xnor U4345 (N_4345,N_1899,N_415);
xnor U4346 (N_4346,N_2206,N_1687);
nand U4347 (N_4347,N_1741,N_2188);
and U4348 (N_4348,N_1465,N_2356);
and U4349 (N_4349,N_980,N_1978);
or U4350 (N_4350,N_822,N_452);
nor U4351 (N_4351,N_1141,N_117);
xor U4352 (N_4352,N_1648,N_2440);
nor U4353 (N_4353,N_704,N_1671);
nor U4354 (N_4354,N_2150,N_164);
nand U4355 (N_4355,N_600,N_1812);
nor U4356 (N_4356,N_2403,N_963);
nand U4357 (N_4357,N_996,N_504);
or U4358 (N_4358,N_946,N_1976);
xnor U4359 (N_4359,N_1652,N_1399);
nand U4360 (N_4360,N_607,N_2014);
nor U4361 (N_4361,N_363,N_200);
and U4362 (N_4362,N_1749,N_1807);
or U4363 (N_4363,N_1745,N_2219);
nor U4364 (N_4364,N_1668,N_1354);
and U4365 (N_4365,N_190,N_2424);
nand U4366 (N_4366,N_159,N_863);
and U4367 (N_4367,N_1059,N_890);
or U4368 (N_4368,N_1158,N_373);
nand U4369 (N_4369,N_2475,N_2107);
nand U4370 (N_4370,N_215,N_1230);
and U4371 (N_4371,N_2226,N_1568);
nand U4372 (N_4372,N_398,N_935);
and U4373 (N_4373,N_2451,N_2376);
nor U4374 (N_4374,N_2353,N_934);
nand U4375 (N_4375,N_75,N_178);
nor U4376 (N_4376,N_472,N_1193);
or U4377 (N_4377,N_191,N_2386);
xnor U4378 (N_4378,N_1713,N_689);
and U4379 (N_4379,N_1749,N_2497);
xor U4380 (N_4380,N_2360,N_127);
and U4381 (N_4381,N_2485,N_1047);
or U4382 (N_4382,N_473,N_1468);
or U4383 (N_4383,N_1563,N_763);
or U4384 (N_4384,N_2235,N_1823);
and U4385 (N_4385,N_615,N_1998);
and U4386 (N_4386,N_1293,N_108);
or U4387 (N_4387,N_2367,N_14);
nand U4388 (N_4388,N_1243,N_602);
and U4389 (N_4389,N_564,N_1525);
or U4390 (N_4390,N_1062,N_999);
nand U4391 (N_4391,N_2061,N_1301);
nor U4392 (N_4392,N_1746,N_2147);
nor U4393 (N_4393,N_934,N_764);
nor U4394 (N_4394,N_1408,N_923);
and U4395 (N_4395,N_848,N_972);
nor U4396 (N_4396,N_785,N_588);
xnor U4397 (N_4397,N_1639,N_1073);
nand U4398 (N_4398,N_1875,N_976);
nand U4399 (N_4399,N_861,N_1359);
nand U4400 (N_4400,N_566,N_258);
nand U4401 (N_4401,N_783,N_879);
nand U4402 (N_4402,N_393,N_1262);
nor U4403 (N_4403,N_1054,N_1895);
nand U4404 (N_4404,N_1342,N_558);
or U4405 (N_4405,N_708,N_769);
and U4406 (N_4406,N_1411,N_2428);
nand U4407 (N_4407,N_1175,N_2165);
nor U4408 (N_4408,N_964,N_2421);
or U4409 (N_4409,N_1412,N_1665);
or U4410 (N_4410,N_1287,N_76);
nor U4411 (N_4411,N_1357,N_112);
or U4412 (N_4412,N_1907,N_406);
nand U4413 (N_4413,N_975,N_137);
or U4414 (N_4414,N_2075,N_1669);
and U4415 (N_4415,N_654,N_1827);
nor U4416 (N_4416,N_295,N_450);
or U4417 (N_4417,N_1617,N_336);
nor U4418 (N_4418,N_2018,N_283);
or U4419 (N_4419,N_949,N_224);
or U4420 (N_4420,N_1811,N_1472);
nand U4421 (N_4421,N_1797,N_1916);
nor U4422 (N_4422,N_1081,N_1107);
xor U4423 (N_4423,N_1435,N_2055);
nor U4424 (N_4424,N_1142,N_351);
nor U4425 (N_4425,N_2469,N_123);
or U4426 (N_4426,N_2455,N_1136);
nand U4427 (N_4427,N_1488,N_2436);
nand U4428 (N_4428,N_1840,N_196);
nor U4429 (N_4429,N_2462,N_595);
nor U4430 (N_4430,N_163,N_1567);
nand U4431 (N_4431,N_1686,N_2450);
or U4432 (N_4432,N_592,N_997);
or U4433 (N_4433,N_1922,N_3);
and U4434 (N_4434,N_1745,N_71);
xnor U4435 (N_4435,N_613,N_2228);
nor U4436 (N_4436,N_2266,N_1357);
nor U4437 (N_4437,N_2422,N_2101);
nor U4438 (N_4438,N_472,N_2372);
or U4439 (N_4439,N_1004,N_2176);
nand U4440 (N_4440,N_1059,N_1272);
nand U4441 (N_4441,N_2045,N_2346);
or U4442 (N_4442,N_844,N_522);
nor U4443 (N_4443,N_854,N_189);
nand U4444 (N_4444,N_1141,N_1462);
nor U4445 (N_4445,N_1829,N_771);
nand U4446 (N_4446,N_1559,N_1542);
xnor U4447 (N_4447,N_2330,N_1636);
nand U4448 (N_4448,N_325,N_1113);
or U4449 (N_4449,N_867,N_1501);
and U4450 (N_4450,N_1078,N_98);
and U4451 (N_4451,N_1001,N_316);
and U4452 (N_4452,N_2246,N_1211);
or U4453 (N_4453,N_2183,N_180);
xnor U4454 (N_4454,N_1533,N_1757);
xor U4455 (N_4455,N_1580,N_1144);
nand U4456 (N_4456,N_1184,N_1965);
nand U4457 (N_4457,N_1694,N_611);
or U4458 (N_4458,N_313,N_812);
nor U4459 (N_4459,N_2406,N_884);
and U4460 (N_4460,N_1547,N_2213);
nand U4461 (N_4461,N_2298,N_2418);
nor U4462 (N_4462,N_267,N_1130);
nor U4463 (N_4463,N_463,N_952);
nor U4464 (N_4464,N_2025,N_2462);
nand U4465 (N_4465,N_1404,N_820);
and U4466 (N_4466,N_2278,N_2444);
or U4467 (N_4467,N_1706,N_351);
or U4468 (N_4468,N_662,N_1241);
xnor U4469 (N_4469,N_737,N_831);
nand U4470 (N_4470,N_1798,N_429);
or U4471 (N_4471,N_693,N_20);
nor U4472 (N_4472,N_1825,N_1669);
or U4473 (N_4473,N_1377,N_1570);
nor U4474 (N_4474,N_1992,N_702);
and U4475 (N_4475,N_2255,N_1768);
nor U4476 (N_4476,N_2377,N_220);
nand U4477 (N_4477,N_2274,N_1584);
and U4478 (N_4478,N_1177,N_1311);
or U4479 (N_4479,N_2306,N_891);
nor U4480 (N_4480,N_1850,N_542);
and U4481 (N_4481,N_1495,N_1236);
nor U4482 (N_4482,N_1750,N_885);
nor U4483 (N_4483,N_1146,N_1041);
or U4484 (N_4484,N_431,N_1972);
nor U4485 (N_4485,N_2106,N_1571);
nor U4486 (N_4486,N_521,N_193);
xor U4487 (N_4487,N_1570,N_954);
nand U4488 (N_4488,N_838,N_1164);
nor U4489 (N_4489,N_264,N_1444);
and U4490 (N_4490,N_157,N_900);
and U4491 (N_4491,N_2000,N_1512);
nand U4492 (N_4492,N_944,N_278);
xor U4493 (N_4493,N_1654,N_1823);
and U4494 (N_4494,N_2053,N_1616);
or U4495 (N_4495,N_612,N_2429);
and U4496 (N_4496,N_538,N_363);
nand U4497 (N_4497,N_1966,N_517);
or U4498 (N_4498,N_728,N_302);
or U4499 (N_4499,N_39,N_112);
or U4500 (N_4500,N_2399,N_83);
or U4501 (N_4501,N_2281,N_2225);
xnor U4502 (N_4502,N_2323,N_689);
or U4503 (N_4503,N_1178,N_2365);
nor U4504 (N_4504,N_964,N_1455);
and U4505 (N_4505,N_130,N_1350);
nand U4506 (N_4506,N_2204,N_1628);
xnor U4507 (N_4507,N_60,N_2160);
or U4508 (N_4508,N_1115,N_1730);
nor U4509 (N_4509,N_1564,N_1394);
nor U4510 (N_4510,N_377,N_234);
nor U4511 (N_4511,N_2320,N_610);
nand U4512 (N_4512,N_1355,N_916);
nor U4513 (N_4513,N_2356,N_669);
and U4514 (N_4514,N_349,N_520);
or U4515 (N_4515,N_2067,N_1987);
nor U4516 (N_4516,N_1578,N_1703);
or U4517 (N_4517,N_937,N_448);
nand U4518 (N_4518,N_2249,N_972);
nand U4519 (N_4519,N_933,N_607);
xnor U4520 (N_4520,N_2323,N_2101);
and U4521 (N_4521,N_9,N_303);
nor U4522 (N_4522,N_2272,N_631);
nand U4523 (N_4523,N_149,N_979);
nor U4524 (N_4524,N_1165,N_512);
nor U4525 (N_4525,N_258,N_540);
nand U4526 (N_4526,N_798,N_191);
nand U4527 (N_4527,N_677,N_834);
nor U4528 (N_4528,N_986,N_267);
and U4529 (N_4529,N_2497,N_763);
nand U4530 (N_4530,N_1511,N_1879);
nand U4531 (N_4531,N_1535,N_1843);
and U4532 (N_4532,N_1140,N_310);
nand U4533 (N_4533,N_1017,N_1479);
nor U4534 (N_4534,N_2239,N_1608);
nor U4535 (N_4535,N_986,N_386);
and U4536 (N_4536,N_2496,N_1657);
or U4537 (N_4537,N_628,N_2357);
or U4538 (N_4538,N_118,N_932);
nand U4539 (N_4539,N_156,N_1796);
nand U4540 (N_4540,N_1203,N_2018);
nand U4541 (N_4541,N_1535,N_426);
and U4542 (N_4542,N_1840,N_564);
nor U4543 (N_4543,N_785,N_1331);
and U4544 (N_4544,N_1653,N_489);
nand U4545 (N_4545,N_461,N_801);
nand U4546 (N_4546,N_302,N_1999);
or U4547 (N_4547,N_1927,N_1322);
and U4548 (N_4548,N_468,N_1774);
nor U4549 (N_4549,N_1266,N_1508);
or U4550 (N_4550,N_1585,N_664);
xnor U4551 (N_4551,N_1246,N_273);
or U4552 (N_4552,N_1392,N_2450);
or U4553 (N_4553,N_1284,N_1444);
and U4554 (N_4554,N_1646,N_1680);
nand U4555 (N_4555,N_1877,N_1607);
nand U4556 (N_4556,N_2015,N_755);
nor U4557 (N_4557,N_612,N_2286);
xor U4558 (N_4558,N_853,N_447);
nand U4559 (N_4559,N_1439,N_358);
nand U4560 (N_4560,N_2322,N_1448);
and U4561 (N_4561,N_2436,N_1965);
nand U4562 (N_4562,N_79,N_590);
or U4563 (N_4563,N_487,N_1358);
and U4564 (N_4564,N_9,N_442);
and U4565 (N_4565,N_449,N_2114);
nand U4566 (N_4566,N_1188,N_1755);
nand U4567 (N_4567,N_877,N_1480);
and U4568 (N_4568,N_1813,N_1341);
xnor U4569 (N_4569,N_1230,N_1346);
and U4570 (N_4570,N_1971,N_1570);
or U4571 (N_4571,N_1133,N_133);
or U4572 (N_4572,N_792,N_2133);
or U4573 (N_4573,N_768,N_679);
xnor U4574 (N_4574,N_395,N_1447);
or U4575 (N_4575,N_1278,N_146);
nor U4576 (N_4576,N_1253,N_1938);
or U4577 (N_4577,N_1104,N_1584);
xor U4578 (N_4578,N_1299,N_401);
and U4579 (N_4579,N_2101,N_1428);
nor U4580 (N_4580,N_1178,N_1614);
xor U4581 (N_4581,N_215,N_54);
nor U4582 (N_4582,N_1869,N_1502);
and U4583 (N_4583,N_480,N_2014);
nand U4584 (N_4584,N_357,N_1595);
nor U4585 (N_4585,N_1875,N_2349);
and U4586 (N_4586,N_103,N_1271);
nor U4587 (N_4587,N_911,N_1815);
nor U4588 (N_4588,N_1976,N_1879);
xor U4589 (N_4589,N_1428,N_49);
or U4590 (N_4590,N_148,N_360);
or U4591 (N_4591,N_861,N_2244);
or U4592 (N_4592,N_1477,N_168);
nand U4593 (N_4593,N_1490,N_1774);
nand U4594 (N_4594,N_303,N_337);
nor U4595 (N_4595,N_1258,N_2298);
nand U4596 (N_4596,N_1075,N_1652);
and U4597 (N_4597,N_1222,N_2440);
nor U4598 (N_4598,N_1788,N_1029);
and U4599 (N_4599,N_483,N_2138);
or U4600 (N_4600,N_923,N_1634);
or U4601 (N_4601,N_224,N_218);
nor U4602 (N_4602,N_2146,N_745);
and U4603 (N_4603,N_328,N_840);
or U4604 (N_4604,N_1097,N_7);
and U4605 (N_4605,N_1339,N_2273);
nand U4606 (N_4606,N_572,N_994);
or U4607 (N_4607,N_996,N_977);
nor U4608 (N_4608,N_674,N_1693);
or U4609 (N_4609,N_1168,N_1761);
or U4610 (N_4610,N_891,N_1236);
or U4611 (N_4611,N_2129,N_1758);
nand U4612 (N_4612,N_900,N_1582);
or U4613 (N_4613,N_76,N_100);
nand U4614 (N_4614,N_1877,N_2472);
xnor U4615 (N_4615,N_1816,N_1106);
and U4616 (N_4616,N_247,N_849);
nor U4617 (N_4617,N_1799,N_2103);
nand U4618 (N_4618,N_2010,N_1020);
and U4619 (N_4619,N_1179,N_510);
nand U4620 (N_4620,N_1618,N_1938);
nand U4621 (N_4621,N_2306,N_561);
and U4622 (N_4622,N_1485,N_2172);
and U4623 (N_4623,N_1321,N_24);
nand U4624 (N_4624,N_1970,N_2043);
xor U4625 (N_4625,N_212,N_1699);
or U4626 (N_4626,N_1524,N_1122);
nor U4627 (N_4627,N_1590,N_105);
nand U4628 (N_4628,N_1742,N_2222);
nor U4629 (N_4629,N_1647,N_1689);
nor U4630 (N_4630,N_1561,N_130);
or U4631 (N_4631,N_1747,N_2275);
nor U4632 (N_4632,N_299,N_852);
nand U4633 (N_4633,N_2138,N_825);
or U4634 (N_4634,N_1529,N_1693);
or U4635 (N_4635,N_289,N_448);
nand U4636 (N_4636,N_2050,N_2317);
or U4637 (N_4637,N_269,N_2437);
and U4638 (N_4638,N_1284,N_2183);
xor U4639 (N_4639,N_995,N_1);
nor U4640 (N_4640,N_949,N_1686);
and U4641 (N_4641,N_2426,N_728);
xnor U4642 (N_4642,N_1115,N_475);
nand U4643 (N_4643,N_755,N_356);
nor U4644 (N_4644,N_1821,N_259);
nand U4645 (N_4645,N_2434,N_2370);
xor U4646 (N_4646,N_1400,N_2087);
xor U4647 (N_4647,N_1618,N_311);
nand U4648 (N_4648,N_2402,N_34);
nand U4649 (N_4649,N_1202,N_1991);
nor U4650 (N_4650,N_76,N_605);
nor U4651 (N_4651,N_2082,N_1411);
nor U4652 (N_4652,N_158,N_2261);
nand U4653 (N_4653,N_2183,N_2227);
nand U4654 (N_4654,N_2426,N_71);
nand U4655 (N_4655,N_1418,N_1347);
and U4656 (N_4656,N_1983,N_840);
and U4657 (N_4657,N_2273,N_322);
and U4658 (N_4658,N_1158,N_150);
nand U4659 (N_4659,N_1177,N_1413);
nand U4660 (N_4660,N_735,N_170);
or U4661 (N_4661,N_1405,N_280);
or U4662 (N_4662,N_2144,N_782);
and U4663 (N_4663,N_276,N_165);
or U4664 (N_4664,N_1857,N_2087);
and U4665 (N_4665,N_1544,N_1641);
and U4666 (N_4666,N_1641,N_1410);
nor U4667 (N_4667,N_497,N_1459);
and U4668 (N_4668,N_517,N_619);
nand U4669 (N_4669,N_1415,N_2074);
nand U4670 (N_4670,N_405,N_141);
and U4671 (N_4671,N_806,N_1465);
and U4672 (N_4672,N_919,N_1117);
and U4673 (N_4673,N_1947,N_985);
and U4674 (N_4674,N_1026,N_462);
or U4675 (N_4675,N_757,N_597);
nor U4676 (N_4676,N_2168,N_2042);
or U4677 (N_4677,N_973,N_422);
or U4678 (N_4678,N_1780,N_2334);
or U4679 (N_4679,N_1386,N_1554);
nor U4680 (N_4680,N_891,N_394);
and U4681 (N_4681,N_1590,N_146);
or U4682 (N_4682,N_2265,N_290);
and U4683 (N_4683,N_139,N_1073);
nor U4684 (N_4684,N_2432,N_1255);
or U4685 (N_4685,N_2099,N_704);
xor U4686 (N_4686,N_1913,N_265);
nor U4687 (N_4687,N_1876,N_113);
and U4688 (N_4688,N_871,N_777);
nand U4689 (N_4689,N_1619,N_566);
nor U4690 (N_4690,N_818,N_2264);
or U4691 (N_4691,N_2283,N_716);
nand U4692 (N_4692,N_2259,N_1663);
nand U4693 (N_4693,N_359,N_730);
nand U4694 (N_4694,N_313,N_1007);
nor U4695 (N_4695,N_2262,N_514);
or U4696 (N_4696,N_2003,N_811);
or U4697 (N_4697,N_805,N_1929);
and U4698 (N_4698,N_261,N_1362);
nand U4699 (N_4699,N_1705,N_1059);
or U4700 (N_4700,N_31,N_526);
or U4701 (N_4701,N_1926,N_1260);
nor U4702 (N_4702,N_510,N_960);
nor U4703 (N_4703,N_616,N_107);
nand U4704 (N_4704,N_1611,N_1523);
and U4705 (N_4705,N_2404,N_884);
and U4706 (N_4706,N_137,N_307);
and U4707 (N_4707,N_2366,N_957);
nand U4708 (N_4708,N_182,N_908);
nor U4709 (N_4709,N_1525,N_1073);
or U4710 (N_4710,N_651,N_1977);
or U4711 (N_4711,N_523,N_14);
and U4712 (N_4712,N_1023,N_668);
and U4713 (N_4713,N_2373,N_1713);
nor U4714 (N_4714,N_754,N_2212);
nor U4715 (N_4715,N_52,N_694);
xnor U4716 (N_4716,N_856,N_831);
and U4717 (N_4717,N_2228,N_1099);
and U4718 (N_4718,N_1867,N_2049);
or U4719 (N_4719,N_1027,N_733);
xnor U4720 (N_4720,N_201,N_1910);
or U4721 (N_4721,N_1293,N_548);
nand U4722 (N_4722,N_449,N_2470);
and U4723 (N_4723,N_556,N_1736);
and U4724 (N_4724,N_1985,N_811);
and U4725 (N_4725,N_1415,N_1143);
or U4726 (N_4726,N_1179,N_1110);
and U4727 (N_4727,N_952,N_162);
nor U4728 (N_4728,N_2100,N_250);
nor U4729 (N_4729,N_1938,N_554);
xnor U4730 (N_4730,N_929,N_106);
and U4731 (N_4731,N_1427,N_1816);
or U4732 (N_4732,N_685,N_1827);
nand U4733 (N_4733,N_241,N_838);
or U4734 (N_4734,N_2083,N_2293);
and U4735 (N_4735,N_2496,N_1510);
nand U4736 (N_4736,N_1852,N_345);
xor U4737 (N_4737,N_1196,N_1332);
nand U4738 (N_4738,N_1505,N_182);
nor U4739 (N_4739,N_1962,N_1398);
or U4740 (N_4740,N_161,N_2310);
or U4741 (N_4741,N_1123,N_310);
xor U4742 (N_4742,N_246,N_1289);
xor U4743 (N_4743,N_783,N_1373);
nor U4744 (N_4744,N_2261,N_924);
or U4745 (N_4745,N_1900,N_1339);
nor U4746 (N_4746,N_1078,N_781);
nor U4747 (N_4747,N_1251,N_416);
and U4748 (N_4748,N_2495,N_517);
nand U4749 (N_4749,N_1929,N_1600);
nor U4750 (N_4750,N_2213,N_614);
or U4751 (N_4751,N_570,N_1473);
and U4752 (N_4752,N_2405,N_631);
xor U4753 (N_4753,N_801,N_2226);
nor U4754 (N_4754,N_2018,N_2294);
nor U4755 (N_4755,N_1379,N_2376);
or U4756 (N_4756,N_1373,N_1227);
and U4757 (N_4757,N_2426,N_631);
and U4758 (N_4758,N_343,N_723);
and U4759 (N_4759,N_1991,N_1156);
nand U4760 (N_4760,N_1107,N_971);
nand U4761 (N_4761,N_2390,N_2133);
xor U4762 (N_4762,N_2005,N_451);
xor U4763 (N_4763,N_108,N_203);
xnor U4764 (N_4764,N_899,N_970);
or U4765 (N_4765,N_1398,N_1926);
xnor U4766 (N_4766,N_447,N_912);
or U4767 (N_4767,N_1440,N_579);
nor U4768 (N_4768,N_786,N_1552);
nand U4769 (N_4769,N_2054,N_1184);
xnor U4770 (N_4770,N_58,N_1270);
xor U4771 (N_4771,N_1791,N_16);
nor U4772 (N_4772,N_2474,N_663);
nand U4773 (N_4773,N_699,N_1562);
nand U4774 (N_4774,N_917,N_409);
xnor U4775 (N_4775,N_2374,N_1129);
and U4776 (N_4776,N_798,N_1580);
or U4777 (N_4777,N_2428,N_2123);
nor U4778 (N_4778,N_13,N_2423);
nor U4779 (N_4779,N_782,N_943);
nor U4780 (N_4780,N_687,N_128);
nand U4781 (N_4781,N_782,N_1589);
nor U4782 (N_4782,N_2371,N_1515);
xnor U4783 (N_4783,N_116,N_674);
or U4784 (N_4784,N_2009,N_1425);
or U4785 (N_4785,N_42,N_1500);
or U4786 (N_4786,N_1829,N_935);
nand U4787 (N_4787,N_1816,N_1772);
nand U4788 (N_4788,N_259,N_1905);
nand U4789 (N_4789,N_2397,N_2241);
nor U4790 (N_4790,N_665,N_1814);
nand U4791 (N_4791,N_367,N_2071);
nor U4792 (N_4792,N_2428,N_554);
nor U4793 (N_4793,N_2232,N_1254);
and U4794 (N_4794,N_2220,N_1550);
and U4795 (N_4795,N_1471,N_297);
nor U4796 (N_4796,N_260,N_2411);
and U4797 (N_4797,N_689,N_1785);
or U4798 (N_4798,N_2330,N_192);
or U4799 (N_4799,N_1983,N_1711);
xor U4800 (N_4800,N_1486,N_936);
nor U4801 (N_4801,N_498,N_982);
xnor U4802 (N_4802,N_668,N_1434);
xor U4803 (N_4803,N_479,N_74);
nor U4804 (N_4804,N_1777,N_1204);
nand U4805 (N_4805,N_2386,N_2405);
and U4806 (N_4806,N_1866,N_2023);
nor U4807 (N_4807,N_670,N_1609);
or U4808 (N_4808,N_617,N_1853);
nor U4809 (N_4809,N_1067,N_1251);
or U4810 (N_4810,N_1803,N_968);
nor U4811 (N_4811,N_1598,N_104);
nor U4812 (N_4812,N_1487,N_341);
and U4813 (N_4813,N_1389,N_2397);
xor U4814 (N_4814,N_1447,N_537);
xnor U4815 (N_4815,N_1703,N_324);
and U4816 (N_4816,N_388,N_1985);
nand U4817 (N_4817,N_1336,N_1171);
nand U4818 (N_4818,N_2452,N_1555);
nor U4819 (N_4819,N_507,N_1941);
nor U4820 (N_4820,N_1346,N_322);
nand U4821 (N_4821,N_746,N_1428);
nand U4822 (N_4822,N_661,N_1545);
and U4823 (N_4823,N_1903,N_1600);
and U4824 (N_4824,N_431,N_425);
xnor U4825 (N_4825,N_2030,N_2417);
nand U4826 (N_4826,N_2114,N_1536);
nor U4827 (N_4827,N_2036,N_68);
nor U4828 (N_4828,N_512,N_708);
or U4829 (N_4829,N_243,N_55);
nand U4830 (N_4830,N_1467,N_531);
xnor U4831 (N_4831,N_130,N_289);
xor U4832 (N_4832,N_1666,N_791);
nand U4833 (N_4833,N_313,N_2121);
or U4834 (N_4834,N_967,N_1826);
and U4835 (N_4835,N_2222,N_1868);
and U4836 (N_4836,N_1838,N_1297);
nor U4837 (N_4837,N_1879,N_1241);
nor U4838 (N_4838,N_894,N_174);
nor U4839 (N_4839,N_2209,N_1521);
and U4840 (N_4840,N_2283,N_2076);
or U4841 (N_4841,N_891,N_1233);
or U4842 (N_4842,N_270,N_2146);
or U4843 (N_4843,N_1875,N_1253);
nand U4844 (N_4844,N_2243,N_1166);
nor U4845 (N_4845,N_541,N_2195);
nor U4846 (N_4846,N_1136,N_1138);
nand U4847 (N_4847,N_2071,N_2045);
nand U4848 (N_4848,N_1514,N_2127);
or U4849 (N_4849,N_1520,N_2259);
nor U4850 (N_4850,N_2169,N_1503);
xor U4851 (N_4851,N_1303,N_2235);
nor U4852 (N_4852,N_7,N_2110);
and U4853 (N_4853,N_2301,N_1531);
nor U4854 (N_4854,N_1525,N_1333);
nand U4855 (N_4855,N_2110,N_1549);
or U4856 (N_4856,N_2495,N_1496);
or U4857 (N_4857,N_1755,N_555);
and U4858 (N_4858,N_1220,N_2118);
nand U4859 (N_4859,N_422,N_702);
or U4860 (N_4860,N_1617,N_1590);
and U4861 (N_4861,N_2330,N_1020);
or U4862 (N_4862,N_310,N_1397);
or U4863 (N_4863,N_2294,N_18);
and U4864 (N_4864,N_1861,N_1510);
or U4865 (N_4865,N_1402,N_1980);
nand U4866 (N_4866,N_112,N_242);
or U4867 (N_4867,N_1725,N_681);
nand U4868 (N_4868,N_2240,N_2034);
nor U4869 (N_4869,N_1464,N_675);
nor U4870 (N_4870,N_1403,N_821);
or U4871 (N_4871,N_1893,N_2147);
nor U4872 (N_4872,N_478,N_2431);
nand U4873 (N_4873,N_2036,N_2446);
nor U4874 (N_4874,N_1601,N_1559);
nand U4875 (N_4875,N_2054,N_393);
or U4876 (N_4876,N_2180,N_246);
and U4877 (N_4877,N_2113,N_950);
or U4878 (N_4878,N_416,N_786);
and U4879 (N_4879,N_1149,N_1633);
or U4880 (N_4880,N_287,N_718);
or U4881 (N_4881,N_1041,N_2328);
nor U4882 (N_4882,N_2100,N_2377);
and U4883 (N_4883,N_912,N_787);
nand U4884 (N_4884,N_875,N_649);
nor U4885 (N_4885,N_1236,N_794);
nand U4886 (N_4886,N_1719,N_355);
or U4887 (N_4887,N_1475,N_1095);
or U4888 (N_4888,N_1914,N_1524);
nand U4889 (N_4889,N_759,N_1285);
and U4890 (N_4890,N_513,N_265);
or U4891 (N_4891,N_105,N_419);
nor U4892 (N_4892,N_184,N_1062);
and U4893 (N_4893,N_1829,N_1212);
and U4894 (N_4894,N_317,N_402);
xnor U4895 (N_4895,N_1020,N_572);
nor U4896 (N_4896,N_1221,N_616);
and U4897 (N_4897,N_139,N_2380);
nor U4898 (N_4898,N_1520,N_2373);
and U4899 (N_4899,N_1531,N_858);
and U4900 (N_4900,N_728,N_1709);
and U4901 (N_4901,N_1955,N_1363);
nand U4902 (N_4902,N_1591,N_605);
nor U4903 (N_4903,N_1547,N_349);
xnor U4904 (N_4904,N_796,N_545);
nor U4905 (N_4905,N_831,N_1932);
and U4906 (N_4906,N_1556,N_1927);
nand U4907 (N_4907,N_653,N_1031);
nand U4908 (N_4908,N_1493,N_632);
or U4909 (N_4909,N_1716,N_1913);
or U4910 (N_4910,N_813,N_1580);
nand U4911 (N_4911,N_859,N_530);
and U4912 (N_4912,N_314,N_1310);
nand U4913 (N_4913,N_1202,N_489);
nor U4914 (N_4914,N_2469,N_2182);
xnor U4915 (N_4915,N_2189,N_2451);
and U4916 (N_4916,N_2440,N_2231);
nor U4917 (N_4917,N_1595,N_422);
or U4918 (N_4918,N_1123,N_1548);
nand U4919 (N_4919,N_13,N_1245);
or U4920 (N_4920,N_2120,N_1261);
or U4921 (N_4921,N_1862,N_676);
nand U4922 (N_4922,N_1812,N_1421);
or U4923 (N_4923,N_753,N_2465);
nand U4924 (N_4924,N_2247,N_2329);
or U4925 (N_4925,N_925,N_1615);
and U4926 (N_4926,N_1138,N_2375);
nor U4927 (N_4927,N_1308,N_18);
xnor U4928 (N_4928,N_1923,N_626);
xnor U4929 (N_4929,N_1268,N_1794);
nand U4930 (N_4930,N_2144,N_1636);
nor U4931 (N_4931,N_2185,N_547);
or U4932 (N_4932,N_1558,N_621);
and U4933 (N_4933,N_2300,N_1410);
nand U4934 (N_4934,N_306,N_178);
and U4935 (N_4935,N_1217,N_717);
and U4936 (N_4936,N_2115,N_453);
nand U4937 (N_4937,N_12,N_235);
and U4938 (N_4938,N_1749,N_1374);
nor U4939 (N_4939,N_2496,N_1930);
and U4940 (N_4940,N_363,N_1538);
nand U4941 (N_4941,N_1292,N_1699);
nor U4942 (N_4942,N_2385,N_487);
and U4943 (N_4943,N_1856,N_2058);
nand U4944 (N_4944,N_1795,N_2395);
xor U4945 (N_4945,N_1757,N_1744);
nor U4946 (N_4946,N_490,N_33);
nor U4947 (N_4947,N_242,N_728);
nor U4948 (N_4948,N_685,N_1193);
and U4949 (N_4949,N_899,N_321);
nor U4950 (N_4950,N_1329,N_1263);
or U4951 (N_4951,N_1084,N_871);
nor U4952 (N_4952,N_1133,N_661);
nor U4953 (N_4953,N_452,N_2321);
or U4954 (N_4954,N_2395,N_1882);
nand U4955 (N_4955,N_1330,N_150);
nand U4956 (N_4956,N_1974,N_62);
nand U4957 (N_4957,N_2318,N_2426);
and U4958 (N_4958,N_1811,N_1835);
or U4959 (N_4959,N_2149,N_1109);
nand U4960 (N_4960,N_728,N_1229);
nor U4961 (N_4961,N_2230,N_2450);
and U4962 (N_4962,N_1692,N_607);
nor U4963 (N_4963,N_1404,N_1098);
nand U4964 (N_4964,N_182,N_244);
nand U4965 (N_4965,N_2402,N_447);
nor U4966 (N_4966,N_1395,N_102);
nor U4967 (N_4967,N_1355,N_2197);
nand U4968 (N_4968,N_1858,N_951);
or U4969 (N_4969,N_1721,N_1563);
and U4970 (N_4970,N_1873,N_1930);
and U4971 (N_4971,N_481,N_1839);
nand U4972 (N_4972,N_917,N_2092);
or U4973 (N_4973,N_572,N_162);
or U4974 (N_4974,N_1505,N_1081);
or U4975 (N_4975,N_515,N_2160);
and U4976 (N_4976,N_340,N_175);
nand U4977 (N_4977,N_2359,N_960);
nor U4978 (N_4978,N_882,N_1396);
or U4979 (N_4979,N_1028,N_106);
or U4980 (N_4980,N_640,N_2054);
nor U4981 (N_4981,N_1713,N_590);
or U4982 (N_4982,N_502,N_509);
and U4983 (N_4983,N_193,N_415);
and U4984 (N_4984,N_399,N_1529);
and U4985 (N_4985,N_2048,N_2349);
nand U4986 (N_4986,N_1134,N_2221);
or U4987 (N_4987,N_147,N_1137);
nand U4988 (N_4988,N_655,N_63);
nand U4989 (N_4989,N_2169,N_535);
and U4990 (N_4990,N_1867,N_1060);
and U4991 (N_4991,N_1342,N_2454);
nand U4992 (N_4992,N_1780,N_2293);
nand U4993 (N_4993,N_1906,N_367);
nor U4994 (N_4994,N_1641,N_2321);
and U4995 (N_4995,N_641,N_796);
nand U4996 (N_4996,N_1553,N_919);
and U4997 (N_4997,N_1732,N_2294);
nor U4998 (N_4998,N_1967,N_130);
xor U4999 (N_4999,N_167,N_2300);
and UO_0 (O_0,N_3866,N_3392);
and UO_1 (O_1,N_4364,N_4995);
and UO_2 (O_2,N_3921,N_4814);
nand UO_3 (O_3,N_3028,N_3374);
or UO_4 (O_4,N_4394,N_3357);
or UO_5 (O_5,N_4152,N_3430);
and UO_6 (O_6,N_3301,N_4699);
nor UO_7 (O_7,N_4883,N_3247);
or UO_8 (O_8,N_3932,N_4062);
or UO_9 (O_9,N_3704,N_2706);
nand UO_10 (O_10,N_4164,N_4983);
or UO_11 (O_11,N_3369,N_3012);
and UO_12 (O_12,N_3300,N_3626);
and UO_13 (O_13,N_3187,N_4874);
or UO_14 (O_14,N_4269,N_4620);
nand UO_15 (O_15,N_2507,N_4854);
and UO_16 (O_16,N_2901,N_3585);
and UO_17 (O_17,N_4585,N_3328);
nand UO_18 (O_18,N_4968,N_2638);
nand UO_19 (O_19,N_3894,N_3453);
and UO_20 (O_20,N_3423,N_3077);
or UO_21 (O_21,N_4352,N_3755);
nand UO_22 (O_22,N_4050,N_4093);
nand UO_23 (O_23,N_3769,N_2511);
xor UO_24 (O_24,N_4345,N_2929);
nor UO_25 (O_25,N_2877,N_3182);
nor UO_26 (O_26,N_4197,N_4135);
or UO_27 (O_27,N_4010,N_4675);
and UO_28 (O_28,N_4739,N_4310);
and UO_29 (O_29,N_4711,N_4268);
nor UO_30 (O_30,N_3327,N_4542);
or UO_31 (O_31,N_3779,N_2547);
or UO_32 (O_32,N_2839,N_3587);
nand UO_33 (O_33,N_2920,N_4970);
nand UO_34 (O_34,N_3641,N_4733);
or UO_35 (O_35,N_4791,N_4473);
nor UO_36 (O_36,N_3265,N_3771);
nand UO_37 (O_37,N_4304,N_4602);
or UO_38 (O_38,N_4499,N_4119);
nor UO_39 (O_39,N_4833,N_4834);
xnor UO_40 (O_40,N_3025,N_4392);
and UO_41 (O_41,N_2767,N_3426);
nor UO_42 (O_42,N_4785,N_3526);
nand UO_43 (O_43,N_2912,N_3211);
and UO_44 (O_44,N_4934,N_3765);
or UO_45 (O_45,N_3793,N_4303);
nor UO_46 (O_46,N_4242,N_4336);
xnor UO_47 (O_47,N_3570,N_3097);
and UO_48 (O_48,N_2632,N_3183);
nor UO_49 (O_49,N_2945,N_2809);
and UO_50 (O_50,N_4532,N_3829);
or UO_51 (O_51,N_3917,N_2512);
or UO_52 (O_52,N_4745,N_4090);
nand UO_53 (O_53,N_3719,N_3498);
or UO_54 (O_54,N_3472,N_3997);
nand UO_55 (O_55,N_4491,N_4348);
nor UO_56 (O_56,N_4070,N_4153);
or UO_57 (O_57,N_3937,N_4965);
and UO_58 (O_58,N_2539,N_2663);
or UO_59 (O_59,N_4341,N_4755);
or UO_60 (O_60,N_4158,N_3216);
nor UO_61 (O_61,N_4233,N_4969);
and UO_62 (O_62,N_3804,N_4365);
or UO_63 (O_63,N_2986,N_4860);
nand UO_64 (O_64,N_4537,N_2600);
and UO_65 (O_65,N_4820,N_4801);
nor UO_66 (O_66,N_4068,N_2922);
and UO_67 (O_67,N_3344,N_3745);
or UO_68 (O_68,N_3321,N_4942);
and UO_69 (O_69,N_2722,N_3831);
and UO_70 (O_70,N_4492,N_4004);
nand UO_71 (O_71,N_4538,N_3574);
and UO_72 (O_72,N_3819,N_4139);
or UO_73 (O_73,N_3249,N_4835);
xor UO_74 (O_74,N_4754,N_4555);
or UO_75 (O_75,N_2564,N_4918);
or UO_76 (O_76,N_2674,N_3001);
nand UO_77 (O_77,N_2536,N_4525);
nand UO_78 (O_78,N_4401,N_4950);
or UO_79 (O_79,N_4940,N_2644);
nand UO_80 (O_80,N_3161,N_4148);
or UO_81 (O_81,N_3555,N_2956);
or UO_82 (O_82,N_3029,N_4727);
or UO_83 (O_83,N_3064,N_3881);
or UO_84 (O_84,N_4150,N_3586);
nor UO_85 (O_85,N_2574,N_3640);
nor UO_86 (O_86,N_3036,N_3254);
nand UO_87 (O_87,N_4608,N_4363);
nor UO_88 (O_88,N_3938,N_3980);
and UO_89 (O_89,N_2907,N_3910);
or UO_90 (O_90,N_3946,N_4359);
or UO_91 (O_91,N_3490,N_4101);
nor UO_92 (O_92,N_3709,N_3062);
nand UO_93 (O_93,N_3055,N_4122);
nor UO_94 (O_94,N_3575,N_2629);
nor UO_95 (O_95,N_4816,N_4159);
or UO_96 (O_96,N_4889,N_3609);
nor UO_97 (O_97,N_3571,N_4893);
or UO_98 (O_98,N_3646,N_3164);
and UO_99 (O_99,N_4081,N_3772);
nor UO_100 (O_100,N_2903,N_2789);
nor UO_101 (O_101,N_4099,N_4992);
nand UO_102 (O_102,N_2870,N_3876);
xnor UO_103 (O_103,N_3972,N_3875);
xnor UO_104 (O_104,N_3583,N_4966);
or UO_105 (O_105,N_4910,N_3468);
nand UO_106 (O_106,N_4662,N_2637);
and UO_107 (O_107,N_2826,N_3904);
nor UO_108 (O_108,N_4779,N_4432);
nor UO_109 (O_109,N_4650,N_3326);
nand UO_110 (O_110,N_4904,N_2689);
or UO_111 (O_111,N_4631,N_3172);
xor UO_112 (O_112,N_2891,N_3761);
nand UO_113 (O_113,N_2636,N_3965);
and UO_114 (O_114,N_3415,N_4614);
nand UO_115 (O_115,N_3722,N_3501);
or UO_116 (O_116,N_4705,N_4858);
nand UO_117 (O_117,N_3653,N_4597);
nor UO_118 (O_118,N_3568,N_4147);
or UO_119 (O_119,N_4223,N_2727);
and UO_120 (O_120,N_4327,N_3027);
nor UO_121 (O_121,N_3451,N_2801);
or UO_122 (O_122,N_3237,N_3457);
nor UO_123 (O_123,N_3970,N_3126);
nand UO_124 (O_124,N_4057,N_3337);
nand UO_125 (O_125,N_4674,N_4815);
and UO_126 (O_126,N_3456,N_3219);
or UO_127 (O_127,N_2944,N_3802);
or UO_128 (O_128,N_4493,N_4418);
and UO_129 (O_129,N_4249,N_3106);
or UO_130 (O_130,N_3417,N_3458);
nand UO_131 (O_131,N_3289,N_3309);
and UO_132 (O_132,N_4257,N_3869);
nand UO_133 (O_133,N_3146,N_4251);
nand UO_134 (O_134,N_4873,N_3669);
or UO_135 (O_135,N_3422,N_2677);
and UO_136 (O_136,N_2571,N_4747);
xnor UO_137 (O_137,N_4741,N_4427);
nand UO_138 (O_138,N_3947,N_4775);
or UO_139 (O_139,N_2947,N_2911);
and UO_140 (O_140,N_2508,N_3162);
and UO_141 (O_141,N_2572,N_4017);
and UO_142 (O_142,N_3079,N_3403);
nand UO_143 (O_143,N_4353,N_4592);
and UO_144 (O_144,N_4431,N_3144);
xor UO_145 (O_145,N_3788,N_2633);
and UO_146 (O_146,N_4137,N_2685);
xnor UO_147 (O_147,N_2994,N_3630);
nor UO_148 (O_148,N_4191,N_4766);
or UO_149 (O_149,N_3205,N_4959);
nor UO_150 (O_150,N_3308,N_4607);
or UO_151 (O_151,N_2893,N_3974);
or UO_152 (O_152,N_3148,N_3203);
and UO_153 (O_153,N_3399,N_4928);
or UO_154 (O_154,N_4316,N_3979);
or UO_155 (O_155,N_4558,N_4804);
nand UO_156 (O_156,N_4465,N_2860);
and UO_157 (O_157,N_3277,N_4051);
and UO_158 (O_158,N_2737,N_2518);
or UO_159 (O_159,N_4045,N_2748);
nand UO_160 (O_160,N_3074,N_4714);
nor UO_161 (O_161,N_2866,N_2898);
nand UO_162 (O_162,N_3338,N_3112);
or UO_163 (O_163,N_2509,N_4925);
or UO_164 (O_164,N_4701,N_3695);
nor UO_165 (O_165,N_3879,N_2762);
nand UO_166 (O_166,N_2981,N_2560);
and UO_167 (O_167,N_3293,N_3836);
nand UO_168 (O_168,N_3660,N_3753);
nor UO_169 (O_169,N_4808,N_3141);
and UO_170 (O_170,N_3091,N_4519);
nor UO_171 (O_171,N_3882,N_4563);
xor UO_172 (O_172,N_4182,N_2720);
nand UO_173 (O_173,N_3957,N_4937);
or UO_174 (O_174,N_4020,N_3523);
nand UO_175 (O_175,N_3533,N_4187);
nand UO_176 (O_176,N_3410,N_3952);
or UO_177 (O_177,N_4520,N_3313);
xnor UO_178 (O_178,N_4027,N_4870);
xor UO_179 (O_179,N_3940,N_3234);
xnor UO_180 (O_180,N_4855,N_3803);
and UO_181 (O_181,N_4377,N_3936);
and UO_182 (O_182,N_3414,N_4121);
or UO_183 (O_183,N_3381,N_3839);
or UO_184 (O_184,N_3143,N_3998);
nand UO_185 (O_185,N_2621,N_4702);
nor UO_186 (O_186,N_4795,N_3748);
and UO_187 (O_187,N_3732,N_3136);
and UO_188 (O_188,N_3636,N_3964);
and UO_189 (O_189,N_4978,N_3220);
or UO_190 (O_190,N_4611,N_3082);
nor UO_191 (O_191,N_2590,N_4312);
or UO_192 (O_192,N_2613,N_2889);
and UO_193 (O_193,N_4688,N_4480);
xnor UO_194 (O_194,N_2589,N_4417);
and UO_195 (O_195,N_2745,N_3877);
and UO_196 (O_196,N_3198,N_4239);
and UO_197 (O_197,N_3513,N_2575);
and UO_198 (O_198,N_4515,N_4192);
or UO_199 (O_199,N_3235,N_2607);
nor UO_200 (O_200,N_2717,N_4939);
nand UO_201 (O_201,N_4037,N_3253);
nand UO_202 (O_202,N_4570,N_3784);
nand UO_203 (O_203,N_3287,N_4508);
and UO_204 (O_204,N_3967,N_3508);
nor UO_205 (O_205,N_3837,N_4504);
nand UO_206 (O_206,N_2824,N_2854);
and UO_207 (O_207,N_3380,N_4550);
and UO_208 (O_208,N_4198,N_2608);
nand UO_209 (O_209,N_4709,N_4758);
or UO_210 (O_210,N_3024,N_4990);
nand UO_211 (O_211,N_2808,N_3482);
nor UO_212 (O_212,N_2946,N_4576);
nand UO_213 (O_213,N_2822,N_2939);
or UO_214 (O_214,N_4656,N_4916);
xor UO_215 (O_215,N_2915,N_3376);
or UO_216 (O_216,N_3231,N_2934);
nor UO_217 (O_217,N_3212,N_4548);
and UO_218 (O_218,N_3576,N_4079);
or UO_219 (O_219,N_3774,N_2960);
nand UO_220 (O_220,N_4529,N_2610);
nor UO_221 (O_221,N_3604,N_3133);
xor UO_222 (O_222,N_2884,N_3888);
or UO_223 (O_223,N_3191,N_2993);
xnor UO_224 (O_224,N_3725,N_4193);
nand UO_225 (O_225,N_4488,N_4810);
and UO_226 (O_226,N_4530,N_4218);
and UO_227 (O_227,N_4593,N_3816);
nor UO_228 (O_228,N_3514,N_4234);
nor UO_229 (O_229,N_2868,N_4993);
and UO_230 (O_230,N_3645,N_3935);
nand UO_231 (O_231,N_4658,N_2549);
nor UO_232 (O_232,N_3778,N_4423);
xnor UO_233 (O_233,N_3297,N_3580);
nor UO_234 (O_234,N_3045,N_4456);
and UO_235 (O_235,N_3923,N_3085);
and UO_236 (O_236,N_3657,N_4664);
or UO_237 (O_237,N_4266,N_4205);
nor UO_238 (O_238,N_4975,N_3007);
or UO_239 (O_239,N_3462,N_4771);
nand UO_240 (O_240,N_3233,N_4385);
nand UO_241 (O_241,N_4219,N_4178);
nor UO_242 (O_242,N_4071,N_4095);
or UO_243 (O_243,N_3620,N_2730);
or UO_244 (O_244,N_3086,N_3274);
nand UO_245 (O_245,N_3763,N_3209);
nor UO_246 (O_246,N_4438,N_3132);
and UO_247 (O_247,N_4435,N_4737);
nand UO_248 (O_248,N_3221,N_3539);
and UO_249 (O_249,N_3632,N_4824);
nand UO_250 (O_250,N_4635,N_4684);
nand UO_251 (O_251,N_4856,N_3515);
nand UO_252 (O_252,N_3049,N_3375);
nor UO_253 (O_253,N_4472,N_2928);
nand UO_254 (O_254,N_3895,N_4466);
nand UO_255 (O_255,N_2517,N_3113);
and UO_256 (O_256,N_4653,N_3003);
or UO_257 (O_257,N_4938,N_4357);
or UO_258 (O_258,N_4666,N_2842);
nand UO_259 (O_259,N_3500,N_2702);
nor UO_260 (O_260,N_4948,N_3638);
nor UO_261 (O_261,N_4370,N_3127);
nand UO_262 (O_262,N_3084,N_3675);
nand UO_263 (O_263,N_3858,N_4536);
nand UO_264 (O_264,N_3723,N_4819);
or UO_265 (O_265,N_4003,N_2527);
or UO_266 (O_266,N_4946,N_3915);
nor UO_267 (O_267,N_2611,N_3118);
nor UO_268 (O_268,N_3928,N_3782);
or UO_269 (O_269,N_3487,N_2501);
or UO_270 (O_270,N_4778,N_3008);
nor UO_271 (O_271,N_3033,N_3087);
and UO_272 (O_272,N_3976,N_3822);
nor UO_273 (O_273,N_3873,N_2859);
nand UO_274 (O_274,N_3081,N_4474);
and UO_275 (O_275,N_4358,N_4102);
nand UO_276 (O_276,N_3443,N_4084);
nand UO_277 (O_277,N_4246,N_2793);
nand UO_278 (O_278,N_3990,N_3749);
and UO_279 (O_279,N_4328,N_4749);
nor UO_280 (O_280,N_4034,N_2559);
nor UO_281 (O_281,N_4588,N_4513);
and UO_282 (O_282,N_3404,N_3269);
and UO_283 (O_283,N_3465,N_4279);
nand UO_284 (O_284,N_3961,N_4203);
and UO_285 (O_285,N_3945,N_3125);
or UO_286 (O_286,N_4183,N_4172);
or UO_287 (O_287,N_3581,N_3529);
nand UO_288 (O_288,N_3032,N_4988);
or UO_289 (O_289,N_2792,N_2863);
nor UO_290 (O_290,N_3090,N_4374);
and UO_291 (O_291,N_4619,N_3827);
or UO_292 (O_292,N_3859,N_4490);
nor UO_293 (O_293,N_4461,N_3264);
nand UO_294 (O_294,N_3322,N_2688);
nor UO_295 (O_295,N_4228,N_2710);
and UO_296 (O_296,N_3861,N_4403);
or UO_297 (O_297,N_4272,N_3018);
and UO_298 (O_298,N_3378,N_4902);
xor UO_299 (O_299,N_4997,N_4391);
or UO_300 (O_300,N_4444,N_4921);
nand UO_301 (O_301,N_4603,N_3181);
nor UO_302 (O_302,N_3846,N_2645);
or UO_303 (O_303,N_4307,N_4752);
and UO_304 (O_304,N_4292,N_3654);
or UO_305 (O_305,N_2563,N_4895);
and UO_306 (O_306,N_4022,N_4072);
nor UO_307 (O_307,N_3053,N_3848);
nor UO_308 (O_308,N_4764,N_3121);
or UO_309 (O_309,N_3232,N_3178);
and UO_310 (O_310,N_3532,N_4894);
and UO_311 (O_311,N_2704,N_3359);
nor UO_312 (O_312,N_3093,N_2502);
xnor UO_313 (O_313,N_2627,N_4163);
or UO_314 (O_314,N_4331,N_4704);
nor UO_315 (O_315,N_4964,N_2926);
or UO_316 (O_316,N_4897,N_4094);
or UO_317 (O_317,N_4606,N_4201);
and UO_318 (O_318,N_3444,N_3809);
and UO_319 (O_319,N_4977,N_4241);
nand UO_320 (O_320,N_4890,N_3336);
and UO_321 (O_321,N_4335,N_2510);
nor UO_322 (O_322,N_4076,N_2634);
nand UO_323 (O_323,N_4923,N_4097);
nor UO_324 (O_324,N_3527,N_4954);
and UO_325 (O_325,N_3275,N_4397);
xnor UO_326 (O_326,N_2558,N_3785);
or UO_327 (O_327,N_4086,N_4100);
or UO_328 (O_328,N_4540,N_2949);
nand UO_329 (O_329,N_2974,N_2665);
and UO_330 (O_330,N_4317,N_2953);
or UO_331 (O_331,N_4278,N_3726);
nand UO_332 (O_332,N_2871,N_3628);
nand UO_333 (O_333,N_2778,N_4282);
or UO_334 (O_334,N_4692,N_2913);
nand UO_335 (O_335,N_2612,N_4533);
nor UO_336 (O_336,N_3613,N_2513);
and UO_337 (O_337,N_4210,N_3467);
or UO_338 (O_338,N_4309,N_4960);
nand UO_339 (O_339,N_3849,N_3993);
nand UO_340 (O_340,N_4837,N_4790);
nand UO_341 (O_341,N_4584,N_2978);
and UO_342 (O_342,N_2855,N_3606);
and UO_343 (O_343,N_4974,N_3907);
xnor UO_344 (O_344,N_4355,N_2882);
nor UO_345 (O_345,N_4445,N_4373);
nor UO_346 (O_346,N_2763,N_3806);
nor UO_347 (O_347,N_4270,N_2967);
or UO_348 (O_348,N_2697,N_2817);
nand UO_349 (O_349,N_4443,N_3582);
or UO_350 (O_350,N_2583,N_2551);
and UO_351 (O_351,N_3637,N_4497);
or UO_352 (O_352,N_3180,N_3329);
xor UO_353 (O_353,N_4792,N_2544);
nand UO_354 (O_354,N_2602,N_4982);
or UO_355 (O_355,N_2721,N_3507);
nor UO_356 (O_356,N_2941,N_3379);
or UO_357 (O_357,N_4545,N_2681);
or UO_358 (O_358,N_4767,N_3599);
nand UO_359 (O_359,N_4012,N_2692);
nor UO_360 (O_360,N_2887,N_3944);
nor UO_361 (O_361,N_4188,N_4769);
nor UO_362 (O_362,N_4750,N_4404);
xor UO_363 (O_363,N_4168,N_3536);
nand UO_364 (O_364,N_4484,N_4609);
nor UO_365 (O_365,N_2711,N_3729);
or UO_366 (O_366,N_3715,N_2682);
and UO_367 (O_367,N_4721,N_2599);
nand UO_368 (O_368,N_4574,N_4481);
xor UO_369 (O_369,N_4615,N_3102);
and UO_370 (O_370,N_3929,N_4787);
nor UO_371 (O_371,N_2528,N_4464);
nor UO_372 (O_372,N_4784,N_3629);
and UO_373 (O_373,N_4526,N_3311);
nand UO_374 (O_374,N_3366,N_3908);
xor UO_375 (O_375,N_3286,N_2862);
or UO_376 (O_376,N_3728,N_3439);
and UO_377 (O_377,N_2795,N_4697);
nand UO_378 (O_378,N_4457,N_2503);
nand UO_379 (O_379,N_4479,N_3706);
xor UO_380 (O_380,N_3543,N_3511);
nor UO_381 (O_381,N_4594,N_2938);
or UO_382 (O_382,N_3663,N_4468);
xnor UO_383 (O_383,N_3190,N_3506);
nor UO_384 (O_384,N_4387,N_3683);
or UO_385 (O_385,N_4332,N_4628);
nor UO_386 (O_386,N_4334,N_4958);
nor UO_387 (O_387,N_2923,N_3095);
or UO_388 (O_388,N_3140,N_4275);
or UO_389 (O_389,N_3271,N_3792);
nand UO_390 (O_390,N_4906,N_3202);
nor UO_391 (O_391,N_4326,N_4612);
and UO_392 (O_392,N_3898,N_4596);
nand UO_393 (O_393,N_2931,N_3996);
nand UO_394 (O_394,N_4586,N_3207);
xor UO_395 (O_395,N_3349,N_4676);
and UO_396 (O_396,N_2740,N_3396);
nor UO_397 (O_397,N_4753,N_3578);
or UO_398 (O_398,N_4802,N_3798);
and UO_399 (O_399,N_4315,N_4565);
or UO_400 (O_400,N_2880,N_4112);
nor UO_401 (O_401,N_4030,N_2714);
and UO_402 (O_402,N_3483,N_4896);
or UO_403 (O_403,N_3259,N_3489);
or UO_404 (O_404,N_3988,N_4277);
nor UO_405 (O_405,N_4759,N_4425);
or UO_406 (O_406,N_4987,N_3165);
xnor UO_407 (O_407,N_3664,N_3222);
nor UO_408 (O_408,N_3931,N_4621);
or UO_409 (O_409,N_3777,N_3612);
and UO_410 (O_410,N_2684,N_4276);
or UO_411 (O_411,N_4681,N_3324);
nor UO_412 (O_412,N_3939,N_3554);
and UO_413 (O_413,N_2875,N_4294);
nand UO_414 (O_414,N_3610,N_3995);
nor UO_415 (O_415,N_3546,N_2617);
nand UO_416 (O_416,N_4259,N_4366);
xor UO_417 (O_417,N_4780,N_4250);
and UO_418 (O_418,N_3335,N_2834);
or UO_419 (O_419,N_2892,N_2883);
nor UO_420 (O_420,N_3246,N_3851);
xnor UO_421 (O_421,N_2819,N_3720);
and UO_422 (O_422,N_3762,N_4669);
nor UO_423 (O_423,N_4673,N_4715);
nor UO_424 (O_424,N_3276,N_2969);
xor UO_425 (O_425,N_4067,N_4695);
and UO_426 (O_426,N_2741,N_3975);
and UO_427 (O_427,N_3953,N_3325);
nor UO_428 (O_428,N_3295,N_2752);
or UO_429 (O_429,N_4065,N_2904);
or UO_430 (O_430,N_4629,N_4013);
xor UO_431 (O_431,N_3649,N_4283);
or UO_432 (O_432,N_2786,N_2615);
nand UO_433 (O_433,N_4587,N_4770);
nor UO_434 (O_434,N_2972,N_3671);
or UO_435 (O_435,N_4381,N_2768);
and UO_436 (O_436,N_2985,N_4862);
and UO_437 (O_437,N_4285,N_3495);
nand UO_438 (O_438,N_2744,N_3054);
nor UO_439 (O_439,N_4175,N_3016);
and UO_440 (O_440,N_2900,N_2917);
and UO_441 (O_441,N_3841,N_3962);
or UO_442 (O_442,N_2918,N_2977);
and UO_443 (O_443,N_2707,N_4248);
nand UO_444 (O_444,N_4165,N_3432);
and UO_445 (O_445,N_4040,N_4299);
and UO_446 (O_446,N_3454,N_2802);
nand UO_447 (O_447,N_4557,N_4826);
xnor UO_448 (O_448,N_2647,N_4722);
and UO_449 (O_449,N_2604,N_3666);
nand UO_450 (O_450,N_2759,N_2995);
or UO_451 (O_451,N_2642,N_2650);
and UO_452 (O_452,N_4630,N_3890);
nor UO_453 (O_453,N_4849,N_3059);
or UO_454 (O_454,N_4124,N_4734);
nor UO_455 (O_455,N_3272,N_2970);
nor UO_456 (O_456,N_3022,N_4793);
and UO_457 (O_457,N_3885,N_3238);
nand UO_458 (O_458,N_3884,N_2691);
or UO_459 (O_459,N_3566,N_4986);
nor UO_460 (O_460,N_3331,N_2516);
xor UO_461 (O_461,N_4679,N_2568);
xnor UO_462 (O_462,N_2800,N_2553);
nor UO_463 (O_463,N_4469,N_2896);
or UO_464 (O_464,N_4340,N_2548);
and UO_465 (O_465,N_3731,N_4642);
or UO_466 (O_466,N_4413,N_4825);
nor UO_467 (O_467,N_4478,N_4598);
or UO_468 (O_468,N_4571,N_4350);
nor UO_469 (O_469,N_4568,N_3052);
and UO_470 (O_470,N_3678,N_4209);
or UO_471 (O_471,N_2631,N_4349);
nor UO_472 (O_472,N_4405,N_4255);
nor UO_473 (O_473,N_4700,N_3364);
nor UO_474 (O_474,N_3201,N_3948);
or UO_475 (O_475,N_4996,N_3355);
nand UO_476 (O_476,N_2648,N_2705);
or UO_477 (O_477,N_3519,N_2971);
nor UO_478 (O_478,N_4410,N_2961);
nand UO_479 (O_479,N_3577,N_3796);
xor UO_480 (O_480,N_3004,N_4195);
and UO_481 (O_481,N_2620,N_4729);
nor UO_482 (O_482,N_3176,N_4196);
nand UO_483 (O_483,N_3579,N_4524);
or UO_484 (O_484,N_3870,N_2690);
and UO_485 (O_485,N_3441,N_2506);
nor UO_486 (O_486,N_4898,N_4117);
xnor UO_487 (O_487,N_3909,N_4516);
or UO_488 (O_488,N_2761,N_4393);
or UO_489 (O_489,N_4724,N_2905);
and UO_490 (O_490,N_2500,N_3983);
and UO_491 (O_491,N_4470,N_3933);
or UO_492 (O_492,N_4634,N_4038);
nand UO_493 (O_493,N_4286,N_3204);
nand UO_494 (O_494,N_4088,N_4177);
nor UO_495 (O_495,N_4610,N_3294);
nor UO_496 (O_496,N_4144,N_2592);
or UO_497 (O_497,N_3832,N_4971);
nand UO_498 (O_498,N_3384,N_4202);
xnor UO_499 (O_499,N_3290,N_3460);
nor UO_500 (O_500,N_3281,N_2990);
or UO_501 (O_501,N_3305,N_4952);
nand UO_502 (O_502,N_2587,N_2818);
nor UO_503 (O_503,N_3367,N_4797);
or UO_504 (O_504,N_2959,N_3548);
xor UO_505 (O_505,N_4738,N_2760);
nand UO_506 (O_506,N_4006,N_3538);
or UO_507 (O_507,N_3900,N_3236);
nand UO_508 (O_508,N_3405,N_4967);
nor UO_509 (O_509,N_3170,N_3789);
and UO_510 (O_510,N_2543,N_3438);
xnor UO_511 (O_511,N_2750,N_3499);
and UO_512 (O_512,N_3020,N_3479);
or UO_513 (O_513,N_4936,N_2666);
and UO_514 (O_514,N_3065,N_4096);
and UO_515 (O_515,N_2878,N_3682);
nand UO_516 (O_516,N_2850,N_3193);
and UO_517 (O_517,N_2683,N_2746);
and UO_518 (O_518,N_2669,N_2872);
nor UO_519 (O_519,N_4092,N_4235);
or UO_520 (O_520,N_3230,N_4798);
nor UO_521 (O_521,N_4932,N_4399);
and UO_522 (O_522,N_4136,N_2708);
nor UO_523 (O_523,N_3502,N_3215);
or UO_524 (O_524,N_3014,N_2529);
and UO_525 (O_525,N_4463,N_3494);
or UO_526 (O_526,N_2897,N_3595);
xnor UO_527 (O_527,N_2521,N_4616);
or UO_528 (O_528,N_2989,N_2739);
nor UO_529 (O_529,N_4746,N_4637);
xnor UO_530 (O_530,N_3484,N_4254);
xnor UO_531 (O_531,N_4760,N_4947);
or UO_532 (O_532,N_4174,N_4229);
nor UO_533 (O_533,N_4221,N_3166);
or UO_534 (O_534,N_3333,N_3185);
and UO_535 (O_535,N_4871,N_4339);
nand UO_536 (O_536,N_3371,N_4569);
nand UO_537 (O_537,N_3710,N_3893);
or UO_538 (O_538,N_3372,N_3061);
or UO_539 (O_539,N_4931,N_4301);
xor UO_540 (O_540,N_4604,N_4929);
xnor UO_541 (O_541,N_3316,N_2925);
nor UO_542 (O_542,N_2832,N_4703);
and UO_543 (O_543,N_2865,N_4049);
xnor UO_544 (O_544,N_4000,N_3089);
and UO_545 (O_545,N_4440,N_2948);
nand UO_546 (O_546,N_3692,N_2921);
nor UO_547 (O_547,N_4212,N_3518);
and UO_548 (O_548,N_2555,N_4560);
or UO_549 (O_549,N_3362,N_2844);
and UO_550 (O_550,N_4728,N_3214);
and UO_551 (O_551,N_4305,N_2606);
nor UO_552 (O_552,N_3863,N_3547);
nand UO_553 (O_553,N_3244,N_4761);
and UO_554 (O_554,N_4252,N_2540);
and UO_555 (O_555,N_2525,N_3889);
and UO_556 (O_556,N_3716,N_2841);
nor UO_557 (O_557,N_2873,N_3797);
nand UO_558 (O_558,N_4510,N_2566);
and UO_559 (O_559,N_3830,N_3056);
and UO_560 (O_560,N_3874,N_3189);
xor UO_561 (O_561,N_4380,N_3680);
or UO_562 (O_562,N_3280,N_2601);
nand UO_563 (O_563,N_4415,N_4115);
and UO_564 (O_564,N_4781,N_4439);
and UO_565 (O_565,N_4909,N_4496);
and UO_566 (O_566,N_3013,N_4878);
or UO_567 (O_567,N_3534,N_2916);
nand UO_568 (O_568,N_4306,N_2794);
or UO_569 (O_569,N_2954,N_3847);
nor UO_570 (O_570,N_2902,N_4337);
and UO_571 (O_571,N_4023,N_2630);
nor UO_572 (O_572,N_2626,N_3843);
and UO_573 (O_573,N_3330,N_3994);
nor UO_574 (O_574,N_2580,N_3044);
and UO_575 (O_575,N_4765,N_4262);
nor UO_576 (O_576,N_3242,N_3662);
and UO_577 (O_577,N_3734,N_4409);
and UO_578 (O_578,N_3174,N_2775);
and UO_579 (O_579,N_4926,N_4919);
or UO_580 (O_580,N_4821,N_4436);
and UO_581 (O_581,N_3696,N_3677);
xor UO_582 (O_582,N_3383,N_4786);
nand UO_583 (O_583,N_3196,N_4073);
nor UO_584 (O_584,N_3751,N_2890);
nor UO_585 (O_585,N_2687,N_3744);
nor UO_586 (O_586,N_3206,N_3622);
or UO_587 (O_587,N_2676,N_4589);
or UO_588 (O_588,N_4053,N_3838);
nor UO_589 (O_589,N_4544,N_4591);
and UO_590 (O_590,N_4846,N_3530);
xnor UO_591 (O_591,N_4400,N_4421);
and UO_592 (O_592,N_4535,N_2686);
nor UO_593 (O_593,N_3340,N_2654);
nor UO_594 (O_594,N_3083,N_3913);
nand UO_595 (O_595,N_3553,N_3169);
nand UO_596 (O_596,N_4141,N_2914);
and UO_597 (O_597,N_4857,N_3155);
nand UO_598 (O_598,N_3918,N_2991);
and UO_599 (O_599,N_3119,N_3466);
or UO_600 (O_600,N_3266,N_2591);
or UO_601 (O_601,N_3063,N_4726);
nor UO_602 (O_602,N_4655,N_3590);
nand UO_603 (O_603,N_2790,N_3999);
nand UO_604 (O_604,N_3868,N_3179);
nor UO_605 (O_605,N_2820,N_4617);
nand UO_606 (O_606,N_4123,N_3634);
nor UO_607 (O_607,N_3051,N_4087);
nand UO_608 (O_608,N_3627,N_4998);
xor UO_609 (O_609,N_3986,N_2950);
nand UO_610 (O_610,N_2523,N_3407);
and UO_611 (O_611,N_4216,N_2738);
and UO_612 (O_612,N_3959,N_3150);
nor UO_613 (O_613,N_3039,N_3592);
and UO_614 (O_614,N_2791,N_4732);
nor UO_615 (O_615,N_4131,N_3824);
or UO_616 (O_616,N_4955,N_3700);
xnor UO_617 (O_617,N_4379,N_3985);
or UO_618 (O_618,N_4980,N_2726);
or UO_619 (O_619,N_2532,N_2699);
nand UO_620 (O_620,N_4859,N_3123);
nor UO_621 (O_621,N_4103,N_2671);
and UO_622 (O_622,N_4371,N_3002);
nand UO_623 (O_623,N_3363,N_3428);
nor UO_624 (O_624,N_3026,N_4803);
nand UO_625 (O_625,N_4031,N_3920);
nor UO_626 (O_626,N_4956,N_4748);
and UO_627 (O_627,N_4712,N_3356);
and UO_628 (O_628,N_3120,N_4302);
or UO_629 (O_629,N_3891,N_3623);
and UO_630 (O_630,N_4194,N_3228);
and UO_631 (O_631,N_4173,N_4880);
or UO_632 (O_632,N_3694,N_2579);
or UO_633 (O_633,N_3815,N_4028);
nor UO_634 (O_634,N_3307,N_3350);
xnor UO_635 (O_635,N_4184,N_2906);
and UO_636 (O_636,N_3122,N_2806);
nor UO_637 (O_637,N_3124,N_3208);
nor UO_638 (O_638,N_4521,N_2680);
or UO_639 (O_639,N_3887,N_4138);
xor UO_640 (O_640,N_3852,N_3252);
nor UO_641 (O_641,N_4200,N_3111);
and UO_642 (O_642,N_4868,N_3758);
nor UO_643 (O_643,N_4145,N_4807);
and UO_644 (O_644,N_4224,N_3665);
or UO_645 (O_645,N_2655,N_4116);
nand UO_646 (O_646,N_4408,N_4927);
nor UO_647 (O_647,N_3302,N_3160);
or UO_648 (O_648,N_4579,N_3319);
and UO_649 (O_649,N_4886,N_3746);
nand UO_650 (O_650,N_3070,N_3411);
nand UO_651 (O_651,N_4429,N_4523);
and UO_652 (O_652,N_3541,N_3615);
xor UO_653 (O_653,N_4344,N_2570);
or UO_654 (O_654,N_3619,N_2951);
nand UO_655 (O_655,N_3435,N_2924);
and UO_656 (O_656,N_2640,N_3702);
or UO_657 (O_657,N_4742,N_2588);
xor UO_658 (O_658,N_3365,N_3315);
nand UO_659 (O_659,N_4128,N_4411);
nand UO_660 (O_660,N_3078,N_3512);
nor UO_661 (O_661,N_3005,N_3941);
nor UO_662 (O_662,N_3129,N_4032);
nor UO_663 (O_663,N_3717,N_3268);
nand UO_664 (O_664,N_3041,N_3429);
nand UO_665 (O_665,N_2764,N_4851);
or UO_666 (O_666,N_4190,N_3000);
xor UO_667 (O_667,N_3223,N_2673);
and UO_668 (O_668,N_4672,N_3200);
nand UO_669 (O_669,N_3047,N_3332);
nor UO_670 (O_670,N_3473,N_3624);
nor UO_671 (O_671,N_4338,N_4052);
or UO_672 (O_672,N_3387,N_4501);
and UO_673 (O_673,N_3562,N_3471);
or UO_674 (O_674,N_4696,N_3616);
nor UO_675 (O_675,N_4333,N_2825);
and UO_676 (O_676,N_4541,N_4624);
nand UO_677 (O_677,N_4866,N_2609);
nor UO_678 (O_678,N_3245,N_4109);
xnor UO_679 (O_679,N_3919,N_2675);
xor UO_680 (O_680,N_2732,N_4170);
xor UO_681 (O_681,N_2874,N_3737);
or UO_682 (O_682,N_4452,N_3603);
or UO_683 (O_683,N_2962,N_4066);
or UO_684 (O_684,N_3672,N_4716);
and UO_685 (O_685,N_2821,N_3420);
nand UO_686 (O_686,N_3794,N_3707);
and UO_687 (O_687,N_2933,N_2881);
and UO_688 (O_688,N_4323,N_3862);
nor UO_689 (O_689,N_2940,N_4503);
nand UO_690 (O_690,N_3299,N_4204);
nor UO_691 (O_691,N_4222,N_4693);
or UO_692 (O_692,N_2576,N_4450);
nand UO_693 (O_693,N_4830,N_3896);
xnor UO_694 (O_694,N_2996,N_3727);
and UO_695 (O_695,N_2766,N_3775);
or UO_696 (O_696,N_3989,N_3810);
nor UO_697 (O_697,N_4626,N_4646);
and UO_698 (O_698,N_3470,N_3821);
nand UO_699 (O_699,N_4442,N_4590);
nand UO_700 (O_700,N_3828,N_4911);
or UO_701 (O_701,N_3130,N_4437);
and UO_702 (O_702,N_2838,N_3413);
and UO_703 (O_703,N_4308,N_3845);
nor UO_704 (O_704,N_3854,N_4402);
nor UO_705 (O_705,N_3283,N_4290);
and UO_706 (O_706,N_3273,N_3602);
nand UO_707 (O_707,N_3304,N_4133);
or UO_708 (O_708,N_4552,N_4459);
and UO_709 (O_709,N_3469,N_2958);
or UO_710 (O_710,N_3416,N_4321);
and UO_711 (O_711,N_3030,N_4645);
nand UO_712 (O_712,N_4685,N_3157);
nand UO_713 (O_713,N_2830,N_4976);
or UO_714 (O_714,N_3525,N_2678);
and UO_715 (O_715,N_4061,N_3912);
nand UO_716 (O_716,N_3795,N_3425);
and UO_717 (O_717,N_2813,N_3625);
nand UO_718 (O_718,N_3255,N_4509);
nand UO_719 (O_719,N_3104,N_4818);
xor UO_720 (O_720,N_2853,N_3676);
nand UO_721 (O_721,N_4018,N_2552);
and UO_722 (O_722,N_4318,N_4517);
nor UO_723 (O_723,N_4021,N_4324);
xor UO_724 (O_724,N_3835,N_3486);
nor UO_725 (O_725,N_2781,N_4245);
and UO_726 (O_726,N_3618,N_4458);
nor UO_727 (O_727,N_2803,N_3872);
nand UO_728 (O_728,N_3377,N_4026);
and UO_729 (O_729,N_3524,N_3496);
and UO_730 (O_730,N_4118,N_2584);
and UO_731 (O_731,N_4300,N_3447);
and UO_732 (O_732,N_4199,N_4367);
nor UO_733 (O_733,N_2899,N_4157);
or UO_734 (O_734,N_4325,N_3043);
or UO_735 (O_735,N_3973,N_2827);
nand UO_736 (O_736,N_3840,N_3485);
or UO_737 (O_737,N_3969,N_4813);
and UO_738 (O_738,N_4056,N_3551);
and UO_739 (O_739,N_4014,N_4089);
nand UO_740 (O_740,N_3768,N_2639);
nor UO_741 (O_741,N_4448,N_3225);
nor UO_742 (O_742,N_3037,N_4651);
nor UO_743 (O_743,N_4206,N_3427);
nor UO_744 (O_744,N_2742,N_3880);
and UO_745 (O_745,N_4689,N_3424);
or UO_746 (O_746,N_2798,N_4449);
or UO_747 (O_747,N_2983,N_2534);
or UO_748 (O_748,N_3564,N_4042);
and UO_749 (O_749,N_4812,N_4098);
or UO_750 (O_750,N_3072,N_4382);
or UO_751 (O_751,N_4130,N_2829);
and UO_752 (O_752,N_4207,N_4146);
nand UO_753 (O_753,N_3192,N_4236);
nand UO_754 (O_754,N_2733,N_4110);
nand UO_755 (O_755,N_4369,N_4063);
or UO_756 (O_756,N_4762,N_3504);
nor UO_757 (O_757,N_3134,N_2846);
nor UO_758 (O_758,N_4476,N_3459);
nor UO_759 (O_759,N_4407,N_4330);
nor UO_760 (O_760,N_4789,N_3023);
nor UO_761 (O_761,N_3341,N_3241);
or UO_762 (O_762,N_3151,N_2888);
xnor UO_763 (O_763,N_3914,N_3323);
and UO_764 (O_764,N_3464,N_4477);
nor UO_765 (O_765,N_3901,N_2538);
and UO_766 (O_766,N_3864,N_3698);
nand UO_767 (O_767,N_4211,N_3926);
or UO_768 (O_768,N_4396,N_3248);
and UO_769 (O_769,N_4531,N_3559);
or UO_770 (O_770,N_2943,N_2505);
or UO_771 (O_771,N_2625,N_2799);
and UO_772 (O_772,N_4774,N_4961);
and UO_773 (O_773,N_2784,N_3463);
or UO_774 (O_774,N_4454,N_4263);
nor UO_775 (O_775,N_2614,N_3048);
nor UO_776 (O_776,N_4368,N_3288);
nor UO_777 (O_777,N_2894,N_4281);
nor UO_778 (O_778,N_3942,N_3171);
nand UO_779 (O_779,N_4329,N_2716);
or UO_780 (O_780,N_3398,N_4238);
xnor UO_781 (O_781,N_3927,N_3757);
nor UO_782 (O_782,N_3034,N_4313);
xnor UO_783 (O_783,N_3450,N_2703);
or UO_784 (O_784,N_2533,N_3137);
or UO_785 (O_785,N_4107,N_2596);
and UO_786 (O_786,N_2782,N_3184);
nand UO_787 (O_787,N_3477,N_2652);
nor UO_788 (O_788,N_3594,N_3905);
nor UO_789 (O_789,N_3668,N_3135);
nor UO_790 (O_790,N_4743,N_4599);
or UO_791 (O_791,N_4618,N_4572);
nor UO_792 (O_792,N_2908,N_3567);
or UO_793 (O_793,N_4075,N_2770);
nand UO_794 (O_794,N_2656,N_3721);
nor UO_795 (O_795,N_3684,N_4085);
and UO_796 (O_796,N_2837,N_2849);
nand UO_797 (O_797,N_4639,N_4884);
or UO_798 (O_798,N_4395,N_2679);
and UO_799 (O_799,N_3565,N_2557);
and UO_800 (O_800,N_4120,N_2812);
and UO_801 (O_801,N_4149,N_3589);
nor UO_802 (O_802,N_2725,N_3046);
or UO_803 (O_803,N_2930,N_3094);
nor UO_804 (O_804,N_3394,N_4744);
nand UO_805 (O_805,N_4105,N_4930);
and UO_806 (O_806,N_3658,N_4941);
and UO_807 (O_807,N_2701,N_4867);
nand UO_808 (O_808,N_2999,N_3773);
and UO_809 (O_809,N_3431,N_3535);
nor UO_810 (O_810,N_4372,N_3310);
nor UO_811 (O_811,N_2582,N_3239);
and UO_812 (O_812,N_4708,N_2585);
nand UO_813 (O_813,N_4273,N_4360);
or UO_814 (O_814,N_2963,N_2594);
and UO_815 (O_815,N_2698,N_4505);
nand UO_816 (O_816,N_3611,N_3736);
nand UO_817 (O_817,N_3418,N_4773);
nor UO_818 (O_818,N_2845,N_4796);
or UO_819 (O_819,N_4872,N_3038);
nor UO_820 (O_820,N_2852,N_3517);
and UO_821 (O_821,N_4577,N_4047);
nand UO_822 (O_822,N_4422,N_3673);
and UO_823 (O_823,N_3739,N_3436);
xor UO_824 (O_824,N_3865,N_3210);
and UO_825 (O_825,N_4573,N_2561);
nor UO_826 (O_826,N_4643,N_4035);
nor UO_827 (O_827,N_3871,N_4487);
and UO_828 (O_828,N_4719,N_4033);
nor UO_829 (O_829,N_4295,N_3303);
nor UO_830 (O_830,N_2661,N_3270);
or UO_831 (O_831,N_2955,N_4944);
and UO_832 (O_832,N_2927,N_3674);
nor UO_833 (O_833,N_3117,N_3569);
and UO_834 (O_834,N_4581,N_2857);
xnor UO_835 (O_835,N_3250,N_4426);
or UO_836 (O_836,N_3218,N_4134);
xnor UO_837 (O_837,N_3224,N_3651);
nand UO_838 (O_838,N_4671,N_4667);
or UO_839 (O_839,N_4414,N_4311);
nand UO_840 (O_840,N_3449,N_3899);
and UO_841 (O_841,N_3291,N_4682);
and UO_842 (O_842,N_4768,N_3258);
or UO_843 (O_843,N_3659,N_3783);
nand UO_844 (O_844,N_4046,N_4915);
or UO_845 (O_845,N_3714,N_3491);
or UO_846 (O_846,N_3388,N_4111);
and UO_847 (O_847,N_3621,N_4864);
xor UO_848 (O_848,N_3261,N_3100);
nor UO_849 (O_849,N_3092,N_3542);
or UO_850 (O_850,N_3516,N_3968);
nand UO_851 (O_851,N_4832,N_2757);
and UO_852 (O_852,N_3760,N_4660);
nor UO_853 (O_853,N_4957,N_4420);
and UO_854 (O_854,N_3661,N_3818);
nand UO_855 (O_855,N_4788,N_4126);
and UO_856 (O_856,N_4253,N_4546);
and UO_857 (O_857,N_4828,N_4419);
nand UO_858 (O_858,N_2728,N_3114);
and UO_859 (O_859,N_4725,N_4008);
nor UO_860 (O_860,N_2641,N_4140);
or UO_861 (O_861,N_4723,N_2519);
or UO_862 (O_862,N_2734,N_4514);
xor UO_863 (O_863,N_4949,N_3679);
nand UO_864 (O_864,N_3296,N_2514);
nor UO_865 (O_865,N_3770,N_4561);
xnor UO_866 (O_866,N_3591,N_4822);
nor UO_867 (O_867,N_2937,N_3334);
nand UO_868 (O_868,N_2651,N_2593);
or UO_869 (O_869,N_4154,N_3747);
nor UO_870 (O_870,N_4686,N_3991);
and UO_871 (O_871,N_3455,N_3573);
nor UO_872 (O_872,N_3312,N_3409);
nand UO_873 (O_873,N_2876,N_4657);
and UO_874 (O_874,N_4215,N_2788);
nand UO_875 (O_875,N_2597,N_3598);
or UO_876 (O_876,N_4917,N_3560);
or UO_877 (O_877,N_2772,N_2504);
nand UO_878 (O_878,N_4580,N_4838);
or UO_879 (O_879,N_4888,N_3080);
nand UO_880 (O_880,N_4455,N_3397);
nor UO_881 (O_881,N_2556,N_3930);
or UO_882 (O_882,N_4829,N_3099);
nand UO_883 (O_883,N_3558,N_3826);
nand UO_884 (O_884,N_4060,N_4865);
nand UO_885 (O_885,N_3361,N_3878);
or UO_886 (O_886,N_3883,N_3855);
and UO_887 (O_887,N_4735,N_3886);
nand UO_888 (O_888,N_3790,N_2932);
or UO_889 (O_889,N_3742,N_2758);
nand UO_890 (O_890,N_3596,N_2709);
xor UO_891 (O_891,N_3787,N_4161);
and UO_892 (O_892,N_2987,N_4267);
nand UO_893 (O_893,N_3856,N_3138);
nand UO_894 (O_894,N_4489,N_4984);
nor UO_895 (O_895,N_4836,N_4189);
and UO_896 (O_896,N_4763,N_2522);
nand UO_897 (O_897,N_2550,N_3195);
nor UO_898 (O_898,N_3346,N_4091);
nand UO_899 (O_899,N_4843,N_2628);
xnor UO_900 (O_900,N_2848,N_4962);
and UO_901 (O_901,N_2724,N_4055);
or UO_902 (O_902,N_2851,N_4740);
nand UO_903 (O_903,N_2624,N_2535);
nand UO_904 (O_904,N_4717,N_3544);
or UO_905 (O_905,N_3738,N_4074);
and UO_906 (O_906,N_4549,N_2771);
or UO_907 (O_907,N_2618,N_3992);
nand UO_908 (O_908,N_4756,N_4892);
nand UO_909 (O_909,N_3186,N_3650);
or UO_910 (O_910,N_3814,N_2695);
nand UO_911 (O_911,N_2753,N_4291);
and UO_912 (O_912,N_4424,N_2520);
nor UO_913 (O_913,N_3042,N_2805);
xor UO_914 (O_914,N_3492,N_4258);
nand UO_915 (O_915,N_3475,N_4142);
nand UO_916 (O_916,N_4048,N_2957);
or UO_917 (O_917,N_4498,N_3767);
or UO_918 (O_918,N_3520,N_4914);
and UO_919 (O_919,N_2836,N_3173);
nor UO_920 (O_920,N_4288,N_4127);
or UO_921 (O_921,N_4839,N_3067);
and UO_922 (O_922,N_3556,N_4451);
nand UO_923 (O_923,N_4876,N_4462);
nand UO_924 (O_924,N_3954,N_4652);
and UO_925 (O_925,N_2658,N_2810);
nand UO_926 (O_926,N_2936,N_2619);
nand UO_927 (O_927,N_4554,N_3897);
nand UO_928 (O_928,N_4217,N_3101);
and UO_929 (O_929,N_4847,N_3385);
xnor UO_930 (O_930,N_3373,N_2700);
or UO_931 (O_931,N_4649,N_3531);
nand UO_932 (O_932,N_2886,N_4891);
and UO_933 (O_933,N_2646,N_3647);
nand UO_934 (O_934,N_4935,N_3754);
xor UO_935 (O_935,N_3440,N_4361);
nor UO_936 (O_936,N_4640,N_4225);
and UO_937 (O_937,N_2562,N_3648);
nor UO_938 (O_938,N_4644,N_2595);
nand UO_939 (O_939,N_3687,N_4156);
or UO_940 (O_940,N_3693,N_2659);
nor UO_941 (O_941,N_4208,N_4230);
nor UO_942 (O_942,N_3057,N_4885);
and UO_943 (O_943,N_3386,N_4600);
or UO_944 (O_944,N_2997,N_4665);
xnor UO_945 (O_945,N_3493,N_4794);
nor UO_946 (O_946,N_3358,N_3510);
nor UO_947 (O_947,N_2975,N_3949);
nand UO_948 (O_948,N_4882,N_2581);
or UO_949 (O_949,N_4113,N_2796);
or UO_950 (O_950,N_3035,N_3412);
nand UO_951 (O_951,N_4434,N_4730);
or UO_952 (O_952,N_4256,N_2546);
nor UO_953 (O_953,N_4687,N_3766);
or UO_954 (O_954,N_4706,N_3759);
and UO_955 (O_955,N_4483,N_2530);
and UO_956 (O_956,N_4559,N_3811);
nand UO_957 (O_957,N_4680,N_4543);
or UO_958 (O_958,N_3368,N_3701);
or UO_959 (O_959,N_3262,N_3408);
nand UO_960 (O_960,N_3892,N_3145);
nand UO_961 (O_961,N_3712,N_3488);
nand UO_962 (O_962,N_4578,N_3561);
nor UO_963 (O_963,N_3474,N_4920);
and UO_964 (O_964,N_4467,N_2569);
nor UO_965 (O_965,N_3478,N_4677);
nor UO_966 (O_966,N_2973,N_3860);
nand UO_967 (O_967,N_3391,N_4632);
xnor UO_968 (O_968,N_4388,N_4678);
or UO_969 (O_969,N_4736,N_3393);
xor UO_970 (O_970,N_4082,N_3823);
and UO_971 (O_971,N_4289,N_3552);
nand UO_972 (O_972,N_4899,N_2747);
and UO_973 (O_973,N_4416,N_3635);
or UO_974 (O_974,N_4973,N_4231);
or UO_975 (O_975,N_4601,N_3528);
nand UO_976 (O_976,N_3922,N_4636);
or UO_977 (O_977,N_3756,N_2982);
nand UO_978 (O_978,N_2984,N_3448);
and UO_979 (O_979,N_4005,N_4319);
nand UO_980 (O_980,N_4024,N_2616);
nand UO_981 (O_981,N_4293,N_2776);
and UO_982 (O_982,N_4817,N_4226);
nor UO_983 (O_983,N_3685,N_4166);
nor UO_984 (O_984,N_4633,N_4167);
nand UO_985 (O_985,N_3107,N_4176);
and UO_986 (O_986,N_2935,N_2831);
xor UO_987 (O_987,N_4691,N_3292);
nand UO_988 (O_988,N_4029,N_3040);
and UO_989 (O_989,N_3689,N_4482);
xor UO_990 (O_990,N_3402,N_2864);
nand UO_991 (O_991,N_4875,N_4375);
nor UO_992 (O_992,N_4991,N_3667);
and UO_993 (O_993,N_2696,N_4213);
nor UO_994 (O_994,N_3461,N_2729);
or UO_995 (O_995,N_3382,N_2749);
nand UO_996 (O_996,N_3400,N_4782);
nor UO_997 (O_997,N_3699,N_4011);
nor UO_998 (O_998,N_4908,N_3110);
nand UO_999 (O_999,N_4777,N_3801);
endmodule