module basic_2000_20000_2500_125_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
nand U0 (N_0,In_515,In_232);
nand U1 (N_1,In_1323,In_1186);
xnor U2 (N_2,In_1355,In_859);
xnor U3 (N_3,In_730,In_425);
xnor U4 (N_4,In_1661,In_694);
or U5 (N_5,In_581,In_1689);
nor U6 (N_6,In_907,In_982);
and U7 (N_7,In_672,In_1195);
nor U8 (N_8,In_605,In_1966);
and U9 (N_9,In_1053,In_1573);
nand U10 (N_10,In_973,In_1506);
nand U11 (N_11,In_1578,In_1990);
or U12 (N_12,In_870,In_1556);
and U13 (N_13,In_1308,In_1534);
and U14 (N_14,In_229,In_616);
nor U15 (N_15,In_849,In_1244);
or U16 (N_16,In_501,In_1895);
xor U17 (N_17,In_540,In_1223);
and U18 (N_18,In_562,In_1013);
or U19 (N_19,In_794,In_144);
xnor U20 (N_20,In_202,In_134);
nor U21 (N_21,In_594,In_436);
and U22 (N_22,In_1154,In_758);
nand U23 (N_23,In_409,In_1944);
and U24 (N_24,In_1294,In_847);
and U25 (N_25,In_856,In_27);
or U26 (N_26,In_1466,In_863);
and U27 (N_27,In_1872,In_102);
nor U28 (N_28,In_572,In_897);
or U29 (N_29,In_1645,In_11);
xnor U30 (N_30,In_206,In_323);
xor U31 (N_31,In_159,In_807);
or U32 (N_32,In_80,In_1394);
and U33 (N_33,In_1473,In_1911);
xnor U34 (N_34,In_1765,In_1601);
nand U35 (N_35,In_840,In_377);
xor U36 (N_36,In_753,In_1399);
nand U37 (N_37,In_125,In_135);
and U38 (N_38,In_435,In_661);
xor U39 (N_39,In_68,In_1107);
or U40 (N_40,In_1433,In_61);
xor U41 (N_41,In_189,In_1015);
or U42 (N_42,In_218,In_1258);
or U43 (N_43,In_846,In_398);
xor U44 (N_44,In_1742,In_404);
and U45 (N_45,In_1286,In_440);
nor U46 (N_46,In_414,In_615);
xor U47 (N_47,In_604,In_1364);
or U48 (N_48,In_1167,In_1896);
xnor U49 (N_49,In_529,In_983);
nand U50 (N_50,In_32,In_1315);
or U51 (N_51,In_410,In_1325);
and U52 (N_52,In_785,In_8);
or U53 (N_53,In_1986,In_1347);
xnor U54 (N_54,In_1392,In_1362);
and U55 (N_55,In_1881,In_1090);
xor U56 (N_56,In_561,In_344);
and U57 (N_57,In_1117,In_1659);
or U58 (N_58,In_1611,In_1733);
nor U59 (N_59,In_340,In_1841);
xor U60 (N_60,In_691,In_1828);
or U61 (N_61,In_76,In_1310);
nor U62 (N_62,In_1129,In_1031);
xor U63 (N_63,In_1997,In_1288);
or U64 (N_64,In_486,In_1257);
nand U65 (N_65,In_654,In_383);
nand U66 (N_66,In_1920,In_993);
nand U67 (N_67,In_838,In_1837);
or U68 (N_68,In_136,In_1151);
nand U69 (N_69,In_50,In_1800);
or U70 (N_70,In_1089,In_402);
nor U71 (N_71,In_1538,In_545);
xnor U72 (N_72,In_1839,In_1835);
nor U73 (N_73,In_348,In_213);
and U74 (N_74,In_1946,In_362);
and U75 (N_75,In_1823,In_1813);
nor U76 (N_76,In_505,In_1735);
or U77 (N_77,In_1239,In_818);
and U78 (N_78,In_667,In_595);
nor U79 (N_79,In_1351,In_685);
or U80 (N_80,In_1846,In_1383);
or U81 (N_81,In_1280,In_551);
nand U82 (N_82,In_502,In_156);
xor U83 (N_83,In_1577,In_857);
nor U84 (N_84,In_795,In_1642);
or U85 (N_85,In_1822,In_1328);
and U86 (N_86,In_231,In_1220);
nor U87 (N_87,In_1023,In_895);
nand U88 (N_88,In_861,In_368);
nor U89 (N_89,In_220,In_416);
and U90 (N_90,In_291,In_1728);
and U91 (N_91,In_1268,In_560);
nand U92 (N_92,In_1868,In_1134);
xor U93 (N_93,In_511,In_602);
and U94 (N_94,In_728,In_592);
nand U95 (N_95,In_179,In_1546);
or U96 (N_96,In_1348,In_279);
and U97 (N_97,In_3,In_89);
and U98 (N_98,In_428,In_471);
xor U99 (N_99,In_1853,In_523);
xnor U100 (N_100,In_166,In_723);
nor U101 (N_101,In_482,In_152);
xnor U102 (N_102,In_632,In_272);
or U103 (N_103,In_1201,In_656);
and U104 (N_104,In_1003,In_1641);
or U105 (N_105,In_1575,In_1713);
or U106 (N_106,In_1729,In_1811);
and U107 (N_107,In_1775,In_939);
or U108 (N_108,In_1673,In_1247);
xor U109 (N_109,In_673,In_874);
nor U110 (N_110,In_1361,In_1617);
nor U111 (N_111,In_621,In_934);
nor U112 (N_112,In_1806,In_1378);
nand U113 (N_113,In_210,In_328);
or U114 (N_114,In_1763,In_1740);
xor U115 (N_115,In_70,In_1372);
nand U116 (N_116,In_254,In_1629);
xor U117 (N_117,In_1767,In_381);
or U118 (N_118,In_677,In_1588);
xor U119 (N_119,In_974,In_1598);
xor U120 (N_120,In_1382,In_520);
nor U121 (N_121,In_652,In_1357);
xor U122 (N_122,In_1236,In_205);
or U123 (N_123,In_451,In_885);
or U124 (N_124,In_1530,In_784);
or U125 (N_125,In_651,In_40);
nand U126 (N_126,In_536,In_603);
xnor U127 (N_127,In_868,In_1485);
and U128 (N_128,In_106,In_413);
nor U129 (N_129,In_1798,In_269);
and U130 (N_130,In_1254,In_1663);
or U131 (N_131,In_777,In_1679);
xnor U132 (N_132,In_1861,In_1829);
xor U133 (N_133,In_1396,In_437);
nor U134 (N_134,In_1698,In_1381);
or U135 (N_135,In_1252,In_330);
xnor U136 (N_136,In_763,In_1675);
nand U137 (N_137,In_1709,In_608);
or U138 (N_138,In_949,In_53);
nor U139 (N_139,In_1924,In_493);
nor U140 (N_140,In_1519,In_16);
nand U141 (N_141,In_1316,In_812);
or U142 (N_142,In_717,In_732);
and U143 (N_143,In_107,In_1904);
xnor U144 (N_144,In_1340,In_1736);
nand U145 (N_145,In_1754,In_1799);
and U146 (N_146,In_312,In_1739);
nand U147 (N_147,In_832,In_517);
nor U148 (N_148,In_1513,In_1307);
nor U149 (N_149,In_792,In_1342);
xor U150 (N_150,In_1533,In_464);
and U151 (N_151,In_1836,In_1779);
or U152 (N_152,In_56,In_1052);
or U153 (N_153,In_1523,In_507);
nor U154 (N_154,In_375,In_252);
or U155 (N_155,In_1241,In_1177);
xnor U156 (N_156,In_1464,In_681);
or U157 (N_157,In_975,In_1501);
xnor U158 (N_158,In_1259,In_802);
nor U159 (N_159,In_343,In_1613);
or U160 (N_160,In_1769,In_187);
nand U161 (N_161,In_990,In_1934);
or U162 (N_162,In_1414,In_1237);
nor U163 (N_163,In_678,In_193);
nor U164 (N_164,In_565,In_1737);
or U165 (N_165,In_1520,In_913);
nand U166 (N_166,In_1266,N_106);
nand U167 (N_167,In_1522,In_1845);
or U168 (N_168,In_467,In_1141);
or U169 (N_169,In_825,In_1084);
and U170 (N_170,In_1616,In_44);
and U171 (N_171,In_492,In_1424);
and U172 (N_172,In_1517,In_514);
and U173 (N_173,In_1745,In_359);
or U174 (N_174,In_1043,In_242);
or U175 (N_175,N_30,In_1336);
xnor U176 (N_176,In_1370,N_93);
nand U177 (N_177,In_1283,In_1889);
nand U178 (N_178,In_755,In_979);
xnor U179 (N_179,In_313,In_542);
and U180 (N_180,In_995,In_688);
nor U181 (N_181,In_1373,In_1599);
xnor U182 (N_182,In_237,In_1181);
xnor U183 (N_183,N_70,In_1435);
xnor U184 (N_184,In_162,In_1486);
or U185 (N_185,In_1918,N_129);
nor U186 (N_186,In_347,In_1233);
nand U187 (N_187,In_790,In_1393);
or U188 (N_188,In_587,In_1993);
nor U189 (N_189,In_441,In_88);
nand U190 (N_190,In_947,N_115);
or U191 (N_191,In_966,In_1048);
nor U192 (N_192,In_1834,In_1312);
nand U193 (N_193,In_1019,In_1029);
and U194 (N_194,In_1744,In_124);
and U195 (N_195,In_662,In_558);
xnor U196 (N_196,N_2,In_532);
xnor U197 (N_197,In_1388,In_1009);
or U198 (N_198,N_68,In_1772);
nand U199 (N_199,In_1144,In_816);
nand U200 (N_200,In_1873,In_251);
or U201 (N_201,In_1380,In_1858);
or U202 (N_202,N_86,In_97);
nor U203 (N_203,In_1278,N_17);
and U204 (N_204,In_1768,In_1262);
nor U205 (N_205,In_851,In_260);
and U206 (N_206,In_637,In_1438);
nor U207 (N_207,In_619,In_692);
nor U208 (N_208,In_423,In_1625);
and U209 (N_209,In_512,In_1985);
nor U210 (N_210,In_130,In_165);
or U211 (N_211,In_376,In_760);
nand U212 (N_212,In_133,In_1717);
nand U213 (N_213,In_396,In_1002);
and U214 (N_214,In_1874,In_697);
and U215 (N_215,In_268,In_235);
and U216 (N_216,In_58,In_1660);
xnor U217 (N_217,In_199,In_890);
and U218 (N_218,N_26,In_1113);
or U219 (N_219,In_1421,In_972);
nand U220 (N_220,In_568,In_439);
or U221 (N_221,In_420,In_1569);
or U222 (N_222,In_964,In_828);
nand U223 (N_223,N_114,In_71);
and U224 (N_224,In_1630,In_1665);
nor U225 (N_225,In_1825,In_1752);
nor U226 (N_226,N_139,In_1657);
or U227 (N_227,In_498,In_483);
or U228 (N_228,In_894,In_1069);
xnor U229 (N_229,In_690,In_1564);
or U230 (N_230,In_99,N_117);
nor U231 (N_231,In_48,In_20);
or U232 (N_232,In_1008,In_1260);
or U233 (N_233,In_278,In_683);
xor U234 (N_234,In_249,In_1809);
and U235 (N_235,In_223,In_702);
or U236 (N_236,N_24,In_841);
xnor U237 (N_237,In_294,In_1844);
xnor U238 (N_238,N_88,In_765);
nand U239 (N_239,In_487,In_174);
or U240 (N_240,In_1275,In_1116);
nand U241 (N_241,In_324,In_1509);
nand U242 (N_242,In_447,In_1781);
nand U243 (N_243,In_920,In_1391);
or U244 (N_244,In_41,In_1408);
and U245 (N_245,In_1389,In_742);
nand U246 (N_246,In_570,In_1916);
and U247 (N_247,In_1593,In_1410);
or U248 (N_248,In_1995,In_1851);
and U249 (N_249,In_622,In_17);
xnor U250 (N_250,In_518,N_84);
xor U251 (N_251,In_837,In_746);
or U252 (N_252,In_1969,In_1138);
or U253 (N_253,In_1855,N_96);
and U254 (N_254,In_1727,In_1771);
nand U255 (N_255,N_138,In_1610);
or U256 (N_256,In_1819,In_1687);
nand U257 (N_257,In_1796,In_1367);
or U258 (N_258,In_1927,In_1037);
nand U259 (N_259,In_712,In_450);
xnor U260 (N_260,In_298,In_877);
and U261 (N_261,In_1234,In_1576);
xor U262 (N_262,In_1132,In_1815);
nor U263 (N_263,In_941,In_1743);
and U264 (N_264,In_642,In_118);
nor U265 (N_265,In_1021,In_1992);
or U266 (N_266,In_1489,In_829);
and U267 (N_267,In_564,N_94);
and U268 (N_268,In_1640,In_1301);
nand U269 (N_269,In_1544,In_567);
nor U270 (N_270,In_687,In_1704);
xnor U271 (N_271,In_1719,In_1476);
and U272 (N_272,In_1417,In_1016);
nand U273 (N_273,In_554,In_1165);
nand U274 (N_274,In_1792,In_142);
nor U275 (N_275,In_817,In_761);
or U276 (N_276,In_121,In_1535);
or U277 (N_277,In_1297,In_1725);
or U278 (N_278,N_156,In_468);
nand U279 (N_279,In_1386,In_1602);
or U280 (N_280,In_1959,In_109);
nor U281 (N_281,In_918,In_117);
xnor U282 (N_282,N_41,In_1963);
and U283 (N_283,In_1991,In_1354);
or U284 (N_284,In_1160,In_1216);
nand U285 (N_285,In_304,In_6);
nor U286 (N_286,In_748,In_475);
nor U287 (N_287,In_844,In_1860);
or U288 (N_288,In_609,In_1179);
xnor U289 (N_289,In_1095,In_591);
xnor U290 (N_290,In_1202,In_1017);
nor U291 (N_291,N_59,In_886);
nor U292 (N_292,In_1453,In_1912);
nor U293 (N_293,In_1962,In_28);
nand U294 (N_294,N_73,In_705);
nand U295 (N_295,In_1831,In_393);
nor U296 (N_296,In_1108,In_1537);
nor U297 (N_297,In_1060,In_1528);
or U298 (N_298,In_1333,In_1757);
nor U299 (N_299,N_8,In_356);
and U300 (N_300,In_1490,In_1353);
or U301 (N_301,In_224,In_9);
and U302 (N_302,In_1667,In_1941);
and U303 (N_303,In_1859,In_752);
xnor U304 (N_304,In_1209,In_415);
xor U305 (N_305,In_1203,In_354);
and U306 (N_306,In_700,In_1931);
or U307 (N_307,In_850,In_1526);
xnor U308 (N_308,In_341,N_20);
or U309 (N_309,In_1812,In_528);
or U310 (N_310,In_1748,In_49);
nor U311 (N_311,In_819,In_198);
and U312 (N_312,In_1020,In_45);
xor U313 (N_313,In_30,In_1892);
xnor U314 (N_314,In_1979,In_31);
and U315 (N_315,In_1746,N_90);
nand U316 (N_316,In_1804,In_1279);
xnor U317 (N_317,In_855,In_1552);
nor U318 (N_318,N_110,In_927);
and U319 (N_319,In_1913,In_1906);
and U320 (N_320,In_525,In_1035);
and U321 (N_321,In_127,In_876);
nor U322 (N_322,In_452,In_146);
xnor U323 (N_323,In_801,In_984);
nor U324 (N_324,In_1334,In_896);
or U325 (N_325,In_1405,In_1605);
and U326 (N_326,In_1933,In_353);
nand U327 (N_327,In_333,In_1567);
and U328 (N_328,In_317,N_150);
or U329 (N_329,In_1558,In_137);
nor U330 (N_330,In_1720,In_39);
nand U331 (N_331,In_1402,In_971);
or U332 (N_332,In_1448,N_233);
nor U333 (N_333,In_209,N_183);
or U334 (N_334,In_1885,In_1936);
and U335 (N_335,In_780,In_1762);
or U336 (N_336,In_860,In_1432);
nand U337 (N_337,In_29,In_620);
nand U338 (N_338,In_881,In_981);
or U339 (N_339,In_960,In_1193);
nor U340 (N_340,In_1390,In_1568);
or U341 (N_341,In_1358,In_1994);
or U342 (N_342,In_1122,In_1409);
nand U343 (N_343,In_1637,In_131);
nor U344 (N_344,In_1945,In_1256);
nand U345 (N_345,N_123,In_1882);
nor U346 (N_346,In_1098,In_950);
nor U347 (N_347,In_287,In_1721);
or U348 (N_348,In_1524,In_586);
nor U349 (N_349,In_1621,In_762);
and U350 (N_350,In_1150,In_650);
nor U351 (N_351,In_1755,In_1542);
xor U352 (N_352,In_1680,In_611);
xnor U353 (N_353,N_52,N_28);
nand U354 (N_354,In_546,In_1724);
nor U355 (N_355,In_744,In_1696);
or U356 (N_356,In_1469,In_1505);
nand U357 (N_357,In_1968,In_756);
and U358 (N_358,In_1042,In_132);
nand U359 (N_359,N_275,N_44);
nor U360 (N_360,In_1341,In_1922);
nand U361 (N_361,In_1480,In_956);
xnor U362 (N_362,In_95,In_1974);
nand U363 (N_363,In_1726,In_314);
nand U364 (N_364,In_1488,In_1975);
nand U365 (N_365,In_519,In_1718);
xnor U366 (N_366,In_938,In_55);
or U367 (N_367,N_169,In_1478);
nand U368 (N_368,In_365,N_189);
xor U369 (N_369,In_789,In_614);
or U370 (N_370,N_299,In_434);
xor U371 (N_371,In_965,In_1143);
nand U372 (N_372,In_1311,N_248);
or U373 (N_373,In_1014,N_104);
or U374 (N_374,In_924,In_285);
nor U375 (N_375,N_250,In_770);
or U376 (N_376,In_963,N_170);
or U377 (N_377,In_1776,In_833);
or U378 (N_378,In_657,In_1110);
or U379 (N_379,In_1527,N_132);
and U380 (N_380,N_126,In_454);
and U381 (N_381,In_1289,In_1497);
and U382 (N_382,In_1038,N_6);
nand U383 (N_383,In_1958,In_1228);
or U384 (N_384,In_1884,In_1187);
and U385 (N_385,In_1600,N_53);
nand U386 (N_386,In_1159,In_1224);
nand U387 (N_387,In_823,In_989);
and U388 (N_388,In_98,N_11);
and U389 (N_389,In_1555,In_1112);
nand U390 (N_390,In_1253,In_1764);
xor U391 (N_391,In_479,In_186);
or U392 (N_392,N_277,In_1040);
and U393 (N_393,In_1604,In_1547);
nor U394 (N_394,In_1903,In_176);
xnor U395 (N_395,In_954,In_81);
or U396 (N_396,N_147,In_976);
nand U397 (N_397,In_830,In_676);
nand U398 (N_398,In_1705,N_318);
and U399 (N_399,In_1624,In_1777);
and U400 (N_400,In_103,In_574);
xnor U401 (N_401,In_1240,In_1644);
xor U402 (N_402,N_305,N_79);
nand U403 (N_403,N_82,In_1914);
nand U404 (N_404,N_71,In_1820);
and U405 (N_405,In_793,N_98);
nand U406 (N_406,N_167,N_272);
or U407 (N_407,N_294,In_1971);
xnor U408 (N_408,N_315,In_2);
xor U409 (N_409,N_221,In_1658);
or U410 (N_410,In_786,In_164);
nand U411 (N_411,In_945,N_282);
nand U412 (N_412,In_1034,In_1221);
and U413 (N_413,In_438,N_197);
or U414 (N_414,In_1147,In_715);
nand U415 (N_415,N_247,In_1423);
or U416 (N_416,In_1425,In_1007);
or U417 (N_417,In_942,In_480);
nor U418 (N_418,In_1073,In_1319);
nor U419 (N_419,In_496,In_810);
or U420 (N_420,In_1440,In_711);
and U421 (N_421,N_151,In_1212);
xor U422 (N_422,In_1632,In_1207);
nor U423 (N_423,In_1051,In_704);
xnor U424 (N_424,In_1715,In_1981);
nand U425 (N_425,In_1429,In_258);
nand U426 (N_426,In_433,In_1120);
nand U427 (N_427,In_549,In_1226);
xor U428 (N_428,In_1699,In_1371);
xor U429 (N_429,In_1338,In_1024);
xor U430 (N_430,In_1937,N_279);
xnor U431 (N_431,In_951,N_195);
and U432 (N_432,In_303,In_573);
xor U433 (N_433,In_47,N_16);
nand U434 (N_434,In_276,In_955);
or U435 (N_435,In_0,In_1824);
or U436 (N_436,In_1570,In_1452);
nand U437 (N_437,N_130,In_403);
nor U438 (N_438,In_1407,In_443);
xnor U439 (N_439,In_494,In_814);
or U440 (N_440,In_296,In_871);
xnor U441 (N_441,In_1267,In_1263);
or U442 (N_442,In_1470,N_280);
xnor U443 (N_443,In_1843,In_537);
or U444 (N_444,In_1586,In_26);
and U445 (N_445,In_1036,In_630);
xor U446 (N_446,In_783,In_1905);
xnor U447 (N_447,In_733,In_1897);
nand U448 (N_448,In_644,In_980);
or U449 (N_449,In_289,In_576);
nor U450 (N_450,In_588,N_9);
nor U451 (N_451,N_278,In_448);
xnor U452 (N_452,In_245,In_1456);
or U453 (N_453,In_1988,In_1046);
xnor U454 (N_454,In_1938,In_301);
and U455 (N_455,In_1001,In_1580);
nand U456 (N_456,In_1594,In_684);
or U457 (N_457,N_145,In_1070);
xnor U458 (N_458,In_66,In_1888);
and U459 (N_459,In_1591,In_1296);
xor U460 (N_460,In_1634,In_288);
and U461 (N_461,N_103,In_722);
or U462 (N_462,N_260,In_1503);
xor U463 (N_463,N_213,In_977);
and U464 (N_464,In_1379,In_476);
or U465 (N_465,In_599,N_246);
xor U466 (N_466,N_237,In_1947);
or U467 (N_467,In_153,In_310);
xor U468 (N_468,In_1374,In_1862);
nand U469 (N_469,In_360,In_1655);
nand U470 (N_470,N_257,In_509);
xnor U471 (N_471,N_236,N_109);
or U472 (N_472,In_1025,In_1635);
xnor U473 (N_473,In_638,In_788);
and U474 (N_474,N_100,In_320);
or U475 (N_475,In_326,In_87);
and U476 (N_476,N_242,In_195);
nor U477 (N_477,N_172,In_1281);
nor U478 (N_478,In_1075,In_370);
xnor U479 (N_479,N_165,In_1208);
and U480 (N_480,N_293,In_1619);
nand U481 (N_481,In_932,In_906);
or U482 (N_482,In_1697,In_1142);
nand U483 (N_483,In_1161,In_1428);
nand U484 (N_484,In_1529,In_250);
nor U485 (N_485,N_1,In_811);
nor U486 (N_486,N_419,N_10);
nand U487 (N_487,N_54,In_110);
nand U488 (N_488,In_1551,In_1230);
xnor U489 (N_489,In_332,In_1264);
nand U490 (N_490,N_56,N_251);
or U491 (N_491,In_612,In_265);
and U492 (N_492,N_373,In_1784);
or U493 (N_493,In_1996,N_453);
nor U494 (N_494,In_481,N_348);
nor U495 (N_495,In_1190,In_1086);
nor U496 (N_496,In_1079,In_1787);
xnor U497 (N_497,N_424,In_1077);
nor U498 (N_498,N_395,In_805);
xnor U499 (N_499,N_451,In_719);
nor U500 (N_500,N_381,N_19);
nand U501 (N_501,In_391,In_834);
and U502 (N_502,In_226,In_18);
xnor U503 (N_503,N_302,In_726);
and U504 (N_504,In_300,In_34);
and U505 (N_505,In_893,N_166);
xnor U506 (N_506,N_48,N_316);
nand U507 (N_507,In_367,In_1649);
or U508 (N_508,In_1178,In_357);
nand U509 (N_509,N_330,N_162);
or U510 (N_510,In_1443,In_1153);
and U511 (N_511,N_235,In_1676);
and U512 (N_512,In_1302,In_1545);
and U513 (N_513,In_1910,In_171);
xor U514 (N_514,In_1747,In_1869);
and U515 (N_515,In_1250,In_259);
and U516 (N_516,In_764,In_295);
and U517 (N_517,In_506,In_1574);
nand U518 (N_518,In_1303,In_815);
and U519 (N_519,In_577,In_1864);
nor U520 (N_520,In_1695,N_358);
nand U521 (N_521,N_286,In_1398);
nor U522 (N_522,N_378,In_858);
nand U523 (N_523,In_946,N_258);
or U524 (N_524,N_352,In_1612);
xor U525 (N_525,In_334,In_1801);
or U526 (N_526,In_161,In_899);
and U527 (N_527,In_203,N_436);
nand U528 (N_528,N_264,In_633);
nand U529 (N_529,In_1006,N_127);
and U530 (N_530,In_1397,N_267);
and U531 (N_531,In_1437,In_46);
xor U532 (N_532,N_332,In_826);
or U533 (N_533,N_469,In_1797);
nand U534 (N_534,In_339,In_503);
nand U535 (N_535,In_1387,N_448);
nand U536 (N_536,In_925,N_124);
xor U537 (N_537,N_34,In_1265);
and U538 (N_538,N_365,In_101);
nor U539 (N_539,In_212,N_152);
and U540 (N_540,N_339,In_1483);
or U541 (N_541,In_358,In_191);
xor U542 (N_542,In_1318,In_986);
or U543 (N_543,In_1989,In_1033);
xor U544 (N_544,In_670,In_1273);
or U545 (N_545,In_665,N_58);
and U546 (N_546,In_898,In_147);
nand U547 (N_547,N_4,In_1541);
nand U548 (N_548,N_65,In_1515);
nor U549 (N_549,In_1314,In_521);
xor U550 (N_550,In_275,N_382);
nor U551 (N_551,N_392,In_1465);
nand U552 (N_552,N_383,N_325);
nor U553 (N_553,In_411,N_83);
or U554 (N_554,N_427,In_1401);
nor U555 (N_555,N_335,N_60);
nor U556 (N_556,N_418,N_292);
nor U557 (N_557,In_1180,N_323);
or U558 (N_558,N_470,N_35);
or U559 (N_559,In_104,In_392);
nor U560 (N_560,In_781,In_831);
and U561 (N_561,N_283,In_194);
nor U562 (N_562,N_429,In_1162);
xnor U563 (N_563,In_1901,In_769);
or U564 (N_564,In_1450,In_1088);
xor U565 (N_565,In_757,N_406);
xor U566 (N_566,In_1074,In_1044);
and U567 (N_567,In_1842,In_914);
nor U568 (N_568,In_1140,In_227);
and U569 (N_569,In_1214,In_1907);
nor U570 (N_570,In_1346,In_129);
xnor U571 (N_571,N_426,In_455);
or U572 (N_572,In_571,In_1217);
xor U573 (N_573,In_1317,In_1706);
and U574 (N_574,In_1572,N_475);
and U575 (N_575,In_1514,In_1475);
nor U576 (N_576,In_418,In_880);
or U577 (N_577,In_1786,N_161);
and U578 (N_578,In_112,In_580);
xnor U579 (N_579,In_337,In_996);
and U580 (N_580,In_419,N_174);
or U581 (N_581,In_1951,In_1231);
and U582 (N_582,In_550,N_380);
xnor U583 (N_583,In_1919,In_634);
or U584 (N_584,In_1157,N_238);
and U585 (N_585,In_1849,In_1106);
nor U586 (N_586,In_1136,In_1877);
nor U587 (N_587,In_1553,In_1270);
nand U588 (N_588,In_373,N_43);
or U589 (N_589,N_160,In_1083);
nand U590 (N_590,N_66,In_773);
and U591 (N_591,In_163,In_1335);
nand U592 (N_592,In_141,N_254);
nor U593 (N_593,In_1977,In_852);
nor U594 (N_594,In_1647,In_384);
xnor U595 (N_595,In_1005,In_1929);
xor U596 (N_596,In_1306,N_344);
nand U597 (N_597,In_1352,In_1510);
xnor U598 (N_598,N_255,In_1536);
nand U599 (N_599,N_321,N_449);
xor U600 (N_600,In_1540,N_210);
nor U601 (N_601,In_1415,In_1902);
nor U602 (N_602,In_539,N_439);
nand U603 (N_603,In_1539,In_342);
and U604 (N_604,In_1554,N_200);
nor U605 (N_605,In_994,In_1690);
nor U606 (N_606,N_412,In_335);
xor U607 (N_607,In_910,N_456);
xnor U608 (N_608,In_836,In_190);
nand U609 (N_609,In_297,In_1299);
nand U610 (N_610,N_120,N_135);
or U611 (N_611,In_372,N_438);
or U612 (N_612,In_1434,N_241);
or U613 (N_613,In_504,In_1427);
xor U614 (N_614,In_1838,In_578);
or U615 (N_615,In_1674,N_112);
xor U616 (N_616,N_455,N_408);
and U617 (N_617,In_1620,In_111);
and U618 (N_618,N_21,N_403);
xor U619 (N_619,In_225,N_303);
xor U620 (N_620,In_318,In_944);
nor U621 (N_621,In_65,In_626);
and U622 (N_622,In_1218,In_566);
nand U623 (N_623,In_222,N_240);
or U624 (N_624,N_196,In_935);
nand U625 (N_625,In_901,In_221);
nor U626 (N_626,In_1418,N_89);
and U627 (N_627,N_217,N_108);
nor U628 (N_628,N_304,In_1511);
or U629 (N_629,In_706,In_601);
xor U630 (N_630,In_1416,N_266);
xor U631 (N_631,N_346,N_0);
and U632 (N_632,In_1194,In_401);
nand U633 (N_633,In_624,In_1700);
nor U634 (N_634,In_1976,In_386);
nand U635 (N_635,In_1973,In_444);
nand U636 (N_636,In_1562,N_99);
xor U637 (N_637,In_1350,In_740);
or U638 (N_638,In_1928,In_1760);
xnor U639 (N_639,In_1961,N_309);
nor U640 (N_640,In_1500,N_508);
or U641 (N_641,In_992,In_182);
and U642 (N_642,In_1245,N_45);
xor U643 (N_643,N_192,In_64);
or U644 (N_644,N_212,In_1852);
nor U645 (N_645,In_1549,N_425);
or U646 (N_646,In_600,In_526);
or U647 (N_647,In_987,In_1065);
xor U648 (N_648,In_1,N_559);
xor U649 (N_649,N_354,In_1707);
xor U650 (N_650,In_698,In_1731);
nand U651 (N_651,In_1206,In_1479);
or U652 (N_652,N_541,In_14);
xor U653 (N_653,In_1163,In_183);
xor U654 (N_654,In_1880,N_369);
nor U655 (N_655,In_782,In_640);
or U656 (N_656,In_1356,In_290);
nor U657 (N_657,In_1189,N_599);
nor U658 (N_658,In_741,In_864);
and U659 (N_659,In_721,In_1284);
nand U660 (N_660,In_585,In_1955);
xor U661 (N_661,In_1670,In_631);
or U662 (N_662,In_1790,N_75);
xnor U663 (N_663,In_607,N_592);
nor U664 (N_664,In_197,In_1908);
or U665 (N_665,N_624,In_1344);
and U666 (N_666,In_22,In_727);
or U667 (N_667,In_635,In_845);
nand U668 (N_668,In_1238,In_1909);
nand U669 (N_669,In_1948,In_749);
and U670 (N_670,In_1451,N_281);
nor U671 (N_671,N_284,In_36);
nor U672 (N_672,In_933,In_139);
or U673 (N_673,In_1329,In_1255);
xnor U674 (N_674,In_660,In_655);
nand U675 (N_675,In_364,In_422);
nor U676 (N_676,In_674,N_588);
nor U677 (N_677,N_466,N_131);
and U678 (N_678,In_552,In_736);
or U679 (N_679,In_1710,In_462);
xnor U680 (N_680,N_320,N_533);
and U681 (N_681,In_1494,In_929);
xnor U682 (N_682,N_18,In_1814);
nand U683 (N_683,N_495,In_1980);
or U684 (N_684,In_1688,In_463);
or U685 (N_685,In_274,In_469);
xnor U686 (N_686,N_603,In_1215);
or U687 (N_687,N_597,In_378);
nand U688 (N_688,In_1761,N_634);
or U689 (N_689,In_1692,N_459);
nor U690 (N_690,In_77,In_820);
xnor U691 (N_691,N_450,In_1213);
nor U692 (N_692,In_1204,N_62);
or U693 (N_693,N_228,N_567);
nor U694 (N_694,In_1926,In_369);
nand U695 (N_695,N_76,In_1596);
xor U696 (N_696,N_173,In_921);
and U697 (N_697,In_430,In_1833);
and U698 (N_698,In_1293,In_1512);
and U699 (N_699,N_128,In_1166);
or U700 (N_700,N_400,In_1626);
nor U701 (N_701,In_1682,N_612);
nand U702 (N_702,N_133,N_572);
or U703 (N_703,N_548,In_477);
or U704 (N_704,N_421,In_590);
and U705 (N_705,In_1363,In_912);
nor U706 (N_706,In_1171,In_489);
and U707 (N_707,In_1368,In_1210);
nand U708 (N_708,In_1460,N_598);
and U709 (N_709,In_1087,N_33);
xor U710 (N_710,N_523,N_374);
nand U711 (N_711,In_891,In_1652);
and U712 (N_712,N_7,In_1271);
nand U713 (N_713,N_61,In_485);
and U714 (N_714,N_556,In_473);
xnor U715 (N_715,In_1518,In_445);
nor U716 (N_716,In_1100,N_385);
xnor U717 (N_717,N_190,In_446);
or U718 (N_718,In_1282,In_488);
or U719 (N_719,N_494,N_394);
nor U720 (N_720,In_1385,In_809);
xnor U721 (N_721,In_1431,In_1173);
and U722 (N_722,N_518,In_754);
or U723 (N_723,In_126,In_1045);
or U724 (N_724,N_506,In_1091);
and U725 (N_725,In_1059,In_1691);
nor U726 (N_726,In_96,In_882);
or U727 (N_727,In_1714,In_1751);
xor U728 (N_728,N_356,In_412);
and U729 (N_729,In_1939,In_230);
xor U730 (N_730,N_199,In_116);
nand U731 (N_731,In_196,In_1442);
or U732 (N_732,In_1121,N_410);
xnor U733 (N_733,In_387,In_647);
or U734 (N_734,In_74,N_589);
nand U735 (N_735,N_566,In_884);
and U736 (N_736,N_140,In_796);
xor U737 (N_737,N_85,N_639);
nor U738 (N_738,In_1246,In_556);
xor U739 (N_739,In_1694,In_1915);
and U740 (N_740,In_1782,N_143);
xnor U741 (N_741,N_532,N_491);
and U742 (N_742,In_1366,In_466);
nand U743 (N_743,In_1345,In_371);
nor U744 (N_744,N_413,N_440);
and U745 (N_745,In_113,In_157);
and U746 (N_746,In_1999,In_1932);
nand U747 (N_747,In_1672,N_476);
or U748 (N_748,In_255,N_136);
and U749 (N_749,N_606,In_1004);
xor U750 (N_750,N_564,In_915);
and U751 (N_751,In_1826,In_916);
nor U752 (N_752,In_67,In_1496);
and U753 (N_753,In_1592,N_573);
nor U754 (N_754,In_1750,In_653);
xor U755 (N_755,In_82,N_265);
xnor U756 (N_756,In_725,In_668);
or U757 (N_757,In_928,In_1493);
or U758 (N_758,N_252,In_345);
nand U759 (N_759,In_1463,N_537);
or U760 (N_760,N_333,In_904);
nor U761 (N_761,In_1956,In_1816);
or U762 (N_762,N_544,In_905);
xor U763 (N_763,In_1708,In_735);
and U764 (N_764,In_598,N_479);
xor U765 (N_765,N_273,In_217);
nand U766 (N_766,N_524,In_1251);
xor U767 (N_767,In_1054,N_306);
or U768 (N_768,In_94,N_307);
or U769 (N_769,In_1810,N_347);
or U770 (N_770,In_1712,N_458);
and U771 (N_771,In_267,In_853);
nor U772 (N_772,In_1322,N_142);
nand U773 (N_773,In_37,In_1830);
and U774 (N_774,In_686,In_1656);
nand U775 (N_775,N_405,In_1285);
nand U776 (N_776,In_1648,In_424);
and U777 (N_777,In_405,In_1891);
xor U778 (N_778,In_449,N_338);
xnor U779 (N_779,In_843,N_342);
nor U780 (N_780,In_1148,In_671);
xor U781 (N_781,N_622,N_411);
nor U782 (N_782,In_240,In_1917);
or U783 (N_783,N_467,In_1788);
nor U784 (N_784,N_371,In_1439);
nand U785 (N_785,In_597,In_872);
xnor U786 (N_786,N_78,In_1584);
and U787 (N_787,In_1807,In_534);
nor U788 (N_788,In_170,In_1359);
xor U789 (N_789,In_1300,In_1061);
or U790 (N_790,In_1609,In_92);
or U791 (N_791,In_1734,N_474);
or U792 (N_792,N_341,N_525);
and U793 (N_793,In_1597,In_234);
or U794 (N_794,In_1866,N_638);
xnor U795 (N_795,N_501,In_1693);
nor U796 (N_796,In_1468,In_169);
or U797 (N_797,N_328,In_724);
nand U798 (N_798,N_636,In_1185);
or U799 (N_799,In_246,In_490);
nand U800 (N_800,In_470,In_596);
nor U801 (N_801,N_661,In_842);
or U802 (N_802,In_12,N_397);
nor U803 (N_803,In_1313,N_640);
or U804 (N_804,In_120,N_692);
nor U805 (N_805,In_1115,In_1198);
nor U806 (N_806,N_389,In_1894);
nand U807 (N_807,In_527,N_92);
and U808 (N_808,In_457,N_685);
nand U809 (N_809,In_1942,In_1732);
or U810 (N_810,In_1738,In_1133);
xnor U811 (N_811,In_930,N_445);
and U812 (N_812,N_617,In_799);
nand U813 (N_813,N_40,In_959);
and U814 (N_814,In_1272,In_178);
nand U815 (N_815,In_1227,N_297);
or U816 (N_816,In_659,N_550);
and U817 (N_817,N_175,In_1030);
and U818 (N_818,In_1235,In_666);
nor U819 (N_819,In_1332,N_704);
xor U820 (N_820,N_722,In_822);
xor U821 (N_821,In_1276,In_1375);
or U822 (N_822,In_699,N_596);
nor U823 (N_823,N_547,N_37);
xnor U824 (N_824,In_1484,In_869);
and U825 (N_825,In_937,In_1124);
nand U826 (N_826,N_349,In_1105);
nand U827 (N_827,In_1965,In_936);
xnor U828 (N_828,In_1865,N_500);
or U829 (N_829,In_1454,In_900);
nand U830 (N_830,In_366,In_1191);
or U831 (N_831,In_1504,N_668);
nand U832 (N_832,N_757,In_926);
or U833 (N_833,N_12,N_579);
nand U834 (N_834,In_1793,In_1890);
nor U835 (N_835,N_77,In_961);
xor U836 (N_836,N_509,N_665);
nand U837 (N_837,In_172,N_717);
and U838 (N_838,In_1949,N_326);
nor U839 (N_839,N_361,N_765);
nor U840 (N_840,In_93,N_313);
nand U841 (N_841,In_1176,N_621);
xor U842 (N_842,In_1805,N_631);
or U843 (N_843,In_1384,In_1950);
and U844 (N_844,N_488,N_289);
nand U845 (N_845,In_873,In_1606);
nor U846 (N_846,N_202,N_205);
or U847 (N_847,N_464,N_608);
and U848 (N_848,N_64,N_185);
xor U849 (N_849,In_1730,In_484);
nor U850 (N_850,In_331,In_663);
nor U851 (N_851,N_271,In_1197);
nand U852 (N_852,N_274,In_361);
nor U853 (N_853,In_800,N_702);
and U854 (N_854,In_889,In_750);
or U855 (N_855,N_775,In_140);
and U856 (N_856,In_997,In_679);
xor U857 (N_857,N_336,N_719);
xor U858 (N_858,N_510,In_641);
xor U859 (N_859,N_489,N_5);
and U860 (N_860,N_288,In_1298);
xnor U861 (N_861,N_357,N_276);
and U862 (N_862,N_504,In_669);
and U863 (N_863,In_306,N_153);
nor U864 (N_864,In_985,In_804);
nor U865 (N_865,In_1498,N_317);
nor U866 (N_866,N_119,In_1403);
and U867 (N_867,In_713,N_234);
nand U868 (N_868,In_1261,In_91);
nand U869 (N_869,N_582,In_1802);
or U870 (N_870,In_286,In_940);
and U871 (N_871,In_1560,In_575);
or U872 (N_872,In_718,In_508);
nor U873 (N_873,In_105,In_1225);
nor U874 (N_874,N_673,N_270);
or U875 (N_875,N_515,N_615);
or U876 (N_876,N_180,In_1508);
nand U877 (N_877,In_1455,In_1277);
nand U878 (N_878,N_746,In_400);
and U879 (N_879,N_443,In_273);
or U880 (N_880,N_249,In_1111);
nand U881 (N_881,In_1164,In_1615);
or U882 (N_882,In_239,In_262);
or U883 (N_883,N_461,N_676);
nor U884 (N_884,N_710,In_1078);
xnor U885 (N_885,N_674,N_345);
xor U886 (N_886,N_186,In_543);
nand U887 (N_887,In_892,N_530);
xor U888 (N_888,N_343,In_1330);
and U889 (N_889,N_15,N_396);
nand U890 (N_890,In_1188,In_617);
nor U891 (N_891,In_1062,In_1158);
or U892 (N_892,In_923,In_1703);
and U893 (N_893,In_1952,In_1794);
xnor U894 (N_894,N_261,In_1935);
and U895 (N_895,In_729,N_122);
nand U896 (N_896,N_428,N_462);
nor U897 (N_897,N_563,In_1900);
nor U898 (N_898,N_786,In_649);
or U899 (N_899,In_1183,N_13);
nand U900 (N_900,In_158,In_1152);
or U901 (N_901,N_788,N_363);
or U902 (N_902,N_756,N_727);
nor U903 (N_903,In_316,In_1654);
or U904 (N_904,In_968,N_620);
nand U905 (N_905,In_1563,In_1766);
xnor U906 (N_906,N_670,In_1650);
xor U907 (N_907,N_107,In_1770);
xor U908 (N_908,N_613,In_1651);
and U909 (N_909,In_1039,N_791);
nor U910 (N_910,N_159,N_774);
nor U911 (N_911,In_1589,In_1085);
nand U912 (N_912,N_574,In_1066);
nor U913 (N_913,N_375,In_510);
nand U914 (N_914,In_627,In_559);
nor U915 (N_915,N_80,In_1686);
nor U916 (N_916,In_516,In_1791);
xor U917 (N_917,In_1064,N_780);
nand U918 (N_918,In_613,N_753);
or U919 (N_919,In_211,N_535);
and U920 (N_920,N_514,N_519);
xor U921 (N_921,N_367,N_468);
or U922 (N_922,In_1628,In_458);
nor U923 (N_923,N_253,In_150);
and U924 (N_924,N_497,In_1170);
nor U925 (N_925,N_675,N_762);
xor U926 (N_926,In_321,N_713);
or U927 (N_927,N_370,In_100);
nand U928 (N_928,In_293,N_460);
nor U929 (N_929,N_67,N_498);
or U930 (N_930,N_415,In_382);
xor U931 (N_931,In_1155,In_465);
xnor U932 (N_932,In_72,In_708);
and U933 (N_933,N_231,N_680);
or U934 (N_934,In_1172,In_1970);
or U935 (N_935,N_198,N_662);
and U936 (N_936,N_552,In_145);
nand U937 (N_937,In_1411,In_261);
or U938 (N_938,In_1139,In_1412);
and U939 (N_939,In_1446,In_1192);
nand U940 (N_940,In_908,N_434);
xnor U941 (N_941,In_1103,N_148);
or U942 (N_942,N_721,In_707);
or U943 (N_943,N_81,In_535);
or U944 (N_944,In_772,In_776);
or U945 (N_945,N_296,N_679);
and U946 (N_946,In_42,In_1339);
or U947 (N_947,N_546,N_102);
or U948 (N_948,N_739,In_108);
nand U949 (N_949,In_407,In_374);
nand U950 (N_950,In_1093,In_1243);
or U951 (N_951,In_175,N_794);
nor U952 (N_952,N_643,In_618);
nand U953 (N_953,N_472,N_14);
and U954 (N_954,In_119,In_497);
nor U955 (N_955,In_696,In_1199);
and U956 (N_956,In_461,In_51);
or U957 (N_957,N_3,N_219);
or U958 (N_958,In_389,In_1487);
xor U959 (N_959,In_208,N_372);
xnor U960 (N_960,N_600,N_310);
or U961 (N_961,N_898,N_946);
nand U962 (N_962,N_819,N_947);
and U963 (N_963,N_181,N_667);
nor U964 (N_964,In_1972,In_13);
or U965 (N_965,N_843,N_626);
nor U966 (N_966,In_909,N_194);
xnor U967 (N_967,N_430,N_890);
xnor U968 (N_968,In_478,In_1047);
and U969 (N_969,N_390,N_857);
xor U970 (N_970,In_1773,In_1027);
and U971 (N_971,N_571,N_203);
and U972 (N_972,In_1248,In_204);
nor U973 (N_973,In_453,In_887);
and U974 (N_974,In_215,N_940);
or U975 (N_975,N_637,N_790);
xnor U976 (N_976,In_1603,In_625);
or U977 (N_977,N_593,In_664);
or U978 (N_978,In_1847,N_576);
and U979 (N_979,N_929,N_672);
or U980 (N_980,In_1076,In_1467);
or U981 (N_981,In_1643,N_329);
nor U982 (N_982,N_209,N_955);
and U983 (N_983,In_1128,N_730);
nand U984 (N_984,N_184,In_138);
nand U985 (N_985,In_970,N_134);
nor U986 (N_986,In_1169,N_645);
nand U987 (N_987,N_301,In_1774);
and U988 (N_988,N_377,N_854);
xor U989 (N_989,N_287,N_611);
nand U990 (N_990,In_69,N_740);
or U991 (N_991,In_1978,In_1585);
nand U992 (N_992,In_1964,N_268);
and U993 (N_993,N_401,N_919);
nand U994 (N_994,N_732,In_1821);
nand U995 (N_995,N_759,In_1491);
or U996 (N_996,In_429,In_1114);
xor U997 (N_997,In_1331,N_555);
nand U998 (N_998,In_417,N_889);
and U999 (N_999,In_406,N_912);
or U1000 (N_1000,In_1983,In_1987);
nand U1001 (N_1001,In_149,In_491);
xor U1002 (N_1002,N_379,In_379);
nor U1003 (N_1003,N_393,N_838);
nand U1004 (N_1004,N_892,N_324);
and U1005 (N_1005,In_1702,N_243);
xnor U1006 (N_1006,In_472,In_284);
and U1007 (N_1007,N_211,N_931);
xor U1008 (N_1008,In_1011,In_1222);
nor U1009 (N_1009,In_1507,N_825);
xor U1010 (N_1010,In_257,In_1472);
xnor U1011 (N_1011,N_543,In_248);
nand U1012 (N_1012,In_1631,N_649);
nor U1013 (N_1013,N_945,N_768);
and U1014 (N_1014,N_862,N_853);
nor U1015 (N_1015,In_883,In_952);
xnor U1016 (N_1016,In_1582,N_527);
nor U1017 (N_1017,N_844,N_602);
or U1018 (N_1018,N_577,N_734);
xor U1019 (N_1019,In_75,In_180);
nor U1020 (N_1020,N_42,In_1930);
or U1021 (N_1021,N_118,In_808);
and U1022 (N_1022,N_485,In_1287);
nor U1023 (N_1023,N_568,In_1304);
or U1024 (N_1024,N_641,In_821);
and U1025 (N_1025,N_229,N_737);
and U1026 (N_1026,N_747,In_1422);
and U1027 (N_1027,In_1471,In_848);
nor U1028 (N_1028,N_290,N_879);
nand U1029 (N_1029,In_244,In_394);
nor U1030 (N_1030,N_630,N_669);
and U1031 (N_1031,In_606,N_594);
and U1032 (N_1032,In_767,In_1080);
and U1033 (N_1033,In_1196,In_270);
and U1034 (N_1034,In_1681,N_591);
xnor U1035 (N_1035,In_1671,In_432);
or U1036 (N_1036,In_238,N_867);
and U1037 (N_1037,In_1943,N_864);
nand U1038 (N_1038,N_331,N_881);
nand U1039 (N_1039,N_549,N_74);
nand U1040 (N_1040,In_1646,N_480);
nor U1041 (N_1041,N_540,N_214);
or U1042 (N_1042,In_280,In_953);
and U1043 (N_1043,N_55,In_390);
xnor U1044 (N_1044,N_644,N_863);
nor U1045 (N_1045,In_1071,N_957);
nor U1046 (N_1046,N_141,N_832);
or U1047 (N_1047,N_870,In_1548);
and U1048 (N_1048,N_876,In_998);
nand U1049 (N_1049,N_726,N_51);
nor U1050 (N_1050,In_553,In_219);
nand U1051 (N_1051,N_220,In_228);
and U1052 (N_1052,In_247,In_21);
or U1053 (N_1053,In_1957,In_1780);
xnor U1054 (N_1054,N_91,N_828);
nand U1055 (N_1055,N_386,In_456);
or U1056 (N_1056,N_50,In_1249);
xnor U1057 (N_1057,In_1579,In_999);
nor U1058 (N_1058,In_639,N_913);
xnor U1059 (N_1059,N_918,In_1557);
and U1060 (N_1060,In_408,N_835);
nand U1061 (N_1061,In_1683,N_650);
and U1062 (N_1062,N_351,N_677);
and U1063 (N_1063,N_789,In_579);
nor U1064 (N_1064,In_1516,In_214);
or U1065 (N_1065,In_185,In_1662);
or U1066 (N_1066,In_1229,N_452);
nor U1067 (N_1067,N_471,N_793);
or U1068 (N_1068,N_745,N_298);
and U1069 (N_1069,N_949,N_952);
and U1070 (N_1070,In_1459,In_1184);
and U1071 (N_1071,N_922,In_336);
or U1072 (N_1072,In_1883,In_1723);
and U1073 (N_1073,N_285,N_366);
xnor U1074 (N_1074,N_778,N_796);
xor U1075 (N_1075,In_1067,In_311);
or U1076 (N_1076,N_736,In_299);
and U1077 (N_1077,In_1960,N_842);
nor U1078 (N_1078,N_417,In_1360);
and U1079 (N_1079,N_880,N_911);
or U1080 (N_1080,N_664,N_826);
xnor U1081 (N_1081,N_182,N_805);
nor U1082 (N_1082,N_125,In_1921);
nor U1083 (N_1083,In_1175,N_291);
nor U1084 (N_1084,N_785,In_315);
or U1085 (N_1085,In_1899,In_967);
nand U1086 (N_1086,In_734,N_792);
nand U1087 (N_1087,N_821,In_1876);
and U1088 (N_1088,N_941,In_154);
nor U1089 (N_1089,N_811,In_1295);
nand U1090 (N_1090,In_629,N_795);
xnor U1091 (N_1091,In_1581,N_761);
xor U1092 (N_1092,N_529,In_803);
xnor U1093 (N_1093,In_1778,N_681);
and U1094 (N_1094,In_1783,N_388);
and U1095 (N_1095,N_893,In_1135);
or U1096 (N_1096,N_755,In_584);
nor U1097 (N_1097,In_731,In_1413);
and U1098 (N_1098,N_711,In_948);
and U1099 (N_1099,In_33,In_1309);
nand U1100 (N_1100,N_729,N_808);
xor U1101 (N_1101,In_1954,N_463);
and U1102 (N_1102,In_188,N_944);
nand U1103 (N_1103,In_1669,In_1326);
nand U1104 (N_1104,N_206,In_779);
or U1105 (N_1105,In_1550,N_245);
xor U1106 (N_1106,N_715,N_697);
xor U1107 (N_1107,In_865,In_623);
xnor U1108 (N_1108,N_860,N_575);
xor U1109 (N_1109,In_78,In_329);
xnor U1110 (N_1110,In_957,N_49);
xor U1111 (N_1111,N_25,In_531);
or U1112 (N_1112,N_750,In_349);
nor U1113 (N_1113,N_553,N_771);
nand U1114 (N_1114,N_505,N_551);
or U1115 (N_1115,N_822,In_73);
nand U1116 (N_1116,N_660,In_1666);
xnor U1117 (N_1117,N_502,N_215);
or U1118 (N_1118,In_1010,N_168);
nor U1119 (N_1119,N_473,N_743);
nand U1120 (N_1120,N_814,N_1087);
or U1121 (N_1121,N_1108,N_1055);
xor U1122 (N_1122,N_1078,In_19);
xnor U1123 (N_1123,N_295,In_1898);
nor U1124 (N_1124,N_1109,N_437);
nor U1125 (N_1125,N_223,In_1940);
and U1126 (N_1126,N_868,In_589);
or U1127 (N_1127,N_787,In_1875);
or U1128 (N_1128,N_404,N_908);
nor U1129 (N_1129,In_988,In_530);
nor U1130 (N_1130,N_1049,In_308);
and U1131 (N_1131,In_1305,In_1094);
and U1132 (N_1132,In_866,In_431);
and U1133 (N_1133,N_486,N_812);
and U1134 (N_1134,In_1863,In_1854);
nor U1135 (N_1135,N_187,In_1871);
nor U1136 (N_1136,N_623,N_1043);
nand U1137 (N_1137,N_885,In_1622);
xnor U1138 (N_1138,N_1050,In_1109);
nand U1139 (N_1139,N_1119,N_262);
nand U1140 (N_1140,N_849,In_1832);
and U1141 (N_1141,N_482,N_968);
nand U1142 (N_1142,In_59,In_1499);
or U1143 (N_1143,N_609,In_399);
or U1144 (N_1144,In_541,N_815);
xor U1145 (N_1145,N_1086,In_703);
and U1146 (N_1146,N_635,In_1711);
nor U1147 (N_1147,N_688,N_1063);
nand U1148 (N_1148,In_241,In_1145);
and U1149 (N_1149,In_1753,In_813);
nor U1150 (N_1150,N_927,N_744);
xnor U1151 (N_1151,N_995,N_1071);
or U1152 (N_1152,N_772,In_1870);
xor U1153 (N_1153,In_173,N_416);
nor U1154 (N_1154,N_610,N_1081);
xor U1155 (N_1155,In_43,N_188);
nand U1156 (N_1156,N_97,In_771);
nand U1157 (N_1157,In_806,N_1036);
and U1158 (N_1158,In_538,In_1984);
or U1159 (N_1159,N_1080,N_935);
and U1160 (N_1160,N_801,In_495);
nor U1161 (N_1161,In_85,In_1406);
or U1162 (N_1162,N_554,N_962);
nand U1163 (N_1163,N_604,N_781);
or U1164 (N_1164,In_1102,In_1716);
nor U1165 (N_1165,N_678,N_1083);
nand U1166 (N_1166,In_1174,N_938);
nor U1167 (N_1167,N_31,In_1449);
or U1168 (N_1168,In_363,N_176);
or U1169 (N_1169,In_555,N_866);
or U1170 (N_1170,N_259,In_114);
and U1171 (N_1171,In_385,N_872);
nor U1172 (N_1172,N_738,N_671);
and U1173 (N_1173,In_1664,In_745);
xor U1174 (N_1174,N_784,N_993);
or U1175 (N_1175,In_1785,N_724);
nand U1176 (N_1176,N_226,N_531);
nor U1177 (N_1177,N_1011,In_1092);
and U1178 (N_1178,N_1112,N_820);
nor U1179 (N_1179,In_253,N_769);
or U1180 (N_1180,N_779,N_1032);
and U1181 (N_1181,N_901,In_283);
or U1182 (N_1182,In_1571,N_706);
and U1183 (N_1183,N_951,In_200);
and U1184 (N_1184,N_985,In_646);
or U1185 (N_1185,In_1349,N_457);
or U1186 (N_1186,In_716,N_1040);
or U1187 (N_1187,N_658,In_583);
nand U1188 (N_1188,In_1057,N_958);
nor U1189 (N_1189,N_1052,In_292);
nand U1190 (N_1190,N_1013,N_886);
and U1191 (N_1191,N_855,In_1684);
xnor U1192 (N_1192,N_694,In_1041);
xor U1193 (N_1193,N_163,N_714);
and U1194 (N_1194,N_431,N_848);
and U1195 (N_1195,N_539,N_1058);
and U1196 (N_1196,In_1081,N_850);
or U1197 (N_1197,In_500,N_896);
and U1198 (N_1198,N_322,N_806);
nor U1199 (N_1199,In_1818,In_1639);
nand U1200 (N_1200,N_873,In_888);
and U1201 (N_1201,N_492,N_1065);
nand U1202 (N_1202,In_277,N_1085);
and U1203 (N_1203,N_542,N_964);
xor U1204 (N_1204,N_882,N_1031);
xnor U1205 (N_1205,N_813,N_818);
nor U1206 (N_1206,N_1098,N_391);
xnor U1207 (N_1207,N_783,N_707);
xnor U1208 (N_1208,In_1595,In_1324);
and U1209 (N_1209,In_1817,N_1017);
or U1210 (N_1210,N_222,In_1365);
xor U1211 (N_1211,N_939,In_739);
xnor U1212 (N_1212,N_350,N_1103);
nor U1213 (N_1213,In_1998,N_689);
and U1214 (N_1214,In_1096,N_399);
or U1215 (N_1215,N_364,In_1758);
or U1216 (N_1216,N_942,N_311);
or U1217 (N_1217,In_1722,N_628);
and U1218 (N_1218,In_1827,N_191);
and U1219 (N_1219,N_686,N_992);
nor U1220 (N_1220,N_903,N_232);
nor U1221 (N_1221,N_1110,N_384);
or U1222 (N_1222,In_1377,N_1064);
nand U1223 (N_1223,N_585,N_178);
nor U1224 (N_1224,N_1095,In_151);
and U1225 (N_1225,N_967,N_1026);
nand U1226 (N_1226,In_1886,N_725);
and U1227 (N_1227,In_148,N_659);
nand U1228 (N_1228,N_1059,In_499);
nor U1229 (N_1229,In_184,N_1027);
nand U1230 (N_1230,In_1395,In_1561);
and U1231 (N_1231,N_218,In_236);
nand U1232 (N_1232,In_524,N_22);
nand U1233 (N_1233,N_1073,In_1146);
or U1234 (N_1234,N_154,In_207);
nand U1235 (N_1235,N_914,N_751);
and U1236 (N_1236,In_1131,N_1090);
xnor U1237 (N_1237,N_923,In_264);
nor U1238 (N_1238,N_982,N_760);
nand U1239 (N_1239,N_368,N_46);
nor U1240 (N_1240,N_1106,N_522);
or U1241 (N_1241,N_875,N_1102);
nand U1242 (N_1242,N_987,In_1741);
or U1243 (N_1243,N_646,In_1749);
and U1244 (N_1244,N_936,N_1047);
nor U1245 (N_1245,In_1050,N_915);
or U1246 (N_1246,In_878,In_1967);
and U1247 (N_1247,In_1369,N_149);
nand U1248 (N_1248,In_38,In_1182);
or U1249 (N_1249,In_1608,In_1614);
nor U1250 (N_1250,N_146,N_63);
or U1251 (N_1251,N_193,N_442);
nand U1252 (N_1252,N_971,N_709);
or U1253 (N_1253,N_959,In_1532);
nand U1254 (N_1254,N_627,N_932);
or U1255 (N_1255,N_690,In_1426);
xnor U1256 (N_1256,N_1054,N_718);
or U1257 (N_1257,In_397,In_658);
and U1258 (N_1258,In_917,N_865);
nand U1259 (N_1259,N_948,In_1461);
xnor U1260 (N_1260,In_787,In_25);
xnor U1261 (N_1261,In_1633,N_845);
xnor U1262 (N_1262,In_427,In_919);
or U1263 (N_1263,N_605,N_619);
and U1264 (N_1264,N_1089,N_907);
and U1265 (N_1265,N_444,N_629);
nand U1266 (N_1266,N_1074,N_1053);
or U1267 (N_1267,In_474,In_319);
xnor U1268 (N_1268,In_766,In_115);
nor U1269 (N_1269,N_409,In_1543);
xor U1270 (N_1270,N_834,In_1492);
nand U1271 (N_1271,N_703,In_63);
nand U1272 (N_1272,In_643,N_560);
nand U1273 (N_1273,N_981,In_1242);
nor U1274 (N_1274,N_965,In_1101);
nor U1275 (N_1275,In_1701,N_269);
nor U1276 (N_1276,In_1982,In_1028);
or U1277 (N_1277,In_1058,N_569);
xor U1278 (N_1278,N_1104,N_871);
or U1279 (N_1279,N_1006,In_1376);
and U1280 (N_1280,N_824,In_701);
nand U1281 (N_1281,N_1163,N_816);
xnor U1282 (N_1282,N_1272,In_309);
and U1283 (N_1283,N_1220,In_256);
or U1284 (N_1284,In_774,In_1291);
nor U1285 (N_1285,N_1111,N_648);
nand U1286 (N_1286,In_1618,In_1232);
nor U1287 (N_1287,N_859,In_15);
nor U1288 (N_1288,In_1447,N_1174);
or U1289 (N_1289,N_1132,N_666);
or U1290 (N_1290,N_749,N_698);
or U1291 (N_1291,In_798,N_733);
xnor U1292 (N_1292,N_1237,In_1759);
nand U1293 (N_1293,N_1105,N_1183);
nand U1294 (N_1294,N_656,N_1208);
or U1295 (N_1295,N_595,N_1179);
nand U1296 (N_1296,N_155,N_969);
and U1297 (N_1297,N_586,N_764);
or U1298 (N_1298,In_791,In_23);
nand U1299 (N_1299,N_1259,N_490);
nor U1300 (N_1300,N_928,In_648);
nand U1301 (N_1301,N_735,In_1327);
and U1302 (N_1302,N_557,In_233);
nand U1303 (N_1303,In_824,N_976);
nor U1304 (N_1304,In_1012,N_116);
or U1305 (N_1305,N_477,N_1121);
and U1306 (N_1306,N_933,N_1155);
nand U1307 (N_1307,In_751,N_1010);
and U1308 (N_1308,N_695,In_426);
and U1309 (N_1309,In_862,In_1430);
or U1310 (N_1310,N_1021,N_999);
and U1311 (N_1311,N_1159,N_1162);
nor U1312 (N_1312,N_1124,N_720);
and U1313 (N_1313,N_804,N_1255);
or U1314 (N_1314,N_113,N_990);
xor U1315 (N_1315,In_1878,In_1856);
nand U1316 (N_1316,In_263,N_831);
and U1317 (N_1317,N_1115,In_351);
or U1318 (N_1318,N_1070,In_160);
nand U1319 (N_1319,N_841,N_956);
and U1320 (N_1320,In_978,In_628);
nand U1321 (N_1321,N_300,In_52);
nor U1322 (N_1322,N_137,N_984);
nand U1323 (N_1323,In_1072,N_513);
or U1324 (N_1324,N_1096,N_1266);
xor U1325 (N_1325,N_934,In_775);
nand U1326 (N_1326,N_225,N_111);
nand U1327 (N_1327,N_1185,N_1212);
nor U1328 (N_1328,In_1343,In_1893);
xnor U1329 (N_1329,N_1199,N_989);
or U1330 (N_1330,N_164,N_970);
and U1331 (N_1331,N_1037,N_1188);
nor U1332 (N_1332,In_714,N_950);
and U1333 (N_1333,N_1100,N_1149);
or U1334 (N_1334,N_712,In_1531);
or U1335 (N_1335,In_1018,N_700);
nand U1336 (N_1336,N_1168,N_693);
or U1337 (N_1337,N_1254,In_1477);
nor U1338 (N_1338,N_1206,In_738);
or U1339 (N_1339,N_742,In_902);
and U1340 (N_1340,N_902,N_1129);
and U1341 (N_1341,N_930,In_177);
xor U1342 (N_1342,N_516,N_1015);
and U1343 (N_1343,In_778,In_867);
xor U1344 (N_1344,N_1051,N_1008);
nand U1345 (N_1345,N_1094,N_1215);
and U1346 (N_1346,In_7,N_1033);
xnor U1347 (N_1347,In_682,In_1653);
or U1348 (N_1348,N_1161,In_879);
nor U1349 (N_1349,In_991,N_1262);
nand U1350 (N_1350,N_1197,N_1091);
nand U1351 (N_1351,In_54,N_708);
xnor U1352 (N_1352,In_1525,In_922);
nor U1353 (N_1353,N_57,N_1278);
xor U1354 (N_1354,In_1420,N_1125);
nand U1355 (N_1355,N_359,In_1168);
xnor U1356 (N_1356,N_1146,N_208);
nand U1357 (N_1357,In_513,In_460);
and U1358 (N_1358,N_1007,N_1048);
nor U1359 (N_1359,N_1225,N_1133);
or U1360 (N_1360,N_607,In_1923);
nand U1361 (N_1361,In_1808,N_960);
and U1362 (N_1362,N_1019,In_931);
or U1363 (N_1363,N_69,N_526);
or U1364 (N_1364,N_38,N_1114);
nand U1365 (N_1365,N_1204,N_1150);
xor U1366 (N_1366,N_1226,N_1099);
xnor U1367 (N_1367,In_352,In_282);
and U1368 (N_1368,N_263,N_906);
or U1369 (N_1369,In_1953,N_1195);
or U1370 (N_1370,In_243,In_1502);
and U1371 (N_1371,N_1257,N_983);
or U1372 (N_1372,In_1097,N_1228);
nor U1373 (N_1373,N_798,N_517);
nand U1374 (N_1374,N_1256,N_481);
nor U1375 (N_1375,N_1137,N_731);
or U1376 (N_1376,In_346,N_1144);
nor U1377 (N_1377,N_899,N_1209);
or U1378 (N_1378,In_854,N_974);
and U1379 (N_1379,N_601,N_1093);
xnor U1380 (N_1380,In_192,In_1049);
or U1381 (N_1381,N_691,N_625);
or U1382 (N_1382,N_1139,In_1137);
nor U1383 (N_1383,N_312,N_179);
nor U1384 (N_1384,N_925,N_891);
xor U1385 (N_1385,N_1030,N_767);
xnor U1386 (N_1386,In_1404,N_823);
xnor U1387 (N_1387,N_1219,N_1140);
xnor U1388 (N_1388,In_4,N_171);
or U1389 (N_1389,N_1077,N_632);
or U1390 (N_1390,In_533,In_35);
and U1391 (N_1391,N_1252,In_557);
or U1392 (N_1392,N_423,In_1887);
and U1393 (N_1393,In_1756,N_1041);
xor U1394 (N_1394,In_1269,N_1193);
or U1395 (N_1395,N_101,N_748);
xor U1396 (N_1396,N_642,N_1147);
xor U1397 (N_1397,N_1152,N_360);
nand U1398 (N_1398,N_1233,N_797);
nand U1399 (N_1399,N_654,In_1840);
xor U1400 (N_1400,N_1218,N_1243);
or U1401 (N_1401,N_1241,In_875);
and U1402 (N_1402,N_874,In_1623);
xnor U1403 (N_1403,N_478,In_1104);
nor U1404 (N_1404,N_1260,In_83);
nand U1405 (N_1405,In_1205,N_1275);
xor U1406 (N_1406,N_1224,N_1069);
and U1407 (N_1407,N_829,In_1219);
and U1408 (N_1408,In_1419,N_1191);
nor U1409 (N_1409,In_1789,N_777);
nor U1410 (N_1410,In_355,N_827);
or U1411 (N_1411,In_1082,In_1055);
nor U1412 (N_1412,N_1128,N_1184);
and U1413 (N_1413,In_442,N_534);
or U1414 (N_1414,N_1062,In_1925);
nand U1415 (N_1415,N_1061,N_1038);
or U1416 (N_1416,N_121,N_1171);
nor U1417 (N_1417,N_327,N_1142);
nand U1418 (N_1418,In_216,N_1214);
nor U1419 (N_1419,N_910,In_962);
nor U1420 (N_1420,In_1063,N_1239);
or U1421 (N_1421,In_5,N_1170);
and U1422 (N_1422,N_1117,N_926);
nand U1423 (N_1423,N_614,N_583);
nor U1424 (N_1424,N_1263,N_1097);
and U1425 (N_1425,N_1028,In_797);
nand U1426 (N_1426,In_737,N_651);
and U1427 (N_1427,N_1004,N_705);
nand U1428 (N_1428,In_1156,N_1165);
and U1429 (N_1429,In_680,N_570);
and U1430 (N_1430,N_652,In_1481);
and U1431 (N_1431,In_1026,N_72);
or U1432 (N_1432,In_1848,N_1205);
xnor U1433 (N_1433,N_741,In_57);
or U1434 (N_1434,In_327,N_1231);
xor U1435 (N_1435,In_544,N_177);
nor U1436 (N_1436,N_895,In_1482);
and U1437 (N_1437,In_1678,N_1221);
nand U1438 (N_1438,N_1250,N_1060);
nand U1439 (N_1439,N_447,N_39);
xor U1440 (N_1440,N_420,N_1432);
and U1441 (N_1441,N_1316,N_1294);
nor U1442 (N_1442,N_1056,N_1330);
nand U1443 (N_1443,N_1265,N_1201);
nand U1444 (N_1444,N_435,N_917);
nand U1445 (N_1445,N_973,N_963);
nor U1446 (N_1446,In_689,In_1850);
nor U1447 (N_1447,N_682,N_581);
or U1448 (N_1448,N_1284,In_350);
or U1449 (N_1449,N_1393,N_1292);
or U1450 (N_1450,N_565,N_1034);
and U1451 (N_1451,N_1419,In_1211);
nor U1452 (N_1452,N_1368,N_446);
or U1453 (N_1453,N_1302,N_1340);
and U1454 (N_1454,N_1075,N_528);
or U1455 (N_1455,N_684,In_710);
xnor U1456 (N_1456,N_1391,N_1076);
or U1457 (N_1457,N_1192,N_1012);
nor U1458 (N_1458,N_1135,In_569);
xor U1459 (N_1459,N_1082,N_1312);
nand U1460 (N_1460,In_563,N_1046);
or U1461 (N_1461,N_422,N_1386);
nor U1462 (N_1462,N_1067,N_1157);
and U1463 (N_1463,N_1268,In_1457);
and U1464 (N_1464,N_32,In_1292);
and U1465 (N_1465,In_302,In_1867);
or U1466 (N_1466,N_1180,N_1421);
xor U1467 (N_1467,N_362,N_1251);
or U1468 (N_1468,N_1194,N_1313);
or U1469 (N_1469,N_1308,N_47);
xor U1470 (N_1470,In_1565,In_181);
nand U1471 (N_1471,N_1002,N_1392);
or U1472 (N_1472,N_1406,N_1164);
or U1473 (N_1473,N_584,In_1521);
or U1474 (N_1474,N_1234,N_1359);
or U1475 (N_1475,In_1441,N_201);
xor U1476 (N_1476,N_687,N_996);
nor U1477 (N_1477,N_1323,In_86);
nand U1478 (N_1478,In_548,N_1230);
nor U1479 (N_1479,N_1305,In_1118);
nor U1480 (N_1480,N_1127,N_836);
nor U1481 (N_1481,N_810,N_1022);
or U1482 (N_1482,N_1299,N_244);
or U1483 (N_1483,N_1186,N_1236);
and U1484 (N_1484,N_1270,N_800);
nand U1485 (N_1485,N_1409,In_1099);
nor U1486 (N_1486,N_1280,N_1113);
or U1487 (N_1487,N_1177,In_1590);
or U1488 (N_1488,N_1375,In_1149);
or U1489 (N_1489,N_904,N_776);
nor U1490 (N_1490,N_1154,N_1235);
xor U1491 (N_1491,N_1153,N_1329);
or U1492 (N_1492,N_536,N_856);
nand U1493 (N_1493,N_696,In_839);
and U1494 (N_1494,N_770,N_1283);
nor U1495 (N_1495,N_545,N_1342);
and U1496 (N_1496,In_10,N_980);
nor U1497 (N_1497,In_128,N_1405);
or U1498 (N_1498,N_1317,N_998);
or U1499 (N_1499,N_975,N_782);
xnor U1500 (N_1500,N_978,In_1000);
nor U1501 (N_1501,N_878,N_1287);
or U1502 (N_1502,N_1143,N_1227);
and U1503 (N_1503,N_1203,In_266);
nor U1504 (N_1504,N_308,N_1309);
and U1505 (N_1505,N_766,N_1361);
and U1506 (N_1506,N_1176,N_802);
xor U1507 (N_1507,N_1399,N_1383);
or U1508 (N_1508,N_1417,N_1079);
xnor U1509 (N_1509,N_1356,In_1583);
nor U1510 (N_1510,In_1566,N_1424);
or U1511 (N_1511,N_897,N_1404);
nor U1512 (N_1512,N_900,N_1295);
or U1513 (N_1513,N_1300,N_1246);
xor U1514 (N_1514,N_1337,N_507);
and U1515 (N_1515,N_1365,N_1148);
xnor U1516 (N_1516,N_1364,N_877);
or U1517 (N_1517,N_1187,N_538);
or U1518 (N_1518,N_578,N_1369);
xor U1519 (N_1519,N_763,N_1293);
nor U1520 (N_1520,In_395,N_809);
or U1521 (N_1521,In_759,N_1437);
xnor U1522 (N_1522,N_465,N_1151);
xnor U1523 (N_1523,In_1445,N_580);
or U1524 (N_1524,N_1269,N_884);
nor U1525 (N_1525,N_846,N_1311);
nor U1526 (N_1526,N_1285,In_1200);
nand U1527 (N_1527,N_1242,N_1247);
xor U1528 (N_1528,In_827,N_402);
nor U1529 (N_1529,N_1003,N_1381);
nor U1530 (N_1530,N_1101,N_1331);
xor U1531 (N_1531,In_1474,N_1264);
or U1532 (N_1532,N_1354,N_943);
nand U1533 (N_1533,In_1627,N_483);
nand U1534 (N_1534,N_1326,N_1018);
nand U1535 (N_1535,N_204,In_522);
nor U1536 (N_1536,N_1222,N_887);
and U1537 (N_1537,N_23,N_1315);
or U1538 (N_1538,N_728,N_1118);
nor U1539 (N_1539,N_1261,N_29);
or U1540 (N_1540,N_839,N_1360);
nor U1541 (N_1541,N_618,N_256);
nand U1542 (N_1542,N_493,N_773);
nor U1543 (N_1543,N_1370,N_723);
and U1544 (N_1544,N_1190,N_1286);
and U1545 (N_1545,N_954,N_1145);
xnor U1546 (N_1546,N_227,In_1056);
nor U1547 (N_1547,In_281,N_1352);
xor U1548 (N_1548,In_720,N_1423);
nand U1549 (N_1549,N_1000,N_87);
xnor U1550 (N_1550,N_512,N_1439);
and U1551 (N_1551,N_991,N_994);
xnor U1552 (N_1552,In_1290,N_1122);
or U1553 (N_1553,N_1173,N_1435);
nand U1554 (N_1554,N_1092,N_334);
and U1555 (N_1555,N_1244,N_920);
xor U1556 (N_1556,N_1023,N_1213);
or U1557 (N_1557,N_817,N_966);
xor U1558 (N_1558,N_414,N_1289);
nand U1559 (N_1559,In_675,N_1267);
and U1560 (N_1560,N_701,N_1318);
and U1561 (N_1561,N_1175,In_155);
and U1562 (N_1562,N_1130,In_1126);
xor U1563 (N_1563,N_376,N_432);
nand U1564 (N_1564,N_852,In_322);
xnor U1565 (N_1565,In_1857,N_986);
nand U1566 (N_1566,In_582,N_752);
or U1567 (N_1567,N_1281,In_709);
xor U1568 (N_1568,N_1277,N_663);
or U1569 (N_1569,In_168,N_1428);
and U1570 (N_1570,N_407,N_1346);
xnor U1571 (N_1571,In_1130,In_903);
and U1572 (N_1572,N_699,In_943);
and U1573 (N_1573,N_1353,N_1290);
xor U1574 (N_1574,N_1068,N_1088);
nand U1575 (N_1575,N_1211,N_36);
nor U1576 (N_1576,N_1158,In_747);
xor U1577 (N_1577,N_1288,N_562);
or U1578 (N_1578,N_503,N_496);
nor U1579 (N_1579,In_167,In_1636);
xor U1580 (N_1580,N_1351,N_916);
nor U1581 (N_1581,N_1232,N_1357);
nand U1582 (N_1582,In_79,In_459);
or U1583 (N_1583,N_861,N_1382);
or U1584 (N_1584,N_1045,N_1380);
xnor U1585 (N_1585,In_636,N_1001);
nand U1586 (N_1586,N_1426,N_1401);
or U1587 (N_1587,N_851,N_1413);
xor U1588 (N_1588,In_547,N_1282);
nand U1589 (N_1589,N_1372,N_1198);
nor U1590 (N_1590,In_84,N_1416);
and U1591 (N_1591,In_958,N_953);
nand U1592 (N_1592,N_1397,In_307);
and U1593 (N_1593,N_1350,N_27);
xnor U1594 (N_1594,N_1291,N_1328);
nand U1595 (N_1595,N_1297,N_1116);
nor U1596 (N_1596,N_314,N_1366);
or U1597 (N_1597,N_1304,N_1307);
nand U1598 (N_1598,N_1274,N_1379);
nor U1599 (N_1599,N_1396,N_1182);
or U1600 (N_1600,N_1507,N_799);
and U1601 (N_1601,N_1485,N_1494);
nor U1602 (N_1602,N_1547,N_1454);
nand U1603 (N_1603,In_1587,N_1332);
or U1604 (N_1604,N_1552,N_1245);
nor U1605 (N_1605,N_647,N_1321);
nor U1606 (N_1606,N_1553,In_911);
nand U1607 (N_1607,N_1296,N_716);
xor U1608 (N_1608,N_1450,N_1472);
and U1609 (N_1609,In_201,N_207);
xor U1610 (N_1610,N_1592,N_1503);
nand U1611 (N_1611,N_1434,N_869);
or U1612 (N_1612,N_1476,N_1298);
nand U1613 (N_1613,N_1310,N_1169);
xnor U1614 (N_1614,N_511,N_616);
and U1615 (N_1615,N_1590,In_1123);
xnor U1616 (N_1616,N_1279,N_1166);
nor U1617 (N_1617,N_883,N_1493);
nor U1618 (N_1618,N_1599,N_988);
xnor U1619 (N_1619,N_1594,N_1207);
nor U1620 (N_1620,In_388,N_972);
xnor U1621 (N_1621,N_398,N_1410);
nand U1622 (N_1622,N_1181,N_1107);
or U1623 (N_1623,N_1394,N_1373);
nand U1624 (N_1624,N_1385,N_337);
and U1625 (N_1625,N_1474,N_653);
and U1626 (N_1626,N_655,N_1516);
xnor U1627 (N_1627,N_758,N_1456);
nand U1628 (N_1628,N_1447,N_1537);
xor U1629 (N_1629,N_1377,N_1202);
or U1630 (N_1630,N_1558,N_1515);
nor U1631 (N_1631,N_1526,In_338);
nand U1632 (N_1632,N_590,N_1389);
xnor U1633 (N_1633,N_1545,N_657);
nor U1634 (N_1634,N_1572,N_1319);
nand U1635 (N_1635,N_1530,N_1480);
nand U1636 (N_1636,N_1527,In_1458);
or U1637 (N_1637,N_1443,N_1249);
or U1638 (N_1638,N_1597,N_1473);
nor U1639 (N_1639,In_24,N_1533);
nor U1640 (N_1640,N_1057,N_1483);
and U1641 (N_1641,N_1303,In_1119);
and U1642 (N_1642,In_693,N_1591);
nand U1643 (N_1643,N_157,N_1581);
or U1644 (N_1644,N_1470,N_1570);
xor U1645 (N_1645,N_1523,N_1349);
and U1646 (N_1646,N_1544,N_1495);
nand U1647 (N_1647,N_1468,In_835);
nand U1648 (N_1648,In_1125,N_1324);
or U1649 (N_1649,N_1528,N_961);
or U1650 (N_1650,N_1334,N_230);
nor U1651 (N_1651,N_1024,N_1522);
or U1652 (N_1652,N_1398,In_1436);
and U1653 (N_1653,N_1189,N_837);
or U1654 (N_1654,N_1444,In_969);
or U1655 (N_1655,N_1535,N_1562);
nor U1656 (N_1656,N_144,N_353);
xor U1657 (N_1657,N_1458,N_1248);
nand U1658 (N_1658,N_1014,N_561);
nor U1659 (N_1659,In_1638,N_1498);
xnor U1660 (N_1660,In_325,N_1229);
nor U1661 (N_1661,N_909,N_1568);
and U1662 (N_1662,In_1668,In_90);
and U1663 (N_1663,N_1338,N_1448);
nor U1664 (N_1664,N_1546,N_1598);
and U1665 (N_1665,N_1025,In_143);
or U1666 (N_1666,N_1567,N_1460);
and U1667 (N_1667,N_1487,N_1301);
and U1668 (N_1668,N_1425,N_433);
nand U1669 (N_1669,N_1347,N_1376);
xor U1670 (N_1670,N_754,N_1459);
nand U1671 (N_1671,N_937,N_1238);
nand U1672 (N_1672,N_1540,N_1543);
nand U1673 (N_1673,In_271,N_1440);
and U1674 (N_1674,N_1463,N_1596);
xor U1675 (N_1675,N_1481,N_1066);
xnor U1676 (N_1676,N_387,N_558);
nor U1677 (N_1677,N_216,N_1240);
and U1678 (N_1678,N_1314,N_1510);
and U1679 (N_1679,N_484,N_1134);
nor U1680 (N_1680,N_1449,N_1210);
and U1681 (N_1681,N_921,N_1196);
xor U1682 (N_1682,N_158,N_1491);
or U1683 (N_1683,N_1455,N_1589);
nand U1684 (N_1684,N_1327,N_1358);
xnor U1685 (N_1685,N_1501,N_977);
or U1686 (N_1686,N_1560,N_1514);
or U1687 (N_1687,N_1519,N_1577);
xor U1688 (N_1688,N_487,N_1580);
nand U1689 (N_1689,In_1685,N_1084);
nand U1690 (N_1690,In_1400,N_1422);
nand U1691 (N_1691,N_1541,N_997);
and U1692 (N_1692,N_1569,N_1430);
or U1693 (N_1693,N_1407,N_1529);
xor U1694 (N_1694,N_1411,In_1274);
nand U1695 (N_1695,N_1511,N_1565);
and U1696 (N_1696,N_807,N_1072);
or U1697 (N_1697,N_1573,N_1588);
xnor U1698 (N_1698,N_1387,In_1803);
or U1699 (N_1699,N_840,N_1595);
xor U1700 (N_1700,N_1469,N_1388);
nor U1701 (N_1701,N_1016,N_1555);
nor U1702 (N_1702,N_1475,N_1551);
nand U1703 (N_1703,N_1178,N_1502);
and U1704 (N_1704,N_1585,N_340);
nor U1705 (N_1705,N_1156,In_768);
or U1706 (N_1706,N_1253,N_1427);
nor U1707 (N_1707,N_1039,N_1446);
nor U1708 (N_1708,In_60,In_1462);
nor U1709 (N_1709,N_1512,N_1464);
nor U1710 (N_1710,N_803,In_305);
nand U1711 (N_1711,N_1420,N_1564);
and U1712 (N_1712,N_1574,In_695);
and U1713 (N_1713,N_1525,N_1395);
and U1714 (N_1714,N_1484,N_1566);
or U1715 (N_1715,N_633,In_645);
and U1716 (N_1716,N_1445,In_1321);
nor U1717 (N_1717,N_1363,N_1172);
nand U1718 (N_1718,In_421,N_888);
xnor U1719 (N_1719,N_1489,N_1123);
nor U1720 (N_1720,N_1486,N_1374);
nand U1721 (N_1721,N_1273,In_1022);
nor U1722 (N_1722,N_1335,N_1539);
nor U1723 (N_1723,N_1471,N_1348);
xnor U1724 (N_1724,N_1500,N_1517);
and U1725 (N_1725,N_858,N_1452);
xor U1726 (N_1726,N_833,N_1343);
and U1727 (N_1727,N_1042,N_1520);
nor U1728 (N_1728,N_1400,N_1333);
nand U1729 (N_1729,N_1587,N_1532);
and U1730 (N_1730,N_1499,N_1408);
xnor U1731 (N_1731,In_1127,N_1513);
or U1732 (N_1732,N_1524,N_1223);
or U1733 (N_1733,N_1505,N_830);
or U1734 (N_1734,N_224,N_1345);
or U1735 (N_1735,In_1032,N_521);
or U1736 (N_1736,N_894,N_1550);
xnor U1737 (N_1737,In_1677,In_1320);
nand U1738 (N_1738,N_1402,N_1378);
xnor U1739 (N_1739,N_1339,N_1322);
xor U1740 (N_1740,N_1136,In_123);
and U1741 (N_1741,N_1506,N_1431);
xor U1742 (N_1742,N_1336,N_1451);
xor U1743 (N_1743,N_1571,N_1477);
xnor U1744 (N_1744,In_1495,N_319);
and U1745 (N_1745,N_1583,N_1466);
xnor U1746 (N_1746,N_1557,N_1341);
and U1747 (N_1747,N_1258,N_1436);
xnor U1748 (N_1748,N_1579,N_1216);
and U1749 (N_1749,N_847,In_1879);
or U1750 (N_1750,N_1518,N_1009);
and U1751 (N_1751,N_1461,N_1005);
and U1752 (N_1752,N_1429,N_1367);
or U1753 (N_1753,N_1325,N_683);
nand U1754 (N_1754,In_1444,N_1414);
xnor U1755 (N_1755,N_1160,N_1457);
xor U1756 (N_1756,N_1563,In_1795);
nand U1757 (N_1757,N_1554,N_1548);
nand U1758 (N_1758,N_1593,N_1415);
nand U1759 (N_1759,N_1479,N_979);
xor U1760 (N_1760,N_1674,N_1663);
nor U1761 (N_1761,N_1743,N_924);
and U1762 (N_1762,N_1584,N_1665);
nor U1763 (N_1763,N_1035,N_1651);
or U1764 (N_1764,N_1712,N_1640);
xor U1765 (N_1765,N_1680,N_1667);
nand U1766 (N_1766,N_1664,N_1654);
and U1767 (N_1767,N_1706,N_1613);
nand U1768 (N_1768,N_1684,N_95);
nand U1769 (N_1769,N_1497,N_1742);
nand U1770 (N_1770,N_1738,N_1627);
nor U1771 (N_1771,N_1731,N_1647);
or U1772 (N_1772,N_1693,N_1747);
nand U1773 (N_1773,N_1734,N_1126);
and U1774 (N_1774,N_1600,N_1619);
xnor U1775 (N_1775,N_1753,N_1636);
xor U1776 (N_1776,N_1670,N_1716);
and U1777 (N_1777,N_1362,N_1739);
or U1778 (N_1778,N_1531,In_1559);
nand U1779 (N_1779,N_1698,N_1614);
nor U1780 (N_1780,N_1749,N_1603);
or U1781 (N_1781,N_1650,In_1607);
nor U1782 (N_1782,N_1120,N_1658);
or U1783 (N_1783,N_1692,N_1714);
or U1784 (N_1784,N_1586,N_1642);
nand U1785 (N_1785,N_1631,N_1733);
nor U1786 (N_1786,N_1559,N_1390);
xor U1787 (N_1787,N_1724,N_1639);
and U1788 (N_1788,N_1621,N_1695);
or U1789 (N_1789,N_1715,N_1741);
xnor U1790 (N_1790,N_1672,N_1200);
or U1791 (N_1791,N_1453,In_62);
nand U1792 (N_1792,N_1646,N_1612);
or U1793 (N_1793,N_1732,N_1605);
nor U1794 (N_1794,N_1608,N_499);
xnor U1795 (N_1795,In_380,N_1276);
nor U1796 (N_1796,N_1656,N_1536);
nand U1797 (N_1797,N_1534,N_1635);
or U1798 (N_1798,N_1538,N_1678);
or U1799 (N_1799,N_1442,N_1607);
or U1800 (N_1800,N_1138,N_1637);
nor U1801 (N_1801,N_1710,N_454);
nor U1802 (N_1802,N_1660,N_1609);
nor U1803 (N_1803,N_1217,N_1689);
or U1804 (N_1804,N_1748,N_1683);
or U1805 (N_1805,N_1320,N_1750);
xnor U1806 (N_1806,N_1721,N_1628);
and U1807 (N_1807,In_1337,N_1725);
xor U1808 (N_1808,N_1029,N_1673);
xnor U1809 (N_1809,N_1634,N_1711);
nand U1810 (N_1810,N_1610,N_1709);
and U1811 (N_1811,N_1713,N_1729);
nand U1812 (N_1812,N_1438,N_1433);
and U1813 (N_1813,N_1576,In_610);
nand U1814 (N_1814,N_1685,N_1549);
or U1815 (N_1815,N_1611,N_1638);
nand U1816 (N_1816,N_1271,In_593);
and U1817 (N_1817,N_1467,N_1746);
or U1818 (N_1818,N_1655,N_1735);
and U1819 (N_1819,N_1726,N_1504);
nand U1820 (N_1820,N_1652,N_1705);
xnor U1821 (N_1821,N_1633,N_1625);
xnor U1822 (N_1822,N_1623,N_441);
xor U1823 (N_1823,N_1718,N_1492);
nor U1824 (N_1824,N_1694,N_1488);
nor U1825 (N_1825,N_1691,N_1542);
xor U1826 (N_1826,N_1582,N_1697);
and U1827 (N_1827,N_1622,N_1708);
or U1828 (N_1828,N_1701,N_587);
nor U1829 (N_1829,N_1418,N_1384);
nand U1830 (N_1830,N_1578,N_1044);
and U1831 (N_1831,N_1630,N_1490);
xor U1832 (N_1832,N_1690,N_1688);
xnor U1833 (N_1833,N_1671,N_1641);
or U1834 (N_1834,N_1645,N_239);
xnor U1835 (N_1835,N_1758,N_1626);
nor U1836 (N_1836,N_1653,N_1648);
nor U1837 (N_1837,N_1620,N_1759);
or U1838 (N_1838,N_1754,N_1666);
nor U1839 (N_1839,N_1668,N_1141);
nand U1840 (N_1840,N_1167,N_1681);
and U1841 (N_1841,N_1344,N_1720);
xor U1842 (N_1842,N_1657,N_1736);
and U1843 (N_1843,N_1131,N_1659);
or U1844 (N_1844,N_1727,In_743);
nand U1845 (N_1845,N_1371,N_1306);
and U1846 (N_1846,In_122,N_1755);
and U1847 (N_1847,N_1687,N_1737);
or U1848 (N_1848,In_1068,N_1703);
nand U1849 (N_1849,N_1556,N_355);
nand U1850 (N_1850,N_1740,N_1508);
and U1851 (N_1851,N_1616,N_1462);
nor U1852 (N_1852,N_1496,N_1717);
xor U1853 (N_1853,N_1679,N_1661);
xnor U1854 (N_1854,N_1602,N_1704);
nand U1855 (N_1855,N_1751,N_1618);
nand U1856 (N_1856,N_1601,N_1744);
or U1857 (N_1857,N_1707,N_1756);
nor U1858 (N_1858,N_1644,N_905);
or U1859 (N_1859,N_1020,N_520);
and U1860 (N_1860,N_1752,N_1745);
or U1861 (N_1861,N_1403,N_1662);
or U1862 (N_1862,N_1675,N_1757);
nand U1863 (N_1863,N_105,N_1730);
nand U1864 (N_1864,N_1686,N_1723);
and U1865 (N_1865,N_1561,N_1677);
nand U1866 (N_1866,N_1521,N_1696);
or U1867 (N_1867,N_1700,N_1629);
nor U1868 (N_1868,N_1478,N_1482);
nor U1869 (N_1869,N_1465,N_1617);
xor U1870 (N_1870,N_1669,N_1676);
xor U1871 (N_1871,N_1722,N_1509);
and U1872 (N_1872,N_1615,N_1643);
nor U1873 (N_1873,N_1441,N_1632);
xor U1874 (N_1874,N_1575,N_1606);
or U1875 (N_1875,N_1702,N_1649);
xnor U1876 (N_1876,N_1719,N_1624);
nor U1877 (N_1877,N_1604,N_1355);
xor U1878 (N_1878,N_1728,N_1682);
and U1879 (N_1879,N_1699,N_1412);
xnor U1880 (N_1880,N_1679,N_1508);
nand U1881 (N_1881,N_1344,N_1746);
xor U1882 (N_1882,In_610,N_1684);
or U1883 (N_1883,N_1675,In_743);
xnor U1884 (N_1884,N_1669,N_1538);
nor U1885 (N_1885,N_1687,N_1670);
or U1886 (N_1886,N_1674,N_1657);
nand U1887 (N_1887,N_1582,N_1497);
and U1888 (N_1888,N_1465,N_1616);
nand U1889 (N_1889,N_1344,N_1693);
nor U1890 (N_1890,N_1627,In_62);
or U1891 (N_1891,N_1749,In_1068);
nor U1892 (N_1892,N_1714,N_1742);
and U1893 (N_1893,N_454,N_1615);
xnor U1894 (N_1894,N_520,N_1636);
and U1895 (N_1895,N_1371,N_239);
or U1896 (N_1896,In_122,In_1068);
or U1897 (N_1897,N_1412,N_1708);
or U1898 (N_1898,N_1739,N_1710);
nand U1899 (N_1899,N_1674,N_1605);
nand U1900 (N_1900,N_1702,N_1742);
or U1901 (N_1901,N_1418,N_1680);
and U1902 (N_1902,N_1634,N_1691);
nor U1903 (N_1903,N_1689,N_454);
or U1904 (N_1904,N_1442,N_1616);
nand U1905 (N_1905,N_1418,N_95);
and U1906 (N_1906,N_1634,N_1743);
nor U1907 (N_1907,N_1717,In_122);
or U1908 (N_1908,N_1671,N_1035);
or U1909 (N_1909,N_1695,N_1747);
nand U1910 (N_1910,N_1618,N_1649);
and U1911 (N_1911,N_1700,N_1719);
or U1912 (N_1912,N_1752,N_1750);
and U1913 (N_1913,In_610,N_1044);
or U1914 (N_1914,N_1734,N_1667);
nand U1915 (N_1915,N_1675,N_1549);
or U1916 (N_1916,N_454,N_1713);
nor U1917 (N_1917,N_1531,N_1750);
xnor U1918 (N_1918,N_1630,N_1613);
nand U1919 (N_1919,N_1658,N_1600);
xnor U1920 (N_1920,N_1792,N_1763);
nor U1921 (N_1921,N_1908,N_1832);
nor U1922 (N_1922,N_1807,N_1840);
nand U1923 (N_1923,N_1827,N_1876);
and U1924 (N_1924,N_1914,N_1772);
nand U1925 (N_1925,N_1859,N_1773);
xnor U1926 (N_1926,N_1852,N_1764);
nor U1927 (N_1927,N_1879,N_1891);
nor U1928 (N_1928,N_1873,N_1881);
nand U1929 (N_1929,N_1819,N_1779);
nor U1930 (N_1930,N_1865,N_1886);
nor U1931 (N_1931,N_1877,N_1902);
nor U1932 (N_1932,N_1861,N_1871);
xnor U1933 (N_1933,N_1862,N_1836);
or U1934 (N_1934,N_1813,N_1849);
xnor U1935 (N_1935,N_1899,N_1817);
or U1936 (N_1936,N_1889,N_1794);
xnor U1937 (N_1937,N_1782,N_1787);
or U1938 (N_1938,N_1805,N_1784);
or U1939 (N_1939,N_1913,N_1896);
nor U1940 (N_1940,N_1834,N_1780);
xor U1941 (N_1941,N_1766,N_1903);
nor U1942 (N_1942,N_1797,N_1838);
nand U1943 (N_1943,N_1863,N_1761);
and U1944 (N_1944,N_1848,N_1833);
or U1945 (N_1945,N_1812,N_1919);
or U1946 (N_1946,N_1905,N_1882);
nor U1947 (N_1947,N_1771,N_1781);
or U1948 (N_1948,N_1866,N_1769);
nand U1949 (N_1949,N_1799,N_1770);
or U1950 (N_1950,N_1897,N_1808);
xor U1951 (N_1951,N_1904,N_1785);
or U1952 (N_1952,N_1850,N_1890);
and U1953 (N_1953,N_1801,N_1847);
nor U1954 (N_1954,N_1822,N_1884);
nand U1955 (N_1955,N_1893,N_1892);
nor U1956 (N_1956,N_1906,N_1762);
nand U1957 (N_1957,N_1790,N_1844);
xor U1958 (N_1958,N_1845,N_1869);
nor U1959 (N_1959,N_1831,N_1851);
or U1960 (N_1960,N_1900,N_1868);
nand U1961 (N_1961,N_1765,N_1880);
nor U1962 (N_1962,N_1802,N_1870);
xnor U1963 (N_1963,N_1835,N_1867);
nor U1964 (N_1964,N_1774,N_1778);
nand U1965 (N_1965,N_1918,N_1775);
or U1966 (N_1966,N_1909,N_1818);
nand U1967 (N_1967,N_1795,N_1768);
nor U1968 (N_1968,N_1894,N_1796);
xor U1969 (N_1969,N_1789,N_1830);
nor U1970 (N_1970,N_1916,N_1826);
nor U1971 (N_1971,N_1878,N_1917);
nand U1972 (N_1972,N_1824,N_1791);
and U1973 (N_1973,N_1829,N_1872);
nand U1974 (N_1974,N_1806,N_1901);
or U1975 (N_1975,N_1839,N_1842);
nand U1976 (N_1976,N_1816,N_1883);
nor U1977 (N_1977,N_1912,N_1810);
xor U1978 (N_1978,N_1858,N_1887);
nor U1979 (N_1979,N_1895,N_1767);
nor U1980 (N_1980,N_1854,N_1804);
nand U1981 (N_1981,N_1800,N_1864);
xor U1982 (N_1982,N_1898,N_1788);
or U1983 (N_1983,N_1793,N_1885);
and U1984 (N_1984,N_1910,N_1777);
nor U1985 (N_1985,N_1875,N_1821);
and U1986 (N_1986,N_1786,N_1837);
nand U1987 (N_1987,N_1855,N_1776);
and U1988 (N_1988,N_1815,N_1798);
xor U1989 (N_1989,N_1843,N_1915);
xnor U1990 (N_1990,N_1760,N_1888);
nor U1991 (N_1991,N_1825,N_1783);
xor U1992 (N_1992,N_1907,N_1853);
nand U1993 (N_1993,N_1856,N_1803);
nand U1994 (N_1994,N_1809,N_1860);
or U1995 (N_1995,N_1811,N_1857);
and U1996 (N_1996,N_1828,N_1823);
xnor U1997 (N_1997,N_1820,N_1911);
nand U1998 (N_1998,N_1841,N_1874);
xor U1999 (N_1999,N_1814,N_1846);
and U2000 (N_2000,N_1866,N_1842);
and U2001 (N_2001,N_1902,N_1889);
nor U2002 (N_2002,N_1760,N_1777);
and U2003 (N_2003,N_1881,N_1784);
nor U2004 (N_2004,N_1845,N_1794);
xor U2005 (N_2005,N_1876,N_1767);
or U2006 (N_2006,N_1852,N_1913);
or U2007 (N_2007,N_1858,N_1859);
or U2008 (N_2008,N_1884,N_1799);
nor U2009 (N_2009,N_1890,N_1762);
and U2010 (N_2010,N_1858,N_1908);
or U2011 (N_2011,N_1766,N_1880);
nor U2012 (N_2012,N_1893,N_1910);
nor U2013 (N_2013,N_1914,N_1786);
nor U2014 (N_2014,N_1858,N_1867);
nand U2015 (N_2015,N_1836,N_1767);
and U2016 (N_2016,N_1851,N_1839);
nor U2017 (N_2017,N_1909,N_1793);
xor U2018 (N_2018,N_1810,N_1814);
and U2019 (N_2019,N_1807,N_1805);
nor U2020 (N_2020,N_1866,N_1790);
or U2021 (N_2021,N_1777,N_1835);
xnor U2022 (N_2022,N_1767,N_1774);
nor U2023 (N_2023,N_1798,N_1768);
and U2024 (N_2024,N_1913,N_1844);
nand U2025 (N_2025,N_1820,N_1898);
nand U2026 (N_2026,N_1910,N_1901);
or U2027 (N_2027,N_1814,N_1767);
and U2028 (N_2028,N_1881,N_1795);
and U2029 (N_2029,N_1884,N_1762);
xor U2030 (N_2030,N_1846,N_1779);
nor U2031 (N_2031,N_1893,N_1828);
nand U2032 (N_2032,N_1868,N_1800);
and U2033 (N_2033,N_1773,N_1805);
nor U2034 (N_2034,N_1769,N_1876);
nand U2035 (N_2035,N_1873,N_1899);
xnor U2036 (N_2036,N_1911,N_1834);
nor U2037 (N_2037,N_1809,N_1834);
xnor U2038 (N_2038,N_1892,N_1771);
and U2039 (N_2039,N_1826,N_1807);
xor U2040 (N_2040,N_1884,N_1856);
and U2041 (N_2041,N_1764,N_1797);
xnor U2042 (N_2042,N_1814,N_1872);
nor U2043 (N_2043,N_1898,N_1799);
or U2044 (N_2044,N_1777,N_1815);
xor U2045 (N_2045,N_1867,N_1771);
nand U2046 (N_2046,N_1819,N_1808);
and U2047 (N_2047,N_1805,N_1863);
and U2048 (N_2048,N_1834,N_1872);
xor U2049 (N_2049,N_1861,N_1832);
nor U2050 (N_2050,N_1814,N_1837);
nor U2051 (N_2051,N_1800,N_1794);
and U2052 (N_2052,N_1846,N_1870);
or U2053 (N_2053,N_1845,N_1895);
or U2054 (N_2054,N_1843,N_1773);
or U2055 (N_2055,N_1861,N_1801);
xnor U2056 (N_2056,N_1896,N_1832);
or U2057 (N_2057,N_1792,N_1918);
nand U2058 (N_2058,N_1846,N_1777);
xor U2059 (N_2059,N_1880,N_1858);
or U2060 (N_2060,N_1834,N_1918);
nor U2061 (N_2061,N_1788,N_1860);
or U2062 (N_2062,N_1915,N_1771);
or U2063 (N_2063,N_1867,N_1788);
and U2064 (N_2064,N_1837,N_1900);
or U2065 (N_2065,N_1815,N_1766);
nand U2066 (N_2066,N_1880,N_1813);
nand U2067 (N_2067,N_1772,N_1768);
nor U2068 (N_2068,N_1813,N_1797);
or U2069 (N_2069,N_1842,N_1790);
or U2070 (N_2070,N_1887,N_1826);
or U2071 (N_2071,N_1763,N_1779);
xnor U2072 (N_2072,N_1779,N_1823);
xnor U2073 (N_2073,N_1847,N_1795);
nand U2074 (N_2074,N_1890,N_1866);
nand U2075 (N_2075,N_1906,N_1772);
or U2076 (N_2076,N_1896,N_1905);
xnor U2077 (N_2077,N_1784,N_1793);
nand U2078 (N_2078,N_1914,N_1915);
or U2079 (N_2079,N_1792,N_1838);
nor U2080 (N_2080,N_2044,N_1998);
nor U2081 (N_2081,N_1942,N_2065);
nor U2082 (N_2082,N_1925,N_1964);
nand U2083 (N_2083,N_1930,N_2056);
nor U2084 (N_2084,N_1971,N_1940);
nand U2085 (N_2085,N_1977,N_1986);
and U2086 (N_2086,N_2028,N_1950);
and U2087 (N_2087,N_1934,N_1980);
nand U2088 (N_2088,N_1999,N_1962);
or U2089 (N_2089,N_1988,N_2018);
or U2090 (N_2090,N_2071,N_2047);
nand U2091 (N_2091,N_2051,N_1939);
nor U2092 (N_2092,N_1961,N_1973);
xnor U2093 (N_2093,N_1927,N_2050);
nor U2094 (N_2094,N_1920,N_2068);
and U2095 (N_2095,N_1926,N_1997);
and U2096 (N_2096,N_1929,N_2003);
nor U2097 (N_2097,N_2064,N_2045);
nor U2098 (N_2098,N_2013,N_2029);
xor U2099 (N_2099,N_1921,N_1969);
xnor U2100 (N_2100,N_1975,N_2053);
or U2101 (N_2101,N_2076,N_1978);
nor U2102 (N_2102,N_1953,N_2016);
nor U2103 (N_2103,N_1923,N_1968);
and U2104 (N_2104,N_1957,N_1935);
nand U2105 (N_2105,N_2033,N_1965);
or U2106 (N_2106,N_2000,N_2059);
nor U2107 (N_2107,N_1931,N_2021);
nor U2108 (N_2108,N_2061,N_2011);
xor U2109 (N_2109,N_1944,N_1958);
and U2110 (N_2110,N_2046,N_2042);
nand U2111 (N_2111,N_2075,N_2009);
or U2112 (N_2112,N_2077,N_2031);
nand U2113 (N_2113,N_1992,N_2069);
or U2114 (N_2114,N_2060,N_2073);
nor U2115 (N_2115,N_2007,N_2058);
xnor U2116 (N_2116,N_2037,N_1955);
or U2117 (N_2117,N_1933,N_1946);
xor U2118 (N_2118,N_1943,N_2025);
and U2119 (N_2119,N_2019,N_1981);
nor U2120 (N_2120,N_2078,N_2067);
xor U2121 (N_2121,N_2072,N_1982);
and U2122 (N_2122,N_1959,N_1970);
and U2123 (N_2123,N_1996,N_2020);
or U2124 (N_2124,N_1938,N_2049);
and U2125 (N_2125,N_1994,N_1928);
xnor U2126 (N_2126,N_1967,N_1932);
and U2127 (N_2127,N_1924,N_2027);
nand U2128 (N_2128,N_2057,N_2017);
nand U2129 (N_2129,N_1945,N_1966);
xor U2130 (N_2130,N_2054,N_2063);
and U2131 (N_2131,N_1991,N_2038);
xor U2132 (N_2132,N_1947,N_2062);
and U2133 (N_2133,N_1995,N_2008);
nand U2134 (N_2134,N_1960,N_2022);
nand U2135 (N_2135,N_1993,N_1983);
and U2136 (N_2136,N_1937,N_2070);
nand U2137 (N_2137,N_2014,N_2032);
nor U2138 (N_2138,N_1985,N_2023);
nor U2139 (N_2139,N_2043,N_2074);
xnor U2140 (N_2140,N_1974,N_2012);
and U2141 (N_2141,N_2040,N_2026);
nand U2142 (N_2142,N_2035,N_1972);
and U2143 (N_2143,N_2052,N_1951);
and U2144 (N_2144,N_2002,N_2041);
nor U2145 (N_2145,N_2034,N_2004);
and U2146 (N_2146,N_2066,N_2055);
nand U2147 (N_2147,N_1990,N_2024);
or U2148 (N_2148,N_2048,N_1963);
nand U2149 (N_2149,N_2079,N_2001);
nand U2150 (N_2150,N_2006,N_2039);
nand U2151 (N_2151,N_2030,N_2036);
nor U2152 (N_2152,N_1984,N_1948);
and U2153 (N_2153,N_1952,N_1987);
nand U2154 (N_2154,N_1949,N_1956);
or U2155 (N_2155,N_1976,N_2005);
nor U2156 (N_2156,N_1979,N_1936);
or U2157 (N_2157,N_2010,N_1954);
nand U2158 (N_2158,N_1989,N_1941);
or U2159 (N_2159,N_2015,N_1922);
and U2160 (N_2160,N_1948,N_1985);
or U2161 (N_2161,N_1979,N_2051);
or U2162 (N_2162,N_1975,N_1964);
xor U2163 (N_2163,N_1968,N_2018);
nand U2164 (N_2164,N_1933,N_2073);
nand U2165 (N_2165,N_2009,N_2022);
nand U2166 (N_2166,N_2053,N_1990);
or U2167 (N_2167,N_2021,N_1993);
nor U2168 (N_2168,N_1936,N_1922);
nor U2169 (N_2169,N_2027,N_1974);
and U2170 (N_2170,N_2065,N_1933);
xor U2171 (N_2171,N_2008,N_1954);
nor U2172 (N_2172,N_2052,N_1921);
nor U2173 (N_2173,N_2036,N_1965);
or U2174 (N_2174,N_2024,N_2054);
nor U2175 (N_2175,N_1952,N_1948);
and U2176 (N_2176,N_2057,N_2077);
and U2177 (N_2177,N_2047,N_1973);
nor U2178 (N_2178,N_2066,N_2053);
and U2179 (N_2179,N_1974,N_1943);
or U2180 (N_2180,N_2071,N_1970);
xor U2181 (N_2181,N_1979,N_2063);
nand U2182 (N_2182,N_1945,N_2057);
and U2183 (N_2183,N_1965,N_2049);
and U2184 (N_2184,N_2054,N_1970);
nor U2185 (N_2185,N_2068,N_2047);
xor U2186 (N_2186,N_2039,N_2058);
xnor U2187 (N_2187,N_1983,N_1943);
nor U2188 (N_2188,N_2042,N_2008);
nand U2189 (N_2189,N_2005,N_1936);
nand U2190 (N_2190,N_2010,N_1973);
nor U2191 (N_2191,N_2078,N_2012);
and U2192 (N_2192,N_2018,N_2021);
nand U2193 (N_2193,N_1969,N_1946);
nand U2194 (N_2194,N_1943,N_1988);
xnor U2195 (N_2195,N_1978,N_2028);
and U2196 (N_2196,N_2042,N_2076);
and U2197 (N_2197,N_2048,N_2045);
or U2198 (N_2198,N_1987,N_2033);
nor U2199 (N_2199,N_2029,N_1958);
nor U2200 (N_2200,N_1935,N_1980);
or U2201 (N_2201,N_1977,N_2009);
xnor U2202 (N_2202,N_1986,N_1966);
nand U2203 (N_2203,N_1922,N_2018);
xor U2204 (N_2204,N_2013,N_2036);
nor U2205 (N_2205,N_2015,N_1948);
nand U2206 (N_2206,N_2017,N_2016);
and U2207 (N_2207,N_1994,N_1976);
xnor U2208 (N_2208,N_1991,N_1955);
nor U2209 (N_2209,N_1972,N_2009);
nand U2210 (N_2210,N_1996,N_1953);
or U2211 (N_2211,N_1987,N_1947);
or U2212 (N_2212,N_2014,N_1926);
and U2213 (N_2213,N_1972,N_2069);
and U2214 (N_2214,N_2018,N_2036);
nand U2215 (N_2215,N_2007,N_2018);
nor U2216 (N_2216,N_2037,N_1928);
or U2217 (N_2217,N_2008,N_1986);
or U2218 (N_2218,N_1975,N_1965);
or U2219 (N_2219,N_1931,N_2053);
and U2220 (N_2220,N_2049,N_2046);
xnor U2221 (N_2221,N_1958,N_2025);
xnor U2222 (N_2222,N_2030,N_2068);
nand U2223 (N_2223,N_2045,N_2073);
or U2224 (N_2224,N_2021,N_2005);
nand U2225 (N_2225,N_1926,N_2030);
xor U2226 (N_2226,N_1985,N_2059);
nand U2227 (N_2227,N_2022,N_1957);
nor U2228 (N_2228,N_2015,N_2033);
and U2229 (N_2229,N_2037,N_2040);
or U2230 (N_2230,N_1931,N_1965);
xor U2231 (N_2231,N_2064,N_2052);
or U2232 (N_2232,N_1957,N_1929);
nor U2233 (N_2233,N_2048,N_2014);
and U2234 (N_2234,N_2079,N_2005);
nand U2235 (N_2235,N_1931,N_2055);
and U2236 (N_2236,N_1931,N_1951);
and U2237 (N_2237,N_2051,N_2030);
xnor U2238 (N_2238,N_2028,N_1975);
nand U2239 (N_2239,N_2002,N_1931);
nor U2240 (N_2240,N_2117,N_2239);
or U2241 (N_2241,N_2169,N_2108);
or U2242 (N_2242,N_2198,N_2188);
and U2243 (N_2243,N_2204,N_2110);
or U2244 (N_2244,N_2091,N_2154);
or U2245 (N_2245,N_2084,N_2214);
xor U2246 (N_2246,N_2185,N_2109);
nor U2247 (N_2247,N_2162,N_2202);
nand U2248 (N_2248,N_2149,N_2176);
xnor U2249 (N_2249,N_2163,N_2126);
and U2250 (N_2250,N_2199,N_2222);
nor U2251 (N_2251,N_2205,N_2148);
or U2252 (N_2252,N_2226,N_2127);
or U2253 (N_2253,N_2229,N_2141);
and U2254 (N_2254,N_2088,N_2100);
and U2255 (N_2255,N_2219,N_2147);
nor U2256 (N_2256,N_2080,N_2167);
nor U2257 (N_2257,N_2142,N_2178);
nor U2258 (N_2258,N_2216,N_2232);
nor U2259 (N_2259,N_2129,N_2112);
and U2260 (N_2260,N_2119,N_2128);
nand U2261 (N_2261,N_2140,N_2101);
or U2262 (N_2262,N_2168,N_2209);
and U2263 (N_2263,N_2238,N_2134);
or U2264 (N_2264,N_2139,N_2131);
nor U2265 (N_2265,N_2107,N_2184);
or U2266 (N_2266,N_2113,N_2160);
nor U2267 (N_2267,N_2106,N_2200);
nor U2268 (N_2268,N_2193,N_2146);
and U2269 (N_2269,N_2187,N_2118);
nor U2270 (N_2270,N_2130,N_2235);
xor U2271 (N_2271,N_2081,N_2208);
and U2272 (N_2272,N_2190,N_2236);
nand U2273 (N_2273,N_2159,N_2195);
nand U2274 (N_2274,N_2221,N_2179);
nor U2275 (N_2275,N_2172,N_2121);
or U2276 (N_2276,N_2098,N_2231);
nand U2277 (N_2277,N_2180,N_2153);
xor U2278 (N_2278,N_2201,N_2150);
xnor U2279 (N_2279,N_2207,N_2224);
nor U2280 (N_2280,N_2124,N_2152);
or U2281 (N_2281,N_2234,N_2095);
nand U2282 (N_2282,N_2197,N_2096);
nand U2283 (N_2283,N_2237,N_2083);
or U2284 (N_2284,N_2155,N_2133);
and U2285 (N_2285,N_2173,N_2090);
xnor U2286 (N_2286,N_2136,N_2210);
nor U2287 (N_2287,N_2123,N_2186);
or U2288 (N_2288,N_2227,N_2099);
xnor U2289 (N_2289,N_2217,N_2138);
nand U2290 (N_2290,N_2104,N_2203);
nor U2291 (N_2291,N_2143,N_2191);
or U2292 (N_2292,N_2087,N_2206);
or U2293 (N_2293,N_2102,N_2223);
nand U2294 (N_2294,N_2183,N_2114);
nor U2295 (N_2295,N_2165,N_2228);
or U2296 (N_2296,N_2158,N_2111);
or U2297 (N_2297,N_2082,N_2092);
or U2298 (N_2298,N_2103,N_2174);
or U2299 (N_2299,N_2220,N_2175);
nand U2300 (N_2300,N_2120,N_2156);
or U2301 (N_2301,N_2144,N_2218);
or U2302 (N_2302,N_2097,N_2233);
and U2303 (N_2303,N_2089,N_2105);
and U2304 (N_2304,N_2211,N_2225);
nor U2305 (N_2305,N_2170,N_2094);
or U2306 (N_2306,N_2116,N_2115);
nor U2307 (N_2307,N_2166,N_2151);
or U2308 (N_2308,N_2157,N_2164);
or U2309 (N_2309,N_2125,N_2132);
xor U2310 (N_2310,N_2189,N_2215);
or U2311 (N_2311,N_2196,N_2177);
xnor U2312 (N_2312,N_2212,N_2171);
nor U2313 (N_2313,N_2230,N_2194);
or U2314 (N_2314,N_2161,N_2085);
nor U2315 (N_2315,N_2181,N_2192);
or U2316 (N_2316,N_2145,N_2086);
and U2317 (N_2317,N_2135,N_2182);
and U2318 (N_2318,N_2122,N_2137);
and U2319 (N_2319,N_2093,N_2213);
or U2320 (N_2320,N_2131,N_2097);
and U2321 (N_2321,N_2159,N_2105);
nand U2322 (N_2322,N_2160,N_2194);
nand U2323 (N_2323,N_2114,N_2133);
or U2324 (N_2324,N_2129,N_2174);
xnor U2325 (N_2325,N_2084,N_2212);
nor U2326 (N_2326,N_2089,N_2148);
xnor U2327 (N_2327,N_2139,N_2186);
nand U2328 (N_2328,N_2189,N_2170);
and U2329 (N_2329,N_2158,N_2163);
or U2330 (N_2330,N_2175,N_2117);
xor U2331 (N_2331,N_2185,N_2234);
and U2332 (N_2332,N_2151,N_2199);
nand U2333 (N_2333,N_2103,N_2226);
and U2334 (N_2334,N_2083,N_2096);
nor U2335 (N_2335,N_2145,N_2190);
nor U2336 (N_2336,N_2201,N_2184);
nand U2337 (N_2337,N_2186,N_2159);
and U2338 (N_2338,N_2140,N_2164);
xor U2339 (N_2339,N_2189,N_2160);
or U2340 (N_2340,N_2130,N_2205);
nand U2341 (N_2341,N_2219,N_2152);
nor U2342 (N_2342,N_2134,N_2188);
xnor U2343 (N_2343,N_2115,N_2104);
or U2344 (N_2344,N_2216,N_2116);
nor U2345 (N_2345,N_2129,N_2184);
nand U2346 (N_2346,N_2221,N_2188);
or U2347 (N_2347,N_2213,N_2082);
nand U2348 (N_2348,N_2237,N_2112);
xnor U2349 (N_2349,N_2223,N_2174);
nor U2350 (N_2350,N_2148,N_2161);
nand U2351 (N_2351,N_2177,N_2084);
xnor U2352 (N_2352,N_2155,N_2159);
nand U2353 (N_2353,N_2189,N_2208);
and U2354 (N_2354,N_2179,N_2152);
or U2355 (N_2355,N_2189,N_2205);
nand U2356 (N_2356,N_2210,N_2086);
nor U2357 (N_2357,N_2164,N_2130);
xnor U2358 (N_2358,N_2167,N_2230);
nor U2359 (N_2359,N_2209,N_2110);
nor U2360 (N_2360,N_2198,N_2081);
and U2361 (N_2361,N_2151,N_2093);
or U2362 (N_2362,N_2081,N_2124);
and U2363 (N_2363,N_2117,N_2223);
nand U2364 (N_2364,N_2197,N_2201);
or U2365 (N_2365,N_2100,N_2234);
and U2366 (N_2366,N_2125,N_2086);
and U2367 (N_2367,N_2083,N_2203);
xnor U2368 (N_2368,N_2119,N_2220);
xnor U2369 (N_2369,N_2235,N_2126);
and U2370 (N_2370,N_2176,N_2207);
xnor U2371 (N_2371,N_2131,N_2092);
xor U2372 (N_2372,N_2177,N_2140);
nand U2373 (N_2373,N_2206,N_2121);
nand U2374 (N_2374,N_2127,N_2148);
nand U2375 (N_2375,N_2145,N_2112);
nand U2376 (N_2376,N_2088,N_2130);
nand U2377 (N_2377,N_2222,N_2192);
nor U2378 (N_2378,N_2159,N_2178);
nor U2379 (N_2379,N_2235,N_2084);
nor U2380 (N_2380,N_2089,N_2137);
nor U2381 (N_2381,N_2165,N_2232);
nand U2382 (N_2382,N_2111,N_2117);
and U2383 (N_2383,N_2181,N_2187);
nor U2384 (N_2384,N_2187,N_2183);
or U2385 (N_2385,N_2157,N_2116);
nand U2386 (N_2386,N_2119,N_2165);
or U2387 (N_2387,N_2089,N_2115);
xnor U2388 (N_2388,N_2125,N_2182);
or U2389 (N_2389,N_2127,N_2121);
xnor U2390 (N_2390,N_2099,N_2129);
nor U2391 (N_2391,N_2229,N_2139);
or U2392 (N_2392,N_2134,N_2173);
and U2393 (N_2393,N_2115,N_2157);
nand U2394 (N_2394,N_2097,N_2095);
xnor U2395 (N_2395,N_2213,N_2198);
and U2396 (N_2396,N_2080,N_2149);
nor U2397 (N_2397,N_2137,N_2191);
xor U2398 (N_2398,N_2226,N_2161);
and U2399 (N_2399,N_2199,N_2193);
nor U2400 (N_2400,N_2296,N_2317);
nand U2401 (N_2401,N_2246,N_2272);
nand U2402 (N_2402,N_2281,N_2319);
xor U2403 (N_2403,N_2352,N_2341);
xnor U2404 (N_2404,N_2273,N_2282);
or U2405 (N_2405,N_2264,N_2315);
nand U2406 (N_2406,N_2338,N_2265);
or U2407 (N_2407,N_2335,N_2377);
xnor U2408 (N_2408,N_2367,N_2299);
nor U2409 (N_2409,N_2386,N_2244);
xnor U2410 (N_2410,N_2275,N_2388);
nand U2411 (N_2411,N_2358,N_2331);
and U2412 (N_2412,N_2261,N_2340);
nor U2413 (N_2413,N_2287,N_2277);
nand U2414 (N_2414,N_2314,N_2267);
nand U2415 (N_2415,N_2361,N_2344);
nand U2416 (N_2416,N_2284,N_2389);
or U2417 (N_2417,N_2330,N_2271);
xor U2418 (N_2418,N_2280,N_2398);
nand U2419 (N_2419,N_2323,N_2247);
xor U2420 (N_2420,N_2321,N_2392);
nand U2421 (N_2421,N_2337,N_2380);
and U2422 (N_2422,N_2241,N_2290);
nand U2423 (N_2423,N_2351,N_2240);
nor U2424 (N_2424,N_2374,N_2257);
or U2425 (N_2425,N_2366,N_2256);
nand U2426 (N_2426,N_2322,N_2385);
or U2427 (N_2427,N_2268,N_2378);
or U2428 (N_2428,N_2263,N_2288);
nand U2429 (N_2429,N_2260,N_2350);
xnor U2430 (N_2430,N_2276,N_2245);
or U2431 (N_2431,N_2312,N_2253);
xor U2432 (N_2432,N_2254,N_2311);
xnor U2433 (N_2433,N_2250,N_2307);
nand U2434 (N_2434,N_2370,N_2309);
or U2435 (N_2435,N_2302,N_2304);
nand U2436 (N_2436,N_2397,N_2318);
nand U2437 (N_2437,N_2286,N_2376);
or U2438 (N_2438,N_2291,N_2258);
nand U2439 (N_2439,N_2362,N_2279);
nand U2440 (N_2440,N_2289,N_2363);
nor U2441 (N_2441,N_2334,N_2354);
xor U2442 (N_2442,N_2305,N_2310);
and U2443 (N_2443,N_2262,N_2255);
or U2444 (N_2444,N_2249,N_2266);
nor U2445 (N_2445,N_2274,N_2359);
nand U2446 (N_2446,N_2298,N_2329);
or U2447 (N_2447,N_2399,N_2332);
and U2448 (N_2448,N_2364,N_2259);
and U2449 (N_2449,N_2357,N_2379);
nor U2450 (N_2450,N_2303,N_2383);
nand U2451 (N_2451,N_2285,N_2269);
xnor U2452 (N_2452,N_2333,N_2300);
nand U2453 (N_2453,N_2356,N_2375);
xnor U2454 (N_2454,N_2393,N_2252);
and U2455 (N_2455,N_2368,N_2297);
or U2456 (N_2456,N_2390,N_2327);
nand U2457 (N_2457,N_2355,N_2243);
xor U2458 (N_2458,N_2345,N_2396);
xor U2459 (N_2459,N_2308,N_2371);
xor U2460 (N_2460,N_2292,N_2369);
nor U2461 (N_2461,N_2293,N_2295);
or U2462 (N_2462,N_2339,N_2326);
nor U2463 (N_2463,N_2336,N_2248);
and U2464 (N_2464,N_2360,N_2320);
nand U2465 (N_2465,N_2251,N_2353);
and U2466 (N_2466,N_2342,N_2343);
or U2467 (N_2467,N_2384,N_2301);
nor U2468 (N_2468,N_2325,N_2328);
nand U2469 (N_2469,N_2395,N_2382);
nor U2470 (N_2470,N_2313,N_2306);
or U2471 (N_2471,N_2294,N_2391);
or U2472 (N_2472,N_2365,N_2270);
or U2473 (N_2473,N_2372,N_2381);
xor U2474 (N_2474,N_2348,N_2242);
or U2475 (N_2475,N_2316,N_2324);
nand U2476 (N_2476,N_2278,N_2387);
xnor U2477 (N_2477,N_2349,N_2346);
or U2478 (N_2478,N_2394,N_2283);
and U2479 (N_2479,N_2373,N_2347);
xor U2480 (N_2480,N_2333,N_2315);
and U2481 (N_2481,N_2384,N_2352);
nor U2482 (N_2482,N_2317,N_2356);
xnor U2483 (N_2483,N_2324,N_2368);
or U2484 (N_2484,N_2240,N_2243);
xnor U2485 (N_2485,N_2246,N_2243);
or U2486 (N_2486,N_2396,N_2328);
nand U2487 (N_2487,N_2276,N_2345);
and U2488 (N_2488,N_2321,N_2268);
and U2489 (N_2489,N_2324,N_2349);
xnor U2490 (N_2490,N_2282,N_2320);
and U2491 (N_2491,N_2371,N_2267);
nand U2492 (N_2492,N_2247,N_2330);
or U2493 (N_2493,N_2313,N_2333);
and U2494 (N_2494,N_2284,N_2275);
xnor U2495 (N_2495,N_2286,N_2353);
xor U2496 (N_2496,N_2292,N_2382);
or U2497 (N_2497,N_2328,N_2257);
nand U2498 (N_2498,N_2365,N_2345);
xor U2499 (N_2499,N_2278,N_2307);
nor U2500 (N_2500,N_2293,N_2351);
xnor U2501 (N_2501,N_2252,N_2300);
nor U2502 (N_2502,N_2377,N_2380);
nand U2503 (N_2503,N_2354,N_2304);
nand U2504 (N_2504,N_2351,N_2267);
xnor U2505 (N_2505,N_2243,N_2337);
nor U2506 (N_2506,N_2240,N_2245);
and U2507 (N_2507,N_2269,N_2268);
nand U2508 (N_2508,N_2282,N_2245);
nand U2509 (N_2509,N_2290,N_2369);
or U2510 (N_2510,N_2299,N_2348);
xor U2511 (N_2511,N_2386,N_2301);
xnor U2512 (N_2512,N_2323,N_2383);
nor U2513 (N_2513,N_2300,N_2271);
nor U2514 (N_2514,N_2255,N_2264);
nand U2515 (N_2515,N_2304,N_2359);
and U2516 (N_2516,N_2385,N_2240);
nor U2517 (N_2517,N_2254,N_2276);
and U2518 (N_2518,N_2361,N_2251);
nand U2519 (N_2519,N_2383,N_2336);
or U2520 (N_2520,N_2350,N_2343);
nand U2521 (N_2521,N_2352,N_2361);
and U2522 (N_2522,N_2251,N_2387);
xnor U2523 (N_2523,N_2273,N_2332);
nor U2524 (N_2524,N_2305,N_2250);
nor U2525 (N_2525,N_2279,N_2322);
and U2526 (N_2526,N_2369,N_2240);
nand U2527 (N_2527,N_2297,N_2381);
and U2528 (N_2528,N_2323,N_2277);
xor U2529 (N_2529,N_2341,N_2344);
xor U2530 (N_2530,N_2322,N_2388);
xnor U2531 (N_2531,N_2249,N_2396);
and U2532 (N_2532,N_2254,N_2351);
and U2533 (N_2533,N_2397,N_2251);
or U2534 (N_2534,N_2324,N_2397);
xnor U2535 (N_2535,N_2308,N_2337);
nor U2536 (N_2536,N_2316,N_2240);
nand U2537 (N_2537,N_2382,N_2246);
nor U2538 (N_2538,N_2332,N_2300);
nor U2539 (N_2539,N_2305,N_2393);
or U2540 (N_2540,N_2368,N_2346);
and U2541 (N_2541,N_2379,N_2269);
nand U2542 (N_2542,N_2397,N_2299);
nor U2543 (N_2543,N_2318,N_2371);
nor U2544 (N_2544,N_2271,N_2321);
xnor U2545 (N_2545,N_2274,N_2375);
or U2546 (N_2546,N_2315,N_2283);
xor U2547 (N_2547,N_2275,N_2338);
nor U2548 (N_2548,N_2352,N_2315);
or U2549 (N_2549,N_2324,N_2356);
nor U2550 (N_2550,N_2318,N_2356);
xnor U2551 (N_2551,N_2289,N_2323);
nor U2552 (N_2552,N_2247,N_2299);
or U2553 (N_2553,N_2397,N_2249);
or U2554 (N_2554,N_2340,N_2326);
nand U2555 (N_2555,N_2240,N_2341);
and U2556 (N_2556,N_2368,N_2350);
or U2557 (N_2557,N_2309,N_2354);
xnor U2558 (N_2558,N_2262,N_2391);
or U2559 (N_2559,N_2389,N_2379);
and U2560 (N_2560,N_2438,N_2536);
nor U2561 (N_2561,N_2423,N_2485);
and U2562 (N_2562,N_2500,N_2541);
xor U2563 (N_2563,N_2402,N_2429);
nand U2564 (N_2564,N_2419,N_2455);
xor U2565 (N_2565,N_2421,N_2498);
nand U2566 (N_2566,N_2463,N_2453);
nor U2567 (N_2567,N_2442,N_2473);
nor U2568 (N_2568,N_2412,N_2471);
nor U2569 (N_2569,N_2430,N_2443);
or U2570 (N_2570,N_2556,N_2496);
nor U2571 (N_2571,N_2464,N_2492);
or U2572 (N_2572,N_2459,N_2417);
nand U2573 (N_2573,N_2512,N_2504);
nand U2574 (N_2574,N_2418,N_2528);
or U2575 (N_2575,N_2415,N_2416);
xnor U2576 (N_2576,N_2448,N_2405);
nor U2577 (N_2577,N_2523,N_2439);
nand U2578 (N_2578,N_2431,N_2493);
xnor U2579 (N_2579,N_2553,N_2529);
and U2580 (N_2580,N_2467,N_2478);
xor U2581 (N_2581,N_2446,N_2537);
and U2582 (N_2582,N_2451,N_2457);
and U2583 (N_2583,N_2458,N_2411);
nor U2584 (N_2584,N_2520,N_2517);
xor U2585 (N_2585,N_2505,N_2497);
or U2586 (N_2586,N_2456,N_2551);
nand U2587 (N_2587,N_2489,N_2532);
xnor U2588 (N_2588,N_2491,N_2499);
or U2589 (N_2589,N_2518,N_2539);
nand U2590 (N_2590,N_2522,N_2490);
nand U2591 (N_2591,N_2555,N_2527);
and U2592 (N_2592,N_2447,N_2538);
and U2593 (N_2593,N_2428,N_2508);
xor U2594 (N_2594,N_2544,N_2432);
nor U2595 (N_2595,N_2542,N_2433);
nand U2596 (N_2596,N_2481,N_2449);
nor U2597 (N_2597,N_2410,N_2445);
and U2598 (N_2598,N_2404,N_2409);
and U2599 (N_2599,N_2531,N_2510);
and U2600 (N_2600,N_2488,N_2540);
or U2601 (N_2601,N_2552,N_2436);
nand U2602 (N_2602,N_2511,N_2514);
xnor U2603 (N_2603,N_2484,N_2407);
nor U2604 (N_2604,N_2557,N_2452);
or U2605 (N_2605,N_2554,N_2475);
nor U2606 (N_2606,N_2503,N_2547);
xor U2607 (N_2607,N_2486,N_2440);
and U2608 (N_2608,N_2502,N_2549);
nand U2609 (N_2609,N_2509,N_2450);
xor U2610 (N_2610,N_2545,N_2516);
and U2611 (N_2611,N_2495,N_2480);
nand U2612 (N_2612,N_2530,N_2435);
nand U2613 (N_2613,N_2461,N_2482);
or U2614 (N_2614,N_2526,N_2507);
nand U2615 (N_2615,N_2441,N_2466);
nor U2616 (N_2616,N_2513,N_2426);
nor U2617 (N_2617,N_2472,N_2437);
and U2618 (N_2618,N_2521,N_2460);
nand U2619 (N_2619,N_2474,N_2519);
xnor U2620 (N_2620,N_2468,N_2414);
and U2621 (N_2621,N_2479,N_2550);
nor U2622 (N_2622,N_2515,N_2408);
nor U2623 (N_2623,N_2506,N_2501);
xnor U2624 (N_2624,N_2525,N_2543);
and U2625 (N_2625,N_2400,N_2469);
nand U2626 (N_2626,N_2559,N_2425);
or U2627 (N_2627,N_2420,N_2465);
and U2628 (N_2628,N_2444,N_2558);
nor U2629 (N_2629,N_2546,N_2494);
nor U2630 (N_2630,N_2535,N_2470);
or U2631 (N_2631,N_2548,N_2454);
or U2632 (N_2632,N_2476,N_2462);
and U2633 (N_2633,N_2477,N_2524);
nand U2634 (N_2634,N_2403,N_2434);
nor U2635 (N_2635,N_2424,N_2401);
xor U2636 (N_2636,N_2533,N_2422);
and U2637 (N_2637,N_2406,N_2487);
xor U2638 (N_2638,N_2427,N_2534);
or U2639 (N_2639,N_2413,N_2483);
or U2640 (N_2640,N_2558,N_2539);
nand U2641 (N_2641,N_2453,N_2548);
nor U2642 (N_2642,N_2427,N_2407);
and U2643 (N_2643,N_2439,N_2437);
nor U2644 (N_2644,N_2546,N_2545);
nand U2645 (N_2645,N_2452,N_2424);
xor U2646 (N_2646,N_2445,N_2534);
nor U2647 (N_2647,N_2447,N_2427);
and U2648 (N_2648,N_2499,N_2496);
and U2649 (N_2649,N_2489,N_2502);
and U2650 (N_2650,N_2447,N_2534);
or U2651 (N_2651,N_2554,N_2472);
xor U2652 (N_2652,N_2403,N_2486);
or U2653 (N_2653,N_2534,N_2511);
or U2654 (N_2654,N_2486,N_2537);
and U2655 (N_2655,N_2445,N_2502);
nor U2656 (N_2656,N_2519,N_2446);
and U2657 (N_2657,N_2478,N_2401);
xnor U2658 (N_2658,N_2490,N_2414);
xor U2659 (N_2659,N_2402,N_2496);
or U2660 (N_2660,N_2417,N_2452);
xnor U2661 (N_2661,N_2435,N_2532);
nand U2662 (N_2662,N_2475,N_2499);
xor U2663 (N_2663,N_2483,N_2478);
and U2664 (N_2664,N_2414,N_2512);
and U2665 (N_2665,N_2427,N_2406);
nor U2666 (N_2666,N_2463,N_2470);
xnor U2667 (N_2667,N_2544,N_2506);
or U2668 (N_2668,N_2494,N_2502);
xnor U2669 (N_2669,N_2535,N_2424);
and U2670 (N_2670,N_2404,N_2430);
nand U2671 (N_2671,N_2455,N_2412);
and U2672 (N_2672,N_2498,N_2419);
nor U2673 (N_2673,N_2485,N_2407);
and U2674 (N_2674,N_2499,N_2419);
nor U2675 (N_2675,N_2470,N_2476);
or U2676 (N_2676,N_2529,N_2420);
nand U2677 (N_2677,N_2410,N_2411);
xor U2678 (N_2678,N_2494,N_2518);
and U2679 (N_2679,N_2440,N_2531);
xor U2680 (N_2680,N_2505,N_2539);
and U2681 (N_2681,N_2514,N_2487);
xor U2682 (N_2682,N_2523,N_2411);
xor U2683 (N_2683,N_2421,N_2442);
xor U2684 (N_2684,N_2522,N_2455);
and U2685 (N_2685,N_2419,N_2471);
nor U2686 (N_2686,N_2444,N_2441);
or U2687 (N_2687,N_2510,N_2457);
nor U2688 (N_2688,N_2532,N_2546);
and U2689 (N_2689,N_2530,N_2520);
and U2690 (N_2690,N_2410,N_2448);
or U2691 (N_2691,N_2438,N_2558);
nand U2692 (N_2692,N_2491,N_2433);
nor U2693 (N_2693,N_2498,N_2520);
nand U2694 (N_2694,N_2477,N_2522);
nand U2695 (N_2695,N_2535,N_2482);
and U2696 (N_2696,N_2500,N_2411);
nand U2697 (N_2697,N_2481,N_2559);
nor U2698 (N_2698,N_2532,N_2419);
nand U2699 (N_2699,N_2465,N_2523);
xnor U2700 (N_2700,N_2529,N_2532);
nor U2701 (N_2701,N_2514,N_2452);
xnor U2702 (N_2702,N_2550,N_2426);
or U2703 (N_2703,N_2528,N_2529);
xor U2704 (N_2704,N_2431,N_2479);
nand U2705 (N_2705,N_2443,N_2500);
xor U2706 (N_2706,N_2452,N_2475);
or U2707 (N_2707,N_2412,N_2464);
and U2708 (N_2708,N_2469,N_2470);
or U2709 (N_2709,N_2516,N_2455);
nand U2710 (N_2710,N_2540,N_2471);
nor U2711 (N_2711,N_2400,N_2450);
xnor U2712 (N_2712,N_2412,N_2409);
and U2713 (N_2713,N_2448,N_2487);
nand U2714 (N_2714,N_2518,N_2418);
or U2715 (N_2715,N_2550,N_2483);
and U2716 (N_2716,N_2549,N_2420);
nand U2717 (N_2717,N_2499,N_2501);
nor U2718 (N_2718,N_2423,N_2408);
nand U2719 (N_2719,N_2460,N_2436);
nand U2720 (N_2720,N_2690,N_2639);
nor U2721 (N_2721,N_2664,N_2624);
and U2722 (N_2722,N_2687,N_2583);
nor U2723 (N_2723,N_2603,N_2691);
nor U2724 (N_2724,N_2628,N_2668);
and U2725 (N_2725,N_2636,N_2714);
or U2726 (N_2726,N_2606,N_2672);
xnor U2727 (N_2727,N_2702,N_2574);
xnor U2728 (N_2728,N_2635,N_2645);
nor U2729 (N_2729,N_2698,N_2671);
xor U2730 (N_2730,N_2646,N_2713);
and U2731 (N_2731,N_2586,N_2594);
xor U2732 (N_2732,N_2654,N_2611);
or U2733 (N_2733,N_2595,N_2622);
nor U2734 (N_2734,N_2700,N_2695);
nand U2735 (N_2735,N_2616,N_2648);
nand U2736 (N_2736,N_2696,N_2697);
and U2737 (N_2737,N_2598,N_2661);
and U2738 (N_2738,N_2647,N_2681);
xnor U2739 (N_2739,N_2563,N_2568);
nand U2740 (N_2740,N_2629,N_2683);
or U2741 (N_2741,N_2680,N_2564);
xnor U2742 (N_2742,N_2686,N_2585);
or U2743 (N_2743,N_2625,N_2660);
nand U2744 (N_2744,N_2631,N_2581);
xor U2745 (N_2745,N_2708,N_2705);
or U2746 (N_2746,N_2621,N_2615);
xor U2747 (N_2747,N_2623,N_2573);
or U2748 (N_2748,N_2608,N_2718);
nor U2749 (N_2749,N_2685,N_2665);
and U2750 (N_2750,N_2675,N_2716);
or U2751 (N_2751,N_2694,N_2711);
nand U2752 (N_2752,N_2601,N_2580);
nor U2753 (N_2753,N_2650,N_2619);
and U2754 (N_2754,N_2617,N_2659);
nor U2755 (N_2755,N_2592,N_2676);
and U2756 (N_2756,N_2599,N_2704);
nor U2757 (N_2757,N_2658,N_2637);
and U2758 (N_2758,N_2589,N_2667);
and U2759 (N_2759,N_2642,N_2673);
nand U2760 (N_2760,N_2677,N_2689);
and U2761 (N_2761,N_2633,N_2652);
nor U2762 (N_2762,N_2679,N_2715);
xor U2763 (N_2763,N_2587,N_2706);
xor U2764 (N_2764,N_2600,N_2684);
xnor U2765 (N_2765,N_2566,N_2644);
or U2766 (N_2766,N_2693,N_2662);
nor U2767 (N_2767,N_2649,N_2602);
nand U2768 (N_2768,N_2582,N_2666);
nand U2769 (N_2769,N_2707,N_2578);
or U2770 (N_2770,N_2655,N_2567);
and U2771 (N_2771,N_2641,N_2591);
nand U2772 (N_2772,N_2562,N_2620);
nor U2773 (N_2773,N_2709,N_2653);
nor U2774 (N_2774,N_2579,N_2618);
nand U2775 (N_2775,N_2607,N_2670);
xor U2776 (N_2776,N_2597,N_2638);
or U2777 (N_2777,N_2571,N_2710);
nand U2778 (N_2778,N_2630,N_2577);
nand U2779 (N_2779,N_2576,N_2656);
or U2780 (N_2780,N_2590,N_2569);
nand U2781 (N_2781,N_2663,N_2560);
nor U2782 (N_2782,N_2612,N_2678);
and U2783 (N_2783,N_2719,N_2593);
or U2784 (N_2784,N_2613,N_2609);
and U2785 (N_2785,N_2669,N_2640);
nand U2786 (N_2786,N_2614,N_2627);
nor U2787 (N_2787,N_2712,N_2610);
nand U2788 (N_2788,N_2604,N_2605);
nand U2789 (N_2789,N_2682,N_2634);
and U2790 (N_2790,N_2692,N_2572);
nor U2791 (N_2791,N_2717,N_2651);
nor U2792 (N_2792,N_2561,N_2596);
xnor U2793 (N_2793,N_2657,N_2584);
nor U2794 (N_2794,N_2632,N_2674);
or U2795 (N_2795,N_2570,N_2565);
and U2796 (N_2796,N_2688,N_2643);
or U2797 (N_2797,N_2701,N_2588);
nand U2798 (N_2798,N_2626,N_2703);
nand U2799 (N_2799,N_2575,N_2699);
xor U2800 (N_2800,N_2701,N_2634);
nor U2801 (N_2801,N_2712,N_2699);
xor U2802 (N_2802,N_2692,N_2645);
and U2803 (N_2803,N_2616,N_2585);
nor U2804 (N_2804,N_2628,N_2638);
nor U2805 (N_2805,N_2570,N_2663);
nand U2806 (N_2806,N_2706,N_2679);
nand U2807 (N_2807,N_2659,N_2690);
nor U2808 (N_2808,N_2686,N_2566);
and U2809 (N_2809,N_2670,N_2620);
and U2810 (N_2810,N_2710,N_2707);
nor U2811 (N_2811,N_2616,N_2715);
xnor U2812 (N_2812,N_2580,N_2669);
and U2813 (N_2813,N_2656,N_2650);
nor U2814 (N_2814,N_2680,N_2634);
or U2815 (N_2815,N_2688,N_2609);
nand U2816 (N_2816,N_2666,N_2717);
xnor U2817 (N_2817,N_2695,N_2672);
and U2818 (N_2818,N_2641,N_2700);
and U2819 (N_2819,N_2619,N_2614);
nor U2820 (N_2820,N_2665,N_2577);
and U2821 (N_2821,N_2707,N_2657);
nor U2822 (N_2822,N_2636,N_2637);
nand U2823 (N_2823,N_2703,N_2584);
and U2824 (N_2824,N_2610,N_2592);
or U2825 (N_2825,N_2642,N_2611);
or U2826 (N_2826,N_2664,N_2666);
or U2827 (N_2827,N_2697,N_2632);
and U2828 (N_2828,N_2718,N_2610);
nor U2829 (N_2829,N_2652,N_2703);
xor U2830 (N_2830,N_2595,N_2566);
or U2831 (N_2831,N_2567,N_2665);
nor U2832 (N_2832,N_2591,N_2706);
xor U2833 (N_2833,N_2673,N_2664);
xor U2834 (N_2834,N_2561,N_2597);
nor U2835 (N_2835,N_2560,N_2708);
nand U2836 (N_2836,N_2566,N_2710);
and U2837 (N_2837,N_2624,N_2585);
and U2838 (N_2838,N_2573,N_2601);
nand U2839 (N_2839,N_2709,N_2702);
nor U2840 (N_2840,N_2566,N_2705);
nand U2841 (N_2841,N_2719,N_2582);
or U2842 (N_2842,N_2632,N_2637);
and U2843 (N_2843,N_2679,N_2650);
xor U2844 (N_2844,N_2659,N_2635);
xnor U2845 (N_2845,N_2584,N_2709);
and U2846 (N_2846,N_2589,N_2604);
nand U2847 (N_2847,N_2645,N_2669);
xor U2848 (N_2848,N_2629,N_2684);
xnor U2849 (N_2849,N_2560,N_2684);
and U2850 (N_2850,N_2616,N_2668);
xnor U2851 (N_2851,N_2583,N_2689);
or U2852 (N_2852,N_2682,N_2649);
or U2853 (N_2853,N_2583,N_2614);
nand U2854 (N_2854,N_2675,N_2646);
nand U2855 (N_2855,N_2635,N_2610);
nor U2856 (N_2856,N_2705,N_2637);
nor U2857 (N_2857,N_2560,N_2710);
or U2858 (N_2858,N_2668,N_2618);
xor U2859 (N_2859,N_2572,N_2698);
xor U2860 (N_2860,N_2690,N_2642);
or U2861 (N_2861,N_2578,N_2574);
or U2862 (N_2862,N_2576,N_2661);
nand U2863 (N_2863,N_2637,N_2599);
nand U2864 (N_2864,N_2632,N_2593);
xor U2865 (N_2865,N_2603,N_2702);
or U2866 (N_2866,N_2595,N_2562);
xnor U2867 (N_2867,N_2560,N_2579);
nor U2868 (N_2868,N_2664,N_2621);
nand U2869 (N_2869,N_2569,N_2704);
nand U2870 (N_2870,N_2648,N_2626);
nor U2871 (N_2871,N_2562,N_2636);
nand U2872 (N_2872,N_2710,N_2583);
nor U2873 (N_2873,N_2674,N_2693);
and U2874 (N_2874,N_2671,N_2706);
nor U2875 (N_2875,N_2605,N_2671);
xnor U2876 (N_2876,N_2599,N_2711);
xnor U2877 (N_2877,N_2717,N_2679);
nor U2878 (N_2878,N_2655,N_2640);
or U2879 (N_2879,N_2608,N_2571);
nand U2880 (N_2880,N_2729,N_2838);
and U2881 (N_2881,N_2865,N_2753);
xnor U2882 (N_2882,N_2778,N_2863);
nor U2883 (N_2883,N_2874,N_2794);
nand U2884 (N_2884,N_2805,N_2786);
and U2885 (N_2885,N_2746,N_2806);
nand U2886 (N_2886,N_2798,N_2809);
and U2887 (N_2887,N_2781,N_2857);
nand U2888 (N_2888,N_2800,N_2818);
xnor U2889 (N_2889,N_2722,N_2854);
nand U2890 (N_2890,N_2769,N_2772);
nand U2891 (N_2891,N_2733,N_2754);
xor U2892 (N_2892,N_2732,N_2723);
and U2893 (N_2893,N_2742,N_2825);
nand U2894 (N_2894,N_2749,N_2728);
nand U2895 (N_2895,N_2835,N_2765);
xor U2896 (N_2896,N_2726,N_2796);
nand U2897 (N_2897,N_2855,N_2851);
or U2898 (N_2898,N_2738,N_2756);
xor U2899 (N_2899,N_2758,N_2802);
or U2900 (N_2900,N_2844,N_2793);
or U2901 (N_2901,N_2832,N_2807);
xor U2902 (N_2902,N_2830,N_2878);
or U2903 (N_2903,N_2811,N_2762);
nor U2904 (N_2904,N_2819,N_2833);
and U2905 (N_2905,N_2760,N_2877);
nor U2906 (N_2906,N_2871,N_2849);
nor U2907 (N_2907,N_2759,N_2731);
or U2908 (N_2908,N_2730,N_2822);
and U2909 (N_2909,N_2839,N_2724);
nand U2910 (N_2910,N_2803,N_2780);
nand U2911 (N_2911,N_2790,N_2840);
nor U2912 (N_2912,N_2873,N_2864);
and U2913 (N_2913,N_2870,N_2770);
nor U2914 (N_2914,N_2824,N_2745);
or U2915 (N_2915,N_2816,N_2842);
or U2916 (N_2916,N_2775,N_2741);
nand U2917 (N_2917,N_2856,N_2783);
xnor U2918 (N_2918,N_2740,N_2829);
nand U2919 (N_2919,N_2737,N_2821);
nand U2920 (N_2920,N_2792,N_2795);
and U2921 (N_2921,N_2766,N_2773);
and U2922 (N_2922,N_2777,N_2748);
nand U2923 (N_2923,N_2812,N_2744);
nor U2924 (N_2924,N_2868,N_2779);
nand U2925 (N_2925,N_2734,N_2866);
nor U2926 (N_2926,N_2834,N_2791);
nand U2927 (N_2927,N_2785,N_2841);
nor U2928 (N_2928,N_2743,N_2727);
xor U2929 (N_2929,N_2847,N_2751);
nor U2930 (N_2930,N_2858,N_2815);
nand U2931 (N_2931,N_2784,N_2767);
or U2932 (N_2932,N_2755,N_2859);
nand U2933 (N_2933,N_2757,N_2860);
or U2934 (N_2934,N_2735,N_2843);
xnor U2935 (N_2935,N_2797,N_2845);
nor U2936 (N_2936,N_2750,N_2768);
and U2937 (N_2937,N_2817,N_2804);
or U2938 (N_2938,N_2771,N_2831);
nand U2939 (N_2939,N_2808,N_2846);
nor U2940 (N_2940,N_2764,N_2761);
nor U2941 (N_2941,N_2747,N_2736);
and U2942 (N_2942,N_2752,N_2869);
nand U2943 (N_2943,N_2872,N_2782);
xnor U2944 (N_2944,N_2850,N_2827);
nand U2945 (N_2945,N_2879,N_2725);
and U2946 (N_2946,N_2799,N_2861);
nor U2947 (N_2947,N_2801,N_2789);
or U2948 (N_2948,N_2828,N_2876);
and U2949 (N_2949,N_2836,N_2810);
or U2950 (N_2950,N_2814,N_2867);
nor U2951 (N_2951,N_2763,N_2848);
xnor U2952 (N_2952,N_2823,N_2820);
and U2953 (N_2953,N_2862,N_2721);
nand U2954 (N_2954,N_2739,N_2852);
nor U2955 (N_2955,N_2720,N_2776);
xor U2956 (N_2956,N_2774,N_2813);
xnor U2957 (N_2957,N_2787,N_2875);
and U2958 (N_2958,N_2837,N_2826);
nand U2959 (N_2959,N_2853,N_2788);
xor U2960 (N_2960,N_2723,N_2792);
and U2961 (N_2961,N_2783,N_2838);
xor U2962 (N_2962,N_2831,N_2811);
and U2963 (N_2963,N_2736,N_2855);
nor U2964 (N_2964,N_2822,N_2792);
nand U2965 (N_2965,N_2825,N_2827);
xnor U2966 (N_2966,N_2768,N_2795);
xor U2967 (N_2967,N_2767,N_2838);
nor U2968 (N_2968,N_2799,N_2835);
nand U2969 (N_2969,N_2784,N_2785);
nand U2970 (N_2970,N_2752,N_2837);
xnor U2971 (N_2971,N_2791,N_2878);
or U2972 (N_2972,N_2854,N_2742);
nand U2973 (N_2973,N_2856,N_2734);
xor U2974 (N_2974,N_2759,N_2839);
xor U2975 (N_2975,N_2760,N_2866);
or U2976 (N_2976,N_2871,N_2723);
or U2977 (N_2977,N_2729,N_2841);
xor U2978 (N_2978,N_2777,N_2819);
or U2979 (N_2979,N_2738,N_2787);
nor U2980 (N_2980,N_2863,N_2793);
or U2981 (N_2981,N_2799,N_2779);
xnor U2982 (N_2982,N_2823,N_2832);
and U2983 (N_2983,N_2817,N_2778);
or U2984 (N_2984,N_2807,N_2870);
nor U2985 (N_2985,N_2851,N_2825);
or U2986 (N_2986,N_2800,N_2798);
nor U2987 (N_2987,N_2823,N_2740);
nand U2988 (N_2988,N_2828,N_2787);
and U2989 (N_2989,N_2852,N_2839);
nand U2990 (N_2990,N_2858,N_2826);
xor U2991 (N_2991,N_2799,N_2762);
nand U2992 (N_2992,N_2787,N_2752);
nand U2993 (N_2993,N_2844,N_2873);
or U2994 (N_2994,N_2839,N_2780);
xnor U2995 (N_2995,N_2821,N_2870);
and U2996 (N_2996,N_2802,N_2842);
and U2997 (N_2997,N_2722,N_2825);
or U2998 (N_2998,N_2813,N_2846);
nor U2999 (N_2999,N_2818,N_2850);
or U3000 (N_3000,N_2835,N_2755);
and U3001 (N_3001,N_2731,N_2857);
and U3002 (N_3002,N_2865,N_2860);
or U3003 (N_3003,N_2831,N_2743);
or U3004 (N_3004,N_2819,N_2774);
nand U3005 (N_3005,N_2736,N_2725);
and U3006 (N_3006,N_2851,N_2804);
nor U3007 (N_3007,N_2873,N_2785);
and U3008 (N_3008,N_2791,N_2824);
nor U3009 (N_3009,N_2830,N_2781);
xor U3010 (N_3010,N_2791,N_2759);
and U3011 (N_3011,N_2834,N_2784);
nor U3012 (N_3012,N_2803,N_2732);
and U3013 (N_3013,N_2853,N_2776);
xnor U3014 (N_3014,N_2856,N_2747);
or U3015 (N_3015,N_2849,N_2801);
or U3016 (N_3016,N_2761,N_2861);
nor U3017 (N_3017,N_2878,N_2869);
nand U3018 (N_3018,N_2750,N_2873);
and U3019 (N_3019,N_2790,N_2854);
or U3020 (N_3020,N_2777,N_2806);
or U3021 (N_3021,N_2804,N_2809);
and U3022 (N_3022,N_2802,N_2845);
and U3023 (N_3023,N_2827,N_2761);
or U3024 (N_3024,N_2770,N_2867);
xnor U3025 (N_3025,N_2802,N_2860);
nand U3026 (N_3026,N_2877,N_2873);
or U3027 (N_3027,N_2787,N_2869);
or U3028 (N_3028,N_2770,N_2756);
nor U3029 (N_3029,N_2797,N_2764);
and U3030 (N_3030,N_2724,N_2844);
nor U3031 (N_3031,N_2749,N_2725);
and U3032 (N_3032,N_2830,N_2859);
or U3033 (N_3033,N_2872,N_2820);
xnor U3034 (N_3034,N_2850,N_2840);
nand U3035 (N_3035,N_2834,N_2837);
nor U3036 (N_3036,N_2773,N_2794);
nand U3037 (N_3037,N_2800,N_2833);
xor U3038 (N_3038,N_2854,N_2876);
nor U3039 (N_3039,N_2726,N_2877);
and U3040 (N_3040,N_3005,N_3007);
nand U3041 (N_3041,N_3010,N_3018);
nor U3042 (N_3042,N_2898,N_3026);
and U3043 (N_3043,N_3012,N_2989);
and U3044 (N_3044,N_3031,N_2950);
xor U3045 (N_3045,N_2887,N_3034);
nor U3046 (N_3046,N_3023,N_2971);
or U3047 (N_3047,N_2993,N_3038);
nand U3048 (N_3048,N_3035,N_2978);
nor U3049 (N_3049,N_3002,N_2920);
or U3050 (N_3050,N_2910,N_2969);
xnor U3051 (N_3051,N_2968,N_2939);
nand U3052 (N_3052,N_2908,N_2930);
xor U3053 (N_3053,N_2980,N_2995);
nor U3054 (N_3054,N_3013,N_2921);
nand U3055 (N_3055,N_2927,N_2943);
nand U3056 (N_3056,N_2900,N_2933);
nand U3057 (N_3057,N_2972,N_3004);
xnor U3058 (N_3058,N_2983,N_3016);
nor U3059 (N_3059,N_2883,N_3039);
or U3060 (N_3060,N_2997,N_2938);
nand U3061 (N_3061,N_2990,N_2952);
nand U3062 (N_3062,N_3009,N_2970);
xor U3063 (N_3063,N_2914,N_3022);
or U3064 (N_3064,N_2988,N_3032);
nor U3065 (N_3065,N_2967,N_3015);
and U3066 (N_3066,N_2891,N_2979);
and U3067 (N_3067,N_2922,N_2884);
nand U3068 (N_3068,N_2940,N_2962);
and U3069 (N_3069,N_2996,N_2893);
xnor U3070 (N_3070,N_2954,N_2941);
or U3071 (N_3071,N_3008,N_2959);
nor U3072 (N_3072,N_2942,N_3000);
xnor U3073 (N_3073,N_2951,N_3028);
nor U3074 (N_3074,N_2966,N_2987);
nand U3075 (N_3075,N_2947,N_2899);
and U3076 (N_3076,N_2961,N_2912);
or U3077 (N_3077,N_2964,N_2886);
and U3078 (N_3078,N_3014,N_2881);
nand U3079 (N_3079,N_2904,N_2896);
xor U3080 (N_3080,N_2902,N_2982);
xnor U3081 (N_3081,N_2919,N_2974);
or U3082 (N_3082,N_3027,N_2999);
xnor U3083 (N_3083,N_2998,N_2931);
nand U3084 (N_3084,N_2885,N_2901);
nor U3085 (N_3085,N_3017,N_2888);
or U3086 (N_3086,N_2975,N_2992);
nand U3087 (N_3087,N_2948,N_2965);
or U3088 (N_3088,N_2981,N_2955);
nor U3089 (N_3089,N_2918,N_2949);
nand U3090 (N_3090,N_3019,N_2906);
or U3091 (N_3091,N_2895,N_2945);
xor U3092 (N_3092,N_3036,N_2958);
nand U3093 (N_3093,N_2911,N_2960);
nand U3094 (N_3094,N_2944,N_2929);
or U3095 (N_3095,N_2925,N_2932);
and U3096 (N_3096,N_2909,N_3003);
or U3097 (N_3097,N_2907,N_3033);
nand U3098 (N_3098,N_2984,N_3001);
nand U3099 (N_3099,N_2915,N_2926);
and U3100 (N_3100,N_2917,N_2905);
nand U3101 (N_3101,N_2937,N_2935);
nor U3102 (N_3102,N_2957,N_3020);
nor U3103 (N_3103,N_3030,N_2936);
nand U3104 (N_3104,N_2986,N_2897);
nor U3105 (N_3105,N_2892,N_2963);
or U3106 (N_3106,N_2991,N_2882);
or U3107 (N_3107,N_2890,N_2894);
and U3108 (N_3108,N_2924,N_3006);
xnor U3109 (N_3109,N_3025,N_2985);
nand U3110 (N_3110,N_2956,N_3011);
xnor U3111 (N_3111,N_2903,N_2934);
and U3112 (N_3112,N_3024,N_2928);
xnor U3113 (N_3113,N_3037,N_2946);
nor U3114 (N_3114,N_2916,N_3021);
xnor U3115 (N_3115,N_2889,N_2913);
nand U3116 (N_3116,N_2880,N_3029);
nand U3117 (N_3117,N_2976,N_2994);
or U3118 (N_3118,N_2923,N_2973);
nand U3119 (N_3119,N_2977,N_2953);
and U3120 (N_3120,N_2955,N_2982);
and U3121 (N_3121,N_2981,N_3011);
nor U3122 (N_3122,N_2941,N_2903);
xnor U3123 (N_3123,N_2989,N_2909);
and U3124 (N_3124,N_3032,N_2903);
or U3125 (N_3125,N_3014,N_2979);
nand U3126 (N_3126,N_3022,N_2940);
xnor U3127 (N_3127,N_2920,N_2978);
nand U3128 (N_3128,N_3000,N_2982);
xnor U3129 (N_3129,N_3035,N_2909);
nand U3130 (N_3130,N_2934,N_3029);
and U3131 (N_3131,N_2967,N_2917);
nor U3132 (N_3132,N_2959,N_2951);
nand U3133 (N_3133,N_2920,N_2884);
nand U3134 (N_3134,N_2898,N_2973);
or U3135 (N_3135,N_3015,N_3038);
nor U3136 (N_3136,N_2998,N_3030);
nor U3137 (N_3137,N_2933,N_2960);
nand U3138 (N_3138,N_2903,N_2963);
or U3139 (N_3139,N_2937,N_2909);
nand U3140 (N_3140,N_3018,N_2993);
and U3141 (N_3141,N_2902,N_2983);
nor U3142 (N_3142,N_3012,N_2956);
nand U3143 (N_3143,N_2896,N_3000);
nor U3144 (N_3144,N_2959,N_2881);
nand U3145 (N_3145,N_2890,N_2935);
nor U3146 (N_3146,N_2903,N_2952);
or U3147 (N_3147,N_2958,N_2945);
xor U3148 (N_3148,N_2893,N_2899);
nor U3149 (N_3149,N_2933,N_2966);
and U3150 (N_3150,N_3035,N_2960);
or U3151 (N_3151,N_2940,N_2991);
xor U3152 (N_3152,N_2919,N_2908);
xnor U3153 (N_3153,N_3014,N_3039);
and U3154 (N_3154,N_3036,N_3037);
and U3155 (N_3155,N_2971,N_2918);
and U3156 (N_3156,N_2888,N_2882);
or U3157 (N_3157,N_2902,N_2891);
and U3158 (N_3158,N_2998,N_3032);
and U3159 (N_3159,N_2982,N_2891);
nand U3160 (N_3160,N_3032,N_3035);
or U3161 (N_3161,N_2999,N_2904);
and U3162 (N_3162,N_2960,N_2956);
nand U3163 (N_3163,N_3004,N_2961);
or U3164 (N_3164,N_2905,N_2961);
nor U3165 (N_3165,N_2998,N_3001);
nand U3166 (N_3166,N_2888,N_2963);
xor U3167 (N_3167,N_3003,N_2963);
or U3168 (N_3168,N_2933,N_2926);
nor U3169 (N_3169,N_2900,N_2956);
nor U3170 (N_3170,N_2949,N_2951);
nor U3171 (N_3171,N_3022,N_2970);
xor U3172 (N_3172,N_2923,N_2963);
nand U3173 (N_3173,N_2918,N_3000);
nor U3174 (N_3174,N_2969,N_2965);
or U3175 (N_3175,N_2906,N_3015);
xnor U3176 (N_3176,N_2881,N_3037);
and U3177 (N_3177,N_2985,N_2931);
nor U3178 (N_3178,N_2933,N_3023);
or U3179 (N_3179,N_3028,N_3019);
xor U3180 (N_3180,N_2929,N_2887);
and U3181 (N_3181,N_2989,N_2992);
nor U3182 (N_3182,N_2932,N_2950);
xor U3183 (N_3183,N_2948,N_2959);
and U3184 (N_3184,N_2998,N_3021);
nand U3185 (N_3185,N_2913,N_2912);
or U3186 (N_3186,N_2990,N_2930);
nor U3187 (N_3187,N_3036,N_2900);
nor U3188 (N_3188,N_3017,N_2983);
and U3189 (N_3189,N_3030,N_2990);
and U3190 (N_3190,N_3029,N_3015);
and U3191 (N_3191,N_2940,N_3038);
and U3192 (N_3192,N_2967,N_3019);
and U3193 (N_3193,N_2880,N_2978);
nor U3194 (N_3194,N_2926,N_2904);
or U3195 (N_3195,N_3034,N_2980);
xor U3196 (N_3196,N_2916,N_2922);
nor U3197 (N_3197,N_2893,N_2977);
nor U3198 (N_3198,N_2996,N_2880);
nor U3199 (N_3199,N_2954,N_2968);
and U3200 (N_3200,N_3065,N_3161);
nor U3201 (N_3201,N_3088,N_3085);
xor U3202 (N_3202,N_3184,N_3192);
xor U3203 (N_3203,N_3074,N_3067);
nor U3204 (N_3204,N_3137,N_3114);
xor U3205 (N_3205,N_3092,N_3090);
nor U3206 (N_3206,N_3094,N_3128);
xnor U3207 (N_3207,N_3191,N_3133);
xnor U3208 (N_3208,N_3140,N_3185);
and U3209 (N_3209,N_3150,N_3080);
nand U3210 (N_3210,N_3145,N_3183);
or U3211 (N_3211,N_3050,N_3170);
nand U3212 (N_3212,N_3047,N_3081);
nand U3213 (N_3213,N_3167,N_3131);
xnor U3214 (N_3214,N_3123,N_3174);
nor U3215 (N_3215,N_3196,N_3112);
xnor U3216 (N_3216,N_3143,N_3043);
nand U3217 (N_3217,N_3181,N_3164);
and U3218 (N_3218,N_3073,N_3125);
xnor U3219 (N_3219,N_3130,N_3177);
xor U3220 (N_3220,N_3101,N_3151);
nor U3221 (N_3221,N_3093,N_3069);
xnor U3222 (N_3222,N_3190,N_3180);
nor U3223 (N_3223,N_3162,N_3046);
xor U3224 (N_3224,N_3102,N_3138);
or U3225 (N_3225,N_3165,N_3105);
nor U3226 (N_3226,N_3115,N_3134);
and U3227 (N_3227,N_3056,N_3097);
nor U3228 (N_3228,N_3111,N_3060);
xnor U3229 (N_3229,N_3045,N_3144);
or U3230 (N_3230,N_3155,N_3197);
xor U3231 (N_3231,N_3091,N_3062);
or U3232 (N_3232,N_3078,N_3157);
or U3233 (N_3233,N_3107,N_3068);
nor U3234 (N_3234,N_3109,N_3173);
nor U3235 (N_3235,N_3049,N_3083);
and U3236 (N_3236,N_3187,N_3059);
or U3237 (N_3237,N_3175,N_3052);
nor U3238 (N_3238,N_3061,N_3042);
or U3239 (N_3239,N_3055,N_3087);
and U3240 (N_3240,N_3072,N_3179);
nor U3241 (N_3241,N_3189,N_3160);
and U3242 (N_3242,N_3178,N_3053);
or U3243 (N_3243,N_3064,N_3166);
xnor U3244 (N_3244,N_3158,N_3117);
nor U3245 (N_3245,N_3195,N_3149);
nor U3246 (N_3246,N_3077,N_3147);
xor U3247 (N_3247,N_3119,N_3186);
nand U3248 (N_3248,N_3126,N_3148);
nand U3249 (N_3249,N_3096,N_3057);
and U3250 (N_3250,N_3118,N_3063);
and U3251 (N_3251,N_3124,N_3122);
nor U3252 (N_3252,N_3108,N_3113);
nand U3253 (N_3253,N_3110,N_3048);
and U3254 (N_3254,N_3044,N_3142);
nand U3255 (N_3255,N_3116,N_3141);
nand U3256 (N_3256,N_3176,N_3082);
or U3257 (N_3257,N_3104,N_3199);
xor U3258 (N_3258,N_3152,N_3194);
or U3259 (N_3259,N_3168,N_3066);
nand U3260 (N_3260,N_3079,N_3106);
nor U3261 (N_3261,N_3156,N_3159);
or U3262 (N_3262,N_3076,N_3139);
nand U3263 (N_3263,N_3198,N_3075);
and U3264 (N_3264,N_3172,N_3163);
nand U3265 (N_3265,N_3099,N_3070);
and U3266 (N_3266,N_3086,N_3041);
xor U3267 (N_3267,N_3040,N_3095);
xor U3268 (N_3268,N_3193,N_3100);
nor U3269 (N_3269,N_3051,N_3054);
nand U3270 (N_3270,N_3103,N_3089);
nor U3271 (N_3271,N_3154,N_3098);
and U3272 (N_3272,N_3135,N_3146);
or U3273 (N_3273,N_3136,N_3084);
nand U3274 (N_3274,N_3169,N_3129);
nand U3275 (N_3275,N_3188,N_3153);
or U3276 (N_3276,N_3171,N_3132);
nand U3277 (N_3277,N_3127,N_3120);
nor U3278 (N_3278,N_3071,N_3058);
and U3279 (N_3279,N_3182,N_3121);
xor U3280 (N_3280,N_3152,N_3140);
xnor U3281 (N_3281,N_3075,N_3049);
and U3282 (N_3282,N_3093,N_3040);
or U3283 (N_3283,N_3061,N_3118);
or U3284 (N_3284,N_3141,N_3164);
nor U3285 (N_3285,N_3113,N_3076);
xor U3286 (N_3286,N_3199,N_3191);
and U3287 (N_3287,N_3041,N_3062);
and U3288 (N_3288,N_3109,N_3097);
nand U3289 (N_3289,N_3181,N_3091);
or U3290 (N_3290,N_3154,N_3106);
xnor U3291 (N_3291,N_3169,N_3157);
and U3292 (N_3292,N_3066,N_3178);
or U3293 (N_3293,N_3118,N_3106);
nand U3294 (N_3294,N_3153,N_3099);
nor U3295 (N_3295,N_3055,N_3141);
nand U3296 (N_3296,N_3154,N_3090);
xor U3297 (N_3297,N_3116,N_3191);
and U3298 (N_3298,N_3196,N_3043);
nand U3299 (N_3299,N_3193,N_3055);
nor U3300 (N_3300,N_3153,N_3182);
or U3301 (N_3301,N_3069,N_3087);
nand U3302 (N_3302,N_3119,N_3097);
or U3303 (N_3303,N_3136,N_3197);
nand U3304 (N_3304,N_3125,N_3081);
nor U3305 (N_3305,N_3197,N_3066);
nand U3306 (N_3306,N_3134,N_3073);
or U3307 (N_3307,N_3075,N_3097);
nor U3308 (N_3308,N_3068,N_3170);
or U3309 (N_3309,N_3107,N_3083);
xor U3310 (N_3310,N_3165,N_3052);
or U3311 (N_3311,N_3117,N_3144);
xor U3312 (N_3312,N_3171,N_3099);
nor U3313 (N_3313,N_3135,N_3147);
and U3314 (N_3314,N_3197,N_3065);
xnor U3315 (N_3315,N_3054,N_3191);
nor U3316 (N_3316,N_3071,N_3148);
or U3317 (N_3317,N_3169,N_3133);
nor U3318 (N_3318,N_3114,N_3130);
nor U3319 (N_3319,N_3065,N_3068);
xnor U3320 (N_3320,N_3073,N_3149);
or U3321 (N_3321,N_3094,N_3132);
xor U3322 (N_3322,N_3116,N_3151);
and U3323 (N_3323,N_3042,N_3082);
and U3324 (N_3324,N_3059,N_3139);
xor U3325 (N_3325,N_3073,N_3174);
nor U3326 (N_3326,N_3113,N_3177);
nor U3327 (N_3327,N_3157,N_3159);
and U3328 (N_3328,N_3105,N_3138);
or U3329 (N_3329,N_3170,N_3114);
nor U3330 (N_3330,N_3145,N_3103);
nor U3331 (N_3331,N_3177,N_3159);
or U3332 (N_3332,N_3080,N_3160);
and U3333 (N_3333,N_3159,N_3189);
xnor U3334 (N_3334,N_3111,N_3179);
and U3335 (N_3335,N_3182,N_3165);
or U3336 (N_3336,N_3176,N_3076);
xor U3337 (N_3337,N_3069,N_3193);
nor U3338 (N_3338,N_3112,N_3111);
nor U3339 (N_3339,N_3148,N_3125);
nand U3340 (N_3340,N_3058,N_3068);
or U3341 (N_3341,N_3091,N_3161);
xnor U3342 (N_3342,N_3065,N_3199);
nor U3343 (N_3343,N_3069,N_3141);
or U3344 (N_3344,N_3183,N_3146);
nand U3345 (N_3345,N_3170,N_3090);
xnor U3346 (N_3346,N_3072,N_3163);
nor U3347 (N_3347,N_3084,N_3196);
or U3348 (N_3348,N_3093,N_3193);
xnor U3349 (N_3349,N_3155,N_3054);
xor U3350 (N_3350,N_3048,N_3096);
nand U3351 (N_3351,N_3161,N_3041);
or U3352 (N_3352,N_3103,N_3095);
nand U3353 (N_3353,N_3119,N_3100);
or U3354 (N_3354,N_3064,N_3115);
nor U3355 (N_3355,N_3157,N_3067);
nand U3356 (N_3356,N_3196,N_3163);
nand U3357 (N_3357,N_3089,N_3160);
nor U3358 (N_3358,N_3096,N_3155);
xnor U3359 (N_3359,N_3057,N_3069);
and U3360 (N_3360,N_3327,N_3359);
xor U3361 (N_3361,N_3277,N_3313);
or U3362 (N_3362,N_3235,N_3206);
xor U3363 (N_3363,N_3226,N_3205);
or U3364 (N_3364,N_3292,N_3320);
and U3365 (N_3365,N_3258,N_3330);
xor U3366 (N_3366,N_3295,N_3311);
or U3367 (N_3367,N_3215,N_3324);
nor U3368 (N_3368,N_3305,N_3221);
nor U3369 (N_3369,N_3231,N_3214);
or U3370 (N_3370,N_3236,N_3293);
or U3371 (N_3371,N_3256,N_3230);
or U3372 (N_3372,N_3309,N_3300);
and U3373 (N_3373,N_3248,N_3259);
or U3374 (N_3374,N_3314,N_3303);
xnor U3375 (N_3375,N_3268,N_3265);
nand U3376 (N_3376,N_3271,N_3253);
xnor U3377 (N_3377,N_3290,N_3229);
or U3378 (N_3378,N_3270,N_3306);
nor U3379 (N_3379,N_3353,N_3242);
and U3380 (N_3380,N_3334,N_3202);
and U3381 (N_3381,N_3257,N_3250);
and U3382 (N_3382,N_3280,N_3341);
and U3383 (N_3383,N_3326,N_3282);
nand U3384 (N_3384,N_3241,N_3217);
or U3385 (N_3385,N_3267,N_3332);
nor U3386 (N_3386,N_3211,N_3266);
xnor U3387 (N_3387,N_3349,N_3247);
nand U3388 (N_3388,N_3336,N_3299);
or U3389 (N_3389,N_3200,N_3335);
nor U3390 (N_3390,N_3203,N_3263);
and U3391 (N_3391,N_3346,N_3232);
or U3392 (N_3392,N_3342,N_3201);
xnor U3393 (N_3393,N_3219,N_3323);
or U3394 (N_3394,N_3224,N_3212);
and U3395 (N_3395,N_3283,N_3262);
xnor U3396 (N_3396,N_3284,N_3358);
and U3397 (N_3397,N_3260,N_3261);
xnor U3398 (N_3398,N_3273,N_3351);
nor U3399 (N_3399,N_3272,N_3298);
or U3400 (N_3400,N_3209,N_3246);
or U3401 (N_3401,N_3315,N_3302);
xor U3402 (N_3402,N_3285,N_3222);
and U3403 (N_3403,N_3274,N_3269);
and U3404 (N_3404,N_3239,N_3333);
nand U3405 (N_3405,N_3223,N_3347);
and U3406 (N_3406,N_3331,N_3301);
nand U3407 (N_3407,N_3343,N_3356);
xnor U3408 (N_3408,N_3238,N_3264);
or U3409 (N_3409,N_3275,N_3319);
nor U3410 (N_3410,N_3318,N_3249);
xnor U3411 (N_3411,N_3339,N_3278);
xnor U3412 (N_3412,N_3310,N_3307);
nand U3413 (N_3413,N_3294,N_3204);
nand U3414 (N_3414,N_3251,N_3207);
xor U3415 (N_3415,N_3254,N_3322);
xor U3416 (N_3416,N_3338,N_3329);
xnor U3417 (N_3417,N_3321,N_3244);
xnor U3418 (N_3418,N_3245,N_3243);
nand U3419 (N_3419,N_3218,N_3297);
or U3420 (N_3420,N_3225,N_3317);
nor U3421 (N_3421,N_3354,N_3316);
nor U3422 (N_3422,N_3355,N_3348);
or U3423 (N_3423,N_3252,N_3237);
nand U3424 (N_3424,N_3240,N_3234);
and U3425 (N_3425,N_3304,N_3357);
xnor U3426 (N_3426,N_3287,N_3281);
and U3427 (N_3427,N_3345,N_3228);
nor U3428 (N_3428,N_3325,N_3337);
nand U3429 (N_3429,N_3233,N_3276);
or U3430 (N_3430,N_3340,N_3255);
or U3431 (N_3431,N_3220,N_3312);
and U3432 (N_3432,N_3328,N_3350);
or U3433 (N_3433,N_3291,N_3352);
nand U3434 (N_3434,N_3208,N_3213);
or U3435 (N_3435,N_3308,N_3210);
and U3436 (N_3436,N_3288,N_3289);
or U3437 (N_3437,N_3344,N_3286);
or U3438 (N_3438,N_3227,N_3216);
xnor U3439 (N_3439,N_3279,N_3296);
or U3440 (N_3440,N_3279,N_3313);
nor U3441 (N_3441,N_3326,N_3313);
and U3442 (N_3442,N_3341,N_3283);
nand U3443 (N_3443,N_3277,N_3206);
nand U3444 (N_3444,N_3296,N_3290);
xor U3445 (N_3445,N_3217,N_3331);
nand U3446 (N_3446,N_3266,N_3220);
nor U3447 (N_3447,N_3299,N_3221);
or U3448 (N_3448,N_3299,N_3357);
and U3449 (N_3449,N_3277,N_3246);
xor U3450 (N_3450,N_3304,N_3228);
nor U3451 (N_3451,N_3339,N_3272);
nand U3452 (N_3452,N_3205,N_3231);
or U3453 (N_3453,N_3301,N_3351);
and U3454 (N_3454,N_3318,N_3303);
or U3455 (N_3455,N_3329,N_3285);
or U3456 (N_3456,N_3288,N_3259);
nor U3457 (N_3457,N_3265,N_3302);
xor U3458 (N_3458,N_3323,N_3251);
nor U3459 (N_3459,N_3335,N_3296);
xnor U3460 (N_3460,N_3213,N_3324);
nand U3461 (N_3461,N_3216,N_3283);
nor U3462 (N_3462,N_3250,N_3349);
nor U3463 (N_3463,N_3282,N_3308);
or U3464 (N_3464,N_3311,N_3209);
or U3465 (N_3465,N_3304,N_3303);
or U3466 (N_3466,N_3268,N_3303);
nand U3467 (N_3467,N_3222,N_3289);
or U3468 (N_3468,N_3311,N_3283);
and U3469 (N_3469,N_3213,N_3283);
and U3470 (N_3470,N_3305,N_3296);
nor U3471 (N_3471,N_3321,N_3319);
or U3472 (N_3472,N_3256,N_3266);
nand U3473 (N_3473,N_3257,N_3290);
nor U3474 (N_3474,N_3291,N_3306);
or U3475 (N_3475,N_3329,N_3282);
or U3476 (N_3476,N_3346,N_3328);
nor U3477 (N_3477,N_3222,N_3256);
and U3478 (N_3478,N_3289,N_3266);
and U3479 (N_3479,N_3297,N_3285);
or U3480 (N_3480,N_3314,N_3232);
nand U3481 (N_3481,N_3344,N_3256);
and U3482 (N_3482,N_3205,N_3214);
or U3483 (N_3483,N_3300,N_3312);
or U3484 (N_3484,N_3307,N_3241);
nand U3485 (N_3485,N_3335,N_3310);
xor U3486 (N_3486,N_3319,N_3274);
nand U3487 (N_3487,N_3318,N_3258);
or U3488 (N_3488,N_3302,N_3285);
xor U3489 (N_3489,N_3260,N_3269);
nor U3490 (N_3490,N_3355,N_3312);
and U3491 (N_3491,N_3272,N_3283);
and U3492 (N_3492,N_3236,N_3313);
nor U3493 (N_3493,N_3209,N_3252);
nand U3494 (N_3494,N_3277,N_3266);
nand U3495 (N_3495,N_3326,N_3222);
xnor U3496 (N_3496,N_3255,N_3260);
or U3497 (N_3497,N_3237,N_3320);
or U3498 (N_3498,N_3340,N_3342);
nor U3499 (N_3499,N_3289,N_3240);
and U3500 (N_3500,N_3342,N_3225);
nor U3501 (N_3501,N_3258,N_3267);
or U3502 (N_3502,N_3243,N_3357);
nor U3503 (N_3503,N_3264,N_3247);
and U3504 (N_3504,N_3237,N_3338);
or U3505 (N_3505,N_3260,N_3254);
and U3506 (N_3506,N_3356,N_3290);
nand U3507 (N_3507,N_3217,N_3312);
nand U3508 (N_3508,N_3287,N_3215);
nor U3509 (N_3509,N_3331,N_3303);
nor U3510 (N_3510,N_3240,N_3239);
nor U3511 (N_3511,N_3329,N_3278);
nor U3512 (N_3512,N_3220,N_3230);
and U3513 (N_3513,N_3304,N_3339);
or U3514 (N_3514,N_3264,N_3352);
xor U3515 (N_3515,N_3233,N_3349);
nand U3516 (N_3516,N_3283,N_3244);
xor U3517 (N_3517,N_3358,N_3224);
nand U3518 (N_3518,N_3317,N_3351);
or U3519 (N_3519,N_3288,N_3299);
nand U3520 (N_3520,N_3503,N_3519);
nand U3521 (N_3521,N_3386,N_3368);
nand U3522 (N_3522,N_3422,N_3482);
or U3523 (N_3523,N_3456,N_3474);
nor U3524 (N_3524,N_3457,N_3518);
or U3525 (N_3525,N_3441,N_3383);
nor U3526 (N_3526,N_3483,N_3453);
xor U3527 (N_3527,N_3431,N_3396);
xor U3528 (N_3528,N_3487,N_3402);
xnor U3529 (N_3529,N_3390,N_3409);
xnor U3530 (N_3530,N_3364,N_3445);
or U3531 (N_3531,N_3363,N_3517);
nor U3532 (N_3532,N_3492,N_3362);
nor U3533 (N_3533,N_3384,N_3378);
and U3534 (N_3534,N_3451,N_3408);
nor U3535 (N_3535,N_3443,N_3476);
and U3536 (N_3536,N_3510,N_3361);
or U3537 (N_3537,N_3400,N_3387);
or U3538 (N_3538,N_3373,N_3395);
or U3539 (N_3539,N_3466,N_3494);
nor U3540 (N_3540,N_3480,N_3394);
nand U3541 (N_3541,N_3458,N_3420);
xnor U3542 (N_3542,N_3506,N_3484);
and U3543 (N_3543,N_3427,N_3432);
and U3544 (N_3544,N_3416,N_3478);
or U3545 (N_3545,N_3514,N_3392);
nand U3546 (N_3546,N_3374,N_3430);
and U3547 (N_3547,N_3398,N_3490);
xor U3548 (N_3548,N_3475,N_3469);
and U3549 (N_3549,N_3450,N_3468);
nand U3550 (N_3550,N_3435,N_3397);
nand U3551 (N_3551,N_3471,N_3455);
or U3552 (N_3552,N_3461,N_3516);
nor U3553 (N_3553,N_3372,N_3404);
or U3554 (N_3554,N_3459,N_3366);
nor U3555 (N_3555,N_3513,N_3485);
nor U3556 (N_3556,N_3470,N_3464);
and U3557 (N_3557,N_3417,N_3375);
xor U3558 (N_3558,N_3454,N_3412);
xnor U3559 (N_3559,N_3437,N_3495);
and U3560 (N_3560,N_3406,N_3436);
xnor U3561 (N_3561,N_3509,N_3410);
nand U3562 (N_3562,N_3380,N_3365);
nor U3563 (N_3563,N_3472,N_3421);
or U3564 (N_3564,N_3446,N_3442);
or U3565 (N_3565,N_3419,N_3389);
or U3566 (N_3566,N_3467,N_3393);
and U3567 (N_3567,N_3497,N_3488);
and U3568 (N_3568,N_3479,N_3415);
or U3569 (N_3569,N_3414,N_3433);
xnor U3570 (N_3570,N_3448,N_3444);
xor U3571 (N_3571,N_3418,N_3462);
or U3572 (N_3572,N_3388,N_3440);
or U3573 (N_3573,N_3411,N_3493);
nor U3574 (N_3574,N_3501,N_3385);
nor U3575 (N_3575,N_3379,N_3371);
xnor U3576 (N_3576,N_3429,N_3491);
and U3577 (N_3577,N_3370,N_3413);
and U3578 (N_3578,N_3481,N_3447);
nor U3579 (N_3579,N_3505,N_3498);
xor U3580 (N_3580,N_3425,N_3399);
nand U3581 (N_3581,N_3405,N_3381);
nor U3582 (N_3582,N_3401,N_3449);
and U3583 (N_3583,N_3507,N_3496);
xnor U3584 (N_3584,N_3403,N_3428);
xnor U3585 (N_3585,N_3376,N_3391);
or U3586 (N_3586,N_3367,N_3489);
and U3587 (N_3587,N_3438,N_3465);
nand U3588 (N_3588,N_3511,N_3407);
nand U3589 (N_3589,N_3504,N_3377);
or U3590 (N_3590,N_3434,N_3424);
and U3591 (N_3591,N_3512,N_3452);
nor U3592 (N_3592,N_3360,N_3460);
nor U3593 (N_3593,N_3499,N_3508);
nand U3594 (N_3594,N_3463,N_3382);
nand U3595 (N_3595,N_3486,N_3426);
nand U3596 (N_3596,N_3473,N_3439);
nor U3597 (N_3597,N_3500,N_3423);
xor U3598 (N_3598,N_3477,N_3515);
or U3599 (N_3599,N_3369,N_3502);
and U3600 (N_3600,N_3501,N_3367);
nor U3601 (N_3601,N_3377,N_3434);
xnor U3602 (N_3602,N_3409,N_3499);
and U3603 (N_3603,N_3384,N_3367);
xor U3604 (N_3604,N_3459,N_3417);
nor U3605 (N_3605,N_3494,N_3472);
or U3606 (N_3606,N_3440,N_3494);
and U3607 (N_3607,N_3389,N_3436);
or U3608 (N_3608,N_3370,N_3497);
and U3609 (N_3609,N_3362,N_3399);
or U3610 (N_3610,N_3375,N_3391);
nor U3611 (N_3611,N_3469,N_3466);
and U3612 (N_3612,N_3457,N_3459);
nand U3613 (N_3613,N_3456,N_3453);
or U3614 (N_3614,N_3505,N_3365);
nor U3615 (N_3615,N_3480,N_3375);
xnor U3616 (N_3616,N_3432,N_3475);
nor U3617 (N_3617,N_3471,N_3519);
nand U3618 (N_3618,N_3393,N_3461);
nand U3619 (N_3619,N_3486,N_3505);
or U3620 (N_3620,N_3379,N_3495);
xnor U3621 (N_3621,N_3440,N_3400);
nor U3622 (N_3622,N_3366,N_3402);
and U3623 (N_3623,N_3397,N_3447);
or U3624 (N_3624,N_3518,N_3477);
nor U3625 (N_3625,N_3383,N_3423);
nor U3626 (N_3626,N_3427,N_3499);
xor U3627 (N_3627,N_3435,N_3422);
and U3628 (N_3628,N_3494,N_3454);
nand U3629 (N_3629,N_3453,N_3407);
xor U3630 (N_3630,N_3430,N_3505);
xor U3631 (N_3631,N_3412,N_3378);
nor U3632 (N_3632,N_3478,N_3392);
and U3633 (N_3633,N_3515,N_3449);
nor U3634 (N_3634,N_3488,N_3412);
nor U3635 (N_3635,N_3507,N_3412);
nand U3636 (N_3636,N_3467,N_3367);
and U3637 (N_3637,N_3451,N_3394);
or U3638 (N_3638,N_3474,N_3473);
or U3639 (N_3639,N_3513,N_3451);
or U3640 (N_3640,N_3395,N_3435);
and U3641 (N_3641,N_3421,N_3365);
and U3642 (N_3642,N_3519,N_3505);
and U3643 (N_3643,N_3430,N_3480);
or U3644 (N_3644,N_3419,N_3423);
nor U3645 (N_3645,N_3409,N_3513);
nor U3646 (N_3646,N_3425,N_3362);
xnor U3647 (N_3647,N_3464,N_3510);
and U3648 (N_3648,N_3380,N_3459);
and U3649 (N_3649,N_3389,N_3382);
nor U3650 (N_3650,N_3396,N_3506);
nor U3651 (N_3651,N_3432,N_3377);
nor U3652 (N_3652,N_3491,N_3477);
or U3653 (N_3653,N_3374,N_3375);
or U3654 (N_3654,N_3504,N_3463);
or U3655 (N_3655,N_3474,N_3416);
xor U3656 (N_3656,N_3394,N_3459);
xor U3657 (N_3657,N_3417,N_3379);
and U3658 (N_3658,N_3432,N_3406);
nand U3659 (N_3659,N_3406,N_3500);
and U3660 (N_3660,N_3459,N_3476);
nand U3661 (N_3661,N_3378,N_3448);
xor U3662 (N_3662,N_3419,N_3404);
and U3663 (N_3663,N_3394,N_3493);
nor U3664 (N_3664,N_3465,N_3505);
and U3665 (N_3665,N_3412,N_3471);
nor U3666 (N_3666,N_3415,N_3396);
nor U3667 (N_3667,N_3480,N_3507);
nand U3668 (N_3668,N_3473,N_3376);
xor U3669 (N_3669,N_3435,N_3409);
or U3670 (N_3670,N_3382,N_3439);
and U3671 (N_3671,N_3378,N_3484);
and U3672 (N_3672,N_3480,N_3389);
nor U3673 (N_3673,N_3369,N_3379);
or U3674 (N_3674,N_3509,N_3432);
xnor U3675 (N_3675,N_3430,N_3490);
nor U3676 (N_3676,N_3403,N_3419);
and U3677 (N_3677,N_3469,N_3450);
or U3678 (N_3678,N_3410,N_3414);
and U3679 (N_3679,N_3452,N_3392);
nor U3680 (N_3680,N_3644,N_3649);
xnor U3681 (N_3681,N_3560,N_3625);
and U3682 (N_3682,N_3614,N_3586);
and U3683 (N_3683,N_3542,N_3606);
nand U3684 (N_3684,N_3627,N_3646);
nor U3685 (N_3685,N_3593,N_3562);
xnor U3686 (N_3686,N_3670,N_3595);
nand U3687 (N_3687,N_3654,N_3634);
nand U3688 (N_3688,N_3527,N_3538);
nand U3689 (N_3689,N_3666,N_3590);
and U3690 (N_3690,N_3569,N_3669);
nor U3691 (N_3691,N_3677,N_3665);
nand U3692 (N_3692,N_3647,N_3581);
or U3693 (N_3693,N_3672,N_3641);
nor U3694 (N_3694,N_3619,N_3667);
xor U3695 (N_3695,N_3628,N_3630);
and U3696 (N_3696,N_3624,N_3632);
nand U3697 (N_3697,N_3596,N_3631);
nor U3698 (N_3698,N_3531,N_3660);
nand U3699 (N_3699,N_3574,N_3663);
nor U3700 (N_3700,N_3570,N_3612);
nor U3701 (N_3701,N_3615,N_3592);
nand U3702 (N_3702,N_3608,N_3546);
and U3703 (N_3703,N_3658,N_3600);
nor U3704 (N_3704,N_3525,N_3544);
or U3705 (N_3705,N_3553,N_3543);
or U3706 (N_3706,N_3640,N_3635);
xnor U3707 (N_3707,N_3638,N_3603);
or U3708 (N_3708,N_3618,N_3626);
nor U3709 (N_3709,N_3617,N_3676);
xnor U3710 (N_3710,N_3583,N_3539);
xor U3711 (N_3711,N_3653,N_3594);
nor U3712 (N_3712,N_3616,N_3645);
xor U3713 (N_3713,N_3529,N_3550);
xnor U3714 (N_3714,N_3559,N_3648);
or U3715 (N_3715,N_3679,N_3637);
nand U3716 (N_3716,N_3673,N_3545);
and U3717 (N_3717,N_3613,N_3656);
nor U3718 (N_3718,N_3607,N_3587);
or U3719 (N_3719,N_3533,N_3573);
nand U3720 (N_3720,N_3530,N_3575);
nand U3721 (N_3721,N_3650,N_3622);
nand U3722 (N_3722,N_3671,N_3652);
or U3723 (N_3723,N_3551,N_3629);
xnor U3724 (N_3724,N_3623,N_3598);
or U3725 (N_3725,N_3566,N_3537);
nor U3726 (N_3726,N_3655,N_3582);
or U3727 (N_3727,N_3556,N_3661);
nor U3728 (N_3728,N_3521,N_3563);
nand U3729 (N_3729,N_3601,N_3534);
xnor U3730 (N_3730,N_3532,N_3651);
nand U3731 (N_3731,N_3675,N_3597);
or U3732 (N_3732,N_3576,N_3548);
nor U3733 (N_3733,N_3633,N_3552);
and U3734 (N_3734,N_3664,N_3540);
nand U3735 (N_3735,N_3659,N_3589);
or U3736 (N_3736,N_3526,N_3535);
and U3737 (N_3737,N_3584,N_3524);
and U3738 (N_3738,N_3528,N_3605);
or U3739 (N_3739,N_3621,N_3602);
xnor U3740 (N_3740,N_3668,N_3571);
or U3741 (N_3741,N_3558,N_3604);
and U3742 (N_3742,N_3636,N_3561);
nor U3743 (N_3743,N_3620,N_3557);
or U3744 (N_3744,N_3549,N_3577);
nor U3745 (N_3745,N_3554,N_3599);
xnor U3746 (N_3746,N_3588,N_3657);
or U3747 (N_3747,N_3610,N_3591);
nand U3748 (N_3748,N_3541,N_3520);
or U3749 (N_3749,N_3547,N_3555);
nand U3750 (N_3750,N_3678,N_3674);
nor U3751 (N_3751,N_3609,N_3585);
xnor U3752 (N_3752,N_3643,N_3639);
or U3753 (N_3753,N_3523,N_3572);
or U3754 (N_3754,N_3536,N_3567);
nor U3755 (N_3755,N_3578,N_3611);
or U3756 (N_3756,N_3522,N_3580);
or U3757 (N_3757,N_3579,N_3565);
and U3758 (N_3758,N_3568,N_3564);
xor U3759 (N_3759,N_3662,N_3642);
xor U3760 (N_3760,N_3666,N_3648);
xnor U3761 (N_3761,N_3525,N_3591);
or U3762 (N_3762,N_3608,N_3609);
or U3763 (N_3763,N_3624,N_3661);
or U3764 (N_3764,N_3637,N_3542);
and U3765 (N_3765,N_3663,N_3606);
and U3766 (N_3766,N_3648,N_3629);
and U3767 (N_3767,N_3569,N_3614);
nand U3768 (N_3768,N_3605,N_3552);
nor U3769 (N_3769,N_3606,N_3594);
nand U3770 (N_3770,N_3661,N_3601);
nand U3771 (N_3771,N_3606,N_3664);
xor U3772 (N_3772,N_3668,N_3589);
nand U3773 (N_3773,N_3575,N_3675);
xor U3774 (N_3774,N_3567,N_3538);
xor U3775 (N_3775,N_3662,N_3640);
xor U3776 (N_3776,N_3550,N_3647);
or U3777 (N_3777,N_3644,N_3662);
or U3778 (N_3778,N_3579,N_3615);
xnor U3779 (N_3779,N_3565,N_3525);
nor U3780 (N_3780,N_3528,N_3570);
and U3781 (N_3781,N_3583,N_3542);
and U3782 (N_3782,N_3644,N_3608);
nand U3783 (N_3783,N_3633,N_3637);
or U3784 (N_3784,N_3533,N_3601);
and U3785 (N_3785,N_3651,N_3618);
and U3786 (N_3786,N_3542,N_3665);
nor U3787 (N_3787,N_3611,N_3639);
nand U3788 (N_3788,N_3590,N_3521);
nor U3789 (N_3789,N_3579,N_3589);
nor U3790 (N_3790,N_3583,N_3659);
nor U3791 (N_3791,N_3676,N_3620);
nor U3792 (N_3792,N_3660,N_3618);
and U3793 (N_3793,N_3596,N_3633);
nor U3794 (N_3794,N_3613,N_3629);
or U3795 (N_3795,N_3626,N_3553);
nand U3796 (N_3796,N_3654,N_3582);
nor U3797 (N_3797,N_3606,N_3629);
xnor U3798 (N_3798,N_3628,N_3677);
or U3799 (N_3799,N_3594,N_3609);
and U3800 (N_3800,N_3662,N_3604);
and U3801 (N_3801,N_3656,N_3529);
nand U3802 (N_3802,N_3523,N_3582);
or U3803 (N_3803,N_3584,N_3551);
or U3804 (N_3804,N_3635,N_3659);
xnor U3805 (N_3805,N_3599,N_3629);
nand U3806 (N_3806,N_3592,N_3636);
xor U3807 (N_3807,N_3598,N_3640);
nand U3808 (N_3808,N_3538,N_3555);
or U3809 (N_3809,N_3677,N_3617);
and U3810 (N_3810,N_3620,N_3634);
xnor U3811 (N_3811,N_3544,N_3633);
nor U3812 (N_3812,N_3597,N_3547);
or U3813 (N_3813,N_3622,N_3662);
xnor U3814 (N_3814,N_3526,N_3540);
or U3815 (N_3815,N_3593,N_3546);
nor U3816 (N_3816,N_3536,N_3652);
or U3817 (N_3817,N_3562,N_3614);
or U3818 (N_3818,N_3589,N_3660);
or U3819 (N_3819,N_3625,N_3533);
xnor U3820 (N_3820,N_3547,N_3661);
or U3821 (N_3821,N_3675,N_3659);
xnor U3822 (N_3822,N_3595,N_3530);
and U3823 (N_3823,N_3520,N_3669);
nand U3824 (N_3824,N_3540,N_3559);
nand U3825 (N_3825,N_3606,N_3553);
or U3826 (N_3826,N_3645,N_3669);
xnor U3827 (N_3827,N_3587,N_3665);
and U3828 (N_3828,N_3650,N_3624);
xor U3829 (N_3829,N_3521,N_3542);
xor U3830 (N_3830,N_3668,N_3634);
nor U3831 (N_3831,N_3572,N_3542);
and U3832 (N_3832,N_3583,N_3647);
and U3833 (N_3833,N_3578,N_3589);
xor U3834 (N_3834,N_3618,N_3555);
nor U3835 (N_3835,N_3676,N_3554);
xor U3836 (N_3836,N_3574,N_3573);
xor U3837 (N_3837,N_3627,N_3534);
nor U3838 (N_3838,N_3594,N_3545);
nor U3839 (N_3839,N_3586,N_3578);
xnor U3840 (N_3840,N_3747,N_3737);
and U3841 (N_3841,N_3782,N_3733);
xnor U3842 (N_3842,N_3731,N_3805);
xnor U3843 (N_3843,N_3738,N_3797);
or U3844 (N_3844,N_3827,N_3777);
and U3845 (N_3845,N_3684,N_3839);
xor U3846 (N_3846,N_3740,N_3734);
nor U3847 (N_3847,N_3722,N_3801);
xnor U3848 (N_3848,N_3695,N_3811);
or U3849 (N_3849,N_3745,N_3688);
and U3850 (N_3850,N_3742,N_3808);
nor U3851 (N_3851,N_3735,N_3820);
and U3852 (N_3852,N_3714,N_3773);
or U3853 (N_3853,N_3824,N_3807);
nand U3854 (N_3854,N_3744,N_3709);
nand U3855 (N_3855,N_3703,N_3763);
nand U3856 (N_3856,N_3817,N_3831);
or U3857 (N_3857,N_3794,N_3757);
and U3858 (N_3858,N_3775,N_3727);
or U3859 (N_3859,N_3704,N_3691);
and U3860 (N_3860,N_3786,N_3761);
xor U3861 (N_3861,N_3739,N_3802);
xor U3862 (N_3862,N_3726,N_3702);
nor U3863 (N_3863,N_3751,N_3723);
or U3864 (N_3864,N_3715,N_3721);
and U3865 (N_3865,N_3810,N_3762);
or U3866 (N_3866,N_3765,N_3836);
and U3867 (N_3867,N_3708,N_3792);
xnor U3868 (N_3868,N_3685,N_3764);
or U3869 (N_3869,N_3711,N_3732);
nand U3870 (N_3870,N_3707,N_3683);
nand U3871 (N_3871,N_3793,N_3804);
xor U3872 (N_3872,N_3832,N_3795);
and U3873 (N_3873,N_3699,N_3686);
nor U3874 (N_3874,N_3717,N_3710);
nand U3875 (N_3875,N_3755,N_3779);
and U3876 (N_3876,N_3796,N_3694);
nor U3877 (N_3877,N_3736,N_3784);
nand U3878 (N_3878,N_3705,N_3692);
nand U3879 (N_3879,N_3799,N_3830);
xor U3880 (N_3880,N_3787,N_3769);
nand U3881 (N_3881,N_3767,N_3696);
or U3882 (N_3882,N_3772,N_3803);
and U3883 (N_3883,N_3785,N_3750);
nor U3884 (N_3884,N_3826,N_3835);
or U3885 (N_3885,N_3770,N_3754);
nand U3886 (N_3886,N_3680,N_3823);
nor U3887 (N_3887,N_3771,N_3806);
nor U3888 (N_3888,N_3838,N_3729);
and U3889 (N_3889,N_3822,N_3718);
or U3890 (N_3890,N_3752,N_3829);
nor U3891 (N_3891,N_3834,N_3816);
xor U3892 (N_3892,N_3706,N_3821);
nand U3893 (N_3893,N_3700,N_3687);
xnor U3894 (N_3894,N_3780,N_3812);
or U3895 (N_3895,N_3789,N_3716);
and U3896 (N_3896,N_3682,N_3701);
xor U3897 (N_3897,N_3809,N_3689);
nor U3898 (N_3898,N_3760,N_3790);
nor U3899 (N_3899,N_3698,N_3725);
or U3900 (N_3900,N_3798,N_3766);
nand U3901 (N_3901,N_3728,N_3758);
xnor U3902 (N_3902,N_3774,N_3720);
or U3903 (N_3903,N_3713,N_3746);
and U3904 (N_3904,N_3814,N_3693);
nor U3905 (N_3905,N_3768,N_3724);
and U3906 (N_3906,N_3833,N_3788);
and U3907 (N_3907,N_3818,N_3756);
and U3908 (N_3908,N_3819,N_3681);
nor U3909 (N_3909,N_3690,N_3815);
nand U3910 (N_3910,N_3837,N_3828);
xor U3911 (N_3911,N_3759,N_3781);
xnor U3912 (N_3912,N_3800,N_3778);
nor U3913 (N_3913,N_3791,N_3741);
nor U3914 (N_3914,N_3748,N_3753);
or U3915 (N_3915,N_3743,N_3719);
xor U3916 (N_3916,N_3813,N_3749);
or U3917 (N_3917,N_3730,N_3825);
nor U3918 (N_3918,N_3783,N_3776);
or U3919 (N_3919,N_3712,N_3697);
or U3920 (N_3920,N_3790,N_3695);
nand U3921 (N_3921,N_3800,N_3796);
xnor U3922 (N_3922,N_3766,N_3796);
nand U3923 (N_3923,N_3720,N_3807);
xnor U3924 (N_3924,N_3735,N_3721);
and U3925 (N_3925,N_3787,N_3754);
nand U3926 (N_3926,N_3749,N_3792);
and U3927 (N_3927,N_3683,N_3831);
nand U3928 (N_3928,N_3801,N_3798);
and U3929 (N_3929,N_3802,N_3681);
xor U3930 (N_3930,N_3782,N_3721);
nor U3931 (N_3931,N_3720,N_3777);
xnor U3932 (N_3932,N_3711,N_3713);
or U3933 (N_3933,N_3800,N_3813);
nor U3934 (N_3934,N_3770,N_3714);
xnor U3935 (N_3935,N_3738,N_3745);
and U3936 (N_3936,N_3739,N_3755);
nand U3937 (N_3937,N_3732,N_3730);
or U3938 (N_3938,N_3791,N_3797);
and U3939 (N_3939,N_3800,N_3821);
or U3940 (N_3940,N_3708,N_3739);
nand U3941 (N_3941,N_3680,N_3702);
nand U3942 (N_3942,N_3767,N_3713);
or U3943 (N_3943,N_3717,N_3737);
or U3944 (N_3944,N_3807,N_3735);
nand U3945 (N_3945,N_3696,N_3813);
xnor U3946 (N_3946,N_3743,N_3817);
or U3947 (N_3947,N_3756,N_3732);
and U3948 (N_3948,N_3701,N_3831);
nand U3949 (N_3949,N_3689,N_3754);
nor U3950 (N_3950,N_3688,N_3724);
or U3951 (N_3951,N_3776,N_3793);
or U3952 (N_3952,N_3705,N_3703);
or U3953 (N_3953,N_3833,N_3682);
and U3954 (N_3954,N_3796,N_3764);
xor U3955 (N_3955,N_3776,N_3731);
nand U3956 (N_3956,N_3727,N_3688);
or U3957 (N_3957,N_3691,N_3819);
nor U3958 (N_3958,N_3815,N_3725);
nand U3959 (N_3959,N_3738,N_3770);
nor U3960 (N_3960,N_3730,N_3804);
xor U3961 (N_3961,N_3824,N_3705);
or U3962 (N_3962,N_3794,N_3773);
xnor U3963 (N_3963,N_3687,N_3692);
or U3964 (N_3964,N_3783,N_3750);
or U3965 (N_3965,N_3721,N_3682);
nand U3966 (N_3966,N_3831,N_3813);
xnor U3967 (N_3967,N_3741,N_3787);
nor U3968 (N_3968,N_3802,N_3750);
or U3969 (N_3969,N_3809,N_3761);
or U3970 (N_3970,N_3818,N_3770);
and U3971 (N_3971,N_3798,N_3695);
xor U3972 (N_3972,N_3746,N_3777);
or U3973 (N_3973,N_3714,N_3732);
xor U3974 (N_3974,N_3695,N_3690);
nand U3975 (N_3975,N_3756,N_3762);
nor U3976 (N_3976,N_3721,N_3783);
and U3977 (N_3977,N_3837,N_3818);
xnor U3978 (N_3978,N_3832,N_3793);
nor U3979 (N_3979,N_3797,N_3688);
or U3980 (N_3980,N_3824,N_3803);
and U3981 (N_3981,N_3813,N_3787);
and U3982 (N_3982,N_3691,N_3777);
and U3983 (N_3983,N_3717,N_3796);
xor U3984 (N_3984,N_3689,N_3764);
and U3985 (N_3985,N_3715,N_3742);
xnor U3986 (N_3986,N_3718,N_3768);
nand U3987 (N_3987,N_3771,N_3780);
nor U3988 (N_3988,N_3690,N_3817);
nand U3989 (N_3989,N_3736,N_3742);
and U3990 (N_3990,N_3810,N_3770);
nor U3991 (N_3991,N_3711,N_3698);
nand U3992 (N_3992,N_3779,N_3696);
xor U3993 (N_3993,N_3683,N_3828);
nand U3994 (N_3994,N_3819,N_3753);
and U3995 (N_3995,N_3817,N_3727);
or U3996 (N_3996,N_3818,N_3715);
nor U3997 (N_3997,N_3707,N_3835);
or U3998 (N_3998,N_3781,N_3760);
nor U3999 (N_3999,N_3794,N_3755);
and U4000 (N_4000,N_3874,N_3965);
nand U4001 (N_4001,N_3876,N_3982);
or U4002 (N_4002,N_3992,N_3906);
or U4003 (N_4003,N_3958,N_3841);
xor U4004 (N_4004,N_3868,N_3864);
nand U4005 (N_4005,N_3998,N_3974);
xor U4006 (N_4006,N_3930,N_3909);
xnor U4007 (N_4007,N_3846,N_3863);
and U4008 (N_4008,N_3994,N_3946);
and U4009 (N_4009,N_3850,N_3987);
and U4010 (N_4010,N_3883,N_3953);
nor U4011 (N_4011,N_3933,N_3960);
and U4012 (N_4012,N_3879,N_3921);
and U4013 (N_4013,N_3967,N_3914);
and U4014 (N_4014,N_3927,N_3975);
nand U4015 (N_4015,N_3870,N_3912);
and U4016 (N_4016,N_3978,N_3949);
nor U4017 (N_4017,N_3993,N_3943);
nand U4018 (N_4018,N_3976,N_3861);
nand U4019 (N_4019,N_3904,N_3897);
nor U4020 (N_4020,N_3971,N_3935);
xor U4021 (N_4021,N_3924,N_3884);
and U4022 (N_4022,N_3881,N_3867);
and U4023 (N_4023,N_3918,N_3979);
nand U4024 (N_4024,N_3968,N_3858);
or U4025 (N_4025,N_3886,N_3937);
and U4026 (N_4026,N_3893,N_3917);
nor U4027 (N_4027,N_3888,N_3931);
nor U4028 (N_4028,N_3847,N_3911);
nand U4029 (N_4029,N_3894,N_3969);
xor U4030 (N_4030,N_3887,N_3980);
or U4031 (N_4031,N_3908,N_3889);
and U4032 (N_4032,N_3973,N_3928);
and U4033 (N_4033,N_3896,N_3860);
xnor U4034 (N_4034,N_3862,N_3986);
and U4035 (N_4035,N_3855,N_3934);
nor U4036 (N_4036,N_3856,N_3916);
nor U4037 (N_4037,N_3952,N_3892);
xor U4038 (N_4038,N_3984,N_3901);
nor U4039 (N_4039,N_3890,N_3851);
or U4040 (N_4040,N_3852,N_3995);
xnor U4041 (N_4041,N_3865,N_3843);
and U4042 (N_4042,N_3880,N_3972);
or U4043 (N_4043,N_3991,N_3942);
nand U4044 (N_4044,N_3898,N_3985);
nor U4045 (N_4045,N_3920,N_3989);
and U4046 (N_4046,N_3966,N_3899);
nand U4047 (N_4047,N_3996,N_3923);
nand U4048 (N_4048,N_3877,N_3866);
and U4049 (N_4049,N_3939,N_3955);
and U4050 (N_4050,N_3945,N_3910);
and U4051 (N_4051,N_3845,N_3873);
nor U4052 (N_4052,N_3957,N_3900);
nor U4053 (N_4053,N_3988,N_3940);
and U4054 (N_4054,N_3956,N_3871);
nor U4055 (N_4055,N_3962,N_3882);
and U4056 (N_4056,N_3961,N_3885);
or U4057 (N_4057,N_3907,N_3891);
nor U4058 (N_4058,N_3936,N_3954);
nand U4059 (N_4059,N_3959,N_3999);
or U4060 (N_4060,N_3950,N_3947);
and U4061 (N_4061,N_3983,N_3857);
and U4062 (N_4062,N_3951,N_3913);
or U4063 (N_4063,N_3922,N_3929);
and U4064 (N_4064,N_3854,N_3840);
nor U4065 (N_4065,N_3948,N_3997);
xor U4066 (N_4066,N_3963,N_3915);
and U4067 (N_4067,N_3970,N_3905);
or U4068 (N_4068,N_3875,N_3919);
nor U4069 (N_4069,N_3926,N_3941);
and U4070 (N_4070,N_3938,N_3859);
xnor U4071 (N_4071,N_3849,N_3932);
xnor U4072 (N_4072,N_3977,N_3848);
xor U4073 (N_4073,N_3844,N_3981);
nor U4074 (N_4074,N_3964,N_3944);
or U4075 (N_4075,N_3869,N_3878);
nor U4076 (N_4076,N_3925,N_3990);
nor U4077 (N_4077,N_3842,N_3902);
xnor U4078 (N_4078,N_3872,N_3903);
nand U4079 (N_4079,N_3853,N_3895);
and U4080 (N_4080,N_3886,N_3985);
xor U4081 (N_4081,N_3976,N_3908);
nand U4082 (N_4082,N_3921,N_3843);
and U4083 (N_4083,N_3976,N_3996);
and U4084 (N_4084,N_3899,N_3901);
and U4085 (N_4085,N_3919,N_3890);
xor U4086 (N_4086,N_3910,N_3959);
or U4087 (N_4087,N_3853,N_3904);
and U4088 (N_4088,N_3991,N_3907);
nand U4089 (N_4089,N_3970,N_3886);
and U4090 (N_4090,N_3868,N_3856);
nand U4091 (N_4091,N_3932,N_3964);
nand U4092 (N_4092,N_3954,N_3962);
nor U4093 (N_4093,N_3973,N_3850);
xnor U4094 (N_4094,N_3864,N_3943);
or U4095 (N_4095,N_3895,N_3974);
nor U4096 (N_4096,N_3884,N_3986);
or U4097 (N_4097,N_3917,N_3928);
or U4098 (N_4098,N_3915,N_3946);
nand U4099 (N_4099,N_3953,N_3874);
nand U4100 (N_4100,N_3876,N_3975);
xor U4101 (N_4101,N_3931,N_3945);
xor U4102 (N_4102,N_3984,N_3877);
nor U4103 (N_4103,N_3921,N_3887);
nor U4104 (N_4104,N_3972,N_3850);
nand U4105 (N_4105,N_3951,N_3974);
or U4106 (N_4106,N_3892,N_3983);
nor U4107 (N_4107,N_3911,N_3979);
xor U4108 (N_4108,N_3990,N_3880);
and U4109 (N_4109,N_3986,N_3892);
nand U4110 (N_4110,N_3912,N_3842);
or U4111 (N_4111,N_3971,N_3890);
or U4112 (N_4112,N_3875,N_3924);
and U4113 (N_4113,N_3939,N_3897);
xor U4114 (N_4114,N_3902,N_3845);
nand U4115 (N_4115,N_3955,N_3896);
xnor U4116 (N_4116,N_3899,N_3847);
or U4117 (N_4117,N_3879,N_3840);
or U4118 (N_4118,N_3921,N_3947);
and U4119 (N_4119,N_3980,N_3848);
or U4120 (N_4120,N_3970,N_3932);
and U4121 (N_4121,N_3844,N_3921);
nor U4122 (N_4122,N_3998,N_3899);
and U4123 (N_4123,N_3846,N_3899);
nand U4124 (N_4124,N_3908,N_3941);
xor U4125 (N_4125,N_3910,N_3971);
or U4126 (N_4126,N_3954,N_3856);
nand U4127 (N_4127,N_3872,N_3846);
xor U4128 (N_4128,N_3935,N_3989);
xor U4129 (N_4129,N_3862,N_3902);
or U4130 (N_4130,N_3851,N_3992);
xor U4131 (N_4131,N_3885,N_3933);
nand U4132 (N_4132,N_3944,N_3993);
or U4133 (N_4133,N_3978,N_3860);
nand U4134 (N_4134,N_3895,N_3971);
nor U4135 (N_4135,N_3888,N_3881);
or U4136 (N_4136,N_3991,N_3957);
and U4137 (N_4137,N_3845,N_3951);
and U4138 (N_4138,N_3971,N_3840);
nor U4139 (N_4139,N_3945,N_3879);
xor U4140 (N_4140,N_3939,N_3937);
or U4141 (N_4141,N_3963,N_3943);
and U4142 (N_4142,N_3982,N_3916);
xor U4143 (N_4143,N_3920,N_3870);
nand U4144 (N_4144,N_3951,N_3843);
or U4145 (N_4145,N_3961,N_3903);
nand U4146 (N_4146,N_3897,N_3989);
xnor U4147 (N_4147,N_3970,N_3927);
or U4148 (N_4148,N_3860,N_3941);
xor U4149 (N_4149,N_3882,N_3892);
nand U4150 (N_4150,N_3852,N_3854);
nor U4151 (N_4151,N_3932,N_3853);
nand U4152 (N_4152,N_3854,N_3977);
or U4153 (N_4153,N_3948,N_3926);
nor U4154 (N_4154,N_3932,N_3984);
xnor U4155 (N_4155,N_3888,N_3922);
and U4156 (N_4156,N_3952,N_3864);
xnor U4157 (N_4157,N_3888,N_3843);
or U4158 (N_4158,N_3966,N_3970);
nand U4159 (N_4159,N_3849,N_3840);
xor U4160 (N_4160,N_4001,N_4029);
and U4161 (N_4161,N_4135,N_4014);
nor U4162 (N_4162,N_4088,N_4136);
xnor U4163 (N_4163,N_4087,N_4049);
or U4164 (N_4164,N_4051,N_4028);
xnor U4165 (N_4165,N_4013,N_4040);
xor U4166 (N_4166,N_4070,N_4124);
nor U4167 (N_4167,N_4101,N_4003);
or U4168 (N_4168,N_4023,N_4039);
nand U4169 (N_4169,N_4033,N_4099);
or U4170 (N_4170,N_4021,N_4133);
nor U4171 (N_4171,N_4153,N_4017);
or U4172 (N_4172,N_4007,N_4060);
or U4173 (N_4173,N_4005,N_4144);
nand U4174 (N_4174,N_4065,N_4147);
xor U4175 (N_4175,N_4116,N_4076);
or U4176 (N_4176,N_4043,N_4139);
nand U4177 (N_4177,N_4159,N_4156);
nor U4178 (N_4178,N_4082,N_4027);
nor U4179 (N_4179,N_4069,N_4015);
xnor U4180 (N_4180,N_4074,N_4010);
nor U4181 (N_4181,N_4091,N_4000);
or U4182 (N_4182,N_4096,N_4157);
and U4183 (N_4183,N_4057,N_4036);
or U4184 (N_4184,N_4058,N_4155);
or U4185 (N_4185,N_4104,N_4146);
nor U4186 (N_4186,N_4067,N_4042);
xnor U4187 (N_4187,N_4075,N_4034);
and U4188 (N_4188,N_4105,N_4110);
nand U4189 (N_4189,N_4011,N_4020);
xor U4190 (N_4190,N_4063,N_4052);
xor U4191 (N_4191,N_4120,N_4064);
and U4192 (N_4192,N_4107,N_4078);
xor U4193 (N_4193,N_4055,N_4123);
and U4194 (N_4194,N_4152,N_4083);
nand U4195 (N_4195,N_4138,N_4031);
or U4196 (N_4196,N_4117,N_4061);
or U4197 (N_4197,N_4080,N_4130);
and U4198 (N_4198,N_4054,N_4046);
nor U4199 (N_4199,N_4103,N_4073);
xor U4200 (N_4200,N_4112,N_4114);
or U4201 (N_4201,N_4094,N_4095);
or U4202 (N_4202,N_4097,N_4149);
or U4203 (N_4203,N_4018,N_4090);
or U4204 (N_4204,N_4012,N_4098);
or U4205 (N_4205,N_4053,N_4071);
and U4206 (N_4206,N_4030,N_4092);
or U4207 (N_4207,N_4038,N_4006);
or U4208 (N_4208,N_4158,N_4068);
xor U4209 (N_4209,N_4131,N_4025);
nand U4210 (N_4210,N_4145,N_4037);
or U4211 (N_4211,N_4143,N_4148);
and U4212 (N_4212,N_4140,N_4128);
and U4213 (N_4213,N_4137,N_4026);
nand U4214 (N_4214,N_4008,N_4016);
xor U4215 (N_4215,N_4121,N_4024);
nand U4216 (N_4216,N_4066,N_4113);
or U4217 (N_4217,N_4141,N_4111);
nor U4218 (N_4218,N_4127,N_4109);
xor U4219 (N_4219,N_4119,N_4059);
nor U4220 (N_4220,N_4079,N_4072);
nor U4221 (N_4221,N_4093,N_4084);
or U4222 (N_4222,N_4041,N_4129);
nand U4223 (N_4223,N_4004,N_4142);
and U4224 (N_4224,N_4032,N_4047);
nand U4225 (N_4225,N_4108,N_4002);
and U4226 (N_4226,N_4115,N_4089);
nand U4227 (N_4227,N_4125,N_4132);
nor U4228 (N_4228,N_4019,N_4077);
nor U4229 (N_4229,N_4081,N_4126);
xnor U4230 (N_4230,N_4118,N_4134);
nor U4231 (N_4231,N_4106,N_4048);
nor U4232 (N_4232,N_4062,N_4044);
or U4233 (N_4233,N_4154,N_4009);
and U4234 (N_4234,N_4086,N_4100);
xor U4235 (N_4235,N_4045,N_4056);
and U4236 (N_4236,N_4022,N_4102);
and U4237 (N_4237,N_4050,N_4035);
nor U4238 (N_4238,N_4150,N_4085);
xor U4239 (N_4239,N_4151,N_4122);
nand U4240 (N_4240,N_4043,N_4131);
and U4241 (N_4241,N_4008,N_4159);
and U4242 (N_4242,N_4051,N_4042);
or U4243 (N_4243,N_4039,N_4047);
xor U4244 (N_4244,N_4028,N_4023);
and U4245 (N_4245,N_4066,N_4135);
or U4246 (N_4246,N_4116,N_4001);
nand U4247 (N_4247,N_4157,N_4080);
or U4248 (N_4248,N_4008,N_4148);
nor U4249 (N_4249,N_4069,N_4071);
xor U4250 (N_4250,N_4082,N_4116);
xnor U4251 (N_4251,N_4008,N_4071);
nand U4252 (N_4252,N_4126,N_4002);
xnor U4253 (N_4253,N_4116,N_4152);
nor U4254 (N_4254,N_4054,N_4117);
nand U4255 (N_4255,N_4075,N_4017);
nor U4256 (N_4256,N_4021,N_4117);
nand U4257 (N_4257,N_4114,N_4068);
or U4258 (N_4258,N_4018,N_4031);
xnor U4259 (N_4259,N_4017,N_4039);
and U4260 (N_4260,N_4118,N_4057);
and U4261 (N_4261,N_4143,N_4155);
and U4262 (N_4262,N_4145,N_4156);
or U4263 (N_4263,N_4059,N_4090);
xor U4264 (N_4264,N_4089,N_4031);
or U4265 (N_4265,N_4010,N_4148);
nand U4266 (N_4266,N_4057,N_4107);
and U4267 (N_4267,N_4157,N_4068);
nand U4268 (N_4268,N_4121,N_4119);
or U4269 (N_4269,N_4073,N_4108);
xor U4270 (N_4270,N_4095,N_4045);
xnor U4271 (N_4271,N_4028,N_4072);
and U4272 (N_4272,N_4004,N_4144);
and U4273 (N_4273,N_4125,N_4063);
xor U4274 (N_4274,N_4080,N_4125);
xor U4275 (N_4275,N_4008,N_4033);
and U4276 (N_4276,N_4096,N_4156);
nand U4277 (N_4277,N_4022,N_4089);
and U4278 (N_4278,N_4009,N_4113);
and U4279 (N_4279,N_4045,N_4104);
and U4280 (N_4280,N_4005,N_4103);
or U4281 (N_4281,N_4025,N_4013);
or U4282 (N_4282,N_4044,N_4066);
nand U4283 (N_4283,N_4000,N_4069);
or U4284 (N_4284,N_4057,N_4149);
nor U4285 (N_4285,N_4051,N_4014);
nor U4286 (N_4286,N_4018,N_4123);
or U4287 (N_4287,N_4064,N_4049);
or U4288 (N_4288,N_4101,N_4002);
nor U4289 (N_4289,N_4082,N_4125);
nand U4290 (N_4290,N_4074,N_4069);
nor U4291 (N_4291,N_4053,N_4095);
nor U4292 (N_4292,N_4068,N_4131);
nor U4293 (N_4293,N_4086,N_4156);
and U4294 (N_4294,N_4008,N_4086);
and U4295 (N_4295,N_4055,N_4064);
and U4296 (N_4296,N_4029,N_4081);
or U4297 (N_4297,N_4004,N_4043);
nand U4298 (N_4298,N_4140,N_4037);
nor U4299 (N_4299,N_4128,N_4139);
nand U4300 (N_4300,N_4047,N_4014);
nor U4301 (N_4301,N_4027,N_4000);
nor U4302 (N_4302,N_4050,N_4010);
and U4303 (N_4303,N_4105,N_4084);
nor U4304 (N_4304,N_4026,N_4146);
nand U4305 (N_4305,N_4131,N_4134);
or U4306 (N_4306,N_4003,N_4059);
xor U4307 (N_4307,N_4139,N_4071);
nand U4308 (N_4308,N_4136,N_4000);
nor U4309 (N_4309,N_4124,N_4091);
or U4310 (N_4310,N_4023,N_4079);
nand U4311 (N_4311,N_4069,N_4059);
nor U4312 (N_4312,N_4078,N_4037);
nor U4313 (N_4313,N_4148,N_4103);
nand U4314 (N_4314,N_4034,N_4086);
and U4315 (N_4315,N_4002,N_4150);
nand U4316 (N_4316,N_4048,N_4081);
and U4317 (N_4317,N_4098,N_4007);
xnor U4318 (N_4318,N_4054,N_4044);
nand U4319 (N_4319,N_4038,N_4095);
xnor U4320 (N_4320,N_4303,N_4170);
nand U4321 (N_4321,N_4188,N_4184);
nor U4322 (N_4322,N_4160,N_4180);
xnor U4323 (N_4323,N_4205,N_4276);
xnor U4324 (N_4324,N_4247,N_4268);
and U4325 (N_4325,N_4306,N_4311);
nor U4326 (N_4326,N_4166,N_4296);
nand U4327 (N_4327,N_4244,N_4187);
nand U4328 (N_4328,N_4213,N_4316);
or U4329 (N_4329,N_4236,N_4194);
nand U4330 (N_4330,N_4183,N_4208);
or U4331 (N_4331,N_4186,N_4231);
and U4332 (N_4332,N_4318,N_4307);
or U4333 (N_4333,N_4210,N_4241);
or U4334 (N_4334,N_4288,N_4227);
nor U4335 (N_4335,N_4298,N_4255);
and U4336 (N_4336,N_4262,N_4193);
xor U4337 (N_4337,N_4226,N_4238);
nand U4338 (N_4338,N_4219,N_4295);
and U4339 (N_4339,N_4237,N_4191);
nor U4340 (N_4340,N_4216,N_4248);
nand U4341 (N_4341,N_4232,N_4289);
and U4342 (N_4342,N_4212,N_4284);
xor U4343 (N_4343,N_4315,N_4286);
or U4344 (N_4344,N_4310,N_4235);
nand U4345 (N_4345,N_4175,N_4196);
nor U4346 (N_4346,N_4275,N_4249);
and U4347 (N_4347,N_4206,N_4274);
xnor U4348 (N_4348,N_4304,N_4234);
nand U4349 (N_4349,N_4280,N_4269);
and U4350 (N_4350,N_4305,N_4259);
nand U4351 (N_4351,N_4181,N_4252);
or U4352 (N_4352,N_4256,N_4228);
nor U4353 (N_4353,N_4198,N_4177);
and U4354 (N_4354,N_4197,N_4242);
and U4355 (N_4355,N_4204,N_4167);
and U4356 (N_4356,N_4199,N_4190);
nand U4357 (N_4357,N_4253,N_4270);
xnor U4358 (N_4358,N_4192,N_4182);
xor U4359 (N_4359,N_4299,N_4287);
xnor U4360 (N_4360,N_4201,N_4265);
xnor U4361 (N_4361,N_4223,N_4277);
nor U4362 (N_4362,N_4300,N_4195);
nand U4363 (N_4363,N_4239,N_4221);
nand U4364 (N_4364,N_4207,N_4220);
nor U4365 (N_4365,N_4251,N_4168);
nand U4366 (N_4366,N_4285,N_4172);
xnor U4367 (N_4367,N_4161,N_4250);
xnor U4368 (N_4368,N_4271,N_4189);
xor U4369 (N_4369,N_4257,N_4282);
or U4370 (N_4370,N_4222,N_4174);
nand U4371 (N_4371,N_4162,N_4245);
and U4372 (N_4372,N_4261,N_4279);
nor U4373 (N_4373,N_4229,N_4246);
nor U4374 (N_4374,N_4293,N_4179);
and U4375 (N_4375,N_4215,N_4165);
nor U4376 (N_4376,N_4173,N_4211);
nor U4377 (N_4377,N_4258,N_4171);
xnor U4378 (N_4378,N_4202,N_4164);
nand U4379 (N_4379,N_4178,N_4176);
nand U4380 (N_4380,N_4209,N_4224);
or U4381 (N_4381,N_4260,N_4281);
or U4382 (N_4382,N_4273,N_4266);
or U4383 (N_4383,N_4264,N_4230);
or U4384 (N_4384,N_4254,N_4200);
or U4385 (N_4385,N_4263,N_4313);
and U4386 (N_4386,N_4309,N_4301);
and U4387 (N_4387,N_4225,N_4243);
nand U4388 (N_4388,N_4214,N_4317);
and U4389 (N_4389,N_4302,N_4312);
nand U4390 (N_4390,N_4297,N_4240);
nor U4391 (N_4391,N_4283,N_4233);
nand U4392 (N_4392,N_4290,N_4217);
and U4393 (N_4393,N_4292,N_4185);
nand U4394 (N_4394,N_4314,N_4308);
and U4395 (N_4395,N_4163,N_4169);
nor U4396 (N_4396,N_4291,N_4267);
nor U4397 (N_4397,N_4272,N_4218);
or U4398 (N_4398,N_4278,N_4319);
and U4399 (N_4399,N_4294,N_4203);
nand U4400 (N_4400,N_4250,N_4252);
or U4401 (N_4401,N_4277,N_4209);
and U4402 (N_4402,N_4200,N_4285);
or U4403 (N_4403,N_4265,N_4242);
nor U4404 (N_4404,N_4192,N_4291);
nand U4405 (N_4405,N_4229,N_4282);
or U4406 (N_4406,N_4233,N_4194);
and U4407 (N_4407,N_4194,N_4213);
xnor U4408 (N_4408,N_4283,N_4216);
xnor U4409 (N_4409,N_4246,N_4165);
nand U4410 (N_4410,N_4281,N_4230);
nand U4411 (N_4411,N_4168,N_4299);
nand U4412 (N_4412,N_4190,N_4181);
nand U4413 (N_4413,N_4302,N_4226);
or U4414 (N_4414,N_4184,N_4228);
or U4415 (N_4415,N_4242,N_4314);
and U4416 (N_4416,N_4222,N_4178);
and U4417 (N_4417,N_4230,N_4195);
and U4418 (N_4418,N_4266,N_4315);
nand U4419 (N_4419,N_4248,N_4249);
and U4420 (N_4420,N_4232,N_4240);
xor U4421 (N_4421,N_4237,N_4272);
or U4422 (N_4422,N_4245,N_4164);
nand U4423 (N_4423,N_4223,N_4197);
nand U4424 (N_4424,N_4228,N_4179);
xnor U4425 (N_4425,N_4232,N_4247);
xnor U4426 (N_4426,N_4207,N_4307);
nor U4427 (N_4427,N_4245,N_4261);
or U4428 (N_4428,N_4318,N_4282);
nor U4429 (N_4429,N_4306,N_4220);
nand U4430 (N_4430,N_4302,N_4221);
or U4431 (N_4431,N_4199,N_4296);
or U4432 (N_4432,N_4175,N_4163);
and U4433 (N_4433,N_4188,N_4181);
nand U4434 (N_4434,N_4178,N_4263);
or U4435 (N_4435,N_4257,N_4184);
and U4436 (N_4436,N_4204,N_4319);
nand U4437 (N_4437,N_4244,N_4197);
xnor U4438 (N_4438,N_4315,N_4244);
nand U4439 (N_4439,N_4220,N_4211);
nand U4440 (N_4440,N_4164,N_4199);
or U4441 (N_4441,N_4179,N_4246);
and U4442 (N_4442,N_4259,N_4207);
nor U4443 (N_4443,N_4246,N_4278);
xor U4444 (N_4444,N_4232,N_4253);
xor U4445 (N_4445,N_4284,N_4296);
nand U4446 (N_4446,N_4314,N_4166);
nand U4447 (N_4447,N_4200,N_4229);
xnor U4448 (N_4448,N_4186,N_4252);
nand U4449 (N_4449,N_4253,N_4317);
nor U4450 (N_4450,N_4213,N_4196);
nor U4451 (N_4451,N_4247,N_4289);
and U4452 (N_4452,N_4249,N_4258);
xor U4453 (N_4453,N_4306,N_4293);
nor U4454 (N_4454,N_4168,N_4301);
nand U4455 (N_4455,N_4284,N_4217);
or U4456 (N_4456,N_4285,N_4244);
xnor U4457 (N_4457,N_4175,N_4208);
and U4458 (N_4458,N_4261,N_4207);
or U4459 (N_4459,N_4249,N_4294);
and U4460 (N_4460,N_4184,N_4206);
xnor U4461 (N_4461,N_4170,N_4193);
nor U4462 (N_4462,N_4308,N_4183);
and U4463 (N_4463,N_4211,N_4291);
nand U4464 (N_4464,N_4300,N_4311);
or U4465 (N_4465,N_4187,N_4178);
nand U4466 (N_4466,N_4223,N_4260);
or U4467 (N_4467,N_4229,N_4299);
nor U4468 (N_4468,N_4184,N_4288);
xnor U4469 (N_4469,N_4281,N_4183);
and U4470 (N_4470,N_4313,N_4255);
nand U4471 (N_4471,N_4253,N_4273);
and U4472 (N_4472,N_4189,N_4303);
nor U4473 (N_4473,N_4295,N_4165);
xnor U4474 (N_4474,N_4319,N_4302);
nor U4475 (N_4475,N_4219,N_4178);
nor U4476 (N_4476,N_4226,N_4277);
nor U4477 (N_4477,N_4187,N_4263);
xor U4478 (N_4478,N_4309,N_4232);
and U4479 (N_4479,N_4267,N_4167);
and U4480 (N_4480,N_4408,N_4320);
xnor U4481 (N_4481,N_4359,N_4327);
nand U4482 (N_4482,N_4354,N_4405);
nand U4483 (N_4483,N_4334,N_4345);
xnor U4484 (N_4484,N_4355,N_4409);
or U4485 (N_4485,N_4365,N_4422);
nand U4486 (N_4486,N_4472,N_4349);
nand U4487 (N_4487,N_4460,N_4437);
and U4488 (N_4488,N_4439,N_4335);
xnor U4489 (N_4489,N_4464,N_4333);
nor U4490 (N_4490,N_4469,N_4465);
nand U4491 (N_4491,N_4398,N_4382);
xnor U4492 (N_4492,N_4364,N_4338);
and U4493 (N_4493,N_4410,N_4376);
nor U4494 (N_4494,N_4384,N_4407);
or U4495 (N_4495,N_4476,N_4462);
and U4496 (N_4496,N_4336,N_4411);
nor U4497 (N_4497,N_4420,N_4323);
and U4498 (N_4498,N_4450,N_4385);
or U4499 (N_4499,N_4377,N_4378);
xnor U4500 (N_4500,N_4325,N_4428);
xor U4501 (N_4501,N_4399,N_4374);
xnor U4502 (N_4502,N_4401,N_4386);
nand U4503 (N_4503,N_4413,N_4415);
and U4504 (N_4504,N_4447,N_4449);
or U4505 (N_4505,N_4458,N_4397);
and U4506 (N_4506,N_4389,N_4388);
xnor U4507 (N_4507,N_4443,N_4412);
xor U4508 (N_4508,N_4416,N_4348);
or U4509 (N_4509,N_4375,N_4463);
nor U4510 (N_4510,N_4356,N_4360);
or U4511 (N_4511,N_4340,N_4326);
xor U4512 (N_4512,N_4442,N_4471);
xor U4513 (N_4513,N_4434,N_4381);
nor U4514 (N_4514,N_4448,N_4431);
nor U4515 (N_4515,N_4372,N_4478);
nand U4516 (N_4516,N_4368,N_4324);
nor U4517 (N_4517,N_4435,N_4454);
or U4518 (N_4518,N_4370,N_4363);
xor U4519 (N_4519,N_4427,N_4466);
xor U4520 (N_4520,N_4351,N_4426);
nor U4521 (N_4521,N_4470,N_4337);
or U4522 (N_4522,N_4475,N_4441);
xnor U4523 (N_4523,N_4383,N_4362);
nand U4524 (N_4524,N_4474,N_4331);
nor U4525 (N_4525,N_4353,N_4379);
and U4526 (N_4526,N_4430,N_4421);
nor U4527 (N_4527,N_4352,N_4446);
nand U4528 (N_4528,N_4371,N_4357);
xnor U4529 (N_4529,N_4429,N_4417);
or U4530 (N_4530,N_4455,N_4402);
or U4531 (N_4531,N_4332,N_4391);
and U4532 (N_4532,N_4328,N_4423);
nand U4533 (N_4533,N_4467,N_4456);
and U4534 (N_4534,N_4321,N_4451);
and U4535 (N_4535,N_4479,N_4461);
nand U4536 (N_4536,N_4392,N_4436);
xor U4537 (N_4537,N_4457,N_4387);
or U4538 (N_4538,N_4322,N_4343);
nor U4539 (N_4539,N_4400,N_4394);
xor U4540 (N_4540,N_4424,N_4433);
nor U4541 (N_4541,N_4473,N_4477);
nand U4542 (N_4542,N_4329,N_4342);
and U4543 (N_4543,N_4367,N_4418);
or U4544 (N_4544,N_4396,N_4393);
nand U4545 (N_4545,N_4344,N_4459);
xor U4546 (N_4546,N_4438,N_4432);
and U4547 (N_4547,N_4373,N_4395);
and U4548 (N_4548,N_4361,N_4419);
or U4549 (N_4549,N_4358,N_4403);
nor U4550 (N_4550,N_4339,N_4404);
or U4551 (N_4551,N_4468,N_4453);
nand U4552 (N_4552,N_4425,N_4445);
or U4553 (N_4553,N_4440,N_4452);
xnor U4554 (N_4554,N_4406,N_4350);
nor U4555 (N_4555,N_4330,N_4390);
and U4556 (N_4556,N_4366,N_4346);
or U4557 (N_4557,N_4369,N_4444);
or U4558 (N_4558,N_4341,N_4347);
nor U4559 (N_4559,N_4414,N_4380);
nor U4560 (N_4560,N_4385,N_4400);
and U4561 (N_4561,N_4447,N_4354);
nor U4562 (N_4562,N_4394,N_4458);
and U4563 (N_4563,N_4469,N_4387);
xnor U4564 (N_4564,N_4341,N_4436);
nor U4565 (N_4565,N_4404,N_4436);
nor U4566 (N_4566,N_4377,N_4455);
and U4567 (N_4567,N_4478,N_4407);
or U4568 (N_4568,N_4465,N_4415);
nor U4569 (N_4569,N_4378,N_4441);
nand U4570 (N_4570,N_4344,N_4405);
nor U4571 (N_4571,N_4371,N_4351);
xnor U4572 (N_4572,N_4328,N_4358);
xnor U4573 (N_4573,N_4419,N_4369);
nand U4574 (N_4574,N_4426,N_4335);
and U4575 (N_4575,N_4324,N_4323);
and U4576 (N_4576,N_4414,N_4321);
nand U4577 (N_4577,N_4375,N_4472);
nor U4578 (N_4578,N_4412,N_4321);
xor U4579 (N_4579,N_4330,N_4432);
and U4580 (N_4580,N_4438,N_4418);
nor U4581 (N_4581,N_4419,N_4427);
or U4582 (N_4582,N_4455,N_4324);
nor U4583 (N_4583,N_4393,N_4324);
and U4584 (N_4584,N_4432,N_4323);
or U4585 (N_4585,N_4353,N_4429);
or U4586 (N_4586,N_4423,N_4347);
xnor U4587 (N_4587,N_4351,N_4435);
or U4588 (N_4588,N_4436,N_4454);
xnor U4589 (N_4589,N_4476,N_4452);
xor U4590 (N_4590,N_4452,N_4470);
nor U4591 (N_4591,N_4426,N_4400);
or U4592 (N_4592,N_4391,N_4341);
or U4593 (N_4593,N_4440,N_4404);
and U4594 (N_4594,N_4439,N_4355);
nor U4595 (N_4595,N_4447,N_4445);
nand U4596 (N_4596,N_4356,N_4389);
xor U4597 (N_4597,N_4362,N_4331);
and U4598 (N_4598,N_4348,N_4326);
nand U4599 (N_4599,N_4380,N_4375);
or U4600 (N_4600,N_4444,N_4420);
and U4601 (N_4601,N_4350,N_4338);
and U4602 (N_4602,N_4417,N_4371);
and U4603 (N_4603,N_4416,N_4412);
or U4604 (N_4604,N_4418,N_4415);
or U4605 (N_4605,N_4412,N_4348);
or U4606 (N_4606,N_4376,N_4479);
xnor U4607 (N_4607,N_4418,N_4417);
nor U4608 (N_4608,N_4372,N_4357);
nand U4609 (N_4609,N_4359,N_4479);
nor U4610 (N_4610,N_4359,N_4477);
nor U4611 (N_4611,N_4431,N_4425);
or U4612 (N_4612,N_4397,N_4370);
nand U4613 (N_4613,N_4458,N_4372);
and U4614 (N_4614,N_4460,N_4435);
or U4615 (N_4615,N_4329,N_4391);
and U4616 (N_4616,N_4460,N_4364);
nand U4617 (N_4617,N_4361,N_4390);
xnor U4618 (N_4618,N_4325,N_4326);
nor U4619 (N_4619,N_4329,N_4332);
nor U4620 (N_4620,N_4425,N_4327);
nor U4621 (N_4621,N_4373,N_4448);
nor U4622 (N_4622,N_4327,N_4391);
or U4623 (N_4623,N_4320,N_4330);
nand U4624 (N_4624,N_4405,N_4361);
nor U4625 (N_4625,N_4428,N_4351);
xnor U4626 (N_4626,N_4369,N_4384);
or U4627 (N_4627,N_4372,N_4416);
or U4628 (N_4628,N_4350,N_4434);
and U4629 (N_4629,N_4392,N_4343);
or U4630 (N_4630,N_4439,N_4479);
nor U4631 (N_4631,N_4392,N_4417);
and U4632 (N_4632,N_4400,N_4459);
nor U4633 (N_4633,N_4345,N_4320);
and U4634 (N_4634,N_4406,N_4347);
or U4635 (N_4635,N_4342,N_4444);
xor U4636 (N_4636,N_4375,N_4438);
xor U4637 (N_4637,N_4461,N_4353);
nand U4638 (N_4638,N_4404,N_4424);
nor U4639 (N_4639,N_4411,N_4431);
nor U4640 (N_4640,N_4574,N_4624);
xor U4641 (N_4641,N_4544,N_4539);
and U4642 (N_4642,N_4553,N_4627);
xnor U4643 (N_4643,N_4616,N_4591);
nand U4644 (N_4644,N_4609,N_4514);
and U4645 (N_4645,N_4583,N_4491);
nand U4646 (N_4646,N_4637,N_4495);
nand U4647 (N_4647,N_4496,N_4596);
and U4648 (N_4648,N_4481,N_4606);
nand U4649 (N_4649,N_4480,N_4618);
xnor U4650 (N_4650,N_4497,N_4633);
nor U4651 (N_4651,N_4562,N_4504);
nand U4652 (N_4652,N_4538,N_4608);
or U4653 (N_4653,N_4517,N_4561);
nor U4654 (N_4654,N_4505,N_4498);
xor U4655 (N_4655,N_4623,N_4625);
xnor U4656 (N_4656,N_4488,N_4537);
or U4657 (N_4657,N_4522,N_4494);
xnor U4658 (N_4658,N_4567,N_4575);
and U4659 (N_4659,N_4592,N_4564);
and U4660 (N_4660,N_4510,N_4565);
and U4661 (N_4661,N_4534,N_4593);
and U4662 (N_4662,N_4587,N_4612);
xor U4663 (N_4663,N_4524,N_4526);
nor U4664 (N_4664,N_4557,N_4548);
xor U4665 (N_4665,N_4519,N_4585);
nand U4666 (N_4666,N_4607,N_4581);
or U4667 (N_4667,N_4571,N_4533);
or U4668 (N_4668,N_4611,N_4525);
and U4669 (N_4669,N_4630,N_4500);
nand U4670 (N_4670,N_4631,N_4604);
or U4671 (N_4671,N_4527,N_4584);
or U4672 (N_4672,N_4489,N_4594);
or U4673 (N_4673,N_4532,N_4547);
and U4674 (N_4674,N_4541,N_4638);
xor U4675 (N_4675,N_4508,N_4490);
xnor U4676 (N_4676,N_4560,N_4511);
nand U4677 (N_4677,N_4580,N_4601);
nor U4678 (N_4678,N_4509,N_4523);
nor U4679 (N_4679,N_4598,N_4577);
nand U4680 (N_4680,N_4566,N_4516);
nor U4681 (N_4681,N_4485,N_4569);
or U4682 (N_4682,N_4529,N_4515);
or U4683 (N_4683,N_4626,N_4503);
nand U4684 (N_4684,N_4563,N_4589);
nand U4685 (N_4685,N_4605,N_4595);
nand U4686 (N_4686,N_4540,N_4482);
and U4687 (N_4687,N_4555,N_4590);
and U4688 (N_4688,N_4542,N_4615);
nand U4689 (N_4689,N_4513,N_4639);
or U4690 (N_4690,N_4549,N_4582);
and U4691 (N_4691,N_4629,N_4603);
nor U4692 (N_4692,N_4502,N_4632);
or U4693 (N_4693,N_4622,N_4530);
nor U4694 (N_4694,N_4528,N_4493);
and U4695 (N_4695,N_4573,N_4492);
nand U4696 (N_4696,N_4578,N_4543);
and U4697 (N_4697,N_4634,N_4520);
or U4698 (N_4698,N_4613,N_4620);
xnor U4699 (N_4699,N_4599,N_4586);
nand U4700 (N_4700,N_4535,N_4487);
nand U4701 (N_4701,N_4621,N_4558);
and U4702 (N_4702,N_4536,N_4597);
nand U4703 (N_4703,N_4617,N_4518);
xnor U4704 (N_4704,N_4570,N_4546);
nor U4705 (N_4705,N_4619,N_4545);
or U4706 (N_4706,N_4579,N_4636);
and U4707 (N_4707,N_4484,N_4600);
or U4708 (N_4708,N_4628,N_4551);
nor U4709 (N_4709,N_4507,N_4572);
nand U4710 (N_4710,N_4614,N_4501);
and U4711 (N_4711,N_4554,N_4550);
nor U4712 (N_4712,N_4483,N_4610);
xnor U4713 (N_4713,N_4512,N_4506);
and U4714 (N_4714,N_4556,N_4568);
or U4715 (N_4715,N_4588,N_4531);
or U4716 (N_4716,N_4559,N_4602);
nand U4717 (N_4717,N_4521,N_4576);
and U4718 (N_4718,N_4635,N_4499);
xor U4719 (N_4719,N_4552,N_4486);
nand U4720 (N_4720,N_4639,N_4494);
or U4721 (N_4721,N_4563,N_4610);
nand U4722 (N_4722,N_4574,N_4612);
and U4723 (N_4723,N_4523,N_4504);
and U4724 (N_4724,N_4627,N_4545);
and U4725 (N_4725,N_4523,N_4590);
nor U4726 (N_4726,N_4503,N_4525);
nor U4727 (N_4727,N_4616,N_4560);
nor U4728 (N_4728,N_4565,N_4548);
and U4729 (N_4729,N_4556,N_4559);
nor U4730 (N_4730,N_4545,N_4612);
and U4731 (N_4731,N_4552,N_4612);
and U4732 (N_4732,N_4590,N_4588);
nand U4733 (N_4733,N_4501,N_4618);
and U4734 (N_4734,N_4627,N_4508);
xnor U4735 (N_4735,N_4636,N_4535);
nand U4736 (N_4736,N_4575,N_4597);
nand U4737 (N_4737,N_4569,N_4638);
or U4738 (N_4738,N_4488,N_4520);
or U4739 (N_4739,N_4536,N_4574);
or U4740 (N_4740,N_4496,N_4587);
xnor U4741 (N_4741,N_4487,N_4493);
or U4742 (N_4742,N_4497,N_4540);
nand U4743 (N_4743,N_4492,N_4565);
nor U4744 (N_4744,N_4515,N_4599);
nor U4745 (N_4745,N_4527,N_4568);
xnor U4746 (N_4746,N_4555,N_4520);
nand U4747 (N_4747,N_4521,N_4622);
or U4748 (N_4748,N_4628,N_4600);
or U4749 (N_4749,N_4542,N_4517);
and U4750 (N_4750,N_4626,N_4489);
or U4751 (N_4751,N_4590,N_4535);
nor U4752 (N_4752,N_4612,N_4601);
nor U4753 (N_4753,N_4537,N_4532);
and U4754 (N_4754,N_4540,N_4623);
nand U4755 (N_4755,N_4605,N_4496);
nand U4756 (N_4756,N_4630,N_4489);
nor U4757 (N_4757,N_4622,N_4528);
nor U4758 (N_4758,N_4635,N_4589);
and U4759 (N_4759,N_4551,N_4496);
nor U4760 (N_4760,N_4593,N_4620);
nor U4761 (N_4761,N_4540,N_4534);
xnor U4762 (N_4762,N_4539,N_4571);
nand U4763 (N_4763,N_4632,N_4626);
or U4764 (N_4764,N_4552,N_4581);
and U4765 (N_4765,N_4509,N_4616);
and U4766 (N_4766,N_4527,N_4529);
nor U4767 (N_4767,N_4578,N_4587);
nor U4768 (N_4768,N_4619,N_4567);
or U4769 (N_4769,N_4526,N_4493);
or U4770 (N_4770,N_4563,N_4597);
nand U4771 (N_4771,N_4539,N_4585);
nor U4772 (N_4772,N_4555,N_4534);
nand U4773 (N_4773,N_4480,N_4505);
or U4774 (N_4774,N_4549,N_4548);
xor U4775 (N_4775,N_4577,N_4516);
xnor U4776 (N_4776,N_4587,N_4530);
and U4777 (N_4777,N_4538,N_4504);
or U4778 (N_4778,N_4621,N_4608);
or U4779 (N_4779,N_4569,N_4550);
or U4780 (N_4780,N_4581,N_4512);
and U4781 (N_4781,N_4490,N_4627);
xnor U4782 (N_4782,N_4638,N_4587);
nor U4783 (N_4783,N_4520,N_4489);
nor U4784 (N_4784,N_4627,N_4581);
nor U4785 (N_4785,N_4602,N_4541);
nand U4786 (N_4786,N_4563,N_4609);
nand U4787 (N_4787,N_4569,N_4614);
xnor U4788 (N_4788,N_4528,N_4526);
nand U4789 (N_4789,N_4527,N_4507);
xor U4790 (N_4790,N_4528,N_4564);
nor U4791 (N_4791,N_4624,N_4524);
xnor U4792 (N_4792,N_4600,N_4505);
nor U4793 (N_4793,N_4506,N_4523);
or U4794 (N_4794,N_4530,N_4494);
xnor U4795 (N_4795,N_4605,N_4532);
and U4796 (N_4796,N_4605,N_4531);
nand U4797 (N_4797,N_4539,N_4490);
xor U4798 (N_4798,N_4635,N_4487);
nor U4799 (N_4799,N_4632,N_4581);
nand U4800 (N_4800,N_4672,N_4669);
nand U4801 (N_4801,N_4795,N_4719);
nand U4802 (N_4802,N_4732,N_4665);
or U4803 (N_4803,N_4670,N_4733);
and U4804 (N_4804,N_4717,N_4794);
nor U4805 (N_4805,N_4780,N_4762);
nor U4806 (N_4806,N_4664,N_4648);
nor U4807 (N_4807,N_4770,N_4680);
nor U4808 (N_4808,N_4775,N_4647);
nand U4809 (N_4809,N_4673,N_4763);
or U4810 (N_4810,N_4728,N_4695);
nand U4811 (N_4811,N_4760,N_4707);
nor U4812 (N_4812,N_4713,N_4744);
nor U4813 (N_4813,N_4653,N_4658);
xor U4814 (N_4814,N_4736,N_4730);
nor U4815 (N_4815,N_4696,N_4750);
or U4816 (N_4816,N_4722,N_4700);
and U4817 (N_4817,N_4789,N_4694);
nand U4818 (N_4818,N_4640,N_4787);
nor U4819 (N_4819,N_4771,N_4688);
xor U4820 (N_4820,N_4738,N_4715);
nor U4821 (N_4821,N_4666,N_4793);
and U4822 (N_4822,N_4788,N_4721);
nor U4823 (N_4823,N_4687,N_4755);
and U4824 (N_4824,N_4756,N_4652);
xor U4825 (N_4825,N_4706,N_4781);
nand U4826 (N_4826,N_4646,N_4727);
and U4827 (N_4827,N_4735,N_4685);
nand U4828 (N_4828,N_4747,N_4778);
and U4829 (N_4829,N_4720,N_4659);
or U4830 (N_4830,N_4708,N_4724);
or U4831 (N_4831,N_4798,N_4797);
nor U4832 (N_4832,N_4681,N_4705);
and U4833 (N_4833,N_4774,N_4679);
nand U4834 (N_4834,N_4644,N_4667);
nor U4835 (N_4835,N_4662,N_4741);
xnor U4836 (N_4836,N_4668,N_4690);
or U4837 (N_4837,N_4758,N_4686);
or U4838 (N_4838,N_4785,N_4742);
or U4839 (N_4839,N_4754,N_4691);
nand U4840 (N_4840,N_4676,N_4649);
xnor U4841 (N_4841,N_4702,N_4726);
xor U4842 (N_4842,N_4779,N_4718);
nor U4843 (N_4843,N_4678,N_4783);
nand U4844 (N_4844,N_4660,N_4697);
and U4845 (N_4845,N_4782,N_4693);
or U4846 (N_4846,N_4739,N_4745);
nand U4847 (N_4847,N_4651,N_4743);
or U4848 (N_4848,N_4799,N_4757);
nor U4849 (N_4849,N_4777,N_4753);
and U4850 (N_4850,N_4684,N_4711);
xnor U4851 (N_4851,N_4645,N_4714);
xor U4852 (N_4852,N_4784,N_4716);
nand U4853 (N_4853,N_4703,N_4769);
nand U4854 (N_4854,N_4766,N_4731);
xor U4855 (N_4855,N_4663,N_4790);
or U4856 (N_4856,N_4796,N_4764);
or U4857 (N_4857,N_4704,N_4725);
xor U4858 (N_4858,N_4675,N_4768);
nand U4859 (N_4859,N_4692,N_4759);
nand U4860 (N_4860,N_4761,N_4773);
nand U4861 (N_4861,N_4650,N_4748);
nor U4862 (N_4862,N_4674,N_4752);
xnor U4863 (N_4863,N_4656,N_4710);
or U4864 (N_4864,N_4740,N_4657);
or U4865 (N_4865,N_4661,N_4671);
and U4866 (N_4866,N_4682,N_4729);
or U4867 (N_4867,N_4776,N_4791);
or U4868 (N_4868,N_4723,N_4642);
and U4869 (N_4869,N_4677,N_4654);
or U4870 (N_4870,N_4786,N_4641);
nor U4871 (N_4871,N_4712,N_4767);
nand U4872 (N_4872,N_4643,N_4683);
nor U4873 (N_4873,N_4749,N_4709);
and U4874 (N_4874,N_4734,N_4655);
nand U4875 (N_4875,N_4701,N_4765);
nand U4876 (N_4876,N_4746,N_4772);
and U4877 (N_4877,N_4698,N_4699);
nand U4878 (N_4878,N_4792,N_4751);
xnor U4879 (N_4879,N_4689,N_4737);
nor U4880 (N_4880,N_4665,N_4792);
xnor U4881 (N_4881,N_4655,N_4776);
nand U4882 (N_4882,N_4733,N_4644);
and U4883 (N_4883,N_4737,N_4653);
nor U4884 (N_4884,N_4656,N_4698);
and U4885 (N_4885,N_4749,N_4779);
nor U4886 (N_4886,N_4681,N_4679);
and U4887 (N_4887,N_4743,N_4753);
nand U4888 (N_4888,N_4643,N_4738);
nand U4889 (N_4889,N_4749,N_4662);
xnor U4890 (N_4890,N_4640,N_4669);
nand U4891 (N_4891,N_4728,N_4792);
xor U4892 (N_4892,N_4665,N_4721);
nor U4893 (N_4893,N_4750,N_4764);
nand U4894 (N_4894,N_4654,N_4730);
nor U4895 (N_4895,N_4731,N_4774);
or U4896 (N_4896,N_4747,N_4677);
xor U4897 (N_4897,N_4647,N_4753);
and U4898 (N_4898,N_4678,N_4706);
nand U4899 (N_4899,N_4658,N_4674);
nor U4900 (N_4900,N_4695,N_4666);
and U4901 (N_4901,N_4775,N_4674);
nand U4902 (N_4902,N_4764,N_4690);
or U4903 (N_4903,N_4682,N_4678);
and U4904 (N_4904,N_4684,N_4663);
and U4905 (N_4905,N_4723,N_4664);
or U4906 (N_4906,N_4730,N_4746);
nor U4907 (N_4907,N_4768,N_4659);
and U4908 (N_4908,N_4653,N_4664);
xor U4909 (N_4909,N_4663,N_4797);
xor U4910 (N_4910,N_4783,N_4648);
and U4911 (N_4911,N_4658,N_4744);
xor U4912 (N_4912,N_4684,N_4666);
or U4913 (N_4913,N_4713,N_4699);
nor U4914 (N_4914,N_4642,N_4742);
xnor U4915 (N_4915,N_4646,N_4686);
and U4916 (N_4916,N_4679,N_4695);
nor U4917 (N_4917,N_4796,N_4698);
xnor U4918 (N_4918,N_4728,N_4749);
and U4919 (N_4919,N_4692,N_4683);
or U4920 (N_4920,N_4714,N_4652);
and U4921 (N_4921,N_4668,N_4684);
nand U4922 (N_4922,N_4706,N_4766);
xor U4923 (N_4923,N_4664,N_4660);
nand U4924 (N_4924,N_4735,N_4719);
nor U4925 (N_4925,N_4663,N_4719);
and U4926 (N_4926,N_4650,N_4672);
nand U4927 (N_4927,N_4690,N_4797);
or U4928 (N_4928,N_4667,N_4697);
and U4929 (N_4929,N_4751,N_4659);
and U4930 (N_4930,N_4709,N_4688);
or U4931 (N_4931,N_4707,N_4770);
xnor U4932 (N_4932,N_4760,N_4783);
or U4933 (N_4933,N_4758,N_4767);
nor U4934 (N_4934,N_4702,N_4660);
and U4935 (N_4935,N_4731,N_4683);
nand U4936 (N_4936,N_4769,N_4677);
xor U4937 (N_4937,N_4779,N_4740);
nand U4938 (N_4938,N_4742,N_4740);
nor U4939 (N_4939,N_4734,N_4644);
and U4940 (N_4940,N_4760,N_4713);
and U4941 (N_4941,N_4662,N_4735);
or U4942 (N_4942,N_4746,N_4703);
and U4943 (N_4943,N_4732,N_4782);
xor U4944 (N_4944,N_4742,N_4688);
or U4945 (N_4945,N_4753,N_4658);
or U4946 (N_4946,N_4726,N_4747);
xnor U4947 (N_4947,N_4647,N_4783);
nand U4948 (N_4948,N_4781,N_4767);
and U4949 (N_4949,N_4784,N_4724);
nand U4950 (N_4950,N_4671,N_4714);
and U4951 (N_4951,N_4680,N_4722);
or U4952 (N_4952,N_4700,N_4796);
and U4953 (N_4953,N_4684,N_4699);
and U4954 (N_4954,N_4644,N_4669);
nor U4955 (N_4955,N_4744,N_4779);
and U4956 (N_4956,N_4760,N_4644);
xnor U4957 (N_4957,N_4648,N_4731);
xnor U4958 (N_4958,N_4757,N_4712);
xnor U4959 (N_4959,N_4654,N_4727);
nand U4960 (N_4960,N_4956,N_4933);
nand U4961 (N_4961,N_4928,N_4898);
or U4962 (N_4962,N_4953,N_4895);
or U4963 (N_4963,N_4856,N_4812);
nand U4964 (N_4964,N_4888,N_4950);
nand U4965 (N_4965,N_4916,N_4848);
nand U4966 (N_4966,N_4818,N_4836);
nor U4967 (N_4967,N_4958,N_4806);
nand U4968 (N_4968,N_4879,N_4834);
xnor U4969 (N_4969,N_4919,N_4827);
and U4970 (N_4970,N_4954,N_4922);
xor U4971 (N_4971,N_4857,N_4808);
or U4972 (N_4972,N_4837,N_4927);
or U4973 (N_4973,N_4894,N_4905);
nor U4974 (N_4974,N_4903,N_4820);
and U4975 (N_4975,N_4801,N_4811);
or U4976 (N_4976,N_4893,N_4830);
xnor U4977 (N_4977,N_4946,N_4809);
and U4978 (N_4978,N_4939,N_4829);
and U4979 (N_4979,N_4911,N_4876);
xor U4980 (N_4980,N_4815,N_4951);
nand U4981 (N_4981,N_4874,N_4904);
xnor U4982 (N_4982,N_4864,N_4841);
xor U4983 (N_4983,N_4936,N_4934);
or U4984 (N_4984,N_4886,N_4900);
xnor U4985 (N_4985,N_4839,N_4855);
nand U4986 (N_4986,N_4920,N_4889);
xnor U4987 (N_4987,N_4882,N_4924);
and U4988 (N_4988,N_4925,N_4878);
xnor U4989 (N_4989,N_4802,N_4943);
nand U4990 (N_4990,N_4947,N_4826);
nor U4991 (N_4991,N_4892,N_4932);
or U4992 (N_4992,N_4938,N_4907);
nand U4993 (N_4993,N_4838,N_4948);
nor U4994 (N_4994,N_4854,N_4923);
nand U4995 (N_4995,N_4828,N_4944);
or U4996 (N_4996,N_4942,N_4896);
or U4997 (N_4997,N_4816,N_4917);
and U4998 (N_4998,N_4859,N_4813);
xor U4999 (N_4999,N_4887,N_4871);
or U5000 (N_5000,N_4868,N_4843);
nand U5001 (N_5001,N_4910,N_4912);
nand U5002 (N_5002,N_4861,N_4897);
nor U5003 (N_5003,N_4862,N_4952);
xnor U5004 (N_5004,N_4810,N_4865);
or U5005 (N_5005,N_4853,N_4822);
xor U5006 (N_5006,N_4842,N_4908);
and U5007 (N_5007,N_4959,N_4872);
nor U5008 (N_5008,N_4825,N_4881);
or U5009 (N_5009,N_4850,N_4805);
nor U5010 (N_5010,N_4835,N_4866);
nand U5011 (N_5011,N_4885,N_4847);
nor U5012 (N_5012,N_4913,N_4931);
or U5013 (N_5013,N_4884,N_4914);
nor U5014 (N_5014,N_4849,N_4831);
and U5015 (N_5015,N_4800,N_4940);
nand U5016 (N_5016,N_4930,N_4863);
xor U5017 (N_5017,N_4844,N_4858);
nor U5018 (N_5018,N_4840,N_4867);
and U5019 (N_5019,N_4918,N_4891);
and U5020 (N_5020,N_4949,N_4902);
nor U5021 (N_5021,N_4929,N_4890);
or U5022 (N_5022,N_4869,N_4852);
nor U5023 (N_5023,N_4957,N_4926);
or U5024 (N_5024,N_4873,N_4883);
and U5025 (N_5025,N_4901,N_4845);
nor U5026 (N_5026,N_4814,N_4833);
and U5027 (N_5027,N_4821,N_4846);
xnor U5028 (N_5028,N_4899,N_4906);
or U5029 (N_5029,N_4935,N_4945);
nand U5030 (N_5030,N_4877,N_4823);
nand U5031 (N_5031,N_4832,N_4851);
xor U5032 (N_5032,N_4819,N_4807);
nor U5033 (N_5033,N_4915,N_4803);
nand U5034 (N_5034,N_4941,N_4955);
and U5035 (N_5035,N_4804,N_4921);
and U5036 (N_5036,N_4817,N_4860);
nor U5037 (N_5037,N_4870,N_4875);
nand U5038 (N_5038,N_4937,N_4880);
nand U5039 (N_5039,N_4824,N_4909);
nor U5040 (N_5040,N_4856,N_4811);
xor U5041 (N_5041,N_4805,N_4854);
or U5042 (N_5042,N_4909,N_4863);
xnor U5043 (N_5043,N_4834,N_4824);
nor U5044 (N_5044,N_4893,N_4934);
xor U5045 (N_5045,N_4881,N_4828);
or U5046 (N_5046,N_4902,N_4814);
or U5047 (N_5047,N_4862,N_4815);
nor U5048 (N_5048,N_4838,N_4891);
nor U5049 (N_5049,N_4897,N_4931);
nand U5050 (N_5050,N_4857,N_4836);
or U5051 (N_5051,N_4877,N_4889);
or U5052 (N_5052,N_4826,N_4945);
xor U5053 (N_5053,N_4903,N_4848);
and U5054 (N_5054,N_4901,N_4931);
or U5055 (N_5055,N_4827,N_4875);
or U5056 (N_5056,N_4899,N_4880);
xor U5057 (N_5057,N_4848,N_4908);
xnor U5058 (N_5058,N_4861,N_4914);
and U5059 (N_5059,N_4940,N_4888);
xnor U5060 (N_5060,N_4825,N_4898);
xnor U5061 (N_5061,N_4845,N_4944);
or U5062 (N_5062,N_4812,N_4858);
or U5063 (N_5063,N_4855,N_4826);
xnor U5064 (N_5064,N_4888,N_4907);
nand U5065 (N_5065,N_4907,N_4910);
xnor U5066 (N_5066,N_4849,N_4824);
nand U5067 (N_5067,N_4924,N_4875);
xnor U5068 (N_5068,N_4947,N_4843);
nor U5069 (N_5069,N_4956,N_4940);
nand U5070 (N_5070,N_4913,N_4946);
nand U5071 (N_5071,N_4901,N_4951);
nand U5072 (N_5072,N_4916,N_4868);
nor U5073 (N_5073,N_4830,N_4806);
nand U5074 (N_5074,N_4843,N_4870);
nand U5075 (N_5075,N_4949,N_4845);
and U5076 (N_5076,N_4942,N_4927);
and U5077 (N_5077,N_4903,N_4827);
nor U5078 (N_5078,N_4959,N_4828);
xnor U5079 (N_5079,N_4909,N_4951);
or U5080 (N_5080,N_4802,N_4836);
or U5081 (N_5081,N_4901,N_4869);
nand U5082 (N_5082,N_4950,N_4846);
nand U5083 (N_5083,N_4865,N_4883);
and U5084 (N_5084,N_4872,N_4925);
and U5085 (N_5085,N_4902,N_4884);
or U5086 (N_5086,N_4807,N_4862);
and U5087 (N_5087,N_4928,N_4956);
and U5088 (N_5088,N_4818,N_4864);
nand U5089 (N_5089,N_4829,N_4888);
nor U5090 (N_5090,N_4874,N_4954);
or U5091 (N_5091,N_4944,N_4936);
and U5092 (N_5092,N_4891,N_4903);
or U5093 (N_5093,N_4911,N_4860);
or U5094 (N_5094,N_4866,N_4892);
xor U5095 (N_5095,N_4909,N_4954);
nand U5096 (N_5096,N_4926,N_4820);
or U5097 (N_5097,N_4860,N_4825);
or U5098 (N_5098,N_4829,N_4818);
and U5099 (N_5099,N_4817,N_4898);
or U5100 (N_5100,N_4806,N_4866);
nand U5101 (N_5101,N_4833,N_4889);
nand U5102 (N_5102,N_4840,N_4885);
xor U5103 (N_5103,N_4904,N_4905);
nor U5104 (N_5104,N_4817,N_4801);
and U5105 (N_5105,N_4803,N_4958);
or U5106 (N_5106,N_4874,N_4898);
and U5107 (N_5107,N_4945,N_4940);
or U5108 (N_5108,N_4816,N_4827);
xnor U5109 (N_5109,N_4894,N_4878);
and U5110 (N_5110,N_4846,N_4882);
xor U5111 (N_5111,N_4804,N_4912);
and U5112 (N_5112,N_4930,N_4949);
xnor U5113 (N_5113,N_4902,N_4878);
xnor U5114 (N_5114,N_4832,N_4909);
nand U5115 (N_5115,N_4863,N_4894);
and U5116 (N_5116,N_4886,N_4932);
nand U5117 (N_5117,N_4901,N_4922);
nor U5118 (N_5118,N_4933,N_4851);
or U5119 (N_5119,N_4930,N_4864);
nor U5120 (N_5120,N_4986,N_4981);
and U5121 (N_5121,N_5014,N_5045);
nand U5122 (N_5122,N_5052,N_5012);
and U5123 (N_5123,N_4970,N_5081);
or U5124 (N_5124,N_5009,N_4991);
or U5125 (N_5125,N_5032,N_4979);
xnor U5126 (N_5126,N_5007,N_4987);
and U5127 (N_5127,N_5102,N_4976);
nand U5128 (N_5128,N_4967,N_5040);
or U5129 (N_5129,N_5088,N_5118);
nor U5130 (N_5130,N_5079,N_5098);
and U5131 (N_5131,N_5071,N_5092);
xnor U5132 (N_5132,N_5113,N_5075);
or U5133 (N_5133,N_5025,N_5089);
xnor U5134 (N_5134,N_5006,N_5105);
nand U5135 (N_5135,N_5049,N_5110);
nor U5136 (N_5136,N_5059,N_5116);
and U5137 (N_5137,N_5020,N_5039);
or U5138 (N_5138,N_4973,N_5076);
xnor U5139 (N_5139,N_5077,N_5107);
nand U5140 (N_5140,N_4995,N_4980);
nor U5141 (N_5141,N_4997,N_5108);
nor U5142 (N_5142,N_5047,N_5060);
or U5143 (N_5143,N_5094,N_4984);
nand U5144 (N_5144,N_5058,N_4977);
and U5145 (N_5145,N_5067,N_5037);
nor U5146 (N_5146,N_5061,N_4993);
xnor U5147 (N_5147,N_4962,N_5099);
or U5148 (N_5148,N_5003,N_5042);
nor U5149 (N_5149,N_5074,N_5086);
or U5150 (N_5150,N_5008,N_5066);
and U5151 (N_5151,N_4965,N_5093);
or U5152 (N_5152,N_5084,N_4971);
xor U5153 (N_5153,N_5034,N_4983);
xor U5154 (N_5154,N_5057,N_4964);
xor U5155 (N_5155,N_5016,N_5023);
or U5156 (N_5156,N_5078,N_5019);
nor U5157 (N_5157,N_5096,N_5097);
and U5158 (N_5158,N_4996,N_5087);
nand U5159 (N_5159,N_4990,N_4999);
and U5160 (N_5160,N_5080,N_5054);
xnor U5161 (N_5161,N_5046,N_4988);
xnor U5162 (N_5162,N_5005,N_5112);
or U5163 (N_5163,N_5106,N_5064);
nand U5164 (N_5164,N_5073,N_5033);
xnor U5165 (N_5165,N_5043,N_5051);
xor U5166 (N_5166,N_5070,N_5055);
nor U5167 (N_5167,N_4992,N_4985);
nand U5168 (N_5168,N_5085,N_5044);
or U5169 (N_5169,N_5117,N_5029);
xnor U5170 (N_5170,N_4978,N_5103);
xor U5171 (N_5171,N_5017,N_5013);
or U5172 (N_5172,N_4982,N_4972);
and U5173 (N_5173,N_5010,N_5082);
and U5174 (N_5174,N_5000,N_5022);
nor U5175 (N_5175,N_5030,N_5015);
nand U5176 (N_5176,N_4975,N_5111);
nand U5177 (N_5177,N_5095,N_4989);
or U5178 (N_5178,N_5072,N_5114);
nand U5179 (N_5179,N_5004,N_5050);
or U5180 (N_5180,N_4994,N_4963);
nor U5181 (N_5181,N_4960,N_5083);
and U5182 (N_5182,N_5002,N_5100);
xnor U5183 (N_5183,N_5063,N_5035);
nor U5184 (N_5184,N_5065,N_4961);
xor U5185 (N_5185,N_5031,N_5011);
xnor U5186 (N_5186,N_5056,N_5090);
nand U5187 (N_5187,N_4974,N_5069);
or U5188 (N_5188,N_5091,N_4968);
and U5189 (N_5189,N_5018,N_5024);
and U5190 (N_5190,N_5036,N_5021);
nand U5191 (N_5191,N_5062,N_5053);
nor U5192 (N_5192,N_5038,N_5109);
xnor U5193 (N_5193,N_5028,N_5041);
xnor U5194 (N_5194,N_5027,N_5001);
and U5195 (N_5195,N_5104,N_5068);
xor U5196 (N_5196,N_5115,N_4998);
nor U5197 (N_5197,N_5119,N_5048);
or U5198 (N_5198,N_5026,N_4969);
and U5199 (N_5199,N_5101,N_4966);
xnor U5200 (N_5200,N_5107,N_4961);
nor U5201 (N_5201,N_5015,N_5038);
or U5202 (N_5202,N_5077,N_5112);
xor U5203 (N_5203,N_5108,N_5030);
or U5204 (N_5204,N_5080,N_5075);
nand U5205 (N_5205,N_4961,N_4999);
and U5206 (N_5206,N_5029,N_5075);
nor U5207 (N_5207,N_5036,N_5078);
and U5208 (N_5208,N_4962,N_5077);
nor U5209 (N_5209,N_5010,N_5036);
or U5210 (N_5210,N_4985,N_5001);
nand U5211 (N_5211,N_4965,N_5025);
and U5212 (N_5212,N_5052,N_5063);
or U5213 (N_5213,N_5081,N_5004);
and U5214 (N_5214,N_5022,N_4998);
or U5215 (N_5215,N_5033,N_4962);
or U5216 (N_5216,N_5114,N_5078);
and U5217 (N_5217,N_5119,N_4981);
nand U5218 (N_5218,N_5097,N_4985);
nand U5219 (N_5219,N_5089,N_5038);
nand U5220 (N_5220,N_5008,N_5018);
and U5221 (N_5221,N_5038,N_5113);
xor U5222 (N_5222,N_4977,N_5082);
xnor U5223 (N_5223,N_5090,N_5083);
nor U5224 (N_5224,N_5021,N_5025);
nor U5225 (N_5225,N_5044,N_5103);
xor U5226 (N_5226,N_5101,N_5039);
xor U5227 (N_5227,N_4982,N_4994);
nand U5228 (N_5228,N_5095,N_5110);
and U5229 (N_5229,N_5041,N_5106);
and U5230 (N_5230,N_4992,N_5002);
and U5231 (N_5231,N_5078,N_5056);
and U5232 (N_5232,N_5100,N_5093);
nor U5233 (N_5233,N_5097,N_5041);
nand U5234 (N_5234,N_5015,N_5073);
xnor U5235 (N_5235,N_5032,N_5029);
nor U5236 (N_5236,N_5108,N_5037);
nor U5237 (N_5237,N_4973,N_4985);
xor U5238 (N_5238,N_5028,N_5033);
or U5239 (N_5239,N_5086,N_5060);
xor U5240 (N_5240,N_5083,N_4981);
and U5241 (N_5241,N_4969,N_5059);
xor U5242 (N_5242,N_4998,N_5025);
xor U5243 (N_5243,N_5039,N_5000);
xnor U5244 (N_5244,N_5025,N_5115);
nor U5245 (N_5245,N_5069,N_5023);
nand U5246 (N_5246,N_4996,N_5115);
or U5247 (N_5247,N_5063,N_5025);
nand U5248 (N_5248,N_5035,N_4962);
or U5249 (N_5249,N_4991,N_4999);
nand U5250 (N_5250,N_4963,N_4993);
and U5251 (N_5251,N_4985,N_4963);
nand U5252 (N_5252,N_5112,N_5035);
nor U5253 (N_5253,N_4984,N_5091);
nand U5254 (N_5254,N_5111,N_5117);
or U5255 (N_5255,N_5104,N_5090);
nor U5256 (N_5256,N_5045,N_4996);
and U5257 (N_5257,N_5085,N_5015);
and U5258 (N_5258,N_5034,N_5084);
or U5259 (N_5259,N_5111,N_5073);
nor U5260 (N_5260,N_5029,N_4988);
xor U5261 (N_5261,N_4961,N_5014);
or U5262 (N_5262,N_5037,N_5023);
nand U5263 (N_5263,N_4978,N_4973);
and U5264 (N_5264,N_4975,N_5080);
and U5265 (N_5265,N_5009,N_5027);
or U5266 (N_5266,N_5072,N_5083);
or U5267 (N_5267,N_5037,N_5081);
nor U5268 (N_5268,N_5011,N_5118);
nand U5269 (N_5269,N_5083,N_5064);
xor U5270 (N_5270,N_5099,N_4991);
nor U5271 (N_5271,N_5008,N_4997);
and U5272 (N_5272,N_5113,N_5116);
xnor U5273 (N_5273,N_5095,N_5106);
xnor U5274 (N_5274,N_5064,N_5057);
nor U5275 (N_5275,N_5100,N_5019);
or U5276 (N_5276,N_5067,N_5082);
nand U5277 (N_5277,N_5109,N_5015);
nand U5278 (N_5278,N_5086,N_4979);
nor U5279 (N_5279,N_5107,N_5029);
or U5280 (N_5280,N_5133,N_5261);
and U5281 (N_5281,N_5249,N_5274);
or U5282 (N_5282,N_5253,N_5273);
xnor U5283 (N_5283,N_5178,N_5163);
and U5284 (N_5284,N_5208,N_5227);
or U5285 (N_5285,N_5159,N_5199);
or U5286 (N_5286,N_5238,N_5168);
xnor U5287 (N_5287,N_5157,N_5129);
xnor U5288 (N_5288,N_5132,N_5179);
nor U5289 (N_5289,N_5175,N_5141);
nand U5290 (N_5290,N_5189,N_5184);
or U5291 (N_5291,N_5166,N_5143);
xnor U5292 (N_5292,N_5228,N_5135);
nor U5293 (N_5293,N_5236,N_5272);
nor U5294 (N_5294,N_5266,N_5194);
nand U5295 (N_5295,N_5220,N_5186);
and U5296 (N_5296,N_5267,N_5125);
or U5297 (N_5297,N_5201,N_5202);
xor U5298 (N_5298,N_5138,N_5187);
nor U5299 (N_5299,N_5185,N_5149);
nor U5300 (N_5300,N_5121,N_5269);
nor U5301 (N_5301,N_5239,N_5247);
and U5302 (N_5302,N_5232,N_5152);
nor U5303 (N_5303,N_5260,N_5172);
or U5304 (N_5304,N_5203,N_5154);
or U5305 (N_5305,N_5130,N_5271);
and U5306 (N_5306,N_5222,N_5206);
or U5307 (N_5307,N_5136,N_5131);
nand U5308 (N_5308,N_5278,N_5140);
xnor U5309 (N_5309,N_5263,N_5195);
nand U5310 (N_5310,N_5259,N_5254);
nor U5311 (N_5311,N_5174,N_5171);
and U5312 (N_5312,N_5204,N_5262);
nand U5313 (N_5313,N_5250,N_5170);
and U5314 (N_5314,N_5167,N_5226);
or U5315 (N_5315,N_5265,N_5241);
xor U5316 (N_5316,N_5235,N_5277);
nor U5317 (N_5317,N_5120,N_5122);
nand U5318 (N_5318,N_5158,N_5214);
nand U5319 (N_5319,N_5237,N_5252);
and U5320 (N_5320,N_5193,N_5180);
or U5321 (N_5321,N_5190,N_5123);
or U5322 (N_5322,N_5146,N_5234);
or U5323 (N_5323,N_5188,N_5233);
or U5324 (N_5324,N_5270,N_5139);
or U5325 (N_5325,N_5245,N_5244);
nor U5326 (N_5326,N_5279,N_5137);
nand U5327 (N_5327,N_5210,N_5224);
nor U5328 (N_5328,N_5275,N_5225);
or U5329 (N_5329,N_5197,N_5191);
and U5330 (N_5330,N_5276,N_5221);
nor U5331 (N_5331,N_5258,N_5150);
nor U5332 (N_5332,N_5264,N_5134);
xnor U5333 (N_5333,N_5155,N_5181);
xor U5334 (N_5334,N_5161,N_5217);
nand U5335 (N_5335,N_5211,N_5126);
nand U5336 (N_5336,N_5165,N_5229);
nand U5337 (N_5337,N_5248,N_5246);
nand U5338 (N_5338,N_5145,N_5242);
and U5339 (N_5339,N_5192,N_5124);
or U5340 (N_5340,N_5212,N_5151);
nor U5341 (N_5341,N_5148,N_5196);
and U5342 (N_5342,N_5142,N_5160);
nor U5343 (N_5343,N_5177,N_5164);
and U5344 (N_5344,N_5223,N_5240);
or U5345 (N_5345,N_5216,N_5207);
nor U5346 (N_5346,N_5257,N_5169);
or U5347 (N_5347,N_5209,N_5183);
xnor U5348 (N_5348,N_5176,N_5162);
or U5349 (N_5349,N_5215,N_5231);
and U5350 (N_5350,N_5147,N_5230);
nor U5351 (N_5351,N_5156,N_5182);
nor U5352 (N_5352,N_5200,N_5127);
nand U5353 (N_5353,N_5213,N_5268);
or U5354 (N_5354,N_5198,N_5255);
xnor U5355 (N_5355,N_5173,N_5128);
nor U5356 (N_5356,N_5144,N_5243);
nor U5357 (N_5357,N_5256,N_5153);
nand U5358 (N_5358,N_5251,N_5218);
xnor U5359 (N_5359,N_5205,N_5219);
nor U5360 (N_5360,N_5215,N_5251);
or U5361 (N_5361,N_5188,N_5179);
nor U5362 (N_5362,N_5176,N_5229);
nor U5363 (N_5363,N_5179,N_5229);
and U5364 (N_5364,N_5221,N_5202);
and U5365 (N_5365,N_5242,N_5266);
or U5366 (N_5366,N_5202,N_5235);
or U5367 (N_5367,N_5171,N_5250);
nor U5368 (N_5368,N_5128,N_5154);
xnor U5369 (N_5369,N_5234,N_5143);
nor U5370 (N_5370,N_5180,N_5128);
nand U5371 (N_5371,N_5194,N_5212);
nand U5372 (N_5372,N_5153,N_5274);
or U5373 (N_5373,N_5168,N_5212);
and U5374 (N_5374,N_5253,N_5156);
nand U5375 (N_5375,N_5247,N_5127);
nand U5376 (N_5376,N_5194,N_5141);
or U5377 (N_5377,N_5260,N_5127);
and U5378 (N_5378,N_5279,N_5230);
or U5379 (N_5379,N_5251,N_5201);
or U5380 (N_5380,N_5215,N_5154);
and U5381 (N_5381,N_5134,N_5235);
nor U5382 (N_5382,N_5196,N_5275);
and U5383 (N_5383,N_5202,N_5229);
or U5384 (N_5384,N_5160,N_5203);
nor U5385 (N_5385,N_5141,N_5149);
xor U5386 (N_5386,N_5148,N_5258);
or U5387 (N_5387,N_5172,N_5174);
xnor U5388 (N_5388,N_5193,N_5268);
or U5389 (N_5389,N_5200,N_5173);
xor U5390 (N_5390,N_5151,N_5253);
and U5391 (N_5391,N_5193,N_5150);
xnor U5392 (N_5392,N_5210,N_5175);
xor U5393 (N_5393,N_5215,N_5200);
nor U5394 (N_5394,N_5264,N_5185);
nor U5395 (N_5395,N_5134,N_5188);
or U5396 (N_5396,N_5225,N_5159);
and U5397 (N_5397,N_5263,N_5142);
and U5398 (N_5398,N_5162,N_5120);
and U5399 (N_5399,N_5256,N_5193);
xor U5400 (N_5400,N_5152,N_5216);
or U5401 (N_5401,N_5163,N_5156);
and U5402 (N_5402,N_5161,N_5224);
nand U5403 (N_5403,N_5225,N_5261);
or U5404 (N_5404,N_5128,N_5244);
nor U5405 (N_5405,N_5157,N_5230);
xnor U5406 (N_5406,N_5131,N_5211);
xnor U5407 (N_5407,N_5186,N_5177);
xnor U5408 (N_5408,N_5254,N_5233);
nor U5409 (N_5409,N_5231,N_5185);
nor U5410 (N_5410,N_5149,N_5262);
xnor U5411 (N_5411,N_5177,N_5279);
nand U5412 (N_5412,N_5215,N_5153);
xor U5413 (N_5413,N_5164,N_5183);
and U5414 (N_5414,N_5216,N_5217);
or U5415 (N_5415,N_5275,N_5130);
xnor U5416 (N_5416,N_5211,N_5261);
or U5417 (N_5417,N_5174,N_5128);
or U5418 (N_5418,N_5214,N_5254);
nand U5419 (N_5419,N_5126,N_5226);
xnor U5420 (N_5420,N_5251,N_5164);
or U5421 (N_5421,N_5274,N_5238);
nand U5422 (N_5422,N_5212,N_5150);
or U5423 (N_5423,N_5264,N_5139);
or U5424 (N_5424,N_5138,N_5250);
or U5425 (N_5425,N_5163,N_5137);
xor U5426 (N_5426,N_5146,N_5208);
xor U5427 (N_5427,N_5188,N_5200);
nand U5428 (N_5428,N_5260,N_5275);
nor U5429 (N_5429,N_5225,N_5239);
xor U5430 (N_5430,N_5247,N_5133);
xnor U5431 (N_5431,N_5122,N_5159);
nand U5432 (N_5432,N_5197,N_5144);
or U5433 (N_5433,N_5225,N_5245);
or U5434 (N_5434,N_5255,N_5153);
xnor U5435 (N_5435,N_5158,N_5227);
or U5436 (N_5436,N_5152,N_5222);
xnor U5437 (N_5437,N_5242,N_5239);
or U5438 (N_5438,N_5191,N_5196);
xnor U5439 (N_5439,N_5128,N_5207);
or U5440 (N_5440,N_5385,N_5343);
and U5441 (N_5441,N_5401,N_5360);
xnor U5442 (N_5442,N_5366,N_5318);
xnor U5443 (N_5443,N_5287,N_5291);
nor U5444 (N_5444,N_5310,N_5341);
nor U5445 (N_5445,N_5280,N_5365);
nor U5446 (N_5446,N_5409,N_5427);
nand U5447 (N_5447,N_5307,N_5285);
and U5448 (N_5448,N_5299,N_5345);
and U5449 (N_5449,N_5305,N_5375);
nor U5450 (N_5450,N_5439,N_5363);
nand U5451 (N_5451,N_5296,N_5425);
nand U5452 (N_5452,N_5426,N_5316);
nor U5453 (N_5453,N_5382,N_5352);
and U5454 (N_5454,N_5388,N_5403);
nand U5455 (N_5455,N_5300,N_5326);
or U5456 (N_5456,N_5325,N_5428);
xnor U5457 (N_5457,N_5301,N_5367);
nor U5458 (N_5458,N_5294,N_5308);
and U5459 (N_5459,N_5364,N_5356);
and U5460 (N_5460,N_5320,N_5391);
xor U5461 (N_5461,N_5306,N_5405);
and U5462 (N_5462,N_5393,N_5361);
nand U5463 (N_5463,N_5348,N_5377);
nand U5464 (N_5464,N_5317,N_5420);
xnor U5465 (N_5465,N_5336,N_5295);
nand U5466 (N_5466,N_5372,N_5286);
xor U5467 (N_5467,N_5432,N_5340);
or U5468 (N_5468,N_5376,N_5400);
nor U5469 (N_5469,N_5378,N_5394);
nor U5470 (N_5470,N_5435,N_5282);
nor U5471 (N_5471,N_5431,N_5438);
xnor U5472 (N_5472,N_5289,N_5293);
nor U5473 (N_5473,N_5353,N_5332);
nor U5474 (N_5474,N_5304,N_5292);
or U5475 (N_5475,N_5407,N_5381);
nand U5476 (N_5476,N_5335,N_5311);
nand U5477 (N_5477,N_5387,N_5354);
or U5478 (N_5478,N_5290,N_5402);
nor U5479 (N_5479,N_5386,N_5371);
nor U5480 (N_5480,N_5437,N_5339);
and U5481 (N_5481,N_5399,N_5397);
xor U5482 (N_5482,N_5414,N_5314);
nor U5483 (N_5483,N_5302,N_5434);
or U5484 (N_5484,N_5412,N_5324);
or U5485 (N_5485,N_5281,N_5380);
xnor U5486 (N_5486,N_5333,N_5369);
or U5487 (N_5487,N_5408,N_5429);
nor U5488 (N_5488,N_5357,N_5379);
or U5489 (N_5489,N_5358,N_5309);
nor U5490 (N_5490,N_5398,N_5392);
or U5491 (N_5491,N_5350,N_5298);
nor U5492 (N_5492,N_5323,N_5322);
and U5493 (N_5493,N_5327,N_5410);
nor U5494 (N_5494,N_5328,N_5319);
and U5495 (N_5495,N_5284,N_5312);
xnor U5496 (N_5496,N_5373,N_5395);
nand U5497 (N_5497,N_5331,N_5338);
xnor U5498 (N_5498,N_5430,N_5384);
and U5499 (N_5499,N_5417,N_5406);
and U5500 (N_5500,N_5303,N_5423);
or U5501 (N_5501,N_5334,N_5421);
and U5502 (N_5502,N_5337,N_5297);
or U5503 (N_5503,N_5413,N_5415);
or U5504 (N_5504,N_5419,N_5424);
or U5505 (N_5505,N_5359,N_5346);
and U5506 (N_5506,N_5313,N_5347);
and U5507 (N_5507,N_5374,N_5351);
nand U5508 (N_5508,N_5370,N_5396);
nor U5509 (N_5509,N_5389,N_5418);
nand U5510 (N_5510,N_5288,N_5329);
or U5511 (N_5511,N_5321,N_5342);
nand U5512 (N_5512,N_5349,N_5436);
or U5513 (N_5513,N_5383,N_5433);
and U5514 (N_5514,N_5390,N_5368);
or U5515 (N_5515,N_5404,N_5315);
or U5516 (N_5516,N_5416,N_5330);
xor U5517 (N_5517,N_5283,N_5411);
nor U5518 (N_5518,N_5344,N_5355);
nand U5519 (N_5519,N_5422,N_5362);
and U5520 (N_5520,N_5282,N_5387);
nor U5521 (N_5521,N_5361,N_5353);
nor U5522 (N_5522,N_5345,N_5435);
xnor U5523 (N_5523,N_5306,N_5399);
and U5524 (N_5524,N_5373,N_5286);
and U5525 (N_5525,N_5313,N_5330);
xnor U5526 (N_5526,N_5347,N_5338);
nand U5527 (N_5527,N_5347,N_5431);
and U5528 (N_5528,N_5364,N_5430);
and U5529 (N_5529,N_5412,N_5317);
or U5530 (N_5530,N_5362,N_5424);
and U5531 (N_5531,N_5338,N_5299);
nand U5532 (N_5532,N_5412,N_5394);
and U5533 (N_5533,N_5434,N_5373);
nand U5534 (N_5534,N_5432,N_5351);
xor U5535 (N_5535,N_5401,N_5413);
xor U5536 (N_5536,N_5421,N_5322);
or U5537 (N_5537,N_5288,N_5392);
nor U5538 (N_5538,N_5404,N_5341);
and U5539 (N_5539,N_5376,N_5342);
and U5540 (N_5540,N_5401,N_5432);
nand U5541 (N_5541,N_5410,N_5378);
nor U5542 (N_5542,N_5321,N_5334);
nand U5543 (N_5543,N_5286,N_5434);
or U5544 (N_5544,N_5293,N_5338);
nor U5545 (N_5545,N_5361,N_5386);
and U5546 (N_5546,N_5327,N_5367);
and U5547 (N_5547,N_5281,N_5375);
and U5548 (N_5548,N_5282,N_5316);
or U5549 (N_5549,N_5406,N_5291);
xnor U5550 (N_5550,N_5304,N_5424);
or U5551 (N_5551,N_5364,N_5374);
or U5552 (N_5552,N_5389,N_5391);
nor U5553 (N_5553,N_5305,N_5355);
xor U5554 (N_5554,N_5342,N_5295);
nand U5555 (N_5555,N_5324,N_5435);
or U5556 (N_5556,N_5382,N_5407);
or U5557 (N_5557,N_5292,N_5282);
xnor U5558 (N_5558,N_5400,N_5307);
or U5559 (N_5559,N_5315,N_5429);
and U5560 (N_5560,N_5422,N_5284);
and U5561 (N_5561,N_5302,N_5397);
or U5562 (N_5562,N_5427,N_5412);
xnor U5563 (N_5563,N_5383,N_5392);
nor U5564 (N_5564,N_5304,N_5322);
xnor U5565 (N_5565,N_5338,N_5313);
nand U5566 (N_5566,N_5300,N_5325);
or U5567 (N_5567,N_5433,N_5354);
nor U5568 (N_5568,N_5318,N_5421);
xor U5569 (N_5569,N_5296,N_5286);
nor U5570 (N_5570,N_5311,N_5424);
nor U5571 (N_5571,N_5408,N_5384);
and U5572 (N_5572,N_5417,N_5334);
xnor U5573 (N_5573,N_5339,N_5400);
or U5574 (N_5574,N_5420,N_5421);
xor U5575 (N_5575,N_5359,N_5317);
or U5576 (N_5576,N_5333,N_5410);
xnor U5577 (N_5577,N_5368,N_5355);
nand U5578 (N_5578,N_5424,N_5282);
and U5579 (N_5579,N_5355,N_5429);
nand U5580 (N_5580,N_5377,N_5428);
or U5581 (N_5581,N_5370,N_5401);
xor U5582 (N_5582,N_5362,N_5387);
nor U5583 (N_5583,N_5321,N_5421);
xor U5584 (N_5584,N_5427,N_5281);
nor U5585 (N_5585,N_5366,N_5317);
nor U5586 (N_5586,N_5337,N_5384);
xor U5587 (N_5587,N_5354,N_5314);
or U5588 (N_5588,N_5401,N_5405);
or U5589 (N_5589,N_5326,N_5344);
or U5590 (N_5590,N_5433,N_5298);
or U5591 (N_5591,N_5325,N_5410);
nand U5592 (N_5592,N_5339,N_5302);
xor U5593 (N_5593,N_5297,N_5415);
or U5594 (N_5594,N_5431,N_5340);
nor U5595 (N_5595,N_5415,N_5291);
nand U5596 (N_5596,N_5309,N_5427);
and U5597 (N_5597,N_5359,N_5338);
and U5598 (N_5598,N_5406,N_5354);
and U5599 (N_5599,N_5312,N_5313);
nand U5600 (N_5600,N_5593,N_5557);
xnor U5601 (N_5601,N_5582,N_5591);
xor U5602 (N_5602,N_5500,N_5449);
xnor U5603 (N_5603,N_5563,N_5466);
nand U5604 (N_5604,N_5541,N_5577);
nand U5605 (N_5605,N_5578,N_5546);
nand U5606 (N_5606,N_5517,N_5553);
nand U5607 (N_5607,N_5492,N_5446);
xor U5608 (N_5608,N_5508,N_5467);
nand U5609 (N_5609,N_5544,N_5540);
nand U5610 (N_5610,N_5512,N_5496);
and U5611 (N_5611,N_5444,N_5549);
and U5612 (N_5612,N_5441,N_5484);
or U5613 (N_5613,N_5531,N_5586);
or U5614 (N_5614,N_5580,N_5583);
xnor U5615 (N_5615,N_5474,N_5471);
nor U5616 (N_5616,N_5548,N_5522);
or U5617 (N_5617,N_5568,N_5463);
nand U5618 (N_5618,N_5559,N_5481);
and U5619 (N_5619,N_5573,N_5485);
xor U5620 (N_5620,N_5585,N_5454);
xnor U5621 (N_5621,N_5489,N_5558);
or U5622 (N_5622,N_5535,N_5459);
and U5623 (N_5623,N_5547,N_5507);
or U5624 (N_5624,N_5543,N_5502);
nor U5625 (N_5625,N_5592,N_5464);
xnor U5626 (N_5626,N_5472,N_5457);
xnor U5627 (N_5627,N_5551,N_5536);
nand U5628 (N_5628,N_5453,N_5598);
nor U5629 (N_5629,N_5462,N_5581);
and U5630 (N_5630,N_5497,N_5560);
nor U5631 (N_5631,N_5482,N_5594);
nand U5632 (N_5632,N_5579,N_5555);
and U5633 (N_5633,N_5509,N_5530);
nand U5634 (N_5634,N_5493,N_5513);
or U5635 (N_5635,N_5554,N_5576);
nand U5636 (N_5636,N_5473,N_5452);
xor U5637 (N_5637,N_5514,N_5488);
xnor U5638 (N_5638,N_5528,N_5504);
nand U5639 (N_5639,N_5519,N_5539);
or U5640 (N_5640,N_5562,N_5440);
xor U5641 (N_5641,N_5498,N_5542);
xnor U5642 (N_5642,N_5589,N_5461);
nor U5643 (N_5643,N_5564,N_5534);
and U5644 (N_5644,N_5458,N_5566);
and U5645 (N_5645,N_5529,N_5584);
and U5646 (N_5646,N_5483,N_5561);
nand U5647 (N_5647,N_5537,N_5516);
nand U5648 (N_5648,N_5468,N_5532);
nor U5649 (N_5649,N_5445,N_5590);
and U5650 (N_5650,N_5490,N_5523);
xnor U5651 (N_5651,N_5491,N_5556);
or U5652 (N_5652,N_5574,N_5477);
nand U5653 (N_5653,N_5518,N_5487);
nor U5654 (N_5654,N_5443,N_5495);
and U5655 (N_5655,N_5569,N_5499);
xnor U5656 (N_5656,N_5501,N_5479);
or U5657 (N_5657,N_5597,N_5476);
or U5658 (N_5658,N_5469,N_5465);
xnor U5659 (N_5659,N_5470,N_5588);
nor U5660 (N_5660,N_5494,N_5521);
nand U5661 (N_5661,N_5455,N_5525);
nand U5662 (N_5662,N_5538,N_5550);
nor U5663 (N_5663,N_5460,N_5599);
xnor U5664 (N_5664,N_5596,N_5526);
nor U5665 (N_5665,N_5527,N_5447);
nor U5666 (N_5666,N_5587,N_5450);
or U5667 (N_5667,N_5475,N_5478);
xor U5668 (N_5668,N_5505,N_5503);
and U5669 (N_5669,N_5510,N_5515);
nor U5670 (N_5670,N_5442,N_5524);
and U5671 (N_5671,N_5480,N_5595);
nand U5672 (N_5672,N_5506,N_5451);
and U5673 (N_5673,N_5456,N_5567);
xnor U5674 (N_5674,N_5533,N_5511);
nor U5675 (N_5675,N_5448,N_5575);
nor U5676 (N_5676,N_5570,N_5545);
or U5677 (N_5677,N_5565,N_5520);
nor U5678 (N_5678,N_5572,N_5552);
xor U5679 (N_5679,N_5571,N_5486);
or U5680 (N_5680,N_5495,N_5594);
and U5681 (N_5681,N_5569,N_5442);
xor U5682 (N_5682,N_5554,N_5465);
and U5683 (N_5683,N_5449,N_5480);
xor U5684 (N_5684,N_5455,N_5596);
nand U5685 (N_5685,N_5529,N_5467);
and U5686 (N_5686,N_5511,N_5577);
nand U5687 (N_5687,N_5571,N_5497);
xnor U5688 (N_5688,N_5485,N_5489);
or U5689 (N_5689,N_5450,N_5584);
xnor U5690 (N_5690,N_5492,N_5487);
and U5691 (N_5691,N_5452,N_5488);
and U5692 (N_5692,N_5519,N_5599);
and U5693 (N_5693,N_5462,N_5563);
nor U5694 (N_5694,N_5537,N_5458);
and U5695 (N_5695,N_5454,N_5536);
and U5696 (N_5696,N_5527,N_5599);
or U5697 (N_5697,N_5496,N_5491);
xnor U5698 (N_5698,N_5581,N_5486);
nand U5699 (N_5699,N_5547,N_5451);
nor U5700 (N_5700,N_5489,N_5594);
xnor U5701 (N_5701,N_5599,N_5490);
nor U5702 (N_5702,N_5452,N_5570);
or U5703 (N_5703,N_5464,N_5530);
nor U5704 (N_5704,N_5528,N_5460);
or U5705 (N_5705,N_5563,N_5459);
nand U5706 (N_5706,N_5562,N_5471);
xnor U5707 (N_5707,N_5511,N_5585);
xnor U5708 (N_5708,N_5574,N_5554);
xnor U5709 (N_5709,N_5519,N_5484);
nand U5710 (N_5710,N_5586,N_5574);
nor U5711 (N_5711,N_5547,N_5462);
and U5712 (N_5712,N_5580,N_5501);
and U5713 (N_5713,N_5539,N_5569);
and U5714 (N_5714,N_5586,N_5549);
nor U5715 (N_5715,N_5550,N_5558);
xor U5716 (N_5716,N_5445,N_5534);
and U5717 (N_5717,N_5493,N_5555);
xnor U5718 (N_5718,N_5460,N_5556);
xnor U5719 (N_5719,N_5547,N_5599);
xor U5720 (N_5720,N_5474,N_5482);
or U5721 (N_5721,N_5509,N_5584);
xor U5722 (N_5722,N_5571,N_5506);
nor U5723 (N_5723,N_5550,N_5503);
xor U5724 (N_5724,N_5541,N_5487);
xor U5725 (N_5725,N_5504,N_5484);
nor U5726 (N_5726,N_5457,N_5477);
nor U5727 (N_5727,N_5445,N_5500);
or U5728 (N_5728,N_5555,N_5537);
and U5729 (N_5729,N_5539,N_5498);
nand U5730 (N_5730,N_5456,N_5524);
or U5731 (N_5731,N_5563,N_5536);
nand U5732 (N_5732,N_5472,N_5542);
and U5733 (N_5733,N_5487,N_5464);
xor U5734 (N_5734,N_5476,N_5504);
and U5735 (N_5735,N_5457,N_5563);
and U5736 (N_5736,N_5576,N_5494);
nand U5737 (N_5737,N_5504,N_5589);
and U5738 (N_5738,N_5481,N_5582);
nor U5739 (N_5739,N_5513,N_5475);
or U5740 (N_5740,N_5535,N_5598);
xor U5741 (N_5741,N_5515,N_5589);
xor U5742 (N_5742,N_5598,N_5464);
nand U5743 (N_5743,N_5494,N_5539);
nor U5744 (N_5744,N_5509,N_5531);
nand U5745 (N_5745,N_5506,N_5563);
or U5746 (N_5746,N_5453,N_5444);
nand U5747 (N_5747,N_5517,N_5546);
nand U5748 (N_5748,N_5506,N_5525);
nand U5749 (N_5749,N_5492,N_5462);
nand U5750 (N_5750,N_5534,N_5543);
and U5751 (N_5751,N_5546,N_5443);
nor U5752 (N_5752,N_5454,N_5566);
and U5753 (N_5753,N_5487,N_5592);
and U5754 (N_5754,N_5463,N_5596);
nor U5755 (N_5755,N_5509,N_5534);
nor U5756 (N_5756,N_5469,N_5583);
or U5757 (N_5757,N_5459,N_5440);
nand U5758 (N_5758,N_5593,N_5520);
nand U5759 (N_5759,N_5590,N_5477);
nor U5760 (N_5760,N_5686,N_5670);
and U5761 (N_5761,N_5642,N_5606);
xnor U5762 (N_5762,N_5632,N_5664);
xor U5763 (N_5763,N_5759,N_5754);
and U5764 (N_5764,N_5658,N_5728);
or U5765 (N_5765,N_5655,N_5740);
xor U5766 (N_5766,N_5648,N_5604);
nor U5767 (N_5767,N_5704,N_5674);
nor U5768 (N_5768,N_5753,N_5628);
nor U5769 (N_5769,N_5603,N_5690);
or U5770 (N_5770,N_5697,N_5739);
and U5771 (N_5771,N_5716,N_5649);
xor U5772 (N_5772,N_5645,N_5668);
and U5773 (N_5773,N_5630,N_5680);
and U5774 (N_5774,N_5676,N_5617);
and U5775 (N_5775,N_5685,N_5640);
nor U5776 (N_5776,N_5743,N_5756);
nor U5777 (N_5777,N_5755,N_5726);
nor U5778 (N_5778,N_5737,N_5602);
xnor U5779 (N_5779,N_5656,N_5695);
nand U5780 (N_5780,N_5675,N_5744);
xnor U5781 (N_5781,N_5652,N_5751);
and U5782 (N_5782,N_5605,N_5727);
nand U5783 (N_5783,N_5644,N_5681);
or U5784 (N_5784,N_5693,N_5738);
nand U5785 (N_5785,N_5663,N_5742);
and U5786 (N_5786,N_5620,N_5608);
nand U5787 (N_5787,N_5752,N_5667);
nor U5788 (N_5788,N_5710,N_5627);
nor U5789 (N_5789,N_5748,N_5747);
nand U5790 (N_5790,N_5700,N_5689);
xor U5791 (N_5791,N_5672,N_5646);
xnor U5792 (N_5792,N_5696,N_5757);
nor U5793 (N_5793,N_5708,N_5724);
xnor U5794 (N_5794,N_5625,N_5731);
and U5795 (N_5795,N_5651,N_5641);
nor U5796 (N_5796,N_5682,N_5707);
nor U5797 (N_5797,N_5687,N_5612);
or U5798 (N_5798,N_5719,N_5673);
and U5799 (N_5799,N_5643,N_5732);
xor U5800 (N_5800,N_5715,N_5611);
and U5801 (N_5801,N_5713,N_5650);
nor U5802 (N_5802,N_5720,N_5709);
or U5803 (N_5803,N_5725,N_5653);
or U5804 (N_5804,N_5698,N_5657);
or U5805 (N_5805,N_5647,N_5691);
nor U5806 (N_5806,N_5679,N_5634);
or U5807 (N_5807,N_5736,N_5749);
or U5808 (N_5808,N_5741,N_5631);
or U5809 (N_5809,N_5619,N_5750);
or U5810 (N_5810,N_5722,N_5692);
nand U5811 (N_5811,N_5626,N_5613);
and U5812 (N_5812,N_5601,N_5729);
and U5813 (N_5813,N_5607,N_5660);
or U5814 (N_5814,N_5671,N_5661);
nand U5815 (N_5815,N_5712,N_5714);
and U5816 (N_5816,N_5614,N_5622);
nand U5817 (N_5817,N_5621,N_5688);
nand U5818 (N_5818,N_5733,N_5677);
xor U5819 (N_5819,N_5702,N_5683);
nand U5820 (N_5820,N_5637,N_5610);
and U5821 (N_5821,N_5735,N_5703);
nand U5822 (N_5822,N_5758,N_5629);
or U5823 (N_5823,N_5624,N_5699);
xor U5824 (N_5824,N_5666,N_5600);
nand U5825 (N_5825,N_5705,N_5718);
xor U5826 (N_5826,N_5706,N_5665);
xnor U5827 (N_5827,N_5684,N_5659);
nor U5828 (N_5828,N_5669,N_5717);
nand U5829 (N_5829,N_5730,N_5615);
or U5830 (N_5830,N_5721,N_5701);
or U5831 (N_5831,N_5623,N_5723);
nand U5832 (N_5832,N_5616,N_5694);
xnor U5833 (N_5833,N_5639,N_5618);
or U5834 (N_5834,N_5636,N_5734);
nor U5835 (N_5835,N_5638,N_5745);
and U5836 (N_5836,N_5633,N_5746);
nor U5837 (N_5837,N_5711,N_5635);
nand U5838 (N_5838,N_5678,N_5609);
nor U5839 (N_5839,N_5662,N_5654);
xnor U5840 (N_5840,N_5670,N_5729);
xor U5841 (N_5841,N_5637,N_5755);
and U5842 (N_5842,N_5636,N_5681);
nor U5843 (N_5843,N_5759,N_5734);
and U5844 (N_5844,N_5743,N_5600);
and U5845 (N_5845,N_5759,N_5706);
nand U5846 (N_5846,N_5611,N_5722);
nor U5847 (N_5847,N_5669,N_5624);
nor U5848 (N_5848,N_5601,N_5619);
nand U5849 (N_5849,N_5644,N_5667);
nand U5850 (N_5850,N_5650,N_5728);
and U5851 (N_5851,N_5750,N_5610);
nand U5852 (N_5852,N_5621,N_5742);
nand U5853 (N_5853,N_5613,N_5753);
xnor U5854 (N_5854,N_5685,N_5749);
nor U5855 (N_5855,N_5723,N_5709);
or U5856 (N_5856,N_5667,N_5753);
or U5857 (N_5857,N_5604,N_5651);
or U5858 (N_5858,N_5625,N_5713);
or U5859 (N_5859,N_5617,N_5724);
xor U5860 (N_5860,N_5747,N_5706);
nand U5861 (N_5861,N_5691,N_5714);
or U5862 (N_5862,N_5740,N_5604);
nor U5863 (N_5863,N_5694,N_5631);
xor U5864 (N_5864,N_5745,N_5691);
and U5865 (N_5865,N_5710,N_5662);
nor U5866 (N_5866,N_5626,N_5686);
nor U5867 (N_5867,N_5607,N_5715);
nand U5868 (N_5868,N_5709,N_5724);
nand U5869 (N_5869,N_5682,N_5635);
nand U5870 (N_5870,N_5675,N_5631);
or U5871 (N_5871,N_5694,N_5660);
nor U5872 (N_5872,N_5741,N_5636);
and U5873 (N_5873,N_5614,N_5692);
or U5874 (N_5874,N_5688,N_5681);
nand U5875 (N_5875,N_5687,N_5710);
nor U5876 (N_5876,N_5730,N_5693);
nor U5877 (N_5877,N_5655,N_5738);
nand U5878 (N_5878,N_5603,N_5622);
xor U5879 (N_5879,N_5633,N_5690);
nand U5880 (N_5880,N_5622,N_5628);
or U5881 (N_5881,N_5643,N_5744);
and U5882 (N_5882,N_5686,N_5652);
and U5883 (N_5883,N_5667,N_5703);
nand U5884 (N_5884,N_5671,N_5665);
and U5885 (N_5885,N_5704,N_5711);
nor U5886 (N_5886,N_5746,N_5664);
nand U5887 (N_5887,N_5611,N_5749);
or U5888 (N_5888,N_5653,N_5742);
nand U5889 (N_5889,N_5650,N_5652);
nand U5890 (N_5890,N_5699,N_5656);
nor U5891 (N_5891,N_5703,N_5717);
and U5892 (N_5892,N_5747,N_5714);
nor U5893 (N_5893,N_5653,N_5680);
nor U5894 (N_5894,N_5676,N_5726);
nor U5895 (N_5895,N_5724,N_5671);
nand U5896 (N_5896,N_5687,N_5759);
and U5897 (N_5897,N_5756,N_5649);
xor U5898 (N_5898,N_5639,N_5675);
or U5899 (N_5899,N_5649,N_5631);
and U5900 (N_5900,N_5664,N_5607);
xnor U5901 (N_5901,N_5642,N_5742);
and U5902 (N_5902,N_5726,N_5735);
or U5903 (N_5903,N_5636,N_5634);
nor U5904 (N_5904,N_5657,N_5755);
nor U5905 (N_5905,N_5616,N_5667);
nor U5906 (N_5906,N_5687,N_5708);
or U5907 (N_5907,N_5675,N_5648);
and U5908 (N_5908,N_5698,N_5639);
nand U5909 (N_5909,N_5735,N_5605);
xor U5910 (N_5910,N_5630,N_5732);
and U5911 (N_5911,N_5669,N_5612);
xor U5912 (N_5912,N_5728,N_5735);
nand U5913 (N_5913,N_5750,N_5646);
nor U5914 (N_5914,N_5671,N_5734);
nor U5915 (N_5915,N_5683,N_5708);
xor U5916 (N_5916,N_5733,N_5608);
and U5917 (N_5917,N_5670,N_5709);
and U5918 (N_5918,N_5677,N_5720);
nor U5919 (N_5919,N_5687,N_5691);
or U5920 (N_5920,N_5781,N_5812);
xnor U5921 (N_5921,N_5860,N_5890);
and U5922 (N_5922,N_5879,N_5824);
or U5923 (N_5923,N_5807,N_5770);
nand U5924 (N_5924,N_5856,N_5853);
xor U5925 (N_5925,N_5771,N_5904);
nand U5926 (N_5926,N_5817,N_5844);
nand U5927 (N_5927,N_5864,N_5836);
or U5928 (N_5928,N_5785,N_5783);
nand U5929 (N_5929,N_5828,N_5786);
or U5930 (N_5930,N_5767,N_5827);
xnor U5931 (N_5931,N_5808,N_5845);
xor U5932 (N_5932,N_5892,N_5862);
xnor U5933 (N_5933,N_5787,N_5800);
nor U5934 (N_5934,N_5766,N_5822);
and U5935 (N_5935,N_5791,N_5867);
or U5936 (N_5936,N_5772,N_5857);
and U5937 (N_5937,N_5778,N_5872);
and U5938 (N_5938,N_5881,N_5790);
nand U5939 (N_5939,N_5915,N_5842);
nand U5940 (N_5940,N_5826,N_5764);
xor U5941 (N_5941,N_5789,N_5810);
nor U5942 (N_5942,N_5788,N_5779);
nand U5943 (N_5943,N_5768,N_5798);
nand U5944 (N_5944,N_5773,N_5899);
nor U5945 (N_5945,N_5849,N_5884);
xor U5946 (N_5946,N_5775,N_5896);
and U5947 (N_5947,N_5792,N_5901);
or U5948 (N_5948,N_5865,N_5820);
xnor U5949 (N_5949,N_5893,N_5762);
nor U5950 (N_5950,N_5910,N_5917);
or U5951 (N_5951,N_5876,N_5794);
nor U5952 (N_5952,N_5804,N_5843);
nand U5953 (N_5953,N_5908,N_5765);
nor U5954 (N_5954,N_5760,N_5914);
and U5955 (N_5955,N_5784,N_5883);
xor U5956 (N_5956,N_5852,N_5913);
nor U5957 (N_5957,N_5868,N_5911);
and U5958 (N_5958,N_5858,N_5895);
nand U5959 (N_5959,N_5796,N_5851);
nor U5960 (N_5960,N_5854,N_5825);
and U5961 (N_5961,N_5906,N_5806);
or U5962 (N_5962,N_5774,N_5912);
nand U5963 (N_5963,N_5894,N_5833);
nor U5964 (N_5964,N_5839,N_5855);
or U5965 (N_5965,N_5863,N_5830);
nand U5966 (N_5966,N_5815,N_5882);
and U5967 (N_5967,N_5837,N_5887);
nand U5968 (N_5968,N_5918,N_5776);
nor U5969 (N_5969,N_5793,N_5885);
and U5970 (N_5970,N_5818,N_5823);
xnor U5971 (N_5971,N_5761,N_5831);
nor U5972 (N_5972,N_5907,N_5900);
and U5973 (N_5973,N_5799,N_5813);
or U5974 (N_5974,N_5834,N_5763);
and U5975 (N_5975,N_5877,N_5847);
and U5976 (N_5976,N_5898,N_5873);
and U5977 (N_5977,N_5841,N_5909);
or U5978 (N_5978,N_5866,N_5874);
and U5979 (N_5979,N_5916,N_5811);
and U5980 (N_5980,N_5919,N_5878);
or U5981 (N_5981,N_5861,N_5903);
or U5982 (N_5982,N_5880,N_5797);
xor U5983 (N_5983,N_5886,N_5805);
or U5984 (N_5984,N_5782,N_5869);
nand U5985 (N_5985,N_5870,N_5809);
xnor U5986 (N_5986,N_5802,N_5897);
xnor U5987 (N_5987,N_5795,N_5888);
and U5988 (N_5988,N_5838,N_5835);
nor U5989 (N_5989,N_5821,N_5840);
or U5990 (N_5990,N_5891,N_5846);
or U5991 (N_5991,N_5848,N_5819);
and U5992 (N_5992,N_5875,N_5780);
xnor U5993 (N_5993,N_5769,N_5814);
xnor U5994 (N_5994,N_5859,N_5777);
and U5995 (N_5995,N_5889,N_5829);
nand U5996 (N_5996,N_5902,N_5871);
xnor U5997 (N_5997,N_5850,N_5832);
and U5998 (N_5998,N_5816,N_5905);
and U5999 (N_5999,N_5801,N_5803);
and U6000 (N_6000,N_5781,N_5884);
and U6001 (N_6001,N_5813,N_5866);
and U6002 (N_6002,N_5888,N_5865);
xor U6003 (N_6003,N_5844,N_5826);
and U6004 (N_6004,N_5770,N_5819);
nand U6005 (N_6005,N_5801,N_5762);
nor U6006 (N_6006,N_5841,N_5767);
nor U6007 (N_6007,N_5802,N_5777);
xor U6008 (N_6008,N_5761,N_5824);
or U6009 (N_6009,N_5909,N_5839);
xor U6010 (N_6010,N_5826,N_5773);
or U6011 (N_6011,N_5917,N_5831);
or U6012 (N_6012,N_5789,N_5840);
xor U6013 (N_6013,N_5794,N_5783);
nor U6014 (N_6014,N_5853,N_5912);
xnor U6015 (N_6015,N_5833,N_5842);
nand U6016 (N_6016,N_5808,N_5846);
or U6017 (N_6017,N_5799,N_5876);
nand U6018 (N_6018,N_5779,N_5859);
nor U6019 (N_6019,N_5779,N_5789);
nand U6020 (N_6020,N_5919,N_5793);
or U6021 (N_6021,N_5886,N_5783);
xnor U6022 (N_6022,N_5772,N_5767);
nand U6023 (N_6023,N_5791,N_5777);
nand U6024 (N_6024,N_5862,N_5805);
and U6025 (N_6025,N_5845,N_5905);
xor U6026 (N_6026,N_5854,N_5781);
nor U6027 (N_6027,N_5873,N_5880);
nor U6028 (N_6028,N_5790,N_5851);
nor U6029 (N_6029,N_5909,N_5910);
nand U6030 (N_6030,N_5860,N_5883);
and U6031 (N_6031,N_5918,N_5852);
nor U6032 (N_6032,N_5765,N_5778);
nand U6033 (N_6033,N_5872,N_5780);
xor U6034 (N_6034,N_5768,N_5825);
and U6035 (N_6035,N_5868,N_5892);
nor U6036 (N_6036,N_5813,N_5905);
nand U6037 (N_6037,N_5917,N_5912);
or U6038 (N_6038,N_5833,N_5829);
nand U6039 (N_6039,N_5912,N_5913);
nand U6040 (N_6040,N_5868,N_5795);
nand U6041 (N_6041,N_5910,N_5857);
or U6042 (N_6042,N_5823,N_5801);
or U6043 (N_6043,N_5800,N_5843);
or U6044 (N_6044,N_5820,N_5915);
and U6045 (N_6045,N_5765,N_5812);
and U6046 (N_6046,N_5886,N_5791);
or U6047 (N_6047,N_5802,N_5842);
xnor U6048 (N_6048,N_5873,N_5917);
nand U6049 (N_6049,N_5785,N_5762);
or U6050 (N_6050,N_5846,N_5816);
nand U6051 (N_6051,N_5789,N_5915);
and U6052 (N_6052,N_5881,N_5763);
xnor U6053 (N_6053,N_5808,N_5893);
and U6054 (N_6054,N_5768,N_5773);
xor U6055 (N_6055,N_5869,N_5773);
and U6056 (N_6056,N_5764,N_5786);
nor U6057 (N_6057,N_5913,N_5860);
or U6058 (N_6058,N_5774,N_5800);
nand U6059 (N_6059,N_5857,N_5882);
or U6060 (N_6060,N_5771,N_5881);
and U6061 (N_6061,N_5896,N_5899);
and U6062 (N_6062,N_5915,N_5888);
and U6063 (N_6063,N_5880,N_5761);
nor U6064 (N_6064,N_5834,N_5821);
nor U6065 (N_6065,N_5760,N_5889);
or U6066 (N_6066,N_5809,N_5802);
nand U6067 (N_6067,N_5783,N_5891);
nor U6068 (N_6068,N_5831,N_5791);
nor U6069 (N_6069,N_5802,N_5878);
nor U6070 (N_6070,N_5843,N_5772);
xor U6071 (N_6071,N_5780,N_5832);
and U6072 (N_6072,N_5822,N_5914);
and U6073 (N_6073,N_5770,N_5827);
or U6074 (N_6074,N_5846,N_5841);
xnor U6075 (N_6075,N_5836,N_5878);
and U6076 (N_6076,N_5791,N_5784);
or U6077 (N_6077,N_5782,N_5795);
nor U6078 (N_6078,N_5894,N_5901);
nand U6079 (N_6079,N_5764,N_5818);
and U6080 (N_6080,N_6028,N_6035);
and U6081 (N_6081,N_6072,N_6046);
xnor U6082 (N_6082,N_6030,N_6049);
xnor U6083 (N_6083,N_6025,N_5959);
nor U6084 (N_6084,N_6020,N_6011);
nor U6085 (N_6085,N_6054,N_5957);
or U6086 (N_6086,N_6068,N_5933);
nand U6087 (N_6087,N_6058,N_5982);
or U6088 (N_6088,N_5925,N_5920);
or U6089 (N_6089,N_5922,N_5943);
nand U6090 (N_6090,N_5953,N_6022);
or U6091 (N_6091,N_6012,N_6055);
nand U6092 (N_6092,N_6036,N_6008);
or U6093 (N_6093,N_5954,N_6015);
xor U6094 (N_6094,N_5991,N_6041);
xor U6095 (N_6095,N_6040,N_5958);
or U6096 (N_6096,N_6067,N_6002);
or U6097 (N_6097,N_6053,N_5992);
nor U6098 (N_6098,N_6018,N_6066);
and U6099 (N_6099,N_6014,N_6075);
nand U6100 (N_6100,N_6038,N_5952);
nor U6101 (N_6101,N_6027,N_5976);
xor U6102 (N_6102,N_5944,N_6061);
nor U6103 (N_6103,N_5989,N_5980);
and U6104 (N_6104,N_5950,N_6048);
xnor U6105 (N_6105,N_5935,N_5940);
nor U6106 (N_6106,N_6043,N_5985);
and U6107 (N_6107,N_5936,N_6039);
or U6108 (N_6108,N_6042,N_5948);
and U6109 (N_6109,N_5968,N_6033);
nand U6110 (N_6110,N_6057,N_6076);
nand U6111 (N_6111,N_6073,N_6047);
or U6112 (N_6112,N_5961,N_5973);
or U6113 (N_6113,N_5941,N_6001);
or U6114 (N_6114,N_5994,N_5966);
nor U6115 (N_6115,N_6071,N_6070);
nand U6116 (N_6116,N_5977,N_6034);
or U6117 (N_6117,N_5962,N_6006);
xnor U6118 (N_6118,N_5956,N_5981);
xor U6119 (N_6119,N_6069,N_5923);
or U6120 (N_6120,N_5937,N_5986);
nor U6121 (N_6121,N_6037,N_6024);
nor U6122 (N_6122,N_5988,N_5947);
xor U6123 (N_6123,N_5975,N_5999);
nor U6124 (N_6124,N_6013,N_5987);
nand U6125 (N_6125,N_5963,N_5932);
or U6126 (N_6126,N_5942,N_5983);
nor U6127 (N_6127,N_5990,N_6009);
or U6128 (N_6128,N_5960,N_6031);
xnor U6129 (N_6129,N_5934,N_5946);
or U6130 (N_6130,N_6063,N_5921);
and U6131 (N_6131,N_5984,N_6032);
nor U6132 (N_6132,N_6017,N_5931);
nor U6133 (N_6133,N_5997,N_5939);
and U6134 (N_6134,N_5928,N_6045);
or U6135 (N_6135,N_6029,N_5971);
nor U6136 (N_6136,N_5926,N_6051);
and U6137 (N_6137,N_6044,N_5998);
and U6138 (N_6138,N_6004,N_6064);
xnor U6139 (N_6139,N_5993,N_5930);
nor U6140 (N_6140,N_5967,N_5965);
xor U6141 (N_6141,N_5924,N_6023);
and U6142 (N_6142,N_6079,N_5995);
nor U6143 (N_6143,N_6010,N_6078);
nand U6144 (N_6144,N_6052,N_5927);
and U6145 (N_6145,N_6050,N_5938);
and U6146 (N_6146,N_6060,N_5951);
and U6147 (N_6147,N_6074,N_6005);
xnor U6148 (N_6148,N_6062,N_6003);
nand U6149 (N_6149,N_6077,N_5964);
and U6150 (N_6150,N_6019,N_6007);
and U6151 (N_6151,N_6026,N_6059);
nor U6152 (N_6152,N_5979,N_6056);
or U6153 (N_6153,N_5972,N_5996);
xnor U6154 (N_6154,N_5978,N_6021);
nor U6155 (N_6155,N_5969,N_5949);
and U6156 (N_6156,N_6016,N_6000);
and U6157 (N_6157,N_5970,N_5955);
nor U6158 (N_6158,N_5974,N_5929);
nand U6159 (N_6159,N_6065,N_5945);
or U6160 (N_6160,N_5968,N_5933);
xnor U6161 (N_6161,N_6043,N_6013);
and U6162 (N_6162,N_5964,N_5935);
nor U6163 (N_6163,N_6066,N_5995);
nand U6164 (N_6164,N_6063,N_5927);
and U6165 (N_6165,N_6034,N_6067);
nor U6166 (N_6166,N_5973,N_5920);
nor U6167 (N_6167,N_6013,N_5989);
nand U6168 (N_6168,N_5975,N_6037);
and U6169 (N_6169,N_6020,N_5977);
and U6170 (N_6170,N_6064,N_5951);
xor U6171 (N_6171,N_5927,N_6074);
xnor U6172 (N_6172,N_6030,N_6058);
and U6173 (N_6173,N_6005,N_5921);
nand U6174 (N_6174,N_6041,N_5953);
and U6175 (N_6175,N_5989,N_6032);
xor U6176 (N_6176,N_5953,N_5941);
nand U6177 (N_6177,N_6062,N_5931);
xor U6178 (N_6178,N_5930,N_5937);
nor U6179 (N_6179,N_6011,N_5973);
nor U6180 (N_6180,N_5938,N_5932);
or U6181 (N_6181,N_6073,N_5931);
and U6182 (N_6182,N_5981,N_5960);
and U6183 (N_6183,N_5956,N_5989);
nand U6184 (N_6184,N_5950,N_5964);
nor U6185 (N_6185,N_6037,N_6033);
nor U6186 (N_6186,N_6028,N_5986);
or U6187 (N_6187,N_6064,N_5995);
nor U6188 (N_6188,N_6002,N_6056);
and U6189 (N_6189,N_6061,N_5968);
nor U6190 (N_6190,N_5947,N_6079);
nor U6191 (N_6191,N_6075,N_6051);
xnor U6192 (N_6192,N_5978,N_5967);
or U6193 (N_6193,N_5953,N_6052);
nand U6194 (N_6194,N_5939,N_6058);
or U6195 (N_6195,N_6035,N_6075);
nand U6196 (N_6196,N_6043,N_6006);
nor U6197 (N_6197,N_6059,N_6013);
xor U6198 (N_6198,N_6057,N_5927);
or U6199 (N_6199,N_6039,N_6031);
or U6200 (N_6200,N_6033,N_5952);
nand U6201 (N_6201,N_5948,N_5988);
nor U6202 (N_6202,N_5944,N_5994);
nor U6203 (N_6203,N_6019,N_5972);
nand U6204 (N_6204,N_5992,N_5934);
nand U6205 (N_6205,N_5966,N_6055);
nor U6206 (N_6206,N_6011,N_6065);
and U6207 (N_6207,N_5973,N_6073);
or U6208 (N_6208,N_5933,N_5938);
and U6209 (N_6209,N_5935,N_5961);
and U6210 (N_6210,N_6079,N_5999);
nor U6211 (N_6211,N_5980,N_6041);
or U6212 (N_6212,N_5997,N_6057);
nand U6213 (N_6213,N_5981,N_5967);
and U6214 (N_6214,N_6013,N_5957);
or U6215 (N_6215,N_5921,N_5930);
xor U6216 (N_6216,N_6010,N_6079);
or U6217 (N_6217,N_5997,N_5920);
and U6218 (N_6218,N_6074,N_5932);
or U6219 (N_6219,N_6012,N_5930);
or U6220 (N_6220,N_6031,N_6079);
nand U6221 (N_6221,N_6054,N_6072);
nor U6222 (N_6222,N_6051,N_5934);
nand U6223 (N_6223,N_5944,N_5925);
and U6224 (N_6224,N_5923,N_6060);
and U6225 (N_6225,N_5979,N_6079);
nand U6226 (N_6226,N_5966,N_5937);
and U6227 (N_6227,N_6011,N_5958);
and U6228 (N_6228,N_6071,N_6043);
xor U6229 (N_6229,N_5998,N_6060);
xor U6230 (N_6230,N_6007,N_6017);
nor U6231 (N_6231,N_5942,N_5948);
or U6232 (N_6232,N_5963,N_5958);
nand U6233 (N_6233,N_5967,N_6021);
nor U6234 (N_6234,N_6031,N_6027);
xnor U6235 (N_6235,N_6026,N_6037);
nor U6236 (N_6236,N_5985,N_6060);
nand U6237 (N_6237,N_5976,N_6015);
or U6238 (N_6238,N_6020,N_6053);
xor U6239 (N_6239,N_5990,N_6069);
xor U6240 (N_6240,N_6160,N_6087);
nand U6241 (N_6241,N_6111,N_6179);
nor U6242 (N_6242,N_6163,N_6101);
xor U6243 (N_6243,N_6177,N_6108);
nor U6244 (N_6244,N_6229,N_6178);
nor U6245 (N_6245,N_6081,N_6188);
nor U6246 (N_6246,N_6225,N_6143);
nor U6247 (N_6247,N_6202,N_6237);
or U6248 (N_6248,N_6086,N_6218);
or U6249 (N_6249,N_6103,N_6094);
and U6250 (N_6250,N_6084,N_6230);
xnor U6251 (N_6251,N_6167,N_6092);
xor U6252 (N_6252,N_6114,N_6110);
xnor U6253 (N_6253,N_6093,N_6161);
nor U6254 (N_6254,N_6159,N_6200);
or U6255 (N_6255,N_6238,N_6236);
and U6256 (N_6256,N_6105,N_6102);
xnor U6257 (N_6257,N_6142,N_6139);
nand U6258 (N_6258,N_6109,N_6239);
nand U6259 (N_6259,N_6234,N_6121);
nor U6260 (N_6260,N_6150,N_6158);
or U6261 (N_6261,N_6164,N_6082);
nor U6262 (N_6262,N_6222,N_6186);
or U6263 (N_6263,N_6232,N_6138);
and U6264 (N_6264,N_6132,N_6195);
nand U6265 (N_6265,N_6080,N_6180);
nor U6266 (N_6266,N_6137,N_6223);
and U6267 (N_6267,N_6209,N_6136);
nor U6268 (N_6268,N_6090,N_6215);
nor U6269 (N_6269,N_6125,N_6192);
nand U6270 (N_6270,N_6154,N_6140);
xnor U6271 (N_6271,N_6211,N_6128);
and U6272 (N_6272,N_6199,N_6126);
nand U6273 (N_6273,N_6193,N_6221);
xnor U6274 (N_6274,N_6205,N_6174);
nand U6275 (N_6275,N_6119,N_6153);
and U6276 (N_6276,N_6187,N_6149);
and U6277 (N_6277,N_6151,N_6115);
nand U6278 (N_6278,N_6217,N_6117);
nand U6279 (N_6279,N_6147,N_6204);
nand U6280 (N_6280,N_6091,N_6213);
and U6281 (N_6281,N_6165,N_6141);
or U6282 (N_6282,N_6198,N_6168);
nor U6283 (N_6283,N_6088,N_6207);
and U6284 (N_6284,N_6226,N_6112);
and U6285 (N_6285,N_6152,N_6104);
or U6286 (N_6286,N_6208,N_6224);
nor U6287 (N_6287,N_6131,N_6176);
nand U6288 (N_6288,N_6184,N_6145);
nor U6289 (N_6289,N_6107,N_6127);
xor U6290 (N_6290,N_6144,N_6175);
nand U6291 (N_6291,N_6220,N_6194);
nor U6292 (N_6292,N_6085,N_6173);
xor U6293 (N_6293,N_6233,N_6172);
nor U6294 (N_6294,N_6162,N_6212);
and U6295 (N_6295,N_6185,N_6166);
and U6296 (N_6296,N_6216,N_6118);
or U6297 (N_6297,N_6191,N_6097);
nand U6298 (N_6298,N_6096,N_6210);
nor U6299 (N_6299,N_6089,N_6203);
nand U6300 (N_6300,N_6235,N_6182);
nor U6301 (N_6301,N_6100,N_6124);
nor U6302 (N_6302,N_6120,N_6219);
or U6303 (N_6303,N_6098,N_6196);
nor U6304 (N_6304,N_6133,N_6190);
xnor U6305 (N_6305,N_6227,N_6181);
nand U6306 (N_6306,N_6155,N_6129);
and U6307 (N_6307,N_6214,N_6106);
and U6308 (N_6308,N_6201,N_6206);
or U6309 (N_6309,N_6183,N_6197);
or U6310 (N_6310,N_6123,N_6099);
nor U6311 (N_6311,N_6231,N_6170);
xnor U6312 (N_6312,N_6083,N_6116);
nor U6313 (N_6313,N_6113,N_6189);
xnor U6314 (N_6314,N_6095,N_6130);
nand U6315 (N_6315,N_6122,N_6135);
nor U6316 (N_6316,N_6171,N_6148);
nor U6317 (N_6317,N_6228,N_6146);
xnor U6318 (N_6318,N_6134,N_6169);
xor U6319 (N_6319,N_6157,N_6156);
nand U6320 (N_6320,N_6225,N_6110);
nor U6321 (N_6321,N_6160,N_6214);
nand U6322 (N_6322,N_6128,N_6155);
xor U6323 (N_6323,N_6096,N_6186);
nand U6324 (N_6324,N_6094,N_6226);
nand U6325 (N_6325,N_6149,N_6180);
xnor U6326 (N_6326,N_6217,N_6197);
or U6327 (N_6327,N_6116,N_6143);
xnor U6328 (N_6328,N_6128,N_6159);
nand U6329 (N_6329,N_6097,N_6128);
xor U6330 (N_6330,N_6111,N_6213);
and U6331 (N_6331,N_6103,N_6156);
nor U6332 (N_6332,N_6148,N_6135);
and U6333 (N_6333,N_6113,N_6194);
nand U6334 (N_6334,N_6172,N_6227);
xnor U6335 (N_6335,N_6217,N_6196);
nand U6336 (N_6336,N_6213,N_6219);
or U6337 (N_6337,N_6172,N_6139);
nand U6338 (N_6338,N_6141,N_6231);
nand U6339 (N_6339,N_6193,N_6236);
or U6340 (N_6340,N_6161,N_6152);
xor U6341 (N_6341,N_6152,N_6126);
and U6342 (N_6342,N_6230,N_6228);
and U6343 (N_6343,N_6200,N_6127);
xor U6344 (N_6344,N_6081,N_6221);
nand U6345 (N_6345,N_6169,N_6235);
and U6346 (N_6346,N_6213,N_6081);
and U6347 (N_6347,N_6207,N_6094);
nand U6348 (N_6348,N_6084,N_6164);
and U6349 (N_6349,N_6210,N_6208);
and U6350 (N_6350,N_6215,N_6140);
and U6351 (N_6351,N_6157,N_6098);
nor U6352 (N_6352,N_6088,N_6181);
xor U6353 (N_6353,N_6085,N_6174);
or U6354 (N_6354,N_6185,N_6109);
xor U6355 (N_6355,N_6160,N_6221);
and U6356 (N_6356,N_6113,N_6105);
and U6357 (N_6357,N_6183,N_6139);
or U6358 (N_6358,N_6102,N_6162);
nand U6359 (N_6359,N_6091,N_6096);
and U6360 (N_6360,N_6211,N_6150);
nand U6361 (N_6361,N_6233,N_6236);
nor U6362 (N_6362,N_6214,N_6221);
xor U6363 (N_6363,N_6212,N_6099);
and U6364 (N_6364,N_6216,N_6222);
or U6365 (N_6365,N_6216,N_6207);
xor U6366 (N_6366,N_6193,N_6163);
or U6367 (N_6367,N_6192,N_6104);
nor U6368 (N_6368,N_6231,N_6146);
nor U6369 (N_6369,N_6102,N_6180);
or U6370 (N_6370,N_6118,N_6211);
and U6371 (N_6371,N_6111,N_6102);
nor U6372 (N_6372,N_6151,N_6190);
and U6373 (N_6373,N_6138,N_6101);
and U6374 (N_6374,N_6098,N_6143);
xor U6375 (N_6375,N_6230,N_6166);
xor U6376 (N_6376,N_6152,N_6143);
xnor U6377 (N_6377,N_6209,N_6172);
nor U6378 (N_6378,N_6209,N_6164);
xnor U6379 (N_6379,N_6153,N_6139);
and U6380 (N_6380,N_6171,N_6131);
nand U6381 (N_6381,N_6167,N_6086);
xor U6382 (N_6382,N_6154,N_6202);
nand U6383 (N_6383,N_6090,N_6107);
xnor U6384 (N_6384,N_6092,N_6087);
nand U6385 (N_6385,N_6138,N_6202);
or U6386 (N_6386,N_6218,N_6208);
or U6387 (N_6387,N_6144,N_6155);
and U6388 (N_6388,N_6133,N_6165);
xor U6389 (N_6389,N_6107,N_6126);
nand U6390 (N_6390,N_6099,N_6135);
xnor U6391 (N_6391,N_6096,N_6232);
nand U6392 (N_6392,N_6127,N_6082);
or U6393 (N_6393,N_6093,N_6225);
nor U6394 (N_6394,N_6095,N_6153);
and U6395 (N_6395,N_6172,N_6151);
nor U6396 (N_6396,N_6098,N_6183);
and U6397 (N_6397,N_6142,N_6145);
xor U6398 (N_6398,N_6192,N_6187);
nor U6399 (N_6399,N_6211,N_6103);
nand U6400 (N_6400,N_6274,N_6341);
and U6401 (N_6401,N_6323,N_6294);
nor U6402 (N_6402,N_6365,N_6279);
nand U6403 (N_6403,N_6361,N_6321);
nand U6404 (N_6404,N_6395,N_6267);
xnor U6405 (N_6405,N_6270,N_6307);
nand U6406 (N_6406,N_6326,N_6310);
xor U6407 (N_6407,N_6278,N_6355);
xor U6408 (N_6408,N_6277,N_6344);
nand U6409 (N_6409,N_6373,N_6370);
or U6410 (N_6410,N_6347,N_6346);
xnor U6411 (N_6411,N_6319,N_6249);
and U6412 (N_6412,N_6322,N_6324);
and U6413 (N_6413,N_6283,N_6259);
xnor U6414 (N_6414,N_6245,N_6396);
nand U6415 (N_6415,N_6386,N_6246);
and U6416 (N_6416,N_6271,N_6254);
or U6417 (N_6417,N_6250,N_6362);
xnor U6418 (N_6418,N_6394,N_6398);
and U6419 (N_6419,N_6262,N_6363);
or U6420 (N_6420,N_6350,N_6313);
and U6421 (N_6421,N_6291,N_6334);
xor U6422 (N_6422,N_6389,N_6377);
and U6423 (N_6423,N_6305,N_6316);
nand U6424 (N_6424,N_6337,N_6383);
nor U6425 (N_6425,N_6295,N_6338);
nand U6426 (N_6426,N_6301,N_6296);
xnor U6427 (N_6427,N_6351,N_6364);
or U6428 (N_6428,N_6331,N_6314);
nor U6429 (N_6429,N_6397,N_6317);
or U6430 (N_6430,N_6357,N_6261);
xnor U6431 (N_6431,N_6244,N_6292);
xor U6432 (N_6432,N_6308,N_6276);
xnor U6433 (N_6433,N_6382,N_6304);
or U6434 (N_6434,N_6315,N_6309);
or U6435 (N_6435,N_6359,N_6286);
and U6436 (N_6436,N_6285,N_6349);
xnor U6437 (N_6437,N_6339,N_6393);
or U6438 (N_6438,N_6311,N_6248);
nor U6439 (N_6439,N_6312,N_6293);
nor U6440 (N_6440,N_6329,N_6273);
or U6441 (N_6441,N_6330,N_6390);
nand U6442 (N_6442,N_6269,N_6399);
nor U6443 (N_6443,N_6384,N_6348);
nand U6444 (N_6444,N_6353,N_6258);
xnor U6445 (N_6445,N_6372,N_6297);
xnor U6446 (N_6446,N_6251,N_6318);
and U6447 (N_6447,N_6268,N_6240);
nor U6448 (N_6448,N_6257,N_6352);
nand U6449 (N_6449,N_6289,N_6281);
nand U6450 (N_6450,N_6366,N_6381);
nor U6451 (N_6451,N_6253,N_6241);
nand U6452 (N_6452,N_6306,N_6299);
nand U6453 (N_6453,N_6335,N_6284);
nor U6454 (N_6454,N_6320,N_6298);
or U6455 (N_6455,N_6303,N_6392);
or U6456 (N_6456,N_6252,N_6367);
and U6457 (N_6457,N_6247,N_6354);
xor U6458 (N_6458,N_6391,N_6255);
xor U6459 (N_6459,N_6345,N_6336);
and U6460 (N_6460,N_6376,N_6327);
nand U6461 (N_6461,N_6256,N_6243);
xor U6462 (N_6462,N_6290,N_6340);
xnor U6463 (N_6463,N_6374,N_6265);
xnor U6464 (N_6464,N_6282,N_6280);
nand U6465 (N_6465,N_6288,N_6369);
nand U6466 (N_6466,N_6358,N_6356);
and U6467 (N_6467,N_6371,N_6360);
xor U6468 (N_6468,N_6333,N_6328);
nor U6469 (N_6469,N_6332,N_6264);
nand U6470 (N_6470,N_6368,N_6385);
xor U6471 (N_6471,N_6387,N_6380);
or U6472 (N_6472,N_6266,N_6325);
and U6473 (N_6473,N_6378,N_6343);
or U6474 (N_6474,N_6302,N_6275);
and U6475 (N_6475,N_6388,N_6287);
xnor U6476 (N_6476,N_6242,N_6375);
and U6477 (N_6477,N_6260,N_6342);
nor U6478 (N_6478,N_6272,N_6263);
and U6479 (N_6479,N_6300,N_6379);
or U6480 (N_6480,N_6269,N_6311);
nand U6481 (N_6481,N_6335,N_6365);
or U6482 (N_6482,N_6317,N_6292);
and U6483 (N_6483,N_6355,N_6399);
and U6484 (N_6484,N_6355,N_6373);
or U6485 (N_6485,N_6263,N_6291);
xor U6486 (N_6486,N_6323,N_6302);
nor U6487 (N_6487,N_6279,N_6374);
xnor U6488 (N_6488,N_6302,N_6385);
nor U6489 (N_6489,N_6316,N_6254);
nor U6490 (N_6490,N_6368,N_6342);
nor U6491 (N_6491,N_6255,N_6339);
and U6492 (N_6492,N_6337,N_6297);
nor U6493 (N_6493,N_6396,N_6249);
xor U6494 (N_6494,N_6303,N_6273);
and U6495 (N_6495,N_6287,N_6350);
or U6496 (N_6496,N_6371,N_6252);
and U6497 (N_6497,N_6299,N_6343);
nor U6498 (N_6498,N_6392,N_6338);
and U6499 (N_6499,N_6275,N_6341);
and U6500 (N_6500,N_6304,N_6245);
or U6501 (N_6501,N_6386,N_6376);
xor U6502 (N_6502,N_6286,N_6303);
nand U6503 (N_6503,N_6245,N_6251);
and U6504 (N_6504,N_6362,N_6344);
and U6505 (N_6505,N_6356,N_6279);
and U6506 (N_6506,N_6346,N_6398);
and U6507 (N_6507,N_6342,N_6298);
nand U6508 (N_6508,N_6359,N_6264);
nor U6509 (N_6509,N_6398,N_6306);
xnor U6510 (N_6510,N_6329,N_6344);
xor U6511 (N_6511,N_6342,N_6370);
nor U6512 (N_6512,N_6307,N_6361);
nor U6513 (N_6513,N_6381,N_6292);
nand U6514 (N_6514,N_6363,N_6289);
nand U6515 (N_6515,N_6387,N_6301);
nand U6516 (N_6516,N_6340,N_6335);
nand U6517 (N_6517,N_6281,N_6345);
nand U6518 (N_6518,N_6270,N_6335);
xnor U6519 (N_6519,N_6352,N_6281);
or U6520 (N_6520,N_6252,N_6274);
xnor U6521 (N_6521,N_6309,N_6304);
xor U6522 (N_6522,N_6377,N_6309);
and U6523 (N_6523,N_6318,N_6267);
nor U6524 (N_6524,N_6280,N_6371);
nor U6525 (N_6525,N_6242,N_6324);
nor U6526 (N_6526,N_6344,N_6242);
or U6527 (N_6527,N_6263,N_6298);
or U6528 (N_6528,N_6277,N_6309);
or U6529 (N_6529,N_6390,N_6263);
or U6530 (N_6530,N_6362,N_6369);
xnor U6531 (N_6531,N_6367,N_6303);
or U6532 (N_6532,N_6295,N_6299);
xnor U6533 (N_6533,N_6248,N_6244);
and U6534 (N_6534,N_6397,N_6341);
nor U6535 (N_6535,N_6385,N_6255);
and U6536 (N_6536,N_6241,N_6340);
nand U6537 (N_6537,N_6368,N_6348);
xor U6538 (N_6538,N_6302,N_6387);
nor U6539 (N_6539,N_6341,N_6242);
and U6540 (N_6540,N_6326,N_6247);
or U6541 (N_6541,N_6255,N_6302);
and U6542 (N_6542,N_6293,N_6314);
nand U6543 (N_6543,N_6311,N_6274);
or U6544 (N_6544,N_6373,N_6245);
and U6545 (N_6545,N_6263,N_6249);
or U6546 (N_6546,N_6341,N_6349);
xnor U6547 (N_6547,N_6262,N_6326);
and U6548 (N_6548,N_6270,N_6244);
nand U6549 (N_6549,N_6309,N_6245);
and U6550 (N_6550,N_6305,N_6332);
nand U6551 (N_6551,N_6336,N_6303);
nand U6552 (N_6552,N_6265,N_6305);
xor U6553 (N_6553,N_6332,N_6379);
nand U6554 (N_6554,N_6283,N_6290);
and U6555 (N_6555,N_6347,N_6373);
nand U6556 (N_6556,N_6256,N_6359);
and U6557 (N_6557,N_6283,N_6385);
nand U6558 (N_6558,N_6247,N_6391);
nor U6559 (N_6559,N_6298,N_6274);
nand U6560 (N_6560,N_6439,N_6438);
and U6561 (N_6561,N_6464,N_6462);
nor U6562 (N_6562,N_6523,N_6444);
or U6563 (N_6563,N_6432,N_6553);
or U6564 (N_6564,N_6440,N_6416);
and U6565 (N_6565,N_6431,N_6518);
nand U6566 (N_6566,N_6470,N_6516);
nor U6567 (N_6567,N_6459,N_6488);
and U6568 (N_6568,N_6451,N_6538);
or U6569 (N_6569,N_6456,N_6517);
or U6570 (N_6570,N_6504,N_6535);
nor U6571 (N_6571,N_6450,N_6507);
xor U6572 (N_6572,N_6437,N_6486);
xor U6573 (N_6573,N_6403,N_6497);
nand U6574 (N_6574,N_6469,N_6474);
nand U6575 (N_6575,N_6402,N_6467);
and U6576 (N_6576,N_6480,N_6545);
xor U6577 (N_6577,N_6550,N_6530);
nor U6578 (N_6578,N_6543,N_6490);
and U6579 (N_6579,N_6420,N_6412);
nand U6580 (N_6580,N_6410,N_6554);
nor U6581 (N_6581,N_6520,N_6427);
and U6582 (N_6582,N_6465,N_6401);
and U6583 (N_6583,N_6468,N_6510);
or U6584 (N_6584,N_6505,N_6524);
nor U6585 (N_6585,N_6548,N_6455);
and U6586 (N_6586,N_6429,N_6483);
or U6587 (N_6587,N_6508,N_6559);
xor U6588 (N_6588,N_6471,N_6442);
xor U6589 (N_6589,N_6526,N_6428);
and U6590 (N_6590,N_6430,N_6532);
or U6591 (N_6591,N_6421,N_6415);
nand U6592 (N_6592,N_6503,N_6542);
or U6593 (N_6593,N_6514,N_6547);
and U6594 (N_6594,N_6413,N_6552);
nor U6595 (N_6595,N_6556,N_6527);
or U6596 (N_6596,N_6452,N_6400);
or U6597 (N_6597,N_6414,N_6434);
and U6598 (N_6598,N_6458,N_6534);
and U6599 (N_6599,N_6519,N_6478);
and U6600 (N_6600,N_6502,N_6436);
nor U6601 (N_6601,N_6453,N_6512);
or U6602 (N_6602,N_6493,N_6406);
nand U6603 (N_6603,N_6522,N_6536);
nor U6604 (N_6604,N_6485,N_6419);
and U6605 (N_6605,N_6558,N_6487);
and U6606 (N_6606,N_6506,N_6418);
or U6607 (N_6607,N_6555,N_6475);
nand U6608 (N_6608,N_6491,N_6495);
and U6609 (N_6609,N_6484,N_6433);
nor U6610 (N_6610,N_6501,N_6481);
nor U6611 (N_6611,N_6482,N_6435);
nor U6612 (N_6612,N_6407,N_6533);
or U6613 (N_6613,N_6411,N_6509);
xnor U6614 (N_6614,N_6551,N_6405);
xor U6615 (N_6615,N_6441,N_6494);
and U6616 (N_6616,N_6546,N_6425);
xnor U6617 (N_6617,N_6539,N_6423);
and U6618 (N_6618,N_6417,N_6472);
or U6619 (N_6619,N_6409,N_6498);
nand U6620 (N_6620,N_6422,N_6511);
nand U6621 (N_6621,N_6489,N_6557);
nand U6622 (N_6622,N_6492,N_6499);
or U6623 (N_6623,N_6513,N_6457);
xnor U6624 (N_6624,N_6528,N_6424);
nor U6625 (N_6625,N_6549,N_6473);
and U6626 (N_6626,N_6426,N_6477);
and U6627 (N_6627,N_6531,N_6476);
and U6628 (N_6628,N_6540,N_6408);
or U6629 (N_6629,N_6446,N_6529);
xor U6630 (N_6630,N_6445,N_6454);
and U6631 (N_6631,N_6443,N_6544);
or U6632 (N_6632,N_6479,N_6541);
nand U6633 (N_6633,N_6463,N_6500);
xor U6634 (N_6634,N_6460,N_6515);
nor U6635 (N_6635,N_6525,N_6449);
or U6636 (N_6636,N_6461,N_6466);
nand U6637 (N_6637,N_6496,N_6447);
xnor U6638 (N_6638,N_6448,N_6521);
and U6639 (N_6639,N_6404,N_6537);
and U6640 (N_6640,N_6487,N_6557);
nand U6641 (N_6641,N_6445,N_6495);
xnor U6642 (N_6642,N_6436,N_6555);
or U6643 (N_6643,N_6461,N_6536);
or U6644 (N_6644,N_6440,N_6473);
xor U6645 (N_6645,N_6460,N_6419);
and U6646 (N_6646,N_6492,N_6510);
nand U6647 (N_6647,N_6530,N_6545);
and U6648 (N_6648,N_6410,N_6489);
nor U6649 (N_6649,N_6472,N_6527);
xor U6650 (N_6650,N_6464,N_6477);
nor U6651 (N_6651,N_6525,N_6464);
and U6652 (N_6652,N_6538,N_6483);
nand U6653 (N_6653,N_6465,N_6487);
and U6654 (N_6654,N_6514,N_6538);
and U6655 (N_6655,N_6486,N_6407);
and U6656 (N_6656,N_6418,N_6492);
xnor U6657 (N_6657,N_6490,N_6466);
or U6658 (N_6658,N_6413,N_6497);
and U6659 (N_6659,N_6537,N_6465);
or U6660 (N_6660,N_6492,N_6456);
and U6661 (N_6661,N_6549,N_6556);
or U6662 (N_6662,N_6451,N_6434);
nand U6663 (N_6663,N_6426,N_6454);
nand U6664 (N_6664,N_6443,N_6428);
or U6665 (N_6665,N_6536,N_6496);
or U6666 (N_6666,N_6510,N_6437);
or U6667 (N_6667,N_6449,N_6517);
and U6668 (N_6668,N_6522,N_6487);
nor U6669 (N_6669,N_6492,N_6554);
xnor U6670 (N_6670,N_6493,N_6498);
nor U6671 (N_6671,N_6498,N_6408);
and U6672 (N_6672,N_6480,N_6504);
nand U6673 (N_6673,N_6460,N_6434);
or U6674 (N_6674,N_6497,N_6453);
xor U6675 (N_6675,N_6439,N_6413);
nor U6676 (N_6676,N_6480,N_6493);
or U6677 (N_6677,N_6542,N_6477);
or U6678 (N_6678,N_6490,N_6401);
nor U6679 (N_6679,N_6462,N_6552);
nor U6680 (N_6680,N_6456,N_6536);
xnor U6681 (N_6681,N_6557,N_6411);
nor U6682 (N_6682,N_6460,N_6556);
xor U6683 (N_6683,N_6485,N_6530);
xnor U6684 (N_6684,N_6402,N_6520);
nor U6685 (N_6685,N_6400,N_6503);
nor U6686 (N_6686,N_6488,N_6509);
and U6687 (N_6687,N_6530,N_6539);
and U6688 (N_6688,N_6513,N_6532);
and U6689 (N_6689,N_6501,N_6496);
or U6690 (N_6690,N_6428,N_6493);
nand U6691 (N_6691,N_6415,N_6449);
and U6692 (N_6692,N_6469,N_6448);
nor U6693 (N_6693,N_6431,N_6493);
nand U6694 (N_6694,N_6465,N_6540);
nand U6695 (N_6695,N_6427,N_6430);
nor U6696 (N_6696,N_6488,N_6427);
xor U6697 (N_6697,N_6489,N_6434);
nand U6698 (N_6698,N_6535,N_6527);
xnor U6699 (N_6699,N_6543,N_6461);
nor U6700 (N_6700,N_6489,N_6536);
nor U6701 (N_6701,N_6430,N_6536);
or U6702 (N_6702,N_6453,N_6504);
and U6703 (N_6703,N_6400,N_6429);
and U6704 (N_6704,N_6483,N_6460);
and U6705 (N_6705,N_6497,N_6433);
nor U6706 (N_6706,N_6451,N_6414);
or U6707 (N_6707,N_6447,N_6418);
xor U6708 (N_6708,N_6521,N_6531);
xnor U6709 (N_6709,N_6502,N_6531);
xnor U6710 (N_6710,N_6510,N_6457);
nand U6711 (N_6711,N_6533,N_6541);
nor U6712 (N_6712,N_6556,N_6416);
or U6713 (N_6713,N_6447,N_6409);
xor U6714 (N_6714,N_6501,N_6528);
or U6715 (N_6715,N_6535,N_6406);
or U6716 (N_6716,N_6487,N_6486);
xnor U6717 (N_6717,N_6471,N_6463);
or U6718 (N_6718,N_6404,N_6416);
xnor U6719 (N_6719,N_6493,N_6411);
nand U6720 (N_6720,N_6696,N_6568);
and U6721 (N_6721,N_6575,N_6679);
nor U6722 (N_6722,N_6580,N_6606);
xor U6723 (N_6723,N_6626,N_6682);
nor U6724 (N_6724,N_6708,N_6663);
nand U6725 (N_6725,N_6608,N_6706);
nor U6726 (N_6726,N_6586,N_6590);
xor U6727 (N_6727,N_6685,N_6659);
xor U6728 (N_6728,N_6646,N_6704);
and U6729 (N_6729,N_6584,N_6700);
xnor U6730 (N_6730,N_6617,N_6604);
and U6731 (N_6731,N_6598,N_6565);
nand U6732 (N_6732,N_6619,N_6623);
nand U6733 (N_6733,N_6688,N_6607);
xnor U6734 (N_6734,N_6703,N_6637);
nand U6735 (N_6735,N_6643,N_6578);
nor U6736 (N_6736,N_6636,N_6667);
nor U6737 (N_6737,N_6563,N_6600);
nand U6738 (N_6738,N_6594,N_6573);
xnor U6739 (N_6739,N_6595,N_6647);
nor U6740 (N_6740,N_6585,N_6673);
and U6741 (N_6741,N_6615,N_6694);
xnor U6742 (N_6742,N_6672,N_6639);
and U6743 (N_6743,N_6664,N_6645);
or U6744 (N_6744,N_6632,N_6709);
nand U6745 (N_6745,N_6705,N_6707);
or U6746 (N_6746,N_6649,N_6641);
and U6747 (N_6747,N_6596,N_6668);
xor U6748 (N_6748,N_6669,N_6711);
nand U6749 (N_6749,N_6652,N_6622);
nand U6750 (N_6750,N_6574,N_6640);
xnor U6751 (N_6751,N_6648,N_6631);
nor U6752 (N_6752,N_6650,N_6658);
nor U6753 (N_6753,N_6665,N_6634);
nand U6754 (N_6754,N_6592,N_6644);
and U6755 (N_6755,N_6689,N_6671);
and U6756 (N_6756,N_6597,N_6674);
or U6757 (N_6757,N_6691,N_6569);
or U6758 (N_6758,N_6562,N_6625);
and U6759 (N_6759,N_6666,N_6603);
xor U6760 (N_6760,N_6630,N_6702);
nor U6761 (N_6761,N_6662,N_6642);
xor U6762 (N_6762,N_6602,N_6692);
nand U6763 (N_6763,N_6616,N_6571);
nand U6764 (N_6764,N_6716,N_6589);
nor U6765 (N_6765,N_6621,N_6693);
nor U6766 (N_6766,N_6567,N_6718);
and U6767 (N_6767,N_6654,N_6628);
nand U6768 (N_6768,N_6588,N_6561);
or U6769 (N_6769,N_6629,N_6612);
nand U6770 (N_6770,N_6697,N_6564);
and U6771 (N_6771,N_6614,N_6678);
xnor U6772 (N_6772,N_6638,N_6591);
nor U6773 (N_6773,N_6566,N_6599);
nand U6774 (N_6774,N_6583,N_6613);
nand U6775 (N_6775,N_6587,N_6593);
nor U6776 (N_6776,N_6605,N_6611);
nor U6777 (N_6777,N_6684,N_6698);
and U6778 (N_6778,N_6635,N_6676);
nand U6779 (N_6779,N_6633,N_6717);
nand U6780 (N_6780,N_6695,N_6627);
nand U6781 (N_6781,N_6719,N_6582);
nor U6782 (N_6782,N_6714,N_6655);
nand U6783 (N_6783,N_6601,N_6656);
xnor U6784 (N_6784,N_6651,N_6570);
xnor U6785 (N_6785,N_6710,N_6675);
nor U6786 (N_6786,N_6657,N_6699);
nor U6787 (N_6787,N_6610,N_6712);
xnor U6788 (N_6788,N_6581,N_6572);
nor U6789 (N_6789,N_6577,N_6618);
and U6790 (N_6790,N_6560,N_6620);
xnor U6791 (N_6791,N_6690,N_6579);
or U6792 (N_6792,N_6686,N_6660);
nor U6793 (N_6793,N_6661,N_6576);
and U6794 (N_6794,N_6701,N_6609);
nor U6795 (N_6795,N_6670,N_6677);
nor U6796 (N_6796,N_6681,N_6624);
xor U6797 (N_6797,N_6715,N_6680);
or U6798 (N_6798,N_6687,N_6713);
xnor U6799 (N_6799,N_6683,N_6653);
xor U6800 (N_6800,N_6561,N_6703);
nor U6801 (N_6801,N_6626,N_6627);
xnor U6802 (N_6802,N_6567,N_6600);
and U6803 (N_6803,N_6655,N_6717);
nor U6804 (N_6804,N_6596,N_6677);
xnor U6805 (N_6805,N_6601,N_6706);
nor U6806 (N_6806,N_6610,N_6710);
nor U6807 (N_6807,N_6606,N_6646);
and U6808 (N_6808,N_6717,N_6561);
and U6809 (N_6809,N_6669,N_6648);
or U6810 (N_6810,N_6599,N_6664);
xor U6811 (N_6811,N_6636,N_6686);
nand U6812 (N_6812,N_6629,N_6718);
xor U6813 (N_6813,N_6567,N_6667);
nand U6814 (N_6814,N_6715,N_6574);
xor U6815 (N_6815,N_6697,N_6592);
xnor U6816 (N_6816,N_6714,N_6648);
and U6817 (N_6817,N_6686,N_6622);
nor U6818 (N_6818,N_6642,N_6699);
and U6819 (N_6819,N_6592,N_6700);
nand U6820 (N_6820,N_6644,N_6662);
or U6821 (N_6821,N_6561,N_6670);
nand U6822 (N_6822,N_6567,N_6618);
or U6823 (N_6823,N_6604,N_6625);
nor U6824 (N_6824,N_6573,N_6563);
and U6825 (N_6825,N_6673,N_6589);
nand U6826 (N_6826,N_6620,N_6640);
and U6827 (N_6827,N_6646,N_6592);
or U6828 (N_6828,N_6581,N_6603);
or U6829 (N_6829,N_6628,N_6563);
nor U6830 (N_6830,N_6659,N_6623);
nand U6831 (N_6831,N_6719,N_6607);
xor U6832 (N_6832,N_6700,N_6637);
xnor U6833 (N_6833,N_6578,N_6689);
or U6834 (N_6834,N_6621,N_6704);
xnor U6835 (N_6835,N_6684,N_6712);
or U6836 (N_6836,N_6591,N_6612);
nand U6837 (N_6837,N_6686,N_6719);
nor U6838 (N_6838,N_6672,N_6604);
nor U6839 (N_6839,N_6584,N_6639);
and U6840 (N_6840,N_6669,N_6619);
xor U6841 (N_6841,N_6578,N_6640);
or U6842 (N_6842,N_6593,N_6648);
or U6843 (N_6843,N_6573,N_6644);
nor U6844 (N_6844,N_6702,N_6704);
xor U6845 (N_6845,N_6577,N_6582);
xnor U6846 (N_6846,N_6624,N_6567);
and U6847 (N_6847,N_6692,N_6607);
nand U6848 (N_6848,N_6672,N_6575);
nor U6849 (N_6849,N_6679,N_6717);
or U6850 (N_6850,N_6715,N_6665);
and U6851 (N_6851,N_6671,N_6612);
or U6852 (N_6852,N_6638,N_6708);
nor U6853 (N_6853,N_6653,N_6624);
xor U6854 (N_6854,N_6617,N_6670);
and U6855 (N_6855,N_6713,N_6598);
xor U6856 (N_6856,N_6685,N_6628);
and U6857 (N_6857,N_6619,N_6632);
or U6858 (N_6858,N_6606,N_6590);
nand U6859 (N_6859,N_6711,N_6667);
or U6860 (N_6860,N_6718,N_6612);
xor U6861 (N_6861,N_6636,N_6631);
nor U6862 (N_6862,N_6715,N_6578);
nand U6863 (N_6863,N_6651,N_6617);
or U6864 (N_6864,N_6569,N_6662);
xor U6865 (N_6865,N_6580,N_6687);
or U6866 (N_6866,N_6646,N_6631);
nand U6867 (N_6867,N_6680,N_6706);
and U6868 (N_6868,N_6571,N_6654);
nor U6869 (N_6869,N_6693,N_6657);
or U6870 (N_6870,N_6650,N_6579);
xnor U6871 (N_6871,N_6622,N_6693);
or U6872 (N_6872,N_6564,N_6583);
xnor U6873 (N_6873,N_6604,N_6684);
nor U6874 (N_6874,N_6663,N_6653);
and U6875 (N_6875,N_6703,N_6602);
nand U6876 (N_6876,N_6682,N_6619);
or U6877 (N_6877,N_6639,N_6649);
xnor U6878 (N_6878,N_6647,N_6609);
or U6879 (N_6879,N_6598,N_6711);
nand U6880 (N_6880,N_6731,N_6795);
xnor U6881 (N_6881,N_6760,N_6878);
or U6882 (N_6882,N_6818,N_6733);
nand U6883 (N_6883,N_6817,N_6789);
nor U6884 (N_6884,N_6831,N_6721);
or U6885 (N_6885,N_6856,N_6737);
or U6886 (N_6886,N_6830,N_6876);
and U6887 (N_6887,N_6751,N_6873);
nand U6888 (N_6888,N_6759,N_6879);
nor U6889 (N_6889,N_6776,N_6812);
xnor U6890 (N_6890,N_6769,N_6848);
or U6891 (N_6891,N_6819,N_6868);
and U6892 (N_6892,N_6768,N_6858);
nand U6893 (N_6893,N_6826,N_6755);
or U6894 (N_6894,N_6854,N_6859);
xnor U6895 (N_6895,N_6862,N_6726);
or U6896 (N_6896,N_6798,N_6732);
xor U6897 (N_6897,N_6839,N_6774);
and U6898 (N_6898,N_6735,N_6727);
and U6899 (N_6899,N_6810,N_6829);
or U6900 (N_6900,N_6746,N_6779);
or U6901 (N_6901,N_6741,N_6750);
or U6902 (N_6902,N_6792,N_6842);
nand U6903 (N_6903,N_6794,N_6747);
nor U6904 (N_6904,N_6877,N_6742);
or U6905 (N_6905,N_6761,N_6806);
and U6906 (N_6906,N_6874,N_6745);
and U6907 (N_6907,N_6836,N_6824);
nor U6908 (N_6908,N_6837,N_6738);
nand U6909 (N_6909,N_6743,N_6823);
and U6910 (N_6910,N_6871,N_6853);
and U6911 (N_6911,N_6803,N_6875);
nand U6912 (N_6912,N_6857,N_6739);
or U6913 (N_6913,N_6787,N_6844);
nand U6914 (N_6914,N_6748,N_6749);
or U6915 (N_6915,N_6834,N_6763);
and U6916 (N_6916,N_6728,N_6822);
or U6917 (N_6917,N_6801,N_6722);
and U6918 (N_6918,N_6861,N_6797);
and U6919 (N_6919,N_6772,N_6734);
nand U6920 (N_6920,N_6838,N_6773);
and U6921 (N_6921,N_6814,N_6869);
or U6922 (N_6922,N_6821,N_6846);
xor U6923 (N_6923,N_6783,N_6725);
xor U6924 (N_6924,N_6793,N_6807);
or U6925 (N_6925,N_6833,N_6729);
and U6926 (N_6926,N_6802,N_6775);
nand U6927 (N_6927,N_6758,N_6799);
xor U6928 (N_6928,N_6840,N_6832);
and U6929 (N_6929,N_6860,N_6757);
nor U6930 (N_6930,N_6796,N_6762);
or U6931 (N_6931,N_6845,N_6850);
or U6932 (N_6932,N_6723,N_6847);
and U6933 (N_6933,N_6730,N_6804);
nor U6934 (N_6934,N_6791,N_6863);
and U6935 (N_6935,N_6867,N_6809);
and U6936 (N_6936,N_6865,N_6771);
xor U6937 (N_6937,N_6827,N_6744);
nand U6938 (N_6938,N_6870,N_6841);
xnor U6939 (N_6939,N_6816,N_6825);
and U6940 (N_6940,N_6753,N_6764);
nand U6941 (N_6941,N_6754,N_6784);
xor U6942 (N_6942,N_6756,N_6800);
and U6943 (N_6943,N_6820,N_6815);
xor U6944 (N_6944,N_6855,N_6786);
xnor U6945 (N_6945,N_6765,N_6766);
or U6946 (N_6946,N_6790,N_6752);
and U6947 (N_6947,N_6782,N_6780);
nor U6948 (N_6948,N_6720,N_6767);
or U6949 (N_6949,N_6843,N_6808);
xor U6950 (N_6950,N_6828,N_6851);
or U6951 (N_6951,N_6785,N_6788);
xor U6952 (N_6952,N_6852,N_6724);
or U6953 (N_6953,N_6813,N_6811);
and U6954 (N_6954,N_6835,N_6866);
nand U6955 (N_6955,N_6740,N_6849);
nand U6956 (N_6956,N_6864,N_6872);
and U6957 (N_6957,N_6778,N_6770);
and U6958 (N_6958,N_6736,N_6805);
nor U6959 (N_6959,N_6777,N_6781);
and U6960 (N_6960,N_6861,N_6820);
or U6961 (N_6961,N_6754,N_6739);
nand U6962 (N_6962,N_6789,N_6815);
and U6963 (N_6963,N_6745,N_6824);
nor U6964 (N_6964,N_6861,N_6799);
nor U6965 (N_6965,N_6739,N_6873);
nand U6966 (N_6966,N_6821,N_6760);
nand U6967 (N_6967,N_6874,N_6797);
and U6968 (N_6968,N_6762,N_6868);
nor U6969 (N_6969,N_6851,N_6804);
xnor U6970 (N_6970,N_6878,N_6819);
and U6971 (N_6971,N_6814,N_6771);
or U6972 (N_6972,N_6762,N_6841);
nand U6973 (N_6973,N_6754,N_6736);
nor U6974 (N_6974,N_6852,N_6842);
and U6975 (N_6975,N_6740,N_6731);
and U6976 (N_6976,N_6813,N_6755);
nor U6977 (N_6977,N_6859,N_6735);
and U6978 (N_6978,N_6764,N_6776);
or U6979 (N_6979,N_6796,N_6815);
xnor U6980 (N_6980,N_6836,N_6759);
and U6981 (N_6981,N_6862,N_6728);
nand U6982 (N_6982,N_6776,N_6847);
or U6983 (N_6983,N_6848,N_6730);
xor U6984 (N_6984,N_6806,N_6753);
or U6985 (N_6985,N_6751,N_6723);
or U6986 (N_6986,N_6749,N_6808);
and U6987 (N_6987,N_6766,N_6768);
nand U6988 (N_6988,N_6793,N_6849);
nand U6989 (N_6989,N_6807,N_6723);
nand U6990 (N_6990,N_6763,N_6871);
and U6991 (N_6991,N_6853,N_6840);
xnor U6992 (N_6992,N_6865,N_6731);
nand U6993 (N_6993,N_6876,N_6732);
xnor U6994 (N_6994,N_6792,N_6814);
or U6995 (N_6995,N_6751,N_6866);
and U6996 (N_6996,N_6738,N_6790);
or U6997 (N_6997,N_6828,N_6868);
nor U6998 (N_6998,N_6877,N_6802);
xor U6999 (N_6999,N_6821,N_6839);
nand U7000 (N_7000,N_6844,N_6793);
nand U7001 (N_7001,N_6875,N_6836);
or U7002 (N_7002,N_6760,N_6748);
xnor U7003 (N_7003,N_6722,N_6846);
nor U7004 (N_7004,N_6814,N_6756);
nor U7005 (N_7005,N_6833,N_6720);
nor U7006 (N_7006,N_6784,N_6874);
nor U7007 (N_7007,N_6805,N_6833);
nand U7008 (N_7008,N_6801,N_6805);
nand U7009 (N_7009,N_6720,N_6848);
xnor U7010 (N_7010,N_6853,N_6775);
nand U7011 (N_7011,N_6831,N_6761);
or U7012 (N_7012,N_6737,N_6785);
or U7013 (N_7013,N_6745,N_6791);
xor U7014 (N_7014,N_6842,N_6849);
nor U7015 (N_7015,N_6759,N_6775);
and U7016 (N_7016,N_6721,N_6741);
nor U7017 (N_7017,N_6876,N_6797);
nor U7018 (N_7018,N_6766,N_6730);
and U7019 (N_7019,N_6774,N_6877);
nor U7020 (N_7020,N_6766,N_6862);
nor U7021 (N_7021,N_6731,N_6804);
xor U7022 (N_7022,N_6819,N_6865);
nand U7023 (N_7023,N_6758,N_6817);
or U7024 (N_7024,N_6790,N_6817);
xnor U7025 (N_7025,N_6756,N_6745);
nor U7026 (N_7026,N_6820,N_6767);
and U7027 (N_7027,N_6768,N_6801);
and U7028 (N_7028,N_6808,N_6794);
or U7029 (N_7029,N_6743,N_6790);
xor U7030 (N_7030,N_6777,N_6729);
nand U7031 (N_7031,N_6739,N_6821);
nand U7032 (N_7032,N_6730,N_6729);
nand U7033 (N_7033,N_6727,N_6788);
xor U7034 (N_7034,N_6877,N_6729);
or U7035 (N_7035,N_6877,N_6728);
nand U7036 (N_7036,N_6769,N_6726);
nand U7037 (N_7037,N_6802,N_6742);
or U7038 (N_7038,N_6873,N_6769);
and U7039 (N_7039,N_6792,N_6727);
or U7040 (N_7040,N_7030,N_6895);
and U7041 (N_7041,N_6998,N_6996);
xor U7042 (N_7042,N_6961,N_7033);
nor U7043 (N_7043,N_6914,N_6956);
nor U7044 (N_7044,N_6966,N_7037);
and U7045 (N_7045,N_6893,N_6910);
nor U7046 (N_7046,N_6986,N_6968);
xor U7047 (N_7047,N_6937,N_6903);
nor U7048 (N_7048,N_7015,N_6987);
nand U7049 (N_7049,N_6926,N_6927);
and U7050 (N_7050,N_6942,N_6881);
nand U7051 (N_7051,N_6905,N_7000);
or U7052 (N_7052,N_6896,N_6899);
nand U7053 (N_7053,N_6975,N_6887);
nand U7054 (N_7054,N_6885,N_7021);
nand U7055 (N_7055,N_6939,N_6979);
or U7056 (N_7056,N_7032,N_6980);
xnor U7057 (N_7057,N_6969,N_6923);
nand U7058 (N_7058,N_6928,N_7002);
nand U7059 (N_7059,N_6891,N_6901);
nand U7060 (N_7060,N_6941,N_6906);
nor U7061 (N_7061,N_6944,N_7001);
nand U7062 (N_7062,N_6940,N_6988);
xor U7063 (N_7063,N_6915,N_7006);
nor U7064 (N_7064,N_6963,N_6938);
xor U7065 (N_7065,N_6889,N_6964);
xnor U7066 (N_7066,N_7008,N_6932);
nand U7067 (N_7067,N_7034,N_7023);
nor U7068 (N_7068,N_6947,N_6897);
and U7069 (N_7069,N_7026,N_6913);
nand U7070 (N_7070,N_6894,N_6970);
nand U7071 (N_7071,N_6892,N_6976);
nor U7072 (N_7072,N_7039,N_6908);
or U7073 (N_7073,N_7011,N_6972);
and U7074 (N_7074,N_6931,N_6990);
xor U7075 (N_7075,N_6922,N_6909);
xor U7076 (N_7076,N_7024,N_6957);
nand U7077 (N_7077,N_6958,N_6991);
or U7078 (N_7078,N_6904,N_6935);
xnor U7079 (N_7079,N_6898,N_6886);
nor U7080 (N_7080,N_6933,N_7016);
or U7081 (N_7081,N_7005,N_6978);
or U7082 (N_7082,N_6930,N_6982);
xnor U7083 (N_7083,N_7013,N_7019);
xor U7084 (N_7084,N_6993,N_6974);
or U7085 (N_7085,N_6967,N_6919);
xnor U7086 (N_7086,N_6981,N_6934);
nand U7087 (N_7087,N_6977,N_7007);
nand U7088 (N_7088,N_6948,N_6989);
nor U7089 (N_7089,N_7025,N_6920);
xor U7090 (N_7090,N_7027,N_6995);
or U7091 (N_7091,N_7022,N_6883);
and U7092 (N_7092,N_6882,N_6907);
and U7093 (N_7093,N_6997,N_6936);
nor U7094 (N_7094,N_6949,N_7003);
nor U7095 (N_7095,N_7012,N_7004);
nand U7096 (N_7096,N_6951,N_7028);
or U7097 (N_7097,N_6946,N_7031);
and U7098 (N_7098,N_7017,N_7029);
nand U7099 (N_7099,N_6912,N_6952);
nor U7100 (N_7100,N_6960,N_6924);
xnor U7101 (N_7101,N_6900,N_7014);
nand U7102 (N_7102,N_6965,N_7009);
nand U7103 (N_7103,N_6890,N_6925);
or U7104 (N_7104,N_7018,N_6959);
and U7105 (N_7105,N_6884,N_6950);
or U7106 (N_7106,N_7038,N_6902);
and U7107 (N_7107,N_6929,N_7020);
nor U7108 (N_7108,N_6973,N_6911);
nand U7109 (N_7109,N_6983,N_6953);
nor U7110 (N_7110,N_6921,N_6955);
nor U7111 (N_7111,N_6943,N_6962);
xnor U7112 (N_7112,N_6945,N_6984);
nand U7113 (N_7113,N_7010,N_6918);
and U7114 (N_7114,N_7035,N_6917);
nand U7115 (N_7115,N_6888,N_6916);
and U7116 (N_7116,N_6954,N_7036);
and U7117 (N_7117,N_6985,N_6994);
and U7118 (N_7118,N_6992,N_6999);
and U7119 (N_7119,N_6880,N_6971);
nor U7120 (N_7120,N_6997,N_7005);
nand U7121 (N_7121,N_6977,N_6915);
nand U7122 (N_7122,N_6911,N_6932);
and U7123 (N_7123,N_7033,N_7031);
xor U7124 (N_7124,N_6955,N_6881);
nand U7125 (N_7125,N_7012,N_6973);
or U7126 (N_7126,N_7033,N_6939);
nand U7127 (N_7127,N_6961,N_6914);
and U7128 (N_7128,N_6986,N_7018);
nand U7129 (N_7129,N_6978,N_6896);
nor U7130 (N_7130,N_6948,N_6917);
nor U7131 (N_7131,N_6921,N_6966);
nand U7132 (N_7132,N_6923,N_7018);
and U7133 (N_7133,N_6912,N_6920);
or U7134 (N_7134,N_6943,N_6952);
nor U7135 (N_7135,N_6897,N_7020);
nor U7136 (N_7136,N_6935,N_6970);
or U7137 (N_7137,N_6917,N_6906);
or U7138 (N_7138,N_6915,N_6931);
nand U7139 (N_7139,N_6963,N_6954);
and U7140 (N_7140,N_6957,N_6886);
nor U7141 (N_7141,N_7038,N_7008);
xnor U7142 (N_7142,N_6946,N_6958);
nand U7143 (N_7143,N_7023,N_7036);
or U7144 (N_7144,N_7038,N_6943);
nor U7145 (N_7145,N_6955,N_6901);
and U7146 (N_7146,N_6905,N_6949);
nor U7147 (N_7147,N_6997,N_6909);
xnor U7148 (N_7148,N_6956,N_7017);
or U7149 (N_7149,N_6990,N_6946);
nand U7150 (N_7150,N_6910,N_7025);
nor U7151 (N_7151,N_6946,N_7019);
and U7152 (N_7152,N_6893,N_6974);
and U7153 (N_7153,N_6963,N_7016);
and U7154 (N_7154,N_6944,N_6997);
nand U7155 (N_7155,N_7007,N_6943);
nand U7156 (N_7156,N_6913,N_6978);
nand U7157 (N_7157,N_7001,N_6926);
or U7158 (N_7158,N_6925,N_7014);
nor U7159 (N_7159,N_6946,N_6964);
or U7160 (N_7160,N_6951,N_6934);
xnor U7161 (N_7161,N_6930,N_6970);
nand U7162 (N_7162,N_6893,N_6993);
xnor U7163 (N_7163,N_6909,N_6923);
or U7164 (N_7164,N_7018,N_6960);
xnor U7165 (N_7165,N_6918,N_6928);
or U7166 (N_7166,N_7032,N_6945);
and U7167 (N_7167,N_6902,N_6880);
xnor U7168 (N_7168,N_6882,N_6949);
and U7169 (N_7169,N_6928,N_6972);
nand U7170 (N_7170,N_7022,N_6946);
xnor U7171 (N_7171,N_7024,N_6895);
and U7172 (N_7172,N_7022,N_6974);
and U7173 (N_7173,N_6951,N_7021);
nor U7174 (N_7174,N_6963,N_7019);
and U7175 (N_7175,N_6948,N_7015);
and U7176 (N_7176,N_6941,N_7039);
and U7177 (N_7177,N_6886,N_7009);
or U7178 (N_7178,N_7013,N_6917);
nand U7179 (N_7179,N_6991,N_6939);
or U7180 (N_7180,N_6957,N_7025);
nand U7181 (N_7181,N_6995,N_6902);
nor U7182 (N_7182,N_6951,N_6950);
nor U7183 (N_7183,N_7037,N_6953);
nor U7184 (N_7184,N_6896,N_6931);
nand U7185 (N_7185,N_6949,N_6934);
nand U7186 (N_7186,N_6900,N_6939);
nor U7187 (N_7187,N_6903,N_6880);
nor U7188 (N_7188,N_6920,N_6982);
or U7189 (N_7189,N_6920,N_6901);
nor U7190 (N_7190,N_6980,N_6887);
nand U7191 (N_7191,N_7029,N_6891);
or U7192 (N_7192,N_6981,N_6892);
xor U7193 (N_7193,N_6899,N_6932);
xnor U7194 (N_7194,N_6899,N_6950);
xor U7195 (N_7195,N_7014,N_6972);
or U7196 (N_7196,N_6924,N_6964);
or U7197 (N_7197,N_7039,N_7000);
xor U7198 (N_7198,N_6986,N_6912);
nand U7199 (N_7199,N_7014,N_6986);
xnor U7200 (N_7200,N_7165,N_7154);
and U7201 (N_7201,N_7122,N_7115);
xor U7202 (N_7202,N_7074,N_7175);
nor U7203 (N_7203,N_7054,N_7088);
xnor U7204 (N_7204,N_7105,N_7119);
or U7205 (N_7205,N_7049,N_7066);
xor U7206 (N_7206,N_7098,N_7104);
nand U7207 (N_7207,N_7082,N_7080);
and U7208 (N_7208,N_7161,N_7063);
nand U7209 (N_7209,N_7140,N_7092);
xor U7210 (N_7210,N_7136,N_7040);
nor U7211 (N_7211,N_7167,N_7148);
nor U7212 (N_7212,N_7060,N_7169);
or U7213 (N_7213,N_7101,N_7069);
and U7214 (N_7214,N_7135,N_7156);
or U7215 (N_7215,N_7193,N_7132);
and U7216 (N_7216,N_7149,N_7095);
nor U7217 (N_7217,N_7081,N_7164);
nand U7218 (N_7218,N_7199,N_7143);
xor U7219 (N_7219,N_7047,N_7113);
xor U7220 (N_7220,N_7152,N_7185);
nor U7221 (N_7221,N_7102,N_7171);
or U7222 (N_7222,N_7050,N_7051);
nand U7223 (N_7223,N_7068,N_7166);
xor U7224 (N_7224,N_7091,N_7116);
and U7225 (N_7225,N_7067,N_7173);
and U7226 (N_7226,N_7071,N_7055);
nand U7227 (N_7227,N_7198,N_7123);
or U7228 (N_7228,N_7073,N_7184);
or U7229 (N_7229,N_7182,N_7094);
nand U7230 (N_7230,N_7183,N_7174);
xnor U7231 (N_7231,N_7170,N_7137);
or U7232 (N_7232,N_7111,N_7042);
xnor U7233 (N_7233,N_7197,N_7053);
nand U7234 (N_7234,N_7126,N_7188);
and U7235 (N_7235,N_7044,N_7117);
and U7236 (N_7236,N_7172,N_7085);
or U7237 (N_7237,N_7138,N_7157);
or U7238 (N_7238,N_7190,N_7191);
nand U7239 (N_7239,N_7176,N_7045);
nor U7240 (N_7240,N_7083,N_7133);
nand U7241 (N_7241,N_7130,N_7192);
nor U7242 (N_7242,N_7155,N_7077);
nor U7243 (N_7243,N_7062,N_7180);
xnor U7244 (N_7244,N_7194,N_7056);
nand U7245 (N_7245,N_7162,N_7112);
nand U7246 (N_7246,N_7186,N_7159);
nand U7247 (N_7247,N_7084,N_7124);
xor U7248 (N_7248,N_7072,N_7127);
nor U7249 (N_7249,N_7163,N_7179);
nand U7250 (N_7250,N_7096,N_7103);
nand U7251 (N_7251,N_7189,N_7150);
xor U7252 (N_7252,N_7196,N_7187);
and U7253 (N_7253,N_7160,N_7086);
nor U7254 (N_7254,N_7118,N_7146);
or U7255 (N_7255,N_7079,N_7093);
and U7256 (N_7256,N_7070,N_7114);
and U7257 (N_7257,N_7046,N_7108);
xor U7258 (N_7258,N_7177,N_7087);
nor U7259 (N_7259,N_7052,N_7195);
or U7260 (N_7260,N_7097,N_7109);
nand U7261 (N_7261,N_7041,N_7128);
or U7262 (N_7262,N_7061,N_7059);
nand U7263 (N_7263,N_7106,N_7099);
nor U7264 (N_7264,N_7134,N_7043);
and U7265 (N_7265,N_7090,N_7153);
nand U7266 (N_7266,N_7168,N_7057);
xnor U7267 (N_7267,N_7075,N_7089);
and U7268 (N_7268,N_7141,N_7121);
and U7269 (N_7269,N_7058,N_7151);
or U7270 (N_7270,N_7139,N_7078);
and U7271 (N_7271,N_7145,N_7125);
and U7272 (N_7272,N_7131,N_7142);
or U7273 (N_7273,N_7147,N_7129);
xor U7274 (N_7274,N_7181,N_7144);
or U7275 (N_7275,N_7107,N_7048);
nor U7276 (N_7276,N_7158,N_7110);
xor U7277 (N_7277,N_7065,N_7120);
or U7278 (N_7278,N_7100,N_7076);
and U7279 (N_7279,N_7178,N_7064);
and U7280 (N_7280,N_7080,N_7184);
or U7281 (N_7281,N_7179,N_7050);
and U7282 (N_7282,N_7045,N_7145);
xor U7283 (N_7283,N_7177,N_7182);
and U7284 (N_7284,N_7177,N_7046);
nand U7285 (N_7285,N_7041,N_7110);
nor U7286 (N_7286,N_7171,N_7047);
nand U7287 (N_7287,N_7059,N_7091);
nor U7288 (N_7288,N_7095,N_7046);
or U7289 (N_7289,N_7079,N_7118);
or U7290 (N_7290,N_7108,N_7138);
or U7291 (N_7291,N_7188,N_7080);
or U7292 (N_7292,N_7043,N_7058);
or U7293 (N_7293,N_7124,N_7061);
nor U7294 (N_7294,N_7087,N_7047);
nand U7295 (N_7295,N_7162,N_7063);
nor U7296 (N_7296,N_7043,N_7189);
and U7297 (N_7297,N_7098,N_7120);
or U7298 (N_7298,N_7101,N_7108);
xnor U7299 (N_7299,N_7130,N_7125);
or U7300 (N_7300,N_7174,N_7061);
nand U7301 (N_7301,N_7114,N_7040);
and U7302 (N_7302,N_7170,N_7192);
xor U7303 (N_7303,N_7199,N_7053);
xnor U7304 (N_7304,N_7089,N_7054);
or U7305 (N_7305,N_7061,N_7163);
nand U7306 (N_7306,N_7196,N_7105);
xor U7307 (N_7307,N_7188,N_7147);
nor U7308 (N_7308,N_7041,N_7067);
nand U7309 (N_7309,N_7050,N_7094);
nor U7310 (N_7310,N_7145,N_7186);
and U7311 (N_7311,N_7192,N_7070);
xnor U7312 (N_7312,N_7105,N_7056);
nand U7313 (N_7313,N_7183,N_7130);
nand U7314 (N_7314,N_7143,N_7095);
and U7315 (N_7315,N_7127,N_7150);
and U7316 (N_7316,N_7139,N_7136);
nor U7317 (N_7317,N_7149,N_7115);
or U7318 (N_7318,N_7066,N_7152);
nor U7319 (N_7319,N_7045,N_7120);
xor U7320 (N_7320,N_7123,N_7131);
or U7321 (N_7321,N_7195,N_7129);
xnor U7322 (N_7322,N_7071,N_7085);
nor U7323 (N_7323,N_7183,N_7192);
xnor U7324 (N_7324,N_7048,N_7071);
or U7325 (N_7325,N_7071,N_7156);
xnor U7326 (N_7326,N_7169,N_7192);
nor U7327 (N_7327,N_7050,N_7089);
nor U7328 (N_7328,N_7165,N_7148);
nor U7329 (N_7329,N_7054,N_7075);
nor U7330 (N_7330,N_7106,N_7192);
xnor U7331 (N_7331,N_7109,N_7177);
and U7332 (N_7332,N_7174,N_7132);
nor U7333 (N_7333,N_7136,N_7107);
and U7334 (N_7334,N_7129,N_7076);
nand U7335 (N_7335,N_7148,N_7114);
nor U7336 (N_7336,N_7127,N_7102);
or U7337 (N_7337,N_7109,N_7133);
and U7338 (N_7338,N_7128,N_7116);
and U7339 (N_7339,N_7092,N_7066);
or U7340 (N_7340,N_7164,N_7097);
and U7341 (N_7341,N_7048,N_7191);
and U7342 (N_7342,N_7042,N_7082);
or U7343 (N_7343,N_7058,N_7198);
and U7344 (N_7344,N_7094,N_7075);
xor U7345 (N_7345,N_7087,N_7190);
nand U7346 (N_7346,N_7199,N_7177);
or U7347 (N_7347,N_7089,N_7161);
or U7348 (N_7348,N_7146,N_7113);
and U7349 (N_7349,N_7075,N_7113);
xor U7350 (N_7350,N_7153,N_7067);
nand U7351 (N_7351,N_7086,N_7100);
and U7352 (N_7352,N_7191,N_7135);
or U7353 (N_7353,N_7140,N_7197);
nor U7354 (N_7354,N_7188,N_7104);
and U7355 (N_7355,N_7173,N_7131);
or U7356 (N_7356,N_7069,N_7048);
nand U7357 (N_7357,N_7065,N_7078);
xor U7358 (N_7358,N_7054,N_7068);
or U7359 (N_7359,N_7080,N_7129);
xor U7360 (N_7360,N_7314,N_7283);
nand U7361 (N_7361,N_7330,N_7222);
nand U7362 (N_7362,N_7333,N_7354);
nand U7363 (N_7363,N_7352,N_7242);
and U7364 (N_7364,N_7350,N_7217);
nor U7365 (N_7365,N_7232,N_7219);
or U7366 (N_7366,N_7267,N_7353);
xnor U7367 (N_7367,N_7235,N_7311);
nor U7368 (N_7368,N_7339,N_7230);
or U7369 (N_7369,N_7218,N_7313);
nand U7370 (N_7370,N_7228,N_7225);
xnor U7371 (N_7371,N_7270,N_7316);
or U7372 (N_7372,N_7293,N_7359);
or U7373 (N_7373,N_7327,N_7212);
xor U7374 (N_7374,N_7261,N_7298);
xnor U7375 (N_7375,N_7325,N_7202);
or U7376 (N_7376,N_7345,N_7266);
and U7377 (N_7377,N_7328,N_7326);
and U7378 (N_7378,N_7205,N_7348);
nor U7379 (N_7379,N_7320,N_7246);
or U7380 (N_7380,N_7337,N_7340);
or U7381 (N_7381,N_7286,N_7201);
or U7382 (N_7382,N_7309,N_7210);
and U7383 (N_7383,N_7216,N_7227);
or U7384 (N_7384,N_7296,N_7253);
nor U7385 (N_7385,N_7310,N_7284);
or U7386 (N_7386,N_7244,N_7317);
or U7387 (N_7387,N_7204,N_7341);
xor U7388 (N_7388,N_7254,N_7272);
and U7389 (N_7389,N_7299,N_7245);
nor U7390 (N_7390,N_7335,N_7291);
nand U7391 (N_7391,N_7236,N_7211);
and U7392 (N_7392,N_7280,N_7241);
and U7393 (N_7393,N_7289,N_7255);
and U7394 (N_7394,N_7221,N_7220);
and U7395 (N_7395,N_7251,N_7297);
nor U7396 (N_7396,N_7269,N_7290);
nor U7397 (N_7397,N_7234,N_7356);
xnor U7398 (N_7398,N_7319,N_7276);
nor U7399 (N_7399,N_7274,N_7268);
and U7400 (N_7400,N_7240,N_7287);
and U7401 (N_7401,N_7342,N_7223);
nor U7402 (N_7402,N_7323,N_7306);
nor U7403 (N_7403,N_7229,N_7252);
and U7404 (N_7404,N_7301,N_7226);
nand U7405 (N_7405,N_7206,N_7332);
xnor U7406 (N_7406,N_7347,N_7358);
nand U7407 (N_7407,N_7346,N_7305);
nor U7408 (N_7408,N_7322,N_7263);
xor U7409 (N_7409,N_7295,N_7334);
xnor U7410 (N_7410,N_7277,N_7258);
or U7411 (N_7411,N_7288,N_7231);
nor U7412 (N_7412,N_7247,N_7213);
or U7413 (N_7413,N_7279,N_7308);
nand U7414 (N_7414,N_7214,N_7250);
nor U7415 (N_7415,N_7278,N_7331);
or U7416 (N_7416,N_7307,N_7304);
nor U7417 (N_7417,N_7312,N_7256);
nand U7418 (N_7418,N_7243,N_7273);
xor U7419 (N_7419,N_7281,N_7237);
nand U7420 (N_7420,N_7264,N_7248);
or U7421 (N_7421,N_7355,N_7292);
xor U7422 (N_7422,N_7318,N_7265);
and U7423 (N_7423,N_7209,N_7349);
nor U7424 (N_7424,N_7257,N_7351);
xnor U7425 (N_7425,N_7357,N_7259);
nand U7426 (N_7426,N_7321,N_7338);
or U7427 (N_7427,N_7302,N_7200);
xor U7428 (N_7428,N_7344,N_7260);
xor U7429 (N_7429,N_7315,N_7215);
or U7430 (N_7430,N_7300,N_7249);
nor U7431 (N_7431,N_7294,N_7303);
xor U7432 (N_7432,N_7208,N_7203);
nor U7433 (N_7433,N_7224,N_7271);
nor U7434 (N_7434,N_7343,N_7233);
xor U7435 (N_7435,N_7336,N_7238);
or U7436 (N_7436,N_7282,N_7275);
and U7437 (N_7437,N_7239,N_7285);
and U7438 (N_7438,N_7262,N_7329);
nand U7439 (N_7439,N_7324,N_7207);
or U7440 (N_7440,N_7344,N_7264);
xor U7441 (N_7441,N_7324,N_7293);
nor U7442 (N_7442,N_7244,N_7323);
nand U7443 (N_7443,N_7207,N_7349);
or U7444 (N_7444,N_7252,N_7287);
nand U7445 (N_7445,N_7241,N_7352);
and U7446 (N_7446,N_7319,N_7328);
and U7447 (N_7447,N_7221,N_7329);
nor U7448 (N_7448,N_7306,N_7281);
and U7449 (N_7449,N_7296,N_7292);
xnor U7450 (N_7450,N_7340,N_7235);
and U7451 (N_7451,N_7209,N_7270);
nand U7452 (N_7452,N_7234,N_7232);
or U7453 (N_7453,N_7276,N_7292);
nor U7454 (N_7454,N_7226,N_7314);
nor U7455 (N_7455,N_7216,N_7322);
xnor U7456 (N_7456,N_7204,N_7237);
xor U7457 (N_7457,N_7301,N_7231);
and U7458 (N_7458,N_7311,N_7333);
xnor U7459 (N_7459,N_7204,N_7203);
nand U7460 (N_7460,N_7240,N_7277);
or U7461 (N_7461,N_7215,N_7222);
xor U7462 (N_7462,N_7336,N_7311);
nand U7463 (N_7463,N_7219,N_7256);
xor U7464 (N_7464,N_7268,N_7338);
nor U7465 (N_7465,N_7348,N_7257);
nor U7466 (N_7466,N_7281,N_7301);
and U7467 (N_7467,N_7324,N_7264);
nor U7468 (N_7468,N_7294,N_7355);
nor U7469 (N_7469,N_7282,N_7357);
and U7470 (N_7470,N_7316,N_7329);
nand U7471 (N_7471,N_7257,N_7247);
nand U7472 (N_7472,N_7290,N_7256);
and U7473 (N_7473,N_7201,N_7296);
nor U7474 (N_7474,N_7232,N_7353);
or U7475 (N_7475,N_7301,N_7283);
or U7476 (N_7476,N_7340,N_7280);
nand U7477 (N_7477,N_7278,N_7216);
nand U7478 (N_7478,N_7274,N_7216);
nor U7479 (N_7479,N_7265,N_7323);
and U7480 (N_7480,N_7268,N_7309);
or U7481 (N_7481,N_7207,N_7240);
and U7482 (N_7482,N_7225,N_7204);
nor U7483 (N_7483,N_7283,N_7315);
nor U7484 (N_7484,N_7327,N_7305);
nand U7485 (N_7485,N_7264,N_7348);
nand U7486 (N_7486,N_7304,N_7330);
nor U7487 (N_7487,N_7260,N_7296);
nand U7488 (N_7488,N_7328,N_7289);
nand U7489 (N_7489,N_7288,N_7280);
nand U7490 (N_7490,N_7357,N_7332);
or U7491 (N_7491,N_7262,N_7232);
xnor U7492 (N_7492,N_7305,N_7315);
nor U7493 (N_7493,N_7357,N_7299);
xnor U7494 (N_7494,N_7319,N_7258);
or U7495 (N_7495,N_7336,N_7357);
nand U7496 (N_7496,N_7343,N_7296);
nor U7497 (N_7497,N_7329,N_7214);
nor U7498 (N_7498,N_7259,N_7249);
and U7499 (N_7499,N_7234,N_7231);
nor U7500 (N_7500,N_7306,N_7269);
and U7501 (N_7501,N_7308,N_7204);
or U7502 (N_7502,N_7261,N_7202);
or U7503 (N_7503,N_7285,N_7258);
and U7504 (N_7504,N_7274,N_7321);
xor U7505 (N_7505,N_7295,N_7264);
or U7506 (N_7506,N_7342,N_7328);
xor U7507 (N_7507,N_7214,N_7284);
nor U7508 (N_7508,N_7230,N_7243);
and U7509 (N_7509,N_7333,N_7267);
and U7510 (N_7510,N_7352,N_7298);
nor U7511 (N_7511,N_7243,N_7280);
nor U7512 (N_7512,N_7248,N_7288);
nand U7513 (N_7513,N_7220,N_7264);
or U7514 (N_7514,N_7304,N_7253);
xnor U7515 (N_7515,N_7334,N_7231);
xnor U7516 (N_7516,N_7211,N_7356);
xnor U7517 (N_7517,N_7326,N_7232);
nand U7518 (N_7518,N_7287,N_7299);
xnor U7519 (N_7519,N_7290,N_7267);
nand U7520 (N_7520,N_7411,N_7464);
or U7521 (N_7521,N_7448,N_7413);
or U7522 (N_7522,N_7425,N_7515);
xor U7523 (N_7523,N_7518,N_7458);
nand U7524 (N_7524,N_7361,N_7468);
xor U7525 (N_7525,N_7439,N_7360);
xnor U7526 (N_7526,N_7457,N_7386);
and U7527 (N_7527,N_7365,N_7442);
and U7528 (N_7528,N_7364,N_7378);
and U7529 (N_7529,N_7429,N_7397);
nand U7530 (N_7530,N_7467,N_7362);
nand U7531 (N_7531,N_7470,N_7499);
or U7532 (N_7532,N_7484,N_7400);
and U7533 (N_7533,N_7434,N_7422);
xnor U7534 (N_7534,N_7431,N_7452);
nor U7535 (N_7535,N_7466,N_7381);
xnor U7536 (N_7536,N_7462,N_7404);
xnor U7537 (N_7537,N_7443,N_7449);
or U7538 (N_7538,N_7367,N_7389);
nand U7539 (N_7539,N_7432,N_7372);
xnor U7540 (N_7540,N_7412,N_7513);
or U7541 (N_7541,N_7454,N_7433);
xor U7542 (N_7542,N_7480,N_7446);
nand U7543 (N_7543,N_7420,N_7504);
and U7544 (N_7544,N_7380,N_7385);
or U7545 (N_7545,N_7419,N_7424);
nand U7546 (N_7546,N_7410,N_7374);
nand U7547 (N_7547,N_7370,N_7415);
nor U7548 (N_7548,N_7398,N_7395);
nor U7549 (N_7549,N_7475,N_7408);
and U7550 (N_7550,N_7407,N_7486);
xor U7551 (N_7551,N_7471,N_7399);
nor U7552 (N_7552,N_7450,N_7498);
xnor U7553 (N_7553,N_7496,N_7519);
nor U7554 (N_7554,N_7376,N_7423);
nand U7555 (N_7555,N_7510,N_7368);
nand U7556 (N_7556,N_7463,N_7490);
nand U7557 (N_7557,N_7384,N_7441);
nand U7558 (N_7558,N_7465,N_7375);
or U7559 (N_7559,N_7500,N_7494);
nor U7560 (N_7560,N_7474,N_7477);
or U7561 (N_7561,N_7507,N_7421);
nor U7562 (N_7562,N_7511,N_7483);
or U7563 (N_7563,N_7377,N_7481);
xor U7564 (N_7564,N_7516,N_7388);
nor U7565 (N_7565,N_7491,N_7461);
or U7566 (N_7566,N_7418,N_7478);
or U7567 (N_7567,N_7438,N_7440);
nand U7568 (N_7568,N_7489,N_7373);
nor U7569 (N_7569,N_7445,N_7479);
xor U7570 (N_7570,N_7492,N_7508);
or U7571 (N_7571,N_7417,N_7488);
or U7572 (N_7572,N_7472,N_7382);
or U7573 (N_7573,N_7460,N_7485);
and U7574 (N_7574,N_7392,N_7509);
xor U7575 (N_7575,N_7453,N_7495);
xor U7576 (N_7576,N_7435,N_7469);
nor U7577 (N_7577,N_7401,N_7493);
xor U7578 (N_7578,N_7447,N_7394);
or U7579 (N_7579,N_7379,N_7393);
and U7580 (N_7580,N_7473,N_7456);
nor U7581 (N_7581,N_7428,N_7427);
nor U7582 (N_7582,N_7403,N_7416);
and U7583 (N_7583,N_7459,N_7371);
nor U7584 (N_7584,N_7437,N_7497);
xnor U7585 (N_7585,N_7436,N_7455);
xor U7586 (N_7586,N_7387,N_7512);
and U7587 (N_7587,N_7501,N_7390);
or U7588 (N_7588,N_7409,N_7482);
nor U7589 (N_7589,N_7476,N_7505);
nor U7590 (N_7590,N_7487,N_7430);
xnor U7591 (N_7591,N_7451,N_7396);
and U7592 (N_7592,N_7405,N_7391);
nand U7593 (N_7593,N_7406,N_7506);
nor U7594 (N_7594,N_7426,N_7444);
nand U7595 (N_7595,N_7503,N_7414);
nor U7596 (N_7596,N_7363,N_7383);
nor U7597 (N_7597,N_7366,N_7502);
or U7598 (N_7598,N_7517,N_7514);
or U7599 (N_7599,N_7402,N_7369);
nand U7600 (N_7600,N_7510,N_7439);
nand U7601 (N_7601,N_7432,N_7402);
and U7602 (N_7602,N_7467,N_7421);
nor U7603 (N_7603,N_7469,N_7431);
nor U7604 (N_7604,N_7473,N_7469);
nor U7605 (N_7605,N_7456,N_7409);
and U7606 (N_7606,N_7467,N_7429);
or U7607 (N_7607,N_7508,N_7467);
xor U7608 (N_7608,N_7376,N_7492);
nand U7609 (N_7609,N_7394,N_7366);
or U7610 (N_7610,N_7387,N_7388);
or U7611 (N_7611,N_7362,N_7391);
xnor U7612 (N_7612,N_7469,N_7491);
nor U7613 (N_7613,N_7395,N_7508);
nor U7614 (N_7614,N_7377,N_7503);
or U7615 (N_7615,N_7390,N_7380);
nand U7616 (N_7616,N_7402,N_7407);
nand U7617 (N_7617,N_7402,N_7496);
and U7618 (N_7618,N_7459,N_7513);
nor U7619 (N_7619,N_7420,N_7516);
xor U7620 (N_7620,N_7362,N_7360);
or U7621 (N_7621,N_7510,N_7487);
nor U7622 (N_7622,N_7415,N_7477);
or U7623 (N_7623,N_7393,N_7476);
xnor U7624 (N_7624,N_7443,N_7406);
nand U7625 (N_7625,N_7505,N_7407);
or U7626 (N_7626,N_7455,N_7368);
xor U7627 (N_7627,N_7501,N_7380);
nand U7628 (N_7628,N_7410,N_7441);
nor U7629 (N_7629,N_7439,N_7517);
or U7630 (N_7630,N_7495,N_7483);
nand U7631 (N_7631,N_7444,N_7406);
xor U7632 (N_7632,N_7486,N_7387);
or U7633 (N_7633,N_7487,N_7470);
and U7634 (N_7634,N_7398,N_7410);
xor U7635 (N_7635,N_7491,N_7442);
nor U7636 (N_7636,N_7504,N_7480);
and U7637 (N_7637,N_7516,N_7448);
or U7638 (N_7638,N_7411,N_7385);
nor U7639 (N_7639,N_7425,N_7415);
nand U7640 (N_7640,N_7444,N_7482);
or U7641 (N_7641,N_7411,N_7366);
and U7642 (N_7642,N_7474,N_7411);
nand U7643 (N_7643,N_7446,N_7401);
nand U7644 (N_7644,N_7503,N_7485);
nand U7645 (N_7645,N_7428,N_7380);
xnor U7646 (N_7646,N_7437,N_7453);
nor U7647 (N_7647,N_7417,N_7466);
nand U7648 (N_7648,N_7507,N_7392);
nand U7649 (N_7649,N_7381,N_7418);
xor U7650 (N_7650,N_7449,N_7400);
and U7651 (N_7651,N_7428,N_7442);
or U7652 (N_7652,N_7387,N_7366);
nor U7653 (N_7653,N_7476,N_7414);
nand U7654 (N_7654,N_7384,N_7463);
and U7655 (N_7655,N_7399,N_7410);
xnor U7656 (N_7656,N_7434,N_7415);
nand U7657 (N_7657,N_7404,N_7487);
and U7658 (N_7658,N_7494,N_7443);
nand U7659 (N_7659,N_7461,N_7372);
nor U7660 (N_7660,N_7364,N_7503);
nor U7661 (N_7661,N_7410,N_7445);
nor U7662 (N_7662,N_7515,N_7446);
or U7663 (N_7663,N_7416,N_7375);
and U7664 (N_7664,N_7488,N_7466);
nand U7665 (N_7665,N_7446,N_7434);
nor U7666 (N_7666,N_7428,N_7403);
and U7667 (N_7667,N_7393,N_7411);
xnor U7668 (N_7668,N_7519,N_7512);
xnor U7669 (N_7669,N_7429,N_7474);
or U7670 (N_7670,N_7463,N_7391);
nand U7671 (N_7671,N_7438,N_7425);
xor U7672 (N_7672,N_7423,N_7377);
or U7673 (N_7673,N_7366,N_7508);
and U7674 (N_7674,N_7399,N_7422);
or U7675 (N_7675,N_7442,N_7404);
and U7676 (N_7676,N_7496,N_7486);
xor U7677 (N_7677,N_7475,N_7428);
xor U7678 (N_7678,N_7480,N_7418);
xor U7679 (N_7679,N_7428,N_7471);
nand U7680 (N_7680,N_7622,N_7632);
nor U7681 (N_7681,N_7593,N_7641);
or U7682 (N_7682,N_7635,N_7678);
nand U7683 (N_7683,N_7557,N_7566);
and U7684 (N_7684,N_7657,N_7651);
or U7685 (N_7685,N_7570,N_7533);
nand U7686 (N_7686,N_7572,N_7523);
and U7687 (N_7687,N_7528,N_7598);
and U7688 (N_7688,N_7628,N_7580);
xor U7689 (N_7689,N_7567,N_7640);
xor U7690 (N_7690,N_7620,N_7574);
nand U7691 (N_7691,N_7627,N_7659);
nand U7692 (N_7692,N_7670,N_7631);
and U7693 (N_7693,N_7526,N_7595);
or U7694 (N_7694,N_7599,N_7653);
xnor U7695 (N_7695,N_7672,N_7527);
and U7696 (N_7696,N_7532,N_7536);
nand U7697 (N_7697,N_7596,N_7551);
and U7698 (N_7698,N_7669,N_7558);
nor U7699 (N_7699,N_7562,N_7529);
or U7700 (N_7700,N_7675,N_7582);
xnor U7701 (N_7701,N_7552,N_7613);
or U7702 (N_7702,N_7619,N_7674);
nor U7703 (N_7703,N_7556,N_7525);
nor U7704 (N_7704,N_7543,N_7667);
or U7705 (N_7705,N_7553,N_7626);
nor U7706 (N_7706,N_7542,N_7521);
xor U7707 (N_7707,N_7600,N_7605);
xnor U7708 (N_7708,N_7573,N_7665);
and U7709 (N_7709,N_7544,N_7643);
xor U7710 (N_7710,N_7637,N_7661);
or U7711 (N_7711,N_7645,N_7671);
xor U7712 (N_7712,N_7537,N_7662);
nor U7713 (N_7713,N_7618,N_7594);
or U7714 (N_7714,N_7548,N_7625);
nor U7715 (N_7715,N_7609,N_7560);
and U7716 (N_7716,N_7629,N_7520);
and U7717 (N_7717,N_7577,N_7581);
or U7718 (N_7718,N_7545,N_7564);
and U7719 (N_7719,N_7656,N_7623);
nand U7720 (N_7720,N_7655,N_7654);
nand U7721 (N_7721,N_7597,N_7559);
or U7722 (N_7722,N_7565,N_7588);
xnor U7723 (N_7723,N_7677,N_7578);
and U7724 (N_7724,N_7571,N_7610);
nand U7725 (N_7725,N_7601,N_7602);
and U7726 (N_7726,N_7647,N_7646);
xnor U7727 (N_7727,N_7584,N_7624);
nand U7728 (N_7728,N_7615,N_7583);
and U7729 (N_7729,N_7534,N_7603);
nand U7730 (N_7730,N_7658,N_7633);
or U7731 (N_7731,N_7634,N_7604);
xor U7732 (N_7732,N_7555,N_7636);
nor U7733 (N_7733,N_7642,N_7550);
and U7734 (N_7734,N_7561,N_7614);
nand U7735 (N_7735,N_7540,N_7538);
and U7736 (N_7736,N_7587,N_7676);
xor U7737 (N_7737,N_7586,N_7576);
and U7738 (N_7738,N_7591,N_7650);
nand U7739 (N_7739,N_7579,N_7649);
and U7740 (N_7740,N_7611,N_7585);
xor U7741 (N_7741,N_7638,N_7679);
or U7742 (N_7742,N_7617,N_7612);
xnor U7743 (N_7743,N_7663,N_7568);
nor U7744 (N_7744,N_7607,N_7668);
and U7745 (N_7745,N_7541,N_7522);
and U7746 (N_7746,N_7589,N_7666);
xnor U7747 (N_7747,N_7630,N_7531);
xnor U7748 (N_7748,N_7621,N_7660);
xor U7749 (N_7749,N_7547,N_7549);
nand U7750 (N_7750,N_7608,N_7575);
nand U7751 (N_7751,N_7535,N_7673);
xor U7752 (N_7752,N_7592,N_7590);
nand U7753 (N_7753,N_7639,N_7539);
nor U7754 (N_7754,N_7569,N_7546);
and U7755 (N_7755,N_7606,N_7616);
or U7756 (N_7756,N_7652,N_7530);
nand U7757 (N_7757,N_7554,N_7563);
and U7758 (N_7758,N_7524,N_7644);
nand U7759 (N_7759,N_7648,N_7664);
xnor U7760 (N_7760,N_7674,N_7566);
xnor U7761 (N_7761,N_7564,N_7521);
nor U7762 (N_7762,N_7585,N_7668);
or U7763 (N_7763,N_7638,N_7549);
nor U7764 (N_7764,N_7614,N_7543);
and U7765 (N_7765,N_7674,N_7568);
and U7766 (N_7766,N_7552,N_7542);
xnor U7767 (N_7767,N_7597,N_7571);
nor U7768 (N_7768,N_7672,N_7641);
and U7769 (N_7769,N_7673,N_7534);
nor U7770 (N_7770,N_7597,N_7620);
or U7771 (N_7771,N_7654,N_7549);
and U7772 (N_7772,N_7609,N_7570);
and U7773 (N_7773,N_7579,N_7557);
and U7774 (N_7774,N_7539,N_7647);
xor U7775 (N_7775,N_7593,N_7664);
and U7776 (N_7776,N_7608,N_7610);
or U7777 (N_7777,N_7649,N_7573);
nor U7778 (N_7778,N_7644,N_7664);
and U7779 (N_7779,N_7678,N_7672);
or U7780 (N_7780,N_7589,N_7602);
or U7781 (N_7781,N_7539,N_7672);
or U7782 (N_7782,N_7584,N_7541);
or U7783 (N_7783,N_7659,N_7600);
nor U7784 (N_7784,N_7637,N_7664);
nand U7785 (N_7785,N_7662,N_7646);
nand U7786 (N_7786,N_7676,N_7664);
and U7787 (N_7787,N_7544,N_7567);
nor U7788 (N_7788,N_7547,N_7551);
nor U7789 (N_7789,N_7546,N_7658);
xnor U7790 (N_7790,N_7658,N_7527);
or U7791 (N_7791,N_7594,N_7559);
xnor U7792 (N_7792,N_7594,N_7535);
and U7793 (N_7793,N_7634,N_7628);
xnor U7794 (N_7794,N_7661,N_7597);
or U7795 (N_7795,N_7536,N_7603);
xor U7796 (N_7796,N_7650,N_7614);
or U7797 (N_7797,N_7557,N_7595);
xnor U7798 (N_7798,N_7672,N_7650);
nand U7799 (N_7799,N_7664,N_7635);
or U7800 (N_7800,N_7679,N_7556);
xnor U7801 (N_7801,N_7537,N_7525);
or U7802 (N_7802,N_7665,N_7624);
nand U7803 (N_7803,N_7665,N_7613);
or U7804 (N_7804,N_7669,N_7679);
nand U7805 (N_7805,N_7585,N_7669);
xor U7806 (N_7806,N_7555,N_7668);
xnor U7807 (N_7807,N_7647,N_7566);
xor U7808 (N_7808,N_7638,N_7675);
or U7809 (N_7809,N_7536,N_7640);
xnor U7810 (N_7810,N_7531,N_7670);
or U7811 (N_7811,N_7632,N_7600);
or U7812 (N_7812,N_7587,N_7572);
xnor U7813 (N_7813,N_7621,N_7568);
nor U7814 (N_7814,N_7614,N_7661);
xnor U7815 (N_7815,N_7545,N_7650);
xor U7816 (N_7816,N_7662,N_7654);
or U7817 (N_7817,N_7661,N_7625);
nand U7818 (N_7818,N_7521,N_7669);
xor U7819 (N_7819,N_7629,N_7590);
nand U7820 (N_7820,N_7567,N_7579);
nor U7821 (N_7821,N_7611,N_7659);
and U7822 (N_7822,N_7590,N_7598);
nand U7823 (N_7823,N_7523,N_7564);
nor U7824 (N_7824,N_7604,N_7644);
nand U7825 (N_7825,N_7675,N_7611);
or U7826 (N_7826,N_7595,N_7596);
nand U7827 (N_7827,N_7636,N_7593);
nor U7828 (N_7828,N_7527,N_7659);
and U7829 (N_7829,N_7592,N_7614);
xor U7830 (N_7830,N_7598,N_7604);
and U7831 (N_7831,N_7648,N_7582);
or U7832 (N_7832,N_7539,N_7600);
nand U7833 (N_7833,N_7660,N_7529);
nand U7834 (N_7834,N_7590,N_7556);
nor U7835 (N_7835,N_7575,N_7666);
nand U7836 (N_7836,N_7638,N_7637);
xor U7837 (N_7837,N_7672,N_7568);
and U7838 (N_7838,N_7609,N_7612);
xor U7839 (N_7839,N_7641,N_7553);
or U7840 (N_7840,N_7692,N_7832);
nor U7841 (N_7841,N_7761,N_7752);
nor U7842 (N_7842,N_7739,N_7793);
nor U7843 (N_7843,N_7811,N_7827);
or U7844 (N_7844,N_7683,N_7729);
and U7845 (N_7845,N_7770,N_7723);
or U7846 (N_7846,N_7753,N_7699);
nor U7847 (N_7847,N_7818,N_7706);
nor U7848 (N_7848,N_7792,N_7786);
or U7849 (N_7849,N_7834,N_7698);
xnor U7850 (N_7850,N_7708,N_7762);
and U7851 (N_7851,N_7791,N_7817);
nand U7852 (N_7852,N_7772,N_7743);
and U7853 (N_7853,N_7815,N_7738);
or U7854 (N_7854,N_7820,N_7730);
nor U7855 (N_7855,N_7731,N_7701);
xnor U7856 (N_7856,N_7798,N_7819);
and U7857 (N_7857,N_7720,N_7705);
and U7858 (N_7858,N_7754,N_7773);
or U7859 (N_7859,N_7800,N_7826);
or U7860 (N_7860,N_7728,N_7778);
and U7861 (N_7861,N_7736,N_7741);
nand U7862 (N_7862,N_7823,N_7745);
and U7863 (N_7863,N_7797,N_7764);
xnor U7864 (N_7864,N_7836,N_7774);
and U7865 (N_7865,N_7771,N_7696);
or U7866 (N_7866,N_7821,N_7837);
nor U7867 (N_7867,N_7765,N_7700);
nand U7868 (N_7868,N_7714,N_7694);
or U7869 (N_7869,N_7751,N_7782);
nor U7870 (N_7870,N_7795,N_7717);
or U7871 (N_7871,N_7803,N_7839);
xnor U7872 (N_7872,N_7732,N_7702);
xnor U7873 (N_7873,N_7830,N_7685);
and U7874 (N_7874,N_7713,N_7733);
nand U7875 (N_7875,N_7822,N_7727);
xnor U7876 (N_7876,N_7788,N_7777);
nand U7877 (N_7877,N_7686,N_7747);
or U7878 (N_7878,N_7718,N_7825);
xor U7879 (N_7879,N_7744,N_7711);
nor U7880 (N_7880,N_7790,N_7828);
xor U7881 (N_7881,N_7735,N_7755);
xor U7882 (N_7882,N_7759,N_7781);
or U7883 (N_7883,N_7681,N_7784);
and U7884 (N_7884,N_7835,N_7707);
nor U7885 (N_7885,N_7726,N_7780);
or U7886 (N_7886,N_7829,N_7783);
or U7887 (N_7887,N_7697,N_7813);
nand U7888 (N_7888,N_7808,N_7721);
and U7889 (N_7889,N_7689,N_7787);
and U7890 (N_7890,N_7758,N_7688);
nand U7891 (N_7891,N_7703,N_7746);
nand U7892 (N_7892,N_7710,N_7682);
and U7893 (N_7893,N_7801,N_7766);
and U7894 (N_7894,N_7734,N_7794);
xor U7895 (N_7895,N_7789,N_7838);
or U7896 (N_7896,N_7814,N_7716);
nor U7897 (N_7897,N_7824,N_7806);
xor U7898 (N_7898,N_7740,N_7693);
and U7899 (N_7899,N_7757,N_7775);
nand U7900 (N_7900,N_7804,N_7805);
nor U7901 (N_7901,N_7799,N_7807);
and U7902 (N_7902,N_7763,N_7680);
nand U7903 (N_7903,N_7704,N_7687);
nor U7904 (N_7904,N_7779,N_7810);
nor U7905 (N_7905,N_7749,N_7724);
xnor U7906 (N_7906,N_7742,N_7709);
or U7907 (N_7907,N_7769,N_7776);
nor U7908 (N_7908,N_7833,N_7816);
xnor U7909 (N_7909,N_7719,N_7768);
nand U7910 (N_7910,N_7691,N_7767);
nand U7911 (N_7911,N_7812,N_7750);
or U7912 (N_7912,N_7756,N_7712);
and U7913 (N_7913,N_7748,N_7725);
xnor U7914 (N_7914,N_7831,N_7722);
xnor U7915 (N_7915,N_7695,N_7760);
nand U7916 (N_7916,N_7785,N_7737);
or U7917 (N_7917,N_7684,N_7690);
or U7918 (N_7918,N_7809,N_7802);
and U7919 (N_7919,N_7796,N_7715);
xor U7920 (N_7920,N_7733,N_7793);
nand U7921 (N_7921,N_7703,N_7749);
nor U7922 (N_7922,N_7777,N_7779);
or U7923 (N_7923,N_7704,N_7755);
or U7924 (N_7924,N_7816,N_7791);
nand U7925 (N_7925,N_7775,N_7787);
and U7926 (N_7926,N_7792,N_7825);
xor U7927 (N_7927,N_7759,N_7783);
and U7928 (N_7928,N_7724,N_7767);
nor U7929 (N_7929,N_7691,N_7716);
xnor U7930 (N_7930,N_7831,N_7833);
or U7931 (N_7931,N_7713,N_7688);
nand U7932 (N_7932,N_7698,N_7799);
xnor U7933 (N_7933,N_7701,N_7706);
and U7934 (N_7934,N_7789,N_7730);
or U7935 (N_7935,N_7775,N_7753);
nand U7936 (N_7936,N_7683,N_7803);
or U7937 (N_7937,N_7790,N_7722);
xnor U7938 (N_7938,N_7731,N_7753);
and U7939 (N_7939,N_7815,N_7773);
and U7940 (N_7940,N_7728,N_7737);
and U7941 (N_7941,N_7681,N_7740);
nand U7942 (N_7942,N_7768,N_7680);
nand U7943 (N_7943,N_7741,N_7756);
nand U7944 (N_7944,N_7785,N_7712);
xor U7945 (N_7945,N_7695,N_7719);
nor U7946 (N_7946,N_7827,N_7714);
or U7947 (N_7947,N_7836,N_7735);
nor U7948 (N_7948,N_7773,N_7837);
or U7949 (N_7949,N_7742,N_7682);
or U7950 (N_7950,N_7752,N_7816);
xnor U7951 (N_7951,N_7715,N_7753);
nand U7952 (N_7952,N_7755,N_7722);
or U7953 (N_7953,N_7690,N_7691);
nand U7954 (N_7954,N_7707,N_7685);
xnor U7955 (N_7955,N_7837,N_7830);
and U7956 (N_7956,N_7820,N_7724);
xor U7957 (N_7957,N_7698,N_7804);
xor U7958 (N_7958,N_7769,N_7830);
nand U7959 (N_7959,N_7807,N_7724);
nand U7960 (N_7960,N_7699,N_7757);
and U7961 (N_7961,N_7778,N_7708);
and U7962 (N_7962,N_7753,N_7748);
and U7963 (N_7963,N_7726,N_7788);
and U7964 (N_7964,N_7771,N_7766);
nand U7965 (N_7965,N_7697,N_7775);
xnor U7966 (N_7966,N_7784,N_7798);
nor U7967 (N_7967,N_7712,N_7741);
or U7968 (N_7968,N_7696,N_7823);
nor U7969 (N_7969,N_7814,N_7770);
xnor U7970 (N_7970,N_7743,N_7702);
or U7971 (N_7971,N_7774,N_7691);
xnor U7972 (N_7972,N_7682,N_7731);
xor U7973 (N_7973,N_7701,N_7691);
and U7974 (N_7974,N_7740,N_7684);
or U7975 (N_7975,N_7681,N_7811);
nand U7976 (N_7976,N_7798,N_7807);
and U7977 (N_7977,N_7823,N_7703);
and U7978 (N_7978,N_7793,N_7755);
or U7979 (N_7979,N_7710,N_7797);
and U7980 (N_7980,N_7736,N_7700);
and U7981 (N_7981,N_7741,N_7819);
nor U7982 (N_7982,N_7697,N_7819);
xor U7983 (N_7983,N_7757,N_7722);
nor U7984 (N_7984,N_7835,N_7818);
or U7985 (N_7985,N_7834,N_7704);
xnor U7986 (N_7986,N_7788,N_7744);
xnor U7987 (N_7987,N_7820,N_7801);
nor U7988 (N_7988,N_7711,N_7781);
or U7989 (N_7989,N_7818,N_7774);
xor U7990 (N_7990,N_7754,N_7779);
or U7991 (N_7991,N_7684,N_7745);
and U7992 (N_7992,N_7714,N_7681);
nand U7993 (N_7993,N_7746,N_7785);
nor U7994 (N_7994,N_7763,N_7727);
nor U7995 (N_7995,N_7780,N_7751);
xor U7996 (N_7996,N_7802,N_7739);
or U7997 (N_7997,N_7691,N_7751);
nor U7998 (N_7998,N_7759,N_7753);
and U7999 (N_7999,N_7725,N_7683);
nand U8000 (N_8000,N_7917,N_7897);
and U8001 (N_8001,N_7985,N_7843);
xnor U8002 (N_8002,N_7852,N_7915);
nor U8003 (N_8003,N_7901,N_7943);
or U8004 (N_8004,N_7841,N_7976);
or U8005 (N_8005,N_7858,N_7942);
nand U8006 (N_8006,N_7940,N_7848);
or U8007 (N_8007,N_7908,N_7885);
xnor U8008 (N_8008,N_7864,N_7883);
nand U8009 (N_8009,N_7990,N_7880);
and U8010 (N_8010,N_7930,N_7863);
nand U8011 (N_8011,N_7980,N_7845);
nor U8012 (N_8012,N_7849,N_7945);
nor U8013 (N_8013,N_7920,N_7861);
or U8014 (N_8014,N_7928,N_7941);
or U8015 (N_8015,N_7904,N_7998);
xnor U8016 (N_8016,N_7936,N_7951);
or U8017 (N_8017,N_7874,N_7869);
or U8018 (N_8018,N_7909,N_7873);
or U8019 (N_8019,N_7854,N_7856);
or U8020 (N_8020,N_7919,N_7857);
or U8021 (N_8021,N_7987,N_7906);
nand U8022 (N_8022,N_7911,N_7887);
nand U8023 (N_8023,N_7844,N_7879);
xor U8024 (N_8024,N_7872,N_7949);
nor U8025 (N_8025,N_7921,N_7865);
nor U8026 (N_8026,N_7960,N_7931);
nor U8027 (N_8027,N_7999,N_7892);
and U8028 (N_8028,N_7914,N_7963);
nand U8029 (N_8029,N_7981,N_7957);
or U8030 (N_8030,N_7958,N_7978);
or U8031 (N_8031,N_7886,N_7929);
xnor U8032 (N_8032,N_7905,N_7891);
and U8033 (N_8033,N_7893,N_7996);
and U8034 (N_8034,N_7953,N_7853);
and U8035 (N_8035,N_7900,N_7934);
or U8036 (N_8036,N_7932,N_7988);
nor U8037 (N_8037,N_7995,N_7875);
nand U8038 (N_8038,N_7989,N_7851);
and U8039 (N_8039,N_7968,N_7884);
and U8040 (N_8040,N_7890,N_7881);
xor U8041 (N_8041,N_7867,N_7860);
xor U8042 (N_8042,N_7946,N_7927);
xnor U8043 (N_8043,N_7916,N_7850);
or U8044 (N_8044,N_7926,N_7952);
xor U8045 (N_8045,N_7876,N_7910);
nor U8046 (N_8046,N_7944,N_7859);
nand U8047 (N_8047,N_7947,N_7882);
nor U8048 (N_8048,N_7913,N_7870);
or U8049 (N_8049,N_7918,N_7888);
xnor U8050 (N_8050,N_7974,N_7898);
nand U8051 (N_8051,N_7871,N_7924);
or U8052 (N_8052,N_7862,N_7842);
nand U8053 (N_8053,N_7984,N_7983);
nand U8054 (N_8054,N_7902,N_7948);
and U8055 (N_8055,N_7840,N_7956);
or U8056 (N_8056,N_7950,N_7969);
nor U8057 (N_8057,N_7972,N_7933);
nand U8058 (N_8058,N_7993,N_7986);
and U8059 (N_8059,N_7991,N_7971);
nand U8060 (N_8060,N_7896,N_7912);
nor U8061 (N_8061,N_7855,N_7970);
xnor U8062 (N_8062,N_7977,N_7922);
and U8063 (N_8063,N_7966,N_7847);
nor U8064 (N_8064,N_7889,N_7973);
nor U8065 (N_8065,N_7965,N_7935);
xnor U8066 (N_8066,N_7994,N_7907);
or U8067 (N_8067,N_7967,N_7899);
nor U8068 (N_8068,N_7975,N_7895);
or U8069 (N_8069,N_7962,N_7903);
xor U8070 (N_8070,N_7982,N_7923);
nand U8071 (N_8071,N_7959,N_7954);
or U8072 (N_8072,N_7894,N_7877);
and U8073 (N_8073,N_7878,N_7925);
nand U8074 (N_8074,N_7939,N_7938);
nand U8075 (N_8075,N_7997,N_7964);
nor U8076 (N_8076,N_7846,N_7992);
nor U8077 (N_8077,N_7955,N_7866);
or U8078 (N_8078,N_7868,N_7979);
xnor U8079 (N_8079,N_7937,N_7961);
nor U8080 (N_8080,N_7956,N_7895);
xor U8081 (N_8081,N_7952,N_7909);
xor U8082 (N_8082,N_7854,N_7945);
xor U8083 (N_8083,N_7925,N_7953);
and U8084 (N_8084,N_7989,N_7906);
or U8085 (N_8085,N_7957,N_7937);
xnor U8086 (N_8086,N_7848,N_7981);
nor U8087 (N_8087,N_7951,N_7946);
and U8088 (N_8088,N_7876,N_7886);
xor U8089 (N_8089,N_7969,N_7890);
or U8090 (N_8090,N_7841,N_7980);
or U8091 (N_8091,N_7952,N_7981);
nand U8092 (N_8092,N_7983,N_7951);
nor U8093 (N_8093,N_7982,N_7964);
and U8094 (N_8094,N_7842,N_7886);
xor U8095 (N_8095,N_7925,N_7944);
nor U8096 (N_8096,N_7986,N_7915);
or U8097 (N_8097,N_7971,N_7857);
xnor U8098 (N_8098,N_7856,N_7843);
and U8099 (N_8099,N_7958,N_7954);
nand U8100 (N_8100,N_7848,N_7925);
or U8101 (N_8101,N_7849,N_7949);
and U8102 (N_8102,N_7944,N_7908);
nand U8103 (N_8103,N_7928,N_7918);
or U8104 (N_8104,N_7985,N_7941);
or U8105 (N_8105,N_7950,N_7956);
and U8106 (N_8106,N_7903,N_7923);
or U8107 (N_8107,N_7880,N_7999);
and U8108 (N_8108,N_7878,N_7873);
or U8109 (N_8109,N_7865,N_7889);
or U8110 (N_8110,N_7940,N_7897);
and U8111 (N_8111,N_7859,N_7924);
or U8112 (N_8112,N_7923,N_7870);
or U8113 (N_8113,N_7887,N_7873);
or U8114 (N_8114,N_7930,N_7963);
or U8115 (N_8115,N_7973,N_7976);
nor U8116 (N_8116,N_7906,N_7967);
xor U8117 (N_8117,N_7844,N_7924);
and U8118 (N_8118,N_7919,N_7940);
and U8119 (N_8119,N_7965,N_7963);
and U8120 (N_8120,N_7957,N_7863);
and U8121 (N_8121,N_7848,N_7997);
or U8122 (N_8122,N_7949,N_7894);
nor U8123 (N_8123,N_7922,N_7862);
nor U8124 (N_8124,N_7861,N_7928);
or U8125 (N_8125,N_7886,N_7956);
nor U8126 (N_8126,N_7889,N_7996);
and U8127 (N_8127,N_7867,N_7845);
nand U8128 (N_8128,N_7986,N_7910);
or U8129 (N_8129,N_7897,N_7907);
nor U8130 (N_8130,N_7915,N_7970);
and U8131 (N_8131,N_7860,N_7974);
or U8132 (N_8132,N_7959,N_7904);
and U8133 (N_8133,N_7982,N_7989);
xor U8134 (N_8134,N_7989,N_7888);
nand U8135 (N_8135,N_7932,N_7867);
xor U8136 (N_8136,N_7917,N_7881);
nand U8137 (N_8137,N_7964,N_7975);
xnor U8138 (N_8138,N_7949,N_7923);
xnor U8139 (N_8139,N_7840,N_7974);
nor U8140 (N_8140,N_7886,N_7946);
xor U8141 (N_8141,N_7991,N_7994);
nand U8142 (N_8142,N_7879,N_7971);
or U8143 (N_8143,N_7853,N_7894);
nand U8144 (N_8144,N_7974,N_7998);
and U8145 (N_8145,N_7921,N_7910);
nand U8146 (N_8146,N_7937,N_7983);
and U8147 (N_8147,N_7949,N_7863);
xor U8148 (N_8148,N_7965,N_7998);
xor U8149 (N_8149,N_7901,N_7845);
and U8150 (N_8150,N_7987,N_7908);
and U8151 (N_8151,N_7988,N_7948);
xor U8152 (N_8152,N_7923,N_7868);
nor U8153 (N_8153,N_7952,N_7944);
xnor U8154 (N_8154,N_7968,N_7879);
xnor U8155 (N_8155,N_7975,N_7891);
xnor U8156 (N_8156,N_7875,N_7951);
nor U8157 (N_8157,N_7961,N_7872);
and U8158 (N_8158,N_7965,N_7975);
nand U8159 (N_8159,N_7912,N_7867);
and U8160 (N_8160,N_8013,N_8055);
or U8161 (N_8161,N_8001,N_8156);
xor U8162 (N_8162,N_8011,N_8135);
nor U8163 (N_8163,N_8074,N_8029);
and U8164 (N_8164,N_8057,N_8121);
nand U8165 (N_8165,N_8139,N_8008);
xnor U8166 (N_8166,N_8152,N_8095);
and U8167 (N_8167,N_8023,N_8035);
nor U8168 (N_8168,N_8090,N_8151);
or U8169 (N_8169,N_8002,N_8058);
xor U8170 (N_8170,N_8012,N_8133);
nand U8171 (N_8171,N_8076,N_8141);
xnor U8172 (N_8172,N_8053,N_8067);
xor U8173 (N_8173,N_8120,N_8144);
xor U8174 (N_8174,N_8089,N_8014);
nor U8175 (N_8175,N_8115,N_8025);
nand U8176 (N_8176,N_8159,N_8078);
and U8177 (N_8177,N_8022,N_8037);
and U8178 (N_8178,N_8009,N_8052);
xor U8179 (N_8179,N_8126,N_8111);
or U8180 (N_8180,N_8044,N_8131);
nand U8181 (N_8181,N_8048,N_8096);
nor U8182 (N_8182,N_8099,N_8024);
or U8183 (N_8183,N_8079,N_8026);
xor U8184 (N_8184,N_8146,N_8043);
nor U8185 (N_8185,N_8006,N_8117);
and U8186 (N_8186,N_8018,N_8085);
or U8187 (N_8187,N_8123,N_8045);
or U8188 (N_8188,N_8068,N_8064);
and U8189 (N_8189,N_8032,N_8038);
xnor U8190 (N_8190,N_8083,N_8030);
and U8191 (N_8191,N_8132,N_8070);
or U8192 (N_8192,N_8080,N_8075);
nand U8193 (N_8193,N_8145,N_8071);
or U8194 (N_8194,N_8114,N_8129);
nand U8195 (N_8195,N_8122,N_8059);
or U8196 (N_8196,N_8056,N_8039);
xor U8197 (N_8197,N_8153,N_8084);
nor U8198 (N_8198,N_8124,N_8154);
nand U8199 (N_8199,N_8158,N_8149);
xor U8200 (N_8200,N_8031,N_8138);
nor U8201 (N_8201,N_8102,N_8118);
nand U8202 (N_8202,N_8000,N_8063);
nor U8203 (N_8203,N_8060,N_8098);
or U8204 (N_8204,N_8104,N_8047);
or U8205 (N_8205,N_8112,N_8130);
nand U8206 (N_8206,N_8157,N_8027);
xnor U8207 (N_8207,N_8142,N_8086);
nor U8208 (N_8208,N_8109,N_8150);
xnor U8209 (N_8209,N_8019,N_8004);
nand U8210 (N_8210,N_8051,N_8028);
or U8211 (N_8211,N_8147,N_8033);
or U8212 (N_8212,N_8061,N_8093);
nand U8213 (N_8213,N_8127,N_8072);
xnor U8214 (N_8214,N_8015,N_8128);
and U8215 (N_8215,N_8049,N_8073);
nor U8216 (N_8216,N_8069,N_8020);
nor U8217 (N_8217,N_8040,N_8091);
xnor U8218 (N_8218,N_8017,N_8062);
xnor U8219 (N_8219,N_8105,N_8054);
nor U8220 (N_8220,N_8143,N_8066);
xnor U8221 (N_8221,N_8110,N_8113);
nor U8222 (N_8222,N_8137,N_8010);
and U8223 (N_8223,N_8107,N_8103);
or U8224 (N_8224,N_8036,N_8106);
or U8225 (N_8225,N_8097,N_8081);
xnor U8226 (N_8226,N_8136,N_8050);
xnor U8227 (N_8227,N_8108,N_8034);
nand U8228 (N_8228,N_8125,N_8021);
or U8229 (N_8229,N_8077,N_8140);
nand U8230 (N_8230,N_8119,N_8155);
or U8231 (N_8231,N_8088,N_8116);
or U8232 (N_8232,N_8101,N_8007);
and U8233 (N_8233,N_8134,N_8003);
and U8234 (N_8234,N_8016,N_8100);
or U8235 (N_8235,N_8082,N_8046);
or U8236 (N_8236,N_8087,N_8042);
or U8237 (N_8237,N_8041,N_8092);
nand U8238 (N_8238,N_8005,N_8065);
xor U8239 (N_8239,N_8094,N_8148);
or U8240 (N_8240,N_8157,N_8049);
xnor U8241 (N_8241,N_8091,N_8107);
xnor U8242 (N_8242,N_8054,N_8136);
nand U8243 (N_8243,N_8019,N_8110);
nor U8244 (N_8244,N_8137,N_8108);
and U8245 (N_8245,N_8033,N_8083);
xor U8246 (N_8246,N_8035,N_8047);
xor U8247 (N_8247,N_8058,N_8081);
or U8248 (N_8248,N_8074,N_8135);
nor U8249 (N_8249,N_8014,N_8063);
nor U8250 (N_8250,N_8009,N_8074);
nor U8251 (N_8251,N_8076,N_8138);
nor U8252 (N_8252,N_8063,N_8127);
nor U8253 (N_8253,N_8109,N_8029);
or U8254 (N_8254,N_8010,N_8148);
nor U8255 (N_8255,N_8031,N_8140);
or U8256 (N_8256,N_8158,N_8142);
nor U8257 (N_8257,N_8095,N_8066);
nand U8258 (N_8258,N_8055,N_8124);
nand U8259 (N_8259,N_8006,N_8046);
nand U8260 (N_8260,N_8076,N_8119);
nor U8261 (N_8261,N_8016,N_8053);
or U8262 (N_8262,N_8064,N_8069);
xnor U8263 (N_8263,N_8099,N_8135);
and U8264 (N_8264,N_8002,N_8140);
nand U8265 (N_8265,N_8054,N_8023);
xor U8266 (N_8266,N_8125,N_8056);
nor U8267 (N_8267,N_8109,N_8084);
nand U8268 (N_8268,N_8065,N_8032);
nor U8269 (N_8269,N_8093,N_8049);
xnor U8270 (N_8270,N_8153,N_8099);
nand U8271 (N_8271,N_8092,N_8007);
and U8272 (N_8272,N_8018,N_8053);
or U8273 (N_8273,N_8081,N_8033);
and U8274 (N_8274,N_8028,N_8103);
nor U8275 (N_8275,N_8118,N_8091);
or U8276 (N_8276,N_8130,N_8002);
and U8277 (N_8277,N_8067,N_8065);
nand U8278 (N_8278,N_8136,N_8051);
xnor U8279 (N_8279,N_8103,N_8078);
nor U8280 (N_8280,N_8159,N_8146);
or U8281 (N_8281,N_8101,N_8015);
nand U8282 (N_8282,N_8150,N_8081);
or U8283 (N_8283,N_8110,N_8089);
nor U8284 (N_8284,N_8087,N_8078);
or U8285 (N_8285,N_8155,N_8005);
nand U8286 (N_8286,N_8031,N_8055);
nor U8287 (N_8287,N_8048,N_8062);
and U8288 (N_8288,N_8146,N_8031);
nand U8289 (N_8289,N_8015,N_8153);
or U8290 (N_8290,N_8001,N_8124);
nor U8291 (N_8291,N_8041,N_8044);
xor U8292 (N_8292,N_8099,N_8062);
nor U8293 (N_8293,N_8131,N_8129);
and U8294 (N_8294,N_8099,N_8066);
nand U8295 (N_8295,N_8125,N_8128);
xnor U8296 (N_8296,N_8053,N_8074);
xor U8297 (N_8297,N_8052,N_8070);
or U8298 (N_8298,N_8103,N_8073);
xnor U8299 (N_8299,N_8008,N_8152);
nand U8300 (N_8300,N_8039,N_8123);
or U8301 (N_8301,N_8000,N_8046);
or U8302 (N_8302,N_8091,N_8057);
and U8303 (N_8303,N_8036,N_8115);
and U8304 (N_8304,N_8101,N_8068);
nand U8305 (N_8305,N_8123,N_8021);
and U8306 (N_8306,N_8000,N_8106);
nor U8307 (N_8307,N_8049,N_8130);
nand U8308 (N_8308,N_8102,N_8146);
xnor U8309 (N_8309,N_8043,N_8047);
and U8310 (N_8310,N_8109,N_8058);
nand U8311 (N_8311,N_8100,N_8046);
nor U8312 (N_8312,N_8084,N_8127);
and U8313 (N_8313,N_8088,N_8070);
nand U8314 (N_8314,N_8026,N_8007);
nor U8315 (N_8315,N_8137,N_8099);
or U8316 (N_8316,N_8042,N_8021);
xnor U8317 (N_8317,N_8090,N_8076);
xor U8318 (N_8318,N_8062,N_8005);
nor U8319 (N_8319,N_8147,N_8027);
or U8320 (N_8320,N_8217,N_8236);
nor U8321 (N_8321,N_8248,N_8192);
xnor U8322 (N_8322,N_8231,N_8164);
nor U8323 (N_8323,N_8182,N_8225);
and U8324 (N_8324,N_8240,N_8302);
xor U8325 (N_8325,N_8269,N_8180);
and U8326 (N_8326,N_8255,N_8163);
nand U8327 (N_8327,N_8268,N_8257);
and U8328 (N_8328,N_8216,N_8183);
nor U8329 (N_8329,N_8218,N_8287);
and U8330 (N_8330,N_8266,N_8209);
nor U8331 (N_8331,N_8283,N_8201);
xnor U8332 (N_8332,N_8271,N_8211);
xor U8333 (N_8333,N_8247,N_8237);
nor U8334 (N_8334,N_8214,N_8250);
nor U8335 (N_8335,N_8242,N_8205);
and U8336 (N_8336,N_8265,N_8303);
and U8337 (N_8337,N_8315,N_8219);
xnor U8338 (N_8338,N_8186,N_8256);
and U8339 (N_8339,N_8316,N_8197);
and U8340 (N_8340,N_8215,N_8304);
xnor U8341 (N_8341,N_8229,N_8312);
nand U8342 (N_8342,N_8233,N_8288);
xnor U8343 (N_8343,N_8244,N_8206);
xnor U8344 (N_8344,N_8223,N_8296);
or U8345 (N_8345,N_8204,N_8175);
or U8346 (N_8346,N_8263,N_8274);
nor U8347 (N_8347,N_8207,N_8230);
nor U8348 (N_8348,N_8319,N_8162);
or U8349 (N_8349,N_8294,N_8270);
nor U8350 (N_8350,N_8165,N_8307);
nand U8351 (N_8351,N_8196,N_8273);
and U8352 (N_8352,N_8221,N_8310);
nor U8353 (N_8353,N_8297,N_8241);
or U8354 (N_8354,N_8189,N_8188);
and U8355 (N_8355,N_8212,N_8278);
nand U8356 (N_8356,N_8202,N_8239);
nor U8357 (N_8357,N_8264,N_8262);
nor U8358 (N_8358,N_8293,N_8258);
nand U8359 (N_8359,N_8166,N_8193);
xnor U8360 (N_8360,N_8245,N_8260);
xor U8361 (N_8361,N_8190,N_8289);
xnor U8362 (N_8362,N_8198,N_8234);
xnor U8363 (N_8363,N_8308,N_8203);
xnor U8364 (N_8364,N_8170,N_8309);
nand U8365 (N_8365,N_8267,N_8282);
xnor U8366 (N_8366,N_8191,N_8185);
or U8367 (N_8367,N_8194,N_8295);
or U8368 (N_8368,N_8279,N_8160);
xnor U8369 (N_8369,N_8311,N_8246);
or U8370 (N_8370,N_8300,N_8318);
nand U8371 (N_8371,N_8227,N_8172);
or U8372 (N_8372,N_8187,N_8252);
and U8373 (N_8373,N_8226,N_8184);
and U8374 (N_8374,N_8210,N_8299);
xnor U8375 (N_8375,N_8243,N_8280);
and U8376 (N_8376,N_8168,N_8277);
nor U8377 (N_8377,N_8275,N_8292);
nor U8378 (N_8378,N_8181,N_8286);
xor U8379 (N_8379,N_8224,N_8161);
xnor U8380 (N_8380,N_8199,N_8232);
nand U8381 (N_8381,N_8272,N_8301);
xnor U8382 (N_8382,N_8208,N_8238);
nor U8383 (N_8383,N_8313,N_8317);
nand U8384 (N_8384,N_8291,N_8213);
nor U8385 (N_8385,N_8314,N_8290);
xnor U8386 (N_8386,N_8306,N_8174);
and U8387 (N_8387,N_8276,N_8220);
nand U8388 (N_8388,N_8195,N_8281);
or U8389 (N_8389,N_8228,N_8249);
nor U8390 (N_8390,N_8251,N_8176);
nor U8391 (N_8391,N_8254,N_8253);
nor U8392 (N_8392,N_8222,N_8179);
nand U8393 (N_8393,N_8200,N_8285);
and U8394 (N_8394,N_8261,N_8305);
or U8395 (N_8395,N_8259,N_8169);
xor U8396 (N_8396,N_8173,N_8284);
and U8397 (N_8397,N_8177,N_8235);
nor U8398 (N_8398,N_8171,N_8298);
xor U8399 (N_8399,N_8167,N_8178);
xnor U8400 (N_8400,N_8257,N_8243);
nand U8401 (N_8401,N_8292,N_8252);
and U8402 (N_8402,N_8242,N_8276);
nand U8403 (N_8403,N_8261,N_8160);
nand U8404 (N_8404,N_8315,N_8278);
nor U8405 (N_8405,N_8281,N_8273);
nor U8406 (N_8406,N_8173,N_8244);
nand U8407 (N_8407,N_8282,N_8188);
nor U8408 (N_8408,N_8276,N_8214);
nor U8409 (N_8409,N_8199,N_8295);
or U8410 (N_8410,N_8171,N_8194);
nor U8411 (N_8411,N_8179,N_8310);
nor U8412 (N_8412,N_8198,N_8167);
nor U8413 (N_8413,N_8186,N_8265);
nand U8414 (N_8414,N_8277,N_8214);
nand U8415 (N_8415,N_8316,N_8178);
nor U8416 (N_8416,N_8310,N_8199);
xor U8417 (N_8417,N_8160,N_8209);
and U8418 (N_8418,N_8191,N_8280);
nand U8419 (N_8419,N_8181,N_8240);
or U8420 (N_8420,N_8278,N_8279);
nor U8421 (N_8421,N_8260,N_8277);
nand U8422 (N_8422,N_8176,N_8175);
and U8423 (N_8423,N_8267,N_8189);
xnor U8424 (N_8424,N_8266,N_8235);
and U8425 (N_8425,N_8202,N_8186);
nand U8426 (N_8426,N_8223,N_8255);
or U8427 (N_8427,N_8236,N_8282);
and U8428 (N_8428,N_8181,N_8174);
or U8429 (N_8429,N_8226,N_8211);
and U8430 (N_8430,N_8269,N_8188);
xor U8431 (N_8431,N_8272,N_8202);
nand U8432 (N_8432,N_8165,N_8170);
nand U8433 (N_8433,N_8199,N_8245);
or U8434 (N_8434,N_8308,N_8202);
nand U8435 (N_8435,N_8257,N_8204);
nor U8436 (N_8436,N_8275,N_8316);
nor U8437 (N_8437,N_8293,N_8215);
xnor U8438 (N_8438,N_8310,N_8308);
xnor U8439 (N_8439,N_8169,N_8288);
nor U8440 (N_8440,N_8315,N_8311);
or U8441 (N_8441,N_8249,N_8307);
xnor U8442 (N_8442,N_8284,N_8281);
or U8443 (N_8443,N_8256,N_8293);
xnor U8444 (N_8444,N_8232,N_8171);
and U8445 (N_8445,N_8203,N_8257);
and U8446 (N_8446,N_8225,N_8167);
or U8447 (N_8447,N_8233,N_8291);
nor U8448 (N_8448,N_8189,N_8302);
xor U8449 (N_8449,N_8236,N_8193);
nand U8450 (N_8450,N_8224,N_8179);
nor U8451 (N_8451,N_8289,N_8220);
or U8452 (N_8452,N_8180,N_8235);
nor U8453 (N_8453,N_8275,N_8308);
xor U8454 (N_8454,N_8247,N_8316);
nor U8455 (N_8455,N_8236,N_8169);
and U8456 (N_8456,N_8208,N_8218);
nand U8457 (N_8457,N_8238,N_8219);
nor U8458 (N_8458,N_8314,N_8296);
nand U8459 (N_8459,N_8173,N_8222);
or U8460 (N_8460,N_8214,N_8263);
nor U8461 (N_8461,N_8276,N_8210);
and U8462 (N_8462,N_8243,N_8209);
nor U8463 (N_8463,N_8176,N_8298);
and U8464 (N_8464,N_8168,N_8243);
nor U8465 (N_8465,N_8318,N_8207);
xnor U8466 (N_8466,N_8248,N_8251);
xor U8467 (N_8467,N_8248,N_8188);
or U8468 (N_8468,N_8182,N_8188);
xor U8469 (N_8469,N_8291,N_8256);
nor U8470 (N_8470,N_8215,N_8160);
nand U8471 (N_8471,N_8307,N_8264);
and U8472 (N_8472,N_8274,N_8250);
or U8473 (N_8473,N_8184,N_8279);
and U8474 (N_8474,N_8282,N_8274);
nand U8475 (N_8475,N_8262,N_8215);
nand U8476 (N_8476,N_8273,N_8208);
or U8477 (N_8477,N_8239,N_8207);
or U8478 (N_8478,N_8177,N_8294);
nor U8479 (N_8479,N_8204,N_8290);
nor U8480 (N_8480,N_8459,N_8368);
xor U8481 (N_8481,N_8466,N_8420);
or U8482 (N_8482,N_8446,N_8355);
and U8483 (N_8483,N_8476,N_8427);
nand U8484 (N_8484,N_8408,N_8340);
xor U8485 (N_8485,N_8469,N_8346);
xnor U8486 (N_8486,N_8383,N_8396);
nor U8487 (N_8487,N_8364,N_8325);
nand U8488 (N_8488,N_8438,N_8333);
nand U8489 (N_8489,N_8419,N_8472);
nor U8490 (N_8490,N_8330,N_8341);
xor U8491 (N_8491,N_8357,N_8415);
and U8492 (N_8492,N_8457,N_8445);
xnor U8493 (N_8493,N_8462,N_8380);
xor U8494 (N_8494,N_8451,N_8455);
xnor U8495 (N_8495,N_8371,N_8361);
xnor U8496 (N_8496,N_8393,N_8414);
nor U8497 (N_8497,N_8407,N_8477);
nand U8498 (N_8498,N_8406,N_8337);
or U8499 (N_8499,N_8391,N_8378);
nand U8500 (N_8500,N_8342,N_8323);
xnor U8501 (N_8501,N_8475,N_8373);
xor U8502 (N_8502,N_8422,N_8335);
and U8503 (N_8503,N_8426,N_8334);
and U8504 (N_8504,N_8351,N_8344);
nand U8505 (N_8505,N_8448,N_8470);
nand U8506 (N_8506,N_8439,N_8417);
nor U8507 (N_8507,N_8348,N_8353);
and U8508 (N_8508,N_8444,N_8442);
xor U8509 (N_8509,N_8405,N_8392);
nand U8510 (N_8510,N_8404,N_8394);
nand U8511 (N_8511,N_8366,N_8349);
nor U8512 (N_8512,N_8377,N_8435);
nor U8513 (N_8513,N_8436,N_8395);
xor U8514 (N_8514,N_8367,N_8345);
xor U8515 (N_8515,N_8429,N_8379);
and U8516 (N_8516,N_8360,N_8376);
nand U8517 (N_8517,N_8467,N_8372);
nand U8518 (N_8518,N_8397,N_8339);
or U8519 (N_8519,N_8464,N_8416);
nand U8520 (N_8520,N_8398,N_8437);
nand U8521 (N_8521,N_8369,N_8441);
xor U8522 (N_8522,N_8460,N_8329);
or U8523 (N_8523,N_8458,N_8425);
xnor U8524 (N_8524,N_8385,N_8389);
nor U8525 (N_8525,N_8365,N_8479);
and U8526 (N_8526,N_8375,N_8399);
or U8527 (N_8527,N_8418,N_8387);
and U8528 (N_8528,N_8463,N_8363);
nand U8529 (N_8529,N_8326,N_8450);
xor U8530 (N_8530,N_8322,N_8402);
and U8531 (N_8531,N_8386,N_8324);
and U8532 (N_8532,N_8382,N_8424);
or U8533 (N_8533,N_8358,N_8440);
and U8534 (N_8534,N_8343,N_8447);
nor U8535 (N_8535,N_8328,N_8411);
nand U8536 (N_8536,N_8362,N_8433);
nor U8537 (N_8537,N_8474,N_8413);
nor U8538 (N_8538,N_8320,N_8352);
xor U8539 (N_8539,N_8390,N_8384);
or U8540 (N_8540,N_8468,N_8434);
or U8541 (N_8541,N_8410,N_8347);
nor U8542 (N_8542,N_8428,N_8409);
nand U8543 (N_8543,N_8461,N_8478);
nand U8544 (N_8544,N_8388,N_8370);
and U8545 (N_8545,N_8431,N_8374);
xor U8546 (N_8546,N_8403,N_8401);
xnor U8547 (N_8547,N_8332,N_8465);
nand U8548 (N_8548,N_8354,N_8452);
and U8549 (N_8549,N_8473,N_8449);
nand U8550 (N_8550,N_8321,N_8359);
or U8551 (N_8551,N_8350,N_8456);
or U8552 (N_8552,N_8454,N_8336);
and U8553 (N_8553,N_8381,N_8432);
and U8554 (N_8554,N_8421,N_8338);
nor U8555 (N_8555,N_8423,N_8453);
or U8556 (N_8556,N_8331,N_8430);
and U8557 (N_8557,N_8400,N_8443);
xor U8558 (N_8558,N_8412,N_8471);
nand U8559 (N_8559,N_8356,N_8327);
nor U8560 (N_8560,N_8472,N_8383);
nor U8561 (N_8561,N_8323,N_8477);
nor U8562 (N_8562,N_8335,N_8472);
nand U8563 (N_8563,N_8413,N_8412);
xnor U8564 (N_8564,N_8353,N_8327);
and U8565 (N_8565,N_8359,N_8461);
and U8566 (N_8566,N_8368,N_8411);
and U8567 (N_8567,N_8440,N_8379);
or U8568 (N_8568,N_8449,N_8373);
xor U8569 (N_8569,N_8354,N_8366);
and U8570 (N_8570,N_8456,N_8448);
or U8571 (N_8571,N_8448,N_8406);
and U8572 (N_8572,N_8451,N_8379);
and U8573 (N_8573,N_8378,N_8351);
and U8574 (N_8574,N_8464,N_8421);
nand U8575 (N_8575,N_8441,N_8378);
xnor U8576 (N_8576,N_8347,N_8346);
nor U8577 (N_8577,N_8386,N_8438);
nand U8578 (N_8578,N_8371,N_8428);
and U8579 (N_8579,N_8467,N_8361);
xnor U8580 (N_8580,N_8399,N_8426);
or U8581 (N_8581,N_8430,N_8326);
or U8582 (N_8582,N_8331,N_8386);
xor U8583 (N_8583,N_8407,N_8426);
or U8584 (N_8584,N_8331,N_8323);
and U8585 (N_8585,N_8350,N_8420);
nor U8586 (N_8586,N_8375,N_8389);
xor U8587 (N_8587,N_8399,N_8345);
nand U8588 (N_8588,N_8450,N_8437);
nand U8589 (N_8589,N_8412,N_8389);
and U8590 (N_8590,N_8476,N_8390);
nand U8591 (N_8591,N_8365,N_8394);
or U8592 (N_8592,N_8375,N_8400);
nor U8593 (N_8593,N_8352,N_8344);
or U8594 (N_8594,N_8418,N_8456);
nand U8595 (N_8595,N_8359,N_8325);
and U8596 (N_8596,N_8359,N_8361);
or U8597 (N_8597,N_8478,N_8350);
nor U8598 (N_8598,N_8445,N_8432);
and U8599 (N_8599,N_8329,N_8368);
or U8600 (N_8600,N_8438,N_8334);
or U8601 (N_8601,N_8452,N_8350);
nor U8602 (N_8602,N_8422,N_8381);
or U8603 (N_8603,N_8410,N_8439);
and U8604 (N_8604,N_8377,N_8428);
xor U8605 (N_8605,N_8350,N_8429);
and U8606 (N_8606,N_8375,N_8476);
nand U8607 (N_8607,N_8390,N_8465);
or U8608 (N_8608,N_8345,N_8339);
and U8609 (N_8609,N_8477,N_8341);
or U8610 (N_8610,N_8469,N_8408);
or U8611 (N_8611,N_8418,N_8402);
and U8612 (N_8612,N_8345,N_8425);
nand U8613 (N_8613,N_8464,N_8379);
nand U8614 (N_8614,N_8470,N_8468);
or U8615 (N_8615,N_8374,N_8369);
nor U8616 (N_8616,N_8322,N_8470);
and U8617 (N_8617,N_8413,N_8408);
xor U8618 (N_8618,N_8429,N_8428);
or U8619 (N_8619,N_8452,N_8407);
nor U8620 (N_8620,N_8451,N_8383);
nor U8621 (N_8621,N_8428,N_8376);
xnor U8622 (N_8622,N_8404,N_8372);
and U8623 (N_8623,N_8378,N_8458);
nor U8624 (N_8624,N_8448,N_8399);
xnor U8625 (N_8625,N_8424,N_8369);
nand U8626 (N_8626,N_8339,N_8391);
nand U8627 (N_8627,N_8338,N_8398);
xor U8628 (N_8628,N_8398,N_8376);
xnor U8629 (N_8629,N_8347,N_8437);
xnor U8630 (N_8630,N_8384,N_8343);
nor U8631 (N_8631,N_8358,N_8357);
and U8632 (N_8632,N_8433,N_8423);
and U8633 (N_8633,N_8395,N_8378);
or U8634 (N_8634,N_8406,N_8353);
nor U8635 (N_8635,N_8428,N_8362);
nor U8636 (N_8636,N_8345,N_8414);
xnor U8637 (N_8637,N_8328,N_8351);
xnor U8638 (N_8638,N_8465,N_8377);
and U8639 (N_8639,N_8437,N_8352);
and U8640 (N_8640,N_8505,N_8488);
nand U8641 (N_8641,N_8545,N_8597);
nor U8642 (N_8642,N_8577,N_8602);
and U8643 (N_8643,N_8626,N_8619);
and U8644 (N_8644,N_8503,N_8537);
or U8645 (N_8645,N_8557,N_8482);
and U8646 (N_8646,N_8535,N_8539);
nand U8647 (N_8647,N_8570,N_8573);
nand U8648 (N_8648,N_8563,N_8636);
or U8649 (N_8649,N_8523,N_8507);
nor U8650 (N_8650,N_8554,N_8498);
nor U8651 (N_8651,N_8632,N_8534);
or U8652 (N_8652,N_8631,N_8603);
xnor U8653 (N_8653,N_8611,N_8569);
nand U8654 (N_8654,N_8559,N_8547);
and U8655 (N_8655,N_8514,N_8500);
and U8656 (N_8656,N_8591,N_8628);
nor U8657 (N_8657,N_8524,N_8624);
nor U8658 (N_8658,N_8553,N_8578);
xnor U8659 (N_8659,N_8574,N_8564);
nand U8660 (N_8660,N_8484,N_8502);
nand U8661 (N_8661,N_8594,N_8606);
nand U8662 (N_8662,N_8561,N_8634);
and U8663 (N_8663,N_8627,N_8584);
xor U8664 (N_8664,N_8635,N_8623);
and U8665 (N_8665,N_8549,N_8633);
nor U8666 (N_8666,N_8552,N_8616);
nor U8667 (N_8667,N_8519,N_8504);
xnor U8668 (N_8668,N_8568,N_8579);
and U8669 (N_8669,N_8497,N_8565);
nor U8670 (N_8670,N_8586,N_8583);
nor U8671 (N_8671,N_8637,N_8639);
xnor U8672 (N_8672,N_8609,N_8527);
xnor U8673 (N_8673,N_8489,N_8520);
and U8674 (N_8674,N_8571,N_8620);
or U8675 (N_8675,N_8582,N_8575);
xor U8676 (N_8676,N_8576,N_8618);
nor U8677 (N_8677,N_8542,N_8533);
and U8678 (N_8678,N_8610,N_8560);
nand U8679 (N_8679,N_8487,N_8496);
nand U8680 (N_8680,N_8546,N_8581);
or U8681 (N_8681,N_8490,N_8567);
and U8682 (N_8682,N_8585,N_8607);
and U8683 (N_8683,N_8543,N_8532);
or U8684 (N_8684,N_8529,N_8521);
and U8685 (N_8685,N_8601,N_8555);
and U8686 (N_8686,N_8558,N_8528);
xor U8687 (N_8687,N_8483,N_8516);
xor U8688 (N_8688,N_8518,N_8599);
and U8689 (N_8689,N_8481,N_8511);
and U8690 (N_8690,N_8536,N_8589);
and U8691 (N_8691,N_8492,N_8508);
nor U8692 (N_8692,N_8526,N_8501);
xor U8693 (N_8693,N_8617,N_8608);
or U8694 (N_8694,N_8538,N_8614);
and U8695 (N_8695,N_8486,N_8515);
nand U8696 (N_8696,N_8604,N_8598);
or U8697 (N_8697,N_8621,N_8592);
nand U8698 (N_8698,N_8629,N_8531);
xor U8699 (N_8699,N_8550,N_8513);
nand U8700 (N_8700,N_8605,N_8541);
xor U8701 (N_8701,N_8600,N_8525);
and U8702 (N_8702,N_8480,N_8580);
and U8703 (N_8703,N_8517,N_8587);
xor U8704 (N_8704,N_8593,N_8551);
nand U8705 (N_8705,N_8615,N_8566);
nor U8706 (N_8706,N_8556,N_8622);
xor U8707 (N_8707,N_8595,N_8506);
xor U8708 (N_8708,N_8491,N_8596);
or U8709 (N_8709,N_8485,N_8540);
or U8710 (N_8710,N_8613,N_8499);
and U8711 (N_8711,N_8572,N_8612);
nor U8712 (N_8712,N_8509,N_8493);
nor U8713 (N_8713,N_8522,N_8495);
nor U8714 (N_8714,N_8590,N_8530);
or U8715 (N_8715,N_8625,N_8638);
or U8716 (N_8716,N_8510,N_8630);
or U8717 (N_8717,N_8562,N_8512);
or U8718 (N_8718,N_8544,N_8548);
nor U8719 (N_8719,N_8588,N_8494);
and U8720 (N_8720,N_8613,N_8620);
nand U8721 (N_8721,N_8556,N_8514);
nand U8722 (N_8722,N_8609,N_8524);
or U8723 (N_8723,N_8596,N_8493);
or U8724 (N_8724,N_8501,N_8484);
and U8725 (N_8725,N_8544,N_8637);
nand U8726 (N_8726,N_8503,N_8556);
xor U8727 (N_8727,N_8487,N_8489);
and U8728 (N_8728,N_8598,N_8544);
or U8729 (N_8729,N_8609,N_8495);
nor U8730 (N_8730,N_8493,N_8586);
or U8731 (N_8731,N_8624,N_8567);
xnor U8732 (N_8732,N_8617,N_8638);
xor U8733 (N_8733,N_8484,N_8525);
and U8734 (N_8734,N_8610,N_8591);
or U8735 (N_8735,N_8547,N_8500);
nor U8736 (N_8736,N_8607,N_8548);
or U8737 (N_8737,N_8513,N_8521);
and U8738 (N_8738,N_8600,N_8599);
xnor U8739 (N_8739,N_8623,N_8599);
nand U8740 (N_8740,N_8582,N_8588);
xnor U8741 (N_8741,N_8605,N_8521);
and U8742 (N_8742,N_8548,N_8525);
or U8743 (N_8743,N_8586,N_8595);
or U8744 (N_8744,N_8583,N_8489);
and U8745 (N_8745,N_8638,N_8540);
nand U8746 (N_8746,N_8511,N_8627);
nor U8747 (N_8747,N_8497,N_8629);
nand U8748 (N_8748,N_8539,N_8586);
or U8749 (N_8749,N_8622,N_8518);
nor U8750 (N_8750,N_8639,N_8621);
nor U8751 (N_8751,N_8603,N_8535);
nand U8752 (N_8752,N_8564,N_8605);
or U8753 (N_8753,N_8547,N_8567);
xnor U8754 (N_8754,N_8572,N_8586);
and U8755 (N_8755,N_8567,N_8525);
nand U8756 (N_8756,N_8511,N_8639);
and U8757 (N_8757,N_8625,N_8512);
xor U8758 (N_8758,N_8551,N_8562);
or U8759 (N_8759,N_8564,N_8543);
nand U8760 (N_8760,N_8557,N_8484);
nor U8761 (N_8761,N_8545,N_8609);
nor U8762 (N_8762,N_8489,N_8524);
and U8763 (N_8763,N_8523,N_8569);
or U8764 (N_8764,N_8542,N_8593);
and U8765 (N_8765,N_8531,N_8588);
or U8766 (N_8766,N_8603,N_8496);
xor U8767 (N_8767,N_8486,N_8599);
and U8768 (N_8768,N_8531,N_8539);
nor U8769 (N_8769,N_8560,N_8488);
nor U8770 (N_8770,N_8572,N_8631);
nor U8771 (N_8771,N_8529,N_8593);
nand U8772 (N_8772,N_8599,N_8529);
xnor U8773 (N_8773,N_8626,N_8509);
or U8774 (N_8774,N_8573,N_8534);
nor U8775 (N_8775,N_8494,N_8570);
nor U8776 (N_8776,N_8590,N_8563);
xor U8777 (N_8777,N_8534,N_8569);
or U8778 (N_8778,N_8481,N_8598);
nand U8779 (N_8779,N_8505,N_8591);
or U8780 (N_8780,N_8556,N_8559);
or U8781 (N_8781,N_8627,N_8544);
xnor U8782 (N_8782,N_8628,N_8639);
nand U8783 (N_8783,N_8575,N_8628);
and U8784 (N_8784,N_8600,N_8632);
xnor U8785 (N_8785,N_8581,N_8528);
and U8786 (N_8786,N_8487,N_8591);
xnor U8787 (N_8787,N_8510,N_8632);
and U8788 (N_8788,N_8613,N_8604);
nor U8789 (N_8789,N_8531,N_8608);
nand U8790 (N_8790,N_8525,N_8591);
xor U8791 (N_8791,N_8616,N_8521);
xor U8792 (N_8792,N_8575,N_8568);
or U8793 (N_8793,N_8581,N_8485);
or U8794 (N_8794,N_8521,N_8637);
or U8795 (N_8795,N_8514,N_8528);
xor U8796 (N_8796,N_8582,N_8486);
nor U8797 (N_8797,N_8489,N_8555);
xor U8798 (N_8798,N_8525,N_8603);
xor U8799 (N_8799,N_8519,N_8483);
or U8800 (N_8800,N_8712,N_8754);
nor U8801 (N_8801,N_8716,N_8696);
or U8802 (N_8802,N_8644,N_8679);
and U8803 (N_8803,N_8643,N_8650);
nand U8804 (N_8804,N_8738,N_8792);
nor U8805 (N_8805,N_8705,N_8749);
or U8806 (N_8806,N_8688,N_8651);
and U8807 (N_8807,N_8704,N_8669);
nor U8808 (N_8808,N_8717,N_8732);
nand U8809 (N_8809,N_8706,N_8791);
nor U8810 (N_8810,N_8740,N_8769);
nor U8811 (N_8811,N_8790,N_8694);
nand U8812 (N_8812,N_8736,N_8662);
and U8813 (N_8813,N_8693,N_8797);
nand U8814 (N_8814,N_8730,N_8780);
or U8815 (N_8815,N_8698,N_8686);
nand U8816 (N_8816,N_8645,N_8655);
nor U8817 (N_8817,N_8786,N_8642);
nor U8818 (N_8818,N_8683,N_8659);
nor U8819 (N_8819,N_8670,N_8793);
nand U8820 (N_8820,N_8702,N_8776);
xnor U8821 (N_8821,N_8646,N_8667);
and U8822 (N_8822,N_8710,N_8666);
nor U8823 (N_8823,N_8779,N_8729);
or U8824 (N_8824,N_8671,N_8746);
nand U8825 (N_8825,N_8684,N_8789);
and U8826 (N_8826,N_8751,N_8763);
or U8827 (N_8827,N_8747,N_8660);
or U8828 (N_8828,N_8759,N_8703);
nand U8829 (N_8829,N_8741,N_8772);
or U8830 (N_8830,N_8678,N_8725);
xor U8831 (N_8831,N_8709,N_8652);
and U8832 (N_8832,N_8734,N_8653);
nor U8833 (N_8833,N_8681,N_8782);
xnor U8834 (N_8834,N_8714,N_8675);
or U8835 (N_8835,N_8723,N_8673);
xor U8836 (N_8836,N_8784,N_8720);
nand U8837 (N_8837,N_8695,N_8798);
nand U8838 (N_8838,N_8743,N_8718);
xnor U8839 (N_8839,N_8777,N_8724);
nand U8840 (N_8840,N_8762,N_8713);
and U8841 (N_8841,N_8689,N_8750);
nand U8842 (N_8842,N_8726,N_8752);
nand U8843 (N_8843,N_8727,N_8641);
and U8844 (N_8844,N_8745,N_8640);
xor U8845 (N_8845,N_8768,N_8672);
nor U8846 (N_8846,N_8766,N_8700);
nand U8847 (N_8847,N_8680,N_8707);
nor U8848 (N_8848,N_8665,N_8661);
or U8849 (N_8849,N_8756,N_8711);
nor U8850 (N_8850,N_8663,N_8674);
or U8851 (N_8851,N_8760,N_8757);
or U8852 (N_8852,N_8722,N_8656);
xnor U8853 (N_8853,N_8647,N_8691);
and U8854 (N_8854,N_8778,N_8649);
nor U8855 (N_8855,N_8676,N_8735);
nor U8856 (N_8856,N_8733,N_8748);
nor U8857 (N_8857,N_8654,N_8682);
and U8858 (N_8858,N_8731,N_8677);
nor U8859 (N_8859,N_8690,N_8657);
and U8860 (N_8860,N_8701,N_8648);
nor U8861 (N_8861,N_8781,N_8697);
xor U8862 (N_8862,N_8715,N_8767);
xor U8863 (N_8863,N_8719,N_8788);
or U8864 (N_8864,N_8770,N_8708);
nor U8865 (N_8865,N_8742,N_8783);
or U8866 (N_8866,N_8664,N_8737);
xnor U8867 (N_8867,N_8771,N_8687);
or U8868 (N_8868,N_8685,N_8794);
nor U8869 (N_8869,N_8758,N_8799);
xor U8870 (N_8870,N_8774,N_8753);
and U8871 (N_8871,N_8795,N_8796);
or U8872 (N_8872,N_8744,N_8764);
and U8873 (N_8873,N_8739,N_8699);
and U8874 (N_8874,N_8668,N_8787);
and U8875 (N_8875,N_8721,N_8773);
xor U8876 (N_8876,N_8765,N_8775);
and U8877 (N_8877,N_8692,N_8658);
and U8878 (N_8878,N_8728,N_8761);
xor U8879 (N_8879,N_8755,N_8785);
xnor U8880 (N_8880,N_8709,N_8672);
and U8881 (N_8881,N_8764,N_8790);
nand U8882 (N_8882,N_8643,N_8773);
or U8883 (N_8883,N_8754,N_8762);
or U8884 (N_8884,N_8691,N_8757);
and U8885 (N_8885,N_8753,N_8698);
and U8886 (N_8886,N_8651,N_8760);
nor U8887 (N_8887,N_8759,N_8673);
xnor U8888 (N_8888,N_8764,N_8694);
and U8889 (N_8889,N_8640,N_8642);
xor U8890 (N_8890,N_8713,N_8742);
or U8891 (N_8891,N_8745,N_8753);
or U8892 (N_8892,N_8774,N_8732);
nand U8893 (N_8893,N_8770,N_8794);
nand U8894 (N_8894,N_8748,N_8676);
nand U8895 (N_8895,N_8640,N_8654);
and U8896 (N_8896,N_8669,N_8710);
nand U8897 (N_8897,N_8784,N_8690);
nand U8898 (N_8898,N_8640,N_8668);
or U8899 (N_8899,N_8642,N_8687);
and U8900 (N_8900,N_8758,N_8739);
xnor U8901 (N_8901,N_8653,N_8708);
xnor U8902 (N_8902,N_8688,N_8658);
nor U8903 (N_8903,N_8706,N_8669);
or U8904 (N_8904,N_8672,N_8689);
or U8905 (N_8905,N_8680,N_8676);
or U8906 (N_8906,N_8784,N_8662);
and U8907 (N_8907,N_8697,N_8793);
and U8908 (N_8908,N_8700,N_8763);
xor U8909 (N_8909,N_8677,N_8688);
nor U8910 (N_8910,N_8777,N_8699);
or U8911 (N_8911,N_8656,N_8672);
and U8912 (N_8912,N_8742,N_8796);
nor U8913 (N_8913,N_8696,N_8668);
nor U8914 (N_8914,N_8771,N_8763);
xnor U8915 (N_8915,N_8792,N_8698);
xnor U8916 (N_8916,N_8643,N_8760);
or U8917 (N_8917,N_8735,N_8770);
and U8918 (N_8918,N_8661,N_8775);
nor U8919 (N_8919,N_8668,N_8738);
or U8920 (N_8920,N_8720,N_8695);
and U8921 (N_8921,N_8791,N_8673);
nand U8922 (N_8922,N_8677,N_8664);
and U8923 (N_8923,N_8735,N_8771);
nand U8924 (N_8924,N_8755,N_8680);
nand U8925 (N_8925,N_8684,N_8651);
or U8926 (N_8926,N_8704,N_8741);
xnor U8927 (N_8927,N_8645,N_8782);
and U8928 (N_8928,N_8793,N_8677);
or U8929 (N_8929,N_8646,N_8743);
and U8930 (N_8930,N_8747,N_8682);
nand U8931 (N_8931,N_8687,N_8710);
nor U8932 (N_8932,N_8650,N_8750);
nor U8933 (N_8933,N_8739,N_8786);
or U8934 (N_8934,N_8717,N_8714);
and U8935 (N_8935,N_8717,N_8678);
nand U8936 (N_8936,N_8697,N_8758);
xnor U8937 (N_8937,N_8698,N_8715);
nand U8938 (N_8938,N_8739,N_8732);
nand U8939 (N_8939,N_8736,N_8730);
nand U8940 (N_8940,N_8690,N_8680);
and U8941 (N_8941,N_8678,N_8673);
or U8942 (N_8942,N_8770,N_8713);
nand U8943 (N_8943,N_8670,N_8739);
xor U8944 (N_8944,N_8680,N_8746);
nand U8945 (N_8945,N_8788,N_8779);
nor U8946 (N_8946,N_8796,N_8731);
nor U8947 (N_8947,N_8722,N_8739);
xor U8948 (N_8948,N_8738,N_8750);
and U8949 (N_8949,N_8659,N_8720);
nor U8950 (N_8950,N_8795,N_8669);
nor U8951 (N_8951,N_8689,N_8742);
nor U8952 (N_8952,N_8753,N_8667);
nand U8953 (N_8953,N_8653,N_8659);
and U8954 (N_8954,N_8764,N_8704);
and U8955 (N_8955,N_8662,N_8711);
nand U8956 (N_8956,N_8715,N_8774);
and U8957 (N_8957,N_8645,N_8770);
or U8958 (N_8958,N_8795,N_8642);
nor U8959 (N_8959,N_8771,N_8690);
or U8960 (N_8960,N_8922,N_8953);
nand U8961 (N_8961,N_8896,N_8852);
or U8962 (N_8962,N_8804,N_8828);
and U8963 (N_8963,N_8865,N_8917);
and U8964 (N_8964,N_8802,N_8809);
xor U8965 (N_8965,N_8807,N_8925);
xnor U8966 (N_8966,N_8803,N_8823);
and U8967 (N_8967,N_8949,N_8891);
xnor U8968 (N_8968,N_8816,N_8857);
nor U8969 (N_8969,N_8872,N_8842);
xnor U8970 (N_8970,N_8819,N_8950);
nand U8971 (N_8971,N_8951,N_8892);
xor U8972 (N_8972,N_8943,N_8874);
xnor U8973 (N_8973,N_8859,N_8937);
nor U8974 (N_8974,N_8879,N_8924);
or U8975 (N_8975,N_8878,N_8821);
and U8976 (N_8976,N_8936,N_8866);
and U8977 (N_8977,N_8831,N_8938);
and U8978 (N_8978,N_8840,N_8808);
and U8979 (N_8979,N_8800,N_8863);
xnor U8980 (N_8980,N_8905,N_8815);
or U8981 (N_8981,N_8884,N_8914);
nor U8982 (N_8982,N_8806,N_8880);
and U8983 (N_8983,N_8837,N_8813);
or U8984 (N_8984,N_8944,N_8919);
nand U8985 (N_8985,N_8945,N_8812);
and U8986 (N_8986,N_8861,N_8886);
and U8987 (N_8987,N_8895,N_8824);
or U8988 (N_8988,N_8894,N_8834);
nor U8989 (N_8989,N_8829,N_8948);
or U8990 (N_8990,N_8830,N_8959);
and U8991 (N_8991,N_8864,N_8875);
nand U8992 (N_8992,N_8897,N_8844);
xor U8993 (N_8993,N_8860,N_8934);
xor U8994 (N_8994,N_8820,N_8923);
or U8995 (N_8995,N_8877,N_8855);
nand U8996 (N_8996,N_8890,N_8825);
nand U8997 (N_8997,N_8918,N_8915);
and U8998 (N_8998,N_8929,N_8900);
nor U8999 (N_8999,N_8827,N_8843);
xor U9000 (N_9000,N_8931,N_8835);
and U9001 (N_9001,N_8871,N_8957);
or U9002 (N_9002,N_8933,N_8913);
xor U9003 (N_9003,N_8836,N_8881);
xor U9004 (N_9004,N_8869,N_8942);
nor U9005 (N_9005,N_8862,N_8845);
xnor U9006 (N_9006,N_8870,N_8805);
and U9007 (N_9007,N_8926,N_8930);
and U9008 (N_9008,N_8903,N_8851);
xnor U9009 (N_9009,N_8946,N_8906);
and U9010 (N_9010,N_8882,N_8801);
nand U9011 (N_9011,N_8958,N_8814);
xor U9012 (N_9012,N_8873,N_8912);
or U9013 (N_9013,N_8940,N_8899);
or U9014 (N_9014,N_8955,N_8904);
and U9015 (N_9015,N_8888,N_8818);
nor U9016 (N_9016,N_8954,N_8952);
nand U9017 (N_9017,N_8921,N_8928);
nor U9018 (N_9018,N_8932,N_8889);
xor U9019 (N_9019,N_8856,N_8817);
nand U9020 (N_9020,N_8841,N_8893);
nor U9021 (N_9021,N_8811,N_8887);
and U9022 (N_9022,N_8839,N_8838);
xor U9023 (N_9023,N_8853,N_8907);
or U9024 (N_9024,N_8810,N_8898);
and U9025 (N_9025,N_8902,N_8846);
xnor U9026 (N_9026,N_8833,N_8868);
nand U9027 (N_9027,N_8927,N_8822);
nor U9028 (N_9028,N_8901,N_8947);
or U9029 (N_9029,N_8858,N_8911);
xor U9030 (N_9030,N_8909,N_8867);
or U9031 (N_9031,N_8849,N_8876);
and U9032 (N_9032,N_8941,N_8848);
or U9033 (N_9033,N_8832,N_8920);
and U9034 (N_9034,N_8908,N_8826);
and U9035 (N_9035,N_8939,N_8910);
nand U9036 (N_9036,N_8854,N_8916);
and U9037 (N_9037,N_8850,N_8885);
nand U9038 (N_9038,N_8935,N_8883);
xor U9039 (N_9039,N_8956,N_8847);
and U9040 (N_9040,N_8843,N_8865);
or U9041 (N_9041,N_8802,N_8829);
nor U9042 (N_9042,N_8918,N_8866);
and U9043 (N_9043,N_8885,N_8927);
or U9044 (N_9044,N_8912,N_8879);
or U9045 (N_9045,N_8916,N_8820);
nand U9046 (N_9046,N_8881,N_8854);
or U9047 (N_9047,N_8913,N_8817);
xnor U9048 (N_9048,N_8848,N_8888);
nand U9049 (N_9049,N_8866,N_8911);
or U9050 (N_9050,N_8837,N_8913);
xnor U9051 (N_9051,N_8851,N_8831);
nand U9052 (N_9052,N_8943,N_8921);
and U9053 (N_9053,N_8800,N_8878);
nand U9054 (N_9054,N_8870,N_8903);
xor U9055 (N_9055,N_8937,N_8887);
or U9056 (N_9056,N_8842,N_8940);
nand U9057 (N_9057,N_8844,N_8869);
nor U9058 (N_9058,N_8910,N_8847);
nand U9059 (N_9059,N_8804,N_8820);
or U9060 (N_9060,N_8880,N_8887);
nand U9061 (N_9061,N_8900,N_8958);
xor U9062 (N_9062,N_8869,N_8883);
nand U9063 (N_9063,N_8922,N_8942);
xnor U9064 (N_9064,N_8873,N_8820);
nor U9065 (N_9065,N_8897,N_8816);
xor U9066 (N_9066,N_8910,N_8852);
nor U9067 (N_9067,N_8939,N_8899);
nand U9068 (N_9068,N_8829,N_8833);
nor U9069 (N_9069,N_8915,N_8927);
and U9070 (N_9070,N_8914,N_8810);
or U9071 (N_9071,N_8888,N_8926);
and U9072 (N_9072,N_8824,N_8802);
xor U9073 (N_9073,N_8948,N_8839);
or U9074 (N_9074,N_8830,N_8835);
xor U9075 (N_9075,N_8839,N_8869);
xor U9076 (N_9076,N_8821,N_8894);
or U9077 (N_9077,N_8953,N_8841);
nor U9078 (N_9078,N_8835,N_8948);
nand U9079 (N_9079,N_8927,N_8835);
nand U9080 (N_9080,N_8811,N_8959);
or U9081 (N_9081,N_8936,N_8872);
nand U9082 (N_9082,N_8857,N_8941);
nor U9083 (N_9083,N_8831,N_8957);
nand U9084 (N_9084,N_8845,N_8848);
or U9085 (N_9085,N_8843,N_8862);
nor U9086 (N_9086,N_8899,N_8814);
and U9087 (N_9087,N_8837,N_8875);
and U9088 (N_9088,N_8933,N_8862);
xnor U9089 (N_9089,N_8938,N_8803);
nand U9090 (N_9090,N_8850,N_8901);
nor U9091 (N_9091,N_8863,N_8816);
and U9092 (N_9092,N_8856,N_8909);
xor U9093 (N_9093,N_8908,N_8916);
and U9094 (N_9094,N_8869,N_8932);
or U9095 (N_9095,N_8813,N_8811);
xnor U9096 (N_9096,N_8872,N_8810);
xnor U9097 (N_9097,N_8926,N_8907);
nor U9098 (N_9098,N_8893,N_8957);
or U9099 (N_9099,N_8948,N_8865);
and U9100 (N_9100,N_8824,N_8917);
and U9101 (N_9101,N_8953,N_8931);
and U9102 (N_9102,N_8866,N_8883);
nor U9103 (N_9103,N_8904,N_8824);
xnor U9104 (N_9104,N_8848,N_8807);
and U9105 (N_9105,N_8829,N_8904);
and U9106 (N_9106,N_8853,N_8833);
nor U9107 (N_9107,N_8825,N_8858);
nand U9108 (N_9108,N_8853,N_8930);
and U9109 (N_9109,N_8911,N_8820);
xnor U9110 (N_9110,N_8882,N_8940);
or U9111 (N_9111,N_8929,N_8864);
xor U9112 (N_9112,N_8926,N_8937);
nand U9113 (N_9113,N_8942,N_8927);
nand U9114 (N_9114,N_8895,N_8943);
nand U9115 (N_9115,N_8944,N_8874);
or U9116 (N_9116,N_8814,N_8801);
or U9117 (N_9117,N_8872,N_8919);
xnor U9118 (N_9118,N_8906,N_8803);
nor U9119 (N_9119,N_8939,N_8859);
and U9120 (N_9120,N_8985,N_8988);
nand U9121 (N_9121,N_9037,N_8986);
nand U9122 (N_9122,N_9102,N_9110);
nor U9123 (N_9123,N_9104,N_9117);
and U9124 (N_9124,N_8977,N_9028);
or U9125 (N_9125,N_9036,N_9054);
xnor U9126 (N_9126,N_9023,N_9013);
nor U9127 (N_9127,N_9017,N_9079);
nand U9128 (N_9128,N_8997,N_8970);
nor U9129 (N_9129,N_9097,N_8978);
or U9130 (N_9130,N_8965,N_9083);
or U9131 (N_9131,N_9098,N_9111);
and U9132 (N_9132,N_9066,N_9020);
and U9133 (N_9133,N_9100,N_9015);
and U9134 (N_9134,N_9034,N_8982);
nand U9135 (N_9135,N_9062,N_9065);
and U9136 (N_9136,N_9118,N_8960);
nand U9137 (N_9137,N_9063,N_8975);
or U9138 (N_9138,N_9059,N_9086);
or U9139 (N_9139,N_9087,N_8994);
nor U9140 (N_9140,N_8974,N_9090);
and U9141 (N_9141,N_9000,N_9095);
nor U9142 (N_9142,N_8981,N_9107);
or U9143 (N_9143,N_9115,N_9113);
or U9144 (N_9144,N_9002,N_8996);
nor U9145 (N_9145,N_9004,N_9003);
nor U9146 (N_9146,N_9119,N_9024);
and U9147 (N_9147,N_9045,N_8967);
xor U9148 (N_9148,N_8969,N_8998);
nor U9149 (N_9149,N_9016,N_8971);
and U9150 (N_9150,N_8976,N_9075);
or U9151 (N_9151,N_8968,N_8993);
and U9152 (N_9152,N_9051,N_9096);
and U9153 (N_9153,N_8989,N_8991);
and U9154 (N_9154,N_9012,N_9052);
and U9155 (N_9155,N_9006,N_9099);
nand U9156 (N_9156,N_9088,N_9008);
xor U9157 (N_9157,N_9085,N_9026);
and U9158 (N_9158,N_9009,N_9093);
and U9159 (N_9159,N_9071,N_9082);
xnor U9160 (N_9160,N_9007,N_8983);
nor U9161 (N_9161,N_9030,N_9040);
xnor U9162 (N_9162,N_8999,N_9072);
xor U9163 (N_9163,N_9035,N_9101);
and U9164 (N_9164,N_8966,N_9080);
nand U9165 (N_9165,N_9010,N_9060);
nand U9166 (N_9166,N_9029,N_8980);
nor U9167 (N_9167,N_9057,N_9055);
nor U9168 (N_9168,N_8987,N_9081);
nand U9169 (N_9169,N_8962,N_9074);
nor U9170 (N_9170,N_8963,N_8995);
or U9171 (N_9171,N_9044,N_9043);
nand U9172 (N_9172,N_9073,N_9031);
nand U9173 (N_9173,N_9061,N_8984);
nor U9174 (N_9174,N_9070,N_9032);
and U9175 (N_9175,N_9116,N_9038);
and U9176 (N_9176,N_9112,N_9039);
nor U9177 (N_9177,N_9018,N_9022);
xnor U9178 (N_9178,N_9011,N_9091);
nor U9179 (N_9179,N_9047,N_9001);
xnor U9180 (N_9180,N_9084,N_9076);
or U9181 (N_9181,N_9114,N_9068);
nand U9182 (N_9182,N_9050,N_9005);
nor U9183 (N_9183,N_9109,N_9041);
nor U9184 (N_9184,N_9094,N_9092);
or U9185 (N_9185,N_9021,N_8979);
nand U9186 (N_9186,N_9058,N_8990);
or U9187 (N_9187,N_8972,N_9089);
nand U9188 (N_9188,N_9025,N_9042);
nand U9189 (N_9189,N_9064,N_9048);
nor U9190 (N_9190,N_9056,N_9067);
nor U9191 (N_9191,N_8992,N_9027);
or U9192 (N_9192,N_8964,N_9108);
nor U9193 (N_9193,N_8973,N_9053);
and U9194 (N_9194,N_9103,N_9014);
nand U9195 (N_9195,N_9069,N_9106);
nor U9196 (N_9196,N_9049,N_9077);
or U9197 (N_9197,N_9019,N_9105);
and U9198 (N_9198,N_9078,N_9033);
nor U9199 (N_9199,N_8961,N_9046);
nor U9200 (N_9200,N_9003,N_9028);
nand U9201 (N_9201,N_9064,N_9079);
or U9202 (N_9202,N_9103,N_9007);
or U9203 (N_9203,N_8975,N_9067);
and U9204 (N_9204,N_9004,N_8993);
or U9205 (N_9205,N_9032,N_8989);
nor U9206 (N_9206,N_8993,N_9068);
xnor U9207 (N_9207,N_9043,N_8988);
xor U9208 (N_9208,N_9107,N_9032);
or U9209 (N_9209,N_9083,N_9018);
xor U9210 (N_9210,N_9114,N_8998);
nor U9211 (N_9211,N_8966,N_8998);
or U9212 (N_9212,N_9097,N_9092);
and U9213 (N_9213,N_8968,N_9056);
nor U9214 (N_9214,N_9015,N_9031);
nand U9215 (N_9215,N_9063,N_8993);
nor U9216 (N_9216,N_9044,N_8994);
and U9217 (N_9217,N_8973,N_8981);
nand U9218 (N_9218,N_9006,N_9074);
or U9219 (N_9219,N_9033,N_9094);
xor U9220 (N_9220,N_8976,N_9054);
xnor U9221 (N_9221,N_9087,N_9067);
or U9222 (N_9222,N_8985,N_9038);
and U9223 (N_9223,N_8968,N_9026);
nor U9224 (N_9224,N_9088,N_9009);
nand U9225 (N_9225,N_9014,N_9082);
xnor U9226 (N_9226,N_8966,N_9039);
nand U9227 (N_9227,N_9077,N_9045);
nor U9228 (N_9228,N_9086,N_8987);
and U9229 (N_9229,N_9004,N_9115);
and U9230 (N_9230,N_9055,N_8963);
nand U9231 (N_9231,N_9076,N_9012);
xor U9232 (N_9232,N_9078,N_9072);
and U9233 (N_9233,N_9093,N_9110);
nor U9234 (N_9234,N_8960,N_9014);
and U9235 (N_9235,N_9057,N_9118);
xor U9236 (N_9236,N_9010,N_9015);
nor U9237 (N_9237,N_9109,N_9073);
nand U9238 (N_9238,N_9015,N_9033);
nand U9239 (N_9239,N_9002,N_8978);
or U9240 (N_9240,N_9084,N_8976);
xor U9241 (N_9241,N_9077,N_9052);
nor U9242 (N_9242,N_9036,N_9068);
xnor U9243 (N_9243,N_8990,N_9006);
nand U9244 (N_9244,N_9043,N_9059);
and U9245 (N_9245,N_9079,N_9097);
or U9246 (N_9246,N_8972,N_8970);
xor U9247 (N_9247,N_9104,N_9058);
or U9248 (N_9248,N_9106,N_8975);
nor U9249 (N_9249,N_9016,N_9021);
or U9250 (N_9250,N_8983,N_9015);
or U9251 (N_9251,N_9088,N_9046);
or U9252 (N_9252,N_8997,N_9009);
and U9253 (N_9253,N_9119,N_8970);
xnor U9254 (N_9254,N_9021,N_9029);
nand U9255 (N_9255,N_8962,N_9073);
nand U9256 (N_9256,N_9076,N_8988);
nand U9257 (N_9257,N_9027,N_9028);
nand U9258 (N_9258,N_9071,N_9115);
xor U9259 (N_9259,N_9044,N_9071);
and U9260 (N_9260,N_9054,N_8982);
nor U9261 (N_9261,N_9048,N_9072);
and U9262 (N_9262,N_9021,N_9104);
nand U9263 (N_9263,N_9073,N_8993);
nor U9264 (N_9264,N_9032,N_9035);
xor U9265 (N_9265,N_9071,N_9054);
nand U9266 (N_9266,N_9060,N_9091);
nand U9267 (N_9267,N_9032,N_9112);
nor U9268 (N_9268,N_9092,N_8979);
or U9269 (N_9269,N_8960,N_8970);
nor U9270 (N_9270,N_9115,N_8999);
xor U9271 (N_9271,N_9011,N_9059);
nand U9272 (N_9272,N_9117,N_9058);
nand U9273 (N_9273,N_8974,N_9097);
nor U9274 (N_9274,N_8994,N_9001);
nor U9275 (N_9275,N_9042,N_8983);
or U9276 (N_9276,N_9049,N_9101);
and U9277 (N_9277,N_9119,N_9034);
nor U9278 (N_9278,N_8984,N_9116);
xor U9279 (N_9279,N_9012,N_8988);
nor U9280 (N_9280,N_9169,N_9203);
nand U9281 (N_9281,N_9201,N_9173);
nor U9282 (N_9282,N_9241,N_9148);
or U9283 (N_9283,N_9145,N_9134);
or U9284 (N_9284,N_9277,N_9265);
nand U9285 (N_9285,N_9136,N_9197);
nor U9286 (N_9286,N_9256,N_9232);
nand U9287 (N_9287,N_9246,N_9174);
nand U9288 (N_9288,N_9222,N_9243);
nand U9289 (N_9289,N_9261,N_9231);
and U9290 (N_9290,N_9138,N_9124);
or U9291 (N_9291,N_9252,N_9210);
xnor U9292 (N_9292,N_9190,N_9238);
nor U9293 (N_9293,N_9123,N_9274);
nand U9294 (N_9294,N_9216,N_9155);
nand U9295 (N_9295,N_9215,N_9166);
nand U9296 (N_9296,N_9275,N_9120);
xor U9297 (N_9297,N_9221,N_9223);
and U9298 (N_9298,N_9147,N_9213);
or U9299 (N_9299,N_9242,N_9260);
xor U9300 (N_9300,N_9244,N_9264);
nand U9301 (N_9301,N_9142,N_9171);
and U9302 (N_9302,N_9158,N_9144);
and U9303 (N_9303,N_9202,N_9168);
nand U9304 (N_9304,N_9245,N_9188);
and U9305 (N_9305,N_9133,N_9248);
nand U9306 (N_9306,N_9154,N_9157);
nor U9307 (N_9307,N_9257,N_9235);
or U9308 (N_9308,N_9278,N_9159);
nor U9309 (N_9309,N_9146,N_9200);
or U9310 (N_9310,N_9205,N_9214);
or U9311 (N_9311,N_9217,N_9187);
nand U9312 (N_9312,N_9163,N_9209);
nand U9313 (N_9313,N_9143,N_9226);
or U9314 (N_9314,N_9270,N_9276);
nand U9315 (N_9315,N_9279,N_9179);
or U9316 (N_9316,N_9227,N_9126);
and U9317 (N_9317,N_9206,N_9189);
nand U9318 (N_9318,N_9152,N_9185);
or U9319 (N_9319,N_9140,N_9170);
xnor U9320 (N_9320,N_9247,N_9269);
nand U9321 (N_9321,N_9131,N_9262);
nand U9322 (N_9322,N_9258,N_9195);
and U9323 (N_9323,N_9250,N_9128);
and U9324 (N_9324,N_9139,N_9164);
xor U9325 (N_9325,N_9150,N_9125);
nand U9326 (N_9326,N_9183,N_9135);
and U9327 (N_9327,N_9160,N_9153);
or U9328 (N_9328,N_9225,N_9259);
nand U9329 (N_9329,N_9228,N_9178);
nor U9330 (N_9330,N_9127,N_9165);
xnor U9331 (N_9331,N_9186,N_9237);
nand U9332 (N_9332,N_9130,N_9268);
and U9333 (N_9333,N_9156,N_9151);
nand U9334 (N_9334,N_9194,N_9172);
nor U9335 (N_9335,N_9184,N_9239);
xnor U9336 (N_9336,N_9193,N_9122);
xor U9337 (N_9337,N_9149,N_9249);
nor U9338 (N_9338,N_9167,N_9129);
nor U9339 (N_9339,N_9191,N_9255);
and U9340 (N_9340,N_9230,N_9132);
and U9341 (N_9341,N_9219,N_9208);
xor U9342 (N_9342,N_9177,N_9229);
xnor U9343 (N_9343,N_9199,N_9182);
and U9344 (N_9344,N_9234,N_9176);
and U9345 (N_9345,N_9180,N_9192);
or U9346 (N_9346,N_9204,N_9273);
nor U9347 (N_9347,N_9121,N_9271);
nor U9348 (N_9348,N_9212,N_9251);
and U9349 (N_9349,N_9267,N_9141);
xnor U9350 (N_9350,N_9220,N_9218);
and U9351 (N_9351,N_9272,N_9137);
xnor U9352 (N_9352,N_9161,N_9240);
and U9353 (N_9353,N_9181,N_9266);
nor U9354 (N_9354,N_9253,N_9162);
and U9355 (N_9355,N_9254,N_9196);
nor U9356 (N_9356,N_9233,N_9211);
xor U9357 (N_9357,N_9175,N_9207);
nand U9358 (N_9358,N_9198,N_9224);
and U9359 (N_9359,N_9263,N_9236);
nand U9360 (N_9360,N_9220,N_9269);
nand U9361 (N_9361,N_9172,N_9278);
and U9362 (N_9362,N_9245,N_9271);
and U9363 (N_9363,N_9242,N_9144);
nor U9364 (N_9364,N_9123,N_9132);
and U9365 (N_9365,N_9193,N_9163);
nor U9366 (N_9366,N_9229,N_9129);
xor U9367 (N_9367,N_9139,N_9190);
nand U9368 (N_9368,N_9126,N_9252);
xor U9369 (N_9369,N_9227,N_9130);
nor U9370 (N_9370,N_9275,N_9237);
nand U9371 (N_9371,N_9206,N_9168);
nand U9372 (N_9372,N_9188,N_9227);
and U9373 (N_9373,N_9133,N_9240);
and U9374 (N_9374,N_9257,N_9241);
and U9375 (N_9375,N_9171,N_9136);
and U9376 (N_9376,N_9231,N_9173);
or U9377 (N_9377,N_9154,N_9188);
nand U9378 (N_9378,N_9174,N_9135);
and U9379 (N_9379,N_9243,N_9163);
nand U9380 (N_9380,N_9261,N_9201);
or U9381 (N_9381,N_9218,N_9171);
or U9382 (N_9382,N_9152,N_9195);
and U9383 (N_9383,N_9160,N_9120);
and U9384 (N_9384,N_9127,N_9201);
nand U9385 (N_9385,N_9122,N_9169);
xnor U9386 (N_9386,N_9196,N_9195);
nand U9387 (N_9387,N_9207,N_9176);
nor U9388 (N_9388,N_9148,N_9261);
or U9389 (N_9389,N_9220,N_9144);
xnor U9390 (N_9390,N_9269,N_9170);
and U9391 (N_9391,N_9143,N_9167);
nand U9392 (N_9392,N_9127,N_9241);
xor U9393 (N_9393,N_9277,N_9133);
or U9394 (N_9394,N_9260,N_9138);
xnor U9395 (N_9395,N_9129,N_9221);
or U9396 (N_9396,N_9238,N_9205);
xnor U9397 (N_9397,N_9124,N_9226);
or U9398 (N_9398,N_9275,N_9149);
or U9399 (N_9399,N_9244,N_9267);
xnor U9400 (N_9400,N_9132,N_9276);
xnor U9401 (N_9401,N_9121,N_9230);
nor U9402 (N_9402,N_9155,N_9137);
and U9403 (N_9403,N_9262,N_9251);
and U9404 (N_9404,N_9222,N_9237);
xnor U9405 (N_9405,N_9133,N_9214);
nand U9406 (N_9406,N_9167,N_9232);
and U9407 (N_9407,N_9200,N_9257);
nand U9408 (N_9408,N_9248,N_9136);
and U9409 (N_9409,N_9256,N_9137);
nand U9410 (N_9410,N_9146,N_9209);
nor U9411 (N_9411,N_9124,N_9206);
nor U9412 (N_9412,N_9164,N_9185);
xnor U9413 (N_9413,N_9224,N_9251);
nor U9414 (N_9414,N_9253,N_9212);
nor U9415 (N_9415,N_9161,N_9262);
and U9416 (N_9416,N_9167,N_9216);
xor U9417 (N_9417,N_9121,N_9197);
xor U9418 (N_9418,N_9230,N_9204);
xnor U9419 (N_9419,N_9210,N_9128);
or U9420 (N_9420,N_9145,N_9268);
nand U9421 (N_9421,N_9202,N_9162);
xnor U9422 (N_9422,N_9143,N_9271);
or U9423 (N_9423,N_9249,N_9236);
and U9424 (N_9424,N_9197,N_9217);
or U9425 (N_9425,N_9155,N_9122);
xor U9426 (N_9426,N_9242,N_9248);
nand U9427 (N_9427,N_9279,N_9156);
nor U9428 (N_9428,N_9139,N_9261);
nand U9429 (N_9429,N_9203,N_9232);
nand U9430 (N_9430,N_9185,N_9144);
or U9431 (N_9431,N_9196,N_9275);
nor U9432 (N_9432,N_9275,N_9184);
and U9433 (N_9433,N_9174,N_9218);
and U9434 (N_9434,N_9169,N_9181);
nand U9435 (N_9435,N_9274,N_9235);
nor U9436 (N_9436,N_9224,N_9247);
nand U9437 (N_9437,N_9213,N_9227);
nand U9438 (N_9438,N_9264,N_9168);
or U9439 (N_9439,N_9130,N_9201);
nor U9440 (N_9440,N_9434,N_9362);
xor U9441 (N_9441,N_9401,N_9391);
nand U9442 (N_9442,N_9392,N_9310);
or U9443 (N_9443,N_9289,N_9319);
and U9444 (N_9444,N_9347,N_9354);
and U9445 (N_9445,N_9378,N_9291);
and U9446 (N_9446,N_9301,N_9369);
xor U9447 (N_9447,N_9387,N_9437);
or U9448 (N_9448,N_9315,N_9406);
or U9449 (N_9449,N_9399,N_9341);
and U9450 (N_9450,N_9323,N_9417);
nand U9451 (N_9451,N_9305,N_9396);
and U9452 (N_9452,N_9394,N_9339);
xnor U9453 (N_9453,N_9357,N_9326);
nand U9454 (N_9454,N_9321,N_9421);
and U9455 (N_9455,N_9390,N_9324);
xnor U9456 (N_9456,N_9404,N_9283);
nand U9457 (N_9457,N_9311,N_9285);
nor U9458 (N_9458,N_9333,N_9355);
or U9459 (N_9459,N_9429,N_9422);
or U9460 (N_9460,N_9334,N_9353);
xnor U9461 (N_9461,N_9436,N_9338);
or U9462 (N_9462,N_9385,N_9423);
or U9463 (N_9463,N_9379,N_9297);
xnor U9464 (N_9464,N_9382,N_9366);
nor U9465 (N_9465,N_9418,N_9359);
or U9466 (N_9466,N_9349,N_9438);
or U9467 (N_9467,N_9304,N_9383);
or U9468 (N_9468,N_9303,N_9416);
and U9469 (N_9469,N_9344,N_9284);
nand U9470 (N_9470,N_9424,N_9282);
xor U9471 (N_9471,N_9415,N_9371);
nor U9472 (N_9472,N_9308,N_9296);
xnor U9473 (N_9473,N_9368,N_9435);
or U9474 (N_9474,N_9425,N_9336);
nor U9475 (N_9475,N_9287,N_9398);
nor U9476 (N_9476,N_9292,N_9340);
xor U9477 (N_9477,N_9306,N_9420);
nand U9478 (N_9478,N_9411,N_9395);
nor U9479 (N_9479,N_9384,N_9428);
and U9480 (N_9480,N_9403,N_9295);
nand U9481 (N_9481,N_9350,N_9363);
or U9482 (N_9482,N_9412,N_9316);
nand U9483 (N_9483,N_9439,N_9309);
xor U9484 (N_9484,N_9367,N_9322);
nor U9485 (N_9485,N_9294,N_9393);
xor U9486 (N_9486,N_9408,N_9325);
xnor U9487 (N_9487,N_9397,N_9370);
and U9488 (N_9488,N_9328,N_9318);
and U9489 (N_9489,N_9409,N_9427);
xor U9490 (N_9490,N_9431,N_9407);
and U9491 (N_9491,N_9312,N_9281);
or U9492 (N_9492,N_9317,N_9430);
and U9493 (N_9493,N_9389,N_9365);
xor U9494 (N_9494,N_9302,N_9419);
xnor U9495 (N_9495,N_9330,N_9402);
nor U9496 (N_9496,N_9331,N_9374);
nor U9497 (N_9497,N_9346,N_9380);
and U9498 (N_9498,N_9360,N_9356);
nor U9499 (N_9499,N_9320,N_9280);
or U9500 (N_9500,N_9290,N_9414);
and U9501 (N_9501,N_9288,N_9329);
or U9502 (N_9502,N_9335,N_9293);
nand U9503 (N_9503,N_9388,N_9313);
nand U9504 (N_9504,N_9364,N_9433);
xnor U9505 (N_9505,N_9337,N_9327);
nor U9506 (N_9506,N_9314,N_9381);
or U9507 (N_9507,N_9352,N_9372);
and U9508 (N_9508,N_9300,N_9400);
nand U9509 (N_9509,N_9298,N_9332);
or U9510 (N_9510,N_9386,N_9375);
or U9511 (N_9511,N_9307,N_9299);
and U9512 (N_9512,N_9343,N_9413);
nand U9513 (N_9513,N_9377,N_9351);
nor U9514 (N_9514,N_9410,N_9348);
nor U9515 (N_9515,N_9405,N_9426);
nor U9516 (N_9516,N_9373,N_9358);
xor U9517 (N_9517,N_9361,N_9342);
or U9518 (N_9518,N_9286,N_9345);
or U9519 (N_9519,N_9376,N_9432);
and U9520 (N_9520,N_9291,N_9287);
xor U9521 (N_9521,N_9307,N_9400);
nand U9522 (N_9522,N_9405,N_9369);
xnor U9523 (N_9523,N_9306,N_9397);
and U9524 (N_9524,N_9399,N_9325);
nor U9525 (N_9525,N_9395,N_9315);
nand U9526 (N_9526,N_9431,N_9307);
nor U9527 (N_9527,N_9386,N_9397);
xor U9528 (N_9528,N_9325,N_9282);
nor U9529 (N_9529,N_9398,N_9314);
and U9530 (N_9530,N_9375,N_9295);
or U9531 (N_9531,N_9423,N_9361);
or U9532 (N_9532,N_9412,N_9286);
nor U9533 (N_9533,N_9423,N_9294);
xor U9534 (N_9534,N_9381,N_9438);
or U9535 (N_9535,N_9409,N_9396);
nor U9536 (N_9536,N_9391,N_9416);
or U9537 (N_9537,N_9364,N_9347);
or U9538 (N_9538,N_9369,N_9409);
nor U9539 (N_9539,N_9432,N_9416);
xor U9540 (N_9540,N_9338,N_9285);
or U9541 (N_9541,N_9410,N_9300);
nor U9542 (N_9542,N_9367,N_9395);
or U9543 (N_9543,N_9384,N_9344);
xor U9544 (N_9544,N_9384,N_9348);
or U9545 (N_9545,N_9283,N_9436);
nand U9546 (N_9546,N_9420,N_9287);
and U9547 (N_9547,N_9403,N_9332);
nand U9548 (N_9548,N_9323,N_9375);
and U9549 (N_9549,N_9426,N_9418);
or U9550 (N_9550,N_9338,N_9411);
or U9551 (N_9551,N_9437,N_9297);
xnor U9552 (N_9552,N_9301,N_9305);
and U9553 (N_9553,N_9340,N_9428);
and U9554 (N_9554,N_9292,N_9414);
xnor U9555 (N_9555,N_9391,N_9332);
nor U9556 (N_9556,N_9427,N_9420);
nand U9557 (N_9557,N_9356,N_9402);
xnor U9558 (N_9558,N_9431,N_9290);
nor U9559 (N_9559,N_9423,N_9326);
or U9560 (N_9560,N_9415,N_9292);
and U9561 (N_9561,N_9434,N_9371);
xnor U9562 (N_9562,N_9340,N_9417);
xnor U9563 (N_9563,N_9328,N_9329);
or U9564 (N_9564,N_9365,N_9417);
or U9565 (N_9565,N_9364,N_9372);
or U9566 (N_9566,N_9284,N_9338);
and U9567 (N_9567,N_9348,N_9313);
nand U9568 (N_9568,N_9380,N_9285);
xor U9569 (N_9569,N_9417,N_9398);
nand U9570 (N_9570,N_9383,N_9345);
nand U9571 (N_9571,N_9322,N_9332);
nand U9572 (N_9572,N_9348,N_9429);
nand U9573 (N_9573,N_9424,N_9353);
or U9574 (N_9574,N_9430,N_9385);
and U9575 (N_9575,N_9313,N_9347);
xor U9576 (N_9576,N_9288,N_9300);
or U9577 (N_9577,N_9424,N_9366);
and U9578 (N_9578,N_9426,N_9358);
and U9579 (N_9579,N_9370,N_9399);
nand U9580 (N_9580,N_9310,N_9307);
nand U9581 (N_9581,N_9322,N_9385);
nand U9582 (N_9582,N_9291,N_9332);
nand U9583 (N_9583,N_9416,N_9383);
xnor U9584 (N_9584,N_9308,N_9376);
xnor U9585 (N_9585,N_9395,N_9420);
or U9586 (N_9586,N_9439,N_9305);
nand U9587 (N_9587,N_9351,N_9313);
nand U9588 (N_9588,N_9402,N_9309);
and U9589 (N_9589,N_9312,N_9378);
or U9590 (N_9590,N_9359,N_9417);
and U9591 (N_9591,N_9334,N_9340);
or U9592 (N_9592,N_9415,N_9428);
xnor U9593 (N_9593,N_9303,N_9338);
or U9594 (N_9594,N_9281,N_9392);
or U9595 (N_9595,N_9420,N_9314);
xor U9596 (N_9596,N_9288,N_9352);
xnor U9597 (N_9597,N_9375,N_9338);
nor U9598 (N_9598,N_9386,N_9421);
and U9599 (N_9599,N_9314,N_9371);
xor U9600 (N_9600,N_9478,N_9587);
or U9601 (N_9601,N_9499,N_9518);
xnor U9602 (N_9602,N_9522,N_9511);
nand U9603 (N_9603,N_9543,N_9541);
nand U9604 (N_9604,N_9467,N_9472);
and U9605 (N_9605,N_9586,N_9537);
nor U9606 (N_9606,N_9597,N_9545);
xor U9607 (N_9607,N_9491,N_9483);
or U9608 (N_9608,N_9521,N_9480);
nand U9609 (N_9609,N_9556,N_9449);
xnor U9610 (N_9610,N_9457,N_9444);
nor U9611 (N_9611,N_9564,N_9539);
or U9612 (N_9612,N_9454,N_9547);
nor U9613 (N_9613,N_9570,N_9589);
nor U9614 (N_9614,N_9523,N_9445);
or U9615 (N_9615,N_9495,N_9554);
or U9616 (N_9616,N_9484,N_9482);
xor U9617 (N_9617,N_9441,N_9575);
or U9618 (N_9618,N_9448,N_9479);
nand U9619 (N_9619,N_9560,N_9507);
xor U9620 (N_9620,N_9548,N_9513);
or U9621 (N_9621,N_9462,N_9474);
nand U9622 (N_9622,N_9534,N_9536);
nor U9623 (N_9623,N_9497,N_9512);
and U9624 (N_9624,N_9580,N_9519);
nand U9625 (N_9625,N_9527,N_9475);
and U9626 (N_9626,N_9487,N_9452);
or U9627 (N_9627,N_9577,N_9465);
nand U9628 (N_9628,N_9451,N_9500);
nand U9629 (N_9629,N_9529,N_9476);
nor U9630 (N_9630,N_9558,N_9594);
and U9631 (N_9631,N_9591,N_9542);
or U9632 (N_9632,N_9466,N_9549);
nand U9633 (N_9633,N_9525,N_9596);
and U9634 (N_9634,N_9471,N_9574);
or U9635 (N_9635,N_9490,N_9486);
or U9636 (N_9636,N_9488,N_9563);
xnor U9637 (N_9637,N_9485,N_9477);
xor U9638 (N_9638,N_9583,N_9515);
xnor U9639 (N_9639,N_9551,N_9559);
and U9640 (N_9640,N_9509,N_9581);
and U9641 (N_9641,N_9463,N_9464);
nor U9642 (N_9642,N_9544,N_9503);
nor U9643 (N_9643,N_9443,N_9598);
or U9644 (N_9644,N_9442,N_9546);
nand U9645 (N_9645,N_9489,N_9568);
or U9646 (N_9646,N_9456,N_9440);
nor U9647 (N_9647,N_9453,N_9550);
nor U9648 (N_9648,N_9526,N_9567);
nand U9649 (N_9649,N_9460,N_9592);
or U9650 (N_9650,N_9504,N_9555);
xnor U9651 (N_9651,N_9455,N_9458);
nand U9652 (N_9652,N_9585,N_9528);
xnor U9653 (N_9653,N_9561,N_9565);
nand U9654 (N_9654,N_9538,N_9505);
nor U9655 (N_9655,N_9566,N_9535);
and U9656 (N_9656,N_9502,N_9595);
nor U9657 (N_9657,N_9493,N_9510);
or U9658 (N_9658,N_9520,N_9557);
xnor U9659 (N_9659,N_9469,N_9590);
or U9660 (N_9660,N_9572,N_9593);
xnor U9661 (N_9661,N_9571,N_9552);
or U9662 (N_9662,N_9540,N_9468);
xnor U9663 (N_9663,N_9492,N_9533);
and U9664 (N_9664,N_9517,N_9578);
nor U9665 (N_9665,N_9599,N_9473);
xnor U9666 (N_9666,N_9524,N_9569);
nor U9667 (N_9667,N_9588,N_9579);
or U9668 (N_9668,N_9531,N_9506);
nand U9669 (N_9669,N_9450,N_9530);
and U9670 (N_9670,N_9501,N_9553);
or U9671 (N_9671,N_9494,N_9481);
nand U9672 (N_9672,N_9582,N_9447);
nand U9673 (N_9673,N_9573,N_9446);
and U9674 (N_9674,N_9461,N_9508);
nand U9675 (N_9675,N_9584,N_9498);
or U9676 (N_9676,N_9532,N_9470);
and U9677 (N_9677,N_9576,N_9562);
xnor U9678 (N_9678,N_9496,N_9459);
and U9679 (N_9679,N_9516,N_9514);
nor U9680 (N_9680,N_9446,N_9494);
nand U9681 (N_9681,N_9485,N_9444);
or U9682 (N_9682,N_9556,N_9521);
or U9683 (N_9683,N_9513,N_9529);
nor U9684 (N_9684,N_9491,N_9565);
and U9685 (N_9685,N_9597,N_9456);
or U9686 (N_9686,N_9473,N_9484);
xnor U9687 (N_9687,N_9494,N_9551);
xnor U9688 (N_9688,N_9442,N_9571);
xnor U9689 (N_9689,N_9469,N_9472);
nor U9690 (N_9690,N_9595,N_9461);
and U9691 (N_9691,N_9545,N_9497);
and U9692 (N_9692,N_9506,N_9511);
and U9693 (N_9693,N_9549,N_9478);
or U9694 (N_9694,N_9527,N_9461);
or U9695 (N_9695,N_9531,N_9576);
nand U9696 (N_9696,N_9579,N_9552);
xnor U9697 (N_9697,N_9474,N_9510);
or U9698 (N_9698,N_9488,N_9526);
and U9699 (N_9699,N_9448,N_9461);
nand U9700 (N_9700,N_9532,N_9566);
and U9701 (N_9701,N_9460,N_9477);
and U9702 (N_9702,N_9500,N_9519);
nand U9703 (N_9703,N_9498,N_9458);
nor U9704 (N_9704,N_9547,N_9545);
nand U9705 (N_9705,N_9584,N_9492);
xnor U9706 (N_9706,N_9492,N_9543);
xnor U9707 (N_9707,N_9595,N_9489);
xnor U9708 (N_9708,N_9489,N_9460);
nand U9709 (N_9709,N_9528,N_9540);
xnor U9710 (N_9710,N_9531,N_9499);
nand U9711 (N_9711,N_9520,N_9494);
or U9712 (N_9712,N_9524,N_9444);
xor U9713 (N_9713,N_9566,N_9574);
xnor U9714 (N_9714,N_9512,N_9501);
nand U9715 (N_9715,N_9470,N_9550);
nor U9716 (N_9716,N_9538,N_9453);
or U9717 (N_9717,N_9518,N_9478);
nor U9718 (N_9718,N_9474,N_9482);
or U9719 (N_9719,N_9564,N_9514);
xnor U9720 (N_9720,N_9598,N_9573);
nor U9721 (N_9721,N_9571,N_9477);
nor U9722 (N_9722,N_9462,N_9546);
nand U9723 (N_9723,N_9588,N_9547);
xor U9724 (N_9724,N_9543,N_9442);
nand U9725 (N_9725,N_9558,N_9478);
nand U9726 (N_9726,N_9502,N_9480);
or U9727 (N_9727,N_9501,N_9507);
or U9728 (N_9728,N_9544,N_9445);
and U9729 (N_9729,N_9549,N_9580);
nor U9730 (N_9730,N_9515,N_9448);
nor U9731 (N_9731,N_9566,N_9587);
nor U9732 (N_9732,N_9476,N_9592);
nand U9733 (N_9733,N_9567,N_9481);
or U9734 (N_9734,N_9449,N_9562);
or U9735 (N_9735,N_9591,N_9463);
nor U9736 (N_9736,N_9574,N_9583);
nor U9737 (N_9737,N_9475,N_9543);
or U9738 (N_9738,N_9458,N_9556);
nor U9739 (N_9739,N_9478,N_9574);
nor U9740 (N_9740,N_9581,N_9534);
and U9741 (N_9741,N_9570,N_9527);
xor U9742 (N_9742,N_9513,N_9497);
nand U9743 (N_9743,N_9535,N_9450);
xnor U9744 (N_9744,N_9507,N_9506);
xnor U9745 (N_9745,N_9523,N_9592);
and U9746 (N_9746,N_9579,N_9509);
xor U9747 (N_9747,N_9556,N_9476);
and U9748 (N_9748,N_9445,N_9502);
or U9749 (N_9749,N_9516,N_9505);
xor U9750 (N_9750,N_9450,N_9469);
nand U9751 (N_9751,N_9572,N_9597);
nor U9752 (N_9752,N_9506,N_9560);
nand U9753 (N_9753,N_9544,N_9502);
or U9754 (N_9754,N_9566,N_9534);
nand U9755 (N_9755,N_9591,N_9576);
and U9756 (N_9756,N_9571,N_9501);
or U9757 (N_9757,N_9567,N_9540);
nand U9758 (N_9758,N_9503,N_9553);
nor U9759 (N_9759,N_9472,N_9495);
nand U9760 (N_9760,N_9643,N_9690);
nor U9761 (N_9761,N_9618,N_9686);
or U9762 (N_9762,N_9645,N_9691);
nand U9763 (N_9763,N_9665,N_9751);
nand U9764 (N_9764,N_9684,N_9699);
and U9765 (N_9765,N_9600,N_9688);
and U9766 (N_9766,N_9725,N_9673);
nor U9767 (N_9767,N_9619,N_9629);
and U9768 (N_9768,N_9612,N_9709);
nand U9769 (N_9769,N_9670,N_9701);
nor U9770 (N_9770,N_9644,N_9624);
or U9771 (N_9771,N_9743,N_9649);
and U9772 (N_9772,N_9747,N_9613);
or U9773 (N_9773,N_9621,N_9755);
nand U9774 (N_9774,N_9666,N_9711);
nor U9775 (N_9775,N_9716,N_9680);
xor U9776 (N_9776,N_9687,N_9605);
nand U9777 (N_9777,N_9733,N_9677);
nor U9778 (N_9778,N_9722,N_9606);
nor U9779 (N_9779,N_9622,N_9635);
or U9780 (N_9780,N_9745,N_9658);
xor U9781 (N_9781,N_9672,N_9671);
xnor U9782 (N_9782,N_9603,N_9655);
and U9783 (N_9783,N_9689,N_9728);
nand U9784 (N_9784,N_9748,N_9726);
xor U9785 (N_9785,N_9668,N_9694);
nand U9786 (N_9786,N_9741,N_9607);
nand U9787 (N_9787,N_9744,N_9610);
nand U9788 (N_9788,N_9702,N_9625);
and U9789 (N_9789,N_9692,N_9674);
or U9790 (N_9790,N_9660,N_9609);
and U9791 (N_9791,N_9700,N_9639);
nor U9792 (N_9792,N_9620,N_9735);
or U9793 (N_9793,N_9710,N_9642);
xor U9794 (N_9794,N_9602,N_9732);
nor U9795 (N_9795,N_9632,N_9614);
or U9796 (N_9796,N_9731,N_9634);
or U9797 (N_9797,N_9752,N_9681);
nand U9798 (N_9798,N_9651,N_9608);
nand U9799 (N_9799,N_9647,N_9640);
nor U9800 (N_9800,N_9682,N_9707);
nor U9801 (N_9801,N_9737,N_9718);
and U9802 (N_9802,N_9636,N_9667);
xor U9803 (N_9803,N_9641,N_9756);
or U9804 (N_9804,N_9715,N_9724);
nor U9805 (N_9805,N_9631,N_9742);
nor U9806 (N_9806,N_9697,N_9730);
and U9807 (N_9807,N_9753,N_9719);
or U9808 (N_9808,N_9738,N_9696);
or U9809 (N_9809,N_9714,N_9661);
xnor U9810 (N_9810,N_9633,N_9617);
or U9811 (N_9811,N_9626,N_9695);
nand U9812 (N_9812,N_9727,N_9615);
or U9813 (N_9813,N_9683,N_9721);
nor U9814 (N_9814,N_9601,N_9705);
or U9815 (N_9815,N_9662,N_9720);
and U9816 (N_9816,N_9703,N_9712);
nand U9817 (N_9817,N_9669,N_9746);
nand U9818 (N_9818,N_9754,N_9650);
and U9819 (N_9819,N_9664,N_9708);
nand U9820 (N_9820,N_9729,N_9627);
xor U9821 (N_9821,N_9704,N_9648);
or U9822 (N_9822,N_9758,N_9623);
and U9823 (N_9823,N_9675,N_9637);
or U9824 (N_9824,N_9638,N_9740);
or U9825 (N_9825,N_9736,N_9646);
nand U9826 (N_9826,N_9693,N_9739);
nor U9827 (N_9827,N_9663,N_9676);
nor U9828 (N_9828,N_9757,N_9657);
nor U9829 (N_9829,N_9653,N_9685);
nand U9830 (N_9830,N_9616,N_9750);
xnor U9831 (N_9831,N_9611,N_9628);
xnor U9832 (N_9832,N_9698,N_9659);
and U9833 (N_9833,N_9713,N_9656);
xnor U9834 (N_9834,N_9749,N_9734);
nand U9835 (N_9835,N_9717,N_9679);
or U9836 (N_9836,N_9706,N_9630);
nor U9837 (N_9837,N_9652,N_9604);
nand U9838 (N_9838,N_9678,N_9759);
and U9839 (N_9839,N_9654,N_9723);
and U9840 (N_9840,N_9724,N_9652);
or U9841 (N_9841,N_9714,N_9731);
and U9842 (N_9842,N_9696,N_9703);
xnor U9843 (N_9843,N_9662,N_9690);
and U9844 (N_9844,N_9699,N_9631);
xor U9845 (N_9845,N_9661,N_9718);
nor U9846 (N_9846,N_9684,N_9718);
nor U9847 (N_9847,N_9654,N_9744);
nand U9848 (N_9848,N_9655,N_9732);
nand U9849 (N_9849,N_9623,N_9655);
xnor U9850 (N_9850,N_9647,N_9745);
nor U9851 (N_9851,N_9622,N_9721);
nor U9852 (N_9852,N_9753,N_9600);
xnor U9853 (N_9853,N_9621,N_9602);
and U9854 (N_9854,N_9731,N_9721);
or U9855 (N_9855,N_9630,N_9755);
xnor U9856 (N_9856,N_9752,N_9657);
and U9857 (N_9857,N_9619,N_9615);
and U9858 (N_9858,N_9604,N_9670);
or U9859 (N_9859,N_9643,N_9607);
nor U9860 (N_9860,N_9661,N_9631);
and U9861 (N_9861,N_9616,N_9723);
or U9862 (N_9862,N_9680,N_9671);
nand U9863 (N_9863,N_9683,N_9700);
and U9864 (N_9864,N_9626,N_9759);
nor U9865 (N_9865,N_9650,N_9688);
nand U9866 (N_9866,N_9693,N_9644);
or U9867 (N_9867,N_9717,N_9619);
xnor U9868 (N_9868,N_9718,N_9744);
and U9869 (N_9869,N_9733,N_9630);
nor U9870 (N_9870,N_9740,N_9635);
nand U9871 (N_9871,N_9686,N_9754);
nor U9872 (N_9872,N_9723,N_9744);
or U9873 (N_9873,N_9665,N_9732);
nand U9874 (N_9874,N_9647,N_9657);
nor U9875 (N_9875,N_9638,N_9646);
nand U9876 (N_9876,N_9706,N_9647);
nor U9877 (N_9877,N_9602,N_9695);
nor U9878 (N_9878,N_9742,N_9739);
nand U9879 (N_9879,N_9754,N_9613);
and U9880 (N_9880,N_9720,N_9747);
nand U9881 (N_9881,N_9759,N_9689);
xor U9882 (N_9882,N_9755,N_9636);
xor U9883 (N_9883,N_9672,N_9642);
xnor U9884 (N_9884,N_9657,N_9758);
xnor U9885 (N_9885,N_9733,N_9708);
xnor U9886 (N_9886,N_9718,N_9629);
xor U9887 (N_9887,N_9661,N_9751);
xor U9888 (N_9888,N_9697,N_9627);
nor U9889 (N_9889,N_9646,N_9735);
nand U9890 (N_9890,N_9637,N_9649);
nand U9891 (N_9891,N_9656,N_9701);
nor U9892 (N_9892,N_9620,N_9605);
nor U9893 (N_9893,N_9627,N_9717);
xor U9894 (N_9894,N_9732,N_9680);
xor U9895 (N_9895,N_9748,N_9658);
xnor U9896 (N_9896,N_9630,N_9727);
nor U9897 (N_9897,N_9672,N_9626);
and U9898 (N_9898,N_9742,N_9646);
nand U9899 (N_9899,N_9606,N_9654);
and U9900 (N_9900,N_9677,N_9748);
nand U9901 (N_9901,N_9659,N_9709);
xnor U9902 (N_9902,N_9627,N_9652);
and U9903 (N_9903,N_9619,N_9667);
nand U9904 (N_9904,N_9637,N_9647);
and U9905 (N_9905,N_9650,N_9730);
xor U9906 (N_9906,N_9677,N_9659);
nor U9907 (N_9907,N_9654,N_9687);
or U9908 (N_9908,N_9636,N_9675);
or U9909 (N_9909,N_9700,N_9658);
xor U9910 (N_9910,N_9747,N_9656);
nor U9911 (N_9911,N_9688,N_9711);
nor U9912 (N_9912,N_9665,N_9727);
and U9913 (N_9913,N_9613,N_9678);
nand U9914 (N_9914,N_9703,N_9612);
and U9915 (N_9915,N_9621,N_9618);
or U9916 (N_9916,N_9706,N_9664);
and U9917 (N_9917,N_9744,N_9694);
nand U9918 (N_9918,N_9646,N_9759);
nand U9919 (N_9919,N_9606,N_9632);
xnor U9920 (N_9920,N_9777,N_9898);
nand U9921 (N_9921,N_9805,N_9764);
and U9922 (N_9922,N_9868,N_9842);
nor U9923 (N_9923,N_9783,N_9811);
or U9924 (N_9924,N_9802,N_9846);
and U9925 (N_9925,N_9801,N_9787);
nand U9926 (N_9926,N_9839,N_9844);
or U9927 (N_9927,N_9911,N_9775);
nand U9928 (N_9928,N_9803,N_9856);
and U9929 (N_9929,N_9828,N_9854);
xnor U9930 (N_9930,N_9873,N_9904);
nand U9931 (N_9931,N_9900,N_9849);
or U9932 (N_9932,N_9793,N_9786);
and U9933 (N_9933,N_9776,N_9913);
xnor U9934 (N_9934,N_9762,N_9788);
or U9935 (N_9935,N_9810,N_9870);
nand U9936 (N_9936,N_9785,N_9878);
nand U9937 (N_9937,N_9822,N_9852);
and U9938 (N_9938,N_9778,N_9864);
xnor U9939 (N_9939,N_9855,N_9899);
nor U9940 (N_9940,N_9851,N_9831);
nor U9941 (N_9941,N_9903,N_9910);
nand U9942 (N_9942,N_9885,N_9848);
nand U9943 (N_9943,N_9876,N_9797);
nor U9944 (N_9944,N_9808,N_9871);
xnor U9945 (N_9945,N_9825,N_9843);
and U9946 (N_9946,N_9845,N_9861);
nor U9947 (N_9947,N_9887,N_9818);
or U9948 (N_9948,N_9795,N_9792);
and U9949 (N_9949,N_9813,N_9765);
xnor U9950 (N_9950,N_9829,N_9826);
and U9951 (N_9951,N_9817,N_9841);
nor U9952 (N_9952,N_9883,N_9880);
and U9953 (N_9953,N_9796,N_9781);
and U9954 (N_9954,N_9890,N_9891);
nand U9955 (N_9955,N_9824,N_9807);
and U9956 (N_9956,N_9820,N_9798);
or U9957 (N_9957,N_9780,N_9760);
nor U9958 (N_9958,N_9832,N_9872);
nor U9959 (N_9959,N_9884,N_9768);
xor U9960 (N_9960,N_9853,N_9874);
or U9961 (N_9961,N_9916,N_9888);
nor U9962 (N_9962,N_9794,N_9830);
xor U9963 (N_9963,N_9827,N_9906);
nor U9964 (N_9964,N_9815,N_9858);
or U9965 (N_9965,N_9879,N_9902);
and U9966 (N_9966,N_9837,N_9833);
nor U9967 (N_9967,N_9909,N_9761);
and U9968 (N_9968,N_9894,N_9770);
nor U9969 (N_9969,N_9919,N_9881);
nand U9970 (N_9970,N_9836,N_9812);
nor U9971 (N_9971,N_9893,N_9819);
nor U9972 (N_9972,N_9774,N_9869);
xnor U9973 (N_9973,N_9866,N_9800);
nand U9974 (N_9974,N_9867,N_9821);
nand U9975 (N_9975,N_9901,N_9882);
and U9976 (N_9976,N_9863,N_9789);
and U9977 (N_9977,N_9877,N_9840);
and U9978 (N_9978,N_9806,N_9865);
xor U9979 (N_9979,N_9769,N_9895);
xor U9980 (N_9980,N_9857,N_9809);
or U9981 (N_9981,N_9799,N_9816);
or U9982 (N_9982,N_9850,N_9766);
nand U9983 (N_9983,N_9790,N_9860);
nor U9984 (N_9984,N_9918,N_9771);
or U9985 (N_9985,N_9897,N_9908);
xnor U9986 (N_9986,N_9917,N_9896);
xor U9987 (N_9987,N_9834,N_9859);
xor U9988 (N_9988,N_9782,N_9823);
xor U9989 (N_9989,N_9779,N_9905);
nor U9990 (N_9990,N_9889,N_9862);
xor U9991 (N_9991,N_9838,N_9784);
nand U9992 (N_9992,N_9914,N_9847);
nor U9993 (N_9993,N_9763,N_9767);
or U9994 (N_9994,N_9886,N_9773);
xor U9995 (N_9995,N_9804,N_9791);
or U9996 (N_9996,N_9907,N_9875);
nor U9997 (N_9997,N_9912,N_9892);
nand U9998 (N_9998,N_9772,N_9915);
and U9999 (N_9999,N_9835,N_9814);
nand U10000 (N_10000,N_9786,N_9910);
nor U10001 (N_10001,N_9784,N_9791);
and U10002 (N_10002,N_9766,N_9917);
nand U10003 (N_10003,N_9783,N_9902);
and U10004 (N_10004,N_9830,N_9914);
nand U10005 (N_10005,N_9875,N_9873);
xnor U10006 (N_10006,N_9911,N_9895);
nand U10007 (N_10007,N_9848,N_9772);
or U10008 (N_10008,N_9777,N_9818);
nand U10009 (N_10009,N_9885,N_9793);
xor U10010 (N_10010,N_9859,N_9780);
nor U10011 (N_10011,N_9835,N_9859);
and U10012 (N_10012,N_9891,N_9809);
or U10013 (N_10013,N_9897,N_9835);
or U10014 (N_10014,N_9877,N_9830);
and U10015 (N_10015,N_9794,N_9902);
and U10016 (N_10016,N_9852,N_9775);
nand U10017 (N_10017,N_9847,N_9768);
nor U10018 (N_10018,N_9762,N_9836);
and U10019 (N_10019,N_9802,N_9821);
nor U10020 (N_10020,N_9841,N_9806);
xnor U10021 (N_10021,N_9787,N_9913);
nor U10022 (N_10022,N_9833,N_9838);
or U10023 (N_10023,N_9811,N_9816);
xnor U10024 (N_10024,N_9845,N_9888);
nand U10025 (N_10025,N_9904,N_9760);
and U10026 (N_10026,N_9896,N_9831);
xor U10027 (N_10027,N_9896,N_9812);
and U10028 (N_10028,N_9780,N_9781);
nand U10029 (N_10029,N_9888,N_9812);
xor U10030 (N_10030,N_9800,N_9844);
and U10031 (N_10031,N_9870,N_9866);
and U10032 (N_10032,N_9786,N_9912);
nand U10033 (N_10033,N_9885,N_9904);
nand U10034 (N_10034,N_9893,N_9919);
and U10035 (N_10035,N_9870,N_9862);
and U10036 (N_10036,N_9877,N_9906);
nand U10037 (N_10037,N_9840,N_9807);
and U10038 (N_10038,N_9793,N_9914);
or U10039 (N_10039,N_9814,N_9842);
nor U10040 (N_10040,N_9762,N_9829);
or U10041 (N_10041,N_9882,N_9853);
xor U10042 (N_10042,N_9866,N_9838);
xor U10043 (N_10043,N_9806,N_9859);
and U10044 (N_10044,N_9802,N_9860);
nor U10045 (N_10045,N_9826,N_9798);
xnor U10046 (N_10046,N_9783,N_9787);
or U10047 (N_10047,N_9896,N_9793);
nor U10048 (N_10048,N_9797,N_9892);
nand U10049 (N_10049,N_9863,N_9779);
xnor U10050 (N_10050,N_9782,N_9913);
nand U10051 (N_10051,N_9768,N_9860);
nand U10052 (N_10052,N_9790,N_9767);
and U10053 (N_10053,N_9813,N_9839);
and U10054 (N_10054,N_9812,N_9879);
and U10055 (N_10055,N_9866,N_9805);
nor U10056 (N_10056,N_9902,N_9770);
or U10057 (N_10057,N_9884,N_9776);
nand U10058 (N_10058,N_9840,N_9811);
or U10059 (N_10059,N_9907,N_9862);
and U10060 (N_10060,N_9836,N_9766);
nor U10061 (N_10061,N_9765,N_9889);
and U10062 (N_10062,N_9914,N_9876);
and U10063 (N_10063,N_9869,N_9777);
and U10064 (N_10064,N_9813,N_9847);
nand U10065 (N_10065,N_9804,N_9827);
or U10066 (N_10066,N_9770,N_9781);
nand U10067 (N_10067,N_9783,N_9913);
or U10068 (N_10068,N_9776,N_9879);
or U10069 (N_10069,N_9793,N_9831);
or U10070 (N_10070,N_9853,N_9810);
xor U10071 (N_10071,N_9803,N_9793);
and U10072 (N_10072,N_9786,N_9832);
xnor U10073 (N_10073,N_9885,N_9792);
nor U10074 (N_10074,N_9811,N_9853);
nand U10075 (N_10075,N_9914,N_9761);
nor U10076 (N_10076,N_9808,N_9830);
and U10077 (N_10077,N_9831,N_9790);
nor U10078 (N_10078,N_9895,N_9897);
and U10079 (N_10079,N_9849,N_9769);
or U10080 (N_10080,N_9961,N_10045);
or U10081 (N_10081,N_9937,N_10050);
nor U10082 (N_10082,N_10017,N_9934);
xnor U10083 (N_10083,N_9921,N_10016);
nand U10084 (N_10084,N_9976,N_10023);
xor U10085 (N_10085,N_9950,N_10035);
and U10086 (N_10086,N_10036,N_9927);
xor U10087 (N_10087,N_9982,N_10066);
nand U10088 (N_10088,N_9971,N_10057);
nor U10089 (N_10089,N_9979,N_10068);
or U10090 (N_10090,N_10056,N_9930);
nand U10091 (N_10091,N_10047,N_9944);
and U10092 (N_10092,N_9959,N_9966);
nor U10093 (N_10093,N_10054,N_10011);
and U10094 (N_10094,N_10002,N_9975);
nand U10095 (N_10095,N_10060,N_9998);
or U10096 (N_10096,N_10029,N_10031);
xor U10097 (N_10097,N_9932,N_10030);
xor U10098 (N_10098,N_10075,N_9926);
or U10099 (N_10099,N_9948,N_10037);
xnor U10100 (N_10100,N_9977,N_10004);
xor U10101 (N_10101,N_9989,N_9957);
nor U10102 (N_10102,N_10043,N_9956);
and U10103 (N_10103,N_10061,N_10027);
and U10104 (N_10104,N_9962,N_10024);
xor U10105 (N_10105,N_9981,N_9920);
and U10106 (N_10106,N_10012,N_9958);
nand U10107 (N_10107,N_9945,N_10063);
nor U10108 (N_10108,N_9974,N_10064);
or U10109 (N_10109,N_10032,N_10009);
nor U10110 (N_10110,N_9960,N_9999);
and U10111 (N_10111,N_9988,N_9946);
xor U10112 (N_10112,N_9924,N_10069);
nand U10113 (N_10113,N_9941,N_10025);
xor U10114 (N_10114,N_9935,N_10052);
xor U10115 (N_10115,N_9949,N_9968);
and U10116 (N_10116,N_9985,N_10018);
xnor U10117 (N_10117,N_10074,N_10049);
or U10118 (N_10118,N_9969,N_9994);
xor U10119 (N_10119,N_10076,N_9990);
nor U10120 (N_10120,N_10014,N_10040);
nand U10121 (N_10121,N_10048,N_9955);
xnor U10122 (N_10122,N_10044,N_9965);
xnor U10123 (N_10123,N_9923,N_9922);
and U10124 (N_10124,N_10008,N_9940);
nand U10125 (N_10125,N_10058,N_10038);
xor U10126 (N_10126,N_9995,N_9947);
and U10127 (N_10127,N_9943,N_9983);
xnor U10128 (N_10128,N_9964,N_9973);
or U10129 (N_10129,N_10006,N_10046);
nor U10130 (N_10130,N_10053,N_10051);
nor U10131 (N_10131,N_9963,N_9929);
and U10132 (N_10132,N_10071,N_10059);
nor U10133 (N_10133,N_10026,N_10077);
and U10134 (N_10134,N_10020,N_9942);
nand U10135 (N_10135,N_10039,N_9933);
nor U10136 (N_10136,N_10073,N_9967);
nor U10137 (N_10137,N_10005,N_9936);
or U10138 (N_10138,N_9970,N_9972);
nand U10139 (N_10139,N_9953,N_9986);
or U10140 (N_10140,N_10065,N_10072);
or U10141 (N_10141,N_9939,N_10070);
and U10142 (N_10142,N_10010,N_10019);
or U10143 (N_10143,N_10021,N_9993);
or U10144 (N_10144,N_9954,N_9996);
nand U10145 (N_10145,N_9984,N_10028);
nor U10146 (N_10146,N_9987,N_10007);
xor U10147 (N_10147,N_9951,N_10067);
or U10148 (N_10148,N_10078,N_9978);
nand U10149 (N_10149,N_10055,N_9928);
xor U10150 (N_10150,N_10000,N_10003);
nand U10151 (N_10151,N_10041,N_9938);
or U10152 (N_10152,N_10022,N_10001);
nor U10153 (N_10153,N_9992,N_9991);
nand U10154 (N_10154,N_9925,N_10013);
and U10155 (N_10155,N_10034,N_10033);
nor U10156 (N_10156,N_9980,N_9997);
xnor U10157 (N_10157,N_9952,N_9931);
nand U10158 (N_10158,N_10015,N_10079);
xnor U10159 (N_10159,N_10062,N_10042);
nand U10160 (N_10160,N_9966,N_9964);
and U10161 (N_10161,N_10079,N_10030);
xnor U10162 (N_10162,N_9990,N_10060);
xor U10163 (N_10163,N_9971,N_10009);
and U10164 (N_10164,N_9925,N_9928);
and U10165 (N_10165,N_10052,N_9981);
and U10166 (N_10166,N_9998,N_10024);
and U10167 (N_10167,N_10065,N_10029);
nand U10168 (N_10168,N_9976,N_10017);
nor U10169 (N_10169,N_9957,N_9952);
nand U10170 (N_10170,N_9965,N_9955);
nand U10171 (N_10171,N_9995,N_9944);
and U10172 (N_10172,N_10054,N_9957);
nand U10173 (N_10173,N_10070,N_10067);
nor U10174 (N_10174,N_10021,N_9994);
xnor U10175 (N_10175,N_10024,N_9952);
or U10176 (N_10176,N_9996,N_10038);
xnor U10177 (N_10177,N_9945,N_9941);
xnor U10178 (N_10178,N_9999,N_9955);
and U10179 (N_10179,N_9951,N_10017);
or U10180 (N_10180,N_10029,N_10002);
xnor U10181 (N_10181,N_9920,N_10005);
and U10182 (N_10182,N_9990,N_10064);
nand U10183 (N_10183,N_9965,N_9979);
nor U10184 (N_10184,N_10019,N_10012);
xnor U10185 (N_10185,N_9971,N_10023);
xor U10186 (N_10186,N_9973,N_10058);
nor U10187 (N_10187,N_10044,N_9968);
xor U10188 (N_10188,N_9995,N_9922);
and U10189 (N_10189,N_9980,N_10012);
or U10190 (N_10190,N_9946,N_10043);
nor U10191 (N_10191,N_9928,N_10057);
and U10192 (N_10192,N_9949,N_10042);
nand U10193 (N_10193,N_9981,N_10044);
nand U10194 (N_10194,N_9988,N_10069);
or U10195 (N_10195,N_10050,N_9967);
or U10196 (N_10196,N_10071,N_9991);
and U10197 (N_10197,N_10020,N_10011);
xnor U10198 (N_10198,N_10058,N_9931);
nand U10199 (N_10199,N_9959,N_9926);
or U10200 (N_10200,N_9987,N_9922);
nand U10201 (N_10201,N_9962,N_10001);
xnor U10202 (N_10202,N_9991,N_9928);
nor U10203 (N_10203,N_10049,N_10052);
or U10204 (N_10204,N_10034,N_9941);
nor U10205 (N_10205,N_9964,N_10003);
or U10206 (N_10206,N_10048,N_9957);
nand U10207 (N_10207,N_9941,N_9938);
nor U10208 (N_10208,N_9922,N_9991);
xor U10209 (N_10209,N_9923,N_10063);
nor U10210 (N_10210,N_10037,N_10028);
nand U10211 (N_10211,N_9994,N_9991);
nor U10212 (N_10212,N_9968,N_10024);
nor U10213 (N_10213,N_9935,N_9941);
xor U10214 (N_10214,N_9923,N_9920);
or U10215 (N_10215,N_10035,N_10013);
xor U10216 (N_10216,N_10067,N_9968);
nor U10217 (N_10217,N_9941,N_10028);
or U10218 (N_10218,N_9974,N_9969);
or U10219 (N_10219,N_10066,N_10010);
nand U10220 (N_10220,N_9930,N_10028);
or U10221 (N_10221,N_10065,N_9947);
xnor U10222 (N_10222,N_9937,N_9981);
xor U10223 (N_10223,N_9926,N_9995);
or U10224 (N_10224,N_9991,N_9971);
xor U10225 (N_10225,N_9971,N_10024);
nand U10226 (N_10226,N_10049,N_10067);
nor U10227 (N_10227,N_10025,N_9928);
nand U10228 (N_10228,N_10059,N_9943);
xnor U10229 (N_10229,N_9999,N_10017);
nor U10230 (N_10230,N_9920,N_9929);
or U10231 (N_10231,N_9932,N_9987);
or U10232 (N_10232,N_10060,N_9932);
or U10233 (N_10233,N_10056,N_10067);
nand U10234 (N_10234,N_9922,N_10007);
or U10235 (N_10235,N_9997,N_9942);
nor U10236 (N_10236,N_10025,N_9971);
and U10237 (N_10237,N_10004,N_9935);
or U10238 (N_10238,N_9931,N_9975);
xnor U10239 (N_10239,N_9973,N_9986);
or U10240 (N_10240,N_10117,N_10127);
nor U10241 (N_10241,N_10186,N_10210);
nor U10242 (N_10242,N_10223,N_10113);
nand U10243 (N_10243,N_10213,N_10196);
or U10244 (N_10244,N_10193,N_10172);
xor U10245 (N_10245,N_10100,N_10156);
and U10246 (N_10246,N_10226,N_10142);
xor U10247 (N_10247,N_10123,N_10209);
nor U10248 (N_10248,N_10237,N_10141);
xor U10249 (N_10249,N_10134,N_10205);
nand U10250 (N_10250,N_10084,N_10129);
or U10251 (N_10251,N_10218,N_10103);
or U10252 (N_10252,N_10102,N_10201);
and U10253 (N_10253,N_10155,N_10121);
and U10254 (N_10254,N_10085,N_10108);
or U10255 (N_10255,N_10116,N_10114);
nor U10256 (N_10256,N_10194,N_10107);
nor U10257 (N_10257,N_10191,N_10128);
nor U10258 (N_10258,N_10200,N_10080);
or U10259 (N_10259,N_10180,N_10119);
and U10260 (N_10260,N_10125,N_10124);
nand U10261 (N_10261,N_10195,N_10207);
nand U10262 (N_10262,N_10190,N_10146);
nand U10263 (N_10263,N_10118,N_10228);
nand U10264 (N_10264,N_10203,N_10173);
or U10265 (N_10265,N_10115,N_10182);
or U10266 (N_10266,N_10143,N_10154);
and U10267 (N_10267,N_10130,N_10235);
nor U10268 (N_10268,N_10167,N_10192);
and U10269 (N_10269,N_10229,N_10139);
nand U10270 (N_10270,N_10144,N_10163);
nand U10271 (N_10271,N_10166,N_10234);
or U10272 (N_10272,N_10110,N_10099);
nand U10273 (N_10273,N_10239,N_10087);
and U10274 (N_10274,N_10090,N_10152);
or U10275 (N_10275,N_10093,N_10225);
and U10276 (N_10276,N_10135,N_10204);
and U10277 (N_10277,N_10160,N_10222);
xnor U10278 (N_10278,N_10089,N_10157);
nand U10279 (N_10279,N_10082,N_10112);
nand U10280 (N_10280,N_10101,N_10238);
nor U10281 (N_10281,N_10158,N_10136);
xor U10282 (N_10282,N_10098,N_10111);
nand U10283 (N_10283,N_10198,N_10197);
nand U10284 (N_10284,N_10177,N_10219);
nor U10285 (N_10285,N_10185,N_10161);
nand U10286 (N_10286,N_10208,N_10137);
or U10287 (N_10287,N_10170,N_10104);
and U10288 (N_10288,N_10159,N_10236);
or U10289 (N_10289,N_10133,N_10122);
and U10290 (N_10290,N_10220,N_10091);
and U10291 (N_10291,N_10216,N_10217);
nand U10292 (N_10292,N_10224,N_10206);
nand U10293 (N_10293,N_10232,N_10126);
or U10294 (N_10294,N_10181,N_10149);
and U10295 (N_10295,N_10164,N_10150);
or U10296 (N_10296,N_10214,N_10151);
and U10297 (N_10297,N_10189,N_10097);
and U10298 (N_10298,N_10120,N_10184);
or U10299 (N_10299,N_10168,N_10233);
nor U10300 (N_10300,N_10162,N_10171);
nor U10301 (N_10301,N_10178,N_10202);
nand U10302 (N_10302,N_10175,N_10165);
nor U10303 (N_10303,N_10106,N_10169);
nor U10304 (N_10304,N_10086,N_10215);
xnor U10305 (N_10305,N_10211,N_10147);
and U10306 (N_10306,N_10230,N_10140);
nor U10307 (N_10307,N_10105,N_10179);
nand U10308 (N_10308,N_10145,N_10231);
nor U10309 (N_10309,N_10083,N_10227);
xnor U10310 (N_10310,N_10095,N_10188);
or U10311 (N_10311,N_10176,N_10148);
xor U10312 (N_10312,N_10131,N_10088);
xnor U10313 (N_10313,N_10109,N_10174);
or U10314 (N_10314,N_10212,N_10094);
or U10315 (N_10315,N_10081,N_10187);
nor U10316 (N_10316,N_10183,N_10199);
nor U10317 (N_10317,N_10092,N_10221);
nor U10318 (N_10318,N_10096,N_10138);
xnor U10319 (N_10319,N_10153,N_10132);
and U10320 (N_10320,N_10127,N_10170);
and U10321 (N_10321,N_10210,N_10201);
or U10322 (N_10322,N_10237,N_10162);
xor U10323 (N_10323,N_10206,N_10098);
or U10324 (N_10324,N_10201,N_10138);
xnor U10325 (N_10325,N_10230,N_10195);
xor U10326 (N_10326,N_10181,N_10176);
nand U10327 (N_10327,N_10212,N_10169);
and U10328 (N_10328,N_10130,N_10206);
or U10329 (N_10329,N_10183,N_10216);
or U10330 (N_10330,N_10166,N_10150);
xnor U10331 (N_10331,N_10139,N_10122);
nor U10332 (N_10332,N_10210,N_10165);
or U10333 (N_10333,N_10138,N_10100);
nand U10334 (N_10334,N_10137,N_10132);
nand U10335 (N_10335,N_10190,N_10156);
xor U10336 (N_10336,N_10104,N_10198);
and U10337 (N_10337,N_10227,N_10201);
xnor U10338 (N_10338,N_10086,N_10093);
nor U10339 (N_10339,N_10216,N_10182);
or U10340 (N_10340,N_10135,N_10239);
nand U10341 (N_10341,N_10131,N_10155);
nor U10342 (N_10342,N_10194,N_10147);
and U10343 (N_10343,N_10207,N_10120);
xor U10344 (N_10344,N_10174,N_10086);
xnor U10345 (N_10345,N_10098,N_10162);
and U10346 (N_10346,N_10165,N_10220);
nor U10347 (N_10347,N_10148,N_10195);
xnor U10348 (N_10348,N_10234,N_10215);
nand U10349 (N_10349,N_10133,N_10107);
or U10350 (N_10350,N_10130,N_10144);
and U10351 (N_10351,N_10171,N_10093);
nor U10352 (N_10352,N_10097,N_10107);
nand U10353 (N_10353,N_10191,N_10195);
xor U10354 (N_10354,N_10132,N_10215);
xnor U10355 (N_10355,N_10222,N_10094);
nor U10356 (N_10356,N_10172,N_10188);
xor U10357 (N_10357,N_10235,N_10106);
or U10358 (N_10358,N_10169,N_10191);
nor U10359 (N_10359,N_10120,N_10224);
xnor U10360 (N_10360,N_10235,N_10200);
or U10361 (N_10361,N_10218,N_10215);
nand U10362 (N_10362,N_10082,N_10230);
nand U10363 (N_10363,N_10239,N_10238);
or U10364 (N_10364,N_10231,N_10113);
or U10365 (N_10365,N_10107,N_10195);
xor U10366 (N_10366,N_10132,N_10187);
or U10367 (N_10367,N_10115,N_10095);
xor U10368 (N_10368,N_10183,N_10096);
and U10369 (N_10369,N_10222,N_10100);
or U10370 (N_10370,N_10120,N_10200);
or U10371 (N_10371,N_10145,N_10115);
nor U10372 (N_10372,N_10205,N_10158);
nor U10373 (N_10373,N_10217,N_10121);
nor U10374 (N_10374,N_10216,N_10108);
and U10375 (N_10375,N_10217,N_10203);
nand U10376 (N_10376,N_10184,N_10115);
xor U10377 (N_10377,N_10125,N_10122);
nor U10378 (N_10378,N_10110,N_10186);
or U10379 (N_10379,N_10085,N_10082);
and U10380 (N_10380,N_10191,N_10151);
xnor U10381 (N_10381,N_10165,N_10204);
xnor U10382 (N_10382,N_10088,N_10083);
or U10383 (N_10383,N_10085,N_10132);
xnor U10384 (N_10384,N_10147,N_10093);
or U10385 (N_10385,N_10096,N_10092);
nor U10386 (N_10386,N_10195,N_10238);
nor U10387 (N_10387,N_10143,N_10166);
xnor U10388 (N_10388,N_10096,N_10152);
or U10389 (N_10389,N_10181,N_10202);
nor U10390 (N_10390,N_10154,N_10113);
or U10391 (N_10391,N_10148,N_10228);
or U10392 (N_10392,N_10123,N_10158);
or U10393 (N_10393,N_10123,N_10178);
or U10394 (N_10394,N_10229,N_10231);
nand U10395 (N_10395,N_10095,N_10111);
xor U10396 (N_10396,N_10221,N_10142);
nor U10397 (N_10397,N_10102,N_10101);
or U10398 (N_10398,N_10095,N_10144);
xor U10399 (N_10399,N_10232,N_10084);
xor U10400 (N_10400,N_10352,N_10266);
nor U10401 (N_10401,N_10304,N_10344);
nor U10402 (N_10402,N_10337,N_10382);
xor U10403 (N_10403,N_10245,N_10347);
or U10404 (N_10404,N_10321,N_10395);
and U10405 (N_10405,N_10380,N_10293);
and U10406 (N_10406,N_10389,N_10392);
nand U10407 (N_10407,N_10251,N_10305);
nor U10408 (N_10408,N_10353,N_10354);
and U10409 (N_10409,N_10390,N_10396);
or U10410 (N_10410,N_10250,N_10265);
xor U10411 (N_10411,N_10334,N_10270);
and U10412 (N_10412,N_10268,N_10296);
nor U10413 (N_10413,N_10246,N_10357);
or U10414 (N_10414,N_10288,N_10342);
xnor U10415 (N_10415,N_10303,N_10370);
or U10416 (N_10416,N_10279,N_10284);
xor U10417 (N_10417,N_10257,N_10322);
or U10418 (N_10418,N_10379,N_10281);
xor U10419 (N_10419,N_10289,N_10325);
nand U10420 (N_10420,N_10394,N_10253);
xnor U10421 (N_10421,N_10367,N_10377);
and U10422 (N_10422,N_10248,N_10328);
xor U10423 (N_10423,N_10378,N_10241);
xor U10424 (N_10424,N_10261,N_10323);
or U10425 (N_10425,N_10286,N_10326);
nor U10426 (N_10426,N_10359,N_10332);
nor U10427 (N_10427,N_10391,N_10329);
xor U10428 (N_10428,N_10276,N_10338);
and U10429 (N_10429,N_10356,N_10311);
and U10430 (N_10430,N_10383,N_10315);
nor U10431 (N_10431,N_10307,N_10282);
nand U10432 (N_10432,N_10361,N_10297);
xor U10433 (N_10433,N_10339,N_10256);
and U10434 (N_10434,N_10277,N_10280);
xor U10435 (N_10435,N_10310,N_10318);
nor U10436 (N_10436,N_10316,N_10317);
nor U10437 (N_10437,N_10386,N_10376);
nand U10438 (N_10438,N_10381,N_10243);
or U10439 (N_10439,N_10292,N_10373);
xnor U10440 (N_10440,N_10341,N_10301);
and U10441 (N_10441,N_10247,N_10385);
and U10442 (N_10442,N_10324,N_10267);
nand U10443 (N_10443,N_10388,N_10327);
and U10444 (N_10444,N_10375,N_10313);
and U10445 (N_10445,N_10308,N_10249);
or U10446 (N_10446,N_10336,N_10252);
or U10447 (N_10447,N_10393,N_10331);
xnor U10448 (N_10448,N_10351,N_10312);
nand U10449 (N_10449,N_10320,N_10369);
xnor U10450 (N_10450,N_10285,N_10355);
or U10451 (N_10451,N_10242,N_10309);
or U10452 (N_10452,N_10299,N_10349);
xor U10453 (N_10453,N_10366,N_10291);
and U10454 (N_10454,N_10374,N_10368);
or U10455 (N_10455,N_10290,N_10263);
and U10456 (N_10456,N_10314,N_10274);
and U10457 (N_10457,N_10371,N_10269);
or U10458 (N_10458,N_10259,N_10255);
nor U10459 (N_10459,N_10262,N_10260);
or U10460 (N_10460,N_10294,N_10302);
nand U10461 (N_10461,N_10346,N_10330);
nand U10462 (N_10462,N_10319,N_10399);
nor U10463 (N_10463,N_10363,N_10275);
and U10464 (N_10464,N_10340,N_10358);
and U10465 (N_10465,N_10273,N_10372);
or U10466 (N_10466,N_10244,N_10365);
or U10467 (N_10467,N_10387,N_10306);
or U10468 (N_10468,N_10335,N_10283);
nor U10469 (N_10469,N_10348,N_10364);
xor U10470 (N_10470,N_10343,N_10240);
nor U10471 (N_10471,N_10272,N_10362);
xnor U10472 (N_10472,N_10254,N_10295);
xnor U10473 (N_10473,N_10360,N_10264);
nand U10474 (N_10474,N_10397,N_10287);
nand U10475 (N_10475,N_10258,N_10298);
and U10476 (N_10476,N_10271,N_10345);
and U10477 (N_10477,N_10278,N_10384);
or U10478 (N_10478,N_10350,N_10333);
nor U10479 (N_10479,N_10300,N_10398);
nand U10480 (N_10480,N_10297,N_10372);
or U10481 (N_10481,N_10351,N_10276);
nor U10482 (N_10482,N_10359,N_10306);
nand U10483 (N_10483,N_10383,N_10385);
and U10484 (N_10484,N_10367,N_10359);
and U10485 (N_10485,N_10267,N_10332);
or U10486 (N_10486,N_10295,N_10353);
and U10487 (N_10487,N_10315,N_10294);
and U10488 (N_10488,N_10389,N_10310);
nor U10489 (N_10489,N_10300,N_10373);
nor U10490 (N_10490,N_10343,N_10364);
xor U10491 (N_10491,N_10398,N_10372);
or U10492 (N_10492,N_10329,N_10281);
nor U10493 (N_10493,N_10399,N_10291);
nand U10494 (N_10494,N_10386,N_10287);
nor U10495 (N_10495,N_10258,N_10259);
nand U10496 (N_10496,N_10263,N_10289);
and U10497 (N_10497,N_10245,N_10312);
nor U10498 (N_10498,N_10385,N_10384);
and U10499 (N_10499,N_10367,N_10257);
nand U10500 (N_10500,N_10398,N_10378);
nand U10501 (N_10501,N_10342,N_10378);
xnor U10502 (N_10502,N_10305,N_10373);
xnor U10503 (N_10503,N_10339,N_10281);
or U10504 (N_10504,N_10310,N_10366);
nor U10505 (N_10505,N_10287,N_10249);
xnor U10506 (N_10506,N_10294,N_10260);
or U10507 (N_10507,N_10243,N_10369);
xor U10508 (N_10508,N_10350,N_10292);
nor U10509 (N_10509,N_10241,N_10272);
nor U10510 (N_10510,N_10279,N_10354);
xor U10511 (N_10511,N_10305,N_10273);
nor U10512 (N_10512,N_10358,N_10259);
nand U10513 (N_10513,N_10383,N_10285);
and U10514 (N_10514,N_10270,N_10346);
nand U10515 (N_10515,N_10307,N_10253);
nor U10516 (N_10516,N_10252,N_10359);
and U10517 (N_10517,N_10358,N_10347);
xnor U10518 (N_10518,N_10249,N_10375);
xor U10519 (N_10519,N_10251,N_10252);
and U10520 (N_10520,N_10376,N_10340);
nor U10521 (N_10521,N_10247,N_10331);
xnor U10522 (N_10522,N_10270,N_10343);
nand U10523 (N_10523,N_10380,N_10357);
nand U10524 (N_10524,N_10356,N_10302);
and U10525 (N_10525,N_10358,N_10280);
and U10526 (N_10526,N_10372,N_10265);
or U10527 (N_10527,N_10310,N_10390);
nor U10528 (N_10528,N_10323,N_10242);
nor U10529 (N_10529,N_10299,N_10297);
or U10530 (N_10530,N_10285,N_10330);
xnor U10531 (N_10531,N_10299,N_10298);
or U10532 (N_10532,N_10255,N_10254);
nand U10533 (N_10533,N_10352,N_10247);
xnor U10534 (N_10534,N_10373,N_10375);
and U10535 (N_10535,N_10387,N_10389);
nand U10536 (N_10536,N_10352,N_10251);
or U10537 (N_10537,N_10367,N_10328);
and U10538 (N_10538,N_10397,N_10252);
xnor U10539 (N_10539,N_10273,N_10306);
nand U10540 (N_10540,N_10274,N_10360);
and U10541 (N_10541,N_10326,N_10244);
nand U10542 (N_10542,N_10353,N_10362);
and U10543 (N_10543,N_10247,N_10272);
and U10544 (N_10544,N_10262,N_10265);
nor U10545 (N_10545,N_10391,N_10338);
and U10546 (N_10546,N_10366,N_10385);
xnor U10547 (N_10547,N_10296,N_10346);
or U10548 (N_10548,N_10257,N_10397);
nor U10549 (N_10549,N_10315,N_10346);
or U10550 (N_10550,N_10312,N_10276);
and U10551 (N_10551,N_10309,N_10284);
nand U10552 (N_10552,N_10327,N_10369);
nand U10553 (N_10553,N_10276,N_10324);
and U10554 (N_10554,N_10242,N_10339);
or U10555 (N_10555,N_10277,N_10275);
nand U10556 (N_10556,N_10372,N_10361);
nor U10557 (N_10557,N_10371,N_10284);
or U10558 (N_10558,N_10335,N_10365);
nand U10559 (N_10559,N_10303,N_10391);
or U10560 (N_10560,N_10429,N_10418);
and U10561 (N_10561,N_10458,N_10546);
nor U10562 (N_10562,N_10547,N_10485);
xnor U10563 (N_10563,N_10466,N_10433);
nor U10564 (N_10564,N_10515,N_10488);
and U10565 (N_10565,N_10413,N_10494);
and U10566 (N_10566,N_10405,N_10506);
nand U10567 (N_10567,N_10513,N_10415);
and U10568 (N_10568,N_10441,N_10412);
xnor U10569 (N_10569,N_10540,N_10554);
xor U10570 (N_10570,N_10519,N_10472);
nand U10571 (N_10571,N_10423,N_10500);
and U10572 (N_10572,N_10460,N_10509);
nor U10573 (N_10573,N_10463,N_10437);
nand U10574 (N_10574,N_10420,N_10447);
or U10575 (N_10575,N_10422,N_10439);
nor U10576 (N_10576,N_10473,N_10409);
nor U10577 (N_10577,N_10480,N_10446);
and U10578 (N_10578,N_10482,N_10402);
and U10579 (N_10579,N_10407,N_10449);
xor U10580 (N_10580,N_10531,N_10529);
or U10581 (N_10581,N_10465,N_10468);
nor U10582 (N_10582,N_10470,N_10455);
or U10583 (N_10583,N_10490,N_10428);
and U10584 (N_10584,N_10448,N_10510);
and U10585 (N_10585,N_10450,N_10533);
xor U10586 (N_10586,N_10404,N_10414);
nand U10587 (N_10587,N_10499,N_10431);
and U10588 (N_10588,N_10477,N_10551);
nand U10589 (N_10589,N_10436,N_10442);
nor U10590 (N_10590,N_10538,N_10524);
or U10591 (N_10591,N_10400,N_10459);
nand U10592 (N_10592,N_10556,N_10421);
and U10593 (N_10593,N_10495,N_10406);
xor U10594 (N_10594,N_10545,N_10511);
or U10595 (N_10595,N_10501,N_10528);
nand U10596 (N_10596,N_10497,N_10474);
and U10597 (N_10597,N_10464,N_10507);
or U10598 (N_10598,N_10539,N_10430);
or U10599 (N_10599,N_10486,N_10557);
or U10600 (N_10600,N_10553,N_10516);
nand U10601 (N_10601,N_10552,N_10536);
or U10602 (N_10602,N_10419,N_10491);
xor U10603 (N_10603,N_10457,N_10445);
and U10604 (N_10604,N_10481,N_10403);
and U10605 (N_10605,N_10503,N_10426);
xnor U10606 (N_10606,N_10549,N_10479);
nor U10607 (N_10607,N_10434,N_10461);
nor U10608 (N_10608,N_10537,N_10526);
and U10609 (N_10609,N_10559,N_10416);
and U10610 (N_10610,N_10514,N_10476);
nand U10611 (N_10611,N_10454,N_10471);
and U10612 (N_10612,N_10462,N_10475);
and U10613 (N_10613,N_10489,N_10492);
and U10614 (N_10614,N_10408,N_10544);
xnor U10615 (N_10615,N_10532,N_10496);
and U10616 (N_10616,N_10487,N_10543);
nand U10617 (N_10617,N_10411,N_10425);
or U10618 (N_10618,N_10484,N_10440);
nor U10619 (N_10619,N_10525,N_10558);
nor U10620 (N_10620,N_10438,N_10530);
and U10621 (N_10621,N_10534,N_10417);
nor U10622 (N_10622,N_10523,N_10444);
or U10623 (N_10623,N_10451,N_10467);
nor U10624 (N_10624,N_10520,N_10410);
xnor U10625 (N_10625,N_10401,N_10508);
or U10626 (N_10626,N_10427,N_10443);
and U10627 (N_10627,N_10527,N_10535);
nand U10628 (N_10628,N_10517,N_10453);
xnor U10629 (N_10629,N_10456,N_10469);
and U10630 (N_10630,N_10483,N_10521);
and U10631 (N_10631,N_10502,N_10555);
or U10632 (N_10632,N_10424,N_10505);
or U10633 (N_10633,N_10542,N_10541);
nand U10634 (N_10634,N_10512,N_10435);
nor U10635 (N_10635,N_10452,N_10518);
and U10636 (N_10636,N_10478,N_10548);
and U10637 (N_10637,N_10522,N_10550);
xor U10638 (N_10638,N_10493,N_10504);
nand U10639 (N_10639,N_10432,N_10498);
or U10640 (N_10640,N_10527,N_10420);
or U10641 (N_10641,N_10413,N_10507);
nor U10642 (N_10642,N_10476,N_10541);
and U10643 (N_10643,N_10445,N_10498);
nor U10644 (N_10644,N_10426,N_10523);
or U10645 (N_10645,N_10450,N_10428);
nor U10646 (N_10646,N_10488,N_10463);
xor U10647 (N_10647,N_10432,N_10491);
and U10648 (N_10648,N_10491,N_10550);
and U10649 (N_10649,N_10415,N_10553);
nand U10650 (N_10650,N_10418,N_10518);
and U10651 (N_10651,N_10476,N_10406);
or U10652 (N_10652,N_10449,N_10442);
and U10653 (N_10653,N_10423,N_10554);
nand U10654 (N_10654,N_10499,N_10519);
and U10655 (N_10655,N_10428,N_10423);
xor U10656 (N_10656,N_10407,N_10524);
nand U10657 (N_10657,N_10472,N_10424);
or U10658 (N_10658,N_10509,N_10499);
nor U10659 (N_10659,N_10450,N_10439);
xor U10660 (N_10660,N_10442,N_10556);
nor U10661 (N_10661,N_10516,N_10489);
or U10662 (N_10662,N_10421,N_10455);
nand U10663 (N_10663,N_10512,N_10404);
and U10664 (N_10664,N_10483,N_10465);
nor U10665 (N_10665,N_10544,N_10543);
nor U10666 (N_10666,N_10450,N_10527);
xor U10667 (N_10667,N_10553,N_10500);
nor U10668 (N_10668,N_10499,N_10546);
or U10669 (N_10669,N_10478,N_10480);
and U10670 (N_10670,N_10448,N_10408);
nor U10671 (N_10671,N_10505,N_10461);
xnor U10672 (N_10672,N_10515,N_10417);
nand U10673 (N_10673,N_10554,N_10402);
or U10674 (N_10674,N_10489,N_10403);
or U10675 (N_10675,N_10437,N_10540);
xor U10676 (N_10676,N_10453,N_10442);
nand U10677 (N_10677,N_10437,N_10556);
nand U10678 (N_10678,N_10535,N_10432);
nor U10679 (N_10679,N_10416,N_10466);
nand U10680 (N_10680,N_10557,N_10501);
nor U10681 (N_10681,N_10463,N_10446);
xnor U10682 (N_10682,N_10414,N_10443);
nor U10683 (N_10683,N_10553,N_10432);
nor U10684 (N_10684,N_10442,N_10407);
nand U10685 (N_10685,N_10529,N_10449);
or U10686 (N_10686,N_10520,N_10482);
or U10687 (N_10687,N_10478,N_10474);
or U10688 (N_10688,N_10447,N_10409);
xnor U10689 (N_10689,N_10428,N_10554);
xnor U10690 (N_10690,N_10450,N_10401);
nand U10691 (N_10691,N_10522,N_10555);
nand U10692 (N_10692,N_10489,N_10538);
nand U10693 (N_10693,N_10545,N_10442);
and U10694 (N_10694,N_10472,N_10446);
xor U10695 (N_10695,N_10470,N_10450);
and U10696 (N_10696,N_10523,N_10538);
nor U10697 (N_10697,N_10435,N_10453);
or U10698 (N_10698,N_10434,N_10538);
xnor U10699 (N_10699,N_10404,N_10495);
or U10700 (N_10700,N_10530,N_10409);
nand U10701 (N_10701,N_10437,N_10499);
or U10702 (N_10702,N_10422,N_10465);
or U10703 (N_10703,N_10475,N_10476);
nor U10704 (N_10704,N_10521,N_10518);
nand U10705 (N_10705,N_10481,N_10413);
nand U10706 (N_10706,N_10529,N_10540);
or U10707 (N_10707,N_10522,N_10536);
or U10708 (N_10708,N_10479,N_10512);
or U10709 (N_10709,N_10408,N_10436);
and U10710 (N_10710,N_10432,N_10508);
nor U10711 (N_10711,N_10545,N_10541);
and U10712 (N_10712,N_10549,N_10539);
xor U10713 (N_10713,N_10512,N_10496);
and U10714 (N_10714,N_10508,N_10529);
nor U10715 (N_10715,N_10501,N_10489);
nand U10716 (N_10716,N_10477,N_10447);
xor U10717 (N_10717,N_10460,N_10449);
xnor U10718 (N_10718,N_10548,N_10432);
xnor U10719 (N_10719,N_10414,N_10415);
or U10720 (N_10720,N_10619,N_10626);
nand U10721 (N_10721,N_10583,N_10591);
nand U10722 (N_10722,N_10633,N_10646);
and U10723 (N_10723,N_10699,N_10610);
or U10724 (N_10724,N_10623,N_10625);
nor U10725 (N_10725,N_10638,N_10664);
nor U10726 (N_10726,N_10644,N_10624);
and U10727 (N_10727,N_10595,N_10585);
nand U10728 (N_10728,N_10598,N_10620);
and U10729 (N_10729,N_10715,N_10695);
and U10730 (N_10730,N_10661,N_10629);
or U10731 (N_10731,N_10580,N_10670);
nor U10732 (N_10732,N_10650,N_10667);
xor U10733 (N_10733,N_10703,N_10679);
nor U10734 (N_10734,N_10600,N_10683);
or U10735 (N_10735,N_10645,N_10608);
or U10736 (N_10736,N_10607,N_10617);
xor U10737 (N_10737,N_10618,N_10631);
nand U10738 (N_10738,N_10665,N_10563);
or U10739 (N_10739,N_10671,N_10592);
and U10740 (N_10740,N_10606,N_10615);
nand U10741 (N_10741,N_10565,N_10637);
nand U10742 (N_10742,N_10704,N_10584);
nor U10743 (N_10743,N_10652,N_10682);
and U10744 (N_10744,N_10604,N_10611);
xnor U10745 (N_10745,N_10696,N_10678);
nor U10746 (N_10746,N_10694,N_10590);
nand U10747 (N_10747,N_10668,N_10709);
nor U10748 (N_10748,N_10711,N_10564);
and U10749 (N_10749,N_10647,N_10675);
nor U10750 (N_10750,N_10577,N_10690);
xnor U10751 (N_10751,N_10573,N_10693);
nand U10752 (N_10752,N_10659,N_10594);
and U10753 (N_10753,N_10685,N_10660);
nand U10754 (N_10754,N_10642,N_10691);
xnor U10755 (N_10755,N_10640,N_10621);
or U10756 (N_10756,N_10614,N_10634);
xnor U10757 (N_10757,N_10578,N_10639);
nor U10758 (N_10758,N_10700,N_10666);
or U10759 (N_10759,N_10609,N_10663);
or U10760 (N_10760,N_10713,N_10651);
nor U10761 (N_10761,N_10605,N_10662);
and U10762 (N_10762,N_10586,N_10576);
nor U10763 (N_10763,N_10687,N_10658);
and U10764 (N_10764,N_10599,N_10697);
xor U10765 (N_10765,N_10574,N_10602);
or U10766 (N_10766,N_10569,N_10648);
or U10767 (N_10767,N_10588,N_10561);
nor U10768 (N_10768,N_10702,N_10701);
nand U10769 (N_10769,N_10688,N_10673);
nand U10770 (N_10770,N_10567,N_10575);
xor U10771 (N_10771,N_10689,N_10601);
nand U10772 (N_10772,N_10714,N_10566);
nor U10773 (N_10773,N_10669,N_10716);
nand U10774 (N_10774,N_10719,N_10692);
or U10775 (N_10775,N_10581,N_10705);
nor U10776 (N_10776,N_10622,N_10657);
or U10777 (N_10777,N_10717,N_10718);
and U10778 (N_10778,N_10636,N_10707);
nor U10779 (N_10779,N_10616,N_10686);
or U10780 (N_10780,N_10649,N_10684);
nand U10781 (N_10781,N_10708,N_10653);
and U10782 (N_10782,N_10572,N_10656);
nor U10783 (N_10783,N_10641,N_10672);
or U10784 (N_10784,N_10560,N_10632);
or U10785 (N_10785,N_10579,N_10712);
nor U10786 (N_10786,N_10643,N_10562);
nand U10787 (N_10787,N_10654,N_10570);
nor U10788 (N_10788,N_10597,N_10677);
nand U10789 (N_10789,N_10613,N_10571);
xor U10790 (N_10790,N_10706,N_10674);
and U10791 (N_10791,N_10582,N_10596);
and U10792 (N_10792,N_10628,N_10698);
nor U10793 (N_10793,N_10710,N_10681);
and U10794 (N_10794,N_10603,N_10627);
or U10795 (N_10795,N_10589,N_10568);
xnor U10796 (N_10796,N_10612,N_10655);
xnor U10797 (N_10797,N_10587,N_10593);
xnor U10798 (N_10798,N_10635,N_10680);
xor U10799 (N_10799,N_10630,N_10676);
or U10800 (N_10800,N_10708,N_10581);
and U10801 (N_10801,N_10700,N_10590);
nand U10802 (N_10802,N_10712,N_10696);
nand U10803 (N_10803,N_10626,N_10709);
xor U10804 (N_10804,N_10691,N_10635);
or U10805 (N_10805,N_10587,N_10573);
and U10806 (N_10806,N_10573,N_10714);
or U10807 (N_10807,N_10585,N_10619);
or U10808 (N_10808,N_10639,N_10667);
and U10809 (N_10809,N_10715,N_10645);
nor U10810 (N_10810,N_10567,N_10607);
or U10811 (N_10811,N_10590,N_10689);
nand U10812 (N_10812,N_10630,N_10642);
nor U10813 (N_10813,N_10716,N_10677);
nor U10814 (N_10814,N_10565,N_10580);
nor U10815 (N_10815,N_10623,N_10597);
xnor U10816 (N_10816,N_10578,N_10615);
nor U10817 (N_10817,N_10659,N_10698);
nor U10818 (N_10818,N_10637,N_10688);
and U10819 (N_10819,N_10699,N_10593);
nor U10820 (N_10820,N_10654,N_10602);
xnor U10821 (N_10821,N_10702,N_10607);
xor U10822 (N_10822,N_10571,N_10674);
nand U10823 (N_10823,N_10706,N_10612);
xnor U10824 (N_10824,N_10571,N_10628);
and U10825 (N_10825,N_10581,N_10696);
and U10826 (N_10826,N_10667,N_10654);
nor U10827 (N_10827,N_10634,N_10701);
nand U10828 (N_10828,N_10632,N_10565);
and U10829 (N_10829,N_10571,N_10704);
or U10830 (N_10830,N_10611,N_10607);
nand U10831 (N_10831,N_10601,N_10684);
xor U10832 (N_10832,N_10577,N_10627);
and U10833 (N_10833,N_10690,N_10695);
nor U10834 (N_10834,N_10572,N_10668);
nor U10835 (N_10835,N_10702,N_10719);
and U10836 (N_10836,N_10563,N_10580);
xnor U10837 (N_10837,N_10702,N_10621);
xnor U10838 (N_10838,N_10635,N_10699);
or U10839 (N_10839,N_10572,N_10613);
nor U10840 (N_10840,N_10616,N_10640);
xnor U10841 (N_10841,N_10635,N_10715);
nor U10842 (N_10842,N_10683,N_10617);
nand U10843 (N_10843,N_10620,N_10633);
nand U10844 (N_10844,N_10563,N_10610);
nand U10845 (N_10845,N_10593,N_10648);
nand U10846 (N_10846,N_10590,N_10668);
xor U10847 (N_10847,N_10671,N_10591);
or U10848 (N_10848,N_10618,N_10676);
xor U10849 (N_10849,N_10659,N_10706);
and U10850 (N_10850,N_10629,N_10711);
nor U10851 (N_10851,N_10600,N_10667);
xor U10852 (N_10852,N_10701,N_10649);
and U10853 (N_10853,N_10697,N_10685);
xnor U10854 (N_10854,N_10688,N_10616);
or U10855 (N_10855,N_10583,N_10589);
nor U10856 (N_10856,N_10634,N_10627);
or U10857 (N_10857,N_10697,N_10705);
and U10858 (N_10858,N_10669,N_10663);
xor U10859 (N_10859,N_10646,N_10650);
nor U10860 (N_10860,N_10651,N_10680);
or U10861 (N_10861,N_10675,N_10570);
or U10862 (N_10862,N_10627,N_10653);
nor U10863 (N_10863,N_10600,N_10588);
nor U10864 (N_10864,N_10627,N_10584);
nor U10865 (N_10865,N_10562,N_10572);
and U10866 (N_10866,N_10651,N_10665);
or U10867 (N_10867,N_10628,N_10693);
xnor U10868 (N_10868,N_10636,N_10580);
or U10869 (N_10869,N_10570,N_10657);
and U10870 (N_10870,N_10636,N_10695);
nor U10871 (N_10871,N_10571,N_10635);
and U10872 (N_10872,N_10581,N_10615);
nor U10873 (N_10873,N_10673,N_10573);
nor U10874 (N_10874,N_10662,N_10595);
and U10875 (N_10875,N_10591,N_10666);
and U10876 (N_10876,N_10714,N_10686);
nand U10877 (N_10877,N_10642,N_10697);
or U10878 (N_10878,N_10682,N_10639);
nor U10879 (N_10879,N_10649,N_10678);
or U10880 (N_10880,N_10812,N_10806);
or U10881 (N_10881,N_10784,N_10803);
nand U10882 (N_10882,N_10732,N_10792);
xnor U10883 (N_10883,N_10870,N_10721);
or U10884 (N_10884,N_10733,N_10727);
nand U10885 (N_10885,N_10864,N_10755);
nor U10886 (N_10886,N_10794,N_10807);
xor U10887 (N_10887,N_10742,N_10796);
xnor U10888 (N_10888,N_10772,N_10723);
or U10889 (N_10889,N_10827,N_10730);
xor U10890 (N_10890,N_10797,N_10722);
or U10891 (N_10891,N_10801,N_10878);
xnor U10892 (N_10892,N_10767,N_10759);
and U10893 (N_10893,N_10778,N_10773);
and U10894 (N_10894,N_10737,N_10833);
nor U10895 (N_10895,N_10775,N_10853);
xor U10896 (N_10896,N_10795,N_10808);
or U10897 (N_10897,N_10758,N_10751);
xnor U10898 (N_10898,N_10877,N_10834);
nand U10899 (N_10899,N_10749,N_10821);
xnor U10900 (N_10900,N_10862,N_10846);
or U10901 (N_10901,N_10843,N_10875);
nor U10902 (N_10902,N_10844,N_10860);
xnor U10903 (N_10903,N_10728,N_10850);
xor U10904 (N_10904,N_10774,N_10817);
nor U10905 (N_10905,N_10836,N_10861);
xor U10906 (N_10906,N_10872,N_10815);
nand U10907 (N_10907,N_10859,N_10819);
and U10908 (N_10908,N_10824,N_10735);
nand U10909 (N_10909,N_10873,N_10771);
nand U10910 (N_10910,N_10828,N_10766);
and U10911 (N_10911,N_10837,N_10804);
xnor U10912 (N_10912,N_10842,N_10743);
nand U10913 (N_10913,N_10813,N_10830);
nor U10914 (N_10914,N_10740,N_10825);
xnor U10915 (N_10915,N_10845,N_10776);
nand U10916 (N_10916,N_10726,N_10805);
xor U10917 (N_10917,N_10770,N_10752);
and U10918 (N_10918,N_10782,N_10764);
xnor U10919 (N_10919,N_10793,N_10777);
xor U10920 (N_10920,N_10851,N_10787);
or U10921 (N_10921,N_10823,N_10832);
nor U10922 (N_10922,N_10754,N_10788);
xor U10923 (N_10923,N_10783,N_10762);
and U10924 (N_10924,N_10857,N_10854);
and U10925 (N_10925,N_10786,N_10798);
or U10926 (N_10926,N_10757,N_10763);
xnor U10927 (N_10927,N_10816,N_10879);
nand U10928 (N_10928,N_10781,N_10856);
or U10929 (N_10929,N_10829,N_10747);
nand U10930 (N_10930,N_10848,N_10741);
xnor U10931 (N_10931,N_10809,N_10820);
nor U10932 (N_10932,N_10736,N_10826);
nand U10933 (N_10933,N_10866,N_10799);
nor U10934 (N_10934,N_10849,N_10818);
and U10935 (N_10935,N_10847,N_10761);
xor U10936 (N_10936,N_10725,N_10756);
or U10937 (N_10937,N_10779,N_10789);
nand U10938 (N_10938,N_10791,N_10852);
xnor U10939 (N_10939,N_10760,N_10768);
nand U10940 (N_10940,N_10876,N_10744);
and U10941 (N_10941,N_10871,N_10748);
xnor U10942 (N_10942,N_10769,N_10811);
xor U10943 (N_10943,N_10822,N_10734);
xor U10944 (N_10944,N_10865,N_10802);
or U10945 (N_10945,N_10731,N_10863);
and U10946 (N_10946,N_10738,N_10858);
nor U10947 (N_10947,N_10800,N_10780);
nand U10948 (N_10948,N_10720,N_10874);
nor U10949 (N_10949,N_10785,N_10868);
nand U10950 (N_10950,N_10724,N_10746);
or U10951 (N_10951,N_10790,N_10814);
nor U10952 (N_10952,N_10835,N_10745);
nand U10953 (N_10953,N_10838,N_10765);
or U10954 (N_10954,N_10729,N_10855);
or U10955 (N_10955,N_10839,N_10831);
and U10956 (N_10956,N_10750,N_10810);
or U10957 (N_10957,N_10840,N_10753);
or U10958 (N_10958,N_10869,N_10841);
nand U10959 (N_10959,N_10867,N_10739);
or U10960 (N_10960,N_10857,N_10749);
nand U10961 (N_10961,N_10857,N_10775);
nand U10962 (N_10962,N_10823,N_10743);
xnor U10963 (N_10963,N_10861,N_10872);
nand U10964 (N_10964,N_10805,N_10817);
xor U10965 (N_10965,N_10831,N_10836);
or U10966 (N_10966,N_10844,N_10746);
nand U10967 (N_10967,N_10787,N_10794);
and U10968 (N_10968,N_10772,N_10796);
and U10969 (N_10969,N_10857,N_10753);
xnor U10970 (N_10970,N_10822,N_10747);
and U10971 (N_10971,N_10757,N_10768);
nor U10972 (N_10972,N_10848,N_10792);
or U10973 (N_10973,N_10773,N_10768);
or U10974 (N_10974,N_10821,N_10817);
or U10975 (N_10975,N_10767,N_10738);
nand U10976 (N_10976,N_10869,N_10874);
nand U10977 (N_10977,N_10788,N_10766);
nand U10978 (N_10978,N_10861,N_10764);
xor U10979 (N_10979,N_10780,N_10721);
and U10980 (N_10980,N_10784,N_10829);
and U10981 (N_10981,N_10820,N_10862);
nor U10982 (N_10982,N_10720,N_10824);
nand U10983 (N_10983,N_10783,N_10724);
nor U10984 (N_10984,N_10771,N_10824);
or U10985 (N_10985,N_10870,N_10835);
or U10986 (N_10986,N_10814,N_10849);
nor U10987 (N_10987,N_10860,N_10825);
nand U10988 (N_10988,N_10796,N_10732);
nor U10989 (N_10989,N_10751,N_10813);
xnor U10990 (N_10990,N_10755,N_10826);
nand U10991 (N_10991,N_10819,N_10845);
and U10992 (N_10992,N_10803,N_10754);
xnor U10993 (N_10993,N_10854,N_10802);
xnor U10994 (N_10994,N_10752,N_10875);
xnor U10995 (N_10995,N_10744,N_10868);
xnor U10996 (N_10996,N_10724,N_10735);
or U10997 (N_10997,N_10839,N_10830);
nor U10998 (N_10998,N_10875,N_10837);
nand U10999 (N_10999,N_10742,N_10741);
xnor U11000 (N_11000,N_10874,N_10870);
nor U11001 (N_11001,N_10855,N_10863);
and U11002 (N_11002,N_10720,N_10810);
and U11003 (N_11003,N_10766,N_10810);
or U11004 (N_11004,N_10850,N_10816);
nand U11005 (N_11005,N_10752,N_10801);
or U11006 (N_11006,N_10874,N_10795);
or U11007 (N_11007,N_10752,N_10831);
nand U11008 (N_11008,N_10826,N_10724);
or U11009 (N_11009,N_10777,N_10823);
or U11010 (N_11010,N_10746,N_10739);
and U11011 (N_11011,N_10801,N_10793);
and U11012 (N_11012,N_10877,N_10734);
nor U11013 (N_11013,N_10746,N_10735);
or U11014 (N_11014,N_10796,N_10840);
or U11015 (N_11015,N_10726,N_10750);
or U11016 (N_11016,N_10855,N_10732);
or U11017 (N_11017,N_10819,N_10744);
or U11018 (N_11018,N_10725,N_10769);
nand U11019 (N_11019,N_10783,N_10853);
xor U11020 (N_11020,N_10827,N_10789);
and U11021 (N_11021,N_10765,N_10858);
and U11022 (N_11022,N_10733,N_10791);
nand U11023 (N_11023,N_10786,N_10754);
or U11024 (N_11024,N_10749,N_10734);
or U11025 (N_11025,N_10751,N_10732);
nand U11026 (N_11026,N_10800,N_10802);
or U11027 (N_11027,N_10830,N_10724);
xor U11028 (N_11028,N_10872,N_10790);
nand U11029 (N_11029,N_10730,N_10871);
xnor U11030 (N_11030,N_10742,N_10788);
xnor U11031 (N_11031,N_10765,N_10863);
or U11032 (N_11032,N_10821,N_10837);
or U11033 (N_11033,N_10744,N_10765);
nor U11034 (N_11034,N_10822,N_10854);
nor U11035 (N_11035,N_10797,N_10838);
nor U11036 (N_11036,N_10870,N_10768);
and U11037 (N_11037,N_10828,N_10844);
and U11038 (N_11038,N_10768,N_10744);
and U11039 (N_11039,N_10806,N_10856);
nor U11040 (N_11040,N_10884,N_10983);
nand U11041 (N_11041,N_10978,N_10968);
nor U11042 (N_11042,N_10885,N_10981);
nor U11043 (N_11043,N_10922,N_10902);
or U11044 (N_11044,N_10934,N_10886);
or U11045 (N_11045,N_10958,N_10985);
or U11046 (N_11046,N_10921,N_10960);
or U11047 (N_11047,N_10991,N_10986);
xor U11048 (N_11048,N_11000,N_11021);
nand U11049 (N_11049,N_11013,N_11014);
xor U11050 (N_11050,N_10989,N_10982);
nand U11051 (N_11051,N_11018,N_10923);
xor U11052 (N_11052,N_10955,N_10995);
and U11053 (N_11053,N_11011,N_10904);
xnor U11054 (N_11054,N_10928,N_10945);
or U11055 (N_11055,N_10905,N_11010);
and U11056 (N_11056,N_10964,N_10994);
xnor U11057 (N_11057,N_10984,N_10999);
nand U11058 (N_11058,N_10912,N_10919);
or U11059 (N_11059,N_11037,N_11001);
nand U11060 (N_11060,N_10942,N_10990);
nor U11061 (N_11061,N_11035,N_11022);
nand U11062 (N_11062,N_10962,N_10938);
or U11063 (N_11063,N_10887,N_11023);
nand U11064 (N_11064,N_10965,N_10917);
xor U11065 (N_11065,N_10931,N_10979);
and U11066 (N_11066,N_11008,N_11002);
nand U11067 (N_11067,N_10889,N_11024);
and U11068 (N_11068,N_10897,N_11004);
nor U11069 (N_11069,N_10988,N_10880);
and U11070 (N_11070,N_10948,N_10924);
xor U11071 (N_11071,N_11030,N_11029);
nand U11072 (N_11072,N_10973,N_10943);
nand U11073 (N_11073,N_11016,N_10947);
xnor U11074 (N_11074,N_10959,N_10957);
and U11075 (N_11075,N_10935,N_10883);
nor U11076 (N_11076,N_10895,N_11015);
xnor U11077 (N_11077,N_10910,N_10888);
and U11078 (N_11078,N_10891,N_10894);
nand U11079 (N_11079,N_10929,N_10956);
or U11080 (N_11080,N_10970,N_10882);
nand U11081 (N_11081,N_10941,N_10974);
or U11082 (N_11082,N_10907,N_10940);
or U11083 (N_11083,N_11020,N_10903);
nor U11084 (N_11084,N_10915,N_10899);
nand U11085 (N_11085,N_10952,N_10949);
xor U11086 (N_11086,N_10998,N_10930);
xor U11087 (N_11087,N_10881,N_10892);
xnor U11088 (N_11088,N_10971,N_10993);
and U11089 (N_11089,N_11032,N_11028);
xnor U11090 (N_11090,N_11005,N_10961);
nand U11091 (N_11091,N_11038,N_10918);
or U11092 (N_11092,N_10963,N_10950);
or U11093 (N_11093,N_11012,N_11031);
nor U11094 (N_11094,N_10939,N_11033);
or U11095 (N_11095,N_10890,N_11039);
nand U11096 (N_11096,N_10975,N_11017);
nor U11097 (N_11097,N_10932,N_10954);
and U11098 (N_11098,N_10927,N_10937);
nand U11099 (N_11099,N_10936,N_10911);
nand U11100 (N_11100,N_11019,N_11003);
nand U11101 (N_11101,N_10976,N_10913);
nand U11102 (N_11102,N_10992,N_11025);
xnor U11103 (N_11103,N_10987,N_10896);
or U11104 (N_11104,N_10951,N_11007);
and U11105 (N_11105,N_10925,N_10900);
nor U11106 (N_11106,N_10906,N_11006);
nor U11107 (N_11107,N_10901,N_10916);
nand U11108 (N_11108,N_10969,N_10914);
or U11109 (N_11109,N_10967,N_10972);
or U11110 (N_11110,N_11036,N_10980);
nand U11111 (N_11111,N_10933,N_10898);
nand U11112 (N_11112,N_10997,N_11009);
or U11113 (N_11113,N_11027,N_10953);
or U11114 (N_11114,N_11026,N_11034);
xnor U11115 (N_11115,N_10946,N_10966);
nand U11116 (N_11116,N_10944,N_10893);
or U11117 (N_11117,N_10977,N_10908);
nor U11118 (N_11118,N_10996,N_10909);
and U11119 (N_11119,N_10926,N_10920);
or U11120 (N_11120,N_10915,N_10945);
or U11121 (N_11121,N_10961,N_10992);
xnor U11122 (N_11122,N_10965,N_10963);
nor U11123 (N_11123,N_10984,N_10887);
xnor U11124 (N_11124,N_10928,N_10930);
or U11125 (N_11125,N_10998,N_10925);
nor U11126 (N_11126,N_11001,N_10886);
and U11127 (N_11127,N_11039,N_11010);
or U11128 (N_11128,N_11031,N_11004);
nand U11129 (N_11129,N_11003,N_10967);
and U11130 (N_11130,N_11013,N_10903);
nand U11131 (N_11131,N_10936,N_11007);
or U11132 (N_11132,N_10944,N_10966);
nor U11133 (N_11133,N_11038,N_10999);
nor U11134 (N_11134,N_10932,N_10880);
nor U11135 (N_11135,N_10996,N_10965);
nor U11136 (N_11136,N_10882,N_11000);
nand U11137 (N_11137,N_10882,N_10886);
nor U11138 (N_11138,N_10941,N_10964);
nand U11139 (N_11139,N_11013,N_10934);
xor U11140 (N_11140,N_10929,N_10992);
or U11141 (N_11141,N_10964,N_10969);
nand U11142 (N_11142,N_10973,N_10923);
nand U11143 (N_11143,N_10893,N_10985);
and U11144 (N_11144,N_10918,N_10961);
and U11145 (N_11145,N_10914,N_11010);
nor U11146 (N_11146,N_11025,N_11012);
nand U11147 (N_11147,N_11010,N_11012);
or U11148 (N_11148,N_11035,N_10991);
or U11149 (N_11149,N_10881,N_10941);
or U11150 (N_11150,N_10894,N_10969);
nor U11151 (N_11151,N_10934,N_10975);
xor U11152 (N_11152,N_10903,N_10977);
nor U11153 (N_11153,N_10937,N_11005);
and U11154 (N_11154,N_10886,N_10950);
xnor U11155 (N_11155,N_11015,N_10986);
and U11156 (N_11156,N_10928,N_10907);
nand U11157 (N_11157,N_10967,N_10995);
nor U11158 (N_11158,N_10958,N_10987);
nand U11159 (N_11159,N_11018,N_10914);
xor U11160 (N_11160,N_10989,N_11023);
and U11161 (N_11161,N_11011,N_10896);
nor U11162 (N_11162,N_11027,N_11013);
and U11163 (N_11163,N_10956,N_11036);
and U11164 (N_11164,N_10911,N_10951);
nor U11165 (N_11165,N_10932,N_10983);
and U11166 (N_11166,N_10983,N_10963);
or U11167 (N_11167,N_10934,N_10970);
xor U11168 (N_11168,N_10952,N_10983);
or U11169 (N_11169,N_10967,N_11033);
nand U11170 (N_11170,N_10905,N_10981);
nor U11171 (N_11171,N_10958,N_10996);
nand U11172 (N_11172,N_11015,N_10926);
nand U11173 (N_11173,N_10908,N_10897);
or U11174 (N_11174,N_10929,N_10907);
xnor U11175 (N_11175,N_10884,N_10896);
xnor U11176 (N_11176,N_10967,N_10954);
xor U11177 (N_11177,N_11039,N_10981);
nor U11178 (N_11178,N_10902,N_11015);
and U11179 (N_11179,N_11004,N_10988);
xnor U11180 (N_11180,N_10937,N_10895);
xnor U11181 (N_11181,N_11028,N_10981);
xnor U11182 (N_11182,N_10975,N_10901);
xnor U11183 (N_11183,N_10898,N_10891);
nor U11184 (N_11184,N_10964,N_10896);
or U11185 (N_11185,N_10957,N_10972);
and U11186 (N_11186,N_10995,N_10974);
nor U11187 (N_11187,N_10961,N_10958);
nand U11188 (N_11188,N_11002,N_10908);
xor U11189 (N_11189,N_10888,N_10953);
and U11190 (N_11190,N_10923,N_11029);
or U11191 (N_11191,N_10955,N_10947);
xor U11192 (N_11192,N_11010,N_10880);
and U11193 (N_11193,N_10896,N_10952);
nand U11194 (N_11194,N_10925,N_10890);
nand U11195 (N_11195,N_11029,N_10932);
xnor U11196 (N_11196,N_10941,N_10992);
nor U11197 (N_11197,N_10944,N_10965);
and U11198 (N_11198,N_10920,N_10968);
or U11199 (N_11199,N_10928,N_10949);
and U11200 (N_11200,N_11051,N_11123);
nor U11201 (N_11201,N_11093,N_11199);
and U11202 (N_11202,N_11057,N_11109);
xnor U11203 (N_11203,N_11130,N_11137);
nand U11204 (N_11204,N_11079,N_11141);
nor U11205 (N_11205,N_11082,N_11155);
nand U11206 (N_11206,N_11177,N_11118);
nand U11207 (N_11207,N_11107,N_11135);
or U11208 (N_11208,N_11142,N_11108);
and U11209 (N_11209,N_11162,N_11043);
nor U11210 (N_11210,N_11105,N_11112);
and U11211 (N_11211,N_11170,N_11185);
nand U11212 (N_11212,N_11047,N_11129);
or U11213 (N_11213,N_11096,N_11140);
nor U11214 (N_11214,N_11110,N_11102);
xnor U11215 (N_11215,N_11103,N_11064);
or U11216 (N_11216,N_11078,N_11157);
nor U11217 (N_11217,N_11117,N_11106);
or U11218 (N_11218,N_11153,N_11191);
nor U11219 (N_11219,N_11190,N_11067);
nand U11220 (N_11220,N_11158,N_11086);
nand U11221 (N_11221,N_11041,N_11136);
and U11222 (N_11222,N_11074,N_11161);
nor U11223 (N_11223,N_11083,N_11111);
xor U11224 (N_11224,N_11100,N_11149);
or U11225 (N_11225,N_11042,N_11168);
nand U11226 (N_11226,N_11148,N_11147);
xnor U11227 (N_11227,N_11048,N_11165);
xor U11228 (N_11228,N_11186,N_11189);
nand U11229 (N_11229,N_11144,N_11193);
xnor U11230 (N_11230,N_11160,N_11120);
and U11231 (N_11231,N_11198,N_11113);
xor U11232 (N_11232,N_11151,N_11089);
nand U11233 (N_11233,N_11055,N_11115);
xnor U11234 (N_11234,N_11090,N_11114);
xnor U11235 (N_11235,N_11045,N_11194);
or U11236 (N_11236,N_11174,N_11104);
or U11237 (N_11237,N_11094,N_11119);
nand U11238 (N_11238,N_11126,N_11134);
nor U11239 (N_11239,N_11087,N_11182);
nor U11240 (N_11240,N_11180,N_11085);
nor U11241 (N_11241,N_11128,N_11184);
or U11242 (N_11242,N_11088,N_11062);
xnor U11243 (N_11243,N_11163,N_11124);
nand U11244 (N_11244,N_11122,N_11150);
and U11245 (N_11245,N_11116,N_11154);
nor U11246 (N_11246,N_11063,N_11197);
or U11247 (N_11247,N_11125,N_11044);
xor U11248 (N_11248,N_11179,N_11080);
xor U11249 (N_11249,N_11059,N_11066);
or U11250 (N_11250,N_11076,N_11138);
nand U11251 (N_11251,N_11098,N_11099);
or U11252 (N_11252,N_11178,N_11071);
and U11253 (N_11253,N_11054,N_11173);
nor U11254 (N_11254,N_11183,N_11046);
nand U11255 (N_11255,N_11187,N_11169);
and U11256 (N_11256,N_11145,N_11061);
and U11257 (N_11257,N_11056,N_11065);
xnor U11258 (N_11258,N_11188,N_11121);
nand U11259 (N_11259,N_11084,N_11049);
nand U11260 (N_11260,N_11133,N_11127);
xnor U11261 (N_11261,N_11068,N_11091);
or U11262 (N_11262,N_11101,N_11181);
or U11263 (N_11263,N_11139,N_11073);
and U11264 (N_11264,N_11081,N_11072);
nor U11265 (N_11265,N_11075,N_11156);
nand U11266 (N_11266,N_11196,N_11171);
nor U11267 (N_11267,N_11131,N_11097);
or U11268 (N_11268,N_11164,N_11167);
or U11269 (N_11269,N_11195,N_11095);
or U11270 (N_11270,N_11143,N_11053);
nor U11271 (N_11271,N_11159,N_11192);
xnor U11272 (N_11272,N_11060,N_11050);
or U11273 (N_11273,N_11152,N_11040);
nor U11274 (N_11274,N_11092,N_11058);
nand U11275 (N_11275,N_11077,N_11176);
xor U11276 (N_11276,N_11070,N_11175);
xnor U11277 (N_11277,N_11172,N_11166);
or U11278 (N_11278,N_11146,N_11069);
and U11279 (N_11279,N_11132,N_11052);
or U11280 (N_11280,N_11132,N_11107);
nor U11281 (N_11281,N_11130,N_11133);
nor U11282 (N_11282,N_11162,N_11063);
nor U11283 (N_11283,N_11172,N_11138);
or U11284 (N_11284,N_11043,N_11065);
xor U11285 (N_11285,N_11193,N_11164);
nor U11286 (N_11286,N_11166,N_11073);
or U11287 (N_11287,N_11064,N_11076);
nor U11288 (N_11288,N_11144,N_11078);
nand U11289 (N_11289,N_11115,N_11197);
nand U11290 (N_11290,N_11098,N_11122);
nand U11291 (N_11291,N_11197,N_11059);
and U11292 (N_11292,N_11058,N_11193);
xnor U11293 (N_11293,N_11181,N_11084);
nor U11294 (N_11294,N_11100,N_11140);
nand U11295 (N_11295,N_11181,N_11093);
nand U11296 (N_11296,N_11171,N_11132);
xnor U11297 (N_11297,N_11077,N_11109);
and U11298 (N_11298,N_11152,N_11079);
and U11299 (N_11299,N_11152,N_11126);
xnor U11300 (N_11300,N_11150,N_11177);
or U11301 (N_11301,N_11199,N_11054);
and U11302 (N_11302,N_11131,N_11149);
nor U11303 (N_11303,N_11115,N_11152);
xnor U11304 (N_11304,N_11086,N_11063);
or U11305 (N_11305,N_11108,N_11084);
nand U11306 (N_11306,N_11189,N_11051);
xor U11307 (N_11307,N_11060,N_11121);
nand U11308 (N_11308,N_11050,N_11185);
xnor U11309 (N_11309,N_11152,N_11100);
and U11310 (N_11310,N_11144,N_11098);
xnor U11311 (N_11311,N_11169,N_11175);
and U11312 (N_11312,N_11133,N_11166);
xnor U11313 (N_11313,N_11181,N_11136);
nand U11314 (N_11314,N_11183,N_11165);
or U11315 (N_11315,N_11157,N_11133);
xor U11316 (N_11316,N_11127,N_11196);
nor U11317 (N_11317,N_11174,N_11184);
or U11318 (N_11318,N_11139,N_11093);
xnor U11319 (N_11319,N_11078,N_11141);
and U11320 (N_11320,N_11045,N_11116);
xnor U11321 (N_11321,N_11068,N_11126);
and U11322 (N_11322,N_11124,N_11194);
or U11323 (N_11323,N_11155,N_11192);
nand U11324 (N_11324,N_11124,N_11056);
and U11325 (N_11325,N_11155,N_11146);
or U11326 (N_11326,N_11124,N_11050);
or U11327 (N_11327,N_11172,N_11088);
nand U11328 (N_11328,N_11174,N_11198);
nor U11329 (N_11329,N_11044,N_11062);
or U11330 (N_11330,N_11064,N_11087);
nor U11331 (N_11331,N_11115,N_11187);
and U11332 (N_11332,N_11105,N_11185);
nand U11333 (N_11333,N_11176,N_11130);
or U11334 (N_11334,N_11112,N_11077);
or U11335 (N_11335,N_11153,N_11166);
nor U11336 (N_11336,N_11196,N_11143);
nand U11337 (N_11337,N_11169,N_11096);
xnor U11338 (N_11338,N_11075,N_11184);
nor U11339 (N_11339,N_11150,N_11160);
nor U11340 (N_11340,N_11101,N_11057);
nand U11341 (N_11341,N_11154,N_11153);
or U11342 (N_11342,N_11170,N_11166);
nand U11343 (N_11343,N_11074,N_11110);
and U11344 (N_11344,N_11196,N_11062);
xor U11345 (N_11345,N_11165,N_11147);
nor U11346 (N_11346,N_11050,N_11187);
nand U11347 (N_11347,N_11130,N_11179);
nand U11348 (N_11348,N_11057,N_11140);
nor U11349 (N_11349,N_11059,N_11076);
nand U11350 (N_11350,N_11194,N_11163);
or U11351 (N_11351,N_11119,N_11185);
and U11352 (N_11352,N_11067,N_11117);
and U11353 (N_11353,N_11199,N_11185);
nor U11354 (N_11354,N_11096,N_11108);
xnor U11355 (N_11355,N_11065,N_11108);
and U11356 (N_11356,N_11160,N_11125);
nor U11357 (N_11357,N_11087,N_11195);
nor U11358 (N_11358,N_11145,N_11054);
xnor U11359 (N_11359,N_11107,N_11062);
nand U11360 (N_11360,N_11326,N_11335);
and U11361 (N_11361,N_11257,N_11304);
nor U11362 (N_11362,N_11353,N_11230);
nand U11363 (N_11363,N_11219,N_11275);
or U11364 (N_11364,N_11356,N_11350);
nor U11365 (N_11365,N_11303,N_11284);
and U11366 (N_11366,N_11292,N_11261);
nor U11367 (N_11367,N_11287,N_11319);
nor U11368 (N_11368,N_11323,N_11225);
nand U11369 (N_11369,N_11224,N_11270);
nor U11370 (N_11370,N_11213,N_11216);
and U11371 (N_11371,N_11315,N_11331);
and U11372 (N_11372,N_11204,N_11222);
and U11373 (N_11373,N_11263,N_11342);
xnor U11374 (N_11374,N_11211,N_11276);
and U11375 (N_11375,N_11321,N_11308);
xnor U11376 (N_11376,N_11264,N_11234);
and U11377 (N_11377,N_11316,N_11291);
nor U11378 (N_11378,N_11357,N_11343);
xor U11379 (N_11379,N_11217,N_11324);
or U11380 (N_11380,N_11289,N_11359);
or U11381 (N_11381,N_11294,N_11220);
and U11382 (N_11382,N_11346,N_11283);
nor U11383 (N_11383,N_11208,N_11277);
or U11384 (N_11384,N_11278,N_11355);
xor U11385 (N_11385,N_11351,N_11310);
nand U11386 (N_11386,N_11313,N_11336);
and U11387 (N_11387,N_11254,N_11273);
xnor U11388 (N_11388,N_11250,N_11228);
or U11389 (N_11389,N_11238,N_11320);
or U11390 (N_11390,N_11229,N_11341);
or U11391 (N_11391,N_11231,N_11332);
or U11392 (N_11392,N_11358,N_11285);
and U11393 (N_11393,N_11242,N_11296);
or U11394 (N_11394,N_11239,N_11271);
nor U11395 (N_11395,N_11297,N_11298);
or U11396 (N_11396,N_11295,N_11318);
nor U11397 (N_11397,N_11251,N_11243);
nand U11398 (N_11398,N_11258,N_11329);
nor U11399 (N_11399,N_11249,N_11256);
nand U11400 (N_11400,N_11209,N_11330);
or U11401 (N_11401,N_11237,N_11337);
and U11402 (N_11402,N_11334,N_11247);
and U11403 (N_11403,N_11223,N_11344);
and U11404 (N_11404,N_11322,N_11207);
xnor U11405 (N_11405,N_11299,N_11354);
or U11406 (N_11406,N_11248,N_11259);
nor U11407 (N_11407,N_11268,N_11267);
xnor U11408 (N_11408,N_11280,N_11290);
nand U11409 (N_11409,N_11236,N_11340);
nand U11410 (N_11410,N_11218,N_11317);
nand U11411 (N_11411,N_11245,N_11281);
or U11412 (N_11412,N_11327,N_11302);
and U11413 (N_11413,N_11311,N_11260);
nand U11414 (N_11414,N_11240,N_11253);
nor U11415 (N_11415,N_11325,N_11274);
nor U11416 (N_11416,N_11333,N_11201);
xor U11417 (N_11417,N_11255,N_11352);
nor U11418 (N_11418,N_11252,N_11203);
nand U11419 (N_11419,N_11266,N_11214);
xor U11420 (N_11420,N_11309,N_11246);
nand U11421 (N_11421,N_11221,N_11293);
and U11422 (N_11422,N_11200,N_11279);
nor U11423 (N_11423,N_11269,N_11210);
nand U11424 (N_11424,N_11286,N_11338);
nor U11425 (N_11425,N_11288,N_11262);
nand U11426 (N_11426,N_11244,N_11347);
and U11427 (N_11427,N_11272,N_11265);
and U11428 (N_11428,N_11282,N_11232);
xor U11429 (N_11429,N_11305,N_11233);
xnor U11430 (N_11430,N_11345,N_11348);
nand U11431 (N_11431,N_11235,N_11226);
or U11432 (N_11432,N_11300,N_11205);
nor U11433 (N_11433,N_11202,N_11215);
or U11434 (N_11434,N_11349,N_11206);
and U11435 (N_11435,N_11312,N_11301);
and U11436 (N_11436,N_11241,N_11339);
nand U11437 (N_11437,N_11328,N_11314);
and U11438 (N_11438,N_11307,N_11306);
nand U11439 (N_11439,N_11212,N_11227);
nor U11440 (N_11440,N_11205,N_11242);
and U11441 (N_11441,N_11313,N_11357);
nand U11442 (N_11442,N_11204,N_11215);
or U11443 (N_11443,N_11217,N_11300);
nand U11444 (N_11444,N_11359,N_11337);
or U11445 (N_11445,N_11217,N_11232);
xnor U11446 (N_11446,N_11289,N_11278);
xor U11447 (N_11447,N_11222,N_11322);
or U11448 (N_11448,N_11347,N_11227);
and U11449 (N_11449,N_11267,N_11354);
xor U11450 (N_11450,N_11246,N_11337);
xor U11451 (N_11451,N_11272,N_11336);
nor U11452 (N_11452,N_11339,N_11203);
nand U11453 (N_11453,N_11292,N_11232);
nor U11454 (N_11454,N_11229,N_11334);
or U11455 (N_11455,N_11278,N_11286);
nor U11456 (N_11456,N_11354,N_11278);
or U11457 (N_11457,N_11258,N_11298);
nand U11458 (N_11458,N_11276,N_11203);
nand U11459 (N_11459,N_11354,N_11276);
nor U11460 (N_11460,N_11337,N_11331);
nand U11461 (N_11461,N_11226,N_11330);
nor U11462 (N_11462,N_11283,N_11280);
and U11463 (N_11463,N_11335,N_11328);
nor U11464 (N_11464,N_11328,N_11333);
nor U11465 (N_11465,N_11240,N_11209);
or U11466 (N_11466,N_11275,N_11297);
or U11467 (N_11467,N_11226,N_11336);
and U11468 (N_11468,N_11309,N_11249);
nor U11469 (N_11469,N_11288,N_11204);
and U11470 (N_11470,N_11314,N_11271);
nand U11471 (N_11471,N_11355,N_11309);
or U11472 (N_11472,N_11222,N_11299);
nor U11473 (N_11473,N_11215,N_11298);
xnor U11474 (N_11474,N_11272,N_11259);
or U11475 (N_11475,N_11349,N_11275);
nor U11476 (N_11476,N_11323,N_11248);
or U11477 (N_11477,N_11289,N_11206);
xor U11478 (N_11478,N_11352,N_11356);
and U11479 (N_11479,N_11252,N_11231);
nor U11480 (N_11480,N_11272,N_11254);
xnor U11481 (N_11481,N_11243,N_11303);
xnor U11482 (N_11482,N_11217,N_11321);
xnor U11483 (N_11483,N_11240,N_11259);
xor U11484 (N_11484,N_11359,N_11306);
nand U11485 (N_11485,N_11289,N_11263);
and U11486 (N_11486,N_11212,N_11255);
nor U11487 (N_11487,N_11355,N_11319);
nand U11488 (N_11488,N_11292,N_11259);
and U11489 (N_11489,N_11333,N_11242);
nand U11490 (N_11490,N_11359,N_11240);
and U11491 (N_11491,N_11216,N_11279);
nor U11492 (N_11492,N_11224,N_11221);
or U11493 (N_11493,N_11302,N_11332);
and U11494 (N_11494,N_11201,N_11296);
nor U11495 (N_11495,N_11253,N_11300);
nand U11496 (N_11496,N_11296,N_11212);
xnor U11497 (N_11497,N_11327,N_11242);
and U11498 (N_11498,N_11223,N_11298);
nand U11499 (N_11499,N_11219,N_11203);
or U11500 (N_11500,N_11313,N_11265);
nand U11501 (N_11501,N_11261,N_11249);
xnor U11502 (N_11502,N_11273,N_11320);
or U11503 (N_11503,N_11344,N_11256);
or U11504 (N_11504,N_11266,N_11210);
nor U11505 (N_11505,N_11295,N_11245);
xor U11506 (N_11506,N_11238,N_11301);
and U11507 (N_11507,N_11317,N_11224);
nand U11508 (N_11508,N_11268,N_11265);
nor U11509 (N_11509,N_11281,N_11235);
and U11510 (N_11510,N_11356,N_11296);
and U11511 (N_11511,N_11245,N_11238);
nand U11512 (N_11512,N_11327,N_11204);
nand U11513 (N_11513,N_11211,N_11338);
and U11514 (N_11514,N_11201,N_11200);
or U11515 (N_11515,N_11304,N_11352);
nand U11516 (N_11516,N_11327,N_11211);
nand U11517 (N_11517,N_11201,N_11208);
or U11518 (N_11518,N_11269,N_11338);
xor U11519 (N_11519,N_11263,N_11324);
nor U11520 (N_11520,N_11409,N_11504);
nor U11521 (N_11521,N_11377,N_11420);
or U11522 (N_11522,N_11398,N_11369);
nor U11523 (N_11523,N_11513,N_11482);
and U11524 (N_11524,N_11440,N_11412);
or U11525 (N_11525,N_11402,N_11435);
nand U11526 (N_11526,N_11383,N_11399);
nand U11527 (N_11527,N_11418,N_11443);
nand U11528 (N_11528,N_11459,N_11458);
nand U11529 (N_11529,N_11462,N_11493);
xnor U11530 (N_11530,N_11421,N_11512);
nor U11531 (N_11531,N_11478,N_11410);
and U11532 (N_11532,N_11386,N_11423);
and U11533 (N_11533,N_11427,N_11479);
nor U11534 (N_11534,N_11509,N_11461);
xor U11535 (N_11535,N_11424,N_11428);
and U11536 (N_11536,N_11450,N_11411);
nand U11537 (N_11537,N_11474,N_11455);
and U11538 (N_11538,N_11470,N_11434);
and U11539 (N_11539,N_11491,N_11516);
and U11540 (N_11540,N_11372,N_11488);
xor U11541 (N_11541,N_11483,N_11413);
or U11542 (N_11542,N_11371,N_11497);
nand U11543 (N_11543,N_11449,N_11519);
or U11544 (N_11544,N_11368,N_11511);
or U11545 (N_11545,N_11490,N_11378);
or U11546 (N_11546,N_11406,N_11433);
nand U11547 (N_11547,N_11460,N_11375);
xnor U11548 (N_11548,N_11388,N_11376);
or U11549 (N_11549,N_11451,N_11415);
xnor U11550 (N_11550,N_11400,N_11405);
or U11551 (N_11551,N_11438,N_11494);
xnor U11552 (N_11552,N_11495,N_11487);
or U11553 (N_11553,N_11475,N_11496);
nor U11554 (N_11554,N_11446,N_11445);
and U11555 (N_11555,N_11444,N_11425);
or U11556 (N_11556,N_11441,N_11469);
nand U11557 (N_11557,N_11515,N_11390);
xnor U11558 (N_11558,N_11382,N_11505);
nor U11559 (N_11559,N_11394,N_11397);
nor U11560 (N_11560,N_11432,N_11426);
xnor U11561 (N_11561,N_11464,N_11456);
nor U11562 (N_11562,N_11499,N_11517);
nor U11563 (N_11563,N_11384,N_11506);
xnor U11564 (N_11564,N_11404,N_11485);
nand U11565 (N_11565,N_11465,N_11436);
nand U11566 (N_11566,N_11508,N_11477);
and U11567 (N_11567,N_11387,N_11489);
nand U11568 (N_11568,N_11492,N_11463);
xnor U11569 (N_11569,N_11395,N_11403);
nand U11570 (N_11570,N_11472,N_11501);
or U11571 (N_11571,N_11471,N_11365);
xnor U11572 (N_11572,N_11447,N_11498);
nor U11573 (N_11573,N_11468,N_11392);
xnor U11574 (N_11574,N_11518,N_11457);
or U11575 (N_11575,N_11453,N_11422);
or U11576 (N_11576,N_11467,N_11373);
or U11577 (N_11577,N_11416,N_11361);
nand U11578 (N_11578,N_11391,N_11385);
or U11579 (N_11579,N_11480,N_11380);
or U11580 (N_11580,N_11442,N_11437);
nand U11581 (N_11581,N_11510,N_11486);
or U11582 (N_11582,N_11454,N_11407);
or U11583 (N_11583,N_11503,N_11473);
nor U11584 (N_11584,N_11430,N_11419);
xnor U11585 (N_11585,N_11362,N_11431);
nand U11586 (N_11586,N_11393,N_11429);
or U11587 (N_11587,N_11374,N_11502);
or U11588 (N_11588,N_11360,N_11379);
nand U11589 (N_11589,N_11401,N_11366);
xor U11590 (N_11590,N_11466,N_11452);
nor U11591 (N_11591,N_11476,N_11484);
nand U11592 (N_11592,N_11414,N_11363);
or U11593 (N_11593,N_11481,N_11367);
xor U11594 (N_11594,N_11514,N_11500);
and U11595 (N_11595,N_11417,N_11381);
nor U11596 (N_11596,N_11408,N_11507);
nand U11597 (N_11597,N_11389,N_11364);
nor U11598 (N_11598,N_11370,N_11396);
nor U11599 (N_11599,N_11439,N_11448);
nor U11600 (N_11600,N_11469,N_11370);
xor U11601 (N_11601,N_11416,N_11406);
xnor U11602 (N_11602,N_11388,N_11480);
and U11603 (N_11603,N_11424,N_11408);
nand U11604 (N_11604,N_11429,N_11398);
and U11605 (N_11605,N_11411,N_11387);
nor U11606 (N_11606,N_11509,N_11391);
nand U11607 (N_11607,N_11486,N_11384);
nor U11608 (N_11608,N_11448,N_11487);
xnor U11609 (N_11609,N_11507,N_11468);
or U11610 (N_11610,N_11383,N_11444);
xor U11611 (N_11611,N_11374,N_11387);
or U11612 (N_11612,N_11512,N_11360);
and U11613 (N_11613,N_11437,N_11439);
and U11614 (N_11614,N_11482,N_11426);
and U11615 (N_11615,N_11430,N_11519);
and U11616 (N_11616,N_11451,N_11421);
or U11617 (N_11617,N_11436,N_11426);
or U11618 (N_11618,N_11510,N_11491);
nand U11619 (N_11619,N_11494,N_11413);
xnor U11620 (N_11620,N_11428,N_11410);
xor U11621 (N_11621,N_11460,N_11440);
xnor U11622 (N_11622,N_11490,N_11458);
xnor U11623 (N_11623,N_11450,N_11456);
nor U11624 (N_11624,N_11436,N_11471);
xor U11625 (N_11625,N_11510,N_11435);
nand U11626 (N_11626,N_11475,N_11375);
or U11627 (N_11627,N_11396,N_11406);
and U11628 (N_11628,N_11473,N_11388);
or U11629 (N_11629,N_11515,N_11422);
or U11630 (N_11630,N_11452,N_11474);
or U11631 (N_11631,N_11495,N_11424);
and U11632 (N_11632,N_11460,N_11373);
nand U11633 (N_11633,N_11460,N_11448);
and U11634 (N_11634,N_11411,N_11507);
xor U11635 (N_11635,N_11446,N_11410);
xnor U11636 (N_11636,N_11367,N_11434);
and U11637 (N_11637,N_11383,N_11445);
xnor U11638 (N_11638,N_11469,N_11473);
nand U11639 (N_11639,N_11514,N_11391);
nand U11640 (N_11640,N_11407,N_11461);
nand U11641 (N_11641,N_11512,N_11488);
or U11642 (N_11642,N_11400,N_11395);
or U11643 (N_11643,N_11480,N_11441);
nor U11644 (N_11644,N_11484,N_11512);
nor U11645 (N_11645,N_11406,N_11448);
nor U11646 (N_11646,N_11515,N_11443);
nand U11647 (N_11647,N_11472,N_11374);
nand U11648 (N_11648,N_11412,N_11443);
nand U11649 (N_11649,N_11444,N_11386);
and U11650 (N_11650,N_11406,N_11397);
nand U11651 (N_11651,N_11412,N_11397);
or U11652 (N_11652,N_11399,N_11374);
or U11653 (N_11653,N_11403,N_11452);
or U11654 (N_11654,N_11446,N_11501);
and U11655 (N_11655,N_11519,N_11417);
or U11656 (N_11656,N_11400,N_11459);
and U11657 (N_11657,N_11381,N_11373);
or U11658 (N_11658,N_11428,N_11435);
nor U11659 (N_11659,N_11426,N_11510);
nand U11660 (N_11660,N_11471,N_11367);
or U11661 (N_11661,N_11419,N_11417);
and U11662 (N_11662,N_11518,N_11389);
nand U11663 (N_11663,N_11479,N_11476);
xnor U11664 (N_11664,N_11444,N_11469);
nand U11665 (N_11665,N_11494,N_11422);
or U11666 (N_11666,N_11456,N_11467);
nand U11667 (N_11667,N_11407,N_11419);
and U11668 (N_11668,N_11378,N_11454);
and U11669 (N_11669,N_11448,N_11378);
nand U11670 (N_11670,N_11485,N_11369);
xor U11671 (N_11671,N_11491,N_11428);
nand U11672 (N_11672,N_11395,N_11429);
and U11673 (N_11673,N_11365,N_11369);
and U11674 (N_11674,N_11461,N_11408);
or U11675 (N_11675,N_11435,N_11513);
nand U11676 (N_11676,N_11440,N_11382);
nor U11677 (N_11677,N_11366,N_11383);
nand U11678 (N_11678,N_11465,N_11489);
and U11679 (N_11679,N_11382,N_11472);
or U11680 (N_11680,N_11580,N_11612);
nor U11681 (N_11681,N_11639,N_11611);
nand U11682 (N_11682,N_11571,N_11617);
or U11683 (N_11683,N_11582,N_11663);
or U11684 (N_11684,N_11554,N_11665);
nand U11685 (N_11685,N_11672,N_11605);
or U11686 (N_11686,N_11583,N_11650);
and U11687 (N_11687,N_11579,N_11602);
nor U11688 (N_11688,N_11556,N_11574);
nand U11689 (N_11689,N_11531,N_11620);
and U11690 (N_11690,N_11645,N_11656);
or U11691 (N_11691,N_11649,N_11591);
and U11692 (N_11692,N_11641,N_11592);
or U11693 (N_11693,N_11593,N_11653);
nand U11694 (N_11694,N_11568,N_11588);
or U11695 (N_11695,N_11601,N_11630);
or U11696 (N_11696,N_11547,N_11659);
nand U11697 (N_11697,N_11589,N_11581);
and U11698 (N_11698,N_11638,N_11561);
nor U11699 (N_11699,N_11626,N_11600);
or U11700 (N_11700,N_11619,N_11569);
nor U11701 (N_11701,N_11530,N_11634);
nand U11702 (N_11702,N_11636,N_11655);
xor U11703 (N_11703,N_11584,N_11564);
nor U11704 (N_11704,N_11660,N_11545);
nor U11705 (N_11705,N_11558,N_11594);
or U11706 (N_11706,N_11538,N_11543);
xnor U11707 (N_11707,N_11657,N_11677);
nor U11708 (N_11708,N_11526,N_11628);
or U11709 (N_11709,N_11675,N_11640);
nor U11710 (N_11710,N_11540,N_11546);
nor U11711 (N_11711,N_11658,N_11666);
or U11712 (N_11712,N_11572,N_11557);
xnor U11713 (N_11713,N_11613,N_11559);
xnor U11714 (N_11714,N_11521,N_11604);
xnor U11715 (N_11715,N_11537,N_11533);
or U11716 (N_11716,N_11646,N_11549);
xor U11717 (N_11717,N_11644,N_11585);
and U11718 (N_11718,N_11586,N_11609);
xnor U11719 (N_11719,N_11671,N_11667);
and U11720 (N_11720,N_11577,N_11535);
or U11721 (N_11721,N_11673,N_11578);
xor U11722 (N_11722,N_11674,N_11614);
nand U11723 (N_11723,N_11542,N_11635);
xnor U11724 (N_11724,N_11532,N_11522);
or U11725 (N_11725,N_11670,N_11573);
nand U11726 (N_11726,N_11529,N_11520);
and U11727 (N_11727,N_11534,N_11527);
or U11728 (N_11728,N_11631,N_11590);
and U11729 (N_11729,N_11587,N_11544);
or U11730 (N_11730,N_11648,N_11679);
and U11731 (N_11731,N_11607,N_11622);
or U11732 (N_11732,N_11621,N_11555);
xor U11733 (N_11733,N_11623,N_11523);
xor U11734 (N_11734,N_11664,N_11565);
or U11735 (N_11735,N_11627,N_11551);
or U11736 (N_11736,N_11595,N_11678);
nand U11737 (N_11737,N_11548,N_11550);
nor U11738 (N_11738,N_11536,N_11651);
nand U11739 (N_11739,N_11570,N_11662);
xnor U11740 (N_11740,N_11629,N_11560);
nand U11741 (N_11741,N_11606,N_11576);
or U11742 (N_11742,N_11598,N_11539);
or U11743 (N_11743,N_11603,N_11524);
nor U11744 (N_11744,N_11633,N_11562);
xnor U11745 (N_11745,N_11552,N_11668);
nor U11746 (N_11746,N_11642,N_11669);
or U11747 (N_11747,N_11599,N_11610);
xor U11748 (N_11748,N_11615,N_11575);
xnor U11749 (N_11749,N_11624,N_11661);
nor U11750 (N_11750,N_11616,N_11618);
xor U11751 (N_11751,N_11643,N_11654);
nor U11752 (N_11752,N_11567,N_11553);
or U11753 (N_11753,N_11637,N_11676);
nand U11754 (N_11754,N_11608,N_11596);
nor U11755 (N_11755,N_11652,N_11632);
nand U11756 (N_11756,N_11563,N_11525);
and U11757 (N_11757,N_11625,N_11541);
and U11758 (N_11758,N_11566,N_11528);
and U11759 (N_11759,N_11647,N_11597);
nand U11760 (N_11760,N_11601,N_11675);
and U11761 (N_11761,N_11655,N_11561);
nand U11762 (N_11762,N_11586,N_11578);
nor U11763 (N_11763,N_11605,N_11606);
nand U11764 (N_11764,N_11556,N_11532);
nand U11765 (N_11765,N_11637,N_11601);
and U11766 (N_11766,N_11641,N_11620);
nand U11767 (N_11767,N_11597,N_11679);
xor U11768 (N_11768,N_11546,N_11603);
and U11769 (N_11769,N_11643,N_11583);
and U11770 (N_11770,N_11571,N_11542);
and U11771 (N_11771,N_11586,N_11615);
and U11772 (N_11772,N_11537,N_11564);
or U11773 (N_11773,N_11650,N_11672);
nor U11774 (N_11774,N_11523,N_11672);
nor U11775 (N_11775,N_11614,N_11532);
xor U11776 (N_11776,N_11621,N_11525);
xnor U11777 (N_11777,N_11587,N_11546);
nand U11778 (N_11778,N_11574,N_11603);
xnor U11779 (N_11779,N_11641,N_11569);
or U11780 (N_11780,N_11541,N_11653);
nor U11781 (N_11781,N_11594,N_11602);
nor U11782 (N_11782,N_11671,N_11618);
xor U11783 (N_11783,N_11570,N_11527);
xnor U11784 (N_11784,N_11555,N_11537);
xnor U11785 (N_11785,N_11597,N_11575);
or U11786 (N_11786,N_11675,N_11623);
and U11787 (N_11787,N_11608,N_11530);
xnor U11788 (N_11788,N_11584,N_11600);
nor U11789 (N_11789,N_11631,N_11651);
xor U11790 (N_11790,N_11563,N_11661);
nand U11791 (N_11791,N_11592,N_11591);
nand U11792 (N_11792,N_11541,N_11526);
or U11793 (N_11793,N_11571,N_11676);
xor U11794 (N_11794,N_11522,N_11597);
nor U11795 (N_11795,N_11662,N_11559);
xnor U11796 (N_11796,N_11581,N_11559);
nor U11797 (N_11797,N_11528,N_11542);
nor U11798 (N_11798,N_11653,N_11637);
or U11799 (N_11799,N_11591,N_11632);
or U11800 (N_11800,N_11558,N_11534);
nand U11801 (N_11801,N_11573,N_11582);
xnor U11802 (N_11802,N_11600,N_11676);
xor U11803 (N_11803,N_11672,N_11533);
xnor U11804 (N_11804,N_11565,N_11576);
xnor U11805 (N_11805,N_11654,N_11576);
and U11806 (N_11806,N_11602,N_11564);
nor U11807 (N_11807,N_11582,N_11631);
xnor U11808 (N_11808,N_11616,N_11570);
or U11809 (N_11809,N_11622,N_11605);
nand U11810 (N_11810,N_11580,N_11591);
nor U11811 (N_11811,N_11549,N_11634);
xnor U11812 (N_11812,N_11571,N_11536);
and U11813 (N_11813,N_11527,N_11649);
xnor U11814 (N_11814,N_11545,N_11576);
or U11815 (N_11815,N_11526,N_11575);
or U11816 (N_11816,N_11672,N_11618);
xnor U11817 (N_11817,N_11542,N_11543);
and U11818 (N_11818,N_11575,N_11577);
nand U11819 (N_11819,N_11572,N_11542);
and U11820 (N_11820,N_11545,N_11630);
nand U11821 (N_11821,N_11526,N_11664);
or U11822 (N_11822,N_11616,N_11602);
or U11823 (N_11823,N_11644,N_11631);
nor U11824 (N_11824,N_11560,N_11671);
nand U11825 (N_11825,N_11625,N_11665);
nand U11826 (N_11826,N_11520,N_11542);
nand U11827 (N_11827,N_11672,N_11626);
or U11828 (N_11828,N_11670,N_11651);
nand U11829 (N_11829,N_11561,N_11671);
and U11830 (N_11830,N_11649,N_11602);
or U11831 (N_11831,N_11601,N_11598);
nor U11832 (N_11832,N_11562,N_11638);
xor U11833 (N_11833,N_11578,N_11595);
xnor U11834 (N_11834,N_11666,N_11644);
nor U11835 (N_11835,N_11587,N_11674);
xor U11836 (N_11836,N_11575,N_11602);
or U11837 (N_11837,N_11562,N_11645);
and U11838 (N_11838,N_11658,N_11671);
xor U11839 (N_11839,N_11536,N_11580);
or U11840 (N_11840,N_11759,N_11731);
xnor U11841 (N_11841,N_11767,N_11774);
and U11842 (N_11842,N_11730,N_11755);
xor U11843 (N_11843,N_11709,N_11716);
nand U11844 (N_11844,N_11700,N_11816);
or U11845 (N_11845,N_11807,N_11782);
nand U11846 (N_11846,N_11682,N_11783);
or U11847 (N_11847,N_11787,N_11693);
xor U11848 (N_11848,N_11809,N_11743);
or U11849 (N_11849,N_11751,N_11690);
nand U11850 (N_11850,N_11778,N_11789);
and U11851 (N_11851,N_11711,N_11754);
xor U11852 (N_11852,N_11707,N_11775);
and U11853 (N_11853,N_11836,N_11696);
nand U11854 (N_11854,N_11806,N_11817);
and U11855 (N_11855,N_11833,N_11829);
and U11856 (N_11856,N_11802,N_11704);
and U11857 (N_11857,N_11748,N_11741);
and U11858 (N_11858,N_11719,N_11753);
nor U11859 (N_11859,N_11835,N_11760);
and U11860 (N_11860,N_11756,N_11819);
xor U11861 (N_11861,N_11712,N_11761);
or U11862 (N_11862,N_11788,N_11834);
nor U11863 (N_11863,N_11791,N_11808);
or U11864 (N_11864,N_11763,N_11769);
nor U11865 (N_11865,N_11824,N_11739);
and U11866 (N_11866,N_11683,N_11747);
xnor U11867 (N_11867,N_11686,N_11758);
or U11868 (N_11868,N_11785,N_11799);
nor U11869 (N_11869,N_11796,N_11745);
and U11870 (N_11870,N_11695,N_11685);
xnor U11871 (N_11871,N_11714,N_11681);
xnor U11872 (N_11872,N_11722,N_11689);
and U11873 (N_11873,N_11780,N_11740);
nor U11874 (N_11874,N_11815,N_11793);
and U11875 (N_11875,N_11801,N_11732);
and U11876 (N_11876,N_11684,N_11823);
nand U11877 (N_11877,N_11728,N_11698);
xor U11878 (N_11878,N_11713,N_11738);
and U11879 (N_11879,N_11691,N_11813);
nor U11880 (N_11880,N_11697,N_11757);
and U11881 (N_11881,N_11826,N_11830);
nand U11882 (N_11882,N_11720,N_11779);
or U11883 (N_11883,N_11770,N_11792);
nor U11884 (N_11884,N_11744,N_11699);
xnor U11885 (N_11885,N_11680,N_11717);
xnor U11886 (N_11886,N_11765,N_11705);
or U11887 (N_11887,N_11781,N_11721);
and U11888 (N_11888,N_11750,N_11790);
xor U11889 (N_11889,N_11771,N_11794);
or U11890 (N_11890,N_11687,N_11768);
nand U11891 (N_11891,N_11837,N_11703);
xor U11892 (N_11892,N_11715,N_11735);
xor U11893 (N_11893,N_11776,N_11827);
and U11894 (N_11894,N_11694,N_11798);
and U11895 (N_11895,N_11724,N_11828);
and U11896 (N_11896,N_11812,N_11692);
nand U11897 (N_11897,N_11688,N_11832);
or U11898 (N_11898,N_11737,N_11710);
nand U11899 (N_11899,N_11764,N_11701);
or U11900 (N_11900,N_11746,N_11718);
and U11901 (N_11901,N_11822,N_11838);
and U11902 (N_11902,N_11777,N_11742);
xnor U11903 (N_11903,N_11800,N_11733);
xnor U11904 (N_11904,N_11821,N_11725);
nand U11905 (N_11905,N_11805,N_11726);
xnor U11906 (N_11906,N_11749,N_11803);
xor U11907 (N_11907,N_11727,N_11752);
and U11908 (N_11908,N_11766,N_11708);
nand U11909 (N_11909,N_11797,N_11795);
or U11910 (N_11910,N_11786,N_11736);
xnor U11911 (N_11911,N_11773,N_11810);
xor U11912 (N_11912,N_11729,N_11839);
xor U11913 (N_11913,N_11723,N_11818);
nand U11914 (N_11914,N_11831,N_11811);
or U11915 (N_11915,N_11772,N_11734);
nor U11916 (N_11916,N_11702,N_11706);
and U11917 (N_11917,N_11825,N_11762);
xor U11918 (N_11918,N_11814,N_11820);
xnor U11919 (N_11919,N_11804,N_11784);
xor U11920 (N_11920,N_11827,N_11812);
xnor U11921 (N_11921,N_11786,N_11773);
xor U11922 (N_11922,N_11812,N_11697);
nand U11923 (N_11923,N_11731,N_11691);
nor U11924 (N_11924,N_11773,N_11777);
nor U11925 (N_11925,N_11771,N_11792);
and U11926 (N_11926,N_11692,N_11709);
nor U11927 (N_11927,N_11697,N_11833);
xor U11928 (N_11928,N_11760,N_11685);
or U11929 (N_11929,N_11733,N_11809);
xor U11930 (N_11930,N_11791,N_11788);
xor U11931 (N_11931,N_11700,N_11775);
and U11932 (N_11932,N_11814,N_11809);
or U11933 (N_11933,N_11731,N_11689);
xnor U11934 (N_11934,N_11776,N_11743);
and U11935 (N_11935,N_11737,N_11802);
or U11936 (N_11936,N_11698,N_11791);
nand U11937 (N_11937,N_11764,N_11697);
nor U11938 (N_11938,N_11756,N_11814);
nand U11939 (N_11939,N_11735,N_11796);
nor U11940 (N_11940,N_11719,N_11837);
nor U11941 (N_11941,N_11725,N_11804);
nand U11942 (N_11942,N_11759,N_11693);
xor U11943 (N_11943,N_11731,N_11739);
and U11944 (N_11944,N_11764,N_11716);
nand U11945 (N_11945,N_11756,N_11775);
or U11946 (N_11946,N_11714,N_11692);
xor U11947 (N_11947,N_11836,N_11831);
nor U11948 (N_11948,N_11724,N_11686);
and U11949 (N_11949,N_11734,N_11702);
nor U11950 (N_11950,N_11756,N_11734);
and U11951 (N_11951,N_11815,N_11762);
nor U11952 (N_11952,N_11774,N_11758);
nor U11953 (N_11953,N_11791,N_11776);
nor U11954 (N_11954,N_11725,N_11770);
nor U11955 (N_11955,N_11683,N_11725);
and U11956 (N_11956,N_11735,N_11758);
nand U11957 (N_11957,N_11759,N_11699);
nand U11958 (N_11958,N_11719,N_11811);
and U11959 (N_11959,N_11807,N_11768);
xor U11960 (N_11960,N_11682,N_11725);
nand U11961 (N_11961,N_11763,N_11767);
or U11962 (N_11962,N_11783,N_11774);
nor U11963 (N_11963,N_11827,N_11808);
nor U11964 (N_11964,N_11683,N_11753);
nand U11965 (N_11965,N_11769,N_11771);
and U11966 (N_11966,N_11784,N_11705);
nor U11967 (N_11967,N_11782,N_11754);
and U11968 (N_11968,N_11766,N_11717);
nand U11969 (N_11969,N_11716,N_11787);
xnor U11970 (N_11970,N_11792,N_11720);
nor U11971 (N_11971,N_11713,N_11757);
nand U11972 (N_11972,N_11697,N_11816);
or U11973 (N_11973,N_11732,N_11730);
nor U11974 (N_11974,N_11787,N_11734);
nor U11975 (N_11975,N_11707,N_11711);
nand U11976 (N_11976,N_11837,N_11806);
nand U11977 (N_11977,N_11802,N_11735);
or U11978 (N_11978,N_11750,N_11783);
or U11979 (N_11979,N_11798,N_11732);
nor U11980 (N_11980,N_11776,N_11810);
nand U11981 (N_11981,N_11830,N_11681);
or U11982 (N_11982,N_11693,N_11827);
nor U11983 (N_11983,N_11774,N_11685);
nand U11984 (N_11984,N_11723,N_11780);
or U11985 (N_11985,N_11815,N_11798);
nor U11986 (N_11986,N_11717,N_11760);
nand U11987 (N_11987,N_11754,N_11757);
nor U11988 (N_11988,N_11827,N_11769);
nor U11989 (N_11989,N_11725,N_11692);
xor U11990 (N_11990,N_11795,N_11828);
or U11991 (N_11991,N_11758,N_11719);
xnor U11992 (N_11992,N_11685,N_11740);
nor U11993 (N_11993,N_11710,N_11768);
nand U11994 (N_11994,N_11825,N_11703);
or U11995 (N_11995,N_11682,N_11825);
nand U11996 (N_11996,N_11762,N_11734);
or U11997 (N_11997,N_11724,N_11726);
nor U11998 (N_11998,N_11774,N_11732);
xor U11999 (N_11999,N_11719,N_11818);
nand U12000 (N_12000,N_11976,N_11861);
and U12001 (N_12001,N_11933,N_11917);
nand U12002 (N_12002,N_11845,N_11866);
nand U12003 (N_12003,N_11881,N_11977);
and U12004 (N_12004,N_11852,N_11944);
nand U12005 (N_12005,N_11997,N_11905);
xnor U12006 (N_12006,N_11900,N_11988);
xor U12007 (N_12007,N_11927,N_11970);
nand U12008 (N_12008,N_11986,N_11850);
nand U12009 (N_12009,N_11871,N_11969);
xnor U12010 (N_12010,N_11912,N_11968);
xor U12011 (N_12011,N_11963,N_11849);
and U12012 (N_12012,N_11909,N_11924);
and U12013 (N_12013,N_11932,N_11956);
or U12014 (N_12014,N_11840,N_11989);
xor U12015 (N_12015,N_11873,N_11978);
or U12016 (N_12016,N_11960,N_11860);
and U12017 (N_12017,N_11863,N_11844);
nand U12018 (N_12018,N_11938,N_11967);
or U12019 (N_12019,N_11858,N_11931);
or U12020 (N_12020,N_11884,N_11954);
xnor U12021 (N_12021,N_11923,N_11918);
nor U12022 (N_12022,N_11922,N_11846);
or U12023 (N_12023,N_11911,N_11972);
nor U12024 (N_12024,N_11957,N_11888);
and U12025 (N_12025,N_11958,N_11897);
or U12026 (N_12026,N_11843,N_11885);
nor U12027 (N_12027,N_11907,N_11984);
xor U12028 (N_12028,N_11889,N_11847);
and U12029 (N_12029,N_11991,N_11891);
nand U12030 (N_12030,N_11929,N_11877);
nor U12031 (N_12031,N_11937,N_11961);
nand U12032 (N_12032,N_11915,N_11955);
or U12033 (N_12033,N_11896,N_11874);
nand U12034 (N_12034,N_11872,N_11892);
and U12035 (N_12035,N_11865,N_11925);
nor U12036 (N_12036,N_11893,N_11980);
or U12037 (N_12037,N_11941,N_11910);
and U12038 (N_12038,N_11981,N_11913);
or U12039 (N_12039,N_11901,N_11982);
xor U12040 (N_12040,N_11953,N_11862);
nand U12041 (N_12041,N_11848,N_11882);
xnor U12042 (N_12042,N_11857,N_11996);
xnor U12043 (N_12043,N_11947,N_11921);
and U12044 (N_12044,N_11964,N_11951);
or U12045 (N_12045,N_11998,N_11959);
or U12046 (N_12046,N_11868,N_11945);
or U12047 (N_12047,N_11920,N_11990);
xor U12048 (N_12048,N_11864,N_11886);
or U12049 (N_12049,N_11887,N_11854);
xnor U12050 (N_12050,N_11946,N_11883);
nand U12051 (N_12051,N_11904,N_11876);
nand U12052 (N_12052,N_11973,N_11841);
or U12053 (N_12053,N_11995,N_11916);
or U12054 (N_12054,N_11939,N_11974);
and U12055 (N_12055,N_11935,N_11926);
xor U12056 (N_12056,N_11943,N_11919);
and U12057 (N_12057,N_11965,N_11908);
nand U12058 (N_12058,N_11870,N_11899);
nand U12059 (N_12059,N_11949,N_11879);
or U12060 (N_12060,N_11906,N_11928);
or U12061 (N_12061,N_11966,N_11993);
or U12062 (N_12062,N_11987,N_11869);
xor U12063 (N_12063,N_11895,N_11936);
nor U12064 (N_12064,N_11898,N_11950);
xor U12065 (N_12065,N_11930,N_11890);
nand U12066 (N_12066,N_11851,N_11855);
and U12067 (N_12067,N_11983,N_11856);
nand U12068 (N_12068,N_11859,N_11962);
nand U12069 (N_12069,N_11999,N_11975);
and U12070 (N_12070,N_11971,N_11842);
and U12071 (N_12071,N_11942,N_11934);
and U12072 (N_12072,N_11985,N_11880);
and U12073 (N_12073,N_11894,N_11853);
or U12074 (N_12074,N_11994,N_11914);
or U12075 (N_12075,N_11992,N_11878);
or U12076 (N_12076,N_11875,N_11948);
and U12077 (N_12077,N_11952,N_11867);
nor U12078 (N_12078,N_11902,N_11903);
xor U12079 (N_12079,N_11940,N_11979);
xor U12080 (N_12080,N_11842,N_11845);
or U12081 (N_12081,N_11894,N_11892);
nand U12082 (N_12082,N_11863,N_11843);
and U12083 (N_12083,N_11851,N_11843);
or U12084 (N_12084,N_11846,N_11898);
xor U12085 (N_12085,N_11893,N_11951);
xor U12086 (N_12086,N_11991,N_11847);
or U12087 (N_12087,N_11980,N_11979);
nor U12088 (N_12088,N_11954,N_11978);
xor U12089 (N_12089,N_11888,N_11850);
nor U12090 (N_12090,N_11969,N_11906);
xor U12091 (N_12091,N_11976,N_11897);
or U12092 (N_12092,N_11983,N_11853);
and U12093 (N_12093,N_11925,N_11893);
nor U12094 (N_12094,N_11883,N_11938);
nand U12095 (N_12095,N_11879,N_11970);
nand U12096 (N_12096,N_11873,N_11953);
nand U12097 (N_12097,N_11935,N_11855);
nand U12098 (N_12098,N_11945,N_11992);
xnor U12099 (N_12099,N_11881,N_11864);
and U12100 (N_12100,N_11932,N_11910);
nand U12101 (N_12101,N_11854,N_11892);
or U12102 (N_12102,N_11877,N_11875);
or U12103 (N_12103,N_11923,N_11989);
xnor U12104 (N_12104,N_11942,N_11915);
or U12105 (N_12105,N_11946,N_11931);
xor U12106 (N_12106,N_11847,N_11934);
xnor U12107 (N_12107,N_11862,N_11915);
nand U12108 (N_12108,N_11897,N_11987);
xnor U12109 (N_12109,N_11901,N_11978);
xnor U12110 (N_12110,N_11853,N_11844);
or U12111 (N_12111,N_11942,N_11950);
and U12112 (N_12112,N_11889,N_11964);
and U12113 (N_12113,N_11932,N_11853);
nor U12114 (N_12114,N_11938,N_11882);
and U12115 (N_12115,N_11979,N_11910);
and U12116 (N_12116,N_11938,N_11849);
or U12117 (N_12117,N_11866,N_11968);
xor U12118 (N_12118,N_11945,N_11865);
xnor U12119 (N_12119,N_11862,N_11887);
or U12120 (N_12120,N_11864,N_11925);
xor U12121 (N_12121,N_11919,N_11965);
nand U12122 (N_12122,N_11986,N_11849);
nor U12123 (N_12123,N_11977,N_11858);
nand U12124 (N_12124,N_11999,N_11955);
nor U12125 (N_12125,N_11908,N_11843);
nand U12126 (N_12126,N_11941,N_11878);
and U12127 (N_12127,N_11975,N_11942);
nor U12128 (N_12128,N_11886,N_11987);
nand U12129 (N_12129,N_11856,N_11959);
nor U12130 (N_12130,N_11899,N_11845);
xnor U12131 (N_12131,N_11944,N_11881);
or U12132 (N_12132,N_11920,N_11958);
nor U12133 (N_12133,N_11968,N_11898);
xnor U12134 (N_12134,N_11871,N_11865);
or U12135 (N_12135,N_11932,N_11901);
and U12136 (N_12136,N_11926,N_11969);
nand U12137 (N_12137,N_11974,N_11960);
or U12138 (N_12138,N_11965,N_11912);
or U12139 (N_12139,N_11933,N_11984);
nor U12140 (N_12140,N_11968,N_11981);
xnor U12141 (N_12141,N_11926,N_11963);
or U12142 (N_12142,N_11892,N_11880);
and U12143 (N_12143,N_11966,N_11858);
xor U12144 (N_12144,N_11851,N_11954);
xor U12145 (N_12145,N_11887,N_11926);
or U12146 (N_12146,N_11959,N_11905);
xnor U12147 (N_12147,N_11985,N_11942);
and U12148 (N_12148,N_11969,N_11927);
or U12149 (N_12149,N_11988,N_11868);
nand U12150 (N_12150,N_11896,N_11880);
xnor U12151 (N_12151,N_11878,N_11934);
and U12152 (N_12152,N_11967,N_11941);
nor U12153 (N_12153,N_11890,N_11996);
or U12154 (N_12154,N_11870,N_11906);
and U12155 (N_12155,N_11946,N_11901);
xnor U12156 (N_12156,N_11943,N_11991);
nor U12157 (N_12157,N_11899,N_11977);
xor U12158 (N_12158,N_11938,N_11945);
and U12159 (N_12159,N_11962,N_11904);
nand U12160 (N_12160,N_12071,N_12122);
nor U12161 (N_12161,N_12107,N_12018);
or U12162 (N_12162,N_12050,N_12114);
nor U12163 (N_12163,N_12126,N_12024);
nor U12164 (N_12164,N_12075,N_12115);
nand U12165 (N_12165,N_12076,N_12105);
or U12166 (N_12166,N_12031,N_12144);
nor U12167 (N_12167,N_12042,N_12027);
or U12168 (N_12168,N_12012,N_12070);
and U12169 (N_12169,N_12061,N_12044);
or U12170 (N_12170,N_12026,N_12096);
nor U12171 (N_12171,N_12055,N_12003);
xnor U12172 (N_12172,N_12052,N_12025);
or U12173 (N_12173,N_12056,N_12116);
nand U12174 (N_12174,N_12088,N_12047);
nor U12175 (N_12175,N_12008,N_12072);
or U12176 (N_12176,N_12128,N_12065);
and U12177 (N_12177,N_12035,N_12112);
nand U12178 (N_12178,N_12131,N_12033);
and U12179 (N_12179,N_12090,N_12133);
nand U12180 (N_12180,N_12023,N_12092);
nor U12181 (N_12181,N_12086,N_12017);
xnor U12182 (N_12182,N_12108,N_12078);
and U12183 (N_12183,N_12104,N_12073);
or U12184 (N_12184,N_12136,N_12053);
and U12185 (N_12185,N_12098,N_12153);
and U12186 (N_12186,N_12041,N_12094);
nand U12187 (N_12187,N_12099,N_12081);
nor U12188 (N_12188,N_12006,N_12000);
nand U12189 (N_12189,N_12020,N_12155);
nor U12190 (N_12190,N_12142,N_12002);
and U12191 (N_12191,N_12015,N_12054);
or U12192 (N_12192,N_12066,N_12151);
nor U12193 (N_12193,N_12080,N_12082);
and U12194 (N_12194,N_12074,N_12148);
and U12195 (N_12195,N_12064,N_12119);
and U12196 (N_12196,N_12117,N_12130);
nand U12197 (N_12197,N_12121,N_12147);
xnor U12198 (N_12198,N_12150,N_12045);
or U12199 (N_12199,N_12125,N_12134);
and U12200 (N_12200,N_12087,N_12143);
xnor U12201 (N_12201,N_12043,N_12158);
or U12202 (N_12202,N_12005,N_12118);
nor U12203 (N_12203,N_12091,N_12101);
nand U12204 (N_12204,N_12046,N_12062);
or U12205 (N_12205,N_12068,N_12010);
and U12206 (N_12206,N_12156,N_12049);
nor U12207 (N_12207,N_12100,N_12146);
nor U12208 (N_12208,N_12109,N_12069);
or U12209 (N_12209,N_12030,N_12097);
nand U12210 (N_12210,N_12021,N_12032);
and U12211 (N_12211,N_12028,N_12157);
and U12212 (N_12212,N_12132,N_12029);
nand U12213 (N_12213,N_12138,N_12120);
nand U12214 (N_12214,N_12083,N_12159);
nor U12215 (N_12215,N_12152,N_12129);
xor U12216 (N_12216,N_12051,N_12137);
nand U12217 (N_12217,N_12001,N_12111);
nand U12218 (N_12218,N_12141,N_12102);
or U12219 (N_12219,N_12014,N_12113);
nor U12220 (N_12220,N_12060,N_12110);
nor U12221 (N_12221,N_12127,N_12058);
nand U12222 (N_12222,N_12140,N_12079);
xor U12223 (N_12223,N_12039,N_12106);
and U12224 (N_12224,N_12034,N_12038);
or U12225 (N_12225,N_12059,N_12009);
xnor U12226 (N_12226,N_12011,N_12095);
xnor U12227 (N_12227,N_12077,N_12004);
nand U12228 (N_12228,N_12007,N_12135);
or U12229 (N_12229,N_12093,N_12123);
or U12230 (N_12230,N_12048,N_12013);
nand U12231 (N_12231,N_12139,N_12019);
and U12232 (N_12232,N_12124,N_12084);
nand U12233 (N_12233,N_12085,N_12037);
and U12234 (N_12234,N_12036,N_12016);
and U12235 (N_12235,N_12057,N_12103);
xor U12236 (N_12236,N_12067,N_12145);
and U12237 (N_12237,N_12063,N_12154);
nand U12238 (N_12238,N_12022,N_12089);
xor U12239 (N_12239,N_12149,N_12040);
xor U12240 (N_12240,N_12136,N_12111);
or U12241 (N_12241,N_12016,N_12039);
or U12242 (N_12242,N_12004,N_12045);
and U12243 (N_12243,N_12156,N_12080);
nand U12244 (N_12244,N_12084,N_12110);
or U12245 (N_12245,N_12061,N_12086);
and U12246 (N_12246,N_12082,N_12051);
xnor U12247 (N_12247,N_12043,N_12015);
xnor U12248 (N_12248,N_12124,N_12129);
xor U12249 (N_12249,N_12035,N_12029);
xnor U12250 (N_12250,N_12122,N_12027);
and U12251 (N_12251,N_12014,N_12143);
xnor U12252 (N_12252,N_12055,N_12113);
nor U12253 (N_12253,N_12059,N_12104);
and U12254 (N_12254,N_12014,N_12048);
nand U12255 (N_12255,N_12121,N_12135);
and U12256 (N_12256,N_12137,N_12044);
and U12257 (N_12257,N_12058,N_12100);
xnor U12258 (N_12258,N_12025,N_12001);
nand U12259 (N_12259,N_12102,N_12154);
or U12260 (N_12260,N_12094,N_12148);
and U12261 (N_12261,N_12005,N_12013);
nand U12262 (N_12262,N_12144,N_12063);
nor U12263 (N_12263,N_12013,N_12025);
nor U12264 (N_12264,N_12132,N_12014);
or U12265 (N_12265,N_12011,N_12063);
nor U12266 (N_12266,N_12030,N_12098);
and U12267 (N_12267,N_12153,N_12009);
nor U12268 (N_12268,N_12106,N_12003);
nand U12269 (N_12269,N_12054,N_12098);
and U12270 (N_12270,N_12098,N_12043);
nor U12271 (N_12271,N_12005,N_12113);
nand U12272 (N_12272,N_12010,N_12029);
nand U12273 (N_12273,N_12087,N_12005);
xor U12274 (N_12274,N_12148,N_12084);
xor U12275 (N_12275,N_12021,N_12069);
xnor U12276 (N_12276,N_12063,N_12085);
or U12277 (N_12277,N_12141,N_12032);
or U12278 (N_12278,N_12112,N_12076);
or U12279 (N_12279,N_12014,N_12064);
nand U12280 (N_12280,N_12016,N_12060);
and U12281 (N_12281,N_12027,N_12081);
or U12282 (N_12282,N_12019,N_12123);
and U12283 (N_12283,N_12134,N_12027);
nor U12284 (N_12284,N_12016,N_12067);
nor U12285 (N_12285,N_12020,N_12063);
and U12286 (N_12286,N_12068,N_12014);
or U12287 (N_12287,N_12113,N_12156);
nand U12288 (N_12288,N_12028,N_12146);
nor U12289 (N_12289,N_12090,N_12092);
xor U12290 (N_12290,N_12105,N_12057);
nor U12291 (N_12291,N_12002,N_12125);
and U12292 (N_12292,N_12061,N_12078);
xnor U12293 (N_12293,N_12062,N_12060);
nor U12294 (N_12294,N_12001,N_12116);
or U12295 (N_12295,N_12097,N_12085);
and U12296 (N_12296,N_12070,N_12058);
or U12297 (N_12297,N_12147,N_12097);
nand U12298 (N_12298,N_12086,N_12003);
nand U12299 (N_12299,N_12041,N_12053);
and U12300 (N_12300,N_12079,N_12097);
nand U12301 (N_12301,N_12056,N_12085);
or U12302 (N_12302,N_12082,N_12000);
nand U12303 (N_12303,N_12096,N_12072);
xnor U12304 (N_12304,N_12071,N_12152);
or U12305 (N_12305,N_12051,N_12001);
or U12306 (N_12306,N_12001,N_12149);
or U12307 (N_12307,N_12128,N_12141);
or U12308 (N_12308,N_12041,N_12042);
nor U12309 (N_12309,N_12052,N_12021);
or U12310 (N_12310,N_12052,N_12063);
nand U12311 (N_12311,N_12152,N_12068);
xnor U12312 (N_12312,N_12069,N_12022);
xnor U12313 (N_12313,N_12073,N_12128);
nor U12314 (N_12314,N_12053,N_12111);
or U12315 (N_12315,N_12010,N_12062);
nand U12316 (N_12316,N_12152,N_12141);
or U12317 (N_12317,N_12065,N_12038);
and U12318 (N_12318,N_12057,N_12124);
nor U12319 (N_12319,N_12037,N_12106);
xor U12320 (N_12320,N_12235,N_12173);
xor U12321 (N_12321,N_12264,N_12196);
xor U12322 (N_12322,N_12168,N_12177);
and U12323 (N_12323,N_12176,N_12259);
or U12324 (N_12324,N_12181,N_12306);
xor U12325 (N_12325,N_12216,N_12283);
nand U12326 (N_12326,N_12313,N_12255);
nand U12327 (N_12327,N_12269,N_12194);
nand U12328 (N_12328,N_12166,N_12172);
nor U12329 (N_12329,N_12284,N_12190);
or U12330 (N_12330,N_12220,N_12222);
nor U12331 (N_12331,N_12160,N_12184);
or U12332 (N_12332,N_12205,N_12265);
or U12333 (N_12333,N_12180,N_12239);
xor U12334 (N_12334,N_12273,N_12211);
and U12335 (N_12335,N_12206,N_12243);
and U12336 (N_12336,N_12192,N_12279);
nand U12337 (N_12337,N_12212,N_12203);
nor U12338 (N_12338,N_12161,N_12167);
xnor U12339 (N_12339,N_12241,N_12179);
or U12340 (N_12340,N_12233,N_12197);
xnor U12341 (N_12341,N_12318,N_12319);
and U12342 (N_12342,N_12217,N_12266);
nor U12343 (N_12343,N_12302,N_12164);
xor U12344 (N_12344,N_12275,N_12246);
and U12345 (N_12345,N_12207,N_12218);
or U12346 (N_12346,N_12200,N_12189);
and U12347 (N_12347,N_12186,N_12303);
xor U12348 (N_12348,N_12256,N_12247);
nand U12349 (N_12349,N_12226,N_12185);
nand U12350 (N_12350,N_12232,N_12209);
nand U12351 (N_12351,N_12162,N_12242);
xnor U12352 (N_12352,N_12278,N_12317);
nand U12353 (N_12353,N_12178,N_12261);
xor U12354 (N_12354,N_12253,N_12204);
nor U12355 (N_12355,N_12295,N_12225);
or U12356 (N_12356,N_12213,N_12298);
nor U12357 (N_12357,N_12231,N_12294);
and U12358 (N_12358,N_12237,N_12287);
nand U12359 (N_12359,N_12300,N_12245);
and U12360 (N_12360,N_12215,N_12268);
nor U12361 (N_12361,N_12260,N_12267);
nand U12362 (N_12362,N_12163,N_12195);
or U12363 (N_12363,N_12271,N_12276);
xor U12364 (N_12364,N_12236,N_12227);
and U12365 (N_12365,N_12296,N_12210);
nand U12366 (N_12366,N_12250,N_12169);
nand U12367 (N_12367,N_12219,N_12274);
nor U12368 (N_12368,N_12263,N_12285);
nor U12369 (N_12369,N_12175,N_12291);
nand U12370 (N_12370,N_12252,N_12208);
or U12371 (N_12371,N_12182,N_12170);
and U12372 (N_12372,N_12223,N_12249);
nor U12373 (N_12373,N_12228,N_12201);
xnor U12374 (N_12374,N_12314,N_12165);
or U12375 (N_12375,N_12299,N_12251);
nand U12376 (N_12376,N_12258,N_12280);
nand U12377 (N_12377,N_12198,N_12221);
xnor U12378 (N_12378,N_12309,N_12183);
xor U12379 (N_12379,N_12293,N_12277);
nor U12380 (N_12380,N_12240,N_12301);
nand U12381 (N_12381,N_12224,N_12282);
nor U12382 (N_12382,N_12290,N_12272);
nor U12383 (N_12383,N_12238,N_12292);
nor U12384 (N_12384,N_12297,N_12304);
or U12385 (N_12385,N_12188,N_12174);
nand U12386 (N_12386,N_12308,N_12254);
nor U12387 (N_12387,N_12262,N_12230);
or U12388 (N_12388,N_12234,N_12171);
xnor U12389 (N_12389,N_12310,N_12248);
nand U12390 (N_12390,N_12311,N_12286);
and U12391 (N_12391,N_12316,N_12289);
nand U12392 (N_12392,N_12288,N_12281);
nand U12393 (N_12393,N_12214,N_12199);
xor U12394 (N_12394,N_12315,N_12187);
or U12395 (N_12395,N_12307,N_12229);
xnor U12396 (N_12396,N_12305,N_12270);
or U12397 (N_12397,N_12257,N_12312);
xnor U12398 (N_12398,N_12244,N_12193);
xnor U12399 (N_12399,N_12191,N_12202);
nand U12400 (N_12400,N_12205,N_12314);
nand U12401 (N_12401,N_12220,N_12269);
xnor U12402 (N_12402,N_12190,N_12286);
or U12403 (N_12403,N_12271,N_12197);
xor U12404 (N_12404,N_12233,N_12234);
nand U12405 (N_12405,N_12316,N_12231);
and U12406 (N_12406,N_12272,N_12175);
and U12407 (N_12407,N_12214,N_12275);
xnor U12408 (N_12408,N_12281,N_12306);
nor U12409 (N_12409,N_12295,N_12278);
nand U12410 (N_12410,N_12284,N_12213);
nand U12411 (N_12411,N_12204,N_12276);
xnor U12412 (N_12412,N_12165,N_12265);
and U12413 (N_12413,N_12228,N_12227);
or U12414 (N_12414,N_12238,N_12185);
nor U12415 (N_12415,N_12231,N_12211);
nand U12416 (N_12416,N_12237,N_12296);
xor U12417 (N_12417,N_12214,N_12293);
nand U12418 (N_12418,N_12281,N_12177);
nand U12419 (N_12419,N_12272,N_12285);
or U12420 (N_12420,N_12285,N_12166);
nand U12421 (N_12421,N_12230,N_12304);
xor U12422 (N_12422,N_12230,N_12300);
nand U12423 (N_12423,N_12223,N_12230);
or U12424 (N_12424,N_12184,N_12244);
nor U12425 (N_12425,N_12294,N_12256);
and U12426 (N_12426,N_12189,N_12178);
nor U12427 (N_12427,N_12243,N_12217);
xor U12428 (N_12428,N_12223,N_12160);
and U12429 (N_12429,N_12240,N_12246);
or U12430 (N_12430,N_12310,N_12270);
or U12431 (N_12431,N_12198,N_12250);
xor U12432 (N_12432,N_12199,N_12300);
nand U12433 (N_12433,N_12270,N_12259);
nand U12434 (N_12434,N_12191,N_12286);
and U12435 (N_12435,N_12210,N_12228);
nor U12436 (N_12436,N_12298,N_12243);
nand U12437 (N_12437,N_12297,N_12232);
nand U12438 (N_12438,N_12295,N_12294);
nor U12439 (N_12439,N_12237,N_12223);
nand U12440 (N_12440,N_12164,N_12208);
xnor U12441 (N_12441,N_12293,N_12316);
nor U12442 (N_12442,N_12231,N_12160);
nand U12443 (N_12443,N_12310,N_12257);
xnor U12444 (N_12444,N_12207,N_12269);
or U12445 (N_12445,N_12176,N_12316);
nand U12446 (N_12446,N_12213,N_12266);
and U12447 (N_12447,N_12171,N_12222);
or U12448 (N_12448,N_12277,N_12230);
nand U12449 (N_12449,N_12240,N_12218);
or U12450 (N_12450,N_12239,N_12295);
or U12451 (N_12451,N_12160,N_12312);
or U12452 (N_12452,N_12290,N_12202);
xnor U12453 (N_12453,N_12294,N_12198);
xnor U12454 (N_12454,N_12223,N_12209);
xor U12455 (N_12455,N_12287,N_12218);
nor U12456 (N_12456,N_12292,N_12242);
or U12457 (N_12457,N_12262,N_12299);
or U12458 (N_12458,N_12286,N_12160);
or U12459 (N_12459,N_12200,N_12308);
xnor U12460 (N_12460,N_12274,N_12214);
or U12461 (N_12461,N_12295,N_12287);
nand U12462 (N_12462,N_12284,N_12250);
nand U12463 (N_12463,N_12209,N_12318);
and U12464 (N_12464,N_12184,N_12181);
xnor U12465 (N_12465,N_12173,N_12244);
and U12466 (N_12466,N_12160,N_12296);
nor U12467 (N_12467,N_12277,N_12268);
xnor U12468 (N_12468,N_12305,N_12250);
xnor U12469 (N_12469,N_12200,N_12312);
and U12470 (N_12470,N_12299,N_12235);
nand U12471 (N_12471,N_12178,N_12310);
xnor U12472 (N_12472,N_12304,N_12286);
and U12473 (N_12473,N_12161,N_12228);
xor U12474 (N_12474,N_12185,N_12174);
or U12475 (N_12475,N_12160,N_12261);
and U12476 (N_12476,N_12268,N_12275);
nand U12477 (N_12477,N_12272,N_12217);
or U12478 (N_12478,N_12284,N_12222);
and U12479 (N_12479,N_12263,N_12209);
and U12480 (N_12480,N_12456,N_12434);
xor U12481 (N_12481,N_12336,N_12357);
and U12482 (N_12482,N_12372,N_12477);
nor U12483 (N_12483,N_12447,N_12425);
or U12484 (N_12484,N_12444,N_12394);
nor U12485 (N_12485,N_12383,N_12362);
or U12486 (N_12486,N_12445,N_12432);
nor U12487 (N_12487,N_12375,N_12359);
or U12488 (N_12488,N_12399,N_12323);
or U12489 (N_12489,N_12395,N_12368);
nor U12490 (N_12490,N_12403,N_12431);
or U12491 (N_12491,N_12389,N_12404);
nor U12492 (N_12492,N_12380,N_12423);
nand U12493 (N_12493,N_12396,N_12386);
and U12494 (N_12494,N_12391,N_12424);
or U12495 (N_12495,N_12350,N_12417);
nand U12496 (N_12496,N_12390,N_12377);
nor U12497 (N_12497,N_12345,N_12439);
and U12498 (N_12498,N_12408,N_12349);
and U12499 (N_12499,N_12363,N_12428);
and U12500 (N_12500,N_12385,N_12388);
xor U12501 (N_12501,N_12321,N_12438);
xor U12502 (N_12502,N_12337,N_12450);
xor U12503 (N_12503,N_12329,N_12387);
xnor U12504 (N_12504,N_12406,N_12418);
nand U12505 (N_12505,N_12440,N_12476);
and U12506 (N_12506,N_12343,N_12448);
and U12507 (N_12507,N_12464,N_12411);
nand U12508 (N_12508,N_12352,N_12351);
and U12509 (N_12509,N_12460,N_12376);
or U12510 (N_12510,N_12401,N_12457);
xnor U12511 (N_12511,N_12346,N_12471);
nor U12512 (N_12512,N_12367,N_12382);
xor U12513 (N_12513,N_12466,N_12433);
and U12514 (N_12514,N_12416,N_12436);
xnor U12515 (N_12515,N_12435,N_12326);
or U12516 (N_12516,N_12333,N_12461);
xnor U12517 (N_12517,N_12437,N_12358);
xor U12518 (N_12518,N_12463,N_12458);
nand U12519 (N_12519,N_12342,N_12327);
nor U12520 (N_12520,N_12378,N_12322);
xnor U12521 (N_12521,N_12465,N_12452);
and U12522 (N_12522,N_12472,N_12470);
xor U12523 (N_12523,N_12338,N_12344);
or U12524 (N_12524,N_12402,N_12468);
or U12525 (N_12525,N_12422,N_12361);
or U12526 (N_12526,N_12479,N_12331);
or U12527 (N_12527,N_12414,N_12455);
or U12528 (N_12528,N_12334,N_12335);
or U12529 (N_12529,N_12409,N_12420);
or U12530 (N_12530,N_12446,N_12407);
nand U12531 (N_12531,N_12347,N_12443);
and U12532 (N_12532,N_12353,N_12429);
or U12533 (N_12533,N_12475,N_12328);
nor U12534 (N_12534,N_12366,N_12467);
xor U12535 (N_12535,N_12330,N_12426);
or U12536 (N_12536,N_12398,N_12413);
and U12537 (N_12537,N_12384,N_12451);
and U12538 (N_12538,N_12365,N_12324);
and U12539 (N_12539,N_12369,N_12325);
nand U12540 (N_12540,N_12462,N_12412);
and U12541 (N_12541,N_12354,N_12355);
and U12542 (N_12542,N_12360,N_12419);
nor U12543 (N_12543,N_12397,N_12400);
or U12544 (N_12544,N_12379,N_12421);
nand U12545 (N_12545,N_12381,N_12459);
nand U12546 (N_12546,N_12348,N_12339);
or U12547 (N_12547,N_12453,N_12478);
or U12548 (N_12548,N_12410,N_12370);
or U12549 (N_12549,N_12332,N_12341);
nand U12550 (N_12550,N_12454,N_12340);
nor U12551 (N_12551,N_12374,N_12405);
nor U12552 (N_12552,N_12430,N_12442);
or U12553 (N_12553,N_12356,N_12427);
or U12554 (N_12554,N_12371,N_12393);
nand U12555 (N_12555,N_12441,N_12449);
nand U12556 (N_12556,N_12474,N_12469);
xnor U12557 (N_12557,N_12392,N_12364);
nand U12558 (N_12558,N_12320,N_12373);
or U12559 (N_12559,N_12415,N_12473);
nor U12560 (N_12560,N_12370,N_12390);
nor U12561 (N_12561,N_12347,N_12346);
nand U12562 (N_12562,N_12349,N_12434);
nor U12563 (N_12563,N_12473,N_12466);
nand U12564 (N_12564,N_12352,N_12374);
nor U12565 (N_12565,N_12327,N_12362);
nor U12566 (N_12566,N_12444,N_12462);
xor U12567 (N_12567,N_12337,N_12455);
xor U12568 (N_12568,N_12412,N_12341);
or U12569 (N_12569,N_12330,N_12400);
or U12570 (N_12570,N_12421,N_12399);
or U12571 (N_12571,N_12424,N_12400);
and U12572 (N_12572,N_12407,N_12335);
and U12573 (N_12573,N_12459,N_12460);
nand U12574 (N_12574,N_12378,N_12476);
and U12575 (N_12575,N_12324,N_12402);
nor U12576 (N_12576,N_12324,N_12343);
nand U12577 (N_12577,N_12356,N_12349);
xor U12578 (N_12578,N_12376,N_12479);
xor U12579 (N_12579,N_12421,N_12326);
and U12580 (N_12580,N_12460,N_12345);
nand U12581 (N_12581,N_12478,N_12470);
nand U12582 (N_12582,N_12472,N_12327);
or U12583 (N_12583,N_12428,N_12444);
xor U12584 (N_12584,N_12408,N_12352);
xor U12585 (N_12585,N_12356,N_12475);
xnor U12586 (N_12586,N_12394,N_12465);
xnor U12587 (N_12587,N_12366,N_12454);
nand U12588 (N_12588,N_12362,N_12372);
nor U12589 (N_12589,N_12431,N_12413);
xnor U12590 (N_12590,N_12397,N_12391);
nor U12591 (N_12591,N_12354,N_12359);
xnor U12592 (N_12592,N_12345,N_12381);
nor U12593 (N_12593,N_12332,N_12462);
or U12594 (N_12594,N_12364,N_12445);
or U12595 (N_12595,N_12431,N_12367);
nand U12596 (N_12596,N_12362,N_12411);
nor U12597 (N_12597,N_12453,N_12461);
and U12598 (N_12598,N_12365,N_12351);
nand U12599 (N_12599,N_12464,N_12332);
nor U12600 (N_12600,N_12323,N_12394);
xor U12601 (N_12601,N_12403,N_12411);
nand U12602 (N_12602,N_12420,N_12399);
nor U12603 (N_12603,N_12387,N_12450);
xor U12604 (N_12604,N_12358,N_12320);
nor U12605 (N_12605,N_12428,N_12442);
nor U12606 (N_12606,N_12479,N_12337);
or U12607 (N_12607,N_12411,N_12428);
or U12608 (N_12608,N_12436,N_12407);
xnor U12609 (N_12609,N_12413,N_12416);
xnor U12610 (N_12610,N_12370,N_12424);
xnor U12611 (N_12611,N_12377,N_12412);
and U12612 (N_12612,N_12448,N_12324);
xor U12613 (N_12613,N_12377,N_12345);
or U12614 (N_12614,N_12379,N_12397);
xor U12615 (N_12615,N_12420,N_12472);
nand U12616 (N_12616,N_12409,N_12433);
xor U12617 (N_12617,N_12462,N_12432);
and U12618 (N_12618,N_12450,N_12384);
nand U12619 (N_12619,N_12406,N_12450);
xnor U12620 (N_12620,N_12436,N_12449);
xnor U12621 (N_12621,N_12353,N_12474);
nand U12622 (N_12622,N_12440,N_12402);
or U12623 (N_12623,N_12447,N_12476);
nor U12624 (N_12624,N_12322,N_12457);
nor U12625 (N_12625,N_12466,N_12382);
xor U12626 (N_12626,N_12351,N_12459);
xor U12627 (N_12627,N_12467,N_12416);
and U12628 (N_12628,N_12399,N_12367);
xor U12629 (N_12629,N_12415,N_12377);
or U12630 (N_12630,N_12449,N_12326);
nor U12631 (N_12631,N_12332,N_12351);
and U12632 (N_12632,N_12449,N_12465);
xor U12633 (N_12633,N_12400,N_12383);
xnor U12634 (N_12634,N_12379,N_12427);
xor U12635 (N_12635,N_12435,N_12363);
or U12636 (N_12636,N_12449,N_12478);
nor U12637 (N_12637,N_12401,N_12438);
or U12638 (N_12638,N_12434,N_12470);
and U12639 (N_12639,N_12389,N_12358);
nor U12640 (N_12640,N_12487,N_12544);
nand U12641 (N_12641,N_12537,N_12545);
nor U12642 (N_12642,N_12609,N_12638);
and U12643 (N_12643,N_12630,N_12504);
and U12644 (N_12644,N_12529,N_12636);
nand U12645 (N_12645,N_12540,N_12521);
or U12646 (N_12646,N_12485,N_12577);
nand U12647 (N_12647,N_12584,N_12551);
nor U12648 (N_12648,N_12536,N_12510);
nand U12649 (N_12649,N_12593,N_12542);
and U12650 (N_12650,N_12580,N_12603);
nor U12651 (N_12651,N_12586,N_12617);
and U12652 (N_12652,N_12483,N_12486);
nand U12653 (N_12653,N_12623,N_12557);
nor U12654 (N_12654,N_12602,N_12624);
xor U12655 (N_12655,N_12533,N_12618);
xnor U12656 (N_12656,N_12500,N_12491);
nand U12657 (N_12657,N_12563,N_12561);
and U12658 (N_12658,N_12524,N_12621);
xnor U12659 (N_12659,N_12488,N_12562);
or U12660 (N_12660,N_12581,N_12626);
nand U12661 (N_12661,N_12637,N_12568);
or U12662 (N_12662,N_12511,N_12614);
or U12663 (N_12663,N_12541,N_12523);
xnor U12664 (N_12664,N_12526,N_12525);
xor U12665 (N_12665,N_12556,N_12496);
or U12666 (N_12666,N_12559,N_12607);
nor U12667 (N_12667,N_12590,N_12600);
xnor U12668 (N_12668,N_12535,N_12605);
xor U12669 (N_12669,N_12480,N_12503);
nor U12670 (N_12670,N_12516,N_12578);
nand U12671 (N_12671,N_12506,N_12601);
nor U12672 (N_12672,N_12518,N_12589);
and U12673 (N_12673,N_12543,N_12595);
and U12674 (N_12674,N_12597,N_12604);
and U12675 (N_12675,N_12547,N_12515);
xnor U12676 (N_12676,N_12552,N_12616);
or U12677 (N_12677,N_12598,N_12558);
nand U12678 (N_12678,N_12615,N_12507);
and U12679 (N_12679,N_12513,N_12564);
or U12680 (N_12680,N_12481,N_12548);
xor U12681 (N_12681,N_12583,N_12530);
or U12682 (N_12682,N_12489,N_12494);
nand U12683 (N_12683,N_12613,N_12512);
nor U12684 (N_12684,N_12592,N_12569);
and U12685 (N_12685,N_12587,N_12499);
nor U12686 (N_12686,N_12629,N_12572);
nor U12687 (N_12687,N_12639,N_12554);
nand U12688 (N_12688,N_12576,N_12575);
and U12689 (N_12689,N_12534,N_12608);
nand U12690 (N_12690,N_12522,N_12514);
or U12691 (N_12691,N_12582,N_12571);
or U12692 (N_12692,N_12591,N_12495);
nand U12693 (N_12693,N_12555,N_12631);
and U12694 (N_12694,N_12625,N_12532);
xnor U12695 (N_12695,N_12492,N_12538);
xnor U12696 (N_12696,N_12505,N_12508);
nor U12697 (N_12697,N_12531,N_12633);
nand U12698 (N_12698,N_12549,N_12627);
and U12699 (N_12699,N_12634,N_12573);
or U12700 (N_12700,N_12611,N_12596);
and U12701 (N_12701,N_12553,N_12622);
xor U12702 (N_12702,N_12493,N_12567);
and U12703 (N_12703,N_12484,N_12546);
nor U12704 (N_12704,N_12490,N_12612);
or U12705 (N_12705,N_12519,N_12497);
nand U12706 (N_12706,N_12501,N_12635);
nand U12707 (N_12707,N_12574,N_12620);
nor U12708 (N_12708,N_12528,N_12482);
nor U12709 (N_12709,N_12585,N_12619);
or U12710 (N_12710,N_12610,N_12527);
and U12711 (N_12711,N_12570,N_12599);
nand U12712 (N_12712,N_12628,N_12517);
nand U12713 (N_12713,N_12566,N_12498);
nand U12714 (N_12714,N_12606,N_12632);
nor U12715 (N_12715,N_12565,N_12539);
and U12716 (N_12716,N_12588,N_12594);
nor U12717 (N_12717,N_12550,N_12502);
nor U12718 (N_12718,N_12520,N_12560);
xor U12719 (N_12719,N_12509,N_12579);
nand U12720 (N_12720,N_12623,N_12571);
nand U12721 (N_12721,N_12634,N_12494);
xnor U12722 (N_12722,N_12537,N_12629);
nand U12723 (N_12723,N_12535,N_12568);
or U12724 (N_12724,N_12607,N_12613);
and U12725 (N_12725,N_12610,N_12565);
or U12726 (N_12726,N_12590,N_12520);
nand U12727 (N_12727,N_12588,N_12632);
nor U12728 (N_12728,N_12598,N_12512);
nand U12729 (N_12729,N_12486,N_12501);
and U12730 (N_12730,N_12615,N_12629);
xnor U12731 (N_12731,N_12480,N_12634);
nor U12732 (N_12732,N_12586,N_12613);
and U12733 (N_12733,N_12495,N_12577);
xor U12734 (N_12734,N_12498,N_12634);
nand U12735 (N_12735,N_12505,N_12589);
or U12736 (N_12736,N_12567,N_12553);
nor U12737 (N_12737,N_12487,N_12617);
or U12738 (N_12738,N_12639,N_12580);
nand U12739 (N_12739,N_12611,N_12628);
nor U12740 (N_12740,N_12588,N_12637);
nand U12741 (N_12741,N_12588,N_12529);
xor U12742 (N_12742,N_12541,N_12577);
nand U12743 (N_12743,N_12555,N_12540);
or U12744 (N_12744,N_12595,N_12604);
and U12745 (N_12745,N_12531,N_12609);
xnor U12746 (N_12746,N_12515,N_12533);
nor U12747 (N_12747,N_12595,N_12627);
nor U12748 (N_12748,N_12534,N_12635);
or U12749 (N_12749,N_12561,N_12540);
or U12750 (N_12750,N_12519,N_12620);
xor U12751 (N_12751,N_12634,N_12515);
nand U12752 (N_12752,N_12532,N_12606);
or U12753 (N_12753,N_12527,N_12556);
and U12754 (N_12754,N_12615,N_12491);
nor U12755 (N_12755,N_12543,N_12492);
or U12756 (N_12756,N_12490,N_12631);
or U12757 (N_12757,N_12569,N_12582);
nor U12758 (N_12758,N_12542,N_12567);
nand U12759 (N_12759,N_12582,N_12590);
nor U12760 (N_12760,N_12586,N_12574);
or U12761 (N_12761,N_12593,N_12610);
or U12762 (N_12762,N_12526,N_12508);
or U12763 (N_12763,N_12512,N_12521);
nor U12764 (N_12764,N_12579,N_12616);
and U12765 (N_12765,N_12567,N_12514);
nor U12766 (N_12766,N_12481,N_12535);
nor U12767 (N_12767,N_12618,N_12582);
or U12768 (N_12768,N_12494,N_12547);
xnor U12769 (N_12769,N_12637,N_12607);
nor U12770 (N_12770,N_12605,N_12596);
or U12771 (N_12771,N_12525,N_12501);
nand U12772 (N_12772,N_12542,N_12541);
xor U12773 (N_12773,N_12503,N_12625);
or U12774 (N_12774,N_12576,N_12483);
xor U12775 (N_12775,N_12532,N_12619);
xor U12776 (N_12776,N_12562,N_12552);
and U12777 (N_12777,N_12583,N_12633);
and U12778 (N_12778,N_12579,N_12604);
nand U12779 (N_12779,N_12613,N_12557);
nand U12780 (N_12780,N_12611,N_12567);
nand U12781 (N_12781,N_12599,N_12487);
or U12782 (N_12782,N_12616,N_12581);
and U12783 (N_12783,N_12631,N_12498);
and U12784 (N_12784,N_12521,N_12599);
xor U12785 (N_12785,N_12614,N_12588);
nand U12786 (N_12786,N_12564,N_12511);
nor U12787 (N_12787,N_12521,N_12551);
or U12788 (N_12788,N_12604,N_12522);
and U12789 (N_12789,N_12537,N_12543);
nand U12790 (N_12790,N_12490,N_12518);
xor U12791 (N_12791,N_12514,N_12616);
or U12792 (N_12792,N_12587,N_12609);
xor U12793 (N_12793,N_12630,N_12559);
or U12794 (N_12794,N_12505,N_12555);
and U12795 (N_12795,N_12636,N_12519);
nor U12796 (N_12796,N_12615,N_12508);
and U12797 (N_12797,N_12522,N_12492);
and U12798 (N_12798,N_12480,N_12611);
and U12799 (N_12799,N_12617,N_12554);
or U12800 (N_12800,N_12658,N_12797);
or U12801 (N_12801,N_12776,N_12774);
nand U12802 (N_12802,N_12681,N_12722);
or U12803 (N_12803,N_12781,N_12720);
and U12804 (N_12804,N_12771,N_12726);
nand U12805 (N_12805,N_12783,N_12696);
nand U12806 (N_12806,N_12685,N_12687);
xor U12807 (N_12807,N_12698,N_12772);
and U12808 (N_12808,N_12659,N_12709);
and U12809 (N_12809,N_12680,N_12728);
nand U12810 (N_12810,N_12782,N_12676);
nand U12811 (N_12811,N_12751,N_12770);
nand U12812 (N_12812,N_12647,N_12725);
or U12813 (N_12813,N_12729,N_12759);
nor U12814 (N_12814,N_12663,N_12796);
nor U12815 (N_12815,N_12778,N_12790);
and U12816 (N_12816,N_12657,N_12747);
and U12817 (N_12817,N_12674,N_12758);
xnor U12818 (N_12818,N_12789,N_12749);
nand U12819 (N_12819,N_12712,N_12718);
nand U12820 (N_12820,N_12703,N_12649);
or U12821 (N_12821,N_12668,N_12692);
nor U12822 (N_12822,N_12742,N_12645);
nor U12823 (N_12823,N_12708,N_12702);
nor U12824 (N_12824,N_12740,N_12661);
nor U12825 (N_12825,N_12727,N_12723);
nor U12826 (N_12826,N_12786,N_12684);
and U12827 (N_12827,N_12799,N_12756);
and U12828 (N_12828,N_12648,N_12646);
xnor U12829 (N_12829,N_12643,N_12675);
and U12830 (N_12830,N_12662,N_12795);
nand U12831 (N_12831,N_12739,N_12752);
or U12832 (N_12832,N_12665,N_12761);
nand U12833 (N_12833,N_12719,N_12679);
nand U12834 (N_12834,N_12715,N_12717);
nor U12835 (N_12835,N_12644,N_12732);
nor U12836 (N_12836,N_12706,N_12653);
or U12837 (N_12837,N_12753,N_12773);
or U12838 (N_12838,N_12656,N_12682);
or U12839 (N_12839,N_12735,N_12699);
nand U12840 (N_12840,N_12677,N_12791);
xnor U12841 (N_12841,N_12784,N_12689);
xnor U12842 (N_12842,N_12678,N_12793);
xnor U12843 (N_12843,N_12711,N_12721);
nand U12844 (N_12844,N_12750,N_12755);
xnor U12845 (N_12845,N_12762,N_12686);
xnor U12846 (N_12846,N_12780,N_12670);
nor U12847 (N_12847,N_12787,N_12650);
and U12848 (N_12848,N_12705,N_12757);
or U12849 (N_12849,N_12764,N_12700);
nor U12850 (N_12850,N_12769,N_12748);
nand U12851 (N_12851,N_12792,N_12736);
or U12852 (N_12852,N_12669,N_12775);
nor U12853 (N_12853,N_12642,N_12743);
and U12854 (N_12854,N_12697,N_12737);
nand U12855 (N_12855,N_12690,N_12651);
nand U12856 (N_12856,N_12741,N_12714);
nand U12857 (N_12857,N_12660,N_12673);
xor U12858 (N_12858,N_12777,N_12754);
or U12859 (N_12859,N_12733,N_12655);
or U12860 (N_12860,N_12652,N_12746);
and U12861 (N_12861,N_12738,N_12734);
nor U12862 (N_12862,N_12767,N_12768);
nor U12863 (N_12863,N_12760,N_12691);
nor U12864 (N_12864,N_12765,N_12779);
or U12865 (N_12865,N_12664,N_12788);
nor U12866 (N_12866,N_12704,N_12724);
and U12867 (N_12867,N_12671,N_12701);
nand U12868 (N_12868,N_12785,N_12667);
xor U12869 (N_12869,N_12654,N_12707);
nand U12870 (N_12870,N_12763,N_12683);
nor U12871 (N_12871,N_12688,N_12798);
nor U12872 (N_12872,N_12730,N_12766);
or U12873 (N_12873,N_12744,N_12640);
nor U12874 (N_12874,N_12794,N_12716);
and U12875 (N_12875,N_12713,N_12710);
xor U12876 (N_12876,N_12666,N_12672);
and U12877 (N_12877,N_12694,N_12693);
xnor U12878 (N_12878,N_12695,N_12745);
nor U12879 (N_12879,N_12731,N_12641);
nor U12880 (N_12880,N_12705,N_12751);
and U12881 (N_12881,N_12738,N_12674);
nand U12882 (N_12882,N_12659,N_12758);
or U12883 (N_12883,N_12651,N_12718);
nand U12884 (N_12884,N_12753,N_12781);
nand U12885 (N_12885,N_12673,N_12785);
nor U12886 (N_12886,N_12699,N_12713);
and U12887 (N_12887,N_12665,N_12759);
and U12888 (N_12888,N_12770,N_12686);
nand U12889 (N_12889,N_12779,N_12737);
and U12890 (N_12890,N_12654,N_12745);
and U12891 (N_12891,N_12721,N_12771);
xnor U12892 (N_12892,N_12737,N_12730);
and U12893 (N_12893,N_12775,N_12688);
nor U12894 (N_12894,N_12749,N_12675);
nand U12895 (N_12895,N_12752,N_12720);
and U12896 (N_12896,N_12645,N_12749);
xor U12897 (N_12897,N_12676,N_12691);
and U12898 (N_12898,N_12745,N_12688);
nor U12899 (N_12899,N_12750,N_12653);
nor U12900 (N_12900,N_12764,N_12741);
and U12901 (N_12901,N_12642,N_12696);
nand U12902 (N_12902,N_12672,N_12660);
or U12903 (N_12903,N_12737,N_12703);
xor U12904 (N_12904,N_12710,N_12783);
xor U12905 (N_12905,N_12756,N_12711);
or U12906 (N_12906,N_12703,N_12760);
and U12907 (N_12907,N_12643,N_12640);
or U12908 (N_12908,N_12760,N_12704);
nor U12909 (N_12909,N_12780,N_12786);
and U12910 (N_12910,N_12657,N_12690);
and U12911 (N_12911,N_12733,N_12738);
nand U12912 (N_12912,N_12688,N_12715);
and U12913 (N_12913,N_12795,N_12766);
and U12914 (N_12914,N_12721,N_12773);
xnor U12915 (N_12915,N_12798,N_12746);
nor U12916 (N_12916,N_12652,N_12797);
nor U12917 (N_12917,N_12742,N_12738);
nor U12918 (N_12918,N_12788,N_12679);
nand U12919 (N_12919,N_12727,N_12695);
nor U12920 (N_12920,N_12719,N_12786);
nor U12921 (N_12921,N_12791,N_12675);
nand U12922 (N_12922,N_12756,N_12699);
nor U12923 (N_12923,N_12744,N_12677);
or U12924 (N_12924,N_12663,N_12643);
xnor U12925 (N_12925,N_12661,N_12796);
nand U12926 (N_12926,N_12650,N_12720);
or U12927 (N_12927,N_12780,N_12647);
or U12928 (N_12928,N_12724,N_12730);
nand U12929 (N_12929,N_12695,N_12710);
nor U12930 (N_12930,N_12739,N_12700);
xor U12931 (N_12931,N_12777,N_12680);
xnor U12932 (N_12932,N_12684,N_12659);
and U12933 (N_12933,N_12679,N_12673);
nand U12934 (N_12934,N_12657,N_12792);
or U12935 (N_12935,N_12692,N_12746);
and U12936 (N_12936,N_12746,N_12674);
nor U12937 (N_12937,N_12709,N_12762);
and U12938 (N_12938,N_12796,N_12669);
nand U12939 (N_12939,N_12770,N_12792);
xor U12940 (N_12940,N_12656,N_12681);
nand U12941 (N_12941,N_12645,N_12757);
nand U12942 (N_12942,N_12777,N_12794);
nor U12943 (N_12943,N_12771,N_12673);
nand U12944 (N_12944,N_12670,N_12698);
and U12945 (N_12945,N_12790,N_12718);
xnor U12946 (N_12946,N_12692,N_12712);
xor U12947 (N_12947,N_12702,N_12726);
xnor U12948 (N_12948,N_12775,N_12757);
or U12949 (N_12949,N_12680,N_12705);
nand U12950 (N_12950,N_12693,N_12710);
nor U12951 (N_12951,N_12687,N_12670);
nand U12952 (N_12952,N_12797,N_12766);
or U12953 (N_12953,N_12687,N_12732);
or U12954 (N_12954,N_12756,N_12643);
nand U12955 (N_12955,N_12714,N_12761);
xor U12956 (N_12956,N_12645,N_12642);
xnor U12957 (N_12957,N_12706,N_12658);
nand U12958 (N_12958,N_12758,N_12787);
nor U12959 (N_12959,N_12779,N_12723);
nor U12960 (N_12960,N_12847,N_12884);
or U12961 (N_12961,N_12887,N_12947);
or U12962 (N_12962,N_12806,N_12914);
and U12963 (N_12963,N_12880,N_12826);
nor U12964 (N_12964,N_12859,N_12916);
xor U12965 (N_12965,N_12902,N_12955);
or U12966 (N_12966,N_12801,N_12839);
or U12967 (N_12967,N_12926,N_12910);
nand U12968 (N_12968,N_12860,N_12900);
xor U12969 (N_12969,N_12848,N_12824);
xnor U12970 (N_12970,N_12869,N_12875);
and U12971 (N_12971,N_12931,N_12933);
nand U12972 (N_12972,N_12903,N_12928);
or U12973 (N_12973,N_12908,N_12845);
and U12974 (N_12974,N_12890,N_12956);
nand U12975 (N_12975,N_12800,N_12936);
or U12976 (N_12976,N_12812,N_12838);
and U12977 (N_12977,N_12924,N_12815);
nor U12978 (N_12978,N_12937,N_12959);
nand U12979 (N_12979,N_12889,N_12823);
and U12980 (N_12980,N_12822,N_12868);
xor U12981 (N_12981,N_12810,N_12940);
and U12982 (N_12982,N_12846,N_12907);
xnor U12983 (N_12983,N_12896,N_12917);
nor U12984 (N_12984,N_12817,N_12865);
or U12985 (N_12985,N_12870,N_12891);
xor U12986 (N_12986,N_12851,N_12909);
nor U12987 (N_12987,N_12912,N_12864);
or U12988 (N_12988,N_12854,N_12813);
or U12989 (N_12989,N_12898,N_12888);
xnor U12990 (N_12990,N_12828,N_12837);
or U12991 (N_12991,N_12836,N_12948);
and U12992 (N_12992,N_12821,N_12877);
xnor U12993 (N_12993,N_12946,N_12951);
nor U12994 (N_12994,N_12952,N_12901);
nand U12995 (N_12995,N_12945,N_12829);
and U12996 (N_12996,N_12930,N_12893);
xnor U12997 (N_12997,N_12881,N_12911);
nand U12998 (N_12998,N_12835,N_12866);
or U12999 (N_12999,N_12805,N_12819);
nor U13000 (N_13000,N_12939,N_12953);
and U13001 (N_13001,N_12905,N_12825);
nor U13002 (N_13002,N_12906,N_12919);
nor U13003 (N_13003,N_12957,N_12904);
xnor U13004 (N_13004,N_12932,N_12941);
xnor U13005 (N_13005,N_12804,N_12915);
nor U13006 (N_13006,N_12850,N_12954);
and U13007 (N_13007,N_12811,N_12934);
and U13008 (N_13008,N_12856,N_12913);
and U13009 (N_13009,N_12925,N_12899);
and U13010 (N_13010,N_12807,N_12886);
or U13011 (N_13011,N_12938,N_12814);
nand U13012 (N_13012,N_12834,N_12927);
nand U13013 (N_13013,N_12853,N_12923);
and U13014 (N_13014,N_12879,N_12894);
and U13015 (N_13015,N_12892,N_12943);
nand U13016 (N_13016,N_12861,N_12885);
and U13017 (N_13017,N_12922,N_12831);
or U13018 (N_13018,N_12882,N_12827);
or U13019 (N_13019,N_12874,N_12840);
nand U13020 (N_13020,N_12832,N_12958);
nor U13021 (N_13021,N_12867,N_12862);
nand U13022 (N_13022,N_12872,N_12802);
nand U13023 (N_13023,N_12942,N_12852);
or U13024 (N_13024,N_12873,N_12844);
nor U13025 (N_13025,N_12833,N_12918);
nand U13026 (N_13026,N_12808,N_12883);
or U13027 (N_13027,N_12871,N_12809);
nand U13028 (N_13028,N_12949,N_12878);
xor U13029 (N_13029,N_12858,N_12950);
nor U13030 (N_13030,N_12849,N_12857);
nor U13031 (N_13031,N_12876,N_12820);
xnor U13032 (N_13032,N_12830,N_12803);
or U13033 (N_13033,N_12816,N_12841);
and U13034 (N_13034,N_12842,N_12935);
and U13035 (N_13035,N_12818,N_12895);
or U13036 (N_13036,N_12929,N_12863);
nor U13037 (N_13037,N_12897,N_12944);
nand U13038 (N_13038,N_12920,N_12843);
and U13039 (N_13039,N_12855,N_12921);
or U13040 (N_13040,N_12861,N_12805);
or U13041 (N_13041,N_12936,N_12875);
xor U13042 (N_13042,N_12854,N_12834);
nand U13043 (N_13043,N_12909,N_12899);
xor U13044 (N_13044,N_12916,N_12924);
nor U13045 (N_13045,N_12803,N_12882);
and U13046 (N_13046,N_12878,N_12810);
and U13047 (N_13047,N_12879,N_12885);
and U13048 (N_13048,N_12846,N_12874);
and U13049 (N_13049,N_12909,N_12866);
xnor U13050 (N_13050,N_12868,N_12947);
and U13051 (N_13051,N_12930,N_12858);
nand U13052 (N_13052,N_12866,N_12956);
or U13053 (N_13053,N_12895,N_12890);
xnor U13054 (N_13054,N_12849,N_12884);
or U13055 (N_13055,N_12934,N_12864);
xor U13056 (N_13056,N_12872,N_12939);
nand U13057 (N_13057,N_12933,N_12908);
nor U13058 (N_13058,N_12875,N_12957);
and U13059 (N_13059,N_12856,N_12896);
and U13060 (N_13060,N_12830,N_12831);
and U13061 (N_13061,N_12831,N_12958);
or U13062 (N_13062,N_12905,N_12942);
xnor U13063 (N_13063,N_12824,N_12882);
or U13064 (N_13064,N_12954,N_12934);
and U13065 (N_13065,N_12802,N_12896);
nor U13066 (N_13066,N_12880,N_12903);
xnor U13067 (N_13067,N_12843,N_12907);
nor U13068 (N_13068,N_12888,N_12807);
or U13069 (N_13069,N_12889,N_12846);
or U13070 (N_13070,N_12843,N_12828);
nand U13071 (N_13071,N_12900,N_12958);
nor U13072 (N_13072,N_12926,N_12827);
xnor U13073 (N_13073,N_12803,N_12814);
nand U13074 (N_13074,N_12876,N_12928);
nand U13075 (N_13075,N_12920,N_12931);
xnor U13076 (N_13076,N_12954,N_12838);
nor U13077 (N_13077,N_12948,N_12834);
or U13078 (N_13078,N_12889,N_12850);
or U13079 (N_13079,N_12812,N_12872);
xor U13080 (N_13080,N_12804,N_12882);
nor U13081 (N_13081,N_12842,N_12875);
and U13082 (N_13082,N_12876,N_12910);
or U13083 (N_13083,N_12818,N_12943);
nor U13084 (N_13084,N_12848,N_12844);
nand U13085 (N_13085,N_12865,N_12827);
xnor U13086 (N_13086,N_12872,N_12907);
and U13087 (N_13087,N_12876,N_12810);
nor U13088 (N_13088,N_12867,N_12817);
xor U13089 (N_13089,N_12867,N_12893);
xor U13090 (N_13090,N_12887,N_12894);
and U13091 (N_13091,N_12945,N_12861);
xnor U13092 (N_13092,N_12844,N_12813);
nor U13093 (N_13093,N_12901,N_12874);
or U13094 (N_13094,N_12810,N_12861);
nand U13095 (N_13095,N_12908,N_12930);
xnor U13096 (N_13096,N_12834,N_12821);
xor U13097 (N_13097,N_12811,N_12832);
nor U13098 (N_13098,N_12909,N_12805);
xor U13099 (N_13099,N_12908,N_12955);
and U13100 (N_13100,N_12911,N_12800);
nand U13101 (N_13101,N_12910,N_12848);
or U13102 (N_13102,N_12895,N_12921);
nor U13103 (N_13103,N_12803,N_12942);
xnor U13104 (N_13104,N_12901,N_12860);
nor U13105 (N_13105,N_12890,N_12889);
nand U13106 (N_13106,N_12917,N_12894);
nor U13107 (N_13107,N_12940,N_12848);
and U13108 (N_13108,N_12944,N_12859);
nand U13109 (N_13109,N_12800,N_12807);
xor U13110 (N_13110,N_12829,N_12822);
or U13111 (N_13111,N_12954,N_12905);
nor U13112 (N_13112,N_12805,N_12902);
or U13113 (N_13113,N_12820,N_12917);
nor U13114 (N_13114,N_12907,N_12802);
or U13115 (N_13115,N_12877,N_12851);
xor U13116 (N_13116,N_12936,N_12917);
or U13117 (N_13117,N_12899,N_12862);
or U13118 (N_13118,N_12889,N_12948);
nand U13119 (N_13119,N_12819,N_12813);
nor U13120 (N_13120,N_13084,N_12964);
nor U13121 (N_13121,N_12992,N_13035);
or U13122 (N_13122,N_13034,N_13073);
or U13123 (N_13123,N_13054,N_13105);
or U13124 (N_13124,N_12975,N_13050);
nand U13125 (N_13125,N_13060,N_13053);
nor U13126 (N_13126,N_13112,N_13024);
xnor U13127 (N_13127,N_13067,N_12998);
or U13128 (N_13128,N_13007,N_13071);
nor U13129 (N_13129,N_12962,N_13052);
xnor U13130 (N_13130,N_13074,N_13109);
xnor U13131 (N_13131,N_12994,N_12966);
nand U13132 (N_13132,N_13029,N_13064);
nand U13133 (N_13133,N_13015,N_13044);
xnor U13134 (N_13134,N_13104,N_12980);
xnor U13135 (N_13135,N_13041,N_13059);
and U13136 (N_13136,N_12986,N_13062);
and U13137 (N_13137,N_13051,N_13099);
nor U13138 (N_13138,N_13010,N_13043);
nor U13139 (N_13139,N_13090,N_12972);
nand U13140 (N_13140,N_13069,N_12974);
xnor U13141 (N_13141,N_13106,N_13068);
nor U13142 (N_13142,N_13097,N_13083);
xor U13143 (N_13143,N_13037,N_13117);
xor U13144 (N_13144,N_13075,N_13081);
or U13145 (N_13145,N_13020,N_13039);
nor U13146 (N_13146,N_13046,N_13008);
nor U13147 (N_13147,N_12995,N_13065);
or U13148 (N_13148,N_13079,N_12982);
nor U13149 (N_13149,N_13049,N_12973);
and U13150 (N_13150,N_12970,N_13005);
nand U13151 (N_13151,N_13110,N_13027);
and U13152 (N_13152,N_13017,N_13061);
xor U13153 (N_13153,N_13002,N_13025);
nand U13154 (N_13154,N_13078,N_13114);
and U13155 (N_13155,N_12960,N_13119);
and U13156 (N_13156,N_13111,N_13019);
xor U13157 (N_13157,N_13047,N_13042);
xnor U13158 (N_13158,N_13108,N_13077);
nor U13159 (N_13159,N_12983,N_13040);
xnor U13160 (N_13160,N_13000,N_13016);
or U13161 (N_13161,N_12990,N_13085);
nand U13162 (N_13162,N_13102,N_13080);
or U13163 (N_13163,N_12967,N_13095);
xnor U13164 (N_13164,N_13004,N_13006);
or U13165 (N_13165,N_13036,N_13056);
nand U13166 (N_13166,N_13014,N_12971);
nand U13167 (N_13167,N_13072,N_12987);
xor U13168 (N_13168,N_13115,N_12999);
nand U13169 (N_13169,N_13058,N_13116);
or U13170 (N_13170,N_13107,N_12981);
nand U13171 (N_13171,N_13031,N_12979);
or U13172 (N_13172,N_13030,N_12989);
and U13173 (N_13173,N_13082,N_13089);
and U13174 (N_13174,N_13100,N_13018);
nor U13175 (N_13175,N_13101,N_12985);
or U13176 (N_13176,N_12968,N_12997);
or U13177 (N_13177,N_13003,N_13066);
or U13178 (N_13178,N_13011,N_13094);
and U13179 (N_13179,N_13086,N_12988);
nor U13180 (N_13180,N_12991,N_13118);
nand U13181 (N_13181,N_13022,N_13033);
and U13182 (N_13182,N_13001,N_13070);
and U13183 (N_13183,N_13009,N_12963);
xor U13184 (N_13184,N_13045,N_13091);
nor U13185 (N_13185,N_13092,N_13012);
and U13186 (N_13186,N_13026,N_13087);
or U13187 (N_13187,N_13023,N_13088);
and U13188 (N_13188,N_13096,N_13032);
nand U13189 (N_13189,N_12984,N_12961);
or U13190 (N_13190,N_12965,N_13076);
xnor U13191 (N_13191,N_13055,N_13093);
or U13192 (N_13192,N_13021,N_13028);
nor U13193 (N_13193,N_13038,N_13063);
xor U13194 (N_13194,N_12978,N_13098);
nand U13195 (N_13195,N_13057,N_12996);
nand U13196 (N_13196,N_12976,N_12977);
and U13197 (N_13197,N_13113,N_12969);
nor U13198 (N_13198,N_13048,N_12993);
nand U13199 (N_13199,N_13013,N_13103);
nand U13200 (N_13200,N_12981,N_13004);
nand U13201 (N_13201,N_13102,N_12987);
nor U13202 (N_13202,N_13086,N_13109);
nand U13203 (N_13203,N_13071,N_13094);
xor U13204 (N_13204,N_13089,N_12988);
nor U13205 (N_13205,N_12969,N_12974);
nand U13206 (N_13206,N_13061,N_12984);
or U13207 (N_13207,N_13079,N_13100);
or U13208 (N_13208,N_13003,N_13113);
or U13209 (N_13209,N_12962,N_13102);
and U13210 (N_13210,N_12976,N_13029);
xnor U13211 (N_13211,N_13081,N_13068);
or U13212 (N_13212,N_13076,N_13119);
nand U13213 (N_13213,N_12986,N_13053);
and U13214 (N_13214,N_13045,N_12967);
nand U13215 (N_13215,N_13076,N_13086);
xor U13216 (N_13216,N_13044,N_13013);
nor U13217 (N_13217,N_12995,N_13019);
and U13218 (N_13218,N_12976,N_13108);
xor U13219 (N_13219,N_13074,N_12981);
nor U13220 (N_13220,N_13048,N_13037);
nor U13221 (N_13221,N_13068,N_13064);
or U13222 (N_13222,N_13008,N_13105);
nor U13223 (N_13223,N_12986,N_13095);
nor U13224 (N_13224,N_13043,N_12962);
nor U13225 (N_13225,N_12997,N_12999);
or U13226 (N_13226,N_13049,N_12986);
and U13227 (N_13227,N_12975,N_13027);
and U13228 (N_13228,N_12984,N_13028);
xor U13229 (N_13229,N_13077,N_13117);
and U13230 (N_13230,N_13016,N_13026);
nand U13231 (N_13231,N_13048,N_13044);
xnor U13232 (N_13232,N_12973,N_12988);
nand U13233 (N_13233,N_13062,N_13014);
and U13234 (N_13234,N_13028,N_13016);
xor U13235 (N_13235,N_13119,N_13063);
or U13236 (N_13236,N_13021,N_13024);
nand U13237 (N_13237,N_13071,N_13030);
xor U13238 (N_13238,N_13100,N_13007);
and U13239 (N_13239,N_12988,N_13030);
or U13240 (N_13240,N_12964,N_12965);
and U13241 (N_13241,N_13032,N_13067);
xor U13242 (N_13242,N_13052,N_12990);
or U13243 (N_13243,N_12982,N_13053);
and U13244 (N_13244,N_13023,N_13005);
or U13245 (N_13245,N_13103,N_13047);
xor U13246 (N_13246,N_12964,N_13109);
xor U13247 (N_13247,N_12983,N_13109);
xor U13248 (N_13248,N_13104,N_13076);
nor U13249 (N_13249,N_13015,N_13039);
or U13250 (N_13250,N_12962,N_12985);
xor U13251 (N_13251,N_13054,N_12990);
or U13252 (N_13252,N_12987,N_13117);
xor U13253 (N_13253,N_13000,N_13028);
or U13254 (N_13254,N_13068,N_13082);
xor U13255 (N_13255,N_12994,N_12982);
nor U13256 (N_13256,N_13057,N_13061);
nor U13257 (N_13257,N_12973,N_13031);
and U13258 (N_13258,N_13029,N_13104);
nor U13259 (N_13259,N_13034,N_13112);
or U13260 (N_13260,N_13087,N_13053);
nor U13261 (N_13261,N_12991,N_13085);
xor U13262 (N_13262,N_12960,N_13024);
xor U13263 (N_13263,N_13031,N_13034);
and U13264 (N_13264,N_12995,N_13063);
xnor U13265 (N_13265,N_13102,N_13096);
nor U13266 (N_13266,N_12995,N_13004);
xnor U13267 (N_13267,N_12960,N_13087);
xor U13268 (N_13268,N_13084,N_12988);
nor U13269 (N_13269,N_12992,N_13014);
and U13270 (N_13270,N_13047,N_13073);
and U13271 (N_13271,N_13049,N_13092);
or U13272 (N_13272,N_12960,N_13057);
nor U13273 (N_13273,N_13088,N_13027);
and U13274 (N_13274,N_13078,N_12960);
nand U13275 (N_13275,N_13042,N_13077);
or U13276 (N_13276,N_13081,N_12990);
or U13277 (N_13277,N_12978,N_13067);
and U13278 (N_13278,N_13004,N_13089);
or U13279 (N_13279,N_13087,N_13047);
nand U13280 (N_13280,N_13254,N_13126);
and U13281 (N_13281,N_13217,N_13139);
nor U13282 (N_13282,N_13136,N_13182);
nor U13283 (N_13283,N_13219,N_13207);
and U13284 (N_13284,N_13195,N_13205);
nor U13285 (N_13285,N_13122,N_13143);
nand U13286 (N_13286,N_13170,N_13245);
or U13287 (N_13287,N_13134,N_13215);
and U13288 (N_13288,N_13222,N_13120);
xor U13289 (N_13289,N_13187,N_13202);
nor U13290 (N_13290,N_13204,N_13151);
nand U13291 (N_13291,N_13121,N_13144);
and U13292 (N_13292,N_13156,N_13232);
nand U13293 (N_13293,N_13211,N_13190);
nand U13294 (N_13294,N_13242,N_13208);
nor U13295 (N_13295,N_13133,N_13234);
or U13296 (N_13296,N_13150,N_13199);
nor U13297 (N_13297,N_13168,N_13224);
xnor U13298 (N_13298,N_13159,N_13175);
or U13299 (N_13299,N_13177,N_13243);
and U13300 (N_13300,N_13181,N_13226);
or U13301 (N_13301,N_13161,N_13130);
and U13302 (N_13302,N_13228,N_13271);
or U13303 (N_13303,N_13153,N_13200);
xor U13304 (N_13304,N_13146,N_13141);
and U13305 (N_13305,N_13174,N_13166);
xor U13306 (N_13306,N_13259,N_13236);
or U13307 (N_13307,N_13192,N_13152);
xor U13308 (N_13308,N_13276,N_13165);
xor U13309 (N_13309,N_13191,N_13258);
nand U13310 (N_13310,N_13266,N_13172);
nand U13311 (N_13311,N_13233,N_13251);
or U13312 (N_13312,N_13273,N_13262);
xnor U13313 (N_13313,N_13230,N_13209);
or U13314 (N_13314,N_13124,N_13220);
nand U13315 (N_13315,N_13196,N_13248);
xor U13316 (N_13316,N_13264,N_13188);
nor U13317 (N_13317,N_13274,N_13162);
and U13318 (N_13318,N_13123,N_13193);
and U13319 (N_13319,N_13127,N_13163);
nand U13320 (N_13320,N_13157,N_13231);
or U13321 (N_13321,N_13149,N_13125);
nand U13322 (N_13322,N_13275,N_13229);
or U13323 (N_13323,N_13221,N_13160);
nand U13324 (N_13324,N_13238,N_13171);
xnor U13325 (N_13325,N_13135,N_13189);
or U13326 (N_13326,N_13272,N_13213);
nor U13327 (N_13327,N_13223,N_13255);
xor U13328 (N_13328,N_13131,N_13206);
nor U13329 (N_13329,N_13216,N_13277);
xor U13330 (N_13330,N_13173,N_13183);
or U13331 (N_13331,N_13180,N_13145);
or U13332 (N_13332,N_13197,N_13218);
nor U13333 (N_13333,N_13278,N_13227);
or U13334 (N_13334,N_13140,N_13142);
and U13335 (N_13335,N_13267,N_13203);
xor U13336 (N_13336,N_13128,N_13179);
xnor U13337 (N_13337,N_13263,N_13270);
nor U13338 (N_13338,N_13214,N_13167);
nand U13339 (N_13339,N_13178,N_13256);
nand U13340 (N_13340,N_13212,N_13155);
and U13341 (N_13341,N_13194,N_13184);
nand U13342 (N_13342,N_13246,N_13137);
and U13343 (N_13343,N_13129,N_13225);
nand U13344 (N_13344,N_13210,N_13148);
nand U13345 (N_13345,N_13252,N_13249);
xnor U13346 (N_13346,N_13261,N_13247);
or U13347 (N_13347,N_13169,N_13147);
and U13348 (N_13348,N_13132,N_13138);
xor U13349 (N_13349,N_13269,N_13239);
or U13350 (N_13350,N_13154,N_13198);
nor U13351 (N_13351,N_13279,N_13241);
xnor U13352 (N_13352,N_13265,N_13237);
nand U13353 (N_13353,N_13244,N_13158);
and U13354 (N_13354,N_13268,N_13250);
or U13355 (N_13355,N_13253,N_13185);
nand U13356 (N_13356,N_13240,N_13235);
nand U13357 (N_13357,N_13176,N_13186);
nand U13358 (N_13358,N_13260,N_13257);
nor U13359 (N_13359,N_13201,N_13164);
or U13360 (N_13360,N_13187,N_13166);
nor U13361 (N_13361,N_13127,N_13126);
or U13362 (N_13362,N_13126,N_13122);
nor U13363 (N_13363,N_13187,N_13193);
or U13364 (N_13364,N_13248,N_13251);
and U13365 (N_13365,N_13192,N_13234);
nor U13366 (N_13366,N_13246,N_13227);
nand U13367 (N_13367,N_13175,N_13237);
nor U13368 (N_13368,N_13275,N_13196);
xnor U13369 (N_13369,N_13260,N_13134);
xor U13370 (N_13370,N_13240,N_13204);
nor U13371 (N_13371,N_13130,N_13199);
xor U13372 (N_13372,N_13161,N_13224);
and U13373 (N_13373,N_13125,N_13185);
or U13374 (N_13374,N_13130,N_13126);
xnor U13375 (N_13375,N_13210,N_13122);
nand U13376 (N_13376,N_13244,N_13212);
xor U13377 (N_13377,N_13168,N_13249);
xnor U13378 (N_13378,N_13122,N_13217);
or U13379 (N_13379,N_13222,N_13159);
or U13380 (N_13380,N_13172,N_13156);
nor U13381 (N_13381,N_13245,N_13157);
nor U13382 (N_13382,N_13175,N_13154);
nand U13383 (N_13383,N_13215,N_13226);
and U13384 (N_13384,N_13206,N_13172);
nand U13385 (N_13385,N_13129,N_13196);
xnor U13386 (N_13386,N_13168,N_13259);
nand U13387 (N_13387,N_13123,N_13190);
xor U13388 (N_13388,N_13240,N_13162);
and U13389 (N_13389,N_13146,N_13219);
nand U13390 (N_13390,N_13221,N_13252);
and U13391 (N_13391,N_13234,N_13254);
and U13392 (N_13392,N_13181,N_13216);
xor U13393 (N_13393,N_13274,N_13135);
xor U13394 (N_13394,N_13124,N_13277);
nor U13395 (N_13395,N_13198,N_13134);
nand U13396 (N_13396,N_13230,N_13271);
or U13397 (N_13397,N_13262,N_13125);
xnor U13398 (N_13398,N_13217,N_13192);
and U13399 (N_13399,N_13209,N_13160);
and U13400 (N_13400,N_13159,N_13258);
xnor U13401 (N_13401,N_13139,N_13266);
and U13402 (N_13402,N_13200,N_13144);
or U13403 (N_13403,N_13123,N_13272);
or U13404 (N_13404,N_13256,N_13169);
xnor U13405 (N_13405,N_13155,N_13278);
nor U13406 (N_13406,N_13269,N_13252);
and U13407 (N_13407,N_13183,N_13130);
nand U13408 (N_13408,N_13237,N_13124);
and U13409 (N_13409,N_13129,N_13141);
xnor U13410 (N_13410,N_13126,N_13273);
and U13411 (N_13411,N_13138,N_13137);
nand U13412 (N_13412,N_13126,N_13192);
xnor U13413 (N_13413,N_13245,N_13172);
nand U13414 (N_13414,N_13152,N_13275);
nor U13415 (N_13415,N_13240,N_13126);
nor U13416 (N_13416,N_13253,N_13227);
xnor U13417 (N_13417,N_13176,N_13181);
nand U13418 (N_13418,N_13277,N_13278);
xnor U13419 (N_13419,N_13242,N_13202);
nand U13420 (N_13420,N_13255,N_13142);
nand U13421 (N_13421,N_13200,N_13217);
nand U13422 (N_13422,N_13246,N_13165);
or U13423 (N_13423,N_13262,N_13129);
or U13424 (N_13424,N_13203,N_13152);
xnor U13425 (N_13425,N_13178,N_13152);
and U13426 (N_13426,N_13170,N_13212);
xor U13427 (N_13427,N_13133,N_13195);
and U13428 (N_13428,N_13218,N_13264);
nand U13429 (N_13429,N_13250,N_13219);
and U13430 (N_13430,N_13196,N_13137);
nand U13431 (N_13431,N_13164,N_13203);
xor U13432 (N_13432,N_13274,N_13167);
nor U13433 (N_13433,N_13172,N_13232);
and U13434 (N_13434,N_13187,N_13213);
or U13435 (N_13435,N_13279,N_13182);
nand U13436 (N_13436,N_13239,N_13142);
or U13437 (N_13437,N_13260,N_13221);
xor U13438 (N_13438,N_13167,N_13222);
nor U13439 (N_13439,N_13198,N_13197);
and U13440 (N_13440,N_13407,N_13439);
and U13441 (N_13441,N_13384,N_13317);
xor U13442 (N_13442,N_13423,N_13352);
or U13443 (N_13443,N_13296,N_13420);
nor U13444 (N_13444,N_13324,N_13340);
nor U13445 (N_13445,N_13343,N_13393);
and U13446 (N_13446,N_13356,N_13285);
and U13447 (N_13447,N_13435,N_13398);
or U13448 (N_13448,N_13344,N_13389);
xor U13449 (N_13449,N_13327,N_13399);
nor U13450 (N_13450,N_13403,N_13417);
xnor U13451 (N_13451,N_13377,N_13336);
and U13452 (N_13452,N_13284,N_13280);
and U13453 (N_13453,N_13319,N_13325);
and U13454 (N_13454,N_13294,N_13429);
nand U13455 (N_13455,N_13363,N_13383);
nor U13456 (N_13456,N_13388,N_13306);
and U13457 (N_13457,N_13304,N_13412);
and U13458 (N_13458,N_13333,N_13282);
and U13459 (N_13459,N_13436,N_13381);
and U13460 (N_13460,N_13307,N_13286);
nor U13461 (N_13461,N_13416,N_13390);
or U13462 (N_13462,N_13359,N_13301);
nand U13463 (N_13463,N_13370,N_13376);
and U13464 (N_13464,N_13322,N_13332);
nand U13465 (N_13465,N_13318,N_13335);
or U13466 (N_13466,N_13334,N_13313);
xor U13467 (N_13467,N_13374,N_13380);
and U13468 (N_13468,N_13297,N_13346);
nor U13469 (N_13469,N_13339,N_13326);
xnor U13470 (N_13470,N_13303,N_13409);
or U13471 (N_13471,N_13310,N_13347);
and U13472 (N_13472,N_13353,N_13316);
and U13473 (N_13473,N_13338,N_13411);
xor U13474 (N_13474,N_13345,N_13350);
xnor U13475 (N_13475,N_13314,N_13361);
nand U13476 (N_13476,N_13298,N_13305);
and U13477 (N_13477,N_13373,N_13372);
nand U13478 (N_13478,N_13364,N_13438);
or U13479 (N_13479,N_13437,N_13424);
or U13480 (N_13480,N_13422,N_13360);
and U13481 (N_13481,N_13369,N_13315);
or U13482 (N_13482,N_13431,N_13378);
nand U13483 (N_13483,N_13329,N_13302);
nand U13484 (N_13484,N_13392,N_13362);
xnor U13485 (N_13485,N_13321,N_13391);
nor U13486 (N_13486,N_13295,N_13426);
nor U13487 (N_13487,N_13367,N_13366);
nor U13488 (N_13488,N_13404,N_13405);
xor U13489 (N_13489,N_13349,N_13331);
and U13490 (N_13490,N_13368,N_13351);
nand U13491 (N_13491,N_13291,N_13348);
and U13492 (N_13492,N_13311,N_13410);
or U13493 (N_13493,N_13402,N_13365);
and U13494 (N_13494,N_13323,N_13421);
xor U13495 (N_13495,N_13418,N_13379);
nor U13496 (N_13496,N_13342,N_13288);
or U13497 (N_13497,N_13292,N_13408);
nand U13498 (N_13498,N_13414,N_13293);
nor U13499 (N_13499,N_13397,N_13427);
or U13500 (N_13500,N_13406,N_13434);
nor U13501 (N_13501,N_13394,N_13309);
nand U13502 (N_13502,N_13396,N_13419);
or U13503 (N_13503,N_13386,N_13283);
or U13504 (N_13504,N_13430,N_13308);
or U13505 (N_13505,N_13299,N_13312);
or U13506 (N_13506,N_13382,N_13395);
nand U13507 (N_13507,N_13428,N_13415);
nor U13508 (N_13508,N_13432,N_13337);
nand U13509 (N_13509,N_13328,N_13375);
nor U13510 (N_13510,N_13413,N_13433);
xnor U13511 (N_13511,N_13320,N_13400);
nand U13512 (N_13512,N_13300,N_13387);
or U13513 (N_13513,N_13354,N_13355);
or U13514 (N_13514,N_13290,N_13357);
or U13515 (N_13515,N_13358,N_13425);
nand U13516 (N_13516,N_13401,N_13289);
and U13517 (N_13517,N_13287,N_13341);
nand U13518 (N_13518,N_13385,N_13281);
xnor U13519 (N_13519,N_13330,N_13371);
nand U13520 (N_13520,N_13282,N_13416);
or U13521 (N_13521,N_13310,N_13331);
nor U13522 (N_13522,N_13372,N_13364);
xor U13523 (N_13523,N_13311,N_13392);
and U13524 (N_13524,N_13390,N_13439);
nand U13525 (N_13525,N_13389,N_13292);
or U13526 (N_13526,N_13316,N_13312);
and U13527 (N_13527,N_13393,N_13339);
xnor U13528 (N_13528,N_13287,N_13399);
xor U13529 (N_13529,N_13437,N_13394);
xor U13530 (N_13530,N_13427,N_13381);
xnor U13531 (N_13531,N_13360,N_13382);
or U13532 (N_13532,N_13335,N_13340);
nor U13533 (N_13533,N_13403,N_13404);
xor U13534 (N_13534,N_13397,N_13432);
nand U13535 (N_13535,N_13381,N_13414);
xor U13536 (N_13536,N_13354,N_13330);
nand U13537 (N_13537,N_13338,N_13294);
nor U13538 (N_13538,N_13308,N_13307);
xnor U13539 (N_13539,N_13402,N_13341);
xnor U13540 (N_13540,N_13283,N_13309);
xnor U13541 (N_13541,N_13423,N_13366);
xor U13542 (N_13542,N_13304,N_13330);
nor U13543 (N_13543,N_13420,N_13318);
and U13544 (N_13544,N_13391,N_13343);
or U13545 (N_13545,N_13435,N_13373);
or U13546 (N_13546,N_13434,N_13350);
xnor U13547 (N_13547,N_13364,N_13402);
nand U13548 (N_13548,N_13314,N_13283);
or U13549 (N_13549,N_13431,N_13288);
nor U13550 (N_13550,N_13322,N_13320);
and U13551 (N_13551,N_13308,N_13303);
and U13552 (N_13552,N_13398,N_13416);
nand U13553 (N_13553,N_13406,N_13307);
nand U13554 (N_13554,N_13404,N_13355);
nand U13555 (N_13555,N_13290,N_13366);
xor U13556 (N_13556,N_13335,N_13408);
nand U13557 (N_13557,N_13365,N_13315);
nor U13558 (N_13558,N_13431,N_13356);
and U13559 (N_13559,N_13357,N_13412);
nand U13560 (N_13560,N_13401,N_13360);
nor U13561 (N_13561,N_13307,N_13429);
nand U13562 (N_13562,N_13395,N_13310);
and U13563 (N_13563,N_13386,N_13332);
nor U13564 (N_13564,N_13350,N_13404);
or U13565 (N_13565,N_13368,N_13339);
xnor U13566 (N_13566,N_13402,N_13434);
nor U13567 (N_13567,N_13438,N_13310);
xor U13568 (N_13568,N_13315,N_13438);
nand U13569 (N_13569,N_13373,N_13425);
and U13570 (N_13570,N_13425,N_13319);
and U13571 (N_13571,N_13309,N_13386);
or U13572 (N_13572,N_13402,N_13385);
nand U13573 (N_13573,N_13411,N_13316);
nor U13574 (N_13574,N_13350,N_13293);
nor U13575 (N_13575,N_13438,N_13405);
and U13576 (N_13576,N_13317,N_13338);
nor U13577 (N_13577,N_13294,N_13434);
xnor U13578 (N_13578,N_13396,N_13295);
or U13579 (N_13579,N_13419,N_13314);
nor U13580 (N_13580,N_13349,N_13287);
xnor U13581 (N_13581,N_13432,N_13311);
or U13582 (N_13582,N_13308,N_13282);
nand U13583 (N_13583,N_13439,N_13344);
nand U13584 (N_13584,N_13364,N_13411);
or U13585 (N_13585,N_13281,N_13388);
and U13586 (N_13586,N_13320,N_13328);
or U13587 (N_13587,N_13331,N_13335);
xnor U13588 (N_13588,N_13391,N_13299);
xnor U13589 (N_13589,N_13334,N_13372);
xnor U13590 (N_13590,N_13358,N_13361);
nand U13591 (N_13591,N_13353,N_13437);
and U13592 (N_13592,N_13413,N_13373);
nor U13593 (N_13593,N_13356,N_13433);
nor U13594 (N_13594,N_13390,N_13405);
or U13595 (N_13595,N_13299,N_13303);
nand U13596 (N_13596,N_13341,N_13347);
nand U13597 (N_13597,N_13324,N_13354);
or U13598 (N_13598,N_13308,N_13286);
and U13599 (N_13599,N_13318,N_13331);
or U13600 (N_13600,N_13557,N_13472);
and U13601 (N_13601,N_13487,N_13460);
xnor U13602 (N_13602,N_13574,N_13570);
xor U13603 (N_13603,N_13554,N_13476);
nand U13604 (N_13604,N_13513,N_13558);
xnor U13605 (N_13605,N_13511,N_13579);
xor U13606 (N_13606,N_13589,N_13446);
and U13607 (N_13607,N_13530,N_13447);
and U13608 (N_13608,N_13525,N_13539);
nand U13609 (N_13609,N_13596,N_13484);
nor U13610 (N_13610,N_13542,N_13466);
or U13611 (N_13611,N_13486,N_13546);
and U13612 (N_13612,N_13568,N_13537);
nand U13613 (N_13613,N_13523,N_13500);
xor U13614 (N_13614,N_13503,N_13505);
nor U13615 (N_13615,N_13441,N_13567);
or U13616 (N_13616,N_13473,N_13440);
or U13617 (N_13617,N_13527,N_13562);
nor U13618 (N_13618,N_13515,N_13518);
nor U13619 (N_13619,N_13470,N_13573);
nand U13620 (N_13620,N_13529,N_13526);
or U13621 (N_13621,N_13520,N_13496);
or U13622 (N_13622,N_13452,N_13492);
nor U13623 (N_13623,N_13549,N_13491);
nand U13624 (N_13624,N_13531,N_13591);
nor U13625 (N_13625,N_13533,N_13507);
or U13626 (N_13626,N_13444,N_13564);
nor U13627 (N_13627,N_13521,N_13458);
or U13628 (N_13628,N_13588,N_13584);
nor U13629 (N_13629,N_13581,N_13455);
nor U13630 (N_13630,N_13469,N_13553);
or U13631 (N_13631,N_13488,N_13597);
and U13632 (N_13632,N_13593,N_13467);
nand U13633 (N_13633,N_13454,N_13550);
nor U13634 (N_13634,N_13540,N_13595);
nor U13635 (N_13635,N_13572,N_13560);
nor U13636 (N_13636,N_13456,N_13544);
nand U13637 (N_13637,N_13543,N_13504);
xor U13638 (N_13638,N_13594,N_13590);
and U13639 (N_13639,N_13580,N_13453);
nor U13640 (N_13640,N_13555,N_13459);
and U13641 (N_13641,N_13463,N_13501);
nand U13642 (N_13642,N_13548,N_13517);
and U13643 (N_13643,N_13510,N_13485);
and U13644 (N_13644,N_13569,N_13516);
xnor U13645 (N_13645,N_13461,N_13443);
nor U13646 (N_13646,N_13475,N_13442);
and U13647 (N_13647,N_13448,N_13490);
nor U13648 (N_13648,N_13598,N_13534);
nand U13649 (N_13649,N_13499,N_13538);
xnor U13650 (N_13650,N_13577,N_13545);
xnor U13651 (N_13651,N_13583,N_13478);
nand U13652 (N_13652,N_13445,N_13509);
xnor U13653 (N_13653,N_13498,N_13462);
nor U13654 (N_13654,N_13582,N_13489);
and U13655 (N_13655,N_13502,N_13457);
or U13656 (N_13656,N_13541,N_13532);
nand U13657 (N_13657,N_13514,N_13468);
xor U13658 (N_13658,N_13585,N_13477);
nand U13659 (N_13659,N_13519,N_13493);
xor U13660 (N_13660,N_13565,N_13465);
nand U13661 (N_13661,N_13566,N_13480);
nor U13662 (N_13662,N_13559,N_13592);
nor U13663 (N_13663,N_13575,N_13451);
or U13664 (N_13664,N_13571,N_13464);
nand U13665 (N_13665,N_13512,N_13506);
nor U13666 (N_13666,N_13495,N_13536);
and U13667 (N_13667,N_13552,N_13450);
xor U13668 (N_13668,N_13535,N_13547);
and U13669 (N_13669,N_13578,N_13497);
nor U13670 (N_13670,N_13587,N_13528);
or U13671 (N_13671,N_13556,N_13563);
nand U13672 (N_13672,N_13474,N_13482);
nor U13673 (N_13673,N_13576,N_13586);
nand U13674 (N_13674,N_13449,N_13479);
nor U13675 (N_13675,N_13508,N_13481);
nor U13676 (N_13676,N_13494,N_13524);
and U13677 (N_13677,N_13561,N_13522);
nor U13678 (N_13678,N_13599,N_13471);
xor U13679 (N_13679,N_13551,N_13483);
nand U13680 (N_13680,N_13526,N_13547);
or U13681 (N_13681,N_13537,N_13527);
or U13682 (N_13682,N_13465,N_13486);
nand U13683 (N_13683,N_13529,N_13584);
nor U13684 (N_13684,N_13592,N_13570);
and U13685 (N_13685,N_13593,N_13496);
nor U13686 (N_13686,N_13513,N_13487);
nor U13687 (N_13687,N_13578,N_13544);
and U13688 (N_13688,N_13540,N_13495);
nand U13689 (N_13689,N_13478,N_13469);
nor U13690 (N_13690,N_13577,N_13495);
nand U13691 (N_13691,N_13442,N_13452);
xnor U13692 (N_13692,N_13535,N_13445);
or U13693 (N_13693,N_13513,N_13571);
nor U13694 (N_13694,N_13481,N_13553);
xor U13695 (N_13695,N_13551,N_13540);
and U13696 (N_13696,N_13595,N_13594);
xor U13697 (N_13697,N_13498,N_13508);
xnor U13698 (N_13698,N_13547,N_13574);
nor U13699 (N_13699,N_13461,N_13451);
or U13700 (N_13700,N_13480,N_13555);
and U13701 (N_13701,N_13528,N_13529);
nor U13702 (N_13702,N_13535,N_13552);
nor U13703 (N_13703,N_13535,N_13441);
xnor U13704 (N_13704,N_13455,N_13520);
nor U13705 (N_13705,N_13520,N_13457);
nor U13706 (N_13706,N_13477,N_13497);
xnor U13707 (N_13707,N_13515,N_13463);
nand U13708 (N_13708,N_13509,N_13543);
or U13709 (N_13709,N_13471,N_13523);
nand U13710 (N_13710,N_13530,N_13536);
xnor U13711 (N_13711,N_13491,N_13448);
nand U13712 (N_13712,N_13528,N_13586);
xnor U13713 (N_13713,N_13457,N_13515);
or U13714 (N_13714,N_13550,N_13566);
nor U13715 (N_13715,N_13520,N_13576);
nor U13716 (N_13716,N_13559,N_13555);
nand U13717 (N_13717,N_13537,N_13493);
or U13718 (N_13718,N_13463,N_13595);
xnor U13719 (N_13719,N_13449,N_13442);
nand U13720 (N_13720,N_13467,N_13536);
xor U13721 (N_13721,N_13443,N_13541);
xor U13722 (N_13722,N_13464,N_13599);
nor U13723 (N_13723,N_13562,N_13597);
or U13724 (N_13724,N_13533,N_13553);
and U13725 (N_13725,N_13454,N_13533);
xnor U13726 (N_13726,N_13484,N_13592);
xnor U13727 (N_13727,N_13515,N_13458);
nor U13728 (N_13728,N_13549,N_13464);
and U13729 (N_13729,N_13454,N_13599);
or U13730 (N_13730,N_13446,N_13554);
or U13731 (N_13731,N_13467,N_13490);
nand U13732 (N_13732,N_13541,N_13534);
xor U13733 (N_13733,N_13442,N_13532);
xnor U13734 (N_13734,N_13595,N_13553);
nand U13735 (N_13735,N_13449,N_13529);
nor U13736 (N_13736,N_13524,N_13539);
xor U13737 (N_13737,N_13513,N_13576);
xnor U13738 (N_13738,N_13582,N_13542);
nand U13739 (N_13739,N_13588,N_13447);
nand U13740 (N_13740,N_13594,N_13585);
and U13741 (N_13741,N_13482,N_13453);
and U13742 (N_13742,N_13589,N_13444);
xnor U13743 (N_13743,N_13598,N_13443);
and U13744 (N_13744,N_13558,N_13593);
xnor U13745 (N_13745,N_13488,N_13538);
and U13746 (N_13746,N_13549,N_13458);
nor U13747 (N_13747,N_13452,N_13487);
xor U13748 (N_13748,N_13552,N_13473);
nor U13749 (N_13749,N_13567,N_13513);
and U13750 (N_13750,N_13525,N_13499);
nor U13751 (N_13751,N_13551,N_13546);
xor U13752 (N_13752,N_13562,N_13578);
or U13753 (N_13753,N_13557,N_13546);
or U13754 (N_13754,N_13590,N_13453);
nand U13755 (N_13755,N_13593,N_13548);
nand U13756 (N_13756,N_13593,N_13533);
and U13757 (N_13757,N_13458,N_13498);
nand U13758 (N_13758,N_13549,N_13477);
and U13759 (N_13759,N_13584,N_13522);
nor U13760 (N_13760,N_13754,N_13742);
nand U13761 (N_13761,N_13613,N_13664);
nor U13762 (N_13762,N_13718,N_13612);
xor U13763 (N_13763,N_13731,N_13735);
or U13764 (N_13764,N_13693,N_13724);
nand U13765 (N_13765,N_13694,N_13601);
and U13766 (N_13766,N_13708,N_13745);
xor U13767 (N_13767,N_13753,N_13711);
nor U13768 (N_13768,N_13671,N_13669);
xor U13769 (N_13769,N_13659,N_13697);
nor U13770 (N_13770,N_13691,N_13704);
and U13771 (N_13771,N_13639,N_13679);
nor U13772 (N_13772,N_13692,N_13625);
nand U13773 (N_13773,N_13681,N_13651);
or U13774 (N_13774,N_13620,N_13732);
or U13775 (N_13775,N_13629,N_13725);
nand U13776 (N_13776,N_13636,N_13638);
or U13777 (N_13777,N_13728,N_13622);
nor U13778 (N_13778,N_13684,N_13686);
xor U13779 (N_13779,N_13600,N_13712);
and U13780 (N_13780,N_13676,N_13609);
and U13781 (N_13781,N_13617,N_13616);
or U13782 (N_13782,N_13663,N_13702);
nand U13783 (N_13783,N_13734,N_13740);
nor U13784 (N_13784,N_13757,N_13665);
nand U13785 (N_13785,N_13668,N_13689);
nor U13786 (N_13786,N_13751,N_13705);
or U13787 (N_13787,N_13759,N_13628);
nand U13788 (N_13788,N_13624,N_13614);
nor U13789 (N_13789,N_13647,N_13621);
nand U13790 (N_13790,N_13756,N_13634);
nor U13791 (N_13791,N_13632,N_13670);
xnor U13792 (N_13792,N_13645,N_13746);
xnor U13793 (N_13793,N_13618,N_13662);
xnor U13794 (N_13794,N_13606,N_13608);
or U13795 (N_13795,N_13737,N_13611);
nor U13796 (N_13796,N_13648,N_13680);
or U13797 (N_13797,N_13672,N_13747);
and U13798 (N_13798,N_13700,N_13619);
or U13799 (N_13799,N_13758,N_13690);
or U13800 (N_13800,N_13673,N_13605);
nor U13801 (N_13801,N_13643,N_13715);
nor U13802 (N_13802,N_13642,N_13710);
and U13803 (N_13803,N_13637,N_13666);
and U13804 (N_13804,N_13675,N_13739);
nor U13805 (N_13805,N_13703,N_13749);
or U13806 (N_13806,N_13730,N_13701);
nand U13807 (N_13807,N_13646,N_13709);
and U13808 (N_13808,N_13652,N_13743);
or U13809 (N_13809,N_13630,N_13657);
nor U13810 (N_13810,N_13744,N_13683);
nand U13811 (N_13811,N_13755,N_13723);
xor U13812 (N_13812,N_13626,N_13603);
or U13813 (N_13813,N_13696,N_13633);
or U13814 (N_13814,N_13748,N_13667);
and U13815 (N_13815,N_13733,N_13736);
nand U13816 (N_13816,N_13655,N_13698);
or U13817 (N_13817,N_13706,N_13654);
and U13818 (N_13818,N_13602,N_13658);
xor U13819 (N_13819,N_13641,N_13623);
xor U13820 (N_13820,N_13650,N_13615);
and U13821 (N_13821,N_13687,N_13682);
and U13822 (N_13822,N_13729,N_13678);
and U13823 (N_13823,N_13714,N_13750);
or U13824 (N_13824,N_13726,N_13677);
and U13825 (N_13825,N_13656,N_13644);
xor U13826 (N_13826,N_13631,N_13685);
nor U13827 (N_13827,N_13635,N_13721);
nor U13828 (N_13828,N_13738,N_13719);
xnor U13829 (N_13829,N_13699,N_13653);
nor U13830 (N_13830,N_13640,N_13727);
nand U13831 (N_13831,N_13604,N_13707);
xnor U13832 (N_13832,N_13688,N_13717);
and U13833 (N_13833,N_13722,N_13627);
or U13834 (N_13834,N_13674,N_13695);
or U13835 (N_13835,N_13713,N_13716);
and U13836 (N_13836,N_13752,N_13741);
nand U13837 (N_13837,N_13610,N_13649);
and U13838 (N_13838,N_13661,N_13720);
nor U13839 (N_13839,N_13660,N_13607);
and U13840 (N_13840,N_13642,N_13679);
and U13841 (N_13841,N_13621,N_13641);
and U13842 (N_13842,N_13698,N_13672);
nor U13843 (N_13843,N_13623,N_13737);
and U13844 (N_13844,N_13673,N_13677);
nand U13845 (N_13845,N_13742,N_13614);
or U13846 (N_13846,N_13701,N_13677);
and U13847 (N_13847,N_13738,N_13690);
or U13848 (N_13848,N_13691,N_13706);
or U13849 (N_13849,N_13736,N_13646);
and U13850 (N_13850,N_13759,N_13608);
nand U13851 (N_13851,N_13753,N_13627);
nand U13852 (N_13852,N_13679,N_13660);
nand U13853 (N_13853,N_13652,N_13744);
nand U13854 (N_13854,N_13725,N_13674);
nand U13855 (N_13855,N_13680,N_13624);
nor U13856 (N_13856,N_13630,N_13622);
or U13857 (N_13857,N_13607,N_13612);
xor U13858 (N_13858,N_13675,N_13686);
or U13859 (N_13859,N_13733,N_13750);
and U13860 (N_13860,N_13646,N_13699);
and U13861 (N_13861,N_13671,N_13689);
and U13862 (N_13862,N_13694,N_13659);
nand U13863 (N_13863,N_13629,N_13704);
and U13864 (N_13864,N_13696,N_13650);
nor U13865 (N_13865,N_13718,N_13698);
nor U13866 (N_13866,N_13735,N_13653);
nand U13867 (N_13867,N_13722,N_13633);
nor U13868 (N_13868,N_13746,N_13663);
xnor U13869 (N_13869,N_13740,N_13747);
nand U13870 (N_13870,N_13681,N_13720);
or U13871 (N_13871,N_13723,N_13674);
nor U13872 (N_13872,N_13726,N_13629);
xor U13873 (N_13873,N_13610,N_13632);
xor U13874 (N_13874,N_13628,N_13720);
xor U13875 (N_13875,N_13712,N_13757);
or U13876 (N_13876,N_13671,N_13617);
xnor U13877 (N_13877,N_13692,N_13629);
nand U13878 (N_13878,N_13720,N_13749);
xnor U13879 (N_13879,N_13721,N_13718);
nor U13880 (N_13880,N_13670,N_13758);
nand U13881 (N_13881,N_13684,N_13646);
nand U13882 (N_13882,N_13668,N_13670);
nor U13883 (N_13883,N_13600,N_13728);
and U13884 (N_13884,N_13641,N_13631);
or U13885 (N_13885,N_13714,N_13660);
nand U13886 (N_13886,N_13665,N_13715);
or U13887 (N_13887,N_13643,N_13681);
and U13888 (N_13888,N_13757,N_13660);
nand U13889 (N_13889,N_13659,N_13650);
and U13890 (N_13890,N_13610,N_13740);
xor U13891 (N_13891,N_13736,N_13703);
nand U13892 (N_13892,N_13688,N_13715);
xor U13893 (N_13893,N_13669,N_13621);
nor U13894 (N_13894,N_13644,N_13725);
nand U13895 (N_13895,N_13624,N_13749);
or U13896 (N_13896,N_13639,N_13660);
xor U13897 (N_13897,N_13734,N_13618);
nand U13898 (N_13898,N_13656,N_13693);
and U13899 (N_13899,N_13611,N_13749);
xor U13900 (N_13900,N_13639,N_13618);
and U13901 (N_13901,N_13664,N_13621);
nor U13902 (N_13902,N_13629,N_13663);
and U13903 (N_13903,N_13714,N_13685);
nand U13904 (N_13904,N_13628,N_13706);
and U13905 (N_13905,N_13634,N_13709);
or U13906 (N_13906,N_13655,N_13626);
and U13907 (N_13907,N_13611,N_13623);
or U13908 (N_13908,N_13693,N_13641);
xor U13909 (N_13909,N_13630,N_13670);
or U13910 (N_13910,N_13614,N_13705);
nor U13911 (N_13911,N_13637,N_13711);
and U13912 (N_13912,N_13612,N_13679);
nand U13913 (N_13913,N_13677,N_13612);
nor U13914 (N_13914,N_13677,N_13708);
nand U13915 (N_13915,N_13654,N_13636);
nand U13916 (N_13916,N_13663,N_13693);
nor U13917 (N_13917,N_13683,N_13721);
nor U13918 (N_13918,N_13620,N_13722);
nor U13919 (N_13919,N_13704,N_13722);
or U13920 (N_13920,N_13871,N_13831);
nand U13921 (N_13921,N_13767,N_13858);
nand U13922 (N_13922,N_13866,N_13789);
and U13923 (N_13923,N_13780,N_13888);
xor U13924 (N_13924,N_13797,N_13819);
or U13925 (N_13925,N_13850,N_13898);
xnor U13926 (N_13926,N_13828,N_13841);
xnor U13927 (N_13927,N_13835,N_13884);
xor U13928 (N_13928,N_13777,N_13769);
xor U13929 (N_13929,N_13790,N_13918);
and U13930 (N_13930,N_13906,N_13834);
and U13931 (N_13931,N_13861,N_13764);
nor U13932 (N_13932,N_13848,N_13879);
xor U13933 (N_13933,N_13904,N_13776);
nor U13934 (N_13934,N_13916,N_13771);
or U13935 (N_13935,N_13813,N_13839);
nor U13936 (N_13936,N_13811,N_13877);
or U13937 (N_13937,N_13791,N_13821);
nor U13938 (N_13938,N_13814,N_13915);
nand U13939 (N_13939,N_13863,N_13919);
or U13940 (N_13940,N_13912,N_13909);
nor U13941 (N_13941,N_13881,N_13775);
or U13942 (N_13942,N_13900,N_13862);
and U13943 (N_13943,N_13760,N_13762);
and U13944 (N_13944,N_13809,N_13860);
or U13945 (N_13945,N_13806,N_13823);
nor U13946 (N_13946,N_13840,N_13778);
nor U13947 (N_13947,N_13854,N_13893);
or U13948 (N_13948,N_13830,N_13901);
nor U13949 (N_13949,N_13903,N_13765);
or U13950 (N_13950,N_13820,N_13770);
xor U13951 (N_13951,N_13805,N_13827);
and U13952 (N_13952,N_13772,N_13895);
or U13953 (N_13953,N_13808,N_13875);
xor U13954 (N_13954,N_13886,N_13773);
nor U13955 (N_13955,N_13796,N_13817);
xnor U13956 (N_13956,N_13907,N_13781);
or U13957 (N_13957,N_13892,N_13917);
and U13958 (N_13958,N_13864,N_13846);
and U13959 (N_13959,N_13802,N_13774);
nand U13960 (N_13960,N_13761,N_13766);
xor U13961 (N_13961,N_13826,N_13807);
and U13962 (N_13962,N_13874,N_13889);
nor U13963 (N_13963,N_13891,N_13783);
nor U13964 (N_13964,N_13793,N_13832);
and U13965 (N_13965,N_13908,N_13782);
nand U13966 (N_13966,N_13800,N_13896);
or U13967 (N_13967,N_13798,N_13799);
and U13968 (N_13968,N_13868,N_13804);
nand U13969 (N_13969,N_13836,N_13882);
or U13970 (N_13970,N_13843,N_13837);
nand U13971 (N_13971,N_13902,N_13870);
and U13972 (N_13972,N_13810,N_13824);
xor U13973 (N_13973,N_13816,N_13853);
and U13974 (N_13974,N_13786,N_13851);
or U13975 (N_13975,N_13867,N_13818);
and U13976 (N_13976,N_13787,N_13897);
xnor U13977 (N_13977,N_13829,N_13887);
nor U13978 (N_13978,N_13803,N_13905);
nand U13979 (N_13979,N_13845,N_13815);
and U13980 (N_13980,N_13856,N_13801);
nor U13981 (N_13981,N_13873,N_13857);
or U13982 (N_13982,N_13869,N_13794);
or U13983 (N_13983,N_13913,N_13910);
xnor U13984 (N_13984,N_13876,N_13865);
nor U13985 (N_13985,N_13784,N_13822);
nor U13986 (N_13986,N_13890,N_13849);
xor U13987 (N_13987,N_13911,N_13825);
xnor U13988 (N_13988,N_13779,N_13833);
nand U13989 (N_13989,N_13792,N_13883);
nor U13990 (N_13990,N_13847,N_13788);
or U13991 (N_13991,N_13844,N_13812);
nand U13992 (N_13992,N_13763,N_13838);
nor U13993 (N_13993,N_13852,N_13785);
and U13994 (N_13994,N_13880,N_13894);
nor U13995 (N_13995,N_13795,N_13878);
and U13996 (N_13996,N_13859,N_13914);
nor U13997 (N_13997,N_13899,N_13842);
and U13998 (N_13998,N_13768,N_13872);
and U13999 (N_13999,N_13855,N_13885);
or U14000 (N_14000,N_13831,N_13812);
xor U14001 (N_14001,N_13762,N_13797);
nand U14002 (N_14002,N_13772,N_13764);
xor U14003 (N_14003,N_13914,N_13873);
xnor U14004 (N_14004,N_13806,N_13842);
or U14005 (N_14005,N_13804,N_13911);
or U14006 (N_14006,N_13833,N_13790);
nand U14007 (N_14007,N_13887,N_13866);
nor U14008 (N_14008,N_13811,N_13761);
nand U14009 (N_14009,N_13760,N_13766);
and U14010 (N_14010,N_13830,N_13823);
xor U14011 (N_14011,N_13820,N_13782);
and U14012 (N_14012,N_13800,N_13886);
xor U14013 (N_14013,N_13842,N_13809);
or U14014 (N_14014,N_13888,N_13864);
or U14015 (N_14015,N_13787,N_13775);
or U14016 (N_14016,N_13783,N_13795);
or U14017 (N_14017,N_13806,N_13811);
nand U14018 (N_14018,N_13881,N_13774);
xor U14019 (N_14019,N_13795,N_13907);
nor U14020 (N_14020,N_13919,N_13840);
or U14021 (N_14021,N_13910,N_13852);
xnor U14022 (N_14022,N_13872,N_13881);
and U14023 (N_14023,N_13761,N_13904);
and U14024 (N_14024,N_13817,N_13801);
and U14025 (N_14025,N_13878,N_13863);
xnor U14026 (N_14026,N_13910,N_13776);
xor U14027 (N_14027,N_13771,N_13792);
nor U14028 (N_14028,N_13777,N_13829);
nand U14029 (N_14029,N_13838,N_13791);
nand U14030 (N_14030,N_13796,N_13788);
or U14031 (N_14031,N_13804,N_13897);
and U14032 (N_14032,N_13873,N_13867);
nand U14033 (N_14033,N_13898,N_13889);
or U14034 (N_14034,N_13782,N_13777);
xor U14035 (N_14035,N_13910,N_13837);
nor U14036 (N_14036,N_13832,N_13773);
or U14037 (N_14037,N_13772,N_13900);
nand U14038 (N_14038,N_13821,N_13914);
xor U14039 (N_14039,N_13858,N_13840);
nand U14040 (N_14040,N_13917,N_13890);
xnor U14041 (N_14041,N_13831,N_13799);
nor U14042 (N_14042,N_13807,N_13811);
xnor U14043 (N_14043,N_13879,N_13876);
nor U14044 (N_14044,N_13810,N_13893);
nand U14045 (N_14045,N_13830,N_13773);
or U14046 (N_14046,N_13864,N_13861);
and U14047 (N_14047,N_13786,N_13848);
or U14048 (N_14048,N_13785,N_13874);
and U14049 (N_14049,N_13819,N_13867);
nor U14050 (N_14050,N_13899,N_13770);
nand U14051 (N_14051,N_13848,N_13850);
or U14052 (N_14052,N_13811,N_13884);
nor U14053 (N_14053,N_13793,N_13865);
nand U14054 (N_14054,N_13834,N_13825);
xor U14055 (N_14055,N_13838,N_13878);
nand U14056 (N_14056,N_13809,N_13858);
xnor U14057 (N_14057,N_13850,N_13770);
or U14058 (N_14058,N_13867,N_13849);
nand U14059 (N_14059,N_13839,N_13880);
and U14060 (N_14060,N_13854,N_13900);
xor U14061 (N_14061,N_13917,N_13885);
xnor U14062 (N_14062,N_13848,N_13824);
xnor U14063 (N_14063,N_13761,N_13771);
xor U14064 (N_14064,N_13762,N_13838);
xor U14065 (N_14065,N_13762,N_13859);
nor U14066 (N_14066,N_13869,N_13838);
xnor U14067 (N_14067,N_13902,N_13791);
and U14068 (N_14068,N_13822,N_13875);
and U14069 (N_14069,N_13843,N_13900);
or U14070 (N_14070,N_13802,N_13888);
nor U14071 (N_14071,N_13816,N_13786);
nor U14072 (N_14072,N_13884,N_13777);
or U14073 (N_14073,N_13807,N_13848);
nor U14074 (N_14074,N_13851,N_13902);
and U14075 (N_14075,N_13855,N_13905);
xor U14076 (N_14076,N_13885,N_13861);
and U14077 (N_14077,N_13887,N_13875);
nand U14078 (N_14078,N_13841,N_13814);
and U14079 (N_14079,N_13815,N_13786);
nand U14080 (N_14080,N_14073,N_13928);
and U14081 (N_14081,N_13976,N_13994);
nor U14082 (N_14082,N_14043,N_13935);
nand U14083 (N_14083,N_14074,N_13937);
or U14084 (N_14084,N_13997,N_14045);
nor U14085 (N_14085,N_13975,N_13924);
nand U14086 (N_14086,N_13946,N_14067);
nor U14087 (N_14087,N_13929,N_13970);
xor U14088 (N_14088,N_14078,N_14039);
or U14089 (N_14089,N_13932,N_13996);
xnor U14090 (N_14090,N_14020,N_13973);
or U14091 (N_14091,N_14075,N_13966);
xor U14092 (N_14092,N_14010,N_13955);
and U14093 (N_14093,N_13962,N_13980);
xnor U14094 (N_14094,N_13930,N_13977);
nand U14095 (N_14095,N_14018,N_13952);
or U14096 (N_14096,N_14031,N_14017);
nor U14097 (N_14097,N_13944,N_13957);
nor U14098 (N_14098,N_13931,N_14057);
xor U14099 (N_14099,N_13961,N_14042);
and U14100 (N_14100,N_14028,N_14059);
nand U14101 (N_14101,N_13983,N_14004);
nand U14102 (N_14102,N_14079,N_13923);
and U14103 (N_14103,N_13956,N_13942);
and U14104 (N_14104,N_14047,N_13941);
xnor U14105 (N_14105,N_13940,N_14063);
or U14106 (N_14106,N_14022,N_13948);
nand U14107 (N_14107,N_13934,N_13985);
nand U14108 (N_14108,N_13998,N_14014);
nor U14109 (N_14109,N_14000,N_13922);
nand U14110 (N_14110,N_14035,N_14055);
nand U14111 (N_14111,N_14015,N_14050);
or U14112 (N_14112,N_13993,N_14006);
and U14113 (N_14113,N_13921,N_14013);
nand U14114 (N_14114,N_14040,N_14009);
or U14115 (N_14115,N_14053,N_14054);
or U14116 (N_14116,N_13992,N_14016);
and U14117 (N_14117,N_13945,N_14048);
xor U14118 (N_14118,N_13965,N_14023);
or U14119 (N_14119,N_14038,N_13989);
xor U14120 (N_14120,N_13986,N_14066);
nor U14121 (N_14121,N_13947,N_13963);
or U14122 (N_14122,N_13999,N_13958);
or U14123 (N_14123,N_13972,N_13971);
nor U14124 (N_14124,N_14005,N_14011);
nor U14125 (N_14125,N_14007,N_14025);
and U14126 (N_14126,N_13995,N_13926);
or U14127 (N_14127,N_14036,N_14068);
nor U14128 (N_14128,N_13959,N_14056);
and U14129 (N_14129,N_14052,N_14046);
or U14130 (N_14130,N_14037,N_14041);
xor U14131 (N_14131,N_14062,N_13951);
nor U14132 (N_14132,N_14061,N_13968);
xnor U14133 (N_14133,N_14064,N_13927);
and U14134 (N_14134,N_13984,N_13990);
and U14135 (N_14135,N_14076,N_14002);
xnor U14136 (N_14136,N_14065,N_13967);
nand U14137 (N_14137,N_13988,N_13964);
or U14138 (N_14138,N_14001,N_14026);
nand U14139 (N_14139,N_14034,N_14030);
xnor U14140 (N_14140,N_14060,N_13950);
and U14141 (N_14141,N_13981,N_14027);
and U14142 (N_14142,N_13939,N_14021);
nand U14143 (N_14143,N_13991,N_14077);
and U14144 (N_14144,N_13974,N_14024);
nor U14145 (N_14145,N_13953,N_14029);
xnor U14146 (N_14146,N_14049,N_14069);
nor U14147 (N_14147,N_14032,N_14019);
xnor U14148 (N_14148,N_14012,N_13943);
nand U14149 (N_14149,N_13925,N_13979);
or U14150 (N_14150,N_14051,N_13954);
nand U14151 (N_14151,N_13920,N_14044);
xor U14152 (N_14152,N_14003,N_14033);
nand U14153 (N_14153,N_13987,N_14008);
nor U14154 (N_14154,N_13969,N_13978);
nor U14155 (N_14155,N_14071,N_13936);
and U14156 (N_14156,N_13938,N_13982);
xnor U14157 (N_14157,N_14072,N_14070);
nand U14158 (N_14158,N_14058,N_13949);
or U14159 (N_14159,N_13933,N_13960);
nor U14160 (N_14160,N_13967,N_13950);
xnor U14161 (N_14161,N_13982,N_14010);
or U14162 (N_14162,N_14009,N_14000);
xor U14163 (N_14163,N_14064,N_14051);
or U14164 (N_14164,N_14020,N_13939);
nor U14165 (N_14165,N_13942,N_13946);
or U14166 (N_14166,N_14061,N_14028);
nor U14167 (N_14167,N_14009,N_13952);
or U14168 (N_14168,N_13924,N_13996);
nor U14169 (N_14169,N_14060,N_14001);
or U14170 (N_14170,N_14066,N_14035);
or U14171 (N_14171,N_13978,N_13988);
and U14172 (N_14172,N_14042,N_14046);
or U14173 (N_14173,N_14026,N_13966);
nand U14174 (N_14174,N_13984,N_14027);
and U14175 (N_14175,N_13930,N_13938);
nand U14176 (N_14176,N_14035,N_14021);
nor U14177 (N_14177,N_14013,N_14015);
and U14178 (N_14178,N_13985,N_13963);
or U14179 (N_14179,N_14049,N_13926);
nor U14180 (N_14180,N_13929,N_13981);
or U14181 (N_14181,N_13949,N_14061);
nor U14182 (N_14182,N_14000,N_14011);
and U14183 (N_14183,N_14062,N_13991);
xor U14184 (N_14184,N_14071,N_14068);
nand U14185 (N_14185,N_13949,N_13974);
nor U14186 (N_14186,N_13997,N_13975);
and U14187 (N_14187,N_13982,N_14030);
or U14188 (N_14188,N_13955,N_14076);
or U14189 (N_14189,N_14025,N_14062);
nand U14190 (N_14190,N_13973,N_13983);
xnor U14191 (N_14191,N_13955,N_14030);
xnor U14192 (N_14192,N_13920,N_13930);
xor U14193 (N_14193,N_13974,N_14051);
xor U14194 (N_14194,N_13978,N_13981);
or U14195 (N_14195,N_14016,N_13980);
nand U14196 (N_14196,N_13962,N_14027);
nand U14197 (N_14197,N_13983,N_13921);
xor U14198 (N_14198,N_14059,N_14072);
nor U14199 (N_14199,N_14046,N_14029);
xnor U14200 (N_14200,N_14029,N_14013);
nor U14201 (N_14201,N_13979,N_14065);
nor U14202 (N_14202,N_14061,N_13964);
and U14203 (N_14203,N_13988,N_13979);
nor U14204 (N_14204,N_13933,N_14020);
and U14205 (N_14205,N_14034,N_13936);
nor U14206 (N_14206,N_13971,N_14056);
and U14207 (N_14207,N_14002,N_14008);
and U14208 (N_14208,N_14036,N_14064);
or U14209 (N_14209,N_13966,N_13938);
or U14210 (N_14210,N_13994,N_14056);
xnor U14211 (N_14211,N_13925,N_14074);
or U14212 (N_14212,N_14040,N_13999);
or U14213 (N_14213,N_14042,N_13927);
xnor U14214 (N_14214,N_13965,N_13964);
and U14215 (N_14215,N_13924,N_14034);
nand U14216 (N_14216,N_13923,N_14064);
xor U14217 (N_14217,N_14007,N_13987);
xnor U14218 (N_14218,N_13934,N_14024);
xnor U14219 (N_14219,N_14068,N_14053);
or U14220 (N_14220,N_13987,N_14061);
xnor U14221 (N_14221,N_13983,N_14009);
or U14222 (N_14222,N_14068,N_14039);
or U14223 (N_14223,N_14011,N_14016);
and U14224 (N_14224,N_13954,N_14016);
nand U14225 (N_14225,N_13978,N_13922);
nand U14226 (N_14226,N_13933,N_13975);
xor U14227 (N_14227,N_14063,N_14029);
nor U14228 (N_14228,N_13937,N_13965);
nand U14229 (N_14229,N_13925,N_13947);
nand U14230 (N_14230,N_14030,N_14052);
xnor U14231 (N_14231,N_14006,N_14036);
or U14232 (N_14232,N_14024,N_13941);
xnor U14233 (N_14233,N_13993,N_13922);
nor U14234 (N_14234,N_14072,N_13933);
nand U14235 (N_14235,N_14024,N_14005);
and U14236 (N_14236,N_13963,N_14009);
or U14237 (N_14237,N_14000,N_14046);
xnor U14238 (N_14238,N_13969,N_13951);
nand U14239 (N_14239,N_14053,N_13989);
or U14240 (N_14240,N_14134,N_14232);
nand U14241 (N_14241,N_14196,N_14168);
nor U14242 (N_14242,N_14195,N_14082);
or U14243 (N_14243,N_14111,N_14095);
or U14244 (N_14244,N_14083,N_14145);
and U14245 (N_14245,N_14157,N_14200);
nand U14246 (N_14246,N_14135,N_14189);
xnor U14247 (N_14247,N_14170,N_14147);
nand U14248 (N_14248,N_14178,N_14204);
xnor U14249 (N_14249,N_14085,N_14238);
nand U14250 (N_14250,N_14202,N_14117);
nor U14251 (N_14251,N_14152,N_14235);
or U14252 (N_14252,N_14151,N_14113);
and U14253 (N_14253,N_14153,N_14239);
and U14254 (N_14254,N_14123,N_14233);
or U14255 (N_14255,N_14190,N_14179);
and U14256 (N_14256,N_14108,N_14175);
nand U14257 (N_14257,N_14120,N_14119);
nand U14258 (N_14258,N_14087,N_14165);
or U14259 (N_14259,N_14208,N_14107);
nand U14260 (N_14260,N_14080,N_14229);
nand U14261 (N_14261,N_14209,N_14230);
nand U14262 (N_14262,N_14096,N_14173);
nor U14263 (N_14263,N_14102,N_14221);
or U14264 (N_14264,N_14187,N_14184);
nor U14265 (N_14265,N_14118,N_14142);
nor U14266 (N_14266,N_14207,N_14138);
xor U14267 (N_14267,N_14150,N_14216);
and U14268 (N_14268,N_14161,N_14234);
nand U14269 (N_14269,N_14163,N_14115);
or U14270 (N_14270,N_14226,N_14188);
xor U14271 (N_14271,N_14106,N_14218);
xnor U14272 (N_14272,N_14162,N_14127);
or U14273 (N_14273,N_14182,N_14211);
nand U14274 (N_14274,N_14220,N_14132);
or U14275 (N_14275,N_14144,N_14097);
xor U14276 (N_14276,N_14236,N_14213);
nor U14277 (N_14277,N_14169,N_14212);
or U14278 (N_14278,N_14104,N_14193);
or U14279 (N_14279,N_14136,N_14086);
and U14280 (N_14280,N_14146,N_14110);
nor U14281 (N_14281,N_14160,N_14126);
xor U14282 (N_14282,N_14092,N_14140);
or U14283 (N_14283,N_14181,N_14197);
or U14284 (N_14284,N_14094,N_14121);
xnor U14285 (N_14285,N_14210,N_14205);
nand U14286 (N_14286,N_14148,N_14093);
and U14287 (N_14287,N_14129,N_14105);
nor U14288 (N_14288,N_14214,N_14116);
nand U14289 (N_14289,N_14203,N_14201);
or U14290 (N_14290,N_14103,N_14098);
and U14291 (N_14291,N_14185,N_14176);
xor U14292 (N_14292,N_14177,N_14171);
and U14293 (N_14293,N_14128,N_14231);
nor U14294 (N_14294,N_14081,N_14137);
and U14295 (N_14295,N_14125,N_14124);
and U14296 (N_14296,N_14143,N_14198);
and U14297 (N_14297,N_14155,N_14167);
xnor U14298 (N_14298,N_14109,N_14133);
nand U14299 (N_14299,N_14217,N_14166);
xnor U14300 (N_14300,N_14219,N_14172);
nor U14301 (N_14301,N_14154,N_14141);
nor U14302 (N_14302,N_14237,N_14225);
or U14303 (N_14303,N_14101,N_14206);
nand U14304 (N_14304,N_14091,N_14130);
xor U14305 (N_14305,N_14149,N_14088);
xnor U14306 (N_14306,N_14139,N_14191);
nand U14307 (N_14307,N_14224,N_14089);
and U14308 (N_14308,N_14228,N_14215);
nor U14309 (N_14309,N_14099,N_14194);
nor U14310 (N_14310,N_14183,N_14174);
nor U14311 (N_14311,N_14112,N_14164);
xor U14312 (N_14312,N_14122,N_14199);
or U14313 (N_14313,N_14192,N_14159);
nor U14314 (N_14314,N_14156,N_14158);
nor U14315 (N_14315,N_14186,N_14223);
and U14316 (N_14316,N_14227,N_14180);
and U14317 (N_14317,N_14090,N_14084);
xnor U14318 (N_14318,N_14131,N_14222);
and U14319 (N_14319,N_14100,N_14114);
and U14320 (N_14320,N_14094,N_14110);
xnor U14321 (N_14321,N_14173,N_14190);
xor U14322 (N_14322,N_14217,N_14237);
xor U14323 (N_14323,N_14185,N_14101);
or U14324 (N_14324,N_14153,N_14225);
or U14325 (N_14325,N_14151,N_14144);
xnor U14326 (N_14326,N_14157,N_14165);
or U14327 (N_14327,N_14105,N_14108);
nand U14328 (N_14328,N_14180,N_14143);
nor U14329 (N_14329,N_14162,N_14117);
and U14330 (N_14330,N_14102,N_14233);
nor U14331 (N_14331,N_14139,N_14216);
and U14332 (N_14332,N_14176,N_14224);
nor U14333 (N_14333,N_14142,N_14185);
or U14334 (N_14334,N_14121,N_14191);
xnor U14335 (N_14335,N_14088,N_14100);
and U14336 (N_14336,N_14200,N_14212);
and U14337 (N_14337,N_14102,N_14134);
and U14338 (N_14338,N_14194,N_14136);
and U14339 (N_14339,N_14158,N_14238);
xnor U14340 (N_14340,N_14151,N_14163);
xor U14341 (N_14341,N_14181,N_14225);
nor U14342 (N_14342,N_14229,N_14090);
nand U14343 (N_14343,N_14205,N_14169);
nand U14344 (N_14344,N_14174,N_14173);
or U14345 (N_14345,N_14235,N_14184);
nand U14346 (N_14346,N_14159,N_14227);
or U14347 (N_14347,N_14171,N_14117);
nor U14348 (N_14348,N_14128,N_14164);
or U14349 (N_14349,N_14138,N_14088);
xnor U14350 (N_14350,N_14232,N_14220);
and U14351 (N_14351,N_14156,N_14091);
nor U14352 (N_14352,N_14165,N_14188);
xnor U14353 (N_14353,N_14128,N_14105);
nor U14354 (N_14354,N_14183,N_14123);
nor U14355 (N_14355,N_14216,N_14217);
nor U14356 (N_14356,N_14089,N_14202);
nand U14357 (N_14357,N_14099,N_14153);
xnor U14358 (N_14358,N_14143,N_14192);
and U14359 (N_14359,N_14090,N_14104);
nor U14360 (N_14360,N_14110,N_14183);
nor U14361 (N_14361,N_14141,N_14206);
or U14362 (N_14362,N_14132,N_14121);
nand U14363 (N_14363,N_14229,N_14213);
or U14364 (N_14364,N_14219,N_14224);
nor U14365 (N_14365,N_14153,N_14234);
and U14366 (N_14366,N_14111,N_14230);
nand U14367 (N_14367,N_14166,N_14175);
and U14368 (N_14368,N_14191,N_14176);
xnor U14369 (N_14369,N_14152,N_14088);
or U14370 (N_14370,N_14239,N_14233);
or U14371 (N_14371,N_14148,N_14173);
nand U14372 (N_14372,N_14182,N_14088);
xor U14373 (N_14373,N_14206,N_14238);
nor U14374 (N_14374,N_14170,N_14150);
nand U14375 (N_14375,N_14107,N_14224);
xor U14376 (N_14376,N_14180,N_14084);
and U14377 (N_14377,N_14201,N_14093);
xor U14378 (N_14378,N_14212,N_14236);
nand U14379 (N_14379,N_14224,N_14125);
or U14380 (N_14380,N_14080,N_14191);
or U14381 (N_14381,N_14191,N_14097);
nand U14382 (N_14382,N_14202,N_14193);
nor U14383 (N_14383,N_14171,N_14099);
or U14384 (N_14384,N_14149,N_14115);
xnor U14385 (N_14385,N_14165,N_14175);
or U14386 (N_14386,N_14110,N_14201);
nand U14387 (N_14387,N_14174,N_14135);
nor U14388 (N_14388,N_14111,N_14146);
or U14389 (N_14389,N_14089,N_14175);
and U14390 (N_14390,N_14124,N_14235);
xnor U14391 (N_14391,N_14189,N_14162);
and U14392 (N_14392,N_14189,N_14223);
or U14393 (N_14393,N_14234,N_14206);
or U14394 (N_14394,N_14174,N_14126);
nand U14395 (N_14395,N_14173,N_14129);
nand U14396 (N_14396,N_14158,N_14126);
and U14397 (N_14397,N_14209,N_14158);
and U14398 (N_14398,N_14186,N_14193);
and U14399 (N_14399,N_14234,N_14217);
nand U14400 (N_14400,N_14248,N_14268);
or U14401 (N_14401,N_14281,N_14319);
nand U14402 (N_14402,N_14359,N_14324);
and U14403 (N_14403,N_14394,N_14303);
xor U14404 (N_14404,N_14371,N_14310);
and U14405 (N_14405,N_14266,N_14337);
nor U14406 (N_14406,N_14399,N_14351);
or U14407 (N_14407,N_14253,N_14367);
nor U14408 (N_14408,N_14328,N_14308);
and U14409 (N_14409,N_14357,N_14270);
nor U14410 (N_14410,N_14372,N_14289);
and U14411 (N_14411,N_14369,N_14284);
and U14412 (N_14412,N_14314,N_14325);
or U14413 (N_14413,N_14356,N_14307);
nand U14414 (N_14414,N_14320,N_14260);
or U14415 (N_14415,N_14244,N_14298);
and U14416 (N_14416,N_14301,N_14304);
nor U14417 (N_14417,N_14322,N_14255);
nor U14418 (N_14418,N_14393,N_14327);
xnor U14419 (N_14419,N_14311,N_14353);
and U14420 (N_14420,N_14283,N_14395);
nor U14421 (N_14421,N_14291,N_14263);
xnor U14422 (N_14422,N_14276,N_14358);
xor U14423 (N_14423,N_14277,N_14398);
xnor U14424 (N_14424,N_14378,N_14347);
nor U14425 (N_14425,N_14247,N_14332);
and U14426 (N_14426,N_14317,N_14312);
xnor U14427 (N_14427,N_14384,N_14379);
xnor U14428 (N_14428,N_14350,N_14279);
nand U14429 (N_14429,N_14245,N_14302);
nor U14430 (N_14430,N_14355,N_14344);
nor U14431 (N_14431,N_14296,N_14264);
and U14432 (N_14432,N_14343,N_14316);
nor U14433 (N_14433,N_14315,N_14396);
nand U14434 (N_14434,N_14282,N_14240);
nand U14435 (N_14435,N_14365,N_14286);
or U14436 (N_14436,N_14330,N_14287);
nor U14437 (N_14437,N_14364,N_14313);
and U14438 (N_14438,N_14285,N_14243);
xor U14439 (N_14439,N_14380,N_14335);
or U14440 (N_14440,N_14388,N_14256);
nor U14441 (N_14441,N_14254,N_14377);
and U14442 (N_14442,N_14251,N_14370);
nor U14443 (N_14443,N_14274,N_14373);
or U14444 (N_14444,N_14306,N_14368);
or U14445 (N_14445,N_14374,N_14280);
and U14446 (N_14446,N_14389,N_14293);
or U14447 (N_14447,N_14339,N_14326);
xnor U14448 (N_14448,N_14262,N_14288);
nor U14449 (N_14449,N_14329,N_14261);
nor U14450 (N_14450,N_14382,N_14361);
or U14451 (N_14451,N_14341,N_14375);
xnor U14452 (N_14452,N_14295,N_14352);
nor U14453 (N_14453,N_14331,N_14290);
and U14454 (N_14454,N_14267,N_14349);
xnor U14455 (N_14455,N_14257,N_14340);
xor U14456 (N_14456,N_14269,N_14242);
nor U14457 (N_14457,N_14249,N_14292);
or U14458 (N_14458,N_14246,N_14354);
and U14459 (N_14459,N_14300,N_14278);
xor U14460 (N_14460,N_14318,N_14386);
nor U14461 (N_14461,N_14250,N_14334);
xor U14462 (N_14462,N_14381,N_14392);
and U14463 (N_14463,N_14383,N_14252);
nand U14464 (N_14464,N_14342,N_14362);
xnor U14465 (N_14465,N_14271,N_14385);
xor U14466 (N_14466,N_14391,N_14309);
or U14467 (N_14467,N_14363,N_14390);
or U14468 (N_14468,N_14294,N_14333);
nand U14469 (N_14469,N_14387,N_14323);
nand U14470 (N_14470,N_14336,N_14297);
and U14471 (N_14471,N_14321,N_14259);
nand U14472 (N_14472,N_14275,N_14345);
nor U14473 (N_14473,N_14241,N_14346);
nor U14474 (N_14474,N_14366,N_14338);
or U14475 (N_14475,N_14376,N_14348);
nor U14476 (N_14476,N_14272,N_14258);
nand U14477 (N_14477,N_14265,N_14273);
nand U14478 (N_14478,N_14305,N_14360);
nand U14479 (N_14479,N_14397,N_14299);
nand U14480 (N_14480,N_14387,N_14249);
or U14481 (N_14481,N_14271,N_14353);
nand U14482 (N_14482,N_14331,N_14394);
nor U14483 (N_14483,N_14377,N_14399);
nand U14484 (N_14484,N_14315,N_14312);
xor U14485 (N_14485,N_14355,N_14349);
xnor U14486 (N_14486,N_14326,N_14360);
xor U14487 (N_14487,N_14368,N_14331);
or U14488 (N_14488,N_14380,N_14342);
and U14489 (N_14489,N_14314,N_14252);
or U14490 (N_14490,N_14381,N_14299);
or U14491 (N_14491,N_14339,N_14267);
nor U14492 (N_14492,N_14304,N_14256);
or U14493 (N_14493,N_14366,N_14264);
or U14494 (N_14494,N_14258,N_14301);
or U14495 (N_14495,N_14295,N_14313);
and U14496 (N_14496,N_14315,N_14368);
nand U14497 (N_14497,N_14344,N_14354);
and U14498 (N_14498,N_14354,N_14296);
xor U14499 (N_14499,N_14373,N_14251);
and U14500 (N_14500,N_14332,N_14361);
or U14501 (N_14501,N_14354,N_14384);
xor U14502 (N_14502,N_14291,N_14372);
or U14503 (N_14503,N_14283,N_14340);
or U14504 (N_14504,N_14346,N_14345);
nor U14505 (N_14505,N_14350,N_14353);
or U14506 (N_14506,N_14341,N_14396);
xor U14507 (N_14507,N_14270,N_14382);
nand U14508 (N_14508,N_14376,N_14244);
xnor U14509 (N_14509,N_14271,N_14297);
xnor U14510 (N_14510,N_14336,N_14391);
nand U14511 (N_14511,N_14361,N_14378);
nor U14512 (N_14512,N_14253,N_14300);
nor U14513 (N_14513,N_14395,N_14253);
or U14514 (N_14514,N_14244,N_14347);
or U14515 (N_14515,N_14295,N_14332);
xor U14516 (N_14516,N_14353,N_14363);
xnor U14517 (N_14517,N_14292,N_14351);
or U14518 (N_14518,N_14266,N_14329);
nor U14519 (N_14519,N_14333,N_14357);
xor U14520 (N_14520,N_14325,N_14281);
and U14521 (N_14521,N_14336,N_14291);
or U14522 (N_14522,N_14317,N_14325);
nand U14523 (N_14523,N_14381,N_14397);
and U14524 (N_14524,N_14389,N_14340);
and U14525 (N_14525,N_14399,N_14314);
xnor U14526 (N_14526,N_14295,N_14328);
nand U14527 (N_14527,N_14359,N_14339);
xor U14528 (N_14528,N_14368,N_14302);
nand U14529 (N_14529,N_14365,N_14326);
or U14530 (N_14530,N_14266,N_14376);
or U14531 (N_14531,N_14342,N_14389);
or U14532 (N_14532,N_14256,N_14387);
nor U14533 (N_14533,N_14316,N_14368);
xor U14534 (N_14534,N_14255,N_14258);
xor U14535 (N_14535,N_14308,N_14296);
nand U14536 (N_14536,N_14293,N_14255);
and U14537 (N_14537,N_14392,N_14247);
and U14538 (N_14538,N_14355,N_14372);
nor U14539 (N_14539,N_14260,N_14251);
xnor U14540 (N_14540,N_14271,N_14298);
nand U14541 (N_14541,N_14274,N_14350);
and U14542 (N_14542,N_14241,N_14254);
and U14543 (N_14543,N_14251,N_14308);
xor U14544 (N_14544,N_14337,N_14255);
and U14545 (N_14545,N_14306,N_14387);
or U14546 (N_14546,N_14289,N_14299);
nand U14547 (N_14547,N_14292,N_14336);
and U14548 (N_14548,N_14247,N_14248);
or U14549 (N_14549,N_14322,N_14374);
nand U14550 (N_14550,N_14295,N_14370);
or U14551 (N_14551,N_14276,N_14279);
or U14552 (N_14552,N_14242,N_14251);
and U14553 (N_14553,N_14307,N_14296);
nand U14554 (N_14554,N_14320,N_14334);
xnor U14555 (N_14555,N_14278,N_14302);
xor U14556 (N_14556,N_14296,N_14397);
and U14557 (N_14557,N_14255,N_14298);
and U14558 (N_14558,N_14258,N_14359);
nand U14559 (N_14559,N_14276,N_14354);
xnor U14560 (N_14560,N_14437,N_14528);
nor U14561 (N_14561,N_14534,N_14429);
xor U14562 (N_14562,N_14443,N_14460);
or U14563 (N_14563,N_14522,N_14499);
and U14564 (N_14564,N_14488,N_14537);
nor U14565 (N_14565,N_14521,N_14517);
nor U14566 (N_14566,N_14549,N_14494);
nor U14567 (N_14567,N_14472,N_14445);
or U14568 (N_14568,N_14553,N_14531);
and U14569 (N_14569,N_14456,N_14506);
nand U14570 (N_14570,N_14431,N_14420);
and U14571 (N_14571,N_14471,N_14547);
xor U14572 (N_14572,N_14473,N_14515);
nand U14573 (N_14573,N_14479,N_14539);
nor U14574 (N_14574,N_14450,N_14412);
and U14575 (N_14575,N_14465,N_14435);
and U14576 (N_14576,N_14557,N_14438);
and U14577 (N_14577,N_14482,N_14533);
nand U14578 (N_14578,N_14426,N_14463);
xnor U14579 (N_14579,N_14470,N_14469);
and U14580 (N_14580,N_14486,N_14483);
nor U14581 (N_14581,N_14406,N_14434);
or U14582 (N_14582,N_14502,N_14449);
and U14583 (N_14583,N_14492,N_14436);
and U14584 (N_14584,N_14545,N_14540);
nor U14585 (N_14585,N_14461,N_14458);
xor U14586 (N_14586,N_14511,N_14548);
nand U14587 (N_14587,N_14414,N_14505);
xnor U14588 (N_14588,N_14466,N_14452);
or U14589 (N_14589,N_14446,N_14524);
xor U14590 (N_14590,N_14556,N_14468);
or U14591 (N_14591,N_14459,N_14497);
or U14592 (N_14592,N_14493,N_14491);
and U14593 (N_14593,N_14447,N_14529);
nor U14594 (N_14594,N_14417,N_14418);
nor U14595 (N_14595,N_14419,N_14409);
or U14596 (N_14596,N_14512,N_14507);
and U14597 (N_14597,N_14421,N_14451);
nand U14598 (N_14598,N_14541,N_14489);
or U14599 (N_14599,N_14474,N_14519);
xnor U14600 (N_14600,N_14530,N_14425);
or U14601 (N_14601,N_14480,N_14427);
nor U14602 (N_14602,N_14424,N_14495);
nor U14603 (N_14603,N_14416,N_14513);
xor U14604 (N_14604,N_14516,N_14485);
and U14605 (N_14605,N_14487,N_14501);
and U14606 (N_14606,N_14546,N_14440);
xor U14607 (N_14607,N_14527,N_14496);
nor U14608 (N_14608,N_14476,N_14430);
or U14609 (N_14609,N_14413,N_14478);
nor U14610 (N_14610,N_14520,N_14518);
nand U14611 (N_14611,N_14404,N_14441);
and U14612 (N_14612,N_14525,N_14464);
nand U14613 (N_14613,N_14535,N_14544);
and U14614 (N_14614,N_14455,N_14402);
or U14615 (N_14615,N_14442,N_14538);
xnor U14616 (N_14616,N_14554,N_14400);
nor U14617 (N_14617,N_14509,N_14523);
and U14618 (N_14618,N_14510,N_14432);
and U14619 (N_14619,N_14462,N_14558);
and U14620 (N_14620,N_14405,N_14526);
xor U14621 (N_14621,N_14552,N_14433);
nand U14622 (N_14622,N_14508,N_14428);
nand U14623 (N_14623,N_14423,N_14551);
and U14624 (N_14624,N_14408,N_14444);
or U14625 (N_14625,N_14504,N_14481);
or U14626 (N_14626,N_14498,N_14457);
nor U14627 (N_14627,N_14422,N_14477);
xor U14628 (N_14628,N_14467,N_14559);
xnor U14629 (N_14629,N_14415,N_14401);
and U14630 (N_14630,N_14542,N_14503);
xor U14631 (N_14631,N_14410,N_14555);
or U14632 (N_14632,N_14407,N_14411);
xor U14633 (N_14633,N_14550,N_14454);
and U14634 (N_14634,N_14543,N_14484);
and U14635 (N_14635,N_14532,N_14536);
nor U14636 (N_14636,N_14448,N_14403);
nand U14637 (N_14637,N_14490,N_14500);
nor U14638 (N_14638,N_14514,N_14453);
and U14639 (N_14639,N_14475,N_14439);
and U14640 (N_14640,N_14559,N_14430);
or U14641 (N_14641,N_14408,N_14503);
nor U14642 (N_14642,N_14451,N_14552);
and U14643 (N_14643,N_14401,N_14556);
nor U14644 (N_14644,N_14550,N_14448);
xnor U14645 (N_14645,N_14508,N_14511);
xor U14646 (N_14646,N_14478,N_14531);
nor U14647 (N_14647,N_14429,N_14490);
xor U14648 (N_14648,N_14428,N_14407);
or U14649 (N_14649,N_14547,N_14531);
nand U14650 (N_14650,N_14524,N_14416);
and U14651 (N_14651,N_14545,N_14474);
nor U14652 (N_14652,N_14437,N_14523);
nor U14653 (N_14653,N_14487,N_14457);
nor U14654 (N_14654,N_14484,N_14417);
and U14655 (N_14655,N_14552,N_14558);
xnor U14656 (N_14656,N_14506,N_14534);
and U14657 (N_14657,N_14531,N_14539);
or U14658 (N_14658,N_14429,N_14401);
or U14659 (N_14659,N_14555,N_14473);
or U14660 (N_14660,N_14405,N_14432);
nand U14661 (N_14661,N_14504,N_14521);
nand U14662 (N_14662,N_14456,N_14544);
nor U14663 (N_14663,N_14469,N_14502);
xor U14664 (N_14664,N_14453,N_14542);
nand U14665 (N_14665,N_14520,N_14442);
xor U14666 (N_14666,N_14468,N_14498);
and U14667 (N_14667,N_14539,N_14559);
xor U14668 (N_14668,N_14479,N_14544);
xnor U14669 (N_14669,N_14485,N_14437);
xor U14670 (N_14670,N_14479,N_14414);
or U14671 (N_14671,N_14411,N_14496);
nand U14672 (N_14672,N_14470,N_14487);
nor U14673 (N_14673,N_14445,N_14414);
nand U14674 (N_14674,N_14455,N_14496);
and U14675 (N_14675,N_14508,N_14433);
or U14676 (N_14676,N_14505,N_14451);
nor U14677 (N_14677,N_14559,N_14525);
and U14678 (N_14678,N_14484,N_14463);
nand U14679 (N_14679,N_14518,N_14465);
xnor U14680 (N_14680,N_14428,N_14544);
or U14681 (N_14681,N_14417,N_14416);
or U14682 (N_14682,N_14547,N_14477);
and U14683 (N_14683,N_14428,N_14470);
nand U14684 (N_14684,N_14458,N_14401);
nor U14685 (N_14685,N_14413,N_14546);
nor U14686 (N_14686,N_14547,N_14516);
nor U14687 (N_14687,N_14537,N_14431);
and U14688 (N_14688,N_14448,N_14489);
nand U14689 (N_14689,N_14516,N_14440);
xor U14690 (N_14690,N_14498,N_14420);
and U14691 (N_14691,N_14525,N_14422);
nor U14692 (N_14692,N_14518,N_14400);
xnor U14693 (N_14693,N_14500,N_14548);
xor U14694 (N_14694,N_14472,N_14455);
xnor U14695 (N_14695,N_14527,N_14521);
nand U14696 (N_14696,N_14439,N_14555);
or U14697 (N_14697,N_14550,N_14400);
or U14698 (N_14698,N_14449,N_14526);
xor U14699 (N_14699,N_14406,N_14516);
and U14700 (N_14700,N_14427,N_14552);
or U14701 (N_14701,N_14538,N_14476);
nor U14702 (N_14702,N_14497,N_14406);
and U14703 (N_14703,N_14417,N_14489);
and U14704 (N_14704,N_14551,N_14484);
or U14705 (N_14705,N_14499,N_14542);
nor U14706 (N_14706,N_14487,N_14520);
nand U14707 (N_14707,N_14463,N_14417);
and U14708 (N_14708,N_14547,N_14474);
nand U14709 (N_14709,N_14509,N_14553);
nor U14710 (N_14710,N_14556,N_14482);
or U14711 (N_14711,N_14498,N_14462);
nor U14712 (N_14712,N_14556,N_14483);
or U14713 (N_14713,N_14479,N_14542);
or U14714 (N_14714,N_14521,N_14530);
and U14715 (N_14715,N_14453,N_14428);
xor U14716 (N_14716,N_14488,N_14453);
nor U14717 (N_14717,N_14432,N_14498);
nor U14718 (N_14718,N_14452,N_14516);
and U14719 (N_14719,N_14400,N_14417);
nand U14720 (N_14720,N_14618,N_14682);
nand U14721 (N_14721,N_14661,N_14598);
nand U14722 (N_14722,N_14631,N_14589);
nor U14723 (N_14723,N_14691,N_14652);
and U14724 (N_14724,N_14625,N_14635);
or U14725 (N_14725,N_14580,N_14595);
and U14726 (N_14726,N_14610,N_14612);
nor U14727 (N_14727,N_14583,N_14639);
and U14728 (N_14728,N_14699,N_14719);
or U14729 (N_14729,N_14672,N_14692);
xor U14730 (N_14730,N_14627,N_14611);
xor U14731 (N_14731,N_14659,N_14614);
nor U14732 (N_14732,N_14696,N_14591);
and U14733 (N_14733,N_14597,N_14686);
xnor U14734 (N_14734,N_14667,N_14579);
or U14735 (N_14735,N_14703,N_14712);
xnor U14736 (N_14736,N_14657,N_14702);
nand U14737 (N_14737,N_14670,N_14704);
or U14738 (N_14738,N_14687,N_14594);
or U14739 (N_14739,N_14706,N_14633);
or U14740 (N_14740,N_14565,N_14563);
nand U14741 (N_14741,N_14684,N_14584);
nand U14742 (N_14742,N_14619,N_14574);
and U14743 (N_14743,N_14650,N_14573);
and U14744 (N_14744,N_14694,N_14567);
nor U14745 (N_14745,N_14581,N_14665);
xor U14746 (N_14746,N_14616,N_14596);
and U14747 (N_14747,N_14623,N_14713);
nand U14748 (N_14748,N_14577,N_14601);
nand U14749 (N_14749,N_14576,N_14709);
and U14750 (N_14750,N_14700,N_14561);
and U14751 (N_14751,N_14675,N_14679);
xor U14752 (N_14752,N_14648,N_14641);
nor U14753 (N_14753,N_14562,N_14697);
nand U14754 (N_14754,N_14599,N_14617);
or U14755 (N_14755,N_14683,N_14643);
xor U14756 (N_14756,N_14621,N_14717);
nor U14757 (N_14757,N_14572,N_14585);
or U14758 (N_14758,N_14613,N_14628);
xor U14759 (N_14759,N_14707,N_14678);
xnor U14760 (N_14760,N_14673,N_14708);
xnor U14761 (N_14761,N_14658,N_14630);
nor U14762 (N_14762,N_14588,N_14666);
nand U14763 (N_14763,N_14676,N_14660);
nand U14764 (N_14764,N_14566,N_14681);
or U14765 (N_14765,N_14671,N_14693);
xnor U14766 (N_14766,N_14622,N_14626);
or U14767 (N_14767,N_14677,N_14674);
or U14768 (N_14768,N_14647,N_14632);
xor U14769 (N_14769,N_14656,N_14638);
nand U14770 (N_14770,N_14602,N_14690);
or U14771 (N_14771,N_14571,N_14695);
or U14772 (N_14772,N_14560,N_14649);
or U14773 (N_14773,N_14592,N_14705);
nor U14774 (N_14774,N_14620,N_14698);
or U14775 (N_14775,N_14609,N_14570);
xor U14776 (N_14776,N_14604,N_14606);
nor U14777 (N_14777,N_14608,N_14685);
or U14778 (N_14778,N_14624,N_14607);
nand U14779 (N_14779,N_14600,N_14637);
xor U14780 (N_14780,N_14710,N_14629);
nand U14781 (N_14781,N_14568,N_14714);
nand U14782 (N_14782,N_14593,N_14662);
and U14783 (N_14783,N_14689,N_14615);
or U14784 (N_14784,N_14664,N_14701);
and U14785 (N_14785,N_14645,N_14634);
nor U14786 (N_14786,N_14718,N_14640);
or U14787 (N_14787,N_14646,N_14582);
or U14788 (N_14788,N_14603,N_14669);
or U14789 (N_14789,N_14586,N_14636);
xor U14790 (N_14790,N_14575,N_14587);
xnor U14791 (N_14791,N_14564,N_14688);
nand U14792 (N_14792,N_14680,N_14578);
xnor U14793 (N_14793,N_14590,N_14651);
and U14794 (N_14794,N_14716,N_14642);
nand U14795 (N_14795,N_14605,N_14715);
nand U14796 (N_14796,N_14654,N_14569);
and U14797 (N_14797,N_14644,N_14655);
nor U14798 (N_14798,N_14668,N_14653);
or U14799 (N_14799,N_14711,N_14663);
nand U14800 (N_14800,N_14566,N_14580);
or U14801 (N_14801,N_14709,N_14674);
nand U14802 (N_14802,N_14646,N_14689);
and U14803 (N_14803,N_14716,N_14629);
or U14804 (N_14804,N_14657,N_14638);
nor U14805 (N_14805,N_14695,N_14567);
nand U14806 (N_14806,N_14617,N_14608);
or U14807 (N_14807,N_14697,N_14568);
xnor U14808 (N_14808,N_14602,N_14709);
and U14809 (N_14809,N_14622,N_14662);
xnor U14810 (N_14810,N_14584,N_14629);
or U14811 (N_14811,N_14623,N_14566);
or U14812 (N_14812,N_14589,N_14609);
xnor U14813 (N_14813,N_14678,N_14708);
nor U14814 (N_14814,N_14603,N_14641);
or U14815 (N_14815,N_14562,N_14609);
xnor U14816 (N_14816,N_14583,N_14703);
or U14817 (N_14817,N_14690,N_14676);
and U14818 (N_14818,N_14701,N_14637);
nor U14819 (N_14819,N_14696,N_14686);
nand U14820 (N_14820,N_14583,N_14625);
nand U14821 (N_14821,N_14653,N_14642);
and U14822 (N_14822,N_14635,N_14660);
nand U14823 (N_14823,N_14560,N_14700);
xnor U14824 (N_14824,N_14702,N_14607);
nor U14825 (N_14825,N_14634,N_14567);
or U14826 (N_14826,N_14622,N_14678);
or U14827 (N_14827,N_14652,N_14644);
and U14828 (N_14828,N_14599,N_14675);
nor U14829 (N_14829,N_14655,N_14706);
xnor U14830 (N_14830,N_14626,N_14693);
xor U14831 (N_14831,N_14641,N_14650);
or U14832 (N_14832,N_14611,N_14642);
or U14833 (N_14833,N_14650,N_14705);
and U14834 (N_14834,N_14655,N_14635);
nor U14835 (N_14835,N_14614,N_14712);
nand U14836 (N_14836,N_14645,N_14561);
nand U14837 (N_14837,N_14599,N_14696);
xor U14838 (N_14838,N_14601,N_14634);
and U14839 (N_14839,N_14618,N_14580);
nand U14840 (N_14840,N_14617,N_14596);
nor U14841 (N_14841,N_14606,N_14649);
xor U14842 (N_14842,N_14563,N_14701);
and U14843 (N_14843,N_14560,N_14695);
and U14844 (N_14844,N_14670,N_14613);
nand U14845 (N_14845,N_14623,N_14683);
xor U14846 (N_14846,N_14714,N_14583);
or U14847 (N_14847,N_14619,N_14652);
and U14848 (N_14848,N_14590,N_14688);
and U14849 (N_14849,N_14596,N_14698);
nand U14850 (N_14850,N_14710,N_14678);
nor U14851 (N_14851,N_14688,N_14611);
xor U14852 (N_14852,N_14712,N_14711);
and U14853 (N_14853,N_14714,N_14567);
and U14854 (N_14854,N_14670,N_14594);
nand U14855 (N_14855,N_14582,N_14605);
xnor U14856 (N_14856,N_14652,N_14623);
and U14857 (N_14857,N_14589,N_14581);
xnor U14858 (N_14858,N_14637,N_14693);
nand U14859 (N_14859,N_14610,N_14673);
nand U14860 (N_14860,N_14666,N_14705);
or U14861 (N_14861,N_14587,N_14688);
nand U14862 (N_14862,N_14691,N_14688);
nand U14863 (N_14863,N_14599,N_14699);
xor U14864 (N_14864,N_14630,N_14671);
nand U14865 (N_14865,N_14694,N_14584);
or U14866 (N_14866,N_14650,N_14616);
and U14867 (N_14867,N_14606,N_14656);
nand U14868 (N_14868,N_14683,N_14695);
or U14869 (N_14869,N_14611,N_14718);
and U14870 (N_14870,N_14694,N_14699);
or U14871 (N_14871,N_14699,N_14614);
xor U14872 (N_14872,N_14627,N_14689);
xor U14873 (N_14873,N_14664,N_14692);
or U14874 (N_14874,N_14604,N_14677);
or U14875 (N_14875,N_14640,N_14564);
xor U14876 (N_14876,N_14569,N_14640);
or U14877 (N_14877,N_14716,N_14661);
and U14878 (N_14878,N_14663,N_14690);
nor U14879 (N_14879,N_14612,N_14708);
nor U14880 (N_14880,N_14747,N_14756);
or U14881 (N_14881,N_14778,N_14846);
and U14882 (N_14882,N_14808,N_14814);
nand U14883 (N_14883,N_14853,N_14727);
xor U14884 (N_14884,N_14771,N_14779);
nor U14885 (N_14885,N_14734,N_14872);
and U14886 (N_14886,N_14757,N_14720);
and U14887 (N_14887,N_14875,N_14824);
and U14888 (N_14888,N_14789,N_14791);
and U14889 (N_14889,N_14800,N_14744);
or U14890 (N_14890,N_14837,N_14838);
xor U14891 (N_14891,N_14855,N_14749);
nor U14892 (N_14892,N_14806,N_14769);
or U14893 (N_14893,N_14879,N_14842);
nand U14894 (N_14894,N_14748,N_14722);
or U14895 (N_14895,N_14728,N_14863);
nor U14896 (N_14896,N_14840,N_14750);
nor U14897 (N_14897,N_14774,N_14831);
and U14898 (N_14898,N_14792,N_14841);
nand U14899 (N_14899,N_14746,N_14821);
xnor U14900 (N_14900,N_14738,N_14819);
nand U14901 (N_14901,N_14844,N_14876);
or U14902 (N_14902,N_14767,N_14812);
and U14903 (N_14903,N_14764,N_14724);
nor U14904 (N_14904,N_14850,N_14818);
xnor U14905 (N_14905,N_14730,N_14828);
and U14906 (N_14906,N_14836,N_14768);
nor U14907 (N_14907,N_14760,N_14731);
and U14908 (N_14908,N_14732,N_14856);
nand U14909 (N_14909,N_14758,N_14874);
nand U14910 (N_14910,N_14823,N_14801);
nand U14911 (N_14911,N_14809,N_14795);
nand U14912 (N_14912,N_14833,N_14857);
nor U14913 (N_14913,N_14725,N_14737);
or U14914 (N_14914,N_14770,N_14766);
and U14915 (N_14915,N_14829,N_14762);
nand U14916 (N_14916,N_14805,N_14733);
and U14917 (N_14917,N_14786,N_14854);
or U14918 (N_14918,N_14765,N_14753);
and U14919 (N_14919,N_14761,N_14807);
nor U14920 (N_14920,N_14845,N_14743);
and U14921 (N_14921,N_14729,N_14859);
and U14922 (N_14922,N_14803,N_14825);
xnor U14923 (N_14923,N_14866,N_14736);
xnor U14924 (N_14924,N_14864,N_14861);
nor U14925 (N_14925,N_14775,N_14868);
nand U14926 (N_14926,N_14759,N_14869);
or U14927 (N_14927,N_14735,N_14843);
nor U14928 (N_14928,N_14790,N_14848);
nor U14929 (N_14929,N_14755,N_14788);
nor U14930 (N_14930,N_14742,N_14751);
nand U14931 (N_14931,N_14797,N_14820);
or U14932 (N_14932,N_14787,N_14810);
and U14933 (N_14933,N_14798,N_14860);
xnor U14934 (N_14934,N_14781,N_14816);
and U14935 (N_14935,N_14776,N_14785);
and U14936 (N_14936,N_14858,N_14871);
nor U14937 (N_14937,N_14754,N_14822);
and U14938 (N_14938,N_14721,N_14782);
nor U14939 (N_14939,N_14784,N_14867);
and U14940 (N_14940,N_14804,N_14847);
nand U14941 (N_14941,N_14794,N_14827);
or U14942 (N_14942,N_14826,N_14878);
or U14943 (N_14943,N_14723,N_14745);
nor U14944 (N_14944,N_14739,N_14852);
xor U14945 (N_14945,N_14870,N_14783);
and U14946 (N_14946,N_14811,N_14865);
xnor U14947 (N_14947,N_14726,N_14796);
or U14948 (N_14948,N_14839,N_14862);
xnor U14949 (N_14949,N_14777,N_14763);
nor U14950 (N_14950,N_14780,N_14813);
xnor U14951 (N_14951,N_14851,N_14830);
nor U14952 (N_14952,N_14849,N_14817);
nor U14953 (N_14953,N_14772,N_14741);
xor U14954 (N_14954,N_14815,N_14877);
xnor U14955 (N_14955,N_14834,N_14773);
and U14956 (N_14956,N_14740,N_14873);
or U14957 (N_14957,N_14799,N_14752);
and U14958 (N_14958,N_14793,N_14835);
nor U14959 (N_14959,N_14802,N_14832);
nand U14960 (N_14960,N_14737,N_14738);
nor U14961 (N_14961,N_14808,N_14803);
and U14962 (N_14962,N_14878,N_14867);
or U14963 (N_14963,N_14864,N_14726);
nand U14964 (N_14964,N_14730,N_14854);
and U14965 (N_14965,N_14746,N_14809);
nand U14966 (N_14966,N_14814,N_14873);
or U14967 (N_14967,N_14736,N_14824);
nor U14968 (N_14968,N_14842,N_14789);
xnor U14969 (N_14969,N_14802,N_14734);
and U14970 (N_14970,N_14839,N_14729);
nand U14971 (N_14971,N_14812,N_14873);
nand U14972 (N_14972,N_14778,N_14729);
xnor U14973 (N_14973,N_14743,N_14732);
nor U14974 (N_14974,N_14721,N_14826);
and U14975 (N_14975,N_14810,N_14747);
nand U14976 (N_14976,N_14863,N_14848);
and U14977 (N_14977,N_14755,N_14744);
and U14978 (N_14978,N_14749,N_14768);
or U14979 (N_14979,N_14819,N_14729);
nor U14980 (N_14980,N_14836,N_14870);
xnor U14981 (N_14981,N_14792,N_14751);
and U14982 (N_14982,N_14732,N_14815);
nor U14983 (N_14983,N_14762,N_14749);
nor U14984 (N_14984,N_14730,N_14827);
and U14985 (N_14985,N_14811,N_14874);
nor U14986 (N_14986,N_14859,N_14826);
and U14987 (N_14987,N_14746,N_14827);
nor U14988 (N_14988,N_14752,N_14845);
or U14989 (N_14989,N_14862,N_14776);
and U14990 (N_14990,N_14816,N_14762);
nand U14991 (N_14991,N_14768,N_14726);
xnor U14992 (N_14992,N_14866,N_14857);
and U14993 (N_14993,N_14774,N_14738);
xor U14994 (N_14994,N_14795,N_14747);
nand U14995 (N_14995,N_14770,N_14852);
nor U14996 (N_14996,N_14735,N_14797);
and U14997 (N_14997,N_14831,N_14752);
xnor U14998 (N_14998,N_14757,N_14813);
nor U14999 (N_14999,N_14786,N_14782);
xor U15000 (N_15000,N_14751,N_14798);
nand U15001 (N_15001,N_14812,N_14737);
xnor U15002 (N_15002,N_14778,N_14802);
nand U15003 (N_15003,N_14825,N_14821);
and U15004 (N_15004,N_14790,N_14805);
and U15005 (N_15005,N_14848,N_14776);
or U15006 (N_15006,N_14746,N_14796);
nor U15007 (N_15007,N_14809,N_14729);
nand U15008 (N_15008,N_14769,N_14797);
and U15009 (N_15009,N_14742,N_14812);
nand U15010 (N_15010,N_14840,N_14866);
nand U15011 (N_15011,N_14876,N_14809);
xnor U15012 (N_15012,N_14871,N_14837);
xnor U15013 (N_15013,N_14820,N_14876);
nand U15014 (N_15014,N_14741,N_14829);
nand U15015 (N_15015,N_14801,N_14852);
nor U15016 (N_15016,N_14837,N_14839);
or U15017 (N_15017,N_14732,N_14788);
nor U15018 (N_15018,N_14776,N_14872);
or U15019 (N_15019,N_14845,N_14838);
nor U15020 (N_15020,N_14873,N_14796);
xnor U15021 (N_15021,N_14733,N_14778);
xor U15022 (N_15022,N_14773,N_14777);
or U15023 (N_15023,N_14827,N_14781);
xor U15024 (N_15024,N_14739,N_14759);
and U15025 (N_15025,N_14746,N_14805);
nor U15026 (N_15026,N_14775,N_14777);
nor U15027 (N_15027,N_14738,N_14744);
and U15028 (N_15028,N_14827,N_14738);
nand U15029 (N_15029,N_14822,N_14782);
and U15030 (N_15030,N_14856,N_14858);
xor U15031 (N_15031,N_14822,N_14762);
nand U15032 (N_15032,N_14791,N_14878);
or U15033 (N_15033,N_14731,N_14840);
nand U15034 (N_15034,N_14814,N_14817);
and U15035 (N_15035,N_14858,N_14755);
and U15036 (N_15036,N_14766,N_14794);
and U15037 (N_15037,N_14744,N_14764);
nor U15038 (N_15038,N_14768,N_14870);
or U15039 (N_15039,N_14827,N_14754);
nor U15040 (N_15040,N_14991,N_15038);
or U15041 (N_15041,N_15023,N_14961);
xor U15042 (N_15042,N_15009,N_14992);
or U15043 (N_15043,N_15035,N_15029);
xnor U15044 (N_15044,N_14996,N_14999);
and U15045 (N_15045,N_14988,N_15007);
xor U15046 (N_15046,N_14913,N_15018);
nor U15047 (N_15047,N_14973,N_15000);
and U15048 (N_15048,N_14933,N_14919);
or U15049 (N_15049,N_14984,N_14974);
nor U15050 (N_15050,N_14883,N_14956);
nand U15051 (N_15051,N_15005,N_14901);
and U15052 (N_15052,N_14920,N_14914);
and U15053 (N_15053,N_14986,N_14911);
xnor U15054 (N_15054,N_14982,N_15006);
nor U15055 (N_15055,N_14975,N_14953);
nand U15056 (N_15056,N_14963,N_14949);
and U15057 (N_15057,N_14929,N_15025);
and U15058 (N_15058,N_14902,N_14959);
and U15059 (N_15059,N_14928,N_14931);
or U15060 (N_15060,N_14990,N_14979);
nor U15061 (N_15061,N_14910,N_15003);
or U15062 (N_15062,N_14970,N_14969);
or U15063 (N_15063,N_14889,N_14941);
nor U15064 (N_15064,N_14947,N_14939);
and U15065 (N_15065,N_14987,N_14932);
or U15066 (N_15066,N_14927,N_14894);
xnor U15067 (N_15067,N_15037,N_15024);
or U15068 (N_15068,N_14917,N_14907);
or U15069 (N_15069,N_14942,N_14938);
or U15070 (N_15070,N_14976,N_14989);
and U15071 (N_15071,N_15030,N_14897);
xnor U15072 (N_15072,N_15020,N_15011);
nor U15073 (N_15073,N_15019,N_14971);
xnor U15074 (N_15074,N_14903,N_14916);
xnor U15075 (N_15075,N_14899,N_14952);
and U15076 (N_15076,N_15008,N_15028);
nor U15077 (N_15077,N_14918,N_14946);
xor U15078 (N_15078,N_14896,N_15027);
nand U15079 (N_15079,N_14882,N_15032);
xor U15080 (N_15080,N_14937,N_14900);
xor U15081 (N_15081,N_14921,N_14922);
nand U15082 (N_15082,N_14925,N_15016);
or U15083 (N_15083,N_14951,N_14985);
nor U15084 (N_15084,N_14964,N_14998);
or U15085 (N_15085,N_14945,N_14967);
nor U15086 (N_15086,N_14977,N_14943);
and U15087 (N_15087,N_14891,N_14978);
nand U15088 (N_15088,N_14958,N_14880);
nand U15089 (N_15089,N_14887,N_15010);
nand U15090 (N_15090,N_14983,N_14935);
nor U15091 (N_15091,N_14915,N_14905);
nor U15092 (N_15092,N_14995,N_14965);
nand U15093 (N_15093,N_14957,N_15015);
nor U15094 (N_15094,N_14923,N_14893);
or U15095 (N_15095,N_14930,N_14966);
nand U15096 (N_15096,N_14934,N_14981);
xnor U15097 (N_15097,N_14912,N_14885);
nand U15098 (N_15098,N_15034,N_15014);
and U15099 (N_15099,N_14994,N_15021);
xor U15100 (N_15100,N_14924,N_14948);
nor U15101 (N_15101,N_14993,N_14954);
nand U15102 (N_15102,N_14950,N_15001);
nand U15103 (N_15103,N_14968,N_14944);
and U15104 (N_15104,N_14906,N_14908);
nor U15105 (N_15105,N_15036,N_14886);
xor U15106 (N_15106,N_14881,N_15004);
nor U15107 (N_15107,N_14909,N_14926);
nand U15108 (N_15108,N_14892,N_14997);
and U15109 (N_15109,N_14962,N_14980);
and U15110 (N_15110,N_14955,N_15012);
and U15111 (N_15111,N_15039,N_14898);
nand U15112 (N_15112,N_14936,N_15002);
nand U15113 (N_15113,N_14884,N_15026);
nor U15114 (N_15114,N_15031,N_14888);
nand U15115 (N_15115,N_15013,N_14972);
xnor U15116 (N_15116,N_15022,N_14960);
nor U15117 (N_15117,N_14904,N_15017);
nand U15118 (N_15118,N_14940,N_15033);
nor U15119 (N_15119,N_14890,N_14895);
nor U15120 (N_15120,N_14996,N_14970);
nor U15121 (N_15121,N_14979,N_14905);
or U15122 (N_15122,N_14932,N_15006);
and U15123 (N_15123,N_15027,N_14960);
nand U15124 (N_15124,N_14912,N_14961);
xor U15125 (N_15125,N_14928,N_14941);
nand U15126 (N_15126,N_15019,N_15035);
nor U15127 (N_15127,N_14882,N_14903);
or U15128 (N_15128,N_14946,N_14953);
nor U15129 (N_15129,N_14969,N_14932);
xnor U15130 (N_15130,N_14887,N_14898);
xor U15131 (N_15131,N_15023,N_14986);
xor U15132 (N_15132,N_15025,N_15003);
xor U15133 (N_15133,N_14968,N_14973);
or U15134 (N_15134,N_14980,N_14986);
and U15135 (N_15135,N_14921,N_14941);
and U15136 (N_15136,N_15038,N_14903);
nand U15137 (N_15137,N_14918,N_14986);
and U15138 (N_15138,N_14958,N_14945);
nor U15139 (N_15139,N_14990,N_14974);
xnor U15140 (N_15140,N_14968,N_14992);
xor U15141 (N_15141,N_14983,N_14917);
nor U15142 (N_15142,N_14883,N_14965);
xnor U15143 (N_15143,N_15022,N_15015);
and U15144 (N_15144,N_14966,N_14916);
nand U15145 (N_15145,N_14910,N_15015);
nor U15146 (N_15146,N_14926,N_14898);
and U15147 (N_15147,N_14947,N_14883);
nand U15148 (N_15148,N_14937,N_14947);
and U15149 (N_15149,N_14981,N_14999);
nand U15150 (N_15150,N_14902,N_14966);
nand U15151 (N_15151,N_14939,N_14963);
xor U15152 (N_15152,N_14943,N_14959);
nand U15153 (N_15153,N_15024,N_14893);
nand U15154 (N_15154,N_14990,N_15039);
xnor U15155 (N_15155,N_14917,N_15021);
xnor U15156 (N_15156,N_14928,N_14989);
nor U15157 (N_15157,N_14941,N_15031);
and U15158 (N_15158,N_15011,N_14888);
nor U15159 (N_15159,N_15007,N_14937);
or U15160 (N_15160,N_14890,N_15027);
nand U15161 (N_15161,N_14935,N_14924);
nand U15162 (N_15162,N_14925,N_14930);
or U15163 (N_15163,N_14894,N_14984);
and U15164 (N_15164,N_14986,N_14938);
xor U15165 (N_15165,N_14989,N_15034);
nand U15166 (N_15166,N_14970,N_14883);
nor U15167 (N_15167,N_15030,N_14990);
and U15168 (N_15168,N_14940,N_14935);
and U15169 (N_15169,N_14918,N_14944);
nand U15170 (N_15170,N_15001,N_15019);
or U15171 (N_15171,N_14914,N_14987);
and U15172 (N_15172,N_14996,N_14925);
and U15173 (N_15173,N_14934,N_15038);
xor U15174 (N_15174,N_15023,N_14930);
and U15175 (N_15175,N_15017,N_14964);
nor U15176 (N_15176,N_14996,N_14940);
xnor U15177 (N_15177,N_14963,N_15005);
xnor U15178 (N_15178,N_15026,N_14898);
nor U15179 (N_15179,N_14902,N_14930);
or U15180 (N_15180,N_14910,N_15032);
and U15181 (N_15181,N_15004,N_14944);
nand U15182 (N_15182,N_14945,N_14906);
and U15183 (N_15183,N_15000,N_15031);
nand U15184 (N_15184,N_15019,N_15023);
or U15185 (N_15185,N_15009,N_14917);
nand U15186 (N_15186,N_15020,N_14923);
and U15187 (N_15187,N_14929,N_14954);
and U15188 (N_15188,N_14996,N_14998);
or U15189 (N_15189,N_14927,N_14951);
nor U15190 (N_15190,N_15026,N_14917);
nor U15191 (N_15191,N_14932,N_14934);
xor U15192 (N_15192,N_14937,N_15004);
and U15193 (N_15193,N_14881,N_14983);
or U15194 (N_15194,N_14886,N_14907);
nand U15195 (N_15195,N_15023,N_14988);
and U15196 (N_15196,N_14949,N_14970);
nor U15197 (N_15197,N_14948,N_14939);
xor U15198 (N_15198,N_14944,N_14921);
nor U15199 (N_15199,N_14921,N_14883);
or U15200 (N_15200,N_15131,N_15049);
nor U15201 (N_15201,N_15136,N_15153);
xor U15202 (N_15202,N_15124,N_15185);
or U15203 (N_15203,N_15171,N_15073);
nand U15204 (N_15204,N_15170,N_15068);
nor U15205 (N_15205,N_15059,N_15168);
or U15206 (N_15206,N_15194,N_15112);
and U15207 (N_15207,N_15106,N_15055);
xor U15208 (N_15208,N_15181,N_15076);
or U15209 (N_15209,N_15145,N_15061);
and U15210 (N_15210,N_15159,N_15167);
xnor U15211 (N_15211,N_15120,N_15161);
and U15212 (N_15212,N_15157,N_15133);
nand U15213 (N_15213,N_15151,N_15066);
and U15214 (N_15214,N_15137,N_15111);
or U15215 (N_15215,N_15116,N_15041);
nor U15216 (N_15216,N_15083,N_15091);
nor U15217 (N_15217,N_15057,N_15075);
or U15218 (N_15218,N_15043,N_15180);
or U15219 (N_15219,N_15177,N_15187);
nor U15220 (N_15220,N_15155,N_15195);
or U15221 (N_15221,N_15045,N_15087);
or U15222 (N_15222,N_15048,N_15152);
xor U15223 (N_15223,N_15064,N_15184);
nand U15224 (N_15224,N_15058,N_15072);
nor U15225 (N_15225,N_15164,N_15085);
and U15226 (N_15226,N_15098,N_15046);
nor U15227 (N_15227,N_15188,N_15050);
or U15228 (N_15228,N_15127,N_15178);
nand U15229 (N_15229,N_15088,N_15162);
and U15230 (N_15230,N_15123,N_15062);
xnor U15231 (N_15231,N_15063,N_15189);
and U15232 (N_15232,N_15154,N_15092);
nand U15233 (N_15233,N_15196,N_15070);
nand U15234 (N_15234,N_15126,N_15069);
or U15235 (N_15235,N_15090,N_15121);
nand U15236 (N_15236,N_15146,N_15093);
xnor U15237 (N_15237,N_15156,N_15165);
and U15238 (N_15238,N_15163,N_15102);
nor U15239 (N_15239,N_15174,N_15089);
nor U15240 (N_15240,N_15147,N_15107);
nor U15241 (N_15241,N_15130,N_15125);
nand U15242 (N_15242,N_15141,N_15110);
or U15243 (N_15243,N_15176,N_15135);
or U15244 (N_15244,N_15139,N_15175);
nand U15245 (N_15245,N_15118,N_15053);
or U15246 (N_15246,N_15074,N_15095);
nand U15247 (N_15247,N_15117,N_15160);
xor U15248 (N_15248,N_15190,N_15079);
or U15249 (N_15249,N_15128,N_15084);
or U15250 (N_15250,N_15179,N_15191);
xnor U15251 (N_15251,N_15056,N_15096);
xnor U15252 (N_15252,N_15101,N_15142);
or U15253 (N_15253,N_15042,N_15182);
and U15254 (N_15254,N_15103,N_15108);
nor U15255 (N_15255,N_15199,N_15054);
nor U15256 (N_15256,N_15094,N_15169);
and U15257 (N_15257,N_15172,N_15122);
and U15258 (N_15258,N_15115,N_15044);
xor U15259 (N_15259,N_15149,N_15158);
or U15260 (N_15260,N_15104,N_15097);
nand U15261 (N_15261,N_15114,N_15040);
or U15262 (N_15262,N_15047,N_15099);
and U15263 (N_15263,N_15060,N_15113);
xor U15264 (N_15264,N_15119,N_15192);
nand U15265 (N_15265,N_15193,N_15197);
or U15266 (N_15266,N_15086,N_15144);
and U15267 (N_15267,N_15109,N_15148);
nor U15268 (N_15268,N_15071,N_15132);
nand U15269 (N_15269,N_15105,N_15052);
nand U15270 (N_15270,N_15143,N_15078);
nor U15271 (N_15271,N_15150,N_15067);
or U15272 (N_15272,N_15138,N_15134);
or U15273 (N_15273,N_15077,N_15065);
nand U15274 (N_15274,N_15080,N_15198);
or U15275 (N_15275,N_15173,N_15129);
or U15276 (N_15276,N_15081,N_15183);
and U15277 (N_15277,N_15100,N_15082);
xor U15278 (N_15278,N_15140,N_15051);
or U15279 (N_15279,N_15166,N_15186);
xor U15280 (N_15280,N_15185,N_15072);
xor U15281 (N_15281,N_15083,N_15183);
xor U15282 (N_15282,N_15049,N_15116);
nor U15283 (N_15283,N_15165,N_15098);
or U15284 (N_15284,N_15173,N_15154);
nor U15285 (N_15285,N_15195,N_15140);
and U15286 (N_15286,N_15190,N_15119);
xnor U15287 (N_15287,N_15190,N_15183);
or U15288 (N_15288,N_15040,N_15199);
xor U15289 (N_15289,N_15045,N_15047);
or U15290 (N_15290,N_15057,N_15170);
nor U15291 (N_15291,N_15091,N_15110);
and U15292 (N_15292,N_15085,N_15134);
and U15293 (N_15293,N_15137,N_15060);
or U15294 (N_15294,N_15081,N_15170);
nand U15295 (N_15295,N_15070,N_15098);
nand U15296 (N_15296,N_15154,N_15197);
and U15297 (N_15297,N_15181,N_15110);
nor U15298 (N_15298,N_15119,N_15181);
or U15299 (N_15299,N_15107,N_15112);
and U15300 (N_15300,N_15195,N_15148);
xor U15301 (N_15301,N_15090,N_15098);
nor U15302 (N_15302,N_15146,N_15088);
xor U15303 (N_15303,N_15135,N_15193);
and U15304 (N_15304,N_15138,N_15152);
nor U15305 (N_15305,N_15137,N_15143);
xnor U15306 (N_15306,N_15092,N_15082);
or U15307 (N_15307,N_15092,N_15197);
or U15308 (N_15308,N_15118,N_15120);
nand U15309 (N_15309,N_15137,N_15073);
nor U15310 (N_15310,N_15123,N_15075);
nor U15311 (N_15311,N_15141,N_15126);
and U15312 (N_15312,N_15172,N_15095);
or U15313 (N_15313,N_15174,N_15153);
or U15314 (N_15314,N_15123,N_15040);
or U15315 (N_15315,N_15172,N_15070);
and U15316 (N_15316,N_15088,N_15095);
nand U15317 (N_15317,N_15153,N_15054);
and U15318 (N_15318,N_15145,N_15050);
and U15319 (N_15319,N_15070,N_15152);
nand U15320 (N_15320,N_15079,N_15134);
or U15321 (N_15321,N_15127,N_15044);
and U15322 (N_15322,N_15125,N_15091);
nand U15323 (N_15323,N_15107,N_15197);
and U15324 (N_15324,N_15047,N_15067);
or U15325 (N_15325,N_15045,N_15168);
or U15326 (N_15326,N_15178,N_15044);
or U15327 (N_15327,N_15182,N_15106);
xor U15328 (N_15328,N_15178,N_15098);
and U15329 (N_15329,N_15090,N_15146);
and U15330 (N_15330,N_15068,N_15143);
nand U15331 (N_15331,N_15099,N_15153);
nor U15332 (N_15332,N_15132,N_15189);
or U15333 (N_15333,N_15070,N_15162);
nor U15334 (N_15334,N_15081,N_15116);
or U15335 (N_15335,N_15140,N_15054);
and U15336 (N_15336,N_15153,N_15190);
and U15337 (N_15337,N_15131,N_15118);
nor U15338 (N_15338,N_15081,N_15110);
xnor U15339 (N_15339,N_15166,N_15098);
xor U15340 (N_15340,N_15097,N_15130);
or U15341 (N_15341,N_15067,N_15186);
xor U15342 (N_15342,N_15178,N_15163);
or U15343 (N_15343,N_15074,N_15135);
and U15344 (N_15344,N_15111,N_15040);
and U15345 (N_15345,N_15056,N_15128);
nand U15346 (N_15346,N_15195,N_15102);
nand U15347 (N_15347,N_15092,N_15044);
nor U15348 (N_15348,N_15110,N_15170);
or U15349 (N_15349,N_15104,N_15076);
xnor U15350 (N_15350,N_15123,N_15069);
xnor U15351 (N_15351,N_15133,N_15055);
nor U15352 (N_15352,N_15153,N_15094);
nor U15353 (N_15353,N_15141,N_15194);
xnor U15354 (N_15354,N_15104,N_15040);
or U15355 (N_15355,N_15152,N_15171);
xnor U15356 (N_15356,N_15107,N_15088);
or U15357 (N_15357,N_15153,N_15111);
nor U15358 (N_15358,N_15165,N_15135);
or U15359 (N_15359,N_15164,N_15065);
or U15360 (N_15360,N_15255,N_15314);
nand U15361 (N_15361,N_15290,N_15240);
or U15362 (N_15362,N_15208,N_15311);
and U15363 (N_15363,N_15348,N_15217);
nor U15364 (N_15364,N_15310,N_15267);
or U15365 (N_15365,N_15296,N_15249);
and U15366 (N_15366,N_15328,N_15315);
xor U15367 (N_15367,N_15346,N_15294);
nand U15368 (N_15368,N_15220,N_15322);
nand U15369 (N_15369,N_15285,N_15237);
xnor U15370 (N_15370,N_15289,N_15352);
or U15371 (N_15371,N_15250,N_15333);
or U15372 (N_15372,N_15308,N_15279);
nor U15373 (N_15373,N_15326,N_15319);
xor U15374 (N_15374,N_15209,N_15235);
nand U15375 (N_15375,N_15339,N_15251);
or U15376 (N_15376,N_15273,N_15280);
xnor U15377 (N_15377,N_15205,N_15212);
or U15378 (N_15378,N_15349,N_15272);
and U15379 (N_15379,N_15295,N_15283);
nand U15380 (N_15380,N_15330,N_15262);
nor U15381 (N_15381,N_15232,N_15317);
and U15382 (N_15382,N_15231,N_15202);
nand U15383 (N_15383,N_15358,N_15284);
and U15384 (N_15384,N_15357,N_15276);
xor U15385 (N_15385,N_15344,N_15312);
and U15386 (N_15386,N_15261,N_15274);
and U15387 (N_15387,N_15281,N_15353);
nor U15388 (N_15388,N_15218,N_15304);
or U15389 (N_15389,N_15313,N_15203);
or U15390 (N_15390,N_15229,N_15236);
or U15391 (N_15391,N_15243,N_15226);
xnor U15392 (N_15392,N_15343,N_15324);
or U15393 (N_15393,N_15297,N_15222);
and U15394 (N_15394,N_15270,N_15221);
and U15395 (N_15395,N_15309,N_15325);
and U15396 (N_15396,N_15327,N_15233);
nor U15397 (N_15397,N_15248,N_15356);
nor U15398 (N_15398,N_15287,N_15265);
xor U15399 (N_15399,N_15345,N_15291);
nand U15400 (N_15400,N_15275,N_15207);
or U15401 (N_15401,N_15245,N_15223);
nand U15402 (N_15402,N_15351,N_15266);
xor U15403 (N_15403,N_15307,N_15268);
or U15404 (N_15404,N_15263,N_15302);
nand U15405 (N_15405,N_15201,N_15225);
or U15406 (N_15406,N_15224,N_15258);
xnor U15407 (N_15407,N_15350,N_15278);
or U15408 (N_15408,N_15323,N_15340);
or U15409 (N_15409,N_15341,N_15216);
xnor U15410 (N_15410,N_15277,N_15305);
or U15411 (N_15411,N_15336,N_15355);
nand U15412 (N_15412,N_15219,N_15299);
xnor U15413 (N_15413,N_15259,N_15354);
nor U15414 (N_15414,N_15329,N_15337);
or U15415 (N_15415,N_15288,N_15227);
or U15416 (N_15416,N_15332,N_15316);
or U15417 (N_15417,N_15234,N_15306);
nor U15418 (N_15418,N_15303,N_15230);
nand U15419 (N_15419,N_15204,N_15253);
xnor U15420 (N_15420,N_15293,N_15241);
xnor U15421 (N_15421,N_15228,N_15215);
xnor U15422 (N_15422,N_15286,N_15359);
nand U15423 (N_15423,N_15256,N_15260);
xnor U15424 (N_15424,N_15252,N_15347);
nor U15425 (N_15425,N_15242,N_15338);
nand U15426 (N_15426,N_15298,N_15246);
nor U15427 (N_15427,N_15335,N_15206);
or U15428 (N_15428,N_15320,N_15334);
nand U15429 (N_15429,N_15264,N_15210);
xnor U15430 (N_15430,N_15247,N_15213);
xor U15431 (N_15431,N_15321,N_15269);
or U15432 (N_15432,N_15244,N_15331);
nand U15433 (N_15433,N_15211,N_15214);
xnor U15434 (N_15434,N_15239,N_15200);
and U15435 (N_15435,N_15292,N_15342);
xor U15436 (N_15436,N_15318,N_15257);
nand U15437 (N_15437,N_15301,N_15238);
and U15438 (N_15438,N_15300,N_15271);
nand U15439 (N_15439,N_15254,N_15282);
nor U15440 (N_15440,N_15247,N_15304);
nor U15441 (N_15441,N_15230,N_15243);
nand U15442 (N_15442,N_15286,N_15348);
nand U15443 (N_15443,N_15214,N_15284);
nor U15444 (N_15444,N_15337,N_15312);
nand U15445 (N_15445,N_15256,N_15255);
nor U15446 (N_15446,N_15358,N_15214);
or U15447 (N_15447,N_15352,N_15253);
nor U15448 (N_15448,N_15348,N_15332);
xnor U15449 (N_15449,N_15267,N_15338);
nor U15450 (N_15450,N_15346,N_15246);
nand U15451 (N_15451,N_15282,N_15339);
and U15452 (N_15452,N_15359,N_15261);
nand U15453 (N_15453,N_15315,N_15299);
nor U15454 (N_15454,N_15293,N_15221);
nor U15455 (N_15455,N_15200,N_15292);
nor U15456 (N_15456,N_15343,N_15357);
xnor U15457 (N_15457,N_15263,N_15272);
nand U15458 (N_15458,N_15257,N_15288);
nor U15459 (N_15459,N_15294,N_15240);
nor U15460 (N_15460,N_15202,N_15247);
nand U15461 (N_15461,N_15200,N_15241);
nor U15462 (N_15462,N_15326,N_15269);
nor U15463 (N_15463,N_15208,N_15246);
or U15464 (N_15464,N_15309,N_15328);
nor U15465 (N_15465,N_15281,N_15357);
or U15466 (N_15466,N_15289,N_15247);
nor U15467 (N_15467,N_15231,N_15219);
nor U15468 (N_15468,N_15302,N_15280);
and U15469 (N_15469,N_15247,N_15358);
nor U15470 (N_15470,N_15291,N_15293);
xnor U15471 (N_15471,N_15343,N_15235);
nor U15472 (N_15472,N_15201,N_15359);
and U15473 (N_15473,N_15256,N_15247);
or U15474 (N_15474,N_15249,N_15217);
nor U15475 (N_15475,N_15243,N_15219);
xor U15476 (N_15476,N_15268,N_15291);
nand U15477 (N_15477,N_15258,N_15291);
nor U15478 (N_15478,N_15297,N_15281);
xor U15479 (N_15479,N_15206,N_15250);
nor U15480 (N_15480,N_15255,N_15310);
xnor U15481 (N_15481,N_15322,N_15296);
and U15482 (N_15482,N_15266,N_15303);
nor U15483 (N_15483,N_15290,N_15351);
xnor U15484 (N_15484,N_15292,N_15344);
or U15485 (N_15485,N_15312,N_15324);
xor U15486 (N_15486,N_15224,N_15335);
xor U15487 (N_15487,N_15316,N_15220);
nand U15488 (N_15488,N_15268,N_15264);
xor U15489 (N_15489,N_15269,N_15288);
and U15490 (N_15490,N_15263,N_15315);
and U15491 (N_15491,N_15301,N_15263);
nand U15492 (N_15492,N_15216,N_15221);
and U15493 (N_15493,N_15260,N_15349);
xnor U15494 (N_15494,N_15340,N_15359);
xnor U15495 (N_15495,N_15341,N_15359);
nor U15496 (N_15496,N_15335,N_15297);
or U15497 (N_15497,N_15289,N_15260);
or U15498 (N_15498,N_15334,N_15202);
nand U15499 (N_15499,N_15205,N_15223);
and U15500 (N_15500,N_15221,N_15275);
nand U15501 (N_15501,N_15271,N_15237);
and U15502 (N_15502,N_15293,N_15257);
or U15503 (N_15503,N_15359,N_15268);
nand U15504 (N_15504,N_15317,N_15230);
and U15505 (N_15505,N_15297,N_15241);
xnor U15506 (N_15506,N_15302,N_15224);
xnor U15507 (N_15507,N_15205,N_15329);
or U15508 (N_15508,N_15341,N_15333);
or U15509 (N_15509,N_15336,N_15325);
and U15510 (N_15510,N_15209,N_15224);
and U15511 (N_15511,N_15329,N_15268);
and U15512 (N_15512,N_15271,N_15249);
or U15513 (N_15513,N_15236,N_15212);
nor U15514 (N_15514,N_15278,N_15322);
and U15515 (N_15515,N_15249,N_15313);
xor U15516 (N_15516,N_15357,N_15286);
or U15517 (N_15517,N_15239,N_15333);
nand U15518 (N_15518,N_15204,N_15221);
nor U15519 (N_15519,N_15239,N_15346);
or U15520 (N_15520,N_15379,N_15409);
or U15521 (N_15521,N_15410,N_15486);
xor U15522 (N_15522,N_15480,N_15456);
or U15523 (N_15523,N_15515,N_15362);
or U15524 (N_15524,N_15504,N_15422);
and U15525 (N_15525,N_15374,N_15412);
xnor U15526 (N_15526,N_15426,N_15494);
nand U15527 (N_15527,N_15376,N_15500);
or U15528 (N_15528,N_15427,N_15478);
or U15529 (N_15529,N_15493,N_15436);
and U15530 (N_15530,N_15508,N_15377);
and U15531 (N_15531,N_15481,N_15461);
nor U15532 (N_15532,N_15503,N_15437);
or U15533 (N_15533,N_15473,N_15511);
or U15534 (N_15534,N_15385,N_15502);
nor U15535 (N_15535,N_15498,N_15397);
or U15536 (N_15536,N_15505,N_15429);
nor U15537 (N_15537,N_15469,N_15491);
or U15538 (N_15538,N_15395,N_15370);
nor U15539 (N_15539,N_15463,N_15390);
nor U15540 (N_15540,N_15518,N_15381);
and U15541 (N_15541,N_15387,N_15372);
and U15542 (N_15542,N_15389,N_15430);
and U15543 (N_15543,N_15432,N_15516);
xnor U15544 (N_15544,N_15440,N_15490);
nor U15545 (N_15545,N_15378,N_15419);
nand U15546 (N_15546,N_15454,N_15363);
nand U15547 (N_15547,N_15401,N_15512);
xnor U15548 (N_15548,N_15452,N_15414);
nand U15549 (N_15549,N_15425,N_15479);
and U15550 (N_15550,N_15509,N_15406);
xnor U15551 (N_15551,N_15392,N_15420);
and U15552 (N_15552,N_15496,N_15448);
nor U15553 (N_15553,N_15472,N_15364);
or U15554 (N_15554,N_15391,N_15441);
or U15555 (N_15555,N_15442,N_15438);
and U15556 (N_15556,N_15433,N_15462);
or U15557 (N_15557,N_15482,N_15371);
nor U15558 (N_15558,N_15475,N_15517);
or U15559 (N_15559,N_15488,N_15449);
or U15560 (N_15560,N_15396,N_15519);
xor U15561 (N_15561,N_15470,N_15402);
xnor U15562 (N_15562,N_15444,N_15418);
xor U15563 (N_15563,N_15484,N_15366);
or U15564 (N_15564,N_15375,N_15487);
nor U15565 (N_15565,N_15380,N_15360);
and U15566 (N_15566,N_15388,N_15439);
and U15567 (N_15567,N_15501,N_15499);
nand U15568 (N_15568,N_15394,N_15453);
or U15569 (N_15569,N_15492,N_15382);
or U15570 (N_15570,N_15495,N_15510);
nor U15571 (N_15571,N_15468,N_15431);
nor U15572 (N_15572,N_15411,N_15455);
xnor U15573 (N_15573,N_15506,N_15365);
xor U15574 (N_15574,N_15458,N_15393);
xnor U15575 (N_15575,N_15383,N_15416);
nand U15576 (N_15576,N_15413,N_15373);
and U15577 (N_15577,N_15368,N_15451);
xor U15578 (N_15578,N_15405,N_15513);
and U15579 (N_15579,N_15404,N_15464);
nor U15580 (N_15580,N_15445,N_15399);
nor U15581 (N_15581,N_15434,N_15384);
or U15582 (N_15582,N_15403,N_15457);
nor U15583 (N_15583,N_15459,N_15408);
nand U15584 (N_15584,N_15386,N_15407);
nand U15585 (N_15585,N_15476,N_15483);
nand U15586 (N_15586,N_15466,N_15507);
or U15587 (N_15587,N_15471,N_15400);
and U15588 (N_15588,N_15424,N_15467);
or U15589 (N_15589,N_15460,N_15450);
or U15590 (N_15590,N_15435,N_15398);
xor U15591 (N_15591,N_15465,N_15423);
nor U15592 (N_15592,N_15489,N_15485);
nand U15593 (N_15593,N_15443,N_15367);
nor U15594 (N_15594,N_15514,N_15447);
nor U15595 (N_15595,N_15497,N_15417);
nor U15596 (N_15596,N_15474,N_15369);
or U15597 (N_15597,N_15446,N_15477);
xor U15598 (N_15598,N_15361,N_15421);
and U15599 (N_15599,N_15428,N_15415);
nand U15600 (N_15600,N_15439,N_15386);
and U15601 (N_15601,N_15516,N_15510);
nor U15602 (N_15602,N_15388,N_15468);
and U15603 (N_15603,N_15459,N_15389);
xor U15604 (N_15604,N_15511,N_15441);
and U15605 (N_15605,N_15416,N_15441);
or U15606 (N_15606,N_15424,N_15458);
xor U15607 (N_15607,N_15493,N_15453);
or U15608 (N_15608,N_15363,N_15480);
and U15609 (N_15609,N_15395,N_15378);
xnor U15610 (N_15610,N_15441,N_15480);
and U15611 (N_15611,N_15464,N_15424);
nor U15612 (N_15612,N_15453,N_15371);
or U15613 (N_15613,N_15372,N_15432);
nor U15614 (N_15614,N_15474,N_15466);
nand U15615 (N_15615,N_15454,N_15507);
nor U15616 (N_15616,N_15496,N_15500);
and U15617 (N_15617,N_15390,N_15448);
nor U15618 (N_15618,N_15379,N_15467);
and U15619 (N_15619,N_15403,N_15507);
nand U15620 (N_15620,N_15418,N_15396);
and U15621 (N_15621,N_15400,N_15466);
nor U15622 (N_15622,N_15415,N_15371);
nand U15623 (N_15623,N_15371,N_15396);
or U15624 (N_15624,N_15388,N_15498);
nand U15625 (N_15625,N_15422,N_15371);
nor U15626 (N_15626,N_15372,N_15456);
and U15627 (N_15627,N_15474,N_15400);
and U15628 (N_15628,N_15467,N_15496);
or U15629 (N_15629,N_15438,N_15374);
xnor U15630 (N_15630,N_15453,N_15423);
xor U15631 (N_15631,N_15420,N_15481);
xnor U15632 (N_15632,N_15366,N_15364);
nor U15633 (N_15633,N_15363,N_15442);
nor U15634 (N_15634,N_15406,N_15402);
nor U15635 (N_15635,N_15507,N_15473);
nand U15636 (N_15636,N_15424,N_15422);
nand U15637 (N_15637,N_15442,N_15475);
or U15638 (N_15638,N_15402,N_15411);
nor U15639 (N_15639,N_15515,N_15389);
and U15640 (N_15640,N_15392,N_15383);
nor U15641 (N_15641,N_15496,N_15427);
nand U15642 (N_15642,N_15507,N_15375);
nor U15643 (N_15643,N_15492,N_15367);
and U15644 (N_15644,N_15401,N_15441);
nand U15645 (N_15645,N_15484,N_15413);
nand U15646 (N_15646,N_15426,N_15502);
or U15647 (N_15647,N_15379,N_15452);
and U15648 (N_15648,N_15492,N_15434);
or U15649 (N_15649,N_15384,N_15448);
xor U15650 (N_15650,N_15416,N_15443);
or U15651 (N_15651,N_15421,N_15441);
nor U15652 (N_15652,N_15373,N_15400);
nand U15653 (N_15653,N_15506,N_15484);
nor U15654 (N_15654,N_15417,N_15421);
or U15655 (N_15655,N_15395,N_15422);
and U15656 (N_15656,N_15446,N_15479);
nor U15657 (N_15657,N_15411,N_15450);
nand U15658 (N_15658,N_15469,N_15468);
nor U15659 (N_15659,N_15377,N_15440);
nor U15660 (N_15660,N_15440,N_15430);
xor U15661 (N_15661,N_15494,N_15375);
nand U15662 (N_15662,N_15367,N_15450);
xor U15663 (N_15663,N_15372,N_15377);
nand U15664 (N_15664,N_15476,N_15421);
xnor U15665 (N_15665,N_15386,N_15460);
nor U15666 (N_15666,N_15366,N_15416);
or U15667 (N_15667,N_15394,N_15469);
or U15668 (N_15668,N_15466,N_15518);
nand U15669 (N_15669,N_15481,N_15366);
nand U15670 (N_15670,N_15363,N_15444);
nand U15671 (N_15671,N_15445,N_15420);
xor U15672 (N_15672,N_15392,N_15471);
nor U15673 (N_15673,N_15511,N_15420);
and U15674 (N_15674,N_15458,N_15363);
or U15675 (N_15675,N_15388,N_15474);
and U15676 (N_15676,N_15381,N_15450);
nor U15677 (N_15677,N_15475,N_15415);
and U15678 (N_15678,N_15480,N_15364);
nand U15679 (N_15679,N_15425,N_15397);
nand U15680 (N_15680,N_15576,N_15634);
xor U15681 (N_15681,N_15567,N_15642);
nor U15682 (N_15682,N_15578,N_15551);
nor U15683 (N_15683,N_15553,N_15591);
and U15684 (N_15684,N_15544,N_15646);
and U15685 (N_15685,N_15561,N_15543);
nor U15686 (N_15686,N_15524,N_15633);
nor U15687 (N_15687,N_15530,N_15556);
xor U15688 (N_15688,N_15638,N_15575);
nor U15689 (N_15689,N_15545,N_15619);
nand U15690 (N_15690,N_15552,N_15639);
xnor U15691 (N_15691,N_15532,N_15573);
nand U15692 (N_15692,N_15621,N_15649);
and U15693 (N_15693,N_15570,N_15527);
nor U15694 (N_15694,N_15669,N_15549);
nor U15695 (N_15695,N_15566,N_15558);
or U15696 (N_15696,N_15632,N_15600);
or U15697 (N_15697,N_15672,N_15577);
nand U15698 (N_15698,N_15550,N_15542);
xnor U15699 (N_15699,N_15562,N_15613);
or U15700 (N_15700,N_15664,N_15528);
or U15701 (N_15701,N_15546,N_15565);
and U15702 (N_15702,N_15523,N_15678);
or U15703 (N_15703,N_15531,N_15661);
nand U15704 (N_15704,N_15622,N_15538);
nor U15705 (N_15705,N_15571,N_15636);
or U15706 (N_15706,N_15588,N_15618);
nand U15707 (N_15707,N_15564,N_15569);
and U15708 (N_15708,N_15597,N_15590);
xor U15709 (N_15709,N_15626,N_15653);
and U15710 (N_15710,N_15677,N_15563);
nor U15711 (N_15711,N_15629,N_15596);
nor U15712 (N_15712,N_15594,N_15660);
nand U15713 (N_15713,N_15595,N_15635);
or U15714 (N_15714,N_15539,N_15628);
nor U15715 (N_15715,N_15587,N_15652);
nand U15716 (N_15716,N_15645,N_15560);
and U15717 (N_15717,N_15657,N_15602);
and U15718 (N_15718,N_15581,N_15593);
or U15719 (N_15719,N_15521,N_15607);
xnor U15720 (N_15720,N_15641,N_15520);
nand U15721 (N_15721,N_15604,N_15643);
and U15722 (N_15722,N_15659,N_15555);
or U15723 (N_15723,N_15579,N_15654);
nand U15724 (N_15724,N_15536,N_15585);
or U15725 (N_15725,N_15534,N_15663);
nor U15726 (N_15726,N_15548,N_15535);
nor U15727 (N_15727,N_15670,N_15611);
xnor U15728 (N_15728,N_15647,N_15614);
or U15729 (N_15729,N_15522,N_15612);
nand U15730 (N_15730,N_15526,N_15616);
nand U15731 (N_15731,N_15609,N_15656);
or U15732 (N_15732,N_15676,N_15671);
nor U15733 (N_15733,N_15525,N_15601);
nor U15734 (N_15734,N_15586,N_15537);
xnor U15735 (N_15735,N_15630,N_15624);
and U15736 (N_15736,N_15533,N_15572);
nand U15737 (N_15737,N_15673,N_15675);
nand U15738 (N_15738,N_15655,N_15667);
and U15739 (N_15739,N_15637,N_15625);
xnor U15740 (N_15740,N_15615,N_15557);
nor U15741 (N_15741,N_15651,N_15640);
nor U15742 (N_15742,N_15574,N_15580);
or U15743 (N_15743,N_15631,N_15627);
xor U15744 (N_15744,N_15584,N_15605);
xor U15745 (N_15745,N_15589,N_15623);
and U15746 (N_15746,N_15599,N_15648);
xnor U15747 (N_15747,N_15666,N_15547);
or U15748 (N_15748,N_15582,N_15668);
xor U15749 (N_15749,N_15617,N_15541);
nor U15750 (N_15750,N_15554,N_15559);
xor U15751 (N_15751,N_15606,N_15583);
nand U15752 (N_15752,N_15598,N_15644);
or U15753 (N_15753,N_15529,N_15662);
and U15754 (N_15754,N_15610,N_15568);
or U15755 (N_15755,N_15592,N_15540);
and U15756 (N_15756,N_15620,N_15603);
nand U15757 (N_15757,N_15674,N_15665);
nand U15758 (N_15758,N_15608,N_15658);
nand U15759 (N_15759,N_15679,N_15650);
nor U15760 (N_15760,N_15665,N_15553);
xor U15761 (N_15761,N_15607,N_15675);
xor U15762 (N_15762,N_15577,N_15596);
nand U15763 (N_15763,N_15559,N_15629);
xnor U15764 (N_15764,N_15599,N_15668);
nor U15765 (N_15765,N_15633,N_15535);
nor U15766 (N_15766,N_15675,N_15596);
or U15767 (N_15767,N_15537,N_15579);
or U15768 (N_15768,N_15521,N_15650);
or U15769 (N_15769,N_15532,N_15521);
xor U15770 (N_15770,N_15633,N_15570);
nor U15771 (N_15771,N_15557,N_15639);
or U15772 (N_15772,N_15615,N_15574);
xor U15773 (N_15773,N_15672,N_15527);
nand U15774 (N_15774,N_15531,N_15622);
xnor U15775 (N_15775,N_15568,N_15597);
and U15776 (N_15776,N_15567,N_15550);
nand U15777 (N_15777,N_15675,N_15533);
nor U15778 (N_15778,N_15617,N_15627);
xor U15779 (N_15779,N_15669,N_15610);
or U15780 (N_15780,N_15529,N_15583);
nor U15781 (N_15781,N_15678,N_15550);
and U15782 (N_15782,N_15553,N_15542);
xor U15783 (N_15783,N_15654,N_15600);
and U15784 (N_15784,N_15534,N_15531);
xnor U15785 (N_15785,N_15528,N_15595);
nor U15786 (N_15786,N_15642,N_15637);
nor U15787 (N_15787,N_15578,N_15539);
and U15788 (N_15788,N_15530,N_15532);
nand U15789 (N_15789,N_15671,N_15586);
nor U15790 (N_15790,N_15587,N_15600);
or U15791 (N_15791,N_15661,N_15625);
xnor U15792 (N_15792,N_15656,N_15637);
nand U15793 (N_15793,N_15542,N_15639);
xnor U15794 (N_15794,N_15633,N_15520);
nor U15795 (N_15795,N_15549,N_15543);
nor U15796 (N_15796,N_15538,N_15555);
nor U15797 (N_15797,N_15615,N_15539);
and U15798 (N_15798,N_15676,N_15603);
xnor U15799 (N_15799,N_15565,N_15615);
and U15800 (N_15800,N_15579,N_15604);
or U15801 (N_15801,N_15579,N_15526);
and U15802 (N_15802,N_15587,N_15523);
nor U15803 (N_15803,N_15669,N_15556);
xnor U15804 (N_15804,N_15658,N_15573);
or U15805 (N_15805,N_15539,N_15533);
and U15806 (N_15806,N_15614,N_15634);
xor U15807 (N_15807,N_15637,N_15653);
xnor U15808 (N_15808,N_15638,N_15659);
and U15809 (N_15809,N_15561,N_15532);
nor U15810 (N_15810,N_15666,N_15601);
nand U15811 (N_15811,N_15651,N_15535);
and U15812 (N_15812,N_15525,N_15649);
xor U15813 (N_15813,N_15523,N_15545);
and U15814 (N_15814,N_15555,N_15621);
xor U15815 (N_15815,N_15555,N_15627);
nand U15816 (N_15816,N_15646,N_15673);
nand U15817 (N_15817,N_15564,N_15595);
nor U15818 (N_15818,N_15602,N_15627);
or U15819 (N_15819,N_15595,N_15653);
or U15820 (N_15820,N_15554,N_15536);
and U15821 (N_15821,N_15588,N_15568);
nor U15822 (N_15822,N_15554,N_15543);
or U15823 (N_15823,N_15666,N_15545);
or U15824 (N_15824,N_15664,N_15663);
and U15825 (N_15825,N_15562,N_15594);
nor U15826 (N_15826,N_15584,N_15596);
nor U15827 (N_15827,N_15561,N_15610);
or U15828 (N_15828,N_15532,N_15578);
nand U15829 (N_15829,N_15597,N_15602);
and U15830 (N_15830,N_15598,N_15647);
nor U15831 (N_15831,N_15579,N_15612);
or U15832 (N_15832,N_15649,N_15642);
or U15833 (N_15833,N_15564,N_15646);
xor U15834 (N_15834,N_15620,N_15653);
and U15835 (N_15835,N_15559,N_15584);
or U15836 (N_15836,N_15617,N_15615);
and U15837 (N_15837,N_15587,N_15555);
or U15838 (N_15838,N_15667,N_15524);
and U15839 (N_15839,N_15648,N_15557);
nand U15840 (N_15840,N_15737,N_15684);
or U15841 (N_15841,N_15715,N_15721);
xnor U15842 (N_15842,N_15690,N_15832);
and U15843 (N_15843,N_15780,N_15803);
and U15844 (N_15844,N_15724,N_15680);
nand U15845 (N_15845,N_15783,N_15766);
xor U15846 (N_15846,N_15807,N_15726);
nor U15847 (N_15847,N_15770,N_15709);
nand U15848 (N_15848,N_15760,N_15686);
and U15849 (N_15849,N_15713,N_15816);
or U15850 (N_15850,N_15794,N_15809);
nand U15851 (N_15851,N_15784,N_15718);
and U15852 (N_15852,N_15827,N_15731);
nor U15853 (N_15853,N_15775,N_15812);
nor U15854 (N_15854,N_15759,N_15758);
and U15855 (N_15855,N_15817,N_15821);
xor U15856 (N_15856,N_15734,N_15723);
nand U15857 (N_15857,N_15838,N_15813);
and U15858 (N_15858,N_15786,N_15756);
nor U15859 (N_15859,N_15742,N_15746);
nor U15860 (N_15860,N_15730,N_15765);
xnor U15861 (N_15861,N_15699,N_15789);
nor U15862 (N_15862,N_15836,N_15739);
xnor U15863 (N_15863,N_15741,N_15693);
xnor U15864 (N_15864,N_15819,N_15762);
and U15865 (N_15865,N_15751,N_15768);
or U15866 (N_15866,N_15777,N_15773);
and U15867 (N_15867,N_15806,N_15705);
xnor U15868 (N_15868,N_15685,N_15771);
nor U15869 (N_15869,N_15797,N_15752);
or U15870 (N_15870,N_15732,N_15736);
or U15871 (N_15871,N_15772,N_15698);
and U15872 (N_15872,N_15703,N_15810);
nor U15873 (N_15873,N_15767,N_15785);
and U15874 (N_15874,N_15837,N_15802);
and U15875 (N_15875,N_15826,N_15834);
xnor U15876 (N_15876,N_15820,N_15788);
nand U15877 (N_15877,N_15687,N_15787);
nor U15878 (N_15878,N_15714,N_15811);
or U15879 (N_15879,N_15757,N_15804);
or U15880 (N_15880,N_15769,N_15750);
nor U15881 (N_15881,N_15808,N_15830);
and U15882 (N_15882,N_15745,N_15829);
or U15883 (N_15883,N_15740,N_15708);
and U15884 (N_15884,N_15798,N_15763);
xor U15885 (N_15885,N_15748,N_15725);
or U15886 (N_15886,N_15704,N_15793);
nand U15887 (N_15887,N_15697,N_15729);
and U15888 (N_15888,N_15683,N_15764);
or U15889 (N_15889,N_15744,N_15696);
nand U15890 (N_15890,N_15743,N_15831);
xor U15891 (N_15891,N_15822,N_15689);
nor U15892 (N_15892,N_15776,N_15728);
or U15893 (N_15893,N_15800,N_15706);
or U15894 (N_15894,N_15755,N_15694);
or U15895 (N_15895,N_15839,N_15738);
xor U15896 (N_15896,N_15707,N_15717);
xnor U15897 (N_15897,N_15735,N_15691);
or U15898 (N_15898,N_15825,N_15828);
nor U15899 (N_15899,N_15747,N_15774);
or U15900 (N_15900,N_15749,N_15716);
and U15901 (N_15901,N_15761,N_15778);
and U15902 (N_15902,N_15799,N_15835);
nor U15903 (N_15903,N_15779,N_15720);
and U15904 (N_15904,N_15824,N_15754);
nand U15905 (N_15905,N_15695,N_15722);
nor U15906 (N_15906,N_15823,N_15833);
and U15907 (N_15907,N_15681,N_15815);
nor U15908 (N_15908,N_15801,N_15782);
and U15909 (N_15909,N_15791,N_15712);
and U15910 (N_15910,N_15781,N_15692);
and U15911 (N_15911,N_15719,N_15701);
nand U15912 (N_15912,N_15710,N_15753);
and U15913 (N_15913,N_15733,N_15727);
nor U15914 (N_15914,N_15790,N_15795);
nor U15915 (N_15915,N_15818,N_15702);
nor U15916 (N_15916,N_15711,N_15700);
and U15917 (N_15917,N_15682,N_15688);
nor U15918 (N_15918,N_15814,N_15805);
nor U15919 (N_15919,N_15796,N_15792);
nand U15920 (N_15920,N_15829,N_15682);
and U15921 (N_15921,N_15747,N_15734);
xor U15922 (N_15922,N_15684,N_15836);
nor U15923 (N_15923,N_15824,N_15773);
and U15924 (N_15924,N_15762,N_15759);
and U15925 (N_15925,N_15698,N_15798);
or U15926 (N_15926,N_15785,N_15819);
nand U15927 (N_15927,N_15694,N_15710);
nand U15928 (N_15928,N_15839,N_15831);
or U15929 (N_15929,N_15837,N_15829);
or U15930 (N_15930,N_15737,N_15750);
nor U15931 (N_15931,N_15808,N_15740);
nor U15932 (N_15932,N_15797,N_15827);
nor U15933 (N_15933,N_15780,N_15715);
xnor U15934 (N_15934,N_15691,N_15752);
nor U15935 (N_15935,N_15693,N_15796);
xnor U15936 (N_15936,N_15806,N_15782);
nor U15937 (N_15937,N_15742,N_15807);
nor U15938 (N_15938,N_15834,N_15767);
nand U15939 (N_15939,N_15750,N_15786);
xnor U15940 (N_15940,N_15724,N_15703);
and U15941 (N_15941,N_15781,N_15775);
and U15942 (N_15942,N_15819,N_15832);
nand U15943 (N_15943,N_15789,N_15753);
nand U15944 (N_15944,N_15796,N_15686);
nor U15945 (N_15945,N_15811,N_15743);
xor U15946 (N_15946,N_15776,N_15825);
and U15947 (N_15947,N_15718,N_15775);
nand U15948 (N_15948,N_15825,N_15815);
xnor U15949 (N_15949,N_15837,N_15809);
or U15950 (N_15950,N_15698,N_15687);
nand U15951 (N_15951,N_15823,N_15749);
or U15952 (N_15952,N_15784,N_15714);
nand U15953 (N_15953,N_15795,N_15767);
xnor U15954 (N_15954,N_15724,N_15750);
and U15955 (N_15955,N_15713,N_15695);
nand U15956 (N_15956,N_15690,N_15808);
or U15957 (N_15957,N_15683,N_15787);
xnor U15958 (N_15958,N_15722,N_15811);
and U15959 (N_15959,N_15786,N_15740);
nand U15960 (N_15960,N_15711,N_15689);
nand U15961 (N_15961,N_15816,N_15805);
and U15962 (N_15962,N_15717,N_15809);
xnor U15963 (N_15963,N_15699,N_15800);
nor U15964 (N_15964,N_15786,N_15819);
xnor U15965 (N_15965,N_15823,N_15739);
and U15966 (N_15966,N_15795,N_15738);
nand U15967 (N_15967,N_15797,N_15804);
and U15968 (N_15968,N_15791,N_15723);
xnor U15969 (N_15969,N_15717,N_15826);
and U15970 (N_15970,N_15698,N_15742);
nand U15971 (N_15971,N_15794,N_15681);
xnor U15972 (N_15972,N_15818,N_15718);
nand U15973 (N_15973,N_15775,N_15805);
or U15974 (N_15974,N_15793,N_15738);
nand U15975 (N_15975,N_15688,N_15745);
or U15976 (N_15976,N_15783,N_15820);
xnor U15977 (N_15977,N_15695,N_15708);
and U15978 (N_15978,N_15825,N_15769);
or U15979 (N_15979,N_15783,N_15767);
nand U15980 (N_15980,N_15738,N_15745);
and U15981 (N_15981,N_15817,N_15684);
nand U15982 (N_15982,N_15757,N_15704);
nor U15983 (N_15983,N_15682,N_15788);
and U15984 (N_15984,N_15768,N_15745);
and U15985 (N_15985,N_15687,N_15717);
and U15986 (N_15986,N_15794,N_15753);
nand U15987 (N_15987,N_15717,N_15686);
nand U15988 (N_15988,N_15721,N_15725);
or U15989 (N_15989,N_15740,N_15835);
or U15990 (N_15990,N_15772,N_15839);
nor U15991 (N_15991,N_15789,N_15762);
or U15992 (N_15992,N_15804,N_15814);
xnor U15993 (N_15993,N_15761,N_15725);
nor U15994 (N_15994,N_15833,N_15747);
and U15995 (N_15995,N_15808,N_15799);
nand U15996 (N_15996,N_15798,N_15728);
nor U15997 (N_15997,N_15795,N_15684);
xnor U15998 (N_15998,N_15734,N_15801);
or U15999 (N_15999,N_15748,N_15735);
xnor U16000 (N_16000,N_15846,N_15875);
and U16001 (N_16001,N_15944,N_15976);
and U16002 (N_16002,N_15862,N_15840);
nor U16003 (N_16003,N_15943,N_15909);
or U16004 (N_16004,N_15893,N_15969);
xnor U16005 (N_16005,N_15891,N_15866);
and U16006 (N_16006,N_15906,N_15973);
or U16007 (N_16007,N_15911,N_15988);
and U16008 (N_16008,N_15850,N_15952);
nand U16009 (N_16009,N_15900,N_15947);
nor U16010 (N_16010,N_15966,N_15902);
xor U16011 (N_16011,N_15908,N_15907);
and U16012 (N_16012,N_15852,N_15896);
xor U16013 (N_16013,N_15937,N_15917);
nor U16014 (N_16014,N_15945,N_15910);
and U16015 (N_16015,N_15935,N_15934);
or U16016 (N_16016,N_15956,N_15881);
nand U16017 (N_16017,N_15984,N_15958);
nand U16018 (N_16018,N_15953,N_15897);
xor U16019 (N_16019,N_15951,N_15904);
xnor U16020 (N_16020,N_15938,N_15992);
xor U16021 (N_16021,N_15977,N_15855);
nor U16022 (N_16022,N_15920,N_15861);
and U16023 (N_16023,N_15931,N_15844);
or U16024 (N_16024,N_15923,N_15962);
xnor U16025 (N_16025,N_15873,N_15925);
or U16026 (N_16026,N_15922,N_15949);
nor U16027 (N_16027,N_15874,N_15971);
or U16028 (N_16028,N_15843,N_15993);
nor U16029 (N_16029,N_15939,N_15946);
nor U16030 (N_16030,N_15880,N_15921);
or U16031 (N_16031,N_15954,N_15960);
nand U16032 (N_16032,N_15978,N_15974);
nand U16033 (N_16033,N_15885,N_15998);
and U16034 (N_16034,N_15851,N_15876);
nand U16035 (N_16035,N_15863,N_15932);
and U16036 (N_16036,N_15936,N_15916);
and U16037 (N_16037,N_15983,N_15868);
nor U16038 (N_16038,N_15869,N_15982);
nand U16039 (N_16039,N_15955,N_15886);
nand U16040 (N_16040,N_15865,N_15899);
and U16041 (N_16041,N_15895,N_15867);
and U16042 (N_16042,N_15887,N_15996);
or U16043 (N_16043,N_15905,N_15961);
and U16044 (N_16044,N_15871,N_15884);
nand U16045 (N_16045,N_15877,N_15980);
or U16046 (N_16046,N_15859,N_15898);
xnor U16047 (N_16047,N_15991,N_15959);
and U16048 (N_16048,N_15995,N_15933);
or U16049 (N_16049,N_15957,N_15990);
nor U16050 (N_16050,N_15964,N_15849);
or U16051 (N_16051,N_15942,N_15894);
nand U16052 (N_16052,N_15930,N_15975);
and U16053 (N_16053,N_15994,N_15882);
xor U16054 (N_16054,N_15989,N_15997);
xnor U16055 (N_16055,N_15903,N_15929);
xnor U16056 (N_16056,N_15914,N_15967);
xor U16057 (N_16057,N_15941,N_15872);
and U16058 (N_16058,N_15889,N_15965);
or U16059 (N_16059,N_15926,N_15972);
nor U16060 (N_16060,N_15963,N_15854);
and U16061 (N_16061,N_15948,N_15853);
nand U16062 (N_16062,N_15919,N_15857);
nand U16063 (N_16063,N_15847,N_15928);
nor U16064 (N_16064,N_15879,N_15878);
xor U16065 (N_16065,N_15860,N_15845);
and U16066 (N_16066,N_15856,N_15981);
and U16067 (N_16067,N_15918,N_15848);
xnor U16068 (N_16068,N_15970,N_15870);
nor U16069 (N_16069,N_15940,N_15915);
xnor U16070 (N_16070,N_15968,N_15979);
nor U16071 (N_16071,N_15842,N_15883);
nor U16072 (N_16072,N_15987,N_15892);
or U16073 (N_16073,N_15888,N_15924);
nor U16074 (N_16074,N_15999,N_15985);
and U16075 (N_16075,N_15986,N_15901);
nor U16076 (N_16076,N_15950,N_15927);
and U16077 (N_16077,N_15890,N_15858);
and U16078 (N_16078,N_15841,N_15864);
and U16079 (N_16079,N_15913,N_15912);
nand U16080 (N_16080,N_15976,N_15979);
or U16081 (N_16081,N_15898,N_15901);
xnor U16082 (N_16082,N_15974,N_15927);
nand U16083 (N_16083,N_15970,N_15966);
xor U16084 (N_16084,N_15938,N_15899);
and U16085 (N_16085,N_15973,N_15865);
nor U16086 (N_16086,N_15935,N_15998);
and U16087 (N_16087,N_15883,N_15898);
xor U16088 (N_16088,N_15862,N_15878);
or U16089 (N_16089,N_15969,N_15995);
nand U16090 (N_16090,N_15871,N_15974);
and U16091 (N_16091,N_15882,N_15934);
or U16092 (N_16092,N_15971,N_15937);
or U16093 (N_16093,N_15934,N_15869);
and U16094 (N_16094,N_15904,N_15957);
nor U16095 (N_16095,N_15868,N_15966);
or U16096 (N_16096,N_15938,N_15880);
nor U16097 (N_16097,N_15933,N_15904);
nand U16098 (N_16098,N_15989,N_15860);
xnor U16099 (N_16099,N_15860,N_15979);
nand U16100 (N_16100,N_15976,N_15865);
xnor U16101 (N_16101,N_15908,N_15905);
and U16102 (N_16102,N_15858,N_15917);
xor U16103 (N_16103,N_15984,N_15988);
or U16104 (N_16104,N_15933,N_15866);
nand U16105 (N_16105,N_15998,N_15863);
xnor U16106 (N_16106,N_15875,N_15911);
and U16107 (N_16107,N_15931,N_15976);
xor U16108 (N_16108,N_15844,N_15978);
nand U16109 (N_16109,N_15902,N_15912);
and U16110 (N_16110,N_15844,N_15990);
nor U16111 (N_16111,N_15948,N_15933);
nor U16112 (N_16112,N_15900,N_15907);
and U16113 (N_16113,N_15945,N_15912);
nand U16114 (N_16114,N_15880,N_15954);
nor U16115 (N_16115,N_15945,N_15957);
or U16116 (N_16116,N_15974,N_15963);
or U16117 (N_16117,N_15963,N_15939);
nor U16118 (N_16118,N_15979,N_15950);
and U16119 (N_16119,N_15880,N_15840);
nand U16120 (N_16120,N_15886,N_15935);
nor U16121 (N_16121,N_15868,N_15885);
and U16122 (N_16122,N_15966,N_15972);
xor U16123 (N_16123,N_15885,N_15982);
nor U16124 (N_16124,N_15982,N_15845);
nand U16125 (N_16125,N_15852,N_15843);
and U16126 (N_16126,N_15923,N_15958);
and U16127 (N_16127,N_15874,N_15882);
or U16128 (N_16128,N_15902,N_15995);
nor U16129 (N_16129,N_15914,N_15961);
nand U16130 (N_16130,N_15983,N_15866);
nand U16131 (N_16131,N_15874,N_15850);
and U16132 (N_16132,N_15849,N_15979);
xnor U16133 (N_16133,N_15918,N_15975);
and U16134 (N_16134,N_15965,N_15942);
nor U16135 (N_16135,N_15953,N_15985);
nor U16136 (N_16136,N_15963,N_15849);
and U16137 (N_16137,N_15864,N_15979);
xnor U16138 (N_16138,N_15857,N_15965);
xnor U16139 (N_16139,N_15856,N_15852);
nand U16140 (N_16140,N_15880,N_15870);
xor U16141 (N_16141,N_15848,N_15937);
xor U16142 (N_16142,N_15905,N_15953);
nor U16143 (N_16143,N_15931,N_15982);
nor U16144 (N_16144,N_15929,N_15956);
and U16145 (N_16145,N_15965,N_15970);
nand U16146 (N_16146,N_15853,N_15851);
and U16147 (N_16147,N_15865,N_15938);
nand U16148 (N_16148,N_15902,N_15989);
and U16149 (N_16149,N_15954,N_15977);
or U16150 (N_16150,N_15854,N_15986);
xor U16151 (N_16151,N_15994,N_15919);
nor U16152 (N_16152,N_15950,N_15878);
and U16153 (N_16153,N_15983,N_15941);
or U16154 (N_16154,N_15983,N_15877);
xnor U16155 (N_16155,N_15920,N_15950);
xor U16156 (N_16156,N_15999,N_15957);
or U16157 (N_16157,N_15879,N_15887);
or U16158 (N_16158,N_15904,N_15958);
and U16159 (N_16159,N_15847,N_15949);
xnor U16160 (N_16160,N_16102,N_16040);
nor U16161 (N_16161,N_16062,N_16046);
nor U16162 (N_16162,N_16012,N_16025);
nor U16163 (N_16163,N_16097,N_16071);
or U16164 (N_16164,N_16092,N_16089);
nand U16165 (N_16165,N_16056,N_16150);
xor U16166 (N_16166,N_16041,N_16005);
nand U16167 (N_16167,N_16120,N_16076);
nand U16168 (N_16168,N_16053,N_16103);
or U16169 (N_16169,N_16007,N_16134);
nand U16170 (N_16170,N_16079,N_16031);
nand U16171 (N_16171,N_16048,N_16125);
and U16172 (N_16172,N_16035,N_16152);
nor U16173 (N_16173,N_16110,N_16123);
or U16174 (N_16174,N_16075,N_16131);
nand U16175 (N_16175,N_16107,N_16118);
and U16176 (N_16176,N_16090,N_16157);
or U16177 (N_16177,N_16070,N_16009);
and U16178 (N_16178,N_16145,N_16060);
and U16179 (N_16179,N_16113,N_16006);
and U16180 (N_16180,N_16121,N_16112);
nor U16181 (N_16181,N_16117,N_16104);
nand U16182 (N_16182,N_16109,N_16032);
nor U16183 (N_16183,N_16140,N_16023);
or U16184 (N_16184,N_16036,N_16017);
nor U16185 (N_16185,N_16085,N_16133);
nand U16186 (N_16186,N_16149,N_16030);
nor U16187 (N_16187,N_16124,N_16051);
xnor U16188 (N_16188,N_16000,N_16037);
nor U16189 (N_16189,N_16135,N_16044);
and U16190 (N_16190,N_16014,N_16141);
or U16191 (N_16191,N_16115,N_16054);
nor U16192 (N_16192,N_16021,N_16015);
and U16193 (N_16193,N_16016,N_16156);
nor U16194 (N_16194,N_16073,N_16147);
and U16195 (N_16195,N_16047,N_16049);
xnor U16196 (N_16196,N_16010,N_16057);
or U16197 (N_16197,N_16126,N_16008);
and U16198 (N_16198,N_16100,N_16096);
xnor U16199 (N_16199,N_16142,N_16063);
or U16200 (N_16200,N_16029,N_16146);
or U16201 (N_16201,N_16072,N_16132);
nand U16202 (N_16202,N_16043,N_16039);
and U16203 (N_16203,N_16129,N_16106);
xnor U16204 (N_16204,N_16093,N_16078);
xor U16205 (N_16205,N_16052,N_16066);
nor U16206 (N_16206,N_16027,N_16004);
and U16207 (N_16207,N_16137,N_16022);
nor U16208 (N_16208,N_16154,N_16011);
nor U16209 (N_16209,N_16159,N_16116);
nand U16210 (N_16210,N_16069,N_16065);
nor U16211 (N_16211,N_16101,N_16158);
or U16212 (N_16212,N_16155,N_16026);
nand U16213 (N_16213,N_16081,N_16002);
xnor U16214 (N_16214,N_16080,N_16119);
xnor U16215 (N_16215,N_16086,N_16038);
and U16216 (N_16216,N_16018,N_16059);
nand U16217 (N_16217,N_16061,N_16024);
and U16218 (N_16218,N_16138,N_16095);
nand U16219 (N_16219,N_16001,N_16108);
nor U16220 (N_16220,N_16055,N_16151);
xor U16221 (N_16221,N_16148,N_16074);
and U16222 (N_16222,N_16094,N_16077);
nand U16223 (N_16223,N_16064,N_16128);
and U16224 (N_16224,N_16136,N_16098);
nand U16225 (N_16225,N_16144,N_16050);
nand U16226 (N_16226,N_16034,N_16067);
xnor U16227 (N_16227,N_16088,N_16042);
or U16228 (N_16228,N_16099,N_16082);
nor U16229 (N_16229,N_16033,N_16084);
and U16230 (N_16230,N_16019,N_16020);
or U16231 (N_16231,N_16028,N_16111);
or U16232 (N_16232,N_16013,N_16087);
nor U16233 (N_16233,N_16153,N_16003);
xor U16234 (N_16234,N_16130,N_16083);
and U16235 (N_16235,N_16143,N_16114);
and U16236 (N_16236,N_16058,N_16091);
and U16237 (N_16237,N_16139,N_16105);
nor U16238 (N_16238,N_16127,N_16045);
and U16239 (N_16239,N_16122,N_16068);
or U16240 (N_16240,N_16033,N_16021);
nor U16241 (N_16241,N_16062,N_16038);
nand U16242 (N_16242,N_16144,N_16104);
or U16243 (N_16243,N_16116,N_16016);
nor U16244 (N_16244,N_16063,N_16112);
nor U16245 (N_16245,N_16063,N_16069);
nand U16246 (N_16246,N_16003,N_16056);
xnor U16247 (N_16247,N_16045,N_16105);
or U16248 (N_16248,N_16068,N_16099);
nand U16249 (N_16249,N_16073,N_16103);
nor U16250 (N_16250,N_16060,N_16157);
and U16251 (N_16251,N_16075,N_16074);
nand U16252 (N_16252,N_16022,N_16106);
xnor U16253 (N_16253,N_16102,N_16063);
nor U16254 (N_16254,N_16119,N_16034);
nor U16255 (N_16255,N_16000,N_16007);
xor U16256 (N_16256,N_16022,N_16129);
nand U16257 (N_16257,N_16000,N_16112);
nand U16258 (N_16258,N_16003,N_16090);
nor U16259 (N_16259,N_16078,N_16083);
nor U16260 (N_16260,N_16095,N_16113);
nand U16261 (N_16261,N_16000,N_16097);
nor U16262 (N_16262,N_16042,N_16048);
nor U16263 (N_16263,N_16082,N_16017);
xnor U16264 (N_16264,N_16122,N_16044);
and U16265 (N_16265,N_16089,N_16001);
and U16266 (N_16266,N_16099,N_16111);
nand U16267 (N_16267,N_16029,N_16077);
and U16268 (N_16268,N_16107,N_16070);
nand U16269 (N_16269,N_16089,N_16058);
nand U16270 (N_16270,N_16051,N_16090);
nor U16271 (N_16271,N_16080,N_16134);
nand U16272 (N_16272,N_16098,N_16043);
or U16273 (N_16273,N_16095,N_16108);
nand U16274 (N_16274,N_16134,N_16123);
or U16275 (N_16275,N_16019,N_16057);
or U16276 (N_16276,N_16140,N_16093);
nor U16277 (N_16277,N_16008,N_16016);
nor U16278 (N_16278,N_16088,N_16102);
nand U16279 (N_16279,N_16032,N_16014);
or U16280 (N_16280,N_16101,N_16135);
and U16281 (N_16281,N_16012,N_16154);
or U16282 (N_16282,N_16066,N_16063);
xor U16283 (N_16283,N_16056,N_16087);
or U16284 (N_16284,N_16023,N_16128);
or U16285 (N_16285,N_16019,N_16120);
nor U16286 (N_16286,N_16069,N_16062);
nor U16287 (N_16287,N_16061,N_16118);
nand U16288 (N_16288,N_16042,N_16013);
xnor U16289 (N_16289,N_16050,N_16047);
or U16290 (N_16290,N_16073,N_16061);
nand U16291 (N_16291,N_16121,N_16088);
nor U16292 (N_16292,N_16090,N_16077);
xor U16293 (N_16293,N_16020,N_16154);
xor U16294 (N_16294,N_16104,N_16155);
nand U16295 (N_16295,N_16081,N_16033);
or U16296 (N_16296,N_16017,N_16130);
nor U16297 (N_16297,N_16078,N_16039);
or U16298 (N_16298,N_16121,N_16137);
and U16299 (N_16299,N_16134,N_16111);
or U16300 (N_16300,N_16118,N_16078);
nor U16301 (N_16301,N_16113,N_16136);
and U16302 (N_16302,N_16082,N_16009);
xnor U16303 (N_16303,N_16154,N_16048);
nor U16304 (N_16304,N_16131,N_16104);
xnor U16305 (N_16305,N_16069,N_16120);
and U16306 (N_16306,N_16095,N_16096);
nand U16307 (N_16307,N_16114,N_16042);
xnor U16308 (N_16308,N_16035,N_16087);
or U16309 (N_16309,N_16101,N_16119);
nand U16310 (N_16310,N_16006,N_16099);
nand U16311 (N_16311,N_16107,N_16018);
and U16312 (N_16312,N_16013,N_16107);
xnor U16313 (N_16313,N_16060,N_16044);
nor U16314 (N_16314,N_16117,N_16085);
nand U16315 (N_16315,N_16083,N_16119);
nor U16316 (N_16316,N_16136,N_16100);
or U16317 (N_16317,N_16070,N_16044);
or U16318 (N_16318,N_16005,N_16087);
nor U16319 (N_16319,N_16134,N_16052);
or U16320 (N_16320,N_16163,N_16313);
nand U16321 (N_16321,N_16261,N_16200);
nor U16322 (N_16322,N_16224,N_16289);
and U16323 (N_16323,N_16298,N_16260);
and U16324 (N_16324,N_16254,N_16236);
xnor U16325 (N_16325,N_16197,N_16170);
and U16326 (N_16326,N_16228,N_16317);
nand U16327 (N_16327,N_16221,N_16262);
and U16328 (N_16328,N_16217,N_16251);
nor U16329 (N_16329,N_16166,N_16250);
or U16330 (N_16330,N_16280,N_16288);
xor U16331 (N_16331,N_16291,N_16245);
xnor U16332 (N_16332,N_16227,N_16173);
or U16333 (N_16333,N_16192,N_16177);
or U16334 (N_16334,N_16306,N_16165);
and U16335 (N_16335,N_16316,N_16161);
nor U16336 (N_16336,N_16293,N_16269);
xor U16337 (N_16337,N_16273,N_16212);
xnor U16338 (N_16338,N_16259,N_16203);
or U16339 (N_16339,N_16241,N_16300);
and U16340 (N_16340,N_16219,N_16171);
or U16341 (N_16341,N_16249,N_16222);
nand U16342 (N_16342,N_16213,N_16215);
nor U16343 (N_16343,N_16195,N_16230);
and U16344 (N_16344,N_16169,N_16193);
and U16345 (N_16345,N_16270,N_16266);
or U16346 (N_16346,N_16202,N_16238);
or U16347 (N_16347,N_16234,N_16319);
or U16348 (N_16348,N_16244,N_16253);
nand U16349 (N_16349,N_16168,N_16223);
and U16350 (N_16350,N_16174,N_16231);
nand U16351 (N_16351,N_16232,N_16233);
or U16352 (N_16352,N_16247,N_16276);
nand U16353 (N_16353,N_16264,N_16308);
nand U16354 (N_16354,N_16175,N_16211);
nor U16355 (N_16355,N_16257,N_16310);
or U16356 (N_16356,N_16242,N_16204);
and U16357 (N_16357,N_16229,N_16243);
xor U16358 (N_16358,N_16210,N_16307);
xor U16359 (N_16359,N_16256,N_16299);
xor U16360 (N_16360,N_16305,N_16178);
nor U16361 (N_16361,N_16272,N_16278);
and U16362 (N_16362,N_16181,N_16297);
or U16363 (N_16363,N_16235,N_16252);
or U16364 (N_16364,N_16201,N_16277);
and U16365 (N_16365,N_16216,N_16176);
and U16366 (N_16366,N_16196,N_16239);
xor U16367 (N_16367,N_16258,N_16189);
nand U16368 (N_16368,N_16290,N_16208);
xor U16369 (N_16369,N_16295,N_16162);
and U16370 (N_16370,N_16198,N_16218);
nand U16371 (N_16371,N_16265,N_16286);
nor U16372 (N_16372,N_16206,N_16281);
nor U16373 (N_16373,N_16185,N_16315);
and U16374 (N_16374,N_16314,N_16186);
nand U16375 (N_16375,N_16191,N_16302);
nor U16376 (N_16376,N_16303,N_16268);
and U16377 (N_16377,N_16292,N_16183);
nor U16378 (N_16378,N_16167,N_16309);
xnor U16379 (N_16379,N_16214,N_16225);
nand U16380 (N_16380,N_16246,N_16240);
and U16381 (N_16381,N_16184,N_16205);
or U16382 (N_16382,N_16207,N_16267);
and U16383 (N_16383,N_16199,N_16179);
nand U16384 (N_16384,N_16180,N_16279);
xor U16385 (N_16385,N_16220,N_16275);
or U16386 (N_16386,N_16164,N_16188);
or U16387 (N_16387,N_16287,N_16285);
or U16388 (N_16388,N_16282,N_16263);
xnor U16389 (N_16389,N_16182,N_16301);
and U16390 (N_16390,N_16283,N_16312);
xor U16391 (N_16391,N_16311,N_16209);
nor U16392 (N_16392,N_16294,N_16190);
nand U16393 (N_16393,N_16255,N_16237);
nand U16394 (N_16394,N_16284,N_16194);
nand U16395 (N_16395,N_16160,N_16318);
or U16396 (N_16396,N_16296,N_16172);
nand U16397 (N_16397,N_16274,N_16187);
or U16398 (N_16398,N_16226,N_16248);
and U16399 (N_16399,N_16271,N_16304);
and U16400 (N_16400,N_16260,N_16239);
or U16401 (N_16401,N_16261,N_16299);
or U16402 (N_16402,N_16255,N_16288);
xnor U16403 (N_16403,N_16263,N_16254);
nand U16404 (N_16404,N_16309,N_16206);
nor U16405 (N_16405,N_16212,N_16306);
nor U16406 (N_16406,N_16230,N_16201);
xnor U16407 (N_16407,N_16246,N_16186);
and U16408 (N_16408,N_16210,N_16219);
and U16409 (N_16409,N_16298,N_16274);
and U16410 (N_16410,N_16293,N_16229);
or U16411 (N_16411,N_16257,N_16194);
or U16412 (N_16412,N_16191,N_16236);
nand U16413 (N_16413,N_16168,N_16263);
nor U16414 (N_16414,N_16177,N_16201);
nor U16415 (N_16415,N_16247,N_16167);
nor U16416 (N_16416,N_16206,N_16169);
nor U16417 (N_16417,N_16289,N_16238);
and U16418 (N_16418,N_16306,N_16315);
nor U16419 (N_16419,N_16268,N_16186);
or U16420 (N_16420,N_16265,N_16193);
and U16421 (N_16421,N_16253,N_16265);
or U16422 (N_16422,N_16189,N_16194);
xnor U16423 (N_16423,N_16169,N_16226);
nand U16424 (N_16424,N_16249,N_16318);
xor U16425 (N_16425,N_16263,N_16269);
or U16426 (N_16426,N_16316,N_16228);
xor U16427 (N_16427,N_16300,N_16206);
nor U16428 (N_16428,N_16260,N_16201);
or U16429 (N_16429,N_16291,N_16163);
nand U16430 (N_16430,N_16262,N_16194);
nand U16431 (N_16431,N_16264,N_16190);
and U16432 (N_16432,N_16200,N_16289);
nand U16433 (N_16433,N_16240,N_16280);
nand U16434 (N_16434,N_16201,N_16246);
nor U16435 (N_16435,N_16257,N_16217);
nor U16436 (N_16436,N_16170,N_16277);
xnor U16437 (N_16437,N_16227,N_16273);
xnor U16438 (N_16438,N_16311,N_16217);
nor U16439 (N_16439,N_16291,N_16247);
and U16440 (N_16440,N_16242,N_16180);
or U16441 (N_16441,N_16186,N_16294);
nor U16442 (N_16442,N_16218,N_16267);
nor U16443 (N_16443,N_16178,N_16170);
and U16444 (N_16444,N_16205,N_16211);
nand U16445 (N_16445,N_16273,N_16263);
or U16446 (N_16446,N_16166,N_16256);
nor U16447 (N_16447,N_16226,N_16241);
nand U16448 (N_16448,N_16295,N_16301);
xor U16449 (N_16449,N_16222,N_16244);
nor U16450 (N_16450,N_16249,N_16252);
nand U16451 (N_16451,N_16303,N_16286);
nor U16452 (N_16452,N_16274,N_16271);
or U16453 (N_16453,N_16190,N_16183);
nor U16454 (N_16454,N_16206,N_16164);
and U16455 (N_16455,N_16166,N_16229);
and U16456 (N_16456,N_16194,N_16308);
nor U16457 (N_16457,N_16198,N_16260);
nand U16458 (N_16458,N_16164,N_16219);
and U16459 (N_16459,N_16232,N_16218);
nand U16460 (N_16460,N_16278,N_16183);
or U16461 (N_16461,N_16274,N_16161);
xnor U16462 (N_16462,N_16278,N_16287);
or U16463 (N_16463,N_16163,N_16185);
nand U16464 (N_16464,N_16311,N_16272);
nor U16465 (N_16465,N_16253,N_16298);
nor U16466 (N_16466,N_16253,N_16300);
and U16467 (N_16467,N_16175,N_16191);
and U16468 (N_16468,N_16180,N_16225);
xor U16469 (N_16469,N_16286,N_16280);
or U16470 (N_16470,N_16236,N_16287);
nand U16471 (N_16471,N_16222,N_16269);
and U16472 (N_16472,N_16226,N_16216);
and U16473 (N_16473,N_16218,N_16264);
or U16474 (N_16474,N_16276,N_16240);
nand U16475 (N_16475,N_16209,N_16192);
and U16476 (N_16476,N_16312,N_16178);
nor U16477 (N_16477,N_16280,N_16312);
xor U16478 (N_16478,N_16317,N_16184);
xnor U16479 (N_16479,N_16276,N_16194);
and U16480 (N_16480,N_16332,N_16347);
nor U16481 (N_16481,N_16384,N_16460);
nand U16482 (N_16482,N_16390,N_16476);
and U16483 (N_16483,N_16325,N_16425);
and U16484 (N_16484,N_16399,N_16404);
or U16485 (N_16485,N_16455,N_16328);
or U16486 (N_16486,N_16381,N_16335);
and U16487 (N_16487,N_16364,N_16477);
or U16488 (N_16488,N_16433,N_16416);
nand U16489 (N_16489,N_16360,N_16383);
nand U16490 (N_16490,N_16453,N_16427);
xor U16491 (N_16491,N_16379,N_16418);
nor U16492 (N_16492,N_16344,N_16391);
nor U16493 (N_16493,N_16422,N_16447);
or U16494 (N_16494,N_16351,N_16397);
and U16495 (N_16495,N_16368,N_16380);
and U16496 (N_16496,N_16388,N_16446);
or U16497 (N_16497,N_16346,N_16412);
xor U16498 (N_16498,N_16378,N_16471);
nor U16499 (N_16499,N_16345,N_16444);
and U16500 (N_16500,N_16428,N_16322);
or U16501 (N_16501,N_16323,N_16366);
nand U16502 (N_16502,N_16452,N_16343);
xnor U16503 (N_16503,N_16372,N_16459);
nor U16504 (N_16504,N_16326,N_16324);
or U16505 (N_16505,N_16406,N_16367);
nor U16506 (N_16506,N_16359,N_16415);
and U16507 (N_16507,N_16400,N_16336);
or U16508 (N_16508,N_16479,N_16348);
xor U16509 (N_16509,N_16411,N_16468);
and U16510 (N_16510,N_16417,N_16478);
and U16511 (N_16511,N_16407,N_16363);
xnor U16512 (N_16512,N_16334,N_16321);
xor U16513 (N_16513,N_16421,N_16450);
and U16514 (N_16514,N_16337,N_16438);
or U16515 (N_16515,N_16475,N_16375);
or U16516 (N_16516,N_16474,N_16405);
nor U16517 (N_16517,N_16426,N_16442);
xor U16518 (N_16518,N_16410,N_16393);
xnor U16519 (N_16519,N_16401,N_16365);
nand U16520 (N_16520,N_16464,N_16386);
or U16521 (N_16521,N_16466,N_16333);
nand U16522 (N_16522,N_16439,N_16362);
or U16523 (N_16523,N_16402,N_16409);
or U16524 (N_16524,N_16419,N_16408);
and U16525 (N_16525,N_16445,N_16472);
or U16526 (N_16526,N_16461,N_16361);
nor U16527 (N_16527,N_16420,N_16430);
and U16528 (N_16528,N_16467,N_16358);
and U16529 (N_16529,N_16354,N_16385);
nand U16530 (N_16530,N_16432,N_16424);
nor U16531 (N_16531,N_16456,N_16440);
and U16532 (N_16532,N_16436,N_16437);
and U16533 (N_16533,N_16395,N_16457);
nand U16534 (N_16534,N_16377,N_16376);
nand U16535 (N_16535,N_16448,N_16353);
nand U16536 (N_16536,N_16394,N_16462);
or U16537 (N_16537,N_16352,N_16374);
and U16538 (N_16538,N_16389,N_16355);
xnor U16539 (N_16539,N_16443,N_16357);
xor U16540 (N_16540,N_16449,N_16434);
nand U16541 (N_16541,N_16330,N_16398);
and U16542 (N_16542,N_16465,N_16429);
or U16543 (N_16543,N_16369,N_16340);
or U16544 (N_16544,N_16463,N_16441);
and U16545 (N_16545,N_16396,N_16327);
nand U16546 (N_16546,N_16329,N_16469);
nor U16547 (N_16547,N_16339,N_16341);
nand U16548 (N_16548,N_16451,N_16356);
xnor U16549 (N_16549,N_16431,N_16320);
or U16550 (N_16550,N_16387,N_16473);
or U16551 (N_16551,N_16413,N_16331);
or U16552 (N_16552,N_16470,N_16370);
or U16553 (N_16553,N_16423,N_16342);
nor U16554 (N_16554,N_16338,N_16454);
nand U16555 (N_16555,N_16373,N_16403);
and U16556 (N_16556,N_16349,N_16392);
nor U16557 (N_16557,N_16458,N_16414);
and U16558 (N_16558,N_16371,N_16435);
or U16559 (N_16559,N_16350,N_16382);
nor U16560 (N_16560,N_16466,N_16454);
xnor U16561 (N_16561,N_16449,N_16414);
nor U16562 (N_16562,N_16430,N_16419);
nor U16563 (N_16563,N_16459,N_16436);
or U16564 (N_16564,N_16358,N_16331);
nor U16565 (N_16565,N_16396,N_16353);
xnor U16566 (N_16566,N_16446,N_16453);
nand U16567 (N_16567,N_16470,N_16388);
xnor U16568 (N_16568,N_16326,N_16362);
xor U16569 (N_16569,N_16444,N_16431);
or U16570 (N_16570,N_16407,N_16409);
and U16571 (N_16571,N_16478,N_16368);
and U16572 (N_16572,N_16416,N_16474);
xor U16573 (N_16573,N_16468,N_16342);
nor U16574 (N_16574,N_16432,N_16406);
or U16575 (N_16575,N_16473,N_16370);
and U16576 (N_16576,N_16333,N_16407);
or U16577 (N_16577,N_16341,N_16349);
xor U16578 (N_16578,N_16474,N_16408);
nor U16579 (N_16579,N_16378,N_16394);
xnor U16580 (N_16580,N_16413,N_16430);
and U16581 (N_16581,N_16369,N_16417);
xor U16582 (N_16582,N_16467,N_16396);
and U16583 (N_16583,N_16397,N_16467);
nor U16584 (N_16584,N_16379,N_16434);
nand U16585 (N_16585,N_16351,N_16453);
xnor U16586 (N_16586,N_16467,N_16436);
nor U16587 (N_16587,N_16456,N_16356);
nor U16588 (N_16588,N_16469,N_16412);
and U16589 (N_16589,N_16396,N_16325);
xnor U16590 (N_16590,N_16460,N_16358);
or U16591 (N_16591,N_16399,N_16405);
nand U16592 (N_16592,N_16441,N_16446);
and U16593 (N_16593,N_16384,N_16477);
nand U16594 (N_16594,N_16377,N_16334);
nor U16595 (N_16595,N_16340,N_16355);
nor U16596 (N_16596,N_16342,N_16366);
or U16597 (N_16597,N_16418,N_16340);
or U16598 (N_16598,N_16443,N_16447);
xor U16599 (N_16599,N_16478,N_16347);
xnor U16600 (N_16600,N_16402,N_16417);
or U16601 (N_16601,N_16323,N_16430);
or U16602 (N_16602,N_16377,N_16460);
or U16603 (N_16603,N_16394,N_16372);
nor U16604 (N_16604,N_16392,N_16382);
and U16605 (N_16605,N_16459,N_16357);
and U16606 (N_16606,N_16362,N_16365);
xnor U16607 (N_16607,N_16407,N_16399);
or U16608 (N_16608,N_16467,N_16447);
xnor U16609 (N_16609,N_16462,N_16439);
nor U16610 (N_16610,N_16423,N_16358);
xnor U16611 (N_16611,N_16327,N_16380);
and U16612 (N_16612,N_16374,N_16419);
and U16613 (N_16613,N_16381,N_16385);
nor U16614 (N_16614,N_16371,N_16329);
or U16615 (N_16615,N_16478,N_16364);
nor U16616 (N_16616,N_16431,N_16398);
or U16617 (N_16617,N_16396,N_16416);
nor U16618 (N_16618,N_16374,N_16433);
nand U16619 (N_16619,N_16368,N_16383);
nand U16620 (N_16620,N_16450,N_16340);
or U16621 (N_16621,N_16325,N_16442);
and U16622 (N_16622,N_16432,N_16379);
xor U16623 (N_16623,N_16320,N_16422);
and U16624 (N_16624,N_16366,N_16405);
and U16625 (N_16625,N_16429,N_16437);
or U16626 (N_16626,N_16375,N_16434);
nor U16627 (N_16627,N_16349,N_16353);
and U16628 (N_16628,N_16437,N_16394);
nor U16629 (N_16629,N_16387,N_16425);
xor U16630 (N_16630,N_16363,N_16353);
xnor U16631 (N_16631,N_16416,N_16467);
xor U16632 (N_16632,N_16336,N_16399);
nand U16633 (N_16633,N_16329,N_16461);
and U16634 (N_16634,N_16351,N_16464);
nor U16635 (N_16635,N_16382,N_16439);
and U16636 (N_16636,N_16469,N_16365);
or U16637 (N_16637,N_16400,N_16443);
xnor U16638 (N_16638,N_16421,N_16331);
nor U16639 (N_16639,N_16323,N_16406);
xor U16640 (N_16640,N_16573,N_16527);
xor U16641 (N_16641,N_16556,N_16605);
xnor U16642 (N_16642,N_16507,N_16518);
xor U16643 (N_16643,N_16628,N_16524);
and U16644 (N_16644,N_16617,N_16530);
nor U16645 (N_16645,N_16516,N_16503);
nor U16646 (N_16646,N_16623,N_16538);
and U16647 (N_16647,N_16522,N_16619);
nand U16648 (N_16648,N_16509,N_16523);
nand U16649 (N_16649,N_16569,N_16580);
nor U16650 (N_16650,N_16563,N_16627);
nand U16651 (N_16651,N_16633,N_16560);
nor U16652 (N_16652,N_16635,N_16535);
and U16653 (N_16653,N_16570,N_16621);
and U16654 (N_16654,N_16618,N_16597);
or U16655 (N_16655,N_16528,N_16636);
nor U16656 (N_16656,N_16547,N_16615);
nor U16657 (N_16657,N_16497,N_16484);
and U16658 (N_16658,N_16625,N_16486);
nand U16659 (N_16659,N_16504,N_16561);
nand U16660 (N_16660,N_16572,N_16493);
and U16661 (N_16661,N_16506,N_16499);
xnor U16662 (N_16662,N_16584,N_16548);
nand U16663 (N_16663,N_16579,N_16488);
nand U16664 (N_16664,N_16559,N_16554);
and U16665 (N_16665,N_16578,N_16490);
nor U16666 (N_16666,N_16510,N_16517);
xnor U16667 (N_16667,N_16541,N_16600);
nor U16668 (N_16668,N_16552,N_16574);
or U16669 (N_16669,N_16601,N_16564);
nor U16670 (N_16670,N_16520,N_16602);
xnor U16671 (N_16671,N_16609,N_16622);
xnor U16672 (N_16672,N_16614,N_16495);
nand U16673 (N_16673,N_16620,N_16582);
or U16674 (N_16674,N_16502,N_16604);
nor U16675 (N_16675,N_16492,N_16546);
xor U16676 (N_16676,N_16611,N_16483);
nor U16677 (N_16677,N_16557,N_16610);
nor U16678 (N_16678,N_16526,N_16489);
nand U16679 (N_16679,N_16632,N_16592);
nand U16680 (N_16680,N_16500,N_16514);
and U16681 (N_16681,N_16629,N_16501);
or U16682 (N_16682,N_16515,N_16529);
nor U16683 (N_16683,N_16599,N_16568);
xnor U16684 (N_16684,N_16511,N_16613);
or U16685 (N_16685,N_16575,N_16630);
nand U16686 (N_16686,N_16505,N_16496);
nand U16687 (N_16687,N_16626,N_16612);
nand U16688 (N_16688,N_16525,N_16487);
and U16689 (N_16689,N_16482,N_16577);
nor U16690 (N_16690,N_16551,N_16550);
xnor U16691 (N_16691,N_16512,N_16540);
xor U16692 (N_16692,N_16607,N_16591);
or U16693 (N_16693,N_16596,N_16594);
nand U16694 (N_16694,N_16587,N_16586);
nand U16695 (N_16695,N_16549,N_16598);
nor U16696 (N_16696,N_16603,N_16536);
and U16697 (N_16697,N_16553,N_16606);
nor U16698 (N_16698,N_16637,N_16519);
nor U16699 (N_16699,N_16571,N_16485);
and U16700 (N_16700,N_16537,N_16565);
or U16701 (N_16701,N_16545,N_16491);
and U16702 (N_16702,N_16631,N_16576);
or U16703 (N_16703,N_16624,N_16585);
and U16704 (N_16704,N_16639,N_16567);
xor U16705 (N_16705,N_16542,N_16558);
and U16706 (N_16706,N_16539,N_16588);
and U16707 (N_16707,N_16616,N_16595);
xor U16708 (N_16708,N_16543,N_16481);
nand U16709 (N_16709,N_16566,N_16531);
nand U16710 (N_16710,N_16494,N_16583);
nor U16711 (N_16711,N_16533,N_16534);
nand U16712 (N_16712,N_16521,N_16634);
or U16713 (N_16713,N_16589,N_16608);
xor U16714 (N_16714,N_16593,N_16508);
xnor U16715 (N_16715,N_16532,N_16590);
and U16716 (N_16716,N_16562,N_16480);
and U16717 (N_16717,N_16581,N_16498);
xor U16718 (N_16718,N_16513,N_16555);
and U16719 (N_16719,N_16544,N_16638);
nor U16720 (N_16720,N_16536,N_16556);
nand U16721 (N_16721,N_16522,N_16581);
nor U16722 (N_16722,N_16542,N_16488);
and U16723 (N_16723,N_16508,N_16553);
or U16724 (N_16724,N_16602,N_16513);
and U16725 (N_16725,N_16482,N_16565);
or U16726 (N_16726,N_16544,N_16580);
or U16727 (N_16727,N_16590,N_16597);
xnor U16728 (N_16728,N_16508,N_16521);
nand U16729 (N_16729,N_16530,N_16552);
nor U16730 (N_16730,N_16548,N_16536);
and U16731 (N_16731,N_16587,N_16637);
and U16732 (N_16732,N_16551,N_16516);
nor U16733 (N_16733,N_16627,N_16623);
nand U16734 (N_16734,N_16557,N_16628);
and U16735 (N_16735,N_16482,N_16541);
xnor U16736 (N_16736,N_16549,N_16514);
or U16737 (N_16737,N_16568,N_16580);
or U16738 (N_16738,N_16564,N_16536);
nand U16739 (N_16739,N_16524,N_16590);
or U16740 (N_16740,N_16570,N_16634);
nand U16741 (N_16741,N_16486,N_16611);
xnor U16742 (N_16742,N_16630,N_16553);
or U16743 (N_16743,N_16548,N_16487);
nand U16744 (N_16744,N_16553,N_16516);
xnor U16745 (N_16745,N_16634,N_16617);
and U16746 (N_16746,N_16595,N_16487);
nand U16747 (N_16747,N_16634,N_16592);
nand U16748 (N_16748,N_16574,N_16606);
nor U16749 (N_16749,N_16506,N_16623);
or U16750 (N_16750,N_16589,N_16587);
and U16751 (N_16751,N_16497,N_16594);
nand U16752 (N_16752,N_16610,N_16622);
or U16753 (N_16753,N_16626,N_16577);
and U16754 (N_16754,N_16547,N_16528);
or U16755 (N_16755,N_16493,N_16505);
and U16756 (N_16756,N_16481,N_16594);
nand U16757 (N_16757,N_16514,N_16623);
nor U16758 (N_16758,N_16485,N_16583);
nor U16759 (N_16759,N_16565,N_16610);
or U16760 (N_16760,N_16586,N_16494);
xor U16761 (N_16761,N_16611,N_16577);
or U16762 (N_16762,N_16483,N_16538);
nand U16763 (N_16763,N_16623,N_16523);
nor U16764 (N_16764,N_16500,N_16523);
xor U16765 (N_16765,N_16614,N_16572);
and U16766 (N_16766,N_16492,N_16566);
nor U16767 (N_16767,N_16600,N_16631);
nor U16768 (N_16768,N_16595,N_16618);
xnor U16769 (N_16769,N_16551,N_16577);
nor U16770 (N_16770,N_16631,N_16540);
or U16771 (N_16771,N_16590,N_16604);
or U16772 (N_16772,N_16628,N_16547);
and U16773 (N_16773,N_16520,N_16544);
xnor U16774 (N_16774,N_16589,N_16583);
nor U16775 (N_16775,N_16567,N_16544);
xor U16776 (N_16776,N_16555,N_16484);
xnor U16777 (N_16777,N_16635,N_16501);
xnor U16778 (N_16778,N_16511,N_16630);
and U16779 (N_16779,N_16617,N_16618);
nand U16780 (N_16780,N_16544,N_16557);
or U16781 (N_16781,N_16582,N_16544);
or U16782 (N_16782,N_16608,N_16547);
nand U16783 (N_16783,N_16487,N_16577);
and U16784 (N_16784,N_16527,N_16634);
nand U16785 (N_16785,N_16599,N_16609);
xor U16786 (N_16786,N_16499,N_16547);
nor U16787 (N_16787,N_16501,N_16486);
xnor U16788 (N_16788,N_16512,N_16485);
nand U16789 (N_16789,N_16605,N_16541);
xnor U16790 (N_16790,N_16582,N_16610);
nand U16791 (N_16791,N_16507,N_16613);
nor U16792 (N_16792,N_16507,N_16584);
nor U16793 (N_16793,N_16518,N_16590);
nand U16794 (N_16794,N_16590,N_16625);
nand U16795 (N_16795,N_16574,N_16495);
or U16796 (N_16796,N_16532,N_16507);
nand U16797 (N_16797,N_16534,N_16491);
xnor U16798 (N_16798,N_16520,N_16576);
xor U16799 (N_16799,N_16501,N_16565);
nand U16800 (N_16800,N_16769,N_16732);
nor U16801 (N_16801,N_16796,N_16641);
nand U16802 (N_16802,N_16761,N_16655);
xor U16803 (N_16803,N_16750,N_16798);
or U16804 (N_16804,N_16702,N_16661);
and U16805 (N_16805,N_16731,N_16680);
xor U16806 (N_16806,N_16727,N_16674);
and U16807 (N_16807,N_16682,N_16756);
nor U16808 (N_16808,N_16724,N_16671);
and U16809 (N_16809,N_16772,N_16746);
nor U16810 (N_16810,N_16691,N_16667);
or U16811 (N_16811,N_16701,N_16759);
or U16812 (N_16812,N_16718,N_16757);
and U16813 (N_16813,N_16766,N_16686);
or U16814 (N_16814,N_16660,N_16743);
nor U16815 (N_16815,N_16696,N_16747);
and U16816 (N_16816,N_16733,N_16687);
xnor U16817 (N_16817,N_16668,N_16797);
nor U16818 (N_16818,N_16762,N_16765);
or U16819 (N_16819,N_16744,N_16665);
and U16820 (N_16820,N_16659,N_16705);
nand U16821 (N_16821,N_16782,N_16719);
xor U16822 (N_16822,N_16740,N_16758);
nand U16823 (N_16823,N_16640,N_16739);
nand U16824 (N_16824,N_16737,N_16730);
nor U16825 (N_16825,N_16794,N_16721);
or U16826 (N_16826,N_16684,N_16642);
nand U16827 (N_16827,N_16692,N_16664);
nor U16828 (N_16828,N_16799,N_16754);
or U16829 (N_16829,N_16658,N_16678);
xor U16830 (N_16830,N_16710,N_16676);
xnor U16831 (N_16831,N_16646,N_16726);
xnor U16832 (N_16832,N_16690,N_16722);
xor U16833 (N_16833,N_16698,N_16657);
nor U16834 (N_16834,N_16697,N_16753);
and U16835 (N_16835,N_16669,N_16656);
xnor U16836 (N_16836,N_16749,N_16653);
or U16837 (N_16837,N_16677,N_16654);
nand U16838 (N_16838,N_16780,N_16688);
nand U16839 (N_16839,N_16742,N_16777);
xor U16840 (N_16840,N_16683,N_16695);
or U16841 (N_16841,N_16707,N_16652);
nor U16842 (N_16842,N_16784,N_16751);
nor U16843 (N_16843,N_16781,N_16649);
nor U16844 (N_16844,N_16778,N_16666);
or U16845 (N_16845,N_16760,N_16725);
xor U16846 (N_16846,N_16789,N_16770);
or U16847 (N_16847,N_16716,N_16648);
and U16848 (N_16848,N_16788,N_16786);
nand U16849 (N_16849,N_16767,N_16755);
xor U16850 (N_16850,N_16679,N_16768);
or U16851 (N_16851,N_16706,N_16709);
xor U16852 (N_16852,N_16787,N_16715);
and U16853 (N_16853,N_16675,N_16795);
and U16854 (N_16854,N_16700,N_16734);
and U16855 (N_16855,N_16693,N_16694);
nand U16856 (N_16856,N_16793,N_16738);
and U16857 (N_16857,N_16672,N_16651);
and U16858 (N_16858,N_16714,N_16704);
nor U16859 (N_16859,N_16779,N_16764);
nor U16860 (N_16860,N_16708,N_16663);
and U16861 (N_16861,N_16763,N_16729);
xor U16862 (N_16862,N_16790,N_16685);
or U16863 (N_16863,N_16775,N_16703);
nand U16864 (N_16864,N_16792,N_16785);
or U16865 (N_16865,N_16712,N_16773);
or U16866 (N_16866,N_16791,N_16647);
nand U16867 (N_16867,N_16776,N_16643);
or U16868 (N_16868,N_16720,N_16681);
xnor U16869 (N_16869,N_16748,N_16774);
nor U16870 (N_16870,N_16644,N_16752);
or U16871 (N_16871,N_16745,N_16736);
nand U16872 (N_16872,N_16717,N_16723);
and U16873 (N_16873,N_16783,N_16645);
xnor U16874 (N_16874,N_16670,N_16662);
and U16875 (N_16875,N_16650,N_16713);
and U16876 (N_16876,N_16741,N_16699);
nor U16877 (N_16877,N_16728,N_16673);
or U16878 (N_16878,N_16735,N_16771);
nor U16879 (N_16879,N_16689,N_16711);
or U16880 (N_16880,N_16648,N_16661);
and U16881 (N_16881,N_16676,N_16648);
xnor U16882 (N_16882,N_16666,N_16670);
and U16883 (N_16883,N_16669,N_16780);
nor U16884 (N_16884,N_16771,N_16758);
or U16885 (N_16885,N_16716,N_16679);
or U16886 (N_16886,N_16790,N_16707);
or U16887 (N_16887,N_16691,N_16720);
or U16888 (N_16888,N_16717,N_16766);
xor U16889 (N_16889,N_16749,N_16738);
nor U16890 (N_16890,N_16781,N_16732);
and U16891 (N_16891,N_16782,N_16665);
and U16892 (N_16892,N_16734,N_16777);
xor U16893 (N_16893,N_16762,N_16645);
nand U16894 (N_16894,N_16733,N_16646);
or U16895 (N_16895,N_16797,N_16673);
nand U16896 (N_16896,N_16737,N_16713);
and U16897 (N_16897,N_16676,N_16788);
and U16898 (N_16898,N_16647,N_16752);
xnor U16899 (N_16899,N_16748,N_16705);
nor U16900 (N_16900,N_16676,N_16799);
and U16901 (N_16901,N_16756,N_16717);
and U16902 (N_16902,N_16767,N_16717);
nor U16903 (N_16903,N_16772,N_16728);
or U16904 (N_16904,N_16665,N_16769);
and U16905 (N_16905,N_16703,N_16757);
nor U16906 (N_16906,N_16746,N_16655);
nand U16907 (N_16907,N_16710,N_16728);
nor U16908 (N_16908,N_16736,N_16719);
nand U16909 (N_16909,N_16736,N_16667);
nand U16910 (N_16910,N_16736,N_16716);
nand U16911 (N_16911,N_16765,N_16696);
and U16912 (N_16912,N_16781,N_16763);
xor U16913 (N_16913,N_16643,N_16703);
or U16914 (N_16914,N_16720,N_16645);
nor U16915 (N_16915,N_16768,N_16675);
and U16916 (N_16916,N_16756,N_16643);
xor U16917 (N_16917,N_16702,N_16689);
nand U16918 (N_16918,N_16662,N_16640);
xnor U16919 (N_16919,N_16732,N_16664);
nand U16920 (N_16920,N_16679,N_16758);
nor U16921 (N_16921,N_16778,N_16752);
nor U16922 (N_16922,N_16657,N_16712);
xnor U16923 (N_16923,N_16644,N_16731);
xor U16924 (N_16924,N_16782,N_16684);
or U16925 (N_16925,N_16722,N_16793);
xor U16926 (N_16926,N_16697,N_16706);
and U16927 (N_16927,N_16769,N_16695);
and U16928 (N_16928,N_16646,N_16685);
nor U16929 (N_16929,N_16654,N_16683);
nand U16930 (N_16930,N_16711,N_16767);
xor U16931 (N_16931,N_16799,N_16725);
and U16932 (N_16932,N_16783,N_16697);
nand U16933 (N_16933,N_16717,N_16650);
nor U16934 (N_16934,N_16793,N_16725);
xnor U16935 (N_16935,N_16692,N_16679);
xnor U16936 (N_16936,N_16759,N_16710);
or U16937 (N_16937,N_16718,N_16712);
nor U16938 (N_16938,N_16749,N_16725);
xnor U16939 (N_16939,N_16670,N_16655);
and U16940 (N_16940,N_16685,N_16716);
nand U16941 (N_16941,N_16716,N_16739);
xor U16942 (N_16942,N_16725,N_16669);
nand U16943 (N_16943,N_16771,N_16646);
nand U16944 (N_16944,N_16641,N_16792);
and U16945 (N_16945,N_16769,N_16731);
or U16946 (N_16946,N_16731,N_16774);
and U16947 (N_16947,N_16694,N_16761);
nand U16948 (N_16948,N_16795,N_16720);
or U16949 (N_16949,N_16674,N_16765);
and U16950 (N_16950,N_16644,N_16720);
and U16951 (N_16951,N_16728,N_16717);
or U16952 (N_16952,N_16727,N_16648);
or U16953 (N_16953,N_16742,N_16675);
nand U16954 (N_16954,N_16668,N_16755);
and U16955 (N_16955,N_16645,N_16665);
nor U16956 (N_16956,N_16641,N_16771);
nand U16957 (N_16957,N_16737,N_16683);
and U16958 (N_16958,N_16719,N_16643);
and U16959 (N_16959,N_16770,N_16734);
nand U16960 (N_16960,N_16848,N_16833);
nor U16961 (N_16961,N_16917,N_16810);
or U16962 (N_16962,N_16872,N_16950);
or U16963 (N_16963,N_16907,N_16928);
nor U16964 (N_16964,N_16891,N_16904);
nand U16965 (N_16965,N_16820,N_16929);
nor U16966 (N_16966,N_16886,N_16817);
or U16967 (N_16967,N_16939,N_16895);
xnor U16968 (N_16968,N_16836,N_16945);
or U16969 (N_16969,N_16857,N_16899);
or U16970 (N_16970,N_16864,N_16953);
xor U16971 (N_16971,N_16839,N_16855);
or U16972 (N_16972,N_16812,N_16959);
or U16973 (N_16973,N_16805,N_16877);
nor U16974 (N_16974,N_16860,N_16896);
and U16975 (N_16975,N_16863,N_16838);
nand U16976 (N_16976,N_16955,N_16876);
nor U16977 (N_16977,N_16865,N_16853);
nor U16978 (N_16978,N_16831,N_16870);
nor U16979 (N_16979,N_16801,N_16800);
nand U16980 (N_16980,N_16909,N_16921);
and U16981 (N_16981,N_16887,N_16845);
and U16982 (N_16982,N_16878,N_16932);
nor U16983 (N_16983,N_16912,N_16911);
and U16984 (N_16984,N_16813,N_16844);
and U16985 (N_16985,N_16931,N_16825);
xor U16986 (N_16986,N_16826,N_16942);
and U16987 (N_16987,N_16867,N_16832);
xnor U16988 (N_16988,N_16819,N_16823);
or U16989 (N_16989,N_16952,N_16874);
and U16990 (N_16990,N_16869,N_16946);
xor U16991 (N_16991,N_16951,N_16940);
nor U16992 (N_16992,N_16814,N_16935);
xnor U16993 (N_16993,N_16829,N_16954);
xor U16994 (N_16994,N_16892,N_16862);
nor U16995 (N_16995,N_16913,N_16908);
nand U16996 (N_16996,N_16824,N_16828);
nand U16997 (N_16997,N_16861,N_16881);
and U16998 (N_16998,N_16875,N_16956);
or U16999 (N_16999,N_16849,N_16850);
nor U17000 (N_17000,N_16901,N_16941);
nand U17001 (N_17001,N_16818,N_16905);
or U17002 (N_17002,N_16802,N_16902);
nand U17003 (N_17003,N_16834,N_16837);
or U17004 (N_17004,N_16918,N_16898);
nor U17005 (N_17005,N_16847,N_16906);
and U17006 (N_17006,N_16811,N_16927);
xor U17007 (N_17007,N_16804,N_16885);
or U17008 (N_17008,N_16854,N_16947);
xnor U17009 (N_17009,N_16882,N_16893);
and U17010 (N_17010,N_16933,N_16936);
and U17011 (N_17011,N_16949,N_16937);
nor U17012 (N_17012,N_16900,N_16821);
xnor U17013 (N_17013,N_16897,N_16809);
nor U17014 (N_17014,N_16883,N_16923);
nand U17015 (N_17015,N_16889,N_16925);
xor U17016 (N_17016,N_16873,N_16915);
and U17017 (N_17017,N_16944,N_16880);
or U17018 (N_17018,N_16948,N_16914);
xor U17019 (N_17019,N_16816,N_16866);
or U17020 (N_17020,N_16884,N_16830);
nor U17021 (N_17021,N_16856,N_16920);
or U17022 (N_17022,N_16815,N_16924);
nor U17023 (N_17023,N_16894,N_16822);
or U17024 (N_17024,N_16922,N_16846);
nand U17025 (N_17025,N_16868,N_16840);
and U17026 (N_17026,N_16957,N_16926);
nand U17027 (N_17027,N_16859,N_16888);
nor U17028 (N_17028,N_16958,N_16858);
nand U17029 (N_17029,N_16827,N_16938);
nand U17030 (N_17030,N_16852,N_16871);
nand U17031 (N_17031,N_16851,N_16835);
nand U17032 (N_17032,N_16934,N_16803);
xnor U17033 (N_17033,N_16807,N_16903);
nand U17034 (N_17034,N_16806,N_16808);
or U17035 (N_17035,N_16890,N_16910);
or U17036 (N_17036,N_16842,N_16919);
nand U17037 (N_17037,N_16916,N_16841);
nor U17038 (N_17038,N_16930,N_16843);
nand U17039 (N_17039,N_16943,N_16879);
or U17040 (N_17040,N_16820,N_16926);
xnor U17041 (N_17041,N_16934,N_16930);
nor U17042 (N_17042,N_16820,N_16865);
or U17043 (N_17043,N_16847,N_16829);
nor U17044 (N_17044,N_16881,N_16906);
xnor U17045 (N_17045,N_16896,N_16824);
or U17046 (N_17046,N_16886,N_16846);
or U17047 (N_17047,N_16892,N_16878);
xnor U17048 (N_17048,N_16817,N_16901);
or U17049 (N_17049,N_16896,N_16845);
nor U17050 (N_17050,N_16811,N_16886);
and U17051 (N_17051,N_16948,N_16913);
xnor U17052 (N_17052,N_16863,N_16899);
nor U17053 (N_17053,N_16809,N_16889);
xnor U17054 (N_17054,N_16805,N_16903);
nand U17055 (N_17055,N_16874,N_16923);
nand U17056 (N_17056,N_16825,N_16873);
and U17057 (N_17057,N_16959,N_16941);
or U17058 (N_17058,N_16890,N_16912);
and U17059 (N_17059,N_16847,N_16874);
nor U17060 (N_17060,N_16944,N_16938);
nor U17061 (N_17061,N_16821,N_16810);
nand U17062 (N_17062,N_16910,N_16858);
or U17063 (N_17063,N_16936,N_16881);
and U17064 (N_17064,N_16825,N_16882);
nand U17065 (N_17065,N_16928,N_16929);
and U17066 (N_17066,N_16840,N_16941);
or U17067 (N_17067,N_16836,N_16849);
nand U17068 (N_17068,N_16950,N_16816);
and U17069 (N_17069,N_16836,N_16901);
xor U17070 (N_17070,N_16932,N_16889);
and U17071 (N_17071,N_16806,N_16878);
nor U17072 (N_17072,N_16958,N_16808);
and U17073 (N_17073,N_16902,N_16942);
xor U17074 (N_17074,N_16871,N_16881);
nand U17075 (N_17075,N_16893,N_16910);
nand U17076 (N_17076,N_16806,N_16957);
or U17077 (N_17077,N_16907,N_16900);
or U17078 (N_17078,N_16940,N_16810);
nand U17079 (N_17079,N_16886,N_16824);
xnor U17080 (N_17080,N_16922,N_16869);
or U17081 (N_17081,N_16954,N_16944);
nor U17082 (N_17082,N_16850,N_16907);
and U17083 (N_17083,N_16852,N_16843);
and U17084 (N_17084,N_16876,N_16800);
nor U17085 (N_17085,N_16945,N_16801);
or U17086 (N_17086,N_16918,N_16832);
nand U17087 (N_17087,N_16910,N_16809);
and U17088 (N_17088,N_16867,N_16864);
nand U17089 (N_17089,N_16916,N_16891);
or U17090 (N_17090,N_16928,N_16883);
xnor U17091 (N_17091,N_16895,N_16858);
nand U17092 (N_17092,N_16851,N_16863);
xor U17093 (N_17093,N_16897,N_16887);
nor U17094 (N_17094,N_16835,N_16955);
and U17095 (N_17095,N_16943,N_16847);
xnor U17096 (N_17096,N_16897,N_16854);
xor U17097 (N_17097,N_16912,N_16821);
nor U17098 (N_17098,N_16834,N_16857);
and U17099 (N_17099,N_16926,N_16876);
nor U17100 (N_17100,N_16957,N_16903);
nand U17101 (N_17101,N_16827,N_16896);
xor U17102 (N_17102,N_16936,N_16860);
and U17103 (N_17103,N_16850,N_16857);
and U17104 (N_17104,N_16903,N_16808);
nor U17105 (N_17105,N_16820,N_16931);
or U17106 (N_17106,N_16875,N_16850);
nand U17107 (N_17107,N_16934,N_16947);
or U17108 (N_17108,N_16844,N_16944);
xnor U17109 (N_17109,N_16839,N_16947);
and U17110 (N_17110,N_16904,N_16954);
nor U17111 (N_17111,N_16928,N_16840);
nor U17112 (N_17112,N_16813,N_16929);
or U17113 (N_17113,N_16824,N_16858);
or U17114 (N_17114,N_16808,N_16897);
and U17115 (N_17115,N_16956,N_16883);
and U17116 (N_17116,N_16835,N_16859);
nand U17117 (N_17117,N_16826,N_16851);
and U17118 (N_17118,N_16888,N_16912);
xnor U17119 (N_17119,N_16898,N_16809);
xnor U17120 (N_17120,N_17072,N_17027);
nor U17121 (N_17121,N_17079,N_17012);
nor U17122 (N_17122,N_17089,N_17116);
nor U17123 (N_17123,N_17074,N_17001);
or U17124 (N_17124,N_16968,N_17064);
or U17125 (N_17125,N_16970,N_16964);
xor U17126 (N_17126,N_17068,N_16967);
and U17127 (N_17127,N_16989,N_16961);
xnor U17128 (N_17128,N_17007,N_17114);
and U17129 (N_17129,N_17015,N_17037);
or U17130 (N_17130,N_17022,N_17021);
xor U17131 (N_17131,N_17110,N_17078);
and U17132 (N_17132,N_17035,N_17067);
nand U17133 (N_17133,N_17094,N_16986);
or U17134 (N_17134,N_16973,N_17005);
xor U17135 (N_17135,N_17034,N_17091);
and U17136 (N_17136,N_17008,N_17002);
xnor U17137 (N_17137,N_17096,N_16971);
xor U17138 (N_17138,N_17055,N_16969);
nor U17139 (N_17139,N_16977,N_17107);
and U17140 (N_17140,N_17070,N_16976);
and U17141 (N_17141,N_17057,N_17024);
xor U17142 (N_17142,N_17090,N_17026);
nand U17143 (N_17143,N_17060,N_17108);
nor U17144 (N_17144,N_17073,N_17031);
and U17145 (N_17145,N_16972,N_17032);
xnor U17146 (N_17146,N_16981,N_17106);
or U17147 (N_17147,N_17084,N_16974);
nor U17148 (N_17148,N_17036,N_17076);
nor U17149 (N_17149,N_16995,N_17099);
nand U17150 (N_17150,N_17100,N_17109);
nand U17151 (N_17151,N_17040,N_17025);
xor U17152 (N_17152,N_16978,N_17097);
nor U17153 (N_17153,N_16965,N_17081);
nand U17154 (N_17154,N_17049,N_16966);
nand U17155 (N_17155,N_17112,N_16996);
or U17156 (N_17156,N_17085,N_16991);
and U17157 (N_17157,N_17029,N_17065);
nor U17158 (N_17158,N_17047,N_17095);
or U17159 (N_17159,N_17080,N_17086);
or U17160 (N_17160,N_16979,N_16988);
nand U17161 (N_17161,N_17030,N_17098);
xnor U17162 (N_17162,N_16993,N_17056);
nor U17163 (N_17163,N_17044,N_17051);
nor U17164 (N_17164,N_17111,N_17006);
nand U17165 (N_17165,N_17103,N_17019);
nor U17166 (N_17166,N_16987,N_17088);
nor U17167 (N_17167,N_17009,N_17016);
nor U17168 (N_17168,N_17041,N_17017);
or U17169 (N_17169,N_17119,N_17014);
or U17170 (N_17170,N_17087,N_17059);
or U17171 (N_17171,N_17113,N_17050);
xnor U17172 (N_17172,N_17052,N_17071);
nor U17173 (N_17173,N_16992,N_16999);
xnor U17174 (N_17174,N_17010,N_17048);
nand U17175 (N_17175,N_17083,N_17058);
nor U17176 (N_17176,N_17043,N_17011);
xor U17177 (N_17177,N_17038,N_17104);
xnor U17178 (N_17178,N_17003,N_17046);
nand U17179 (N_17179,N_17117,N_16994);
and U17180 (N_17180,N_17118,N_16960);
nor U17181 (N_17181,N_17013,N_17039);
nor U17182 (N_17182,N_17066,N_16997);
or U17183 (N_17183,N_17018,N_17101);
and U17184 (N_17184,N_17033,N_16985);
or U17185 (N_17185,N_17105,N_17063);
and U17186 (N_17186,N_16998,N_17028);
and U17187 (N_17187,N_16982,N_16990);
or U17188 (N_17188,N_16975,N_17042);
xor U17189 (N_17189,N_17077,N_17082);
nor U17190 (N_17190,N_17069,N_16984);
nor U17191 (N_17191,N_17075,N_17102);
or U17192 (N_17192,N_17115,N_17061);
or U17193 (N_17193,N_17053,N_16962);
nor U17194 (N_17194,N_17020,N_17000);
xor U17195 (N_17195,N_17093,N_17004);
or U17196 (N_17196,N_17023,N_17054);
or U17197 (N_17197,N_17092,N_17045);
or U17198 (N_17198,N_16983,N_17062);
nand U17199 (N_17199,N_16980,N_16963);
nor U17200 (N_17200,N_17075,N_16977);
nand U17201 (N_17201,N_17111,N_17064);
xor U17202 (N_17202,N_16993,N_17108);
nor U17203 (N_17203,N_17020,N_17056);
xnor U17204 (N_17204,N_17112,N_17077);
or U17205 (N_17205,N_16973,N_17072);
xnor U17206 (N_17206,N_17022,N_17093);
or U17207 (N_17207,N_17043,N_17090);
nand U17208 (N_17208,N_16982,N_17047);
and U17209 (N_17209,N_17051,N_17087);
nand U17210 (N_17210,N_17115,N_17086);
nand U17211 (N_17211,N_17087,N_16981);
nor U17212 (N_17212,N_17020,N_17097);
xnor U17213 (N_17213,N_17086,N_17038);
and U17214 (N_17214,N_17024,N_16999);
and U17215 (N_17215,N_17048,N_16978);
and U17216 (N_17216,N_17048,N_16974);
nor U17217 (N_17217,N_17028,N_16960);
xnor U17218 (N_17218,N_17072,N_17106);
nor U17219 (N_17219,N_17033,N_17078);
nand U17220 (N_17220,N_17103,N_17080);
or U17221 (N_17221,N_16981,N_17048);
and U17222 (N_17222,N_17045,N_17068);
and U17223 (N_17223,N_16979,N_17045);
xnor U17224 (N_17224,N_17101,N_16978);
or U17225 (N_17225,N_17033,N_17097);
or U17226 (N_17226,N_16963,N_17026);
nand U17227 (N_17227,N_17050,N_17008);
xor U17228 (N_17228,N_17091,N_17036);
or U17229 (N_17229,N_17010,N_16999);
and U17230 (N_17230,N_17062,N_17054);
nor U17231 (N_17231,N_17037,N_17075);
nor U17232 (N_17232,N_17075,N_17099);
nor U17233 (N_17233,N_17100,N_17002);
xnor U17234 (N_17234,N_17003,N_17109);
or U17235 (N_17235,N_17052,N_17001);
or U17236 (N_17236,N_17011,N_17118);
nor U17237 (N_17237,N_17109,N_16981);
and U17238 (N_17238,N_17060,N_17096);
nor U17239 (N_17239,N_16988,N_17104);
nor U17240 (N_17240,N_17017,N_17108);
and U17241 (N_17241,N_17119,N_17047);
nor U17242 (N_17242,N_17044,N_17033);
and U17243 (N_17243,N_17072,N_17060);
and U17244 (N_17244,N_17027,N_17071);
xor U17245 (N_17245,N_17101,N_17044);
and U17246 (N_17246,N_17089,N_17075);
nand U17247 (N_17247,N_17114,N_17009);
nand U17248 (N_17248,N_17078,N_17104);
or U17249 (N_17249,N_17038,N_16968);
xor U17250 (N_17250,N_16997,N_17071);
xor U17251 (N_17251,N_16975,N_17022);
nand U17252 (N_17252,N_16993,N_17088);
or U17253 (N_17253,N_17113,N_17114);
nand U17254 (N_17254,N_16991,N_16980);
nor U17255 (N_17255,N_17109,N_16977);
and U17256 (N_17256,N_17072,N_17031);
or U17257 (N_17257,N_16990,N_17044);
nand U17258 (N_17258,N_17096,N_17012);
or U17259 (N_17259,N_17071,N_17001);
and U17260 (N_17260,N_17018,N_16978);
and U17261 (N_17261,N_16986,N_17058);
or U17262 (N_17262,N_17078,N_16971);
or U17263 (N_17263,N_17005,N_17097);
xnor U17264 (N_17264,N_17028,N_17014);
nand U17265 (N_17265,N_17059,N_17028);
or U17266 (N_17266,N_16975,N_17009);
xnor U17267 (N_17267,N_17043,N_17065);
nor U17268 (N_17268,N_17069,N_17025);
and U17269 (N_17269,N_16980,N_17014);
nand U17270 (N_17270,N_16986,N_17045);
or U17271 (N_17271,N_17052,N_17104);
xnor U17272 (N_17272,N_16984,N_17087);
xor U17273 (N_17273,N_16991,N_16960);
and U17274 (N_17274,N_17102,N_17104);
and U17275 (N_17275,N_16964,N_17060);
or U17276 (N_17276,N_17023,N_17076);
xnor U17277 (N_17277,N_17050,N_17112);
xor U17278 (N_17278,N_17023,N_16964);
or U17279 (N_17279,N_17031,N_16985);
xor U17280 (N_17280,N_17126,N_17219);
xnor U17281 (N_17281,N_17125,N_17171);
nor U17282 (N_17282,N_17254,N_17275);
nor U17283 (N_17283,N_17258,N_17140);
xor U17284 (N_17284,N_17210,N_17183);
xnor U17285 (N_17285,N_17278,N_17273);
or U17286 (N_17286,N_17242,N_17224);
xor U17287 (N_17287,N_17132,N_17235);
nand U17288 (N_17288,N_17147,N_17246);
nand U17289 (N_17289,N_17180,N_17267);
nor U17290 (N_17290,N_17265,N_17141);
xor U17291 (N_17291,N_17160,N_17136);
nand U17292 (N_17292,N_17144,N_17270);
nor U17293 (N_17293,N_17233,N_17269);
and U17294 (N_17294,N_17276,N_17191);
xor U17295 (N_17295,N_17240,N_17179);
or U17296 (N_17296,N_17199,N_17260);
nand U17297 (N_17297,N_17268,N_17205);
nand U17298 (N_17298,N_17266,N_17245);
nor U17299 (N_17299,N_17129,N_17128);
or U17300 (N_17300,N_17271,N_17252);
nand U17301 (N_17301,N_17263,N_17256);
and U17302 (N_17302,N_17241,N_17186);
and U17303 (N_17303,N_17124,N_17145);
nor U17304 (N_17304,N_17151,N_17274);
nand U17305 (N_17305,N_17193,N_17135);
nand U17306 (N_17306,N_17175,N_17243);
or U17307 (N_17307,N_17154,N_17190);
nor U17308 (N_17308,N_17178,N_17163);
and U17309 (N_17309,N_17211,N_17214);
nand U17310 (N_17310,N_17225,N_17203);
nor U17311 (N_17311,N_17182,N_17202);
nand U17312 (N_17312,N_17272,N_17277);
and U17313 (N_17313,N_17184,N_17208);
nor U17314 (N_17314,N_17229,N_17255);
nand U17315 (N_17315,N_17253,N_17162);
xor U17316 (N_17316,N_17220,N_17195);
xor U17317 (N_17317,N_17207,N_17216);
and U17318 (N_17318,N_17122,N_17123);
nor U17319 (N_17319,N_17153,N_17169);
nor U17320 (N_17320,N_17127,N_17181);
xnor U17321 (N_17321,N_17121,N_17247);
nor U17322 (N_17322,N_17173,N_17213);
or U17323 (N_17323,N_17222,N_17130);
or U17324 (N_17324,N_17192,N_17152);
xor U17325 (N_17325,N_17198,N_17155);
nor U17326 (N_17326,N_17146,N_17176);
nand U17327 (N_17327,N_17204,N_17164);
nor U17328 (N_17328,N_17218,N_17139);
nor U17329 (N_17329,N_17237,N_17223);
or U17330 (N_17330,N_17212,N_17170);
nand U17331 (N_17331,N_17194,N_17157);
or U17332 (N_17332,N_17239,N_17134);
nand U17333 (N_17333,N_17264,N_17131);
xor U17334 (N_17334,N_17230,N_17200);
xnor U17335 (N_17335,N_17206,N_17172);
xnor U17336 (N_17336,N_17166,N_17226);
nor U17337 (N_17337,N_17148,N_17150);
and U17338 (N_17338,N_17215,N_17231);
or U17339 (N_17339,N_17238,N_17232);
nor U17340 (N_17340,N_17174,N_17188);
or U17341 (N_17341,N_17189,N_17142);
nor U17342 (N_17342,N_17137,N_17244);
or U17343 (N_17343,N_17167,N_17250);
nand U17344 (N_17344,N_17177,N_17161);
xnor U17345 (N_17345,N_17168,N_17251);
or U17346 (N_17346,N_17133,N_17221);
or U17347 (N_17347,N_17201,N_17248);
xor U17348 (N_17348,N_17159,N_17156);
or U17349 (N_17349,N_17228,N_17261);
nor U17350 (N_17350,N_17165,N_17143);
or U17351 (N_17351,N_17279,N_17257);
nand U17352 (N_17352,N_17158,N_17249);
nand U17353 (N_17353,N_17234,N_17262);
and U17354 (N_17354,N_17196,N_17197);
and U17355 (N_17355,N_17120,N_17227);
nor U17356 (N_17356,N_17149,N_17236);
and U17357 (N_17357,N_17217,N_17185);
nand U17358 (N_17358,N_17187,N_17259);
nand U17359 (N_17359,N_17138,N_17209);
nor U17360 (N_17360,N_17230,N_17251);
or U17361 (N_17361,N_17135,N_17140);
or U17362 (N_17362,N_17141,N_17259);
nand U17363 (N_17363,N_17278,N_17217);
xnor U17364 (N_17364,N_17167,N_17222);
xor U17365 (N_17365,N_17279,N_17216);
nand U17366 (N_17366,N_17222,N_17143);
nand U17367 (N_17367,N_17224,N_17226);
and U17368 (N_17368,N_17220,N_17178);
and U17369 (N_17369,N_17170,N_17240);
or U17370 (N_17370,N_17254,N_17161);
nand U17371 (N_17371,N_17130,N_17252);
nand U17372 (N_17372,N_17259,N_17237);
and U17373 (N_17373,N_17206,N_17223);
and U17374 (N_17374,N_17248,N_17268);
nor U17375 (N_17375,N_17145,N_17143);
nand U17376 (N_17376,N_17169,N_17266);
or U17377 (N_17377,N_17232,N_17144);
xnor U17378 (N_17378,N_17203,N_17163);
and U17379 (N_17379,N_17276,N_17206);
and U17380 (N_17380,N_17162,N_17271);
nand U17381 (N_17381,N_17250,N_17177);
xor U17382 (N_17382,N_17197,N_17171);
nand U17383 (N_17383,N_17277,N_17154);
and U17384 (N_17384,N_17272,N_17262);
nor U17385 (N_17385,N_17171,N_17266);
nor U17386 (N_17386,N_17131,N_17268);
xnor U17387 (N_17387,N_17268,N_17167);
and U17388 (N_17388,N_17240,N_17148);
and U17389 (N_17389,N_17246,N_17122);
and U17390 (N_17390,N_17217,N_17258);
nor U17391 (N_17391,N_17247,N_17243);
nand U17392 (N_17392,N_17272,N_17271);
nand U17393 (N_17393,N_17279,N_17274);
or U17394 (N_17394,N_17187,N_17266);
xor U17395 (N_17395,N_17260,N_17180);
nand U17396 (N_17396,N_17162,N_17148);
or U17397 (N_17397,N_17237,N_17129);
nor U17398 (N_17398,N_17266,N_17254);
nor U17399 (N_17399,N_17131,N_17123);
and U17400 (N_17400,N_17176,N_17182);
xor U17401 (N_17401,N_17209,N_17252);
nand U17402 (N_17402,N_17145,N_17236);
or U17403 (N_17403,N_17221,N_17269);
nor U17404 (N_17404,N_17268,N_17238);
xor U17405 (N_17405,N_17126,N_17135);
and U17406 (N_17406,N_17219,N_17171);
nand U17407 (N_17407,N_17147,N_17160);
or U17408 (N_17408,N_17220,N_17256);
nor U17409 (N_17409,N_17151,N_17158);
and U17410 (N_17410,N_17225,N_17160);
or U17411 (N_17411,N_17235,N_17248);
nand U17412 (N_17412,N_17156,N_17232);
and U17413 (N_17413,N_17223,N_17236);
xnor U17414 (N_17414,N_17131,N_17273);
xor U17415 (N_17415,N_17140,N_17275);
nand U17416 (N_17416,N_17182,N_17169);
xor U17417 (N_17417,N_17271,N_17277);
or U17418 (N_17418,N_17204,N_17158);
xor U17419 (N_17419,N_17279,N_17219);
nand U17420 (N_17420,N_17241,N_17198);
xor U17421 (N_17421,N_17162,N_17199);
xor U17422 (N_17422,N_17248,N_17266);
xnor U17423 (N_17423,N_17134,N_17219);
nand U17424 (N_17424,N_17218,N_17175);
or U17425 (N_17425,N_17228,N_17164);
or U17426 (N_17426,N_17236,N_17141);
nor U17427 (N_17427,N_17162,N_17158);
xor U17428 (N_17428,N_17135,N_17221);
and U17429 (N_17429,N_17245,N_17163);
nand U17430 (N_17430,N_17167,N_17183);
nor U17431 (N_17431,N_17234,N_17176);
nor U17432 (N_17432,N_17228,N_17262);
nor U17433 (N_17433,N_17197,N_17234);
or U17434 (N_17434,N_17164,N_17201);
and U17435 (N_17435,N_17145,N_17199);
nand U17436 (N_17436,N_17223,N_17152);
and U17437 (N_17437,N_17205,N_17158);
nand U17438 (N_17438,N_17247,N_17195);
or U17439 (N_17439,N_17269,N_17139);
or U17440 (N_17440,N_17335,N_17379);
nand U17441 (N_17441,N_17344,N_17373);
and U17442 (N_17442,N_17322,N_17426);
or U17443 (N_17443,N_17329,N_17417);
or U17444 (N_17444,N_17309,N_17287);
nor U17445 (N_17445,N_17400,N_17331);
nor U17446 (N_17446,N_17420,N_17352);
nand U17447 (N_17447,N_17356,N_17409);
nand U17448 (N_17448,N_17377,N_17419);
xnor U17449 (N_17449,N_17389,N_17403);
nand U17450 (N_17450,N_17438,N_17401);
or U17451 (N_17451,N_17307,N_17361);
or U17452 (N_17452,N_17293,N_17312);
or U17453 (N_17453,N_17319,N_17434);
or U17454 (N_17454,N_17375,N_17385);
nand U17455 (N_17455,N_17341,N_17428);
nand U17456 (N_17456,N_17324,N_17314);
and U17457 (N_17457,N_17320,N_17342);
or U17458 (N_17458,N_17340,N_17354);
nor U17459 (N_17459,N_17378,N_17355);
nand U17460 (N_17460,N_17422,N_17423);
nor U17461 (N_17461,N_17338,N_17416);
xnor U17462 (N_17462,N_17339,N_17301);
nand U17463 (N_17463,N_17291,N_17316);
xnor U17464 (N_17464,N_17295,N_17418);
xor U17465 (N_17465,N_17386,N_17299);
xor U17466 (N_17466,N_17365,N_17376);
nand U17467 (N_17467,N_17302,N_17292);
nand U17468 (N_17468,N_17437,N_17286);
nand U17469 (N_17469,N_17429,N_17387);
nor U17470 (N_17470,N_17280,N_17405);
and U17471 (N_17471,N_17369,N_17305);
nor U17472 (N_17472,N_17284,N_17433);
nor U17473 (N_17473,N_17435,N_17349);
or U17474 (N_17474,N_17323,N_17282);
or U17475 (N_17475,N_17391,N_17406);
or U17476 (N_17476,N_17285,N_17348);
and U17477 (N_17477,N_17351,N_17415);
xor U17478 (N_17478,N_17388,N_17362);
xor U17479 (N_17479,N_17411,N_17436);
nor U17480 (N_17480,N_17407,N_17371);
nand U17481 (N_17481,N_17396,N_17374);
nand U17482 (N_17482,N_17336,N_17350);
and U17483 (N_17483,N_17390,N_17421);
xor U17484 (N_17484,N_17398,N_17358);
nor U17485 (N_17485,N_17408,N_17306);
or U17486 (N_17486,N_17347,N_17283);
nand U17487 (N_17487,N_17367,N_17333);
nand U17488 (N_17488,N_17363,N_17399);
nor U17489 (N_17489,N_17326,N_17313);
nor U17490 (N_17490,N_17357,N_17412);
xor U17491 (N_17491,N_17334,N_17300);
or U17492 (N_17492,N_17414,N_17393);
nand U17493 (N_17493,N_17360,N_17315);
nor U17494 (N_17494,N_17431,N_17345);
or U17495 (N_17495,N_17427,N_17297);
or U17496 (N_17496,N_17330,N_17397);
and U17497 (N_17497,N_17424,N_17332);
nand U17498 (N_17498,N_17288,N_17368);
nor U17499 (N_17499,N_17380,N_17311);
or U17500 (N_17500,N_17290,N_17325);
nor U17501 (N_17501,N_17298,N_17308);
or U17502 (N_17502,N_17372,N_17402);
nor U17503 (N_17503,N_17364,N_17439);
nor U17504 (N_17504,N_17294,N_17337);
nand U17505 (N_17505,N_17425,N_17381);
xnor U17506 (N_17506,N_17366,N_17296);
nand U17507 (N_17507,N_17328,N_17395);
or U17508 (N_17508,N_17384,N_17317);
or U17509 (N_17509,N_17343,N_17327);
or U17510 (N_17510,N_17382,N_17353);
or U17511 (N_17511,N_17370,N_17359);
and U17512 (N_17512,N_17281,N_17321);
and U17513 (N_17513,N_17310,N_17392);
or U17514 (N_17514,N_17413,N_17289);
or U17515 (N_17515,N_17346,N_17432);
nand U17516 (N_17516,N_17303,N_17404);
and U17517 (N_17517,N_17304,N_17318);
nand U17518 (N_17518,N_17410,N_17430);
xor U17519 (N_17519,N_17394,N_17383);
and U17520 (N_17520,N_17325,N_17365);
xor U17521 (N_17521,N_17411,N_17348);
nor U17522 (N_17522,N_17397,N_17352);
or U17523 (N_17523,N_17431,N_17410);
nand U17524 (N_17524,N_17297,N_17342);
nor U17525 (N_17525,N_17284,N_17312);
xnor U17526 (N_17526,N_17361,N_17285);
xor U17527 (N_17527,N_17325,N_17301);
nand U17528 (N_17528,N_17332,N_17426);
and U17529 (N_17529,N_17411,N_17393);
nand U17530 (N_17530,N_17285,N_17299);
xnor U17531 (N_17531,N_17289,N_17369);
or U17532 (N_17532,N_17294,N_17343);
and U17533 (N_17533,N_17367,N_17294);
nor U17534 (N_17534,N_17343,N_17394);
and U17535 (N_17535,N_17334,N_17411);
xor U17536 (N_17536,N_17377,N_17299);
or U17537 (N_17537,N_17332,N_17312);
or U17538 (N_17538,N_17389,N_17335);
xor U17539 (N_17539,N_17346,N_17294);
nor U17540 (N_17540,N_17375,N_17423);
or U17541 (N_17541,N_17348,N_17362);
or U17542 (N_17542,N_17396,N_17351);
or U17543 (N_17543,N_17345,N_17400);
or U17544 (N_17544,N_17378,N_17385);
xnor U17545 (N_17545,N_17320,N_17417);
or U17546 (N_17546,N_17430,N_17335);
or U17547 (N_17547,N_17300,N_17301);
nor U17548 (N_17548,N_17372,N_17415);
nor U17549 (N_17549,N_17283,N_17369);
nand U17550 (N_17550,N_17436,N_17375);
and U17551 (N_17551,N_17342,N_17411);
nand U17552 (N_17552,N_17402,N_17327);
xnor U17553 (N_17553,N_17336,N_17367);
nor U17554 (N_17554,N_17347,N_17338);
nand U17555 (N_17555,N_17313,N_17314);
nor U17556 (N_17556,N_17390,N_17430);
nand U17557 (N_17557,N_17312,N_17381);
and U17558 (N_17558,N_17325,N_17435);
nor U17559 (N_17559,N_17437,N_17434);
nand U17560 (N_17560,N_17385,N_17349);
and U17561 (N_17561,N_17362,N_17389);
nor U17562 (N_17562,N_17381,N_17356);
and U17563 (N_17563,N_17325,N_17398);
nand U17564 (N_17564,N_17371,N_17306);
and U17565 (N_17565,N_17421,N_17333);
or U17566 (N_17566,N_17295,N_17286);
and U17567 (N_17567,N_17301,N_17401);
xor U17568 (N_17568,N_17324,N_17288);
and U17569 (N_17569,N_17407,N_17308);
and U17570 (N_17570,N_17310,N_17315);
and U17571 (N_17571,N_17381,N_17360);
and U17572 (N_17572,N_17432,N_17345);
xor U17573 (N_17573,N_17435,N_17429);
and U17574 (N_17574,N_17306,N_17351);
or U17575 (N_17575,N_17293,N_17325);
nor U17576 (N_17576,N_17371,N_17365);
and U17577 (N_17577,N_17382,N_17426);
xor U17578 (N_17578,N_17301,N_17398);
nor U17579 (N_17579,N_17305,N_17311);
or U17580 (N_17580,N_17384,N_17386);
nand U17581 (N_17581,N_17355,N_17413);
nand U17582 (N_17582,N_17336,N_17289);
or U17583 (N_17583,N_17295,N_17289);
xnor U17584 (N_17584,N_17390,N_17338);
xor U17585 (N_17585,N_17395,N_17379);
nor U17586 (N_17586,N_17381,N_17282);
nand U17587 (N_17587,N_17383,N_17360);
nor U17588 (N_17588,N_17416,N_17359);
and U17589 (N_17589,N_17297,N_17402);
nand U17590 (N_17590,N_17304,N_17374);
xnor U17591 (N_17591,N_17287,N_17420);
or U17592 (N_17592,N_17327,N_17393);
nand U17593 (N_17593,N_17301,N_17352);
xnor U17594 (N_17594,N_17337,N_17424);
nand U17595 (N_17595,N_17429,N_17285);
nor U17596 (N_17596,N_17296,N_17286);
or U17597 (N_17597,N_17427,N_17403);
nor U17598 (N_17598,N_17410,N_17369);
or U17599 (N_17599,N_17356,N_17352);
nor U17600 (N_17600,N_17513,N_17448);
nor U17601 (N_17601,N_17515,N_17509);
nor U17602 (N_17602,N_17450,N_17455);
nand U17603 (N_17603,N_17477,N_17542);
and U17604 (N_17604,N_17577,N_17528);
or U17605 (N_17605,N_17486,N_17560);
nor U17606 (N_17606,N_17554,N_17573);
or U17607 (N_17607,N_17501,N_17525);
xnor U17608 (N_17608,N_17583,N_17453);
and U17609 (N_17609,N_17510,N_17543);
or U17610 (N_17610,N_17567,N_17483);
or U17611 (N_17611,N_17473,N_17508);
xor U17612 (N_17612,N_17478,N_17481);
nor U17613 (N_17613,N_17586,N_17548);
nand U17614 (N_17614,N_17452,N_17559);
xnor U17615 (N_17615,N_17574,N_17444);
or U17616 (N_17616,N_17512,N_17460);
nand U17617 (N_17617,N_17449,N_17585);
and U17618 (N_17618,N_17589,N_17480);
xor U17619 (N_17619,N_17563,N_17556);
xnor U17620 (N_17620,N_17507,N_17446);
xnor U17621 (N_17621,N_17492,N_17484);
and U17622 (N_17622,N_17474,N_17550);
nor U17623 (N_17623,N_17491,N_17467);
nand U17624 (N_17624,N_17519,N_17594);
or U17625 (N_17625,N_17552,N_17549);
nor U17626 (N_17626,N_17593,N_17523);
nor U17627 (N_17627,N_17584,N_17546);
or U17628 (N_17628,N_17575,N_17476);
and U17629 (N_17629,N_17497,N_17539);
xor U17630 (N_17630,N_17493,N_17470);
xnor U17631 (N_17631,N_17553,N_17535);
or U17632 (N_17632,N_17443,N_17469);
nor U17633 (N_17633,N_17440,N_17498);
nor U17634 (N_17634,N_17524,N_17475);
xnor U17635 (N_17635,N_17578,N_17555);
xnor U17636 (N_17636,N_17487,N_17527);
and U17637 (N_17637,N_17479,N_17530);
and U17638 (N_17638,N_17540,N_17457);
and U17639 (N_17639,N_17572,N_17551);
and U17640 (N_17640,N_17571,N_17482);
nand U17641 (N_17641,N_17505,N_17579);
and U17642 (N_17642,N_17517,N_17516);
nand U17643 (N_17643,N_17468,N_17458);
nor U17644 (N_17644,N_17558,N_17597);
xnor U17645 (N_17645,N_17562,N_17537);
nor U17646 (N_17646,N_17595,N_17488);
and U17647 (N_17647,N_17456,N_17545);
xor U17648 (N_17648,N_17518,N_17544);
and U17649 (N_17649,N_17533,N_17565);
nand U17650 (N_17650,N_17520,N_17511);
or U17651 (N_17651,N_17561,N_17592);
nand U17652 (N_17652,N_17485,N_17590);
nor U17653 (N_17653,N_17463,N_17504);
and U17654 (N_17654,N_17581,N_17588);
xor U17655 (N_17655,N_17557,N_17547);
nor U17656 (N_17656,N_17536,N_17514);
or U17657 (N_17657,N_17489,N_17462);
nor U17658 (N_17658,N_17521,N_17459);
nand U17659 (N_17659,N_17576,N_17534);
or U17660 (N_17660,N_17569,N_17465);
xnor U17661 (N_17661,N_17499,N_17580);
or U17662 (N_17662,N_17442,N_17464);
nor U17663 (N_17663,N_17466,N_17503);
nand U17664 (N_17664,N_17441,N_17591);
and U17665 (N_17665,N_17447,N_17532);
nor U17666 (N_17666,N_17451,N_17502);
and U17667 (N_17667,N_17490,N_17599);
and U17668 (N_17668,N_17471,N_17500);
xnor U17669 (N_17669,N_17472,N_17461);
nand U17670 (N_17670,N_17566,N_17531);
nand U17671 (N_17671,N_17587,N_17596);
nand U17672 (N_17672,N_17506,N_17529);
and U17673 (N_17673,N_17538,N_17526);
nor U17674 (N_17674,N_17541,N_17598);
nand U17675 (N_17675,N_17494,N_17522);
or U17676 (N_17676,N_17454,N_17564);
nand U17677 (N_17677,N_17570,N_17582);
and U17678 (N_17678,N_17495,N_17496);
nand U17679 (N_17679,N_17568,N_17445);
nand U17680 (N_17680,N_17576,N_17480);
xor U17681 (N_17681,N_17574,N_17474);
or U17682 (N_17682,N_17532,N_17471);
and U17683 (N_17683,N_17572,N_17447);
nor U17684 (N_17684,N_17464,N_17517);
nand U17685 (N_17685,N_17533,N_17447);
nand U17686 (N_17686,N_17496,N_17493);
nor U17687 (N_17687,N_17453,N_17482);
or U17688 (N_17688,N_17566,N_17526);
xnor U17689 (N_17689,N_17524,N_17476);
nand U17690 (N_17690,N_17578,N_17595);
and U17691 (N_17691,N_17520,N_17549);
xnor U17692 (N_17692,N_17580,N_17551);
xor U17693 (N_17693,N_17553,N_17582);
or U17694 (N_17694,N_17477,N_17589);
and U17695 (N_17695,N_17462,N_17544);
nand U17696 (N_17696,N_17553,N_17589);
or U17697 (N_17697,N_17452,N_17535);
nor U17698 (N_17698,N_17591,N_17487);
nor U17699 (N_17699,N_17537,N_17546);
nor U17700 (N_17700,N_17573,N_17598);
xnor U17701 (N_17701,N_17535,N_17532);
xor U17702 (N_17702,N_17595,N_17472);
nand U17703 (N_17703,N_17587,N_17449);
xnor U17704 (N_17704,N_17510,N_17575);
xor U17705 (N_17705,N_17562,N_17517);
xnor U17706 (N_17706,N_17502,N_17587);
and U17707 (N_17707,N_17465,N_17477);
nor U17708 (N_17708,N_17523,N_17469);
and U17709 (N_17709,N_17466,N_17508);
or U17710 (N_17710,N_17455,N_17558);
nor U17711 (N_17711,N_17525,N_17519);
nand U17712 (N_17712,N_17509,N_17573);
nor U17713 (N_17713,N_17452,N_17440);
or U17714 (N_17714,N_17469,N_17531);
or U17715 (N_17715,N_17597,N_17512);
and U17716 (N_17716,N_17474,N_17547);
and U17717 (N_17717,N_17470,N_17525);
nand U17718 (N_17718,N_17566,N_17586);
nand U17719 (N_17719,N_17468,N_17500);
and U17720 (N_17720,N_17492,N_17440);
xor U17721 (N_17721,N_17509,N_17517);
xor U17722 (N_17722,N_17559,N_17468);
or U17723 (N_17723,N_17525,N_17520);
nor U17724 (N_17724,N_17520,N_17462);
nor U17725 (N_17725,N_17528,N_17525);
nor U17726 (N_17726,N_17573,N_17447);
nand U17727 (N_17727,N_17568,N_17547);
or U17728 (N_17728,N_17478,N_17572);
or U17729 (N_17729,N_17571,N_17475);
xnor U17730 (N_17730,N_17503,N_17460);
or U17731 (N_17731,N_17440,N_17524);
and U17732 (N_17732,N_17499,N_17503);
xor U17733 (N_17733,N_17550,N_17493);
nor U17734 (N_17734,N_17521,N_17553);
nand U17735 (N_17735,N_17548,N_17462);
and U17736 (N_17736,N_17455,N_17484);
and U17737 (N_17737,N_17472,N_17566);
or U17738 (N_17738,N_17557,N_17579);
xor U17739 (N_17739,N_17552,N_17528);
nand U17740 (N_17740,N_17460,N_17491);
xor U17741 (N_17741,N_17550,N_17585);
nor U17742 (N_17742,N_17549,N_17464);
nor U17743 (N_17743,N_17505,N_17532);
xor U17744 (N_17744,N_17531,N_17586);
or U17745 (N_17745,N_17526,N_17536);
nor U17746 (N_17746,N_17586,N_17519);
or U17747 (N_17747,N_17458,N_17443);
and U17748 (N_17748,N_17465,N_17515);
nor U17749 (N_17749,N_17532,N_17572);
nand U17750 (N_17750,N_17517,N_17474);
nor U17751 (N_17751,N_17479,N_17442);
nand U17752 (N_17752,N_17467,N_17475);
or U17753 (N_17753,N_17512,N_17509);
or U17754 (N_17754,N_17516,N_17477);
xor U17755 (N_17755,N_17541,N_17448);
nor U17756 (N_17756,N_17524,N_17494);
or U17757 (N_17757,N_17592,N_17588);
or U17758 (N_17758,N_17485,N_17581);
or U17759 (N_17759,N_17572,N_17520);
nor U17760 (N_17760,N_17603,N_17701);
and U17761 (N_17761,N_17704,N_17672);
or U17762 (N_17762,N_17645,N_17629);
xnor U17763 (N_17763,N_17635,N_17706);
or U17764 (N_17764,N_17643,N_17605);
xnor U17765 (N_17765,N_17708,N_17740);
and U17766 (N_17766,N_17681,N_17757);
xnor U17767 (N_17767,N_17602,N_17680);
or U17768 (N_17768,N_17642,N_17688);
or U17769 (N_17769,N_17736,N_17695);
or U17770 (N_17770,N_17662,N_17734);
and U17771 (N_17771,N_17639,N_17620);
and U17772 (N_17772,N_17673,N_17697);
nor U17773 (N_17773,N_17666,N_17606);
xnor U17774 (N_17774,N_17721,N_17678);
or U17775 (N_17775,N_17610,N_17711);
or U17776 (N_17776,N_17632,N_17644);
or U17777 (N_17777,N_17607,N_17756);
or U17778 (N_17778,N_17705,N_17739);
xnor U17779 (N_17779,N_17687,N_17731);
or U17780 (N_17780,N_17655,N_17665);
and U17781 (N_17781,N_17646,N_17745);
nand U17782 (N_17782,N_17661,N_17626);
xnor U17783 (N_17783,N_17675,N_17647);
and U17784 (N_17784,N_17611,N_17613);
xor U17785 (N_17785,N_17730,N_17679);
nor U17786 (N_17786,N_17690,N_17722);
or U17787 (N_17787,N_17657,N_17614);
xor U17788 (N_17788,N_17609,N_17732);
nand U17789 (N_17789,N_17653,N_17692);
nand U17790 (N_17790,N_17670,N_17616);
and U17791 (N_17791,N_17649,N_17625);
or U17792 (N_17792,N_17622,N_17751);
or U17793 (N_17793,N_17748,N_17733);
or U17794 (N_17794,N_17601,N_17750);
nor U17795 (N_17795,N_17630,N_17627);
nand U17796 (N_17796,N_17685,N_17719);
and U17797 (N_17797,N_17671,N_17749);
xnor U17798 (N_17798,N_17698,N_17709);
xor U17799 (N_17799,N_17741,N_17752);
nor U17800 (N_17800,N_17638,N_17634);
xor U17801 (N_17801,N_17628,N_17637);
or U17802 (N_17802,N_17659,N_17648);
and U17803 (N_17803,N_17619,N_17720);
and U17804 (N_17804,N_17693,N_17694);
xor U17805 (N_17805,N_17755,N_17641);
xor U17806 (N_17806,N_17728,N_17656);
or U17807 (N_17807,N_17684,N_17623);
xor U17808 (N_17808,N_17669,N_17617);
or U17809 (N_17809,N_17676,N_17683);
nor U17810 (N_17810,N_17725,N_17727);
and U17811 (N_17811,N_17743,N_17726);
nor U17812 (N_17812,N_17652,N_17636);
nand U17813 (N_17813,N_17717,N_17654);
nor U17814 (N_17814,N_17640,N_17718);
xnor U17815 (N_17815,N_17702,N_17707);
and U17816 (N_17816,N_17714,N_17660);
nand U17817 (N_17817,N_17759,N_17664);
nand U17818 (N_17818,N_17713,N_17691);
nor U17819 (N_17819,N_17689,N_17674);
nand U17820 (N_17820,N_17663,N_17618);
nor U17821 (N_17821,N_17737,N_17696);
and U17822 (N_17822,N_17650,N_17712);
xnor U17823 (N_17823,N_17716,N_17612);
xor U17824 (N_17824,N_17723,N_17735);
nor U17825 (N_17825,N_17651,N_17621);
nor U17826 (N_17826,N_17600,N_17738);
or U17827 (N_17827,N_17744,N_17758);
and U17828 (N_17828,N_17677,N_17710);
xnor U17829 (N_17829,N_17703,N_17700);
xnor U17830 (N_17830,N_17699,N_17729);
nor U17831 (N_17831,N_17608,N_17746);
or U17832 (N_17832,N_17715,N_17624);
nor U17833 (N_17833,N_17667,N_17682);
and U17834 (N_17834,N_17633,N_17753);
and U17835 (N_17835,N_17686,N_17658);
or U17836 (N_17836,N_17754,N_17604);
nand U17837 (N_17837,N_17631,N_17742);
and U17838 (N_17838,N_17724,N_17615);
and U17839 (N_17839,N_17747,N_17668);
or U17840 (N_17840,N_17698,N_17612);
nor U17841 (N_17841,N_17683,N_17745);
and U17842 (N_17842,N_17670,N_17624);
or U17843 (N_17843,N_17633,N_17687);
nor U17844 (N_17844,N_17670,N_17726);
or U17845 (N_17845,N_17690,N_17739);
xor U17846 (N_17846,N_17727,N_17622);
nand U17847 (N_17847,N_17651,N_17600);
or U17848 (N_17848,N_17636,N_17613);
xor U17849 (N_17849,N_17704,N_17603);
xnor U17850 (N_17850,N_17663,N_17695);
or U17851 (N_17851,N_17616,N_17602);
xnor U17852 (N_17852,N_17609,N_17602);
xnor U17853 (N_17853,N_17722,N_17710);
xor U17854 (N_17854,N_17636,N_17682);
and U17855 (N_17855,N_17657,N_17610);
nor U17856 (N_17856,N_17741,N_17600);
or U17857 (N_17857,N_17680,N_17676);
and U17858 (N_17858,N_17656,N_17711);
nand U17859 (N_17859,N_17719,N_17758);
xor U17860 (N_17860,N_17672,N_17707);
nor U17861 (N_17861,N_17661,N_17609);
and U17862 (N_17862,N_17696,N_17741);
xnor U17863 (N_17863,N_17733,N_17604);
nand U17864 (N_17864,N_17611,N_17740);
or U17865 (N_17865,N_17703,N_17670);
nand U17866 (N_17866,N_17683,N_17754);
or U17867 (N_17867,N_17703,N_17678);
nor U17868 (N_17868,N_17693,N_17616);
or U17869 (N_17869,N_17739,N_17746);
nand U17870 (N_17870,N_17681,N_17622);
and U17871 (N_17871,N_17646,N_17720);
xor U17872 (N_17872,N_17733,N_17718);
nor U17873 (N_17873,N_17663,N_17738);
nor U17874 (N_17874,N_17707,N_17666);
xnor U17875 (N_17875,N_17620,N_17740);
and U17876 (N_17876,N_17677,N_17756);
nand U17877 (N_17877,N_17731,N_17712);
or U17878 (N_17878,N_17612,N_17639);
xor U17879 (N_17879,N_17650,N_17747);
nor U17880 (N_17880,N_17703,N_17660);
xnor U17881 (N_17881,N_17618,N_17691);
and U17882 (N_17882,N_17690,N_17613);
and U17883 (N_17883,N_17661,N_17714);
nand U17884 (N_17884,N_17603,N_17684);
nor U17885 (N_17885,N_17612,N_17610);
nor U17886 (N_17886,N_17724,N_17697);
xor U17887 (N_17887,N_17697,N_17740);
and U17888 (N_17888,N_17612,N_17669);
or U17889 (N_17889,N_17654,N_17616);
or U17890 (N_17890,N_17645,N_17755);
and U17891 (N_17891,N_17670,N_17613);
xor U17892 (N_17892,N_17636,N_17720);
xor U17893 (N_17893,N_17743,N_17679);
nor U17894 (N_17894,N_17618,N_17748);
and U17895 (N_17895,N_17650,N_17680);
and U17896 (N_17896,N_17690,N_17734);
nor U17897 (N_17897,N_17653,N_17673);
xor U17898 (N_17898,N_17612,N_17755);
or U17899 (N_17899,N_17674,N_17613);
nor U17900 (N_17900,N_17647,N_17648);
or U17901 (N_17901,N_17696,N_17668);
or U17902 (N_17902,N_17651,N_17664);
nor U17903 (N_17903,N_17677,N_17651);
xnor U17904 (N_17904,N_17675,N_17680);
xor U17905 (N_17905,N_17656,N_17607);
nand U17906 (N_17906,N_17607,N_17697);
nand U17907 (N_17907,N_17667,N_17663);
xor U17908 (N_17908,N_17633,N_17609);
nor U17909 (N_17909,N_17755,N_17678);
nor U17910 (N_17910,N_17651,N_17626);
nand U17911 (N_17911,N_17660,N_17642);
nand U17912 (N_17912,N_17744,N_17719);
nor U17913 (N_17913,N_17633,N_17689);
and U17914 (N_17914,N_17606,N_17653);
and U17915 (N_17915,N_17683,N_17714);
nand U17916 (N_17916,N_17640,N_17614);
nor U17917 (N_17917,N_17614,N_17701);
nor U17918 (N_17918,N_17685,N_17716);
nor U17919 (N_17919,N_17677,N_17755);
nor U17920 (N_17920,N_17906,N_17769);
and U17921 (N_17921,N_17791,N_17828);
nand U17922 (N_17922,N_17794,N_17842);
xor U17923 (N_17923,N_17869,N_17871);
nor U17924 (N_17924,N_17810,N_17849);
nor U17925 (N_17925,N_17891,N_17876);
and U17926 (N_17926,N_17861,N_17881);
or U17927 (N_17927,N_17879,N_17904);
and U17928 (N_17928,N_17914,N_17838);
nand U17929 (N_17929,N_17860,N_17847);
xnor U17930 (N_17930,N_17907,N_17837);
nor U17931 (N_17931,N_17826,N_17793);
and U17932 (N_17932,N_17902,N_17859);
xnor U17933 (N_17933,N_17777,N_17762);
xor U17934 (N_17934,N_17882,N_17767);
nand U17935 (N_17935,N_17760,N_17761);
or U17936 (N_17936,N_17835,N_17796);
or U17937 (N_17937,N_17913,N_17877);
and U17938 (N_17938,N_17889,N_17789);
nor U17939 (N_17939,N_17900,N_17809);
nor U17940 (N_17940,N_17856,N_17901);
and U17941 (N_17941,N_17905,N_17819);
or U17942 (N_17942,N_17917,N_17805);
and U17943 (N_17943,N_17795,N_17840);
nand U17944 (N_17944,N_17829,N_17801);
or U17945 (N_17945,N_17909,N_17897);
xnor U17946 (N_17946,N_17804,N_17787);
nor U17947 (N_17947,N_17855,N_17865);
or U17948 (N_17948,N_17784,N_17806);
and U17949 (N_17949,N_17853,N_17823);
and U17950 (N_17950,N_17885,N_17818);
nand U17951 (N_17951,N_17798,N_17803);
and U17952 (N_17952,N_17911,N_17765);
nand U17953 (N_17953,N_17774,N_17832);
nor U17954 (N_17954,N_17822,N_17852);
nand U17955 (N_17955,N_17813,N_17790);
and U17956 (N_17956,N_17772,N_17824);
nand U17957 (N_17957,N_17894,N_17811);
xnor U17958 (N_17958,N_17783,N_17830);
and U17959 (N_17959,N_17820,N_17816);
nand U17960 (N_17960,N_17844,N_17854);
and U17961 (N_17961,N_17896,N_17785);
nand U17962 (N_17962,N_17776,N_17802);
nor U17963 (N_17963,N_17850,N_17878);
nand U17964 (N_17964,N_17780,N_17903);
and U17965 (N_17965,N_17890,N_17880);
nand U17966 (N_17966,N_17786,N_17833);
and U17967 (N_17967,N_17825,N_17918);
or U17968 (N_17968,N_17886,N_17867);
and U17969 (N_17969,N_17763,N_17843);
xnor U17970 (N_17970,N_17764,N_17872);
nand U17971 (N_17971,N_17870,N_17775);
and U17972 (N_17972,N_17895,N_17766);
nor U17973 (N_17973,N_17768,N_17919);
nor U17974 (N_17974,N_17797,N_17888);
xnor U17975 (N_17975,N_17807,N_17892);
or U17976 (N_17976,N_17848,N_17779);
nor U17977 (N_17977,N_17858,N_17875);
or U17978 (N_17978,N_17781,N_17808);
or U17979 (N_17979,N_17831,N_17799);
nand U17980 (N_17980,N_17857,N_17862);
nor U17981 (N_17981,N_17788,N_17778);
xnor U17982 (N_17982,N_17912,N_17887);
and U17983 (N_17983,N_17863,N_17898);
xor U17984 (N_17984,N_17846,N_17874);
nor U17985 (N_17985,N_17821,N_17851);
nor U17986 (N_17986,N_17845,N_17771);
or U17987 (N_17987,N_17873,N_17836);
nand U17988 (N_17988,N_17841,N_17899);
and U17989 (N_17989,N_17834,N_17908);
and U17990 (N_17990,N_17864,N_17812);
and U17991 (N_17991,N_17916,N_17792);
nor U17992 (N_17992,N_17815,N_17883);
xnor U17993 (N_17993,N_17893,N_17782);
xor U17994 (N_17994,N_17817,N_17800);
xnor U17995 (N_17995,N_17827,N_17868);
and U17996 (N_17996,N_17910,N_17814);
and U17997 (N_17997,N_17770,N_17839);
nor U17998 (N_17998,N_17773,N_17884);
nor U17999 (N_17999,N_17866,N_17915);
nor U18000 (N_18000,N_17875,N_17764);
and U18001 (N_18001,N_17848,N_17859);
nor U18002 (N_18002,N_17878,N_17863);
or U18003 (N_18003,N_17881,N_17884);
xnor U18004 (N_18004,N_17861,N_17902);
or U18005 (N_18005,N_17904,N_17809);
xor U18006 (N_18006,N_17846,N_17763);
nor U18007 (N_18007,N_17804,N_17786);
nand U18008 (N_18008,N_17811,N_17797);
or U18009 (N_18009,N_17782,N_17865);
or U18010 (N_18010,N_17837,N_17796);
nand U18011 (N_18011,N_17882,N_17903);
or U18012 (N_18012,N_17833,N_17770);
nand U18013 (N_18013,N_17867,N_17836);
nor U18014 (N_18014,N_17848,N_17885);
or U18015 (N_18015,N_17900,N_17889);
or U18016 (N_18016,N_17800,N_17792);
nand U18017 (N_18017,N_17902,N_17795);
xor U18018 (N_18018,N_17833,N_17827);
or U18019 (N_18019,N_17827,N_17849);
nand U18020 (N_18020,N_17898,N_17761);
or U18021 (N_18021,N_17782,N_17797);
or U18022 (N_18022,N_17810,N_17776);
xnor U18023 (N_18023,N_17801,N_17888);
nand U18024 (N_18024,N_17803,N_17810);
nand U18025 (N_18025,N_17777,N_17899);
nor U18026 (N_18026,N_17853,N_17822);
xor U18027 (N_18027,N_17916,N_17826);
and U18028 (N_18028,N_17825,N_17864);
or U18029 (N_18029,N_17773,N_17842);
or U18030 (N_18030,N_17888,N_17859);
or U18031 (N_18031,N_17875,N_17813);
or U18032 (N_18032,N_17899,N_17864);
xnor U18033 (N_18033,N_17819,N_17869);
or U18034 (N_18034,N_17898,N_17795);
nor U18035 (N_18035,N_17772,N_17822);
nor U18036 (N_18036,N_17861,N_17891);
and U18037 (N_18037,N_17813,N_17803);
and U18038 (N_18038,N_17851,N_17828);
nor U18039 (N_18039,N_17792,N_17798);
xnor U18040 (N_18040,N_17800,N_17805);
and U18041 (N_18041,N_17909,N_17824);
nor U18042 (N_18042,N_17763,N_17906);
or U18043 (N_18043,N_17899,N_17859);
nor U18044 (N_18044,N_17818,N_17842);
or U18045 (N_18045,N_17803,N_17914);
and U18046 (N_18046,N_17852,N_17868);
nand U18047 (N_18047,N_17864,N_17901);
or U18048 (N_18048,N_17880,N_17841);
nor U18049 (N_18049,N_17907,N_17791);
xor U18050 (N_18050,N_17792,N_17892);
and U18051 (N_18051,N_17793,N_17913);
nand U18052 (N_18052,N_17868,N_17874);
and U18053 (N_18053,N_17799,N_17854);
xnor U18054 (N_18054,N_17837,N_17835);
xnor U18055 (N_18055,N_17886,N_17919);
nand U18056 (N_18056,N_17852,N_17911);
nor U18057 (N_18057,N_17881,N_17816);
xnor U18058 (N_18058,N_17772,N_17917);
nor U18059 (N_18059,N_17883,N_17886);
or U18060 (N_18060,N_17791,N_17771);
xor U18061 (N_18061,N_17812,N_17813);
xnor U18062 (N_18062,N_17851,N_17808);
or U18063 (N_18063,N_17768,N_17887);
nand U18064 (N_18064,N_17792,N_17789);
and U18065 (N_18065,N_17817,N_17812);
and U18066 (N_18066,N_17766,N_17775);
xnor U18067 (N_18067,N_17775,N_17910);
nor U18068 (N_18068,N_17885,N_17891);
xor U18069 (N_18069,N_17789,N_17841);
or U18070 (N_18070,N_17898,N_17919);
or U18071 (N_18071,N_17858,N_17814);
xnor U18072 (N_18072,N_17857,N_17775);
nand U18073 (N_18073,N_17890,N_17856);
xnor U18074 (N_18074,N_17918,N_17795);
nor U18075 (N_18075,N_17804,N_17780);
and U18076 (N_18076,N_17849,N_17798);
nand U18077 (N_18077,N_17839,N_17914);
xor U18078 (N_18078,N_17806,N_17849);
or U18079 (N_18079,N_17798,N_17874);
xnor U18080 (N_18080,N_18077,N_18063);
and U18081 (N_18081,N_18070,N_17994);
nand U18082 (N_18082,N_18076,N_17998);
and U18083 (N_18083,N_17997,N_18007);
nor U18084 (N_18084,N_18035,N_18011);
xor U18085 (N_18085,N_18003,N_17965);
nor U18086 (N_18086,N_17985,N_18064);
nand U18087 (N_18087,N_18013,N_18023);
or U18088 (N_18088,N_17986,N_18051);
and U18089 (N_18089,N_18019,N_17927);
and U18090 (N_18090,N_18024,N_18078);
and U18091 (N_18091,N_17969,N_18054);
nand U18092 (N_18092,N_17932,N_17934);
and U18093 (N_18093,N_17936,N_18071);
nand U18094 (N_18094,N_17941,N_18052);
xnor U18095 (N_18095,N_18038,N_17982);
or U18096 (N_18096,N_17926,N_17968);
and U18097 (N_18097,N_17970,N_18001);
nand U18098 (N_18098,N_17981,N_18039);
nand U18099 (N_18099,N_18066,N_17973);
xnor U18100 (N_18100,N_17975,N_17937);
and U18101 (N_18101,N_17991,N_17939);
or U18102 (N_18102,N_18042,N_18058);
or U18103 (N_18103,N_18057,N_18074);
xnor U18104 (N_18104,N_18041,N_18020);
nor U18105 (N_18105,N_18016,N_17952);
nand U18106 (N_18106,N_18073,N_18034);
xnor U18107 (N_18107,N_18055,N_18062);
or U18108 (N_18108,N_17955,N_18032);
nor U18109 (N_18109,N_17929,N_18018);
nor U18110 (N_18110,N_17987,N_17928);
or U18111 (N_18111,N_18008,N_17950);
nor U18112 (N_18112,N_17958,N_17954);
nor U18113 (N_18113,N_17942,N_17977);
and U18114 (N_18114,N_18045,N_18050);
and U18115 (N_18115,N_17978,N_17966);
xnor U18116 (N_18116,N_18014,N_18069);
xor U18117 (N_18117,N_17930,N_18036);
nand U18118 (N_18118,N_17979,N_17940);
nor U18119 (N_18119,N_17996,N_17963);
and U18120 (N_18120,N_17971,N_17974);
or U18121 (N_18121,N_18017,N_17989);
nand U18122 (N_18122,N_18060,N_17925);
xnor U18123 (N_18123,N_18009,N_18030);
nor U18124 (N_18124,N_18040,N_17960);
xnor U18125 (N_18125,N_18010,N_18015);
or U18126 (N_18126,N_18043,N_18037);
nand U18127 (N_18127,N_18065,N_17938);
nor U18128 (N_18128,N_18059,N_17953);
and U18129 (N_18129,N_18025,N_17923);
and U18130 (N_18130,N_17946,N_18033);
xnor U18131 (N_18131,N_18072,N_17972);
xnor U18132 (N_18132,N_18021,N_17957);
and U18133 (N_18133,N_17933,N_18026);
nand U18134 (N_18134,N_18002,N_18068);
or U18135 (N_18135,N_18022,N_18056);
nor U18136 (N_18136,N_17948,N_17944);
nor U18137 (N_18137,N_17959,N_18029);
nor U18138 (N_18138,N_18061,N_17931);
xor U18139 (N_18139,N_17999,N_17980);
or U18140 (N_18140,N_17964,N_18067);
and U18141 (N_18141,N_17935,N_18053);
xnor U18142 (N_18142,N_17983,N_18048);
xor U18143 (N_18143,N_17990,N_18006);
and U18144 (N_18144,N_17921,N_18046);
xnor U18145 (N_18145,N_18005,N_18012);
nor U18146 (N_18146,N_17988,N_18079);
nand U18147 (N_18147,N_17992,N_18049);
nand U18148 (N_18148,N_17961,N_17967);
or U18149 (N_18149,N_17951,N_18004);
or U18150 (N_18150,N_17976,N_18031);
nand U18151 (N_18151,N_17945,N_18027);
nand U18152 (N_18152,N_18028,N_18044);
nor U18153 (N_18153,N_17984,N_17920);
or U18154 (N_18154,N_18047,N_17943);
xnor U18155 (N_18155,N_17962,N_17949);
or U18156 (N_18156,N_17956,N_17924);
xor U18157 (N_18157,N_17995,N_18000);
nand U18158 (N_18158,N_17993,N_17922);
or U18159 (N_18159,N_18075,N_17947);
xor U18160 (N_18160,N_17922,N_18045);
nand U18161 (N_18161,N_18032,N_17971);
and U18162 (N_18162,N_18029,N_17990);
xor U18163 (N_18163,N_17947,N_18055);
nor U18164 (N_18164,N_18065,N_17947);
xnor U18165 (N_18165,N_17946,N_18028);
and U18166 (N_18166,N_18047,N_17932);
or U18167 (N_18167,N_17926,N_17932);
xor U18168 (N_18168,N_17963,N_18021);
nand U18169 (N_18169,N_18017,N_17955);
and U18170 (N_18170,N_18058,N_17965);
nand U18171 (N_18171,N_18008,N_17965);
or U18172 (N_18172,N_18062,N_17984);
xor U18173 (N_18173,N_18073,N_17955);
and U18174 (N_18174,N_17940,N_17968);
xor U18175 (N_18175,N_17965,N_18020);
xor U18176 (N_18176,N_18062,N_18022);
or U18177 (N_18177,N_18000,N_18052);
nand U18178 (N_18178,N_18045,N_18004);
xnor U18179 (N_18179,N_17988,N_18071);
and U18180 (N_18180,N_17939,N_18002);
nand U18181 (N_18181,N_18054,N_17946);
xnor U18182 (N_18182,N_17951,N_17942);
nor U18183 (N_18183,N_18061,N_18020);
nand U18184 (N_18184,N_18061,N_17990);
nand U18185 (N_18185,N_18062,N_18048);
xnor U18186 (N_18186,N_17967,N_17971);
nor U18187 (N_18187,N_18012,N_18040);
xor U18188 (N_18188,N_18031,N_18009);
nand U18189 (N_18189,N_18050,N_18030);
and U18190 (N_18190,N_17978,N_17988);
or U18191 (N_18191,N_17965,N_17921);
nand U18192 (N_18192,N_18046,N_17948);
nand U18193 (N_18193,N_17952,N_18008);
nand U18194 (N_18194,N_17943,N_17931);
or U18195 (N_18195,N_17980,N_18057);
nand U18196 (N_18196,N_17992,N_17988);
nor U18197 (N_18197,N_17971,N_18058);
and U18198 (N_18198,N_17992,N_17996);
xor U18199 (N_18199,N_18003,N_17936);
or U18200 (N_18200,N_18066,N_17971);
nand U18201 (N_18201,N_17948,N_17984);
and U18202 (N_18202,N_17989,N_18000);
xnor U18203 (N_18203,N_17973,N_17942);
or U18204 (N_18204,N_18020,N_18073);
nand U18205 (N_18205,N_17922,N_18002);
nand U18206 (N_18206,N_17988,N_17970);
nor U18207 (N_18207,N_18025,N_18006);
nor U18208 (N_18208,N_17947,N_18051);
nand U18209 (N_18209,N_18064,N_18028);
nand U18210 (N_18210,N_17999,N_17920);
and U18211 (N_18211,N_18059,N_17936);
xnor U18212 (N_18212,N_17951,N_17944);
nand U18213 (N_18213,N_18004,N_18058);
nor U18214 (N_18214,N_18020,N_18051);
and U18215 (N_18215,N_17933,N_18050);
nor U18216 (N_18216,N_18039,N_17987);
xnor U18217 (N_18217,N_18025,N_18054);
or U18218 (N_18218,N_17991,N_17996);
nor U18219 (N_18219,N_18064,N_18020);
nor U18220 (N_18220,N_17991,N_17945);
and U18221 (N_18221,N_18061,N_17926);
and U18222 (N_18222,N_17943,N_17982);
or U18223 (N_18223,N_17954,N_17988);
or U18224 (N_18224,N_18077,N_18016);
and U18225 (N_18225,N_17964,N_18053);
xnor U18226 (N_18226,N_18059,N_18069);
nand U18227 (N_18227,N_18054,N_17934);
nand U18228 (N_18228,N_17978,N_18004);
nand U18229 (N_18229,N_18038,N_18041);
and U18230 (N_18230,N_18074,N_17972);
nor U18231 (N_18231,N_17936,N_18004);
xnor U18232 (N_18232,N_17951,N_18077);
and U18233 (N_18233,N_17980,N_17962);
or U18234 (N_18234,N_18043,N_18069);
nor U18235 (N_18235,N_17949,N_17946);
nand U18236 (N_18236,N_17940,N_18045);
xor U18237 (N_18237,N_18069,N_17959);
nand U18238 (N_18238,N_18077,N_18019);
nor U18239 (N_18239,N_18014,N_18074);
xor U18240 (N_18240,N_18131,N_18195);
nor U18241 (N_18241,N_18116,N_18175);
nand U18242 (N_18242,N_18139,N_18124);
nor U18243 (N_18243,N_18083,N_18089);
and U18244 (N_18244,N_18112,N_18093);
xnor U18245 (N_18245,N_18162,N_18214);
xnor U18246 (N_18246,N_18199,N_18163);
or U18247 (N_18247,N_18166,N_18239);
and U18248 (N_18248,N_18188,N_18187);
xor U18249 (N_18249,N_18227,N_18117);
nor U18250 (N_18250,N_18122,N_18111);
nor U18251 (N_18251,N_18150,N_18103);
nor U18252 (N_18252,N_18109,N_18123);
or U18253 (N_18253,N_18184,N_18129);
or U18254 (N_18254,N_18107,N_18161);
or U18255 (N_18255,N_18233,N_18194);
nand U18256 (N_18256,N_18237,N_18196);
xor U18257 (N_18257,N_18222,N_18105);
xor U18258 (N_18258,N_18095,N_18177);
xor U18259 (N_18259,N_18203,N_18171);
nand U18260 (N_18260,N_18114,N_18091);
and U18261 (N_18261,N_18197,N_18178);
xnor U18262 (N_18262,N_18088,N_18154);
nand U18263 (N_18263,N_18113,N_18145);
xnor U18264 (N_18264,N_18101,N_18208);
and U18265 (N_18265,N_18179,N_18225);
nand U18266 (N_18266,N_18192,N_18229);
nor U18267 (N_18267,N_18102,N_18128);
xnor U18268 (N_18268,N_18118,N_18094);
and U18269 (N_18269,N_18223,N_18115);
and U18270 (N_18270,N_18085,N_18169);
nor U18271 (N_18271,N_18183,N_18164);
or U18272 (N_18272,N_18167,N_18147);
or U18273 (N_18273,N_18104,N_18182);
nor U18274 (N_18274,N_18200,N_18236);
nand U18275 (N_18275,N_18228,N_18159);
nand U18276 (N_18276,N_18216,N_18207);
nor U18277 (N_18277,N_18141,N_18081);
nor U18278 (N_18278,N_18148,N_18120);
nand U18279 (N_18279,N_18098,N_18151);
xnor U18280 (N_18280,N_18137,N_18180);
or U18281 (N_18281,N_18080,N_18209);
or U18282 (N_18282,N_18217,N_18092);
nor U18283 (N_18283,N_18082,N_18153);
and U18284 (N_18284,N_18130,N_18218);
or U18285 (N_18285,N_18173,N_18108);
and U18286 (N_18286,N_18176,N_18143);
and U18287 (N_18287,N_18136,N_18157);
nand U18288 (N_18288,N_18230,N_18186);
nand U18289 (N_18289,N_18125,N_18099);
and U18290 (N_18290,N_18231,N_18174);
xnor U18291 (N_18291,N_18198,N_18205);
or U18292 (N_18292,N_18213,N_18168);
nor U18293 (N_18293,N_18106,N_18096);
and U18294 (N_18294,N_18146,N_18158);
or U18295 (N_18295,N_18155,N_18238);
xor U18296 (N_18296,N_18220,N_18152);
xor U18297 (N_18297,N_18193,N_18086);
xor U18298 (N_18298,N_18189,N_18127);
nor U18299 (N_18299,N_18234,N_18170);
nand U18300 (N_18300,N_18185,N_18206);
nand U18301 (N_18301,N_18165,N_18126);
nor U18302 (N_18302,N_18140,N_18119);
and U18303 (N_18303,N_18211,N_18156);
and U18304 (N_18304,N_18134,N_18160);
nand U18305 (N_18305,N_18138,N_18224);
nand U18306 (N_18306,N_18135,N_18190);
and U18307 (N_18307,N_18144,N_18215);
nand U18308 (N_18308,N_18191,N_18221);
nand U18309 (N_18309,N_18097,N_18133);
or U18310 (N_18310,N_18132,N_18100);
and U18311 (N_18311,N_18235,N_18172);
nand U18312 (N_18312,N_18204,N_18110);
xor U18313 (N_18313,N_18142,N_18181);
or U18314 (N_18314,N_18232,N_18210);
or U18315 (N_18315,N_18212,N_18219);
xor U18316 (N_18316,N_18226,N_18087);
and U18317 (N_18317,N_18090,N_18149);
and U18318 (N_18318,N_18201,N_18202);
and U18319 (N_18319,N_18084,N_18121);
and U18320 (N_18320,N_18189,N_18166);
or U18321 (N_18321,N_18236,N_18145);
and U18322 (N_18322,N_18189,N_18223);
or U18323 (N_18323,N_18139,N_18211);
or U18324 (N_18324,N_18122,N_18198);
or U18325 (N_18325,N_18139,N_18169);
nor U18326 (N_18326,N_18171,N_18176);
nand U18327 (N_18327,N_18157,N_18171);
xnor U18328 (N_18328,N_18165,N_18142);
xor U18329 (N_18329,N_18232,N_18112);
nand U18330 (N_18330,N_18149,N_18151);
nand U18331 (N_18331,N_18089,N_18180);
xor U18332 (N_18332,N_18197,N_18172);
nand U18333 (N_18333,N_18194,N_18161);
and U18334 (N_18334,N_18094,N_18147);
xor U18335 (N_18335,N_18131,N_18113);
or U18336 (N_18336,N_18142,N_18084);
nand U18337 (N_18337,N_18130,N_18217);
or U18338 (N_18338,N_18145,N_18152);
nor U18339 (N_18339,N_18146,N_18215);
nor U18340 (N_18340,N_18163,N_18181);
nand U18341 (N_18341,N_18119,N_18206);
nor U18342 (N_18342,N_18174,N_18135);
xnor U18343 (N_18343,N_18136,N_18084);
and U18344 (N_18344,N_18110,N_18208);
nor U18345 (N_18345,N_18114,N_18220);
nand U18346 (N_18346,N_18145,N_18177);
or U18347 (N_18347,N_18164,N_18143);
or U18348 (N_18348,N_18209,N_18108);
nand U18349 (N_18349,N_18219,N_18142);
nor U18350 (N_18350,N_18164,N_18081);
and U18351 (N_18351,N_18215,N_18225);
and U18352 (N_18352,N_18214,N_18118);
nand U18353 (N_18353,N_18108,N_18092);
nor U18354 (N_18354,N_18150,N_18142);
or U18355 (N_18355,N_18130,N_18171);
or U18356 (N_18356,N_18124,N_18167);
xor U18357 (N_18357,N_18154,N_18184);
or U18358 (N_18358,N_18216,N_18184);
nor U18359 (N_18359,N_18196,N_18186);
nor U18360 (N_18360,N_18095,N_18112);
xnor U18361 (N_18361,N_18232,N_18207);
nand U18362 (N_18362,N_18147,N_18198);
nand U18363 (N_18363,N_18215,N_18162);
and U18364 (N_18364,N_18138,N_18126);
nand U18365 (N_18365,N_18152,N_18182);
nor U18366 (N_18366,N_18224,N_18204);
or U18367 (N_18367,N_18089,N_18090);
xnor U18368 (N_18368,N_18128,N_18233);
nor U18369 (N_18369,N_18129,N_18166);
nor U18370 (N_18370,N_18232,N_18204);
or U18371 (N_18371,N_18107,N_18239);
nand U18372 (N_18372,N_18153,N_18221);
and U18373 (N_18373,N_18106,N_18177);
and U18374 (N_18374,N_18203,N_18118);
nand U18375 (N_18375,N_18177,N_18088);
xnor U18376 (N_18376,N_18224,N_18187);
xor U18377 (N_18377,N_18230,N_18205);
xor U18378 (N_18378,N_18133,N_18177);
or U18379 (N_18379,N_18117,N_18132);
or U18380 (N_18380,N_18160,N_18101);
or U18381 (N_18381,N_18140,N_18157);
and U18382 (N_18382,N_18148,N_18105);
nor U18383 (N_18383,N_18194,N_18162);
and U18384 (N_18384,N_18161,N_18196);
nor U18385 (N_18385,N_18190,N_18092);
nor U18386 (N_18386,N_18235,N_18191);
or U18387 (N_18387,N_18157,N_18170);
nor U18388 (N_18388,N_18133,N_18178);
nand U18389 (N_18389,N_18152,N_18203);
nor U18390 (N_18390,N_18217,N_18097);
and U18391 (N_18391,N_18159,N_18089);
and U18392 (N_18392,N_18177,N_18100);
xnor U18393 (N_18393,N_18117,N_18131);
and U18394 (N_18394,N_18107,N_18216);
xnor U18395 (N_18395,N_18228,N_18238);
xor U18396 (N_18396,N_18103,N_18217);
nor U18397 (N_18397,N_18219,N_18149);
xnor U18398 (N_18398,N_18134,N_18216);
or U18399 (N_18399,N_18142,N_18125);
or U18400 (N_18400,N_18279,N_18321);
nor U18401 (N_18401,N_18386,N_18314);
nand U18402 (N_18402,N_18381,N_18278);
xnor U18403 (N_18403,N_18329,N_18343);
xor U18404 (N_18404,N_18356,N_18241);
xnor U18405 (N_18405,N_18303,N_18277);
and U18406 (N_18406,N_18371,N_18384);
or U18407 (N_18407,N_18360,N_18370);
nand U18408 (N_18408,N_18297,N_18281);
or U18409 (N_18409,N_18262,N_18245);
xor U18410 (N_18410,N_18358,N_18289);
nor U18411 (N_18411,N_18319,N_18292);
or U18412 (N_18412,N_18256,N_18252);
nand U18413 (N_18413,N_18270,N_18246);
xor U18414 (N_18414,N_18389,N_18379);
nor U18415 (N_18415,N_18305,N_18257);
xnor U18416 (N_18416,N_18249,N_18274);
nand U18417 (N_18417,N_18363,N_18337);
xnor U18418 (N_18418,N_18325,N_18380);
or U18419 (N_18419,N_18395,N_18397);
xnor U18420 (N_18420,N_18273,N_18272);
xnor U18421 (N_18421,N_18344,N_18317);
or U18422 (N_18422,N_18383,N_18283);
nor U18423 (N_18423,N_18394,N_18374);
nor U18424 (N_18424,N_18365,N_18318);
xor U18425 (N_18425,N_18250,N_18393);
xor U18426 (N_18426,N_18323,N_18316);
xor U18427 (N_18427,N_18324,N_18280);
nor U18428 (N_18428,N_18275,N_18385);
or U18429 (N_18429,N_18340,N_18351);
nand U18430 (N_18430,N_18296,N_18290);
nand U18431 (N_18431,N_18350,N_18285);
nor U18432 (N_18432,N_18251,N_18352);
and U18433 (N_18433,N_18311,N_18342);
and U18434 (N_18434,N_18254,N_18240);
nor U18435 (N_18435,N_18267,N_18286);
nor U18436 (N_18436,N_18266,N_18331);
and U18437 (N_18437,N_18353,N_18320);
xor U18438 (N_18438,N_18261,N_18333);
or U18439 (N_18439,N_18347,N_18387);
xor U18440 (N_18440,N_18312,N_18396);
or U18441 (N_18441,N_18243,N_18315);
nor U18442 (N_18442,N_18295,N_18359);
xnor U18443 (N_18443,N_18349,N_18302);
nand U18444 (N_18444,N_18260,N_18300);
xor U18445 (N_18445,N_18391,N_18265);
nand U18446 (N_18446,N_18309,N_18377);
nor U18447 (N_18447,N_18287,N_18330);
nor U18448 (N_18448,N_18293,N_18392);
xnor U18449 (N_18449,N_18372,N_18294);
nor U18450 (N_18450,N_18247,N_18264);
or U18451 (N_18451,N_18339,N_18269);
nor U18452 (N_18452,N_18354,N_18334);
or U18453 (N_18453,N_18304,N_18332);
xnor U18454 (N_18454,N_18368,N_18366);
nand U18455 (N_18455,N_18362,N_18284);
and U18456 (N_18456,N_18307,N_18375);
or U18457 (N_18457,N_18306,N_18376);
xnor U18458 (N_18458,N_18364,N_18242);
xnor U18459 (N_18459,N_18336,N_18301);
xnor U18460 (N_18460,N_18382,N_18361);
and U18461 (N_18461,N_18348,N_18345);
and U18462 (N_18462,N_18357,N_18355);
nor U18463 (N_18463,N_18268,N_18369);
xnor U18464 (N_18464,N_18291,N_18378);
xnor U18465 (N_18465,N_18398,N_18341);
nand U18466 (N_18466,N_18248,N_18253);
or U18467 (N_18467,N_18276,N_18298);
nor U18468 (N_18468,N_18367,N_18326);
and U18469 (N_18469,N_18263,N_18322);
and U18470 (N_18470,N_18373,N_18258);
and U18471 (N_18471,N_18299,N_18310);
nand U18472 (N_18472,N_18255,N_18313);
nand U18473 (N_18473,N_18335,N_18338);
nand U18474 (N_18474,N_18346,N_18259);
nor U18475 (N_18475,N_18327,N_18288);
xnor U18476 (N_18476,N_18308,N_18244);
or U18477 (N_18477,N_18390,N_18399);
xnor U18478 (N_18478,N_18282,N_18328);
or U18479 (N_18479,N_18388,N_18271);
nand U18480 (N_18480,N_18339,N_18384);
nor U18481 (N_18481,N_18273,N_18346);
or U18482 (N_18482,N_18392,N_18354);
and U18483 (N_18483,N_18375,N_18330);
and U18484 (N_18484,N_18242,N_18393);
and U18485 (N_18485,N_18325,N_18346);
or U18486 (N_18486,N_18322,N_18256);
and U18487 (N_18487,N_18259,N_18329);
nand U18488 (N_18488,N_18260,N_18259);
nand U18489 (N_18489,N_18340,N_18301);
xnor U18490 (N_18490,N_18312,N_18391);
or U18491 (N_18491,N_18350,N_18363);
nor U18492 (N_18492,N_18299,N_18325);
nor U18493 (N_18493,N_18364,N_18388);
nand U18494 (N_18494,N_18281,N_18305);
and U18495 (N_18495,N_18360,N_18332);
and U18496 (N_18496,N_18365,N_18393);
and U18497 (N_18497,N_18392,N_18289);
nand U18498 (N_18498,N_18327,N_18353);
nand U18499 (N_18499,N_18361,N_18264);
or U18500 (N_18500,N_18332,N_18286);
and U18501 (N_18501,N_18348,N_18350);
and U18502 (N_18502,N_18332,N_18289);
or U18503 (N_18503,N_18355,N_18364);
xor U18504 (N_18504,N_18305,N_18288);
and U18505 (N_18505,N_18361,N_18244);
or U18506 (N_18506,N_18345,N_18248);
nand U18507 (N_18507,N_18324,N_18245);
and U18508 (N_18508,N_18358,N_18354);
nor U18509 (N_18509,N_18302,N_18274);
nand U18510 (N_18510,N_18255,N_18372);
or U18511 (N_18511,N_18304,N_18347);
nor U18512 (N_18512,N_18265,N_18244);
or U18513 (N_18513,N_18341,N_18319);
xor U18514 (N_18514,N_18314,N_18334);
and U18515 (N_18515,N_18272,N_18314);
nor U18516 (N_18516,N_18277,N_18347);
nand U18517 (N_18517,N_18317,N_18318);
xnor U18518 (N_18518,N_18263,N_18313);
nand U18519 (N_18519,N_18342,N_18329);
nor U18520 (N_18520,N_18259,N_18307);
xor U18521 (N_18521,N_18352,N_18343);
nand U18522 (N_18522,N_18271,N_18275);
and U18523 (N_18523,N_18294,N_18350);
xor U18524 (N_18524,N_18250,N_18391);
xnor U18525 (N_18525,N_18349,N_18364);
xor U18526 (N_18526,N_18349,N_18312);
xnor U18527 (N_18527,N_18329,N_18241);
nand U18528 (N_18528,N_18299,N_18323);
nor U18529 (N_18529,N_18370,N_18371);
nor U18530 (N_18530,N_18385,N_18375);
and U18531 (N_18531,N_18337,N_18302);
nor U18532 (N_18532,N_18393,N_18390);
nor U18533 (N_18533,N_18300,N_18313);
nand U18534 (N_18534,N_18381,N_18266);
nand U18535 (N_18535,N_18297,N_18354);
nor U18536 (N_18536,N_18390,N_18275);
or U18537 (N_18537,N_18300,N_18254);
nor U18538 (N_18538,N_18379,N_18386);
nor U18539 (N_18539,N_18266,N_18242);
xnor U18540 (N_18540,N_18258,N_18296);
nand U18541 (N_18541,N_18246,N_18299);
xnor U18542 (N_18542,N_18316,N_18258);
or U18543 (N_18543,N_18348,N_18366);
or U18544 (N_18544,N_18398,N_18266);
nand U18545 (N_18545,N_18246,N_18348);
and U18546 (N_18546,N_18349,N_18287);
nand U18547 (N_18547,N_18359,N_18340);
xor U18548 (N_18548,N_18247,N_18366);
or U18549 (N_18549,N_18293,N_18380);
xnor U18550 (N_18550,N_18315,N_18321);
nand U18551 (N_18551,N_18370,N_18361);
nand U18552 (N_18552,N_18380,N_18306);
nand U18553 (N_18553,N_18348,N_18285);
xnor U18554 (N_18554,N_18374,N_18373);
or U18555 (N_18555,N_18396,N_18395);
xor U18556 (N_18556,N_18274,N_18361);
or U18557 (N_18557,N_18263,N_18257);
or U18558 (N_18558,N_18379,N_18392);
nor U18559 (N_18559,N_18317,N_18336);
and U18560 (N_18560,N_18453,N_18430);
and U18561 (N_18561,N_18439,N_18474);
and U18562 (N_18562,N_18436,N_18419);
and U18563 (N_18563,N_18437,N_18492);
nand U18564 (N_18564,N_18410,N_18432);
xnor U18565 (N_18565,N_18460,N_18417);
or U18566 (N_18566,N_18493,N_18501);
xnor U18567 (N_18567,N_18498,N_18479);
or U18568 (N_18568,N_18495,N_18409);
and U18569 (N_18569,N_18520,N_18444);
or U18570 (N_18570,N_18447,N_18431);
and U18571 (N_18571,N_18523,N_18408);
or U18572 (N_18572,N_18536,N_18557);
nor U18573 (N_18573,N_18477,N_18551);
xor U18574 (N_18574,N_18464,N_18509);
nor U18575 (N_18575,N_18530,N_18525);
nand U18576 (N_18576,N_18438,N_18426);
nand U18577 (N_18577,N_18500,N_18440);
xnor U18578 (N_18578,N_18559,N_18508);
nor U18579 (N_18579,N_18471,N_18484);
xnor U18580 (N_18580,N_18516,N_18405);
nand U18581 (N_18581,N_18402,N_18496);
nand U18582 (N_18582,N_18415,N_18537);
nand U18583 (N_18583,N_18465,N_18543);
and U18584 (N_18584,N_18433,N_18450);
or U18585 (N_18585,N_18485,N_18411);
nor U18586 (N_18586,N_18448,N_18552);
nor U18587 (N_18587,N_18504,N_18519);
nor U18588 (N_18588,N_18442,N_18503);
nor U18589 (N_18589,N_18494,N_18400);
or U18590 (N_18590,N_18497,N_18549);
xnor U18591 (N_18591,N_18434,N_18488);
xnor U18592 (N_18592,N_18429,N_18507);
nand U18593 (N_18593,N_18499,N_18462);
nand U18594 (N_18594,N_18445,N_18540);
or U18595 (N_18595,N_18468,N_18527);
nor U18596 (N_18596,N_18542,N_18534);
and U18597 (N_18597,N_18478,N_18418);
xnor U18598 (N_18598,N_18533,N_18441);
or U18599 (N_18599,N_18451,N_18489);
and U18600 (N_18600,N_18476,N_18443);
and U18601 (N_18601,N_18556,N_18461);
and U18602 (N_18602,N_18452,N_18518);
and U18603 (N_18603,N_18514,N_18469);
nor U18604 (N_18604,N_18463,N_18524);
nor U18605 (N_18605,N_18473,N_18482);
nand U18606 (N_18606,N_18486,N_18475);
xor U18607 (N_18607,N_18406,N_18490);
and U18608 (N_18608,N_18420,N_18456);
nor U18609 (N_18609,N_18548,N_18425);
xor U18610 (N_18610,N_18555,N_18554);
nor U18611 (N_18611,N_18532,N_18428);
xor U18612 (N_18612,N_18422,N_18545);
or U18613 (N_18613,N_18423,N_18459);
xnor U18614 (N_18614,N_18470,N_18421);
nor U18615 (N_18615,N_18412,N_18513);
and U18616 (N_18616,N_18517,N_18487);
and U18617 (N_18617,N_18550,N_18539);
xor U18618 (N_18618,N_18535,N_18491);
or U18619 (N_18619,N_18404,N_18522);
and U18620 (N_18620,N_18512,N_18407);
or U18621 (N_18621,N_18403,N_18414);
or U18622 (N_18622,N_18427,N_18454);
nor U18623 (N_18623,N_18511,N_18413);
nor U18624 (N_18624,N_18424,N_18458);
xor U18625 (N_18625,N_18528,N_18435);
and U18626 (N_18626,N_18521,N_18541);
nand U18627 (N_18627,N_18472,N_18502);
nor U18628 (N_18628,N_18558,N_18505);
and U18629 (N_18629,N_18515,N_18526);
nand U18630 (N_18630,N_18506,N_18481);
and U18631 (N_18631,N_18466,N_18531);
or U18632 (N_18632,N_18483,N_18467);
and U18633 (N_18633,N_18529,N_18446);
nand U18634 (N_18634,N_18480,N_18449);
and U18635 (N_18635,N_18416,N_18544);
nor U18636 (N_18636,N_18553,N_18510);
nand U18637 (N_18637,N_18547,N_18546);
xnor U18638 (N_18638,N_18401,N_18455);
or U18639 (N_18639,N_18538,N_18457);
xor U18640 (N_18640,N_18463,N_18416);
xnor U18641 (N_18641,N_18558,N_18472);
and U18642 (N_18642,N_18513,N_18473);
and U18643 (N_18643,N_18522,N_18519);
or U18644 (N_18644,N_18417,N_18506);
nor U18645 (N_18645,N_18435,N_18530);
or U18646 (N_18646,N_18426,N_18428);
or U18647 (N_18647,N_18402,N_18434);
and U18648 (N_18648,N_18412,N_18497);
or U18649 (N_18649,N_18536,N_18477);
xor U18650 (N_18650,N_18552,N_18453);
nand U18651 (N_18651,N_18451,N_18516);
or U18652 (N_18652,N_18533,N_18415);
nor U18653 (N_18653,N_18485,N_18450);
and U18654 (N_18654,N_18411,N_18502);
xor U18655 (N_18655,N_18423,N_18534);
or U18656 (N_18656,N_18422,N_18434);
nand U18657 (N_18657,N_18555,N_18412);
xor U18658 (N_18658,N_18467,N_18462);
nor U18659 (N_18659,N_18493,N_18414);
nand U18660 (N_18660,N_18412,N_18435);
or U18661 (N_18661,N_18440,N_18496);
nand U18662 (N_18662,N_18438,N_18423);
and U18663 (N_18663,N_18456,N_18507);
and U18664 (N_18664,N_18523,N_18514);
or U18665 (N_18665,N_18529,N_18547);
and U18666 (N_18666,N_18408,N_18437);
or U18667 (N_18667,N_18530,N_18452);
nor U18668 (N_18668,N_18552,N_18540);
nor U18669 (N_18669,N_18437,N_18524);
and U18670 (N_18670,N_18470,N_18505);
xnor U18671 (N_18671,N_18424,N_18400);
and U18672 (N_18672,N_18508,N_18496);
and U18673 (N_18673,N_18524,N_18502);
nand U18674 (N_18674,N_18557,N_18540);
xor U18675 (N_18675,N_18536,N_18450);
or U18676 (N_18676,N_18423,N_18484);
xnor U18677 (N_18677,N_18538,N_18428);
nor U18678 (N_18678,N_18401,N_18506);
or U18679 (N_18679,N_18402,N_18523);
and U18680 (N_18680,N_18547,N_18491);
or U18681 (N_18681,N_18445,N_18535);
xnor U18682 (N_18682,N_18463,N_18499);
nand U18683 (N_18683,N_18455,N_18501);
xor U18684 (N_18684,N_18541,N_18491);
nand U18685 (N_18685,N_18455,N_18534);
nor U18686 (N_18686,N_18559,N_18453);
xor U18687 (N_18687,N_18438,N_18515);
and U18688 (N_18688,N_18434,N_18432);
and U18689 (N_18689,N_18469,N_18509);
or U18690 (N_18690,N_18541,N_18488);
and U18691 (N_18691,N_18520,N_18419);
or U18692 (N_18692,N_18508,N_18549);
nor U18693 (N_18693,N_18427,N_18524);
or U18694 (N_18694,N_18493,N_18465);
nor U18695 (N_18695,N_18407,N_18467);
and U18696 (N_18696,N_18422,N_18499);
or U18697 (N_18697,N_18463,N_18504);
xor U18698 (N_18698,N_18538,N_18499);
xnor U18699 (N_18699,N_18407,N_18410);
nor U18700 (N_18700,N_18535,N_18456);
nor U18701 (N_18701,N_18486,N_18453);
or U18702 (N_18702,N_18455,N_18417);
or U18703 (N_18703,N_18405,N_18518);
or U18704 (N_18704,N_18457,N_18499);
or U18705 (N_18705,N_18411,N_18439);
and U18706 (N_18706,N_18431,N_18492);
and U18707 (N_18707,N_18401,N_18545);
nand U18708 (N_18708,N_18479,N_18456);
xor U18709 (N_18709,N_18544,N_18410);
xor U18710 (N_18710,N_18549,N_18435);
nor U18711 (N_18711,N_18471,N_18546);
nor U18712 (N_18712,N_18543,N_18508);
or U18713 (N_18713,N_18520,N_18431);
or U18714 (N_18714,N_18408,N_18548);
and U18715 (N_18715,N_18525,N_18517);
or U18716 (N_18716,N_18436,N_18555);
nand U18717 (N_18717,N_18410,N_18452);
or U18718 (N_18718,N_18536,N_18521);
xor U18719 (N_18719,N_18482,N_18498);
and U18720 (N_18720,N_18560,N_18589);
nand U18721 (N_18721,N_18713,N_18629);
and U18722 (N_18722,N_18717,N_18664);
nor U18723 (N_18723,N_18668,N_18711);
nand U18724 (N_18724,N_18604,N_18613);
or U18725 (N_18725,N_18635,N_18694);
or U18726 (N_18726,N_18619,N_18638);
nor U18727 (N_18727,N_18714,N_18590);
and U18728 (N_18728,N_18688,N_18612);
nand U18729 (N_18729,N_18696,N_18596);
and U18730 (N_18730,N_18577,N_18636);
or U18731 (N_18731,N_18665,N_18630);
nand U18732 (N_18732,N_18691,N_18655);
nor U18733 (N_18733,N_18606,N_18610);
xor U18734 (N_18734,N_18682,N_18661);
xnor U18735 (N_18735,N_18672,N_18680);
nand U18736 (N_18736,N_18616,N_18637);
or U18737 (N_18737,N_18686,N_18615);
nand U18738 (N_18738,N_18603,N_18670);
nand U18739 (N_18739,N_18667,N_18678);
xor U18740 (N_18740,N_18709,N_18685);
xnor U18741 (N_18741,N_18697,N_18654);
and U18742 (N_18742,N_18622,N_18653);
and U18743 (N_18743,N_18666,N_18611);
nor U18744 (N_18744,N_18689,N_18699);
or U18745 (N_18745,N_18585,N_18657);
xor U18746 (N_18746,N_18671,N_18599);
xnor U18747 (N_18747,N_18675,N_18574);
and U18748 (N_18748,N_18634,N_18624);
or U18749 (N_18749,N_18681,N_18712);
or U18750 (N_18750,N_18598,N_18602);
nand U18751 (N_18751,N_18702,N_18684);
xnor U18752 (N_18752,N_18593,N_18658);
nor U18753 (N_18753,N_18649,N_18707);
and U18754 (N_18754,N_18716,N_18564);
xor U18755 (N_18755,N_18627,N_18625);
nor U18756 (N_18756,N_18705,N_18633);
xnor U18757 (N_18757,N_18631,N_18597);
xor U18758 (N_18758,N_18591,N_18676);
nand U18759 (N_18759,N_18614,N_18663);
nand U18760 (N_18760,N_18648,N_18632);
xor U18761 (N_18761,N_18656,N_18623);
nand U18762 (N_18762,N_18645,N_18583);
nand U18763 (N_18763,N_18642,N_18592);
or U18764 (N_18764,N_18601,N_18572);
and U18765 (N_18765,N_18586,N_18660);
or U18766 (N_18766,N_18640,N_18659);
xnor U18767 (N_18767,N_18695,N_18573);
or U18768 (N_18768,N_18620,N_18690);
and U18769 (N_18769,N_18595,N_18669);
nor U18770 (N_18770,N_18571,N_18609);
nor U18771 (N_18771,N_18701,N_18562);
nand U18772 (N_18772,N_18650,N_18608);
and U18773 (N_18773,N_18567,N_18565);
or U18774 (N_18774,N_18651,N_18588);
or U18775 (N_18775,N_18710,N_18600);
nand U18776 (N_18776,N_18628,N_18706);
nor U18777 (N_18777,N_18580,N_18693);
nor U18778 (N_18778,N_18647,N_18579);
and U18779 (N_18779,N_18582,N_18662);
nand U18780 (N_18780,N_18674,N_18563);
or U18781 (N_18781,N_18584,N_18561);
and U18782 (N_18782,N_18646,N_18715);
nand U18783 (N_18783,N_18652,N_18576);
nor U18784 (N_18784,N_18617,N_18626);
and U18785 (N_18785,N_18692,N_18581);
or U18786 (N_18786,N_18703,N_18687);
or U18787 (N_18787,N_18621,N_18643);
nor U18788 (N_18788,N_18704,N_18569);
nor U18789 (N_18789,N_18618,N_18673);
and U18790 (N_18790,N_18708,N_18677);
and U18791 (N_18791,N_18644,N_18578);
nand U18792 (N_18792,N_18607,N_18566);
nor U18793 (N_18793,N_18594,N_18568);
nor U18794 (N_18794,N_18719,N_18683);
and U18795 (N_18795,N_18587,N_18570);
nor U18796 (N_18796,N_18700,N_18641);
nor U18797 (N_18797,N_18639,N_18718);
nand U18798 (N_18798,N_18679,N_18605);
nand U18799 (N_18799,N_18575,N_18698);
and U18800 (N_18800,N_18561,N_18699);
or U18801 (N_18801,N_18623,N_18673);
xor U18802 (N_18802,N_18632,N_18704);
xnor U18803 (N_18803,N_18683,N_18624);
nand U18804 (N_18804,N_18701,N_18694);
nor U18805 (N_18805,N_18656,N_18571);
and U18806 (N_18806,N_18658,N_18608);
and U18807 (N_18807,N_18709,N_18670);
or U18808 (N_18808,N_18582,N_18616);
and U18809 (N_18809,N_18709,N_18560);
nand U18810 (N_18810,N_18639,N_18626);
and U18811 (N_18811,N_18608,N_18620);
and U18812 (N_18812,N_18701,N_18586);
or U18813 (N_18813,N_18672,N_18649);
nor U18814 (N_18814,N_18683,N_18650);
nor U18815 (N_18815,N_18574,N_18605);
nor U18816 (N_18816,N_18704,N_18614);
or U18817 (N_18817,N_18597,N_18562);
and U18818 (N_18818,N_18648,N_18705);
nor U18819 (N_18819,N_18676,N_18588);
or U18820 (N_18820,N_18591,N_18657);
or U18821 (N_18821,N_18589,N_18641);
and U18822 (N_18822,N_18585,N_18627);
nand U18823 (N_18823,N_18705,N_18572);
nor U18824 (N_18824,N_18664,N_18649);
nor U18825 (N_18825,N_18703,N_18563);
and U18826 (N_18826,N_18635,N_18606);
and U18827 (N_18827,N_18641,N_18601);
or U18828 (N_18828,N_18672,N_18635);
or U18829 (N_18829,N_18574,N_18678);
xnor U18830 (N_18830,N_18691,N_18574);
and U18831 (N_18831,N_18667,N_18657);
or U18832 (N_18832,N_18674,N_18600);
xor U18833 (N_18833,N_18600,N_18670);
nor U18834 (N_18834,N_18645,N_18630);
nor U18835 (N_18835,N_18683,N_18642);
and U18836 (N_18836,N_18627,N_18633);
nand U18837 (N_18837,N_18664,N_18610);
and U18838 (N_18838,N_18649,N_18698);
or U18839 (N_18839,N_18564,N_18706);
nor U18840 (N_18840,N_18575,N_18561);
nor U18841 (N_18841,N_18706,N_18626);
xor U18842 (N_18842,N_18577,N_18612);
xnor U18843 (N_18843,N_18697,N_18638);
and U18844 (N_18844,N_18698,N_18579);
or U18845 (N_18845,N_18689,N_18560);
nor U18846 (N_18846,N_18571,N_18594);
and U18847 (N_18847,N_18697,N_18631);
nor U18848 (N_18848,N_18626,N_18694);
nand U18849 (N_18849,N_18592,N_18693);
or U18850 (N_18850,N_18587,N_18650);
nand U18851 (N_18851,N_18610,N_18671);
nor U18852 (N_18852,N_18684,N_18564);
xnor U18853 (N_18853,N_18654,N_18604);
nand U18854 (N_18854,N_18671,N_18653);
xor U18855 (N_18855,N_18661,N_18642);
nand U18856 (N_18856,N_18596,N_18641);
or U18857 (N_18857,N_18632,N_18609);
or U18858 (N_18858,N_18561,N_18649);
nand U18859 (N_18859,N_18625,N_18586);
or U18860 (N_18860,N_18592,N_18706);
nand U18861 (N_18861,N_18708,N_18580);
and U18862 (N_18862,N_18594,N_18662);
or U18863 (N_18863,N_18700,N_18703);
nand U18864 (N_18864,N_18688,N_18707);
xor U18865 (N_18865,N_18607,N_18575);
or U18866 (N_18866,N_18647,N_18696);
xnor U18867 (N_18867,N_18676,N_18580);
nor U18868 (N_18868,N_18662,N_18702);
and U18869 (N_18869,N_18707,N_18646);
and U18870 (N_18870,N_18560,N_18624);
or U18871 (N_18871,N_18596,N_18678);
xor U18872 (N_18872,N_18638,N_18695);
or U18873 (N_18873,N_18582,N_18585);
or U18874 (N_18874,N_18696,N_18646);
and U18875 (N_18875,N_18601,N_18634);
or U18876 (N_18876,N_18659,N_18623);
xor U18877 (N_18877,N_18610,N_18673);
nor U18878 (N_18878,N_18693,N_18602);
or U18879 (N_18879,N_18623,N_18641);
or U18880 (N_18880,N_18858,N_18786);
nor U18881 (N_18881,N_18765,N_18742);
nand U18882 (N_18882,N_18868,N_18741);
nor U18883 (N_18883,N_18877,N_18840);
and U18884 (N_18884,N_18736,N_18879);
nand U18885 (N_18885,N_18754,N_18874);
and U18886 (N_18886,N_18788,N_18819);
nor U18887 (N_18887,N_18813,N_18846);
nor U18888 (N_18888,N_18756,N_18771);
nor U18889 (N_18889,N_18810,N_18746);
or U18890 (N_18890,N_18811,N_18793);
and U18891 (N_18891,N_18854,N_18739);
xnor U18892 (N_18892,N_18804,N_18814);
or U18893 (N_18893,N_18850,N_18856);
xor U18894 (N_18894,N_18792,N_18835);
and U18895 (N_18895,N_18785,N_18729);
nand U18896 (N_18896,N_18799,N_18873);
nand U18897 (N_18897,N_18762,N_18735);
nor U18898 (N_18898,N_18875,N_18836);
nor U18899 (N_18899,N_18830,N_18767);
or U18900 (N_18900,N_18826,N_18829);
and U18901 (N_18901,N_18801,N_18779);
or U18902 (N_18902,N_18825,N_18800);
or U18903 (N_18903,N_18822,N_18798);
nand U18904 (N_18904,N_18748,N_18781);
and U18905 (N_18905,N_18838,N_18865);
xnor U18906 (N_18906,N_18761,N_18831);
nand U18907 (N_18907,N_18750,N_18720);
or U18908 (N_18908,N_18795,N_18853);
or U18909 (N_18909,N_18864,N_18727);
xnor U18910 (N_18910,N_18747,N_18818);
xor U18911 (N_18911,N_18851,N_18809);
xnor U18912 (N_18912,N_18731,N_18772);
xor U18913 (N_18913,N_18749,N_18844);
or U18914 (N_18914,N_18728,N_18721);
nand U18915 (N_18915,N_18872,N_18783);
nor U18916 (N_18916,N_18869,N_18732);
nor U18917 (N_18917,N_18845,N_18834);
nor U18918 (N_18918,N_18737,N_18808);
and U18919 (N_18919,N_18782,N_18774);
nand U18920 (N_18920,N_18841,N_18802);
xor U18921 (N_18921,N_18820,N_18796);
nand U18922 (N_18922,N_18866,N_18855);
nand U18923 (N_18923,N_18780,N_18862);
nor U18924 (N_18924,N_18770,N_18743);
and U18925 (N_18925,N_18817,N_18828);
or U18926 (N_18926,N_18751,N_18837);
xnor U18927 (N_18927,N_18784,N_18803);
nand U18928 (N_18928,N_18763,N_18876);
nor U18929 (N_18929,N_18753,N_18791);
nand U18930 (N_18930,N_18769,N_18734);
and U18931 (N_18931,N_18773,N_18815);
and U18932 (N_18932,N_18859,N_18733);
and U18933 (N_18933,N_18847,N_18861);
nor U18934 (N_18934,N_18863,N_18823);
nand U18935 (N_18935,N_18768,N_18755);
and U18936 (N_18936,N_18777,N_18775);
or U18937 (N_18937,N_18827,N_18832);
or U18938 (N_18938,N_18857,N_18878);
nor U18939 (N_18939,N_18724,N_18797);
nand U18940 (N_18940,N_18725,N_18760);
xor U18941 (N_18941,N_18849,N_18848);
xor U18942 (N_18942,N_18757,N_18789);
xor U18943 (N_18943,N_18744,N_18870);
xor U18944 (N_18944,N_18787,N_18843);
or U18945 (N_18945,N_18776,N_18812);
xnor U18946 (N_18946,N_18852,N_18758);
nor U18947 (N_18947,N_18726,N_18871);
nand U18948 (N_18948,N_18790,N_18806);
nor U18949 (N_18949,N_18821,N_18860);
nor U18950 (N_18950,N_18766,N_18759);
or U18951 (N_18951,N_18740,N_18867);
and U18952 (N_18952,N_18816,N_18738);
or U18953 (N_18953,N_18824,N_18839);
nand U18954 (N_18954,N_18752,N_18778);
or U18955 (N_18955,N_18723,N_18745);
or U18956 (N_18956,N_18722,N_18794);
nand U18957 (N_18957,N_18807,N_18842);
nor U18958 (N_18958,N_18730,N_18833);
or U18959 (N_18959,N_18764,N_18805);
nand U18960 (N_18960,N_18820,N_18868);
xor U18961 (N_18961,N_18850,N_18826);
nand U18962 (N_18962,N_18745,N_18767);
or U18963 (N_18963,N_18730,N_18793);
and U18964 (N_18964,N_18753,N_18869);
xnor U18965 (N_18965,N_18790,N_18758);
nand U18966 (N_18966,N_18738,N_18791);
xnor U18967 (N_18967,N_18860,N_18724);
and U18968 (N_18968,N_18790,N_18738);
nor U18969 (N_18969,N_18725,N_18776);
nor U18970 (N_18970,N_18839,N_18746);
and U18971 (N_18971,N_18812,N_18762);
and U18972 (N_18972,N_18873,N_18831);
nand U18973 (N_18973,N_18739,N_18844);
xor U18974 (N_18974,N_18867,N_18782);
and U18975 (N_18975,N_18747,N_18756);
xor U18976 (N_18976,N_18765,N_18841);
or U18977 (N_18977,N_18826,N_18746);
xor U18978 (N_18978,N_18804,N_18809);
nand U18979 (N_18979,N_18832,N_18726);
and U18980 (N_18980,N_18738,N_18733);
and U18981 (N_18981,N_18748,N_18877);
and U18982 (N_18982,N_18737,N_18874);
nand U18983 (N_18983,N_18843,N_18833);
and U18984 (N_18984,N_18778,N_18721);
xnor U18985 (N_18985,N_18726,N_18791);
and U18986 (N_18986,N_18720,N_18783);
or U18987 (N_18987,N_18787,N_18732);
or U18988 (N_18988,N_18807,N_18738);
and U18989 (N_18989,N_18820,N_18734);
nand U18990 (N_18990,N_18739,N_18878);
xor U18991 (N_18991,N_18863,N_18853);
nor U18992 (N_18992,N_18838,N_18875);
or U18993 (N_18993,N_18839,N_18869);
nand U18994 (N_18994,N_18858,N_18743);
and U18995 (N_18995,N_18840,N_18824);
nor U18996 (N_18996,N_18864,N_18791);
and U18997 (N_18997,N_18870,N_18802);
nand U18998 (N_18998,N_18818,N_18743);
and U18999 (N_18999,N_18855,N_18788);
xnor U19000 (N_19000,N_18765,N_18847);
xnor U19001 (N_19001,N_18818,N_18869);
or U19002 (N_19002,N_18733,N_18821);
or U19003 (N_19003,N_18783,N_18827);
nand U19004 (N_19004,N_18875,N_18853);
xnor U19005 (N_19005,N_18855,N_18801);
xnor U19006 (N_19006,N_18807,N_18778);
nor U19007 (N_19007,N_18803,N_18807);
or U19008 (N_19008,N_18733,N_18879);
nor U19009 (N_19009,N_18845,N_18798);
nor U19010 (N_19010,N_18727,N_18838);
or U19011 (N_19011,N_18796,N_18730);
or U19012 (N_19012,N_18813,N_18763);
or U19013 (N_19013,N_18769,N_18801);
and U19014 (N_19014,N_18853,N_18816);
xor U19015 (N_19015,N_18735,N_18753);
and U19016 (N_19016,N_18760,N_18818);
or U19017 (N_19017,N_18828,N_18783);
nor U19018 (N_19018,N_18840,N_18727);
xor U19019 (N_19019,N_18806,N_18762);
nor U19020 (N_19020,N_18732,N_18731);
xnor U19021 (N_19021,N_18844,N_18780);
nand U19022 (N_19022,N_18839,N_18868);
or U19023 (N_19023,N_18725,N_18808);
or U19024 (N_19024,N_18735,N_18794);
nor U19025 (N_19025,N_18824,N_18835);
xnor U19026 (N_19026,N_18822,N_18760);
or U19027 (N_19027,N_18844,N_18752);
nand U19028 (N_19028,N_18757,N_18808);
nand U19029 (N_19029,N_18843,N_18803);
xnor U19030 (N_19030,N_18871,N_18730);
nand U19031 (N_19031,N_18855,N_18854);
nand U19032 (N_19032,N_18861,N_18724);
nor U19033 (N_19033,N_18827,N_18838);
nand U19034 (N_19034,N_18856,N_18787);
or U19035 (N_19035,N_18735,N_18804);
and U19036 (N_19036,N_18865,N_18822);
nor U19037 (N_19037,N_18857,N_18802);
and U19038 (N_19038,N_18754,N_18877);
xnor U19039 (N_19039,N_18799,N_18730);
xnor U19040 (N_19040,N_19006,N_18958);
xor U19041 (N_19041,N_19031,N_18912);
nor U19042 (N_19042,N_18913,N_18995);
nor U19043 (N_19043,N_18927,N_18946);
and U19044 (N_19044,N_18979,N_19035);
xnor U19045 (N_19045,N_19033,N_18948);
nand U19046 (N_19046,N_18890,N_18998);
or U19047 (N_19047,N_18929,N_18955);
nand U19048 (N_19048,N_18915,N_19015);
and U19049 (N_19049,N_18885,N_19009);
nor U19050 (N_19050,N_18896,N_18956);
nand U19051 (N_19051,N_19030,N_18977);
xor U19052 (N_19052,N_18962,N_18938);
nor U19053 (N_19053,N_18924,N_19038);
xnor U19054 (N_19054,N_18901,N_18987);
and U19055 (N_19055,N_18966,N_19014);
nand U19056 (N_19056,N_18934,N_18908);
nor U19057 (N_19057,N_18897,N_18982);
xor U19058 (N_19058,N_18944,N_18953);
and U19059 (N_19059,N_18936,N_19007);
or U19060 (N_19060,N_18949,N_18968);
or U19061 (N_19061,N_18976,N_19019);
and U19062 (N_19062,N_18972,N_18952);
nand U19063 (N_19063,N_18898,N_18997);
or U19064 (N_19064,N_18895,N_18900);
or U19065 (N_19065,N_18907,N_18884);
nand U19066 (N_19066,N_18964,N_18894);
nand U19067 (N_19067,N_18926,N_19011);
and U19068 (N_19068,N_19002,N_18881);
and U19069 (N_19069,N_18910,N_18971);
or U19070 (N_19070,N_18947,N_18889);
or U19071 (N_19071,N_19025,N_18965);
xor U19072 (N_19072,N_19034,N_18880);
and U19073 (N_19073,N_18888,N_18957);
or U19074 (N_19074,N_18932,N_18960);
nand U19075 (N_19075,N_18967,N_18970);
nor U19076 (N_19076,N_18904,N_18975);
nand U19077 (N_19077,N_18903,N_19013);
xnor U19078 (N_19078,N_19022,N_18992);
nor U19079 (N_19079,N_19017,N_18939);
nand U19080 (N_19080,N_18981,N_19012);
xnor U19081 (N_19081,N_18996,N_18917);
or U19082 (N_19082,N_19021,N_18999);
or U19083 (N_19083,N_18921,N_19036);
or U19084 (N_19084,N_18920,N_18893);
xor U19085 (N_19085,N_18883,N_18933);
and U19086 (N_19086,N_18930,N_19010);
or U19087 (N_19087,N_18994,N_19000);
or U19088 (N_19088,N_18990,N_18961);
nand U19089 (N_19089,N_19001,N_19027);
nor U19090 (N_19090,N_18882,N_19039);
and U19091 (N_19091,N_18985,N_18941);
nor U19092 (N_19092,N_18902,N_19024);
xor U19093 (N_19093,N_18991,N_19018);
and U19094 (N_19094,N_18905,N_18969);
xnor U19095 (N_19095,N_18980,N_19028);
nor U19096 (N_19096,N_18886,N_19008);
or U19097 (N_19097,N_18931,N_18925);
nor U19098 (N_19098,N_18983,N_19029);
nor U19099 (N_19099,N_18945,N_19037);
nand U19100 (N_19100,N_18922,N_19016);
or U19101 (N_19101,N_18916,N_18937);
xnor U19102 (N_19102,N_18988,N_19026);
nor U19103 (N_19103,N_18918,N_18899);
xnor U19104 (N_19104,N_18963,N_18942);
nand U19105 (N_19105,N_18892,N_18974);
or U19106 (N_19106,N_19005,N_18935);
and U19107 (N_19107,N_18978,N_18943);
nand U19108 (N_19108,N_18887,N_18959);
and U19109 (N_19109,N_18906,N_18989);
and U19110 (N_19110,N_18950,N_18891);
nand U19111 (N_19111,N_19032,N_18986);
and U19112 (N_19112,N_18984,N_18909);
xor U19113 (N_19113,N_18928,N_18923);
and U19114 (N_19114,N_18973,N_18940);
or U19115 (N_19115,N_18993,N_19020);
nor U19116 (N_19116,N_18911,N_19004);
and U19117 (N_19117,N_18954,N_19023);
and U19118 (N_19118,N_18951,N_18919);
nand U19119 (N_19119,N_19003,N_18914);
nand U19120 (N_19120,N_18889,N_18961);
and U19121 (N_19121,N_18921,N_18887);
nor U19122 (N_19122,N_18887,N_18883);
xor U19123 (N_19123,N_18977,N_18905);
and U19124 (N_19124,N_18991,N_18947);
nor U19125 (N_19125,N_19023,N_18921);
nor U19126 (N_19126,N_19005,N_18926);
xor U19127 (N_19127,N_18905,N_18983);
and U19128 (N_19128,N_18915,N_18898);
nor U19129 (N_19129,N_19024,N_18907);
xor U19130 (N_19130,N_18964,N_19022);
nor U19131 (N_19131,N_18973,N_19037);
xor U19132 (N_19132,N_18908,N_18917);
and U19133 (N_19133,N_18898,N_18913);
nand U19134 (N_19134,N_18895,N_18896);
nand U19135 (N_19135,N_18903,N_19027);
nor U19136 (N_19136,N_18989,N_18943);
xor U19137 (N_19137,N_18940,N_18919);
xor U19138 (N_19138,N_19005,N_18905);
and U19139 (N_19139,N_18992,N_19020);
xnor U19140 (N_19140,N_18973,N_18884);
nor U19141 (N_19141,N_18950,N_18925);
and U19142 (N_19142,N_18880,N_19036);
nand U19143 (N_19143,N_18923,N_18995);
or U19144 (N_19144,N_19037,N_19035);
or U19145 (N_19145,N_18936,N_18967);
and U19146 (N_19146,N_18977,N_18880);
and U19147 (N_19147,N_18884,N_18970);
nor U19148 (N_19148,N_19017,N_19000);
or U19149 (N_19149,N_18903,N_18979);
nor U19150 (N_19150,N_18903,N_18904);
and U19151 (N_19151,N_18911,N_18883);
or U19152 (N_19152,N_18891,N_18915);
and U19153 (N_19153,N_18895,N_18898);
and U19154 (N_19154,N_18888,N_19003);
nor U19155 (N_19155,N_19015,N_19006);
nand U19156 (N_19156,N_18950,N_18977);
nor U19157 (N_19157,N_18935,N_18988);
and U19158 (N_19158,N_19012,N_18951);
xnor U19159 (N_19159,N_18888,N_18918);
nand U19160 (N_19160,N_19006,N_18884);
xnor U19161 (N_19161,N_18940,N_18916);
or U19162 (N_19162,N_18921,N_18903);
xnor U19163 (N_19163,N_18957,N_19016);
or U19164 (N_19164,N_19038,N_18935);
nor U19165 (N_19165,N_18957,N_18882);
xnor U19166 (N_19166,N_19039,N_18929);
or U19167 (N_19167,N_18888,N_18995);
xor U19168 (N_19168,N_18903,N_18984);
and U19169 (N_19169,N_18949,N_18950);
xnor U19170 (N_19170,N_18925,N_18990);
nand U19171 (N_19171,N_18909,N_18930);
nand U19172 (N_19172,N_18992,N_18896);
or U19173 (N_19173,N_18961,N_19016);
nor U19174 (N_19174,N_18972,N_18967);
and U19175 (N_19175,N_19007,N_18956);
and U19176 (N_19176,N_18924,N_18956);
or U19177 (N_19177,N_18976,N_19037);
nor U19178 (N_19178,N_18902,N_19015);
or U19179 (N_19179,N_19021,N_18957);
xor U19180 (N_19180,N_18951,N_18912);
xor U19181 (N_19181,N_18934,N_18897);
and U19182 (N_19182,N_18917,N_18960);
nand U19183 (N_19183,N_18936,N_18992);
and U19184 (N_19184,N_18882,N_18881);
nand U19185 (N_19185,N_18886,N_18880);
xor U19186 (N_19186,N_18882,N_18995);
or U19187 (N_19187,N_18996,N_18957);
nor U19188 (N_19188,N_18902,N_19021);
xnor U19189 (N_19189,N_18887,N_18927);
xnor U19190 (N_19190,N_18950,N_18892);
or U19191 (N_19191,N_18993,N_18905);
and U19192 (N_19192,N_18918,N_19005);
nand U19193 (N_19193,N_19004,N_18985);
nor U19194 (N_19194,N_18897,N_18977);
nor U19195 (N_19195,N_18923,N_19034);
nor U19196 (N_19196,N_18969,N_19016);
nand U19197 (N_19197,N_18980,N_18969);
xor U19198 (N_19198,N_18896,N_18978);
or U19199 (N_19199,N_18897,N_18962);
xor U19200 (N_19200,N_19082,N_19047);
xor U19201 (N_19201,N_19061,N_19076);
nor U19202 (N_19202,N_19132,N_19085);
and U19203 (N_19203,N_19097,N_19046);
xor U19204 (N_19204,N_19094,N_19051);
and U19205 (N_19205,N_19152,N_19118);
and U19206 (N_19206,N_19182,N_19058);
and U19207 (N_19207,N_19189,N_19149);
nand U19208 (N_19208,N_19069,N_19145);
and U19209 (N_19209,N_19141,N_19146);
nor U19210 (N_19210,N_19104,N_19126);
or U19211 (N_19211,N_19185,N_19183);
xor U19212 (N_19212,N_19155,N_19055);
nor U19213 (N_19213,N_19103,N_19199);
and U19214 (N_19214,N_19128,N_19043);
nor U19215 (N_19215,N_19044,N_19158);
or U19216 (N_19216,N_19073,N_19190);
xor U19217 (N_19217,N_19113,N_19045);
and U19218 (N_19218,N_19084,N_19102);
xnor U19219 (N_19219,N_19174,N_19101);
or U19220 (N_19220,N_19111,N_19096);
or U19221 (N_19221,N_19140,N_19063);
nor U19222 (N_19222,N_19186,N_19086);
or U19223 (N_19223,N_19064,N_19040);
nor U19224 (N_19224,N_19192,N_19106);
or U19225 (N_19225,N_19195,N_19121);
xnor U19226 (N_19226,N_19169,N_19144);
nand U19227 (N_19227,N_19188,N_19196);
or U19228 (N_19228,N_19135,N_19120);
and U19229 (N_19229,N_19116,N_19052);
and U19230 (N_19230,N_19062,N_19191);
nor U19231 (N_19231,N_19057,N_19095);
or U19232 (N_19232,N_19168,N_19110);
nand U19233 (N_19233,N_19175,N_19108);
nor U19234 (N_19234,N_19122,N_19056);
or U19235 (N_19235,N_19059,N_19161);
nor U19236 (N_19236,N_19176,N_19193);
xor U19237 (N_19237,N_19173,N_19180);
nor U19238 (N_19238,N_19139,N_19081);
xor U19239 (N_19239,N_19067,N_19156);
nand U19240 (N_19240,N_19171,N_19119);
or U19241 (N_19241,N_19071,N_19177);
nand U19242 (N_19242,N_19074,N_19127);
xnor U19243 (N_19243,N_19091,N_19166);
and U19244 (N_19244,N_19184,N_19080);
nand U19245 (N_19245,N_19100,N_19088);
nor U19246 (N_19246,N_19137,N_19083);
xor U19247 (N_19247,N_19197,N_19134);
or U19248 (N_19248,N_19065,N_19165);
nand U19249 (N_19249,N_19143,N_19089);
nand U19250 (N_19250,N_19170,N_19041);
nand U19251 (N_19251,N_19154,N_19099);
nor U19252 (N_19252,N_19187,N_19160);
or U19253 (N_19253,N_19092,N_19167);
or U19254 (N_19254,N_19053,N_19163);
xnor U19255 (N_19255,N_19079,N_19194);
or U19256 (N_19256,N_19157,N_19164);
xor U19257 (N_19257,N_19131,N_19151);
nor U19258 (N_19258,N_19142,N_19130);
nand U19259 (N_19259,N_19124,N_19112);
nor U19260 (N_19260,N_19133,N_19117);
and U19261 (N_19261,N_19107,N_19198);
nand U19262 (N_19262,N_19123,N_19105);
and U19263 (N_19263,N_19098,N_19075);
nand U19264 (N_19264,N_19054,N_19050);
xnor U19265 (N_19265,N_19162,N_19159);
nor U19266 (N_19266,N_19066,N_19136);
nand U19267 (N_19267,N_19093,N_19179);
xnor U19268 (N_19268,N_19087,N_19115);
nand U19269 (N_19269,N_19125,N_19077);
nand U19270 (N_19270,N_19072,N_19147);
or U19271 (N_19271,N_19138,N_19070);
nand U19272 (N_19272,N_19048,N_19181);
nand U19273 (N_19273,N_19150,N_19042);
and U19274 (N_19274,N_19172,N_19148);
nand U19275 (N_19275,N_19060,N_19178);
and U19276 (N_19276,N_19114,N_19090);
nor U19277 (N_19277,N_19068,N_19153);
nor U19278 (N_19278,N_19129,N_19078);
nand U19279 (N_19279,N_19049,N_19109);
and U19280 (N_19280,N_19135,N_19187);
or U19281 (N_19281,N_19083,N_19198);
and U19282 (N_19282,N_19159,N_19180);
xnor U19283 (N_19283,N_19142,N_19050);
and U19284 (N_19284,N_19194,N_19195);
nand U19285 (N_19285,N_19059,N_19074);
xor U19286 (N_19286,N_19161,N_19102);
or U19287 (N_19287,N_19190,N_19055);
nand U19288 (N_19288,N_19132,N_19143);
or U19289 (N_19289,N_19180,N_19155);
nor U19290 (N_19290,N_19185,N_19184);
nor U19291 (N_19291,N_19168,N_19047);
or U19292 (N_19292,N_19084,N_19116);
xnor U19293 (N_19293,N_19100,N_19181);
nand U19294 (N_19294,N_19131,N_19164);
nand U19295 (N_19295,N_19156,N_19108);
xor U19296 (N_19296,N_19101,N_19103);
nor U19297 (N_19297,N_19145,N_19093);
and U19298 (N_19298,N_19183,N_19148);
xor U19299 (N_19299,N_19171,N_19132);
xnor U19300 (N_19300,N_19114,N_19116);
or U19301 (N_19301,N_19171,N_19096);
nand U19302 (N_19302,N_19077,N_19120);
nor U19303 (N_19303,N_19108,N_19094);
nand U19304 (N_19304,N_19159,N_19052);
and U19305 (N_19305,N_19161,N_19184);
xnor U19306 (N_19306,N_19084,N_19082);
or U19307 (N_19307,N_19103,N_19167);
nor U19308 (N_19308,N_19139,N_19100);
xor U19309 (N_19309,N_19132,N_19141);
or U19310 (N_19310,N_19137,N_19198);
nor U19311 (N_19311,N_19102,N_19186);
nand U19312 (N_19312,N_19110,N_19139);
and U19313 (N_19313,N_19133,N_19085);
xor U19314 (N_19314,N_19042,N_19142);
nor U19315 (N_19315,N_19173,N_19158);
nand U19316 (N_19316,N_19125,N_19050);
nand U19317 (N_19317,N_19147,N_19119);
nor U19318 (N_19318,N_19149,N_19171);
xnor U19319 (N_19319,N_19082,N_19119);
xnor U19320 (N_19320,N_19159,N_19071);
nand U19321 (N_19321,N_19157,N_19192);
or U19322 (N_19322,N_19150,N_19079);
or U19323 (N_19323,N_19196,N_19130);
nor U19324 (N_19324,N_19153,N_19059);
nand U19325 (N_19325,N_19127,N_19079);
nor U19326 (N_19326,N_19189,N_19089);
and U19327 (N_19327,N_19050,N_19176);
xor U19328 (N_19328,N_19117,N_19151);
nor U19329 (N_19329,N_19187,N_19108);
xor U19330 (N_19330,N_19137,N_19055);
nor U19331 (N_19331,N_19139,N_19167);
nand U19332 (N_19332,N_19126,N_19175);
or U19333 (N_19333,N_19138,N_19158);
nand U19334 (N_19334,N_19122,N_19041);
xor U19335 (N_19335,N_19135,N_19116);
xnor U19336 (N_19336,N_19051,N_19077);
or U19337 (N_19337,N_19153,N_19128);
or U19338 (N_19338,N_19193,N_19064);
nand U19339 (N_19339,N_19085,N_19041);
nor U19340 (N_19340,N_19097,N_19168);
and U19341 (N_19341,N_19163,N_19125);
nand U19342 (N_19342,N_19168,N_19101);
and U19343 (N_19343,N_19091,N_19078);
xnor U19344 (N_19344,N_19141,N_19114);
xnor U19345 (N_19345,N_19148,N_19089);
and U19346 (N_19346,N_19153,N_19114);
xor U19347 (N_19347,N_19156,N_19197);
nand U19348 (N_19348,N_19194,N_19127);
nand U19349 (N_19349,N_19063,N_19197);
or U19350 (N_19350,N_19062,N_19184);
or U19351 (N_19351,N_19124,N_19151);
and U19352 (N_19352,N_19103,N_19108);
or U19353 (N_19353,N_19107,N_19185);
and U19354 (N_19354,N_19070,N_19185);
and U19355 (N_19355,N_19170,N_19131);
or U19356 (N_19356,N_19159,N_19041);
nor U19357 (N_19357,N_19063,N_19093);
xnor U19358 (N_19358,N_19091,N_19060);
nor U19359 (N_19359,N_19184,N_19195);
or U19360 (N_19360,N_19225,N_19227);
nand U19361 (N_19361,N_19204,N_19348);
or U19362 (N_19362,N_19301,N_19286);
nor U19363 (N_19363,N_19288,N_19250);
nand U19364 (N_19364,N_19340,N_19215);
or U19365 (N_19365,N_19245,N_19350);
nor U19366 (N_19366,N_19216,N_19352);
nand U19367 (N_19367,N_19234,N_19224);
nor U19368 (N_19368,N_19321,N_19326);
nor U19369 (N_19369,N_19243,N_19306);
nand U19370 (N_19370,N_19318,N_19231);
or U19371 (N_19371,N_19226,N_19331);
nand U19372 (N_19372,N_19287,N_19341);
or U19373 (N_19373,N_19240,N_19358);
nand U19374 (N_19374,N_19222,N_19237);
and U19375 (N_19375,N_19357,N_19229);
and U19376 (N_19376,N_19281,N_19300);
xor U19377 (N_19377,N_19228,N_19349);
and U19378 (N_19378,N_19263,N_19283);
and U19379 (N_19379,N_19309,N_19218);
nor U19380 (N_19380,N_19328,N_19285);
xnor U19381 (N_19381,N_19353,N_19271);
nor U19382 (N_19382,N_19217,N_19330);
nand U19383 (N_19383,N_19256,N_19339);
and U19384 (N_19384,N_19268,N_19261);
nand U19385 (N_19385,N_19290,N_19275);
nor U19386 (N_19386,N_19282,N_19253);
nand U19387 (N_19387,N_19270,N_19292);
nand U19388 (N_19388,N_19254,N_19344);
nor U19389 (N_19389,N_19205,N_19316);
nor U19390 (N_19390,N_19265,N_19345);
nor U19391 (N_19391,N_19221,N_19251);
and U19392 (N_19392,N_19320,N_19333);
and U19393 (N_19393,N_19332,N_19299);
and U19394 (N_19394,N_19201,N_19249);
nand U19395 (N_19395,N_19279,N_19272);
nor U19396 (N_19396,N_19317,N_19312);
or U19397 (N_19397,N_19220,N_19308);
xor U19398 (N_19398,N_19329,N_19230);
and U19399 (N_19399,N_19296,N_19239);
nor U19400 (N_19400,N_19310,N_19209);
xnor U19401 (N_19401,N_19325,N_19212);
xor U19402 (N_19402,N_19307,N_19207);
and U19403 (N_19403,N_19257,N_19322);
and U19404 (N_19404,N_19338,N_19232);
nand U19405 (N_19405,N_19200,N_19346);
and U19406 (N_19406,N_19244,N_19314);
nand U19407 (N_19407,N_19323,N_19276);
nor U19408 (N_19408,N_19211,N_19273);
xnor U19409 (N_19409,N_19327,N_19302);
nand U19410 (N_19410,N_19235,N_19334);
and U19411 (N_19411,N_19303,N_19247);
or U19412 (N_19412,N_19294,N_19233);
nand U19413 (N_19413,N_19266,N_19258);
nor U19414 (N_19414,N_19248,N_19238);
nor U19415 (N_19415,N_19336,N_19219);
nor U19416 (N_19416,N_19298,N_19210);
nor U19417 (N_19417,N_19259,N_19241);
and U19418 (N_19418,N_19252,N_19354);
or U19419 (N_19419,N_19236,N_19342);
nand U19420 (N_19420,N_19206,N_19324);
xnor U19421 (N_19421,N_19214,N_19295);
nand U19422 (N_19422,N_19269,N_19319);
or U19423 (N_19423,N_19311,N_19260);
and U19424 (N_19424,N_19335,N_19355);
xor U19425 (N_19425,N_19337,N_19246);
xor U19426 (N_19426,N_19262,N_19315);
and U19427 (N_19427,N_19242,N_19297);
or U19428 (N_19428,N_19278,N_19213);
nand U19429 (N_19429,N_19223,N_19277);
nand U19430 (N_19430,N_19291,N_19343);
and U19431 (N_19431,N_19267,N_19305);
xor U19432 (N_19432,N_19293,N_19203);
nand U19433 (N_19433,N_19255,N_19274);
nor U19434 (N_19434,N_19351,N_19284);
or U19435 (N_19435,N_19280,N_19347);
nand U19436 (N_19436,N_19289,N_19356);
and U19437 (N_19437,N_19359,N_19313);
nand U19438 (N_19438,N_19304,N_19202);
and U19439 (N_19439,N_19264,N_19208);
xor U19440 (N_19440,N_19208,N_19224);
nand U19441 (N_19441,N_19287,N_19356);
or U19442 (N_19442,N_19312,N_19313);
and U19443 (N_19443,N_19320,N_19303);
nor U19444 (N_19444,N_19274,N_19219);
and U19445 (N_19445,N_19269,N_19265);
nand U19446 (N_19446,N_19277,N_19252);
xor U19447 (N_19447,N_19287,N_19353);
nand U19448 (N_19448,N_19332,N_19317);
and U19449 (N_19449,N_19333,N_19321);
nor U19450 (N_19450,N_19352,N_19269);
xnor U19451 (N_19451,N_19263,N_19222);
nand U19452 (N_19452,N_19265,N_19240);
and U19453 (N_19453,N_19201,N_19246);
nand U19454 (N_19454,N_19305,N_19358);
xnor U19455 (N_19455,N_19334,N_19305);
and U19456 (N_19456,N_19352,N_19203);
nand U19457 (N_19457,N_19277,N_19321);
xnor U19458 (N_19458,N_19320,N_19353);
nor U19459 (N_19459,N_19201,N_19261);
xnor U19460 (N_19460,N_19272,N_19258);
and U19461 (N_19461,N_19203,N_19202);
nor U19462 (N_19462,N_19233,N_19308);
nor U19463 (N_19463,N_19237,N_19320);
xnor U19464 (N_19464,N_19271,N_19307);
nand U19465 (N_19465,N_19339,N_19243);
xor U19466 (N_19466,N_19213,N_19344);
nor U19467 (N_19467,N_19316,N_19324);
nand U19468 (N_19468,N_19315,N_19355);
xor U19469 (N_19469,N_19296,N_19245);
and U19470 (N_19470,N_19350,N_19289);
and U19471 (N_19471,N_19268,N_19283);
or U19472 (N_19472,N_19212,N_19254);
and U19473 (N_19473,N_19268,N_19234);
nand U19474 (N_19474,N_19323,N_19309);
and U19475 (N_19475,N_19283,N_19315);
or U19476 (N_19476,N_19276,N_19298);
xor U19477 (N_19477,N_19260,N_19239);
nor U19478 (N_19478,N_19300,N_19257);
nand U19479 (N_19479,N_19253,N_19338);
or U19480 (N_19480,N_19255,N_19251);
or U19481 (N_19481,N_19328,N_19356);
or U19482 (N_19482,N_19207,N_19239);
nor U19483 (N_19483,N_19288,N_19319);
nand U19484 (N_19484,N_19276,N_19271);
xnor U19485 (N_19485,N_19304,N_19208);
nor U19486 (N_19486,N_19301,N_19277);
xnor U19487 (N_19487,N_19280,N_19262);
xor U19488 (N_19488,N_19213,N_19323);
xor U19489 (N_19489,N_19297,N_19207);
xor U19490 (N_19490,N_19251,N_19280);
and U19491 (N_19491,N_19290,N_19354);
and U19492 (N_19492,N_19207,N_19281);
or U19493 (N_19493,N_19206,N_19333);
or U19494 (N_19494,N_19241,N_19233);
or U19495 (N_19495,N_19341,N_19339);
and U19496 (N_19496,N_19235,N_19271);
nand U19497 (N_19497,N_19330,N_19346);
nand U19498 (N_19498,N_19218,N_19296);
xor U19499 (N_19499,N_19277,N_19259);
or U19500 (N_19500,N_19214,N_19243);
and U19501 (N_19501,N_19309,N_19341);
nand U19502 (N_19502,N_19282,N_19271);
or U19503 (N_19503,N_19224,N_19209);
and U19504 (N_19504,N_19259,N_19220);
nand U19505 (N_19505,N_19247,N_19350);
nand U19506 (N_19506,N_19304,N_19327);
xor U19507 (N_19507,N_19284,N_19357);
xor U19508 (N_19508,N_19319,N_19314);
nand U19509 (N_19509,N_19331,N_19265);
and U19510 (N_19510,N_19220,N_19326);
and U19511 (N_19511,N_19274,N_19333);
or U19512 (N_19512,N_19294,N_19310);
and U19513 (N_19513,N_19358,N_19303);
nand U19514 (N_19514,N_19279,N_19300);
xor U19515 (N_19515,N_19212,N_19348);
and U19516 (N_19516,N_19316,N_19215);
or U19517 (N_19517,N_19317,N_19269);
nand U19518 (N_19518,N_19280,N_19316);
xor U19519 (N_19519,N_19249,N_19245);
and U19520 (N_19520,N_19369,N_19383);
and U19521 (N_19521,N_19463,N_19413);
and U19522 (N_19522,N_19434,N_19468);
nand U19523 (N_19523,N_19412,N_19508);
and U19524 (N_19524,N_19481,N_19392);
nand U19525 (N_19525,N_19371,N_19389);
nor U19526 (N_19526,N_19424,N_19406);
xnor U19527 (N_19527,N_19401,N_19414);
and U19528 (N_19528,N_19466,N_19375);
xnor U19529 (N_19529,N_19495,N_19421);
nand U19530 (N_19530,N_19436,N_19433);
nor U19531 (N_19531,N_19446,N_19454);
nand U19532 (N_19532,N_19470,N_19395);
xor U19533 (N_19533,N_19367,N_19407);
nand U19534 (N_19534,N_19469,N_19409);
nor U19535 (N_19535,N_19438,N_19388);
nand U19536 (N_19536,N_19377,N_19426);
xor U19537 (N_19537,N_19465,N_19439);
nand U19538 (N_19538,N_19486,N_19425);
and U19539 (N_19539,N_19471,N_19394);
xor U19540 (N_19540,N_19361,N_19366);
nor U19541 (N_19541,N_19501,N_19497);
and U19542 (N_19542,N_19511,N_19418);
and U19543 (N_19543,N_19419,N_19429);
nor U19544 (N_19544,N_19444,N_19376);
xnor U19545 (N_19545,N_19518,N_19507);
nor U19546 (N_19546,N_19374,N_19442);
xnor U19547 (N_19547,N_19513,N_19482);
nor U19548 (N_19548,N_19472,N_19493);
or U19549 (N_19549,N_19516,N_19475);
xor U19550 (N_19550,N_19423,N_19467);
nand U19551 (N_19551,N_19473,N_19391);
nor U19552 (N_19552,N_19519,N_19386);
xor U19553 (N_19553,N_19450,N_19385);
nor U19554 (N_19554,N_19447,N_19431);
nor U19555 (N_19555,N_19477,N_19448);
xor U19556 (N_19556,N_19500,N_19373);
nand U19557 (N_19557,N_19363,N_19362);
and U19558 (N_19558,N_19505,N_19499);
nor U19559 (N_19559,N_19494,N_19437);
and U19560 (N_19560,N_19420,N_19422);
or U19561 (N_19561,N_19474,N_19380);
nand U19562 (N_19562,N_19498,N_19379);
or U19563 (N_19563,N_19453,N_19514);
and U19564 (N_19564,N_19489,N_19504);
or U19565 (N_19565,N_19459,N_19397);
nor U19566 (N_19566,N_19410,N_19440);
xor U19567 (N_19567,N_19456,N_19443);
nor U19568 (N_19568,N_19502,N_19488);
and U19569 (N_19569,N_19462,N_19485);
and U19570 (N_19570,N_19452,N_19512);
nand U19571 (N_19571,N_19387,N_19372);
nor U19572 (N_19572,N_19364,N_19393);
xnor U19573 (N_19573,N_19390,N_19396);
and U19574 (N_19574,N_19496,N_19378);
and U19575 (N_19575,N_19487,N_19399);
xnor U19576 (N_19576,N_19509,N_19403);
xnor U19577 (N_19577,N_19365,N_19411);
xor U19578 (N_19578,N_19480,N_19515);
or U19579 (N_19579,N_19416,N_19455);
nor U19580 (N_19580,N_19506,N_19400);
and U19581 (N_19581,N_19460,N_19432);
nand U19582 (N_19582,N_19478,N_19398);
and U19583 (N_19583,N_19492,N_19368);
nand U19584 (N_19584,N_19427,N_19503);
nand U19585 (N_19585,N_19381,N_19449);
or U19586 (N_19586,N_19405,N_19417);
xnor U19587 (N_19587,N_19464,N_19461);
and U19588 (N_19588,N_19360,N_19445);
or U19589 (N_19589,N_19510,N_19451);
nand U19590 (N_19590,N_19435,N_19457);
and U19591 (N_19591,N_19402,N_19370);
nor U19592 (N_19592,N_19384,N_19428);
or U19593 (N_19593,N_19484,N_19430);
and U19594 (N_19594,N_19491,N_19458);
nand U19595 (N_19595,N_19483,N_19408);
or U19596 (N_19596,N_19490,N_19476);
nand U19597 (N_19597,N_19404,N_19415);
or U19598 (N_19598,N_19517,N_19441);
or U19599 (N_19599,N_19382,N_19479);
or U19600 (N_19600,N_19427,N_19380);
xor U19601 (N_19601,N_19517,N_19380);
nor U19602 (N_19602,N_19484,N_19479);
or U19603 (N_19603,N_19407,N_19366);
or U19604 (N_19604,N_19425,N_19476);
and U19605 (N_19605,N_19473,N_19373);
nor U19606 (N_19606,N_19360,N_19481);
nand U19607 (N_19607,N_19456,N_19411);
and U19608 (N_19608,N_19507,N_19490);
nor U19609 (N_19609,N_19478,N_19457);
nand U19610 (N_19610,N_19424,N_19384);
nand U19611 (N_19611,N_19465,N_19518);
nand U19612 (N_19612,N_19421,N_19453);
nor U19613 (N_19613,N_19447,N_19444);
and U19614 (N_19614,N_19412,N_19380);
or U19615 (N_19615,N_19513,N_19410);
nor U19616 (N_19616,N_19452,N_19369);
or U19617 (N_19617,N_19381,N_19462);
or U19618 (N_19618,N_19496,N_19504);
nand U19619 (N_19619,N_19492,N_19441);
and U19620 (N_19620,N_19380,N_19415);
nand U19621 (N_19621,N_19479,N_19488);
nor U19622 (N_19622,N_19403,N_19446);
and U19623 (N_19623,N_19458,N_19428);
and U19624 (N_19624,N_19510,N_19485);
xnor U19625 (N_19625,N_19413,N_19506);
nor U19626 (N_19626,N_19492,N_19455);
nand U19627 (N_19627,N_19451,N_19423);
nand U19628 (N_19628,N_19470,N_19415);
nand U19629 (N_19629,N_19383,N_19444);
nor U19630 (N_19630,N_19427,N_19423);
or U19631 (N_19631,N_19420,N_19449);
or U19632 (N_19632,N_19508,N_19512);
nand U19633 (N_19633,N_19432,N_19470);
nand U19634 (N_19634,N_19367,N_19472);
xor U19635 (N_19635,N_19496,N_19467);
nor U19636 (N_19636,N_19510,N_19417);
nor U19637 (N_19637,N_19513,N_19510);
nor U19638 (N_19638,N_19493,N_19363);
and U19639 (N_19639,N_19494,N_19434);
nand U19640 (N_19640,N_19511,N_19420);
xor U19641 (N_19641,N_19399,N_19492);
or U19642 (N_19642,N_19412,N_19503);
and U19643 (N_19643,N_19427,N_19452);
or U19644 (N_19644,N_19466,N_19454);
nand U19645 (N_19645,N_19413,N_19411);
nand U19646 (N_19646,N_19473,N_19507);
nand U19647 (N_19647,N_19433,N_19476);
nand U19648 (N_19648,N_19519,N_19411);
nand U19649 (N_19649,N_19438,N_19471);
xnor U19650 (N_19650,N_19498,N_19429);
xnor U19651 (N_19651,N_19421,N_19365);
nand U19652 (N_19652,N_19509,N_19382);
nor U19653 (N_19653,N_19458,N_19384);
nor U19654 (N_19654,N_19437,N_19364);
and U19655 (N_19655,N_19494,N_19495);
and U19656 (N_19656,N_19376,N_19405);
or U19657 (N_19657,N_19400,N_19367);
and U19658 (N_19658,N_19365,N_19415);
nand U19659 (N_19659,N_19489,N_19438);
and U19660 (N_19660,N_19385,N_19468);
and U19661 (N_19661,N_19386,N_19469);
xor U19662 (N_19662,N_19401,N_19393);
nand U19663 (N_19663,N_19454,N_19391);
or U19664 (N_19664,N_19453,N_19488);
nand U19665 (N_19665,N_19368,N_19476);
nor U19666 (N_19666,N_19442,N_19452);
or U19667 (N_19667,N_19386,N_19466);
xor U19668 (N_19668,N_19459,N_19467);
nand U19669 (N_19669,N_19476,N_19386);
nor U19670 (N_19670,N_19476,N_19370);
or U19671 (N_19671,N_19491,N_19376);
xor U19672 (N_19672,N_19364,N_19421);
nand U19673 (N_19673,N_19513,N_19485);
and U19674 (N_19674,N_19493,N_19476);
nand U19675 (N_19675,N_19414,N_19459);
or U19676 (N_19676,N_19476,N_19508);
and U19677 (N_19677,N_19439,N_19512);
nor U19678 (N_19678,N_19402,N_19407);
and U19679 (N_19679,N_19395,N_19404);
or U19680 (N_19680,N_19593,N_19650);
nor U19681 (N_19681,N_19581,N_19521);
and U19682 (N_19682,N_19621,N_19605);
xor U19683 (N_19683,N_19638,N_19631);
nor U19684 (N_19684,N_19634,N_19527);
or U19685 (N_19685,N_19660,N_19556);
nor U19686 (N_19686,N_19586,N_19564);
xor U19687 (N_19687,N_19574,N_19542);
nand U19688 (N_19688,N_19657,N_19659);
xnor U19689 (N_19689,N_19569,N_19588);
or U19690 (N_19690,N_19627,N_19545);
or U19691 (N_19691,N_19549,N_19644);
or U19692 (N_19692,N_19664,N_19550);
nor U19693 (N_19693,N_19568,N_19672);
and U19694 (N_19694,N_19599,N_19679);
nor U19695 (N_19695,N_19646,N_19607);
or U19696 (N_19696,N_19663,N_19630);
nand U19697 (N_19697,N_19575,N_19579);
xnor U19698 (N_19698,N_19539,N_19558);
or U19699 (N_19699,N_19554,N_19666);
nand U19700 (N_19700,N_19618,N_19661);
and U19701 (N_19701,N_19538,N_19534);
or U19702 (N_19702,N_19662,N_19598);
and U19703 (N_19703,N_19647,N_19655);
or U19704 (N_19704,N_19637,N_19589);
nand U19705 (N_19705,N_19559,N_19604);
and U19706 (N_19706,N_19602,N_19674);
nand U19707 (N_19707,N_19530,N_19626);
or U19708 (N_19708,N_19528,N_19535);
nand U19709 (N_19709,N_19651,N_19582);
and U19710 (N_19710,N_19536,N_19597);
nand U19711 (N_19711,N_19533,N_19677);
nor U19712 (N_19712,N_19566,N_19654);
and U19713 (N_19713,N_19537,N_19547);
xnor U19714 (N_19714,N_19667,N_19642);
nand U19715 (N_19715,N_19543,N_19608);
xnor U19716 (N_19716,N_19625,N_19531);
nor U19717 (N_19717,N_19572,N_19671);
nor U19718 (N_19718,N_19524,N_19544);
xor U19719 (N_19719,N_19656,N_19552);
nand U19720 (N_19720,N_19557,N_19636);
and U19721 (N_19721,N_19600,N_19648);
and U19722 (N_19722,N_19573,N_19583);
xnor U19723 (N_19723,N_19567,N_19675);
or U19724 (N_19724,N_19609,N_19639);
and U19725 (N_19725,N_19617,N_19529);
xor U19726 (N_19726,N_19526,N_19540);
xnor U19727 (N_19727,N_19670,N_19629);
xnor U19728 (N_19728,N_19596,N_19610);
xor U19729 (N_19729,N_19635,N_19590);
or U19730 (N_19730,N_19669,N_19623);
and U19731 (N_19731,N_19525,N_19548);
nor U19732 (N_19732,N_19652,N_19673);
or U19733 (N_19733,N_19649,N_19668);
and U19734 (N_19734,N_19603,N_19601);
nor U19735 (N_19735,N_19522,N_19594);
nor U19736 (N_19736,N_19587,N_19615);
nand U19737 (N_19737,N_19632,N_19640);
nor U19738 (N_19738,N_19613,N_19624);
and U19739 (N_19739,N_19584,N_19611);
nand U19740 (N_19740,N_19585,N_19551);
nand U19741 (N_19741,N_19565,N_19678);
or U19742 (N_19742,N_19658,N_19580);
xnor U19743 (N_19743,N_19641,N_19643);
and U19744 (N_19744,N_19592,N_19619);
or U19745 (N_19745,N_19532,N_19628);
nand U19746 (N_19746,N_19665,N_19541);
and U19747 (N_19747,N_19616,N_19676);
nand U19748 (N_19748,N_19591,N_19562);
nor U19749 (N_19749,N_19614,N_19523);
and U19750 (N_19750,N_19520,N_19633);
xnor U19751 (N_19751,N_19578,N_19555);
or U19752 (N_19752,N_19577,N_19606);
nand U19753 (N_19753,N_19553,N_19570);
nand U19754 (N_19754,N_19653,N_19622);
nand U19755 (N_19755,N_19620,N_19560);
nand U19756 (N_19756,N_19612,N_19595);
or U19757 (N_19757,N_19576,N_19571);
nand U19758 (N_19758,N_19546,N_19561);
or U19759 (N_19759,N_19645,N_19563);
and U19760 (N_19760,N_19606,N_19618);
nand U19761 (N_19761,N_19543,N_19532);
nand U19762 (N_19762,N_19658,N_19566);
xor U19763 (N_19763,N_19666,N_19637);
or U19764 (N_19764,N_19578,N_19585);
or U19765 (N_19765,N_19563,N_19551);
nand U19766 (N_19766,N_19537,N_19600);
nor U19767 (N_19767,N_19652,N_19603);
and U19768 (N_19768,N_19615,N_19613);
and U19769 (N_19769,N_19554,N_19664);
or U19770 (N_19770,N_19603,N_19629);
or U19771 (N_19771,N_19658,N_19595);
xor U19772 (N_19772,N_19639,N_19539);
nand U19773 (N_19773,N_19616,N_19619);
and U19774 (N_19774,N_19583,N_19616);
nor U19775 (N_19775,N_19662,N_19605);
xor U19776 (N_19776,N_19611,N_19524);
xor U19777 (N_19777,N_19611,N_19539);
or U19778 (N_19778,N_19674,N_19658);
or U19779 (N_19779,N_19520,N_19610);
xnor U19780 (N_19780,N_19525,N_19598);
or U19781 (N_19781,N_19568,N_19533);
nand U19782 (N_19782,N_19561,N_19648);
or U19783 (N_19783,N_19634,N_19651);
or U19784 (N_19784,N_19578,N_19536);
xor U19785 (N_19785,N_19669,N_19530);
nor U19786 (N_19786,N_19667,N_19578);
or U19787 (N_19787,N_19589,N_19669);
nand U19788 (N_19788,N_19604,N_19523);
and U19789 (N_19789,N_19611,N_19652);
xnor U19790 (N_19790,N_19650,N_19522);
xnor U19791 (N_19791,N_19609,N_19543);
xnor U19792 (N_19792,N_19597,N_19558);
or U19793 (N_19793,N_19527,N_19617);
nand U19794 (N_19794,N_19630,N_19652);
or U19795 (N_19795,N_19558,N_19625);
or U19796 (N_19796,N_19585,N_19649);
and U19797 (N_19797,N_19624,N_19657);
xnor U19798 (N_19798,N_19661,N_19636);
nor U19799 (N_19799,N_19577,N_19537);
and U19800 (N_19800,N_19612,N_19523);
nand U19801 (N_19801,N_19524,N_19533);
nand U19802 (N_19802,N_19653,N_19581);
or U19803 (N_19803,N_19570,N_19670);
or U19804 (N_19804,N_19605,N_19587);
xnor U19805 (N_19805,N_19637,N_19602);
nor U19806 (N_19806,N_19615,N_19536);
nand U19807 (N_19807,N_19592,N_19530);
nor U19808 (N_19808,N_19642,N_19652);
and U19809 (N_19809,N_19587,N_19574);
or U19810 (N_19810,N_19552,N_19660);
and U19811 (N_19811,N_19654,N_19648);
xor U19812 (N_19812,N_19585,N_19615);
nand U19813 (N_19813,N_19610,N_19657);
or U19814 (N_19814,N_19576,N_19625);
nand U19815 (N_19815,N_19603,N_19615);
nor U19816 (N_19816,N_19542,N_19587);
xnor U19817 (N_19817,N_19618,N_19627);
xnor U19818 (N_19818,N_19625,N_19632);
xor U19819 (N_19819,N_19650,N_19540);
or U19820 (N_19820,N_19599,N_19538);
xnor U19821 (N_19821,N_19650,N_19609);
nor U19822 (N_19822,N_19641,N_19675);
nor U19823 (N_19823,N_19526,N_19594);
nor U19824 (N_19824,N_19648,N_19639);
or U19825 (N_19825,N_19647,N_19635);
nand U19826 (N_19826,N_19539,N_19620);
or U19827 (N_19827,N_19609,N_19619);
and U19828 (N_19828,N_19561,N_19622);
xor U19829 (N_19829,N_19557,N_19576);
nand U19830 (N_19830,N_19530,N_19646);
nand U19831 (N_19831,N_19627,N_19648);
xor U19832 (N_19832,N_19540,N_19536);
and U19833 (N_19833,N_19661,N_19521);
xnor U19834 (N_19834,N_19611,N_19535);
nand U19835 (N_19835,N_19673,N_19553);
and U19836 (N_19836,N_19551,N_19672);
or U19837 (N_19837,N_19659,N_19565);
or U19838 (N_19838,N_19558,N_19575);
xnor U19839 (N_19839,N_19618,N_19590);
xnor U19840 (N_19840,N_19816,N_19700);
nand U19841 (N_19841,N_19718,N_19835);
nor U19842 (N_19842,N_19712,N_19733);
nor U19843 (N_19843,N_19826,N_19773);
or U19844 (N_19844,N_19754,N_19704);
and U19845 (N_19845,N_19734,N_19731);
or U19846 (N_19846,N_19811,N_19694);
xnor U19847 (N_19847,N_19832,N_19805);
nand U19848 (N_19848,N_19744,N_19772);
nand U19849 (N_19849,N_19807,N_19748);
nor U19850 (N_19850,N_19758,N_19793);
xor U19851 (N_19851,N_19692,N_19720);
and U19852 (N_19852,N_19695,N_19818);
or U19853 (N_19853,N_19723,N_19741);
nor U19854 (N_19854,N_19781,N_19710);
and U19855 (N_19855,N_19770,N_19735);
nand U19856 (N_19856,N_19795,N_19697);
xnor U19857 (N_19857,N_19813,N_19761);
nand U19858 (N_19858,N_19787,N_19764);
or U19859 (N_19859,N_19681,N_19698);
xor U19860 (N_19860,N_19750,N_19738);
nor U19861 (N_19861,N_19782,N_19831);
or U19862 (N_19862,N_19737,N_19736);
nand U19863 (N_19863,N_19684,N_19766);
xnor U19864 (N_19864,N_19828,N_19707);
nor U19865 (N_19865,N_19716,N_19685);
or U19866 (N_19866,N_19804,N_19699);
nand U19867 (N_19867,N_19834,N_19774);
and U19868 (N_19868,N_19709,N_19839);
nand U19869 (N_19869,N_19812,N_19719);
nor U19870 (N_19870,N_19760,N_19686);
or U19871 (N_19871,N_19703,N_19799);
nand U19872 (N_19872,N_19753,N_19696);
and U19873 (N_19873,N_19775,N_19759);
nor U19874 (N_19874,N_19808,N_19780);
nor U19875 (N_19875,N_19825,N_19743);
or U19876 (N_19876,N_19767,N_19765);
or U19877 (N_19877,N_19814,N_19838);
nand U19878 (N_19878,N_19728,N_19803);
xor U19879 (N_19879,N_19745,N_19796);
nor U19880 (N_19880,N_19791,N_19730);
nand U19881 (N_19881,N_19794,N_19806);
xor U19882 (N_19882,N_19827,N_19815);
xnor U19883 (N_19883,N_19769,N_19800);
xnor U19884 (N_19884,N_19726,N_19749);
xor U19885 (N_19885,N_19727,N_19790);
nand U19886 (N_19886,N_19763,N_19777);
and U19887 (N_19887,N_19705,N_19789);
or U19888 (N_19888,N_19756,N_19746);
nand U19889 (N_19889,N_19801,N_19690);
and U19890 (N_19890,N_19768,N_19689);
xnor U19891 (N_19891,N_19740,N_19823);
or U19892 (N_19892,N_19691,N_19797);
xnor U19893 (N_19893,N_19798,N_19810);
and U19894 (N_19894,N_19817,N_19792);
and U19895 (N_19895,N_19739,N_19820);
xnor U19896 (N_19896,N_19715,N_19722);
and U19897 (N_19897,N_19802,N_19701);
or U19898 (N_19898,N_19682,N_19725);
and U19899 (N_19899,N_19819,N_19751);
or U19900 (N_19900,N_19708,N_19829);
nand U19901 (N_19901,N_19757,N_19836);
xor U19902 (N_19902,N_19711,N_19683);
or U19903 (N_19903,N_19687,N_19776);
xor U19904 (N_19904,N_19778,N_19824);
xor U19905 (N_19905,N_19747,N_19830);
nand U19906 (N_19906,N_19693,N_19729);
xor U19907 (N_19907,N_19702,N_19837);
xor U19908 (N_19908,N_19784,N_19821);
and U19909 (N_19909,N_19755,N_19779);
xor U19910 (N_19910,N_19809,N_19833);
or U19911 (N_19911,N_19771,N_19721);
nand U19912 (N_19912,N_19680,N_19714);
and U19913 (N_19913,N_19752,N_19717);
and U19914 (N_19914,N_19706,N_19822);
nor U19915 (N_19915,N_19785,N_19713);
or U19916 (N_19916,N_19742,N_19788);
nand U19917 (N_19917,N_19783,N_19724);
xnor U19918 (N_19918,N_19762,N_19786);
nor U19919 (N_19919,N_19732,N_19688);
xor U19920 (N_19920,N_19755,N_19705);
nor U19921 (N_19921,N_19832,N_19732);
xor U19922 (N_19922,N_19690,N_19770);
and U19923 (N_19923,N_19681,N_19781);
nor U19924 (N_19924,N_19819,N_19699);
xor U19925 (N_19925,N_19716,N_19696);
nand U19926 (N_19926,N_19836,N_19799);
nand U19927 (N_19927,N_19755,N_19778);
xnor U19928 (N_19928,N_19760,N_19691);
nand U19929 (N_19929,N_19774,N_19719);
nand U19930 (N_19930,N_19721,N_19790);
and U19931 (N_19931,N_19750,N_19720);
or U19932 (N_19932,N_19719,N_19820);
nor U19933 (N_19933,N_19734,N_19726);
or U19934 (N_19934,N_19692,N_19772);
and U19935 (N_19935,N_19728,N_19817);
nor U19936 (N_19936,N_19691,N_19686);
or U19937 (N_19937,N_19823,N_19797);
xnor U19938 (N_19938,N_19791,N_19746);
nor U19939 (N_19939,N_19823,N_19836);
nand U19940 (N_19940,N_19798,N_19819);
nand U19941 (N_19941,N_19687,N_19734);
or U19942 (N_19942,N_19722,N_19683);
or U19943 (N_19943,N_19725,N_19797);
and U19944 (N_19944,N_19800,N_19749);
nand U19945 (N_19945,N_19723,N_19789);
and U19946 (N_19946,N_19830,N_19813);
and U19947 (N_19947,N_19680,N_19724);
nand U19948 (N_19948,N_19759,N_19686);
nor U19949 (N_19949,N_19695,N_19802);
xor U19950 (N_19950,N_19738,N_19728);
nor U19951 (N_19951,N_19721,N_19767);
nor U19952 (N_19952,N_19761,N_19743);
nor U19953 (N_19953,N_19759,N_19720);
and U19954 (N_19954,N_19688,N_19723);
xor U19955 (N_19955,N_19786,N_19756);
xnor U19956 (N_19956,N_19817,N_19814);
xnor U19957 (N_19957,N_19759,N_19799);
xnor U19958 (N_19958,N_19777,N_19721);
xnor U19959 (N_19959,N_19722,N_19726);
nor U19960 (N_19960,N_19786,N_19685);
xor U19961 (N_19961,N_19731,N_19688);
xor U19962 (N_19962,N_19790,N_19816);
nand U19963 (N_19963,N_19745,N_19720);
and U19964 (N_19964,N_19801,N_19710);
xor U19965 (N_19965,N_19686,N_19789);
or U19966 (N_19966,N_19832,N_19697);
nor U19967 (N_19967,N_19761,N_19726);
xnor U19968 (N_19968,N_19773,N_19834);
or U19969 (N_19969,N_19833,N_19753);
nand U19970 (N_19970,N_19740,N_19743);
nand U19971 (N_19971,N_19720,N_19696);
nor U19972 (N_19972,N_19693,N_19746);
or U19973 (N_19973,N_19771,N_19688);
xor U19974 (N_19974,N_19824,N_19706);
and U19975 (N_19975,N_19683,N_19811);
nand U19976 (N_19976,N_19756,N_19826);
or U19977 (N_19977,N_19815,N_19825);
or U19978 (N_19978,N_19803,N_19792);
nor U19979 (N_19979,N_19734,N_19716);
nor U19980 (N_19980,N_19828,N_19710);
nor U19981 (N_19981,N_19769,N_19785);
xnor U19982 (N_19982,N_19714,N_19835);
nor U19983 (N_19983,N_19684,N_19780);
nand U19984 (N_19984,N_19792,N_19779);
nand U19985 (N_19985,N_19812,N_19728);
nand U19986 (N_19986,N_19707,N_19774);
nand U19987 (N_19987,N_19737,N_19728);
nor U19988 (N_19988,N_19744,N_19750);
or U19989 (N_19989,N_19811,N_19743);
xnor U19990 (N_19990,N_19691,N_19816);
xnor U19991 (N_19991,N_19818,N_19789);
and U19992 (N_19992,N_19798,N_19834);
and U19993 (N_19993,N_19742,N_19782);
nor U19994 (N_19994,N_19791,N_19801);
nand U19995 (N_19995,N_19741,N_19824);
xor U19996 (N_19996,N_19721,N_19822);
nand U19997 (N_19997,N_19754,N_19761);
xor U19998 (N_19998,N_19774,N_19680);
and U19999 (N_19999,N_19771,N_19700);
nand UO_0 (O_0,N_19995,N_19906);
or UO_1 (O_1,N_19880,N_19840);
and UO_2 (O_2,N_19850,N_19990);
or UO_3 (O_3,N_19941,N_19986);
nor UO_4 (O_4,N_19883,N_19930);
or UO_5 (O_5,N_19860,N_19856);
nor UO_6 (O_6,N_19846,N_19894);
nor UO_7 (O_7,N_19965,N_19936);
nor UO_8 (O_8,N_19892,N_19891);
or UO_9 (O_9,N_19976,N_19895);
or UO_10 (O_10,N_19974,N_19984);
or UO_11 (O_11,N_19862,N_19985);
nor UO_12 (O_12,N_19852,N_19954);
xor UO_13 (O_13,N_19983,N_19958);
xnor UO_14 (O_14,N_19933,N_19864);
xnor UO_15 (O_15,N_19901,N_19956);
or UO_16 (O_16,N_19874,N_19938);
nand UO_17 (O_17,N_19996,N_19855);
nand UO_18 (O_18,N_19861,N_19886);
and UO_19 (O_19,N_19848,N_19982);
or UO_20 (O_20,N_19946,N_19866);
nand UO_21 (O_21,N_19966,N_19844);
nor UO_22 (O_22,N_19929,N_19991);
nor UO_23 (O_23,N_19870,N_19942);
nor UO_24 (O_24,N_19911,N_19971);
xor UO_25 (O_25,N_19916,N_19893);
nand UO_26 (O_26,N_19845,N_19947);
nand UO_27 (O_27,N_19913,N_19900);
or UO_28 (O_28,N_19989,N_19853);
or UO_29 (O_29,N_19863,N_19920);
or UO_30 (O_30,N_19994,N_19950);
nand UO_31 (O_31,N_19872,N_19889);
and UO_32 (O_32,N_19960,N_19928);
or UO_33 (O_33,N_19973,N_19961);
and UO_34 (O_34,N_19997,N_19899);
nand UO_35 (O_35,N_19999,N_19857);
and UO_36 (O_36,N_19903,N_19843);
nor UO_37 (O_37,N_19951,N_19910);
and UO_38 (O_38,N_19885,N_19988);
nand UO_39 (O_39,N_19963,N_19915);
xnor UO_40 (O_40,N_19964,N_19878);
or UO_41 (O_41,N_19869,N_19897);
nand UO_42 (O_42,N_19905,N_19959);
or UO_43 (O_43,N_19873,N_19969);
and UO_44 (O_44,N_19858,N_19972);
or UO_45 (O_45,N_19940,N_19884);
or UO_46 (O_46,N_19948,N_19992);
or UO_47 (O_47,N_19887,N_19937);
nand UO_48 (O_48,N_19977,N_19935);
or UO_49 (O_49,N_19842,N_19865);
xor UO_50 (O_50,N_19841,N_19912);
xor UO_51 (O_51,N_19981,N_19854);
or UO_52 (O_52,N_19934,N_19904);
and UO_53 (O_53,N_19949,N_19924);
xnor UO_54 (O_54,N_19867,N_19849);
or UO_55 (O_55,N_19914,N_19952);
and UO_56 (O_56,N_19975,N_19882);
and UO_57 (O_57,N_19993,N_19922);
nor UO_58 (O_58,N_19927,N_19987);
and UO_59 (O_59,N_19909,N_19944);
xnor UO_60 (O_60,N_19888,N_19979);
xnor UO_61 (O_61,N_19881,N_19923);
xor UO_62 (O_62,N_19962,N_19896);
nand UO_63 (O_63,N_19859,N_19945);
nor UO_64 (O_64,N_19939,N_19980);
and UO_65 (O_65,N_19902,N_19925);
nor UO_66 (O_66,N_19919,N_19847);
nor UO_67 (O_67,N_19868,N_19907);
nor UO_68 (O_68,N_19879,N_19926);
xnor UO_69 (O_69,N_19851,N_19877);
nand UO_70 (O_70,N_19970,N_19875);
or UO_71 (O_71,N_19967,N_19955);
xnor UO_72 (O_72,N_19908,N_19978);
nand UO_73 (O_73,N_19968,N_19921);
nor UO_74 (O_74,N_19931,N_19943);
xnor UO_75 (O_75,N_19998,N_19876);
and UO_76 (O_76,N_19918,N_19890);
nand UO_77 (O_77,N_19953,N_19871);
and UO_78 (O_78,N_19932,N_19898);
and UO_79 (O_79,N_19917,N_19957);
and UO_80 (O_80,N_19941,N_19982);
and UO_81 (O_81,N_19873,N_19960);
nor UO_82 (O_82,N_19893,N_19875);
nor UO_83 (O_83,N_19855,N_19867);
nor UO_84 (O_84,N_19862,N_19901);
or UO_85 (O_85,N_19969,N_19975);
nand UO_86 (O_86,N_19998,N_19890);
nand UO_87 (O_87,N_19958,N_19881);
nor UO_88 (O_88,N_19922,N_19971);
nor UO_89 (O_89,N_19924,N_19849);
and UO_90 (O_90,N_19954,N_19944);
and UO_91 (O_91,N_19868,N_19969);
and UO_92 (O_92,N_19914,N_19846);
xor UO_93 (O_93,N_19963,N_19897);
nand UO_94 (O_94,N_19904,N_19849);
and UO_95 (O_95,N_19966,N_19842);
nor UO_96 (O_96,N_19902,N_19853);
or UO_97 (O_97,N_19951,N_19963);
nand UO_98 (O_98,N_19863,N_19870);
or UO_99 (O_99,N_19854,N_19928);
nand UO_100 (O_100,N_19868,N_19994);
nand UO_101 (O_101,N_19925,N_19865);
and UO_102 (O_102,N_19883,N_19936);
xor UO_103 (O_103,N_19936,N_19870);
or UO_104 (O_104,N_19925,N_19983);
or UO_105 (O_105,N_19978,N_19894);
nor UO_106 (O_106,N_19921,N_19902);
and UO_107 (O_107,N_19878,N_19945);
nor UO_108 (O_108,N_19850,N_19909);
and UO_109 (O_109,N_19946,N_19852);
nand UO_110 (O_110,N_19841,N_19885);
and UO_111 (O_111,N_19925,N_19894);
nor UO_112 (O_112,N_19855,N_19898);
xnor UO_113 (O_113,N_19934,N_19916);
and UO_114 (O_114,N_19955,N_19944);
nand UO_115 (O_115,N_19946,N_19896);
or UO_116 (O_116,N_19939,N_19983);
or UO_117 (O_117,N_19956,N_19914);
nor UO_118 (O_118,N_19887,N_19890);
and UO_119 (O_119,N_19979,N_19985);
and UO_120 (O_120,N_19960,N_19859);
or UO_121 (O_121,N_19913,N_19922);
and UO_122 (O_122,N_19971,N_19840);
xor UO_123 (O_123,N_19981,N_19868);
xnor UO_124 (O_124,N_19957,N_19942);
or UO_125 (O_125,N_19860,N_19967);
or UO_126 (O_126,N_19864,N_19963);
and UO_127 (O_127,N_19849,N_19936);
or UO_128 (O_128,N_19896,N_19845);
nor UO_129 (O_129,N_19860,N_19904);
nand UO_130 (O_130,N_19885,N_19976);
nor UO_131 (O_131,N_19954,N_19919);
or UO_132 (O_132,N_19931,N_19865);
nor UO_133 (O_133,N_19995,N_19940);
and UO_134 (O_134,N_19845,N_19999);
and UO_135 (O_135,N_19857,N_19974);
xor UO_136 (O_136,N_19942,N_19926);
nor UO_137 (O_137,N_19934,N_19905);
or UO_138 (O_138,N_19949,N_19867);
or UO_139 (O_139,N_19841,N_19852);
nand UO_140 (O_140,N_19897,N_19902);
xor UO_141 (O_141,N_19871,N_19987);
and UO_142 (O_142,N_19908,N_19910);
xor UO_143 (O_143,N_19985,N_19952);
xnor UO_144 (O_144,N_19938,N_19931);
xnor UO_145 (O_145,N_19916,N_19990);
and UO_146 (O_146,N_19869,N_19905);
or UO_147 (O_147,N_19857,N_19948);
nand UO_148 (O_148,N_19961,N_19874);
nand UO_149 (O_149,N_19909,N_19913);
nand UO_150 (O_150,N_19860,N_19943);
and UO_151 (O_151,N_19966,N_19865);
xor UO_152 (O_152,N_19997,N_19960);
xnor UO_153 (O_153,N_19958,N_19906);
nor UO_154 (O_154,N_19938,N_19918);
and UO_155 (O_155,N_19861,N_19905);
xor UO_156 (O_156,N_19994,N_19899);
xnor UO_157 (O_157,N_19843,N_19896);
nor UO_158 (O_158,N_19994,N_19999);
and UO_159 (O_159,N_19889,N_19897);
xnor UO_160 (O_160,N_19947,N_19992);
and UO_161 (O_161,N_19844,N_19916);
xnor UO_162 (O_162,N_19856,N_19970);
nor UO_163 (O_163,N_19880,N_19913);
nor UO_164 (O_164,N_19978,N_19907);
xor UO_165 (O_165,N_19997,N_19921);
nand UO_166 (O_166,N_19928,N_19991);
xor UO_167 (O_167,N_19958,N_19933);
nand UO_168 (O_168,N_19963,N_19968);
or UO_169 (O_169,N_19854,N_19868);
and UO_170 (O_170,N_19863,N_19850);
xor UO_171 (O_171,N_19956,N_19955);
nor UO_172 (O_172,N_19953,N_19947);
nor UO_173 (O_173,N_19984,N_19921);
and UO_174 (O_174,N_19986,N_19879);
and UO_175 (O_175,N_19912,N_19942);
nand UO_176 (O_176,N_19949,N_19869);
nand UO_177 (O_177,N_19994,N_19861);
or UO_178 (O_178,N_19991,N_19908);
and UO_179 (O_179,N_19910,N_19914);
and UO_180 (O_180,N_19900,N_19973);
nor UO_181 (O_181,N_19995,N_19988);
xor UO_182 (O_182,N_19850,N_19910);
xor UO_183 (O_183,N_19927,N_19906);
and UO_184 (O_184,N_19895,N_19841);
and UO_185 (O_185,N_19883,N_19947);
xnor UO_186 (O_186,N_19967,N_19895);
and UO_187 (O_187,N_19928,N_19845);
or UO_188 (O_188,N_19918,N_19862);
xor UO_189 (O_189,N_19889,N_19866);
nor UO_190 (O_190,N_19981,N_19900);
and UO_191 (O_191,N_19848,N_19902);
nand UO_192 (O_192,N_19884,N_19954);
nor UO_193 (O_193,N_19919,N_19904);
nand UO_194 (O_194,N_19879,N_19935);
and UO_195 (O_195,N_19925,N_19966);
and UO_196 (O_196,N_19877,N_19969);
nand UO_197 (O_197,N_19906,N_19942);
nor UO_198 (O_198,N_19860,N_19911);
and UO_199 (O_199,N_19959,N_19898);
nor UO_200 (O_200,N_19974,N_19921);
nor UO_201 (O_201,N_19851,N_19941);
nand UO_202 (O_202,N_19979,N_19875);
nand UO_203 (O_203,N_19969,N_19871);
xnor UO_204 (O_204,N_19987,N_19933);
xnor UO_205 (O_205,N_19908,N_19960);
and UO_206 (O_206,N_19898,N_19903);
xnor UO_207 (O_207,N_19840,N_19918);
nand UO_208 (O_208,N_19969,N_19847);
nand UO_209 (O_209,N_19929,N_19867);
nor UO_210 (O_210,N_19926,N_19849);
xor UO_211 (O_211,N_19921,N_19886);
nor UO_212 (O_212,N_19999,N_19932);
xnor UO_213 (O_213,N_19877,N_19929);
and UO_214 (O_214,N_19879,N_19942);
xnor UO_215 (O_215,N_19875,N_19980);
nand UO_216 (O_216,N_19842,N_19934);
and UO_217 (O_217,N_19994,N_19974);
or UO_218 (O_218,N_19997,N_19852);
and UO_219 (O_219,N_19900,N_19903);
or UO_220 (O_220,N_19971,N_19964);
or UO_221 (O_221,N_19977,N_19840);
nand UO_222 (O_222,N_19872,N_19946);
nor UO_223 (O_223,N_19973,N_19865);
nand UO_224 (O_224,N_19847,N_19848);
nand UO_225 (O_225,N_19949,N_19845);
xnor UO_226 (O_226,N_19885,N_19899);
nor UO_227 (O_227,N_19862,N_19914);
nand UO_228 (O_228,N_19988,N_19858);
nor UO_229 (O_229,N_19964,N_19922);
xnor UO_230 (O_230,N_19967,N_19907);
nor UO_231 (O_231,N_19974,N_19922);
xor UO_232 (O_232,N_19964,N_19890);
nand UO_233 (O_233,N_19987,N_19953);
nand UO_234 (O_234,N_19904,N_19963);
nand UO_235 (O_235,N_19932,N_19982);
nand UO_236 (O_236,N_19940,N_19943);
xor UO_237 (O_237,N_19916,N_19987);
nand UO_238 (O_238,N_19949,N_19890);
nand UO_239 (O_239,N_19853,N_19929);
nand UO_240 (O_240,N_19946,N_19887);
xnor UO_241 (O_241,N_19975,N_19886);
nor UO_242 (O_242,N_19975,N_19971);
and UO_243 (O_243,N_19986,N_19884);
nor UO_244 (O_244,N_19995,N_19904);
nand UO_245 (O_245,N_19885,N_19849);
nor UO_246 (O_246,N_19980,N_19937);
nor UO_247 (O_247,N_19917,N_19905);
nor UO_248 (O_248,N_19918,N_19989);
or UO_249 (O_249,N_19970,N_19906);
xor UO_250 (O_250,N_19900,N_19867);
nor UO_251 (O_251,N_19845,N_19901);
or UO_252 (O_252,N_19877,N_19919);
nand UO_253 (O_253,N_19936,N_19860);
or UO_254 (O_254,N_19846,N_19926);
nand UO_255 (O_255,N_19956,N_19951);
or UO_256 (O_256,N_19899,N_19887);
xor UO_257 (O_257,N_19981,N_19917);
nor UO_258 (O_258,N_19892,N_19866);
nor UO_259 (O_259,N_19988,N_19846);
and UO_260 (O_260,N_19972,N_19955);
and UO_261 (O_261,N_19938,N_19932);
or UO_262 (O_262,N_19909,N_19914);
and UO_263 (O_263,N_19981,N_19843);
nand UO_264 (O_264,N_19890,N_19959);
nand UO_265 (O_265,N_19983,N_19948);
nor UO_266 (O_266,N_19840,N_19986);
and UO_267 (O_267,N_19902,N_19941);
or UO_268 (O_268,N_19945,N_19910);
and UO_269 (O_269,N_19927,N_19934);
and UO_270 (O_270,N_19842,N_19947);
nor UO_271 (O_271,N_19948,N_19985);
xor UO_272 (O_272,N_19897,N_19923);
nand UO_273 (O_273,N_19993,N_19933);
nor UO_274 (O_274,N_19970,N_19903);
xnor UO_275 (O_275,N_19911,N_19920);
and UO_276 (O_276,N_19899,N_19976);
and UO_277 (O_277,N_19903,N_19883);
nor UO_278 (O_278,N_19864,N_19995);
or UO_279 (O_279,N_19885,N_19997);
nand UO_280 (O_280,N_19981,N_19916);
and UO_281 (O_281,N_19979,N_19950);
or UO_282 (O_282,N_19972,N_19889);
nand UO_283 (O_283,N_19862,N_19953);
nor UO_284 (O_284,N_19926,N_19999);
nand UO_285 (O_285,N_19853,N_19947);
and UO_286 (O_286,N_19970,N_19923);
nor UO_287 (O_287,N_19934,N_19847);
xnor UO_288 (O_288,N_19847,N_19986);
xnor UO_289 (O_289,N_19880,N_19918);
xnor UO_290 (O_290,N_19945,N_19871);
xor UO_291 (O_291,N_19963,N_19959);
and UO_292 (O_292,N_19866,N_19977);
nor UO_293 (O_293,N_19973,N_19873);
nand UO_294 (O_294,N_19877,N_19952);
nor UO_295 (O_295,N_19877,N_19861);
nand UO_296 (O_296,N_19925,N_19922);
nand UO_297 (O_297,N_19901,N_19989);
and UO_298 (O_298,N_19916,N_19909);
or UO_299 (O_299,N_19970,N_19841);
nor UO_300 (O_300,N_19842,N_19962);
or UO_301 (O_301,N_19875,N_19858);
and UO_302 (O_302,N_19933,N_19906);
xnor UO_303 (O_303,N_19847,N_19907);
xor UO_304 (O_304,N_19915,N_19966);
and UO_305 (O_305,N_19903,N_19965);
nand UO_306 (O_306,N_19986,N_19846);
nor UO_307 (O_307,N_19905,N_19907);
xnor UO_308 (O_308,N_19852,N_19956);
nand UO_309 (O_309,N_19900,N_19974);
or UO_310 (O_310,N_19984,N_19862);
and UO_311 (O_311,N_19941,N_19927);
or UO_312 (O_312,N_19986,N_19909);
or UO_313 (O_313,N_19941,N_19865);
or UO_314 (O_314,N_19851,N_19855);
or UO_315 (O_315,N_19860,N_19973);
or UO_316 (O_316,N_19976,N_19959);
or UO_317 (O_317,N_19876,N_19884);
nand UO_318 (O_318,N_19930,N_19975);
and UO_319 (O_319,N_19890,N_19907);
nor UO_320 (O_320,N_19868,N_19944);
and UO_321 (O_321,N_19990,N_19851);
nor UO_322 (O_322,N_19943,N_19885);
nand UO_323 (O_323,N_19889,N_19910);
nor UO_324 (O_324,N_19867,N_19975);
nor UO_325 (O_325,N_19980,N_19975);
or UO_326 (O_326,N_19963,N_19975);
and UO_327 (O_327,N_19841,N_19856);
or UO_328 (O_328,N_19885,N_19871);
xnor UO_329 (O_329,N_19842,N_19907);
nand UO_330 (O_330,N_19933,N_19890);
nand UO_331 (O_331,N_19850,N_19856);
or UO_332 (O_332,N_19999,N_19986);
or UO_333 (O_333,N_19959,N_19846);
or UO_334 (O_334,N_19944,N_19862);
nor UO_335 (O_335,N_19973,N_19985);
nand UO_336 (O_336,N_19910,N_19947);
nor UO_337 (O_337,N_19947,N_19988);
nand UO_338 (O_338,N_19886,N_19894);
and UO_339 (O_339,N_19957,N_19873);
xnor UO_340 (O_340,N_19950,N_19865);
xnor UO_341 (O_341,N_19893,N_19919);
and UO_342 (O_342,N_19974,N_19854);
nor UO_343 (O_343,N_19938,N_19963);
or UO_344 (O_344,N_19897,N_19950);
nor UO_345 (O_345,N_19907,N_19911);
xor UO_346 (O_346,N_19856,N_19990);
nor UO_347 (O_347,N_19970,N_19952);
nand UO_348 (O_348,N_19885,N_19888);
and UO_349 (O_349,N_19909,N_19848);
xor UO_350 (O_350,N_19882,N_19863);
or UO_351 (O_351,N_19978,N_19903);
or UO_352 (O_352,N_19868,N_19954);
or UO_353 (O_353,N_19970,N_19911);
or UO_354 (O_354,N_19917,N_19996);
or UO_355 (O_355,N_19959,N_19943);
nor UO_356 (O_356,N_19911,N_19864);
or UO_357 (O_357,N_19895,N_19940);
nand UO_358 (O_358,N_19997,N_19905);
nand UO_359 (O_359,N_19966,N_19923);
nand UO_360 (O_360,N_19972,N_19913);
nand UO_361 (O_361,N_19989,N_19996);
and UO_362 (O_362,N_19914,N_19979);
and UO_363 (O_363,N_19997,N_19931);
and UO_364 (O_364,N_19915,N_19954);
nor UO_365 (O_365,N_19926,N_19871);
or UO_366 (O_366,N_19873,N_19847);
and UO_367 (O_367,N_19972,N_19890);
nand UO_368 (O_368,N_19871,N_19893);
nand UO_369 (O_369,N_19926,N_19922);
and UO_370 (O_370,N_19977,N_19899);
and UO_371 (O_371,N_19943,N_19889);
xor UO_372 (O_372,N_19987,N_19995);
nand UO_373 (O_373,N_19966,N_19959);
nand UO_374 (O_374,N_19856,N_19846);
nand UO_375 (O_375,N_19975,N_19967);
nor UO_376 (O_376,N_19891,N_19984);
xnor UO_377 (O_377,N_19927,N_19967);
and UO_378 (O_378,N_19889,N_19880);
nor UO_379 (O_379,N_19958,N_19951);
nor UO_380 (O_380,N_19861,N_19850);
or UO_381 (O_381,N_19975,N_19987);
and UO_382 (O_382,N_19954,N_19910);
and UO_383 (O_383,N_19979,N_19862);
nand UO_384 (O_384,N_19902,N_19939);
xor UO_385 (O_385,N_19864,N_19898);
nand UO_386 (O_386,N_19962,N_19977);
and UO_387 (O_387,N_19858,N_19908);
xor UO_388 (O_388,N_19898,N_19972);
nor UO_389 (O_389,N_19899,N_19908);
nor UO_390 (O_390,N_19922,N_19991);
nor UO_391 (O_391,N_19926,N_19881);
xor UO_392 (O_392,N_19936,N_19862);
xor UO_393 (O_393,N_19852,N_19967);
nor UO_394 (O_394,N_19991,N_19969);
xnor UO_395 (O_395,N_19998,N_19945);
or UO_396 (O_396,N_19937,N_19926);
and UO_397 (O_397,N_19855,N_19987);
nor UO_398 (O_398,N_19880,N_19853);
xnor UO_399 (O_399,N_19861,N_19961);
xnor UO_400 (O_400,N_19999,N_19955);
nand UO_401 (O_401,N_19945,N_19970);
nor UO_402 (O_402,N_19853,N_19895);
nor UO_403 (O_403,N_19955,N_19973);
xor UO_404 (O_404,N_19981,N_19982);
xor UO_405 (O_405,N_19864,N_19916);
nand UO_406 (O_406,N_19918,N_19966);
and UO_407 (O_407,N_19896,N_19884);
nor UO_408 (O_408,N_19939,N_19998);
or UO_409 (O_409,N_19869,N_19843);
xor UO_410 (O_410,N_19873,N_19917);
nand UO_411 (O_411,N_19895,N_19881);
and UO_412 (O_412,N_19938,N_19885);
nand UO_413 (O_413,N_19987,N_19991);
nor UO_414 (O_414,N_19851,N_19982);
and UO_415 (O_415,N_19955,N_19855);
nor UO_416 (O_416,N_19840,N_19955);
xnor UO_417 (O_417,N_19943,N_19898);
and UO_418 (O_418,N_19853,N_19955);
xnor UO_419 (O_419,N_19956,N_19881);
nor UO_420 (O_420,N_19922,N_19851);
nor UO_421 (O_421,N_19966,N_19873);
xor UO_422 (O_422,N_19961,N_19932);
and UO_423 (O_423,N_19956,N_19843);
xnor UO_424 (O_424,N_19983,N_19877);
nand UO_425 (O_425,N_19844,N_19891);
nand UO_426 (O_426,N_19965,N_19998);
xnor UO_427 (O_427,N_19934,N_19973);
xor UO_428 (O_428,N_19959,N_19930);
xnor UO_429 (O_429,N_19892,N_19952);
nor UO_430 (O_430,N_19917,N_19907);
nand UO_431 (O_431,N_19941,N_19918);
nand UO_432 (O_432,N_19946,N_19947);
nand UO_433 (O_433,N_19915,N_19973);
or UO_434 (O_434,N_19850,N_19895);
xnor UO_435 (O_435,N_19875,N_19998);
nand UO_436 (O_436,N_19966,N_19909);
nor UO_437 (O_437,N_19857,N_19906);
and UO_438 (O_438,N_19999,N_19934);
and UO_439 (O_439,N_19998,N_19925);
xnor UO_440 (O_440,N_19905,N_19928);
nand UO_441 (O_441,N_19965,N_19910);
or UO_442 (O_442,N_19932,N_19896);
xor UO_443 (O_443,N_19965,N_19854);
and UO_444 (O_444,N_19908,N_19962);
and UO_445 (O_445,N_19859,N_19961);
xnor UO_446 (O_446,N_19975,N_19990);
and UO_447 (O_447,N_19989,N_19864);
and UO_448 (O_448,N_19993,N_19842);
and UO_449 (O_449,N_19966,N_19945);
nor UO_450 (O_450,N_19993,N_19966);
nand UO_451 (O_451,N_19883,N_19989);
and UO_452 (O_452,N_19998,N_19894);
nor UO_453 (O_453,N_19948,N_19902);
xnor UO_454 (O_454,N_19946,N_19975);
and UO_455 (O_455,N_19942,N_19848);
and UO_456 (O_456,N_19950,N_19955);
xor UO_457 (O_457,N_19954,N_19854);
and UO_458 (O_458,N_19964,N_19993);
xnor UO_459 (O_459,N_19891,N_19934);
xor UO_460 (O_460,N_19952,N_19910);
nand UO_461 (O_461,N_19950,N_19921);
nor UO_462 (O_462,N_19956,N_19944);
or UO_463 (O_463,N_19988,N_19919);
nand UO_464 (O_464,N_19870,N_19965);
nor UO_465 (O_465,N_19960,N_19970);
or UO_466 (O_466,N_19995,N_19967);
nor UO_467 (O_467,N_19851,N_19841);
or UO_468 (O_468,N_19937,N_19891);
and UO_469 (O_469,N_19870,N_19842);
or UO_470 (O_470,N_19843,N_19977);
nand UO_471 (O_471,N_19936,N_19880);
and UO_472 (O_472,N_19890,N_19951);
xnor UO_473 (O_473,N_19890,N_19980);
and UO_474 (O_474,N_19859,N_19894);
or UO_475 (O_475,N_19901,N_19977);
xnor UO_476 (O_476,N_19905,N_19859);
or UO_477 (O_477,N_19857,N_19885);
and UO_478 (O_478,N_19914,N_19942);
or UO_479 (O_479,N_19857,N_19841);
nor UO_480 (O_480,N_19943,N_19956);
xor UO_481 (O_481,N_19925,N_19993);
nor UO_482 (O_482,N_19918,N_19937);
nand UO_483 (O_483,N_19998,N_19889);
xor UO_484 (O_484,N_19942,N_19932);
nor UO_485 (O_485,N_19858,N_19963);
or UO_486 (O_486,N_19962,N_19960);
and UO_487 (O_487,N_19973,N_19880);
nor UO_488 (O_488,N_19940,N_19978);
or UO_489 (O_489,N_19931,N_19932);
xor UO_490 (O_490,N_19862,N_19941);
xor UO_491 (O_491,N_19956,N_19877);
nand UO_492 (O_492,N_19872,N_19869);
and UO_493 (O_493,N_19858,N_19952);
xnor UO_494 (O_494,N_19964,N_19859);
nand UO_495 (O_495,N_19927,N_19985);
or UO_496 (O_496,N_19846,N_19971);
and UO_497 (O_497,N_19903,N_19849);
or UO_498 (O_498,N_19986,N_19926);
xor UO_499 (O_499,N_19852,N_19923);
and UO_500 (O_500,N_19859,N_19846);
and UO_501 (O_501,N_19902,N_19970);
nor UO_502 (O_502,N_19868,N_19899);
nor UO_503 (O_503,N_19987,N_19949);
nand UO_504 (O_504,N_19929,N_19985);
and UO_505 (O_505,N_19875,N_19994);
or UO_506 (O_506,N_19902,N_19845);
nor UO_507 (O_507,N_19939,N_19929);
nand UO_508 (O_508,N_19946,N_19941);
or UO_509 (O_509,N_19978,N_19994);
xnor UO_510 (O_510,N_19993,N_19924);
or UO_511 (O_511,N_19899,N_19852);
nand UO_512 (O_512,N_19942,N_19943);
or UO_513 (O_513,N_19952,N_19944);
or UO_514 (O_514,N_19877,N_19872);
and UO_515 (O_515,N_19942,N_19874);
nand UO_516 (O_516,N_19878,N_19900);
xor UO_517 (O_517,N_19905,N_19998);
nand UO_518 (O_518,N_19961,N_19921);
and UO_519 (O_519,N_19887,N_19919);
nor UO_520 (O_520,N_19932,N_19849);
and UO_521 (O_521,N_19869,N_19968);
xor UO_522 (O_522,N_19905,N_19852);
and UO_523 (O_523,N_19883,N_19847);
xor UO_524 (O_524,N_19872,N_19891);
nand UO_525 (O_525,N_19918,N_19928);
and UO_526 (O_526,N_19999,N_19894);
nand UO_527 (O_527,N_19890,N_19898);
nor UO_528 (O_528,N_19953,N_19920);
or UO_529 (O_529,N_19844,N_19860);
xor UO_530 (O_530,N_19927,N_19983);
or UO_531 (O_531,N_19986,N_19889);
and UO_532 (O_532,N_19965,N_19950);
xnor UO_533 (O_533,N_19995,N_19976);
and UO_534 (O_534,N_19847,N_19956);
nand UO_535 (O_535,N_19924,N_19848);
nand UO_536 (O_536,N_19893,N_19917);
or UO_537 (O_537,N_19876,N_19873);
or UO_538 (O_538,N_19895,N_19843);
xnor UO_539 (O_539,N_19899,N_19842);
or UO_540 (O_540,N_19973,N_19896);
xnor UO_541 (O_541,N_19897,N_19857);
or UO_542 (O_542,N_19975,N_19850);
or UO_543 (O_543,N_19933,N_19907);
nor UO_544 (O_544,N_19986,N_19843);
or UO_545 (O_545,N_19854,N_19984);
nand UO_546 (O_546,N_19908,N_19856);
xor UO_547 (O_547,N_19873,N_19880);
nor UO_548 (O_548,N_19996,N_19967);
xnor UO_549 (O_549,N_19931,N_19898);
nand UO_550 (O_550,N_19929,N_19881);
xnor UO_551 (O_551,N_19999,N_19978);
and UO_552 (O_552,N_19897,N_19952);
nor UO_553 (O_553,N_19993,N_19893);
xor UO_554 (O_554,N_19902,N_19932);
nor UO_555 (O_555,N_19917,N_19894);
or UO_556 (O_556,N_19961,N_19856);
nor UO_557 (O_557,N_19879,N_19924);
or UO_558 (O_558,N_19963,N_19856);
xnor UO_559 (O_559,N_19848,N_19934);
and UO_560 (O_560,N_19865,N_19871);
and UO_561 (O_561,N_19897,N_19961);
nand UO_562 (O_562,N_19881,N_19854);
nand UO_563 (O_563,N_19947,N_19939);
nand UO_564 (O_564,N_19954,N_19873);
and UO_565 (O_565,N_19840,N_19872);
xnor UO_566 (O_566,N_19913,N_19997);
nand UO_567 (O_567,N_19855,N_19980);
nand UO_568 (O_568,N_19945,N_19990);
xor UO_569 (O_569,N_19965,N_19869);
or UO_570 (O_570,N_19984,N_19992);
xnor UO_571 (O_571,N_19961,N_19935);
and UO_572 (O_572,N_19907,N_19852);
nor UO_573 (O_573,N_19909,N_19946);
and UO_574 (O_574,N_19886,N_19856);
or UO_575 (O_575,N_19850,N_19878);
xnor UO_576 (O_576,N_19971,N_19903);
and UO_577 (O_577,N_19907,N_19961);
and UO_578 (O_578,N_19938,N_19878);
nand UO_579 (O_579,N_19931,N_19851);
nor UO_580 (O_580,N_19884,N_19883);
nor UO_581 (O_581,N_19914,N_19993);
nand UO_582 (O_582,N_19977,N_19971);
and UO_583 (O_583,N_19917,N_19845);
and UO_584 (O_584,N_19850,N_19906);
and UO_585 (O_585,N_19997,N_19866);
nand UO_586 (O_586,N_19934,N_19876);
nor UO_587 (O_587,N_19883,N_19946);
nand UO_588 (O_588,N_19874,N_19881);
xnor UO_589 (O_589,N_19937,N_19902);
or UO_590 (O_590,N_19843,N_19866);
or UO_591 (O_591,N_19943,N_19920);
xor UO_592 (O_592,N_19906,N_19941);
and UO_593 (O_593,N_19846,N_19913);
nor UO_594 (O_594,N_19867,N_19896);
and UO_595 (O_595,N_19901,N_19865);
nand UO_596 (O_596,N_19954,N_19963);
or UO_597 (O_597,N_19850,N_19849);
nor UO_598 (O_598,N_19896,N_19856);
xor UO_599 (O_599,N_19981,N_19920);
xnor UO_600 (O_600,N_19947,N_19952);
nor UO_601 (O_601,N_19866,N_19846);
or UO_602 (O_602,N_19868,N_19913);
xor UO_603 (O_603,N_19905,N_19992);
nand UO_604 (O_604,N_19929,N_19989);
nand UO_605 (O_605,N_19932,N_19847);
nand UO_606 (O_606,N_19851,N_19934);
xnor UO_607 (O_607,N_19856,N_19926);
or UO_608 (O_608,N_19971,N_19979);
and UO_609 (O_609,N_19933,N_19973);
or UO_610 (O_610,N_19957,N_19922);
or UO_611 (O_611,N_19963,N_19950);
and UO_612 (O_612,N_19850,N_19926);
or UO_613 (O_613,N_19958,N_19910);
or UO_614 (O_614,N_19845,N_19970);
or UO_615 (O_615,N_19860,N_19948);
nor UO_616 (O_616,N_19952,N_19915);
nand UO_617 (O_617,N_19992,N_19987);
nor UO_618 (O_618,N_19887,N_19983);
nand UO_619 (O_619,N_19909,N_19891);
and UO_620 (O_620,N_19902,N_19863);
nor UO_621 (O_621,N_19957,N_19887);
xor UO_622 (O_622,N_19938,N_19877);
and UO_623 (O_623,N_19854,N_19847);
xor UO_624 (O_624,N_19946,N_19952);
xor UO_625 (O_625,N_19944,N_19960);
and UO_626 (O_626,N_19855,N_19885);
and UO_627 (O_627,N_19853,N_19973);
or UO_628 (O_628,N_19995,N_19992);
and UO_629 (O_629,N_19852,N_19876);
nor UO_630 (O_630,N_19996,N_19844);
nor UO_631 (O_631,N_19859,N_19911);
and UO_632 (O_632,N_19911,N_19874);
xnor UO_633 (O_633,N_19921,N_19881);
nor UO_634 (O_634,N_19934,N_19870);
nand UO_635 (O_635,N_19853,N_19936);
nor UO_636 (O_636,N_19858,N_19891);
or UO_637 (O_637,N_19842,N_19990);
xnor UO_638 (O_638,N_19971,N_19937);
nor UO_639 (O_639,N_19872,N_19933);
xor UO_640 (O_640,N_19916,N_19931);
or UO_641 (O_641,N_19858,N_19993);
or UO_642 (O_642,N_19990,N_19857);
and UO_643 (O_643,N_19899,N_19947);
or UO_644 (O_644,N_19881,N_19855);
or UO_645 (O_645,N_19923,N_19860);
nor UO_646 (O_646,N_19934,N_19908);
or UO_647 (O_647,N_19874,N_19974);
nor UO_648 (O_648,N_19982,N_19938);
xor UO_649 (O_649,N_19910,N_19866);
xor UO_650 (O_650,N_19975,N_19970);
nor UO_651 (O_651,N_19848,N_19868);
and UO_652 (O_652,N_19845,N_19967);
nand UO_653 (O_653,N_19966,N_19903);
xnor UO_654 (O_654,N_19919,N_19943);
xor UO_655 (O_655,N_19941,N_19864);
and UO_656 (O_656,N_19861,N_19949);
or UO_657 (O_657,N_19860,N_19862);
xor UO_658 (O_658,N_19889,N_19982);
or UO_659 (O_659,N_19843,N_19940);
or UO_660 (O_660,N_19973,N_19851);
xor UO_661 (O_661,N_19953,N_19911);
xnor UO_662 (O_662,N_19895,N_19930);
and UO_663 (O_663,N_19965,N_19954);
and UO_664 (O_664,N_19899,N_19917);
xor UO_665 (O_665,N_19903,N_19972);
nand UO_666 (O_666,N_19878,N_19954);
or UO_667 (O_667,N_19922,N_19889);
or UO_668 (O_668,N_19980,N_19888);
and UO_669 (O_669,N_19954,N_19885);
xor UO_670 (O_670,N_19927,N_19909);
and UO_671 (O_671,N_19848,N_19901);
and UO_672 (O_672,N_19891,N_19975);
xor UO_673 (O_673,N_19871,N_19997);
nand UO_674 (O_674,N_19859,N_19925);
nand UO_675 (O_675,N_19912,N_19880);
xnor UO_676 (O_676,N_19882,N_19891);
and UO_677 (O_677,N_19999,N_19907);
xnor UO_678 (O_678,N_19974,N_19937);
nand UO_679 (O_679,N_19998,N_19940);
and UO_680 (O_680,N_19999,N_19941);
xor UO_681 (O_681,N_19933,N_19898);
xor UO_682 (O_682,N_19907,N_19925);
nor UO_683 (O_683,N_19925,N_19895);
nand UO_684 (O_684,N_19888,N_19848);
or UO_685 (O_685,N_19986,N_19891);
nand UO_686 (O_686,N_19876,N_19879);
xnor UO_687 (O_687,N_19957,N_19850);
nand UO_688 (O_688,N_19989,N_19891);
nand UO_689 (O_689,N_19926,N_19997);
or UO_690 (O_690,N_19919,N_19846);
nand UO_691 (O_691,N_19966,N_19857);
nor UO_692 (O_692,N_19843,N_19913);
and UO_693 (O_693,N_19877,N_19985);
nor UO_694 (O_694,N_19927,N_19966);
nand UO_695 (O_695,N_19947,N_19969);
xor UO_696 (O_696,N_19973,N_19861);
nand UO_697 (O_697,N_19894,N_19885);
xor UO_698 (O_698,N_19924,N_19843);
xnor UO_699 (O_699,N_19910,N_19960);
and UO_700 (O_700,N_19923,N_19936);
or UO_701 (O_701,N_19847,N_19911);
xnor UO_702 (O_702,N_19876,N_19862);
nor UO_703 (O_703,N_19917,N_19862);
nand UO_704 (O_704,N_19844,N_19873);
nor UO_705 (O_705,N_19981,N_19992);
nand UO_706 (O_706,N_19925,N_19851);
xnor UO_707 (O_707,N_19947,N_19972);
xor UO_708 (O_708,N_19959,N_19903);
xor UO_709 (O_709,N_19947,N_19923);
or UO_710 (O_710,N_19997,N_19888);
and UO_711 (O_711,N_19935,N_19889);
xor UO_712 (O_712,N_19949,N_19911);
and UO_713 (O_713,N_19960,N_19967);
or UO_714 (O_714,N_19973,N_19988);
or UO_715 (O_715,N_19981,N_19875);
or UO_716 (O_716,N_19873,N_19851);
nor UO_717 (O_717,N_19901,N_19997);
and UO_718 (O_718,N_19972,N_19900);
nand UO_719 (O_719,N_19929,N_19844);
or UO_720 (O_720,N_19890,N_19986);
xnor UO_721 (O_721,N_19845,N_19879);
or UO_722 (O_722,N_19842,N_19923);
nor UO_723 (O_723,N_19999,N_19943);
xor UO_724 (O_724,N_19967,N_19894);
and UO_725 (O_725,N_19934,N_19864);
xnor UO_726 (O_726,N_19958,N_19944);
or UO_727 (O_727,N_19864,N_19871);
nand UO_728 (O_728,N_19902,N_19917);
xor UO_729 (O_729,N_19953,N_19954);
and UO_730 (O_730,N_19938,N_19923);
and UO_731 (O_731,N_19893,N_19891);
nand UO_732 (O_732,N_19924,N_19947);
nor UO_733 (O_733,N_19934,N_19917);
xnor UO_734 (O_734,N_19971,N_19962);
and UO_735 (O_735,N_19966,N_19967);
xnor UO_736 (O_736,N_19998,N_19962);
nor UO_737 (O_737,N_19898,N_19840);
xnor UO_738 (O_738,N_19971,N_19919);
or UO_739 (O_739,N_19997,N_19874);
or UO_740 (O_740,N_19862,N_19932);
nor UO_741 (O_741,N_19918,N_19899);
nand UO_742 (O_742,N_19933,N_19875);
xnor UO_743 (O_743,N_19990,N_19954);
xnor UO_744 (O_744,N_19874,N_19919);
nand UO_745 (O_745,N_19974,N_19948);
and UO_746 (O_746,N_19929,N_19963);
and UO_747 (O_747,N_19849,N_19922);
xor UO_748 (O_748,N_19996,N_19994);
xnor UO_749 (O_749,N_19987,N_19863);
or UO_750 (O_750,N_19874,N_19853);
nor UO_751 (O_751,N_19985,N_19841);
or UO_752 (O_752,N_19890,N_19999);
and UO_753 (O_753,N_19972,N_19935);
nor UO_754 (O_754,N_19925,N_19857);
nor UO_755 (O_755,N_19892,N_19983);
xnor UO_756 (O_756,N_19886,N_19884);
xnor UO_757 (O_757,N_19941,N_19875);
and UO_758 (O_758,N_19999,N_19930);
nor UO_759 (O_759,N_19976,N_19999);
nor UO_760 (O_760,N_19930,N_19958);
nor UO_761 (O_761,N_19918,N_19855);
xnor UO_762 (O_762,N_19917,N_19938);
nand UO_763 (O_763,N_19982,N_19879);
xnor UO_764 (O_764,N_19845,N_19939);
nor UO_765 (O_765,N_19880,N_19920);
or UO_766 (O_766,N_19927,N_19890);
or UO_767 (O_767,N_19949,N_19995);
nand UO_768 (O_768,N_19873,N_19932);
nand UO_769 (O_769,N_19970,N_19880);
or UO_770 (O_770,N_19844,N_19885);
and UO_771 (O_771,N_19986,N_19957);
or UO_772 (O_772,N_19858,N_19884);
or UO_773 (O_773,N_19969,N_19979);
and UO_774 (O_774,N_19901,N_19852);
or UO_775 (O_775,N_19947,N_19912);
xor UO_776 (O_776,N_19951,N_19917);
nand UO_777 (O_777,N_19940,N_19864);
and UO_778 (O_778,N_19954,N_19861);
nor UO_779 (O_779,N_19881,N_19996);
nand UO_780 (O_780,N_19996,N_19953);
and UO_781 (O_781,N_19910,N_19948);
or UO_782 (O_782,N_19916,N_19933);
and UO_783 (O_783,N_19920,N_19888);
and UO_784 (O_784,N_19963,N_19857);
xor UO_785 (O_785,N_19878,N_19967);
xor UO_786 (O_786,N_19840,N_19907);
nor UO_787 (O_787,N_19939,N_19881);
nor UO_788 (O_788,N_19922,N_19930);
nand UO_789 (O_789,N_19899,N_19969);
or UO_790 (O_790,N_19889,N_19931);
and UO_791 (O_791,N_19978,N_19979);
and UO_792 (O_792,N_19849,N_19859);
or UO_793 (O_793,N_19850,N_19991);
xor UO_794 (O_794,N_19933,N_19862);
and UO_795 (O_795,N_19970,N_19904);
xnor UO_796 (O_796,N_19977,N_19988);
nand UO_797 (O_797,N_19907,N_19886);
nor UO_798 (O_798,N_19983,N_19995);
nor UO_799 (O_799,N_19982,N_19917);
nor UO_800 (O_800,N_19986,N_19906);
nor UO_801 (O_801,N_19889,N_19849);
and UO_802 (O_802,N_19992,N_19950);
nand UO_803 (O_803,N_19919,N_19855);
or UO_804 (O_804,N_19986,N_19982);
nor UO_805 (O_805,N_19975,N_19982);
or UO_806 (O_806,N_19888,N_19969);
and UO_807 (O_807,N_19960,N_19843);
nor UO_808 (O_808,N_19980,N_19964);
nor UO_809 (O_809,N_19955,N_19934);
xor UO_810 (O_810,N_19934,N_19981);
xor UO_811 (O_811,N_19870,N_19871);
or UO_812 (O_812,N_19989,N_19964);
and UO_813 (O_813,N_19848,N_19899);
nor UO_814 (O_814,N_19959,N_19944);
or UO_815 (O_815,N_19900,N_19982);
and UO_816 (O_816,N_19950,N_19906);
or UO_817 (O_817,N_19857,N_19972);
nand UO_818 (O_818,N_19890,N_19967);
nor UO_819 (O_819,N_19860,N_19841);
nor UO_820 (O_820,N_19905,N_19842);
nand UO_821 (O_821,N_19860,N_19845);
nor UO_822 (O_822,N_19881,N_19894);
nor UO_823 (O_823,N_19931,N_19853);
xor UO_824 (O_824,N_19926,N_19910);
and UO_825 (O_825,N_19917,N_19879);
and UO_826 (O_826,N_19978,N_19842);
or UO_827 (O_827,N_19986,N_19896);
or UO_828 (O_828,N_19881,N_19927);
and UO_829 (O_829,N_19865,N_19945);
and UO_830 (O_830,N_19900,N_19920);
or UO_831 (O_831,N_19905,N_19957);
nand UO_832 (O_832,N_19920,N_19991);
or UO_833 (O_833,N_19933,N_19997);
xor UO_834 (O_834,N_19970,N_19917);
or UO_835 (O_835,N_19931,N_19877);
and UO_836 (O_836,N_19861,N_19978);
or UO_837 (O_837,N_19870,N_19985);
nor UO_838 (O_838,N_19919,N_19907);
xor UO_839 (O_839,N_19893,N_19999);
xnor UO_840 (O_840,N_19843,N_19966);
nand UO_841 (O_841,N_19897,N_19919);
and UO_842 (O_842,N_19918,N_19842);
nand UO_843 (O_843,N_19937,N_19946);
nor UO_844 (O_844,N_19879,N_19856);
or UO_845 (O_845,N_19863,N_19959);
nand UO_846 (O_846,N_19932,N_19958);
xor UO_847 (O_847,N_19866,N_19891);
and UO_848 (O_848,N_19948,N_19870);
xnor UO_849 (O_849,N_19914,N_19887);
and UO_850 (O_850,N_19867,N_19848);
xnor UO_851 (O_851,N_19877,N_19868);
nand UO_852 (O_852,N_19961,N_19942);
nand UO_853 (O_853,N_19940,N_19854);
nor UO_854 (O_854,N_19879,N_19959);
xnor UO_855 (O_855,N_19972,N_19966);
or UO_856 (O_856,N_19960,N_19891);
and UO_857 (O_857,N_19845,N_19842);
or UO_858 (O_858,N_19858,N_19860);
xnor UO_859 (O_859,N_19981,N_19966);
and UO_860 (O_860,N_19889,N_19945);
and UO_861 (O_861,N_19874,N_19999);
and UO_862 (O_862,N_19875,N_19879);
xor UO_863 (O_863,N_19914,N_19844);
nand UO_864 (O_864,N_19952,N_19904);
nand UO_865 (O_865,N_19958,N_19882);
nor UO_866 (O_866,N_19997,N_19940);
xor UO_867 (O_867,N_19855,N_19891);
nand UO_868 (O_868,N_19938,N_19840);
or UO_869 (O_869,N_19984,N_19975);
nor UO_870 (O_870,N_19887,N_19859);
nor UO_871 (O_871,N_19947,N_19974);
or UO_872 (O_872,N_19907,N_19940);
and UO_873 (O_873,N_19928,N_19949);
xnor UO_874 (O_874,N_19866,N_19847);
or UO_875 (O_875,N_19941,N_19922);
and UO_876 (O_876,N_19904,N_19908);
nor UO_877 (O_877,N_19885,N_19925);
or UO_878 (O_878,N_19935,N_19938);
and UO_879 (O_879,N_19890,N_19904);
nand UO_880 (O_880,N_19953,N_19960);
nand UO_881 (O_881,N_19956,N_19907);
nor UO_882 (O_882,N_19976,N_19869);
xor UO_883 (O_883,N_19929,N_19866);
and UO_884 (O_884,N_19931,N_19908);
xnor UO_885 (O_885,N_19999,N_19922);
nand UO_886 (O_886,N_19908,N_19872);
or UO_887 (O_887,N_19895,N_19914);
nor UO_888 (O_888,N_19982,N_19909);
nor UO_889 (O_889,N_19914,N_19989);
nand UO_890 (O_890,N_19929,N_19969);
nand UO_891 (O_891,N_19966,N_19911);
xnor UO_892 (O_892,N_19904,N_19936);
or UO_893 (O_893,N_19916,N_19988);
nand UO_894 (O_894,N_19860,N_19886);
xor UO_895 (O_895,N_19927,N_19861);
and UO_896 (O_896,N_19866,N_19871);
and UO_897 (O_897,N_19998,N_19845);
and UO_898 (O_898,N_19969,N_19933);
or UO_899 (O_899,N_19986,N_19856);
nor UO_900 (O_900,N_19941,N_19873);
xnor UO_901 (O_901,N_19980,N_19994);
or UO_902 (O_902,N_19923,N_19926);
xor UO_903 (O_903,N_19868,N_19879);
and UO_904 (O_904,N_19975,N_19968);
and UO_905 (O_905,N_19841,N_19954);
and UO_906 (O_906,N_19931,N_19962);
nand UO_907 (O_907,N_19925,N_19936);
nor UO_908 (O_908,N_19886,N_19981);
or UO_909 (O_909,N_19989,N_19906);
and UO_910 (O_910,N_19857,N_19996);
or UO_911 (O_911,N_19920,N_19912);
nand UO_912 (O_912,N_19904,N_19851);
and UO_913 (O_913,N_19984,N_19844);
nor UO_914 (O_914,N_19923,N_19959);
or UO_915 (O_915,N_19841,N_19919);
xnor UO_916 (O_916,N_19875,N_19960);
or UO_917 (O_917,N_19865,N_19860);
or UO_918 (O_918,N_19986,N_19853);
and UO_919 (O_919,N_19991,N_19979);
and UO_920 (O_920,N_19887,N_19846);
nor UO_921 (O_921,N_19864,N_19974);
and UO_922 (O_922,N_19867,N_19915);
nand UO_923 (O_923,N_19861,N_19923);
xor UO_924 (O_924,N_19995,N_19934);
nor UO_925 (O_925,N_19937,N_19960);
or UO_926 (O_926,N_19953,N_19975);
nand UO_927 (O_927,N_19917,N_19965);
or UO_928 (O_928,N_19865,N_19968);
nor UO_929 (O_929,N_19852,N_19906);
nand UO_930 (O_930,N_19968,N_19941);
and UO_931 (O_931,N_19943,N_19974);
nand UO_932 (O_932,N_19851,N_19928);
and UO_933 (O_933,N_19857,N_19861);
nand UO_934 (O_934,N_19946,N_19995);
or UO_935 (O_935,N_19964,N_19855);
nor UO_936 (O_936,N_19920,N_19882);
and UO_937 (O_937,N_19923,N_19884);
or UO_938 (O_938,N_19954,N_19891);
nand UO_939 (O_939,N_19971,N_19896);
nor UO_940 (O_940,N_19938,N_19973);
nor UO_941 (O_941,N_19987,N_19950);
or UO_942 (O_942,N_19873,N_19881);
nand UO_943 (O_943,N_19975,N_19966);
or UO_944 (O_944,N_19963,N_19902);
or UO_945 (O_945,N_19987,N_19896);
or UO_946 (O_946,N_19993,N_19864);
nand UO_947 (O_947,N_19874,N_19889);
nand UO_948 (O_948,N_19904,N_19869);
xor UO_949 (O_949,N_19871,N_19954);
nor UO_950 (O_950,N_19854,N_19871);
nand UO_951 (O_951,N_19962,N_19855);
or UO_952 (O_952,N_19962,N_19979);
xor UO_953 (O_953,N_19968,N_19933);
nand UO_954 (O_954,N_19860,N_19852);
xor UO_955 (O_955,N_19934,N_19884);
xor UO_956 (O_956,N_19840,N_19932);
nor UO_957 (O_957,N_19949,N_19899);
nor UO_958 (O_958,N_19937,N_19996);
nand UO_959 (O_959,N_19877,N_19987);
and UO_960 (O_960,N_19982,N_19976);
or UO_961 (O_961,N_19891,N_19949);
xnor UO_962 (O_962,N_19997,N_19986);
and UO_963 (O_963,N_19880,N_19886);
nor UO_964 (O_964,N_19855,N_19927);
and UO_965 (O_965,N_19993,N_19941);
or UO_966 (O_966,N_19917,N_19860);
xor UO_967 (O_967,N_19960,N_19901);
xor UO_968 (O_968,N_19871,N_19923);
or UO_969 (O_969,N_19842,N_19864);
and UO_970 (O_970,N_19852,N_19920);
nand UO_971 (O_971,N_19937,N_19957);
nand UO_972 (O_972,N_19908,N_19943);
or UO_973 (O_973,N_19999,N_19925);
xnor UO_974 (O_974,N_19896,N_19848);
xnor UO_975 (O_975,N_19931,N_19963);
and UO_976 (O_976,N_19929,N_19863);
nor UO_977 (O_977,N_19904,N_19886);
nand UO_978 (O_978,N_19998,N_19910);
xor UO_979 (O_979,N_19892,N_19898);
xnor UO_980 (O_980,N_19913,N_19845);
and UO_981 (O_981,N_19913,N_19875);
nand UO_982 (O_982,N_19868,N_19921);
nor UO_983 (O_983,N_19883,N_19885);
xor UO_984 (O_984,N_19867,N_19846);
nor UO_985 (O_985,N_19985,N_19908);
xor UO_986 (O_986,N_19893,N_19915);
xor UO_987 (O_987,N_19975,N_19895);
or UO_988 (O_988,N_19865,N_19854);
and UO_989 (O_989,N_19948,N_19917);
or UO_990 (O_990,N_19905,N_19945);
xor UO_991 (O_991,N_19909,N_19989);
or UO_992 (O_992,N_19891,N_19939);
and UO_993 (O_993,N_19997,N_19872);
and UO_994 (O_994,N_19860,N_19981);
or UO_995 (O_995,N_19955,N_19976);
nor UO_996 (O_996,N_19840,N_19943);
nand UO_997 (O_997,N_19878,N_19910);
and UO_998 (O_998,N_19897,N_19980);
or UO_999 (O_999,N_19855,N_19856);
nor UO_1000 (O_1000,N_19999,N_19896);
or UO_1001 (O_1001,N_19984,N_19956);
nand UO_1002 (O_1002,N_19995,N_19972);
nand UO_1003 (O_1003,N_19887,N_19875);
and UO_1004 (O_1004,N_19892,N_19954);
and UO_1005 (O_1005,N_19984,N_19913);
nor UO_1006 (O_1006,N_19948,N_19994);
nand UO_1007 (O_1007,N_19985,N_19881);
nand UO_1008 (O_1008,N_19923,N_19981);
or UO_1009 (O_1009,N_19978,N_19918);
xnor UO_1010 (O_1010,N_19883,N_19897);
nand UO_1011 (O_1011,N_19903,N_19937);
and UO_1012 (O_1012,N_19845,N_19885);
xnor UO_1013 (O_1013,N_19856,N_19971);
and UO_1014 (O_1014,N_19986,N_19908);
nand UO_1015 (O_1015,N_19968,N_19879);
nand UO_1016 (O_1016,N_19936,N_19971);
xor UO_1017 (O_1017,N_19936,N_19865);
and UO_1018 (O_1018,N_19993,N_19860);
or UO_1019 (O_1019,N_19963,N_19966);
xor UO_1020 (O_1020,N_19892,N_19889);
xnor UO_1021 (O_1021,N_19953,N_19865);
nor UO_1022 (O_1022,N_19912,N_19921);
and UO_1023 (O_1023,N_19993,N_19905);
xnor UO_1024 (O_1024,N_19993,N_19871);
xor UO_1025 (O_1025,N_19968,N_19892);
nor UO_1026 (O_1026,N_19880,N_19878);
or UO_1027 (O_1027,N_19935,N_19965);
and UO_1028 (O_1028,N_19934,N_19880);
xor UO_1029 (O_1029,N_19957,N_19879);
nand UO_1030 (O_1030,N_19999,N_19937);
xor UO_1031 (O_1031,N_19998,N_19974);
nand UO_1032 (O_1032,N_19864,N_19892);
nor UO_1033 (O_1033,N_19937,N_19848);
xnor UO_1034 (O_1034,N_19958,N_19919);
or UO_1035 (O_1035,N_19864,N_19858);
nor UO_1036 (O_1036,N_19947,N_19882);
xor UO_1037 (O_1037,N_19883,N_19931);
or UO_1038 (O_1038,N_19941,N_19866);
and UO_1039 (O_1039,N_19857,N_19912);
xnor UO_1040 (O_1040,N_19871,N_19951);
and UO_1041 (O_1041,N_19890,N_19988);
and UO_1042 (O_1042,N_19986,N_19950);
or UO_1043 (O_1043,N_19924,N_19864);
or UO_1044 (O_1044,N_19944,N_19911);
and UO_1045 (O_1045,N_19968,N_19942);
nor UO_1046 (O_1046,N_19864,N_19973);
nor UO_1047 (O_1047,N_19936,N_19909);
nand UO_1048 (O_1048,N_19985,N_19847);
xor UO_1049 (O_1049,N_19996,N_19852);
nand UO_1050 (O_1050,N_19991,N_19970);
or UO_1051 (O_1051,N_19931,N_19850);
or UO_1052 (O_1052,N_19882,N_19916);
and UO_1053 (O_1053,N_19843,N_19898);
and UO_1054 (O_1054,N_19845,N_19930);
nand UO_1055 (O_1055,N_19933,N_19878);
nand UO_1056 (O_1056,N_19864,N_19843);
and UO_1057 (O_1057,N_19846,N_19974);
or UO_1058 (O_1058,N_19887,N_19844);
and UO_1059 (O_1059,N_19848,N_19870);
nor UO_1060 (O_1060,N_19867,N_19925);
and UO_1061 (O_1061,N_19933,N_19956);
xnor UO_1062 (O_1062,N_19904,N_19924);
xor UO_1063 (O_1063,N_19924,N_19944);
nand UO_1064 (O_1064,N_19976,N_19941);
nand UO_1065 (O_1065,N_19895,N_19934);
nand UO_1066 (O_1066,N_19982,N_19979);
nor UO_1067 (O_1067,N_19965,N_19840);
and UO_1068 (O_1068,N_19977,N_19918);
xnor UO_1069 (O_1069,N_19982,N_19952);
or UO_1070 (O_1070,N_19926,N_19906);
and UO_1071 (O_1071,N_19854,N_19894);
and UO_1072 (O_1072,N_19926,N_19888);
nor UO_1073 (O_1073,N_19981,N_19926);
and UO_1074 (O_1074,N_19998,N_19848);
or UO_1075 (O_1075,N_19848,N_19915);
nand UO_1076 (O_1076,N_19943,N_19941);
xnor UO_1077 (O_1077,N_19981,N_19991);
and UO_1078 (O_1078,N_19892,N_19975);
or UO_1079 (O_1079,N_19955,N_19921);
and UO_1080 (O_1080,N_19925,N_19959);
nand UO_1081 (O_1081,N_19989,N_19998);
xnor UO_1082 (O_1082,N_19910,N_19869);
xnor UO_1083 (O_1083,N_19918,N_19961);
xnor UO_1084 (O_1084,N_19848,N_19871);
or UO_1085 (O_1085,N_19853,N_19909);
or UO_1086 (O_1086,N_19978,N_19958);
nor UO_1087 (O_1087,N_19974,N_19848);
nor UO_1088 (O_1088,N_19938,N_19949);
xor UO_1089 (O_1089,N_19876,N_19926);
and UO_1090 (O_1090,N_19976,N_19978);
xor UO_1091 (O_1091,N_19882,N_19942);
nand UO_1092 (O_1092,N_19870,N_19943);
or UO_1093 (O_1093,N_19949,N_19887);
or UO_1094 (O_1094,N_19843,N_19874);
nand UO_1095 (O_1095,N_19851,N_19939);
nand UO_1096 (O_1096,N_19963,N_19945);
and UO_1097 (O_1097,N_19999,N_19882);
and UO_1098 (O_1098,N_19878,N_19943);
nor UO_1099 (O_1099,N_19981,N_19969);
or UO_1100 (O_1100,N_19990,N_19863);
xnor UO_1101 (O_1101,N_19877,N_19873);
xnor UO_1102 (O_1102,N_19933,N_19852);
nand UO_1103 (O_1103,N_19971,N_19920);
or UO_1104 (O_1104,N_19920,N_19904);
and UO_1105 (O_1105,N_19878,N_19883);
nor UO_1106 (O_1106,N_19908,N_19948);
nand UO_1107 (O_1107,N_19849,N_19942);
nand UO_1108 (O_1108,N_19968,N_19910);
nor UO_1109 (O_1109,N_19947,N_19902);
nand UO_1110 (O_1110,N_19975,N_19898);
xnor UO_1111 (O_1111,N_19954,N_19982);
and UO_1112 (O_1112,N_19884,N_19921);
nor UO_1113 (O_1113,N_19846,N_19996);
xor UO_1114 (O_1114,N_19883,N_19867);
xnor UO_1115 (O_1115,N_19942,N_19892);
nand UO_1116 (O_1116,N_19964,N_19927);
nand UO_1117 (O_1117,N_19962,N_19888);
xnor UO_1118 (O_1118,N_19988,N_19901);
or UO_1119 (O_1119,N_19887,N_19843);
nand UO_1120 (O_1120,N_19959,N_19911);
or UO_1121 (O_1121,N_19883,N_19851);
nor UO_1122 (O_1122,N_19979,N_19944);
or UO_1123 (O_1123,N_19928,N_19935);
and UO_1124 (O_1124,N_19925,N_19886);
and UO_1125 (O_1125,N_19843,N_19885);
nand UO_1126 (O_1126,N_19848,N_19890);
and UO_1127 (O_1127,N_19974,N_19923);
xor UO_1128 (O_1128,N_19864,N_19841);
and UO_1129 (O_1129,N_19892,N_19996);
nor UO_1130 (O_1130,N_19980,N_19885);
nor UO_1131 (O_1131,N_19840,N_19940);
or UO_1132 (O_1132,N_19939,N_19933);
xnor UO_1133 (O_1133,N_19886,N_19922);
and UO_1134 (O_1134,N_19923,N_19962);
nor UO_1135 (O_1135,N_19902,N_19916);
xor UO_1136 (O_1136,N_19877,N_19852);
and UO_1137 (O_1137,N_19872,N_19880);
xor UO_1138 (O_1138,N_19866,N_19999);
and UO_1139 (O_1139,N_19877,N_19945);
nor UO_1140 (O_1140,N_19871,N_19880);
nand UO_1141 (O_1141,N_19988,N_19904);
and UO_1142 (O_1142,N_19893,N_19887);
and UO_1143 (O_1143,N_19968,N_19908);
or UO_1144 (O_1144,N_19954,N_19862);
xnor UO_1145 (O_1145,N_19889,N_19964);
or UO_1146 (O_1146,N_19848,N_19970);
xnor UO_1147 (O_1147,N_19914,N_19954);
or UO_1148 (O_1148,N_19931,N_19959);
or UO_1149 (O_1149,N_19858,N_19928);
xor UO_1150 (O_1150,N_19891,N_19972);
and UO_1151 (O_1151,N_19903,N_19967);
or UO_1152 (O_1152,N_19935,N_19937);
and UO_1153 (O_1153,N_19994,N_19892);
or UO_1154 (O_1154,N_19941,N_19916);
nor UO_1155 (O_1155,N_19915,N_19857);
or UO_1156 (O_1156,N_19904,N_19978);
xnor UO_1157 (O_1157,N_19995,N_19936);
nand UO_1158 (O_1158,N_19895,N_19871);
or UO_1159 (O_1159,N_19990,N_19931);
xnor UO_1160 (O_1160,N_19858,N_19865);
xor UO_1161 (O_1161,N_19852,N_19851);
nor UO_1162 (O_1162,N_19951,N_19919);
nor UO_1163 (O_1163,N_19848,N_19863);
nand UO_1164 (O_1164,N_19856,N_19862);
nor UO_1165 (O_1165,N_19961,N_19929);
xor UO_1166 (O_1166,N_19861,N_19887);
nor UO_1167 (O_1167,N_19944,N_19882);
nor UO_1168 (O_1168,N_19926,N_19948);
nand UO_1169 (O_1169,N_19963,N_19848);
or UO_1170 (O_1170,N_19965,N_19968);
xnor UO_1171 (O_1171,N_19936,N_19956);
nor UO_1172 (O_1172,N_19921,N_19928);
nor UO_1173 (O_1173,N_19945,N_19880);
nand UO_1174 (O_1174,N_19960,N_19846);
nand UO_1175 (O_1175,N_19989,N_19927);
and UO_1176 (O_1176,N_19919,N_19896);
nor UO_1177 (O_1177,N_19937,N_19893);
xnor UO_1178 (O_1178,N_19911,N_19855);
nor UO_1179 (O_1179,N_19970,N_19895);
nor UO_1180 (O_1180,N_19998,N_19907);
nand UO_1181 (O_1181,N_19855,N_19863);
and UO_1182 (O_1182,N_19987,N_19903);
xnor UO_1183 (O_1183,N_19874,N_19960);
nor UO_1184 (O_1184,N_19982,N_19849);
nor UO_1185 (O_1185,N_19901,N_19979);
or UO_1186 (O_1186,N_19949,N_19888);
nand UO_1187 (O_1187,N_19854,N_19929);
nand UO_1188 (O_1188,N_19963,N_19878);
nand UO_1189 (O_1189,N_19982,N_19861);
nand UO_1190 (O_1190,N_19855,N_19940);
nand UO_1191 (O_1191,N_19995,N_19953);
xnor UO_1192 (O_1192,N_19952,N_19894);
or UO_1193 (O_1193,N_19892,N_19930);
nor UO_1194 (O_1194,N_19987,N_19955);
and UO_1195 (O_1195,N_19844,N_19880);
nor UO_1196 (O_1196,N_19939,N_19923);
nor UO_1197 (O_1197,N_19997,N_19934);
and UO_1198 (O_1198,N_19861,N_19896);
and UO_1199 (O_1199,N_19872,N_19953);
nor UO_1200 (O_1200,N_19988,N_19853);
or UO_1201 (O_1201,N_19933,N_19917);
and UO_1202 (O_1202,N_19914,N_19845);
or UO_1203 (O_1203,N_19973,N_19888);
xor UO_1204 (O_1204,N_19973,N_19962);
nand UO_1205 (O_1205,N_19870,N_19967);
xnor UO_1206 (O_1206,N_19842,N_19967);
and UO_1207 (O_1207,N_19974,N_19853);
nand UO_1208 (O_1208,N_19857,N_19891);
or UO_1209 (O_1209,N_19844,N_19889);
xor UO_1210 (O_1210,N_19957,N_19875);
nand UO_1211 (O_1211,N_19867,N_19902);
or UO_1212 (O_1212,N_19924,N_19920);
or UO_1213 (O_1213,N_19928,N_19863);
or UO_1214 (O_1214,N_19900,N_19965);
nand UO_1215 (O_1215,N_19926,N_19930);
nand UO_1216 (O_1216,N_19984,N_19845);
xor UO_1217 (O_1217,N_19866,N_19860);
and UO_1218 (O_1218,N_19896,N_19997);
xor UO_1219 (O_1219,N_19866,N_19945);
and UO_1220 (O_1220,N_19963,N_19979);
xor UO_1221 (O_1221,N_19925,N_19847);
xnor UO_1222 (O_1222,N_19986,N_19924);
and UO_1223 (O_1223,N_19905,N_19971);
nor UO_1224 (O_1224,N_19841,N_19998);
nor UO_1225 (O_1225,N_19860,N_19938);
xnor UO_1226 (O_1226,N_19924,N_19893);
xor UO_1227 (O_1227,N_19932,N_19881);
or UO_1228 (O_1228,N_19977,N_19948);
nor UO_1229 (O_1229,N_19859,N_19989);
or UO_1230 (O_1230,N_19877,N_19953);
and UO_1231 (O_1231,N_19968,N_19930);
and UO_1232 (O_1232,N_19959,N_19982);
nand UO_1233 (O_1233,N_19936,N_19874);
nor UO_1234 (O_1234,N_19841,N_19916);
nor UO_1235 (O_1235,N_19891,N_19876);
nand UO_1236 (O_1236,N_19922,N_19924);
xnor UO_1237 (O_1237,N_19928,N_19913);
or UO_1238 (O_1238,N_19907,N_19946);
or UO_1239 (O_1239,N_19899,N_19938);
and UO_1240 (O_1240,N_19969,N_19879);
and UO_1241 (O_1241,N_19977,N_19844);
xor UO_1242 (O_1242,N_19930,N_19941);
or UO_1243 (O_1243,N_19967,N_19919);
nor UO_1244 (O_1244,N_19882,N_19881);
and UO_1245 (O_1245,N_19875,N_19840);
xor UO_1246 (O_1246,N_19919,N_19875);
xor UO_1247 (O_1247,N_19978,N_19974);
or UO_1248 (O_1248,N_19968,N_19849);
and UO_1249 (O_1249,N_19955,N_19887);
nor UO_1250 (O_1250,N_19945,N_19944);
nand UO_1251 (O_1251,N_19988,N_19970);
nor UO_1252 (O_1252,N_19934,N_19871);
nor UO_1253 (O_1253,N_19953,N_19989);
xor UO_1254 (O_1254,N_19985,N_19895);
and UO_1255 (O_1255,N_19988,N_19939);
xor UO_1256 (O_1256,N_19873,N_19958);
xnor UO_1257 (O_1257,N_19914,N_19935);
or UO_1258 (O_1258,N_19992,N_19840);
xnor UO_1259 (O_1259,N_19882,N_19912);
and UO_1260 (O_1260,N_19874,N_19844);
nor UO_1261 (O_1261,N_19868,N_19934);
nand UO_1262 (O_1262,N_19843,N_19870);
nand UO_1263 (O_1263,N_19936,N_19948);
xnor UO_1264 (O_1264,N_19915,N_19872);
or UO_1265 (O_1265,N_19862,N_19847);
nand UO_1266 (O_1266,N_19980,N_19922);
or UO_1267 (O_1267,N_19940,N_19991);
or UO_1268 (O_1268,N_19935,N_19882);
xor UO_1269 (O_1269,N_19908,N_19859);
nand UO_1270 (O_1270,N_19961,N_19908);
or UO_1271 (O_1271,N_19954,N_19959);
nor UO_1272 (O_1272,N_19949,N_19971);
xor UO_1273 (O_1273,N_19940,N_19944);
xnor UO_1274 (O_1274,N_19938,N_19848);
nor UO_1275 (O_1275,N_19949,N_19871);
nand UO_1276 (O_1276,N_19876,N_19849);
xor UO_1277 (O_1277,N_19981,N_19976);
xor UO_1278 (O_1278,N_19853,N_19946);
or UO_1279 (O_1279,N_19898,N_19844);
nand UO_1280 (O_1280,N_19902,N_19866);
nand UO_1281 (O_1281,N_19997,N_19873);
xnor UO_1282 (O_1282,N_19941,N_19957);
nand UO_1283 (O_1283,N_19983,N_19854);
xor UO_1284 (O_1284,N_19966,N_19901);
nor UO_1285 (O_1285,N_19950,N_19977);
or UO_1286 (O_1286,N_19927,N_19884);
and UO_1287 (O_1287,N_19972,N_19854);
xnor UO_1288 (O_1288,N_19900,N_19877);
xor UO_1289 (O_1289,N_19987,N_19862);
xor UO_1290 (O_1290,N_19841,N_19888);
nor UO_1291 (O_1291,N_19876,N_19952);
and UO_1292 (O_1292,N_19901,N_19902);
nor UO_1293 (O_1293,N_19951,N_19967);
xor UO_1294 (O_1294,N_19999,N_19998);
or UO_1295 (O_1295,N_19967,N_19871);
and UO_1296 (O_1296,N_19914,N_19966);
or UO_1297 (O_1297,N_19976,N_19876);
xor UO_1298 (O_1298,N_19938,N_19914);
nand UO_1299 (O_1299,N_19957,N_19891);
xor UO_1300 (O_1300,N_19892,N_19977);
xor UO_1301 (O_1301,N_19982,N_19899);
xor UO_1302 (O_1302,N_19921,N_19873);
nand UO_1303 (O_1303,N_19937,N_19928);
nand UO_1304 (O_1304,N_19876,N_19974);
nor UO_1305 (O_1305,N_19857,N_19870);
xnor UO_1306 (O_1306,N_19893,N_19846);
nand UO_1307 (O_1307,N_19848,N_19994);
and UO_1308 (O_1308,N_19989,N_19893);
or UO_1309 (O_1309,N_19843,N_19881);
nand UO_1310 (O_1310,N_19874,N_19917);
nand UO_1311 (O_1311,N_19944,N_19896);
nand UO_1312 (O_1312,N_19931,N_19956);
xnor UO_1313 (O_1313,N_19955,N_19945);
xnor UO_1314 (O_1314,N_19933,N_19991);
nor UO_1315 (O_1315,N_19855,N_19993);
or UO_1316 (O_1316,N_19840,N_19865);
or UO_1317 (O_1317,N_19863,N_19886);
xor UO_1318 (O_1318,N_19992,N_19943);
nor UO_1319 (O_1319,N_19919,N_19916);
and UO_1320 (O_1320,N_19908,N_19921);
or UO_1321 (O_1321,N_19950,N_19879);
or UO_1322 (O_1322,N_19881,N_19984);
or UO_1323 (O_1323,N_19992,N_19881);
or UO_1324 (O_1324,N_19918,N_19932);
and UO_1325 (O_1325,N_19906,N_19938);
or UO_1326 (O_1326,N_19893,N_19964);
or UO_1327 (O_1327,N_19867,N_19955);
nor UO_1328 (O_1328,N_19854,N_19903);
xnor UO_1329 (O_1329,N_19892,N_19911);
or UO_1330 (O_1330,N_19935,N_19865);
or UO_1331 (O_1331,N_19976,N_19889);
xnor UO_1332 (O_1332,N_19886,N_19875);
and UO_1333 (O_1333,N_19941,N_19856);
and UO_1334 (O_1334,N_19866,N_19993);
nand UO_1335 (O_1335,N_19943,N_19926);
nand UO_1336 (O_1336,N_19992,N_19996);
nand UO_1337 (O_1337,N_19948,N_19863);
or UO_1338 (O_1338,N_19855,N_19989);
xor UO_1339 (O_1339,N_19870,N_19962);
nand UO_1340 (O_1340,N_19848,N_19892);
or UO_1341 (O_1341,N_19927,N_19842);
xor UO_1342 (O_1342,N_19999,N_19990);
nand UO_1343 (O_1343,N_19957,N_19919);
nor UO_1344 (O_1344,N_19937,N_19849);
xnor UO_1345 (O_1345,N_19875,N_19963);
nor UO_1346 (O_1346,N_19850,N_19897);
xor UO_1347 (O_1347,N_19844,N_19909);
and UO_1348 (O_1348,N_19968,N_19964);
and UO_1349 (O_1349,N_19978,N_19871);
and UO_1350 (O_1350,N_19930,N_19916);
nor UO_1351 (O_1351,N_19985,N_19866);
xor UO_1352 (O_1352,N_19930,N_19955);
nor UO_1353 (O_1353,N_19934,N_19958);
nand UO_1354 (O_1354,N_19935,N_19962);
or UO_1355 (O_1355,N_19841,N_19878);
or UO_1356 (O_1356,N_19859,N_19995);
nand UO_1357 (O_1357,N_19978,N_19959);
nor UO_1358 (O_1358,N_19852,N_19917);
xnor UO_1359 (O_1359,N_19957,N_19855);
xor UO_1360 (O_1360,N_19952,N_19879);
xor UO_1361 (O_1361,N_19945,N_19926);
xnor UO_1362 (O_1362,N_19866,N_19961);
and UO_1363 (O_1363,N_19901,N_19916);
and UO_1364 (O_1364,N_19918,N_19897);
nor UO_1365 (O_1365,N_19953,N_19994);
and UO_1366 (O_1366,N_19933,N_19858);
xnor UO_1367 (O_1367,N_19932,N_19968);
or UO_1368 (O_1368,N_19942,N_19873);
xnor UO_1369 (O_1369,N_19983,N_19946);
xnor UO_1370 (O_1370,N_19956,N_19848);
nor UO_1371 (O_1371,N_19846,N_19847);
or UO_1372 (O_1372,N_19840,N_19854);
nor UO_1373 (O_1373,N_19929,N_19953);
xor UO_1374 (O_1374,N_19854,N_19998);
xor UO_1375 (O_1375,N_19923,N_19937);
xnor UO_1376 (O_1376,N_19844,N_19875);
or UO_1377 (O_1377,N_19925,N_19994);
nand UO_1378 (O_1378,N_19995,N_19870);
xor UO_1379 (O_1379,N_19921,N_19897);
xor UO_1380 (O_1380,N_19890,N_19856);
nand UO_1381 (O_1381,N_19870,N_19924);
and UO_1382 (O_1382,N_19944,N_19842);
nor UO_1383 (O_1383,N_19934,N_19935);
or UO_1384 (O_1384,N_19886,N_19864);
and UO_1385 (O_1385,N_19921,N_19980);
nand UO_1386 (O_1386,N_19962,N_19852);
nor UO_1387 (O_1387,N_19947,N_19905);
or UO_1388 (O_1388,N_19904,N_19949);
nor UO_1389 (O_1389,N_19965,N_19980);
nor UO_1390 (O_1390,N_19899,N_19971);
nand UO_1391 (O_1391,N_19887,N_19910);
nand UO_1392 (O_1392,N_19867,N_19970);
nor UO_1393 (O_1393,N_19983,N_19998);
or UO_1394 (O_1394,N_19952,N_19993);
xnor UO_1395 (O_1395,N_19866,N_19964);
xor UO_1396 (O_1396,N_19887,N_19975);
nand UO_1397 (O_1397,N_19851,N_19985);
nand UO_1398 (O_1398,N_19958,N_19974);
xor UO_1399 (O_1399,N_19888,N_19883);
and UO_1400 (O_1400,N_19856,N_19884);
xor UO_1401 (O_1401,N_19926,N_19886);
nor UO_1402 (O_1402,N_19927,N_19849);
xor UO_1403 (O_1403,N_19992,N_19949);
or UO_1404 (O_1404,N_19908,N_19895);
and UO_1405 (O_1405,N_19944,N_19928);
nor UO_1406 (O_1406,N_19907,N_19930);
nor UO_1407 (O_1407,N_19963,N_19862);
or UO_1408 (O_1408,N_19846,N_19924);
nand UO_1409 (O_1409,N_19941,N_19901);
and UO_1410 (O_1410,N_19908,N_19897);
xnor UO_1411 (O_1411,N_19977,N_19842);
and UO_1412 (O_1412,N_19976,N_19888);
nand UO_1413 (O_1413,N_19850,N_19952);
and UO_1414 (O_1414,N_19857,N_19918);
nand UO_1415 (O_1415,N_19873,N_19870);
nor UO_1416 (O_1416,N_19952,N_19957);
xor UO_1417 (O_1417,N_19968,N_19898);
or UO_1418 (O_1418,N_19890,N_19912);
nand UO_1419 (O_1419,N_19869,N_19989);
or UO_1420 (O_1420,N_19871,N_19867);
nor UO_1421 (O_1421,N_19999,N_19873);
or UO_1422 (O_1422,N_19915,N_19976);
nand UO_1423 (O_1423,N_19902,N_19974);
or UO_1424 (O_1424,N_19996,N_19880);
or UO_1425 (O_1425,N_19898,N_19907);
nand UO_1426 (O_1426,N_19869,N_19971);
xnor UO_1427 (O_1427,N_19941,N_19893);
or UO_1428 (O_1428,N_19840,N_19889);
and UO_1429 (O_1429,N_19971,N_19907);
nor UO_1430 (O_1430,N_19859,N_19889);
xor UO_1431 (O_1431,N_19981,N_19899);
or UO_1432 (O_1432,N_19886,N_19994);
nor UO_1433 (O_1433,N_19989,N_19897);
nand UO_1434 (O_1434,N_19849,N_19961);
xor UO_1435 (O_1435,N_19993,N_19937);
nor UO_1436 (O_1436,N_19931,N_19885);
nand UO_1437 (O_1437,N_19987,N_19911);
or UO_1438 (O_1438,N_19880,N_19972);
or UO_1439 (O_1439,N_19978,N_19840);
nor UO_1440 (O_1440,N_19877,N_19968);
nor UO_1441 (O_1441,N_19881,N_19867);
nor UO_1442 (O_1442,N_19865,N_19960);
and UO_1443 (O_1443,N_19995,N_19947);
xor UO_1444 (O_1444,N_19846,N_19909);
or UO_1445 (O_1445,N_19961,N_19920);
xor UO_1446 (O_1446,N_19938,N_19970);
xnor UO_1447 (O_1447,N_19922,N_19947);
nand UO_1448 (O_1448,N_19849,N_19953);
xnor UO_1449 (O_1449,N_19928,N_19853);
xnor UO_1450 (O_1450,N_19943,N_19905);
xnor UO_1451 (O_1451,N_19969,N_19880);
xnor UO_1452 (O_1452,N_19992,N_19967);
nand UO_1453 (O_1453,N_19856,N_19893);
nor UO_1454 (O_1454,N_19960,N_19961);
and UO_1455 (O_1455,N_19856,N_19885);
or UO_1456 (O_1456,N_19841,N_19905);
nor UO_1457 (O_1457,N_19869,N_19895);
xor UO_1458 (O_1458,N_19917,N_19975);
or UO_1459 (O_1459,N_19900,N_19985);
nor UO_1460 (O_1460,N_19897,N_19928);
nand UO_1461 (O_1461,N_19860,N_19912);
xor UO_1462 (O_1462,N_19889,N_19933);
nand UO_1463 (O_1463,N_19938,N_19930);
nor UO_1464 (O_1464,N_19880,N_19951);
nor UO_1465 (O_1465,N_19973,N_19852);
xor UO_1466 (O_1466,N_19995,N_19889);
nor UO_1467 (O_1467,N_19975,N_19848);
and UO_1468 (O_1468,N_19996,N_19858);
nor UO_1469 (O_1469,N_19864,N_19921);
and UO_1470 (O_1470,N_19858,N_19903);
or UO_1471 (O_1471,N_19998,N_19946);
and UO_1472 (O_1472,N_19887,N_19941);
xnor UO_1473 (O_1473,N_19906,N_19943);
or UO_1474 (O_1474,N_19907,N_19963);
or UO_1475 (O_1475,N_19914,N_19970);
or UO_1476 (O_1476,N_19878,N_19971);
nand UO_1477 (O_1477,N_19859,N_19842);
xnor UO_1478 (O_1478,N_19918,N_19975);
xor UO_1479 (O_1479,N_19967,N_19850);
nand UO_1480 (O_1480,N_19998,N_19880);
xor UO_1481 (O_1481,N_19886,N_19976);
nor UO_1482 (O_1482,N_19975,N_19880);
or UO_1483 (O_1483,N_19891,N_19956);
and UO_1484 (O_1484,N_19915,N_19980);
and UO_1485 (O_1485,N_19978,N_19856);
nand UO_1486 (O_1486,N_19923,N_19996);
nand UO_1487 (O_1487,N_19979,N_19846);
nand UO_1488 (O_1488,N_19870,N_19919);
nand UO_1489 (O_1489,N_19932,N_19930);
xor UO_1490 (O_1490,N_19902,N_19875);
nand UO_1491 (O_1491,N_19974,N_19954);
xor UO_1492 (O_1492,N_19881,N_19883);
and UO_1493 (O_1493,N_19995,N_19893);
nand UO_1494 (O_1494,N_19924,N_19890);
nand UO_1495 (O_1495,N_19950,N_19860);
xor UO_1496 (O_1496,N_19954,N_19899);
nand UO_1497 (O_1497,N_19952,N_19856);
nand UO_1498 (O_1498,N_19942,N_19936);
and UO_1499 (O_1499,N_19869,N_19859);
nand UO_1500 (O_1500,N_19883,N_19866);
nor UO_1501 (O_1501,N_19875,N_19855);
nand UO_1502 (O_1502,N_19918,N_19983);
or UO_1503 (O_1503,N_19957,N_19951);
xnor UO_1504 (O_1504,N_19989,N_19885);
nand UO_1505 (O_1505,N_19908,N_19864);
and UO_1506 (O_1506,N_19902,N_19995);
nand UO_1507 (O_1507,N_19991,N_19912);
xnor UO_1508 (O_1508,N_19952,N_19926);
nand UO_1509 (O_1509,N_19851,N_19927);
nor UO_1510 (O_1510,N_19885,N_19983);
nand UO_1511 (O_1511,N_19937,N_19845);
nor UO_1512 (O_1512,N_19895,N_19875);
nand UO_1513 (O_1513,N_19896,N_19983);
xnor UO_1514 (O_1514,N_19926,N_19957);
or UO_1515 (O_1515,N_19852,N_19947);
or UO_1516 (O_1516,N_19888,N_19893);
xnor UO_1517 (O_1517,N_19990,N_19849);
or UO_1518 (O_1518,N_19875,N_19927);
or UO_1519 (O_1519,N_19898,N_19928);
nor UO_1520 (O_1520,N_19888,N_19992);
nand UO_1521 (O_1521,N_19987,N_19971);
xor UO_1522 (O_1522,N_19928,N_19950);
nand UO_1523 (O_1523,N_19963,N_19845);
xor UO_1524 (O_1524,N_19953,N_19874);
nor UO_1525 (O_1525,N_19891,N_19868);
or UO_1526 (O_1526,N_19999,N_19915);
nor UO_1527 (O_1527,N_19934,N_19989);
xor UO_1528 (O_1528,N_19914,N_19996);
or UO_1529 (O_1529,N_19979,N_19964);
or UO_1530 (O_1530,N_19863,N_19898);
or UO_1531 (O_1531,N_19874,N_19890);
nor UO_1532 (O_1532,N_19895,N_19939);
nand UO_1533 (O_1533,N_19948,N_19887);
nand UO_1534 (O_1534,N_19933,N_19918);
xor UO_1535 (O_1535,N_19995,N_19927);
xor UO_1536 (O_1536,N_19853,N_19994);
nor UO_1537 (O_1537,N_19853,N_19958);
nor UO_1538 (O_1538,N_19959,N_19938);
and UO_1539 (O_1539,N_19905,N_19868);
nor UO_1540 (O_1540,N_19937,N_19841);
nor UO_1541 (O_1541,N_19887,N_19943);
xor UO_1542 (O_1542,N_19871,N_19863);
nand UO_1543 (O_1543,N_19990,N_19859);
xor UO_1544 (O_1544,N_19981,N_19936);
nor UO_1545 (O_1545,N_19977,N_19941);
or UO_1546 (O_1546,N_19949,N_19856);
nand UO_1547 (O_1547,N_19884,N_19998);
nand UO_1548 (O_1548,N_19907,N_19853);
or UO_1549 (O_1549,N_19994,N_19943);
xnor UO_1550 (O_1550,N_19972,N_19874);
nor UO_1551 (O_1551,N_19925,N_19840);
nor UO_1552 (O_1552,N_19928,N_19857);
nor UO_1553 (O_1553,N_19892,N_19974);
nand UO_1554 (O_1554,N_19861,N_19960);
and UO_1555 (O_1555,N_19915,N_19928);
and UO_1556 (O_1556,N_19879,N_19899);
or UO_1557 (O_1557,N_19928,N_19994);
nand UO_1558 (O_1558,N_19961,N_19972);
nor UO_1559 (O_1559,N_19993,N_19934);
nand UO_1560 (O_1560,N_19945,N_19962);
and UO_1561 (O_1561,N_19995,N_19923);
xor UO_1562 (O_1562,N_19931,N_19900);
nor UO_1563 (O_1563,N_19874,N_19945);
xor UO_1564 (O_1564,N_19913,N_19927);
nor UO_1565 (O_1565,N_19845,N_19989);
nor UO_1566 (O_1566,N_19964,N_19899);
or UO_1567 (O_1567,N_19954,N_19958);
or UO_1568 (O_1568,N_19962,N_19910);
and UO_1569 (O_1569,N_19937,N_19869);
nand UO_1570 (O_1570,N_19935,N_19939);
xor UO_1571 (O_1571,N_19912,N_19889);
xor UO_1572 (O_1572,N_19873,N_19900);
nor UO_1573 (O_1573,N_19889,N_19899);
or UO_1574 (O_1574,N_19936,N_19868);
nand UO_1575 (O_1575,N_19882,N_19979);
or UO_1576 (O_1576,N_19850,N_19971);
xor UO_1577 (O_1577,N_19977,N_19865);
or UO_1578 (O_1578,N_19847,N_19996);
nor UO_1579 (O_1579,N_19955,N_19908);
nor UO_1580 (O_1580,N_19873,N_19862);
nor UO_1581 (O_1581,N_19994,N_19956);
nor UO_1582 (O_1582,N_19942,N_19978);
nand UO_1583 (O_1583,N_19940,N_19857);
nand UO_1584 (O_1584,N_19943,N_19952);
xor UO_1585 (O_1585,N_19880,N_19985);
and UO_1586 (O_1586,N_19934,N_19844);
or UO_1587 (O_1587,N_19894,N_19966);
nand UO_1588 (O_1588,N_19938,N_19849);
xnor UO_1589 (O_1589,N_19936,N_19882);
nor UO_1590 (O_1590,N_19989,N_19842);
nand UO_1591 (O_1591,N_19940,N_19871);
nor UO_1592 (O_1592,N_19944,N_19999);
nor UO_1593 (O_1593,N_19945,N_19876);
nand UO_1594 (O_1594,N_19851,N_19991);
nor UO_1595 (O_1595,N_19886,N_19987);
xnor UO_1596 (O_1596,N_19850,N_19868);
or UO_1597 (O_1597,N_19874,N_19869);
or UO_1598 (O_1598,N_19946,N_19958);
nand UO_1599 (O_1599,N_19973,N_19957);
nand UO_1600 (O_1600,N_19869,N_19981);
nor UO_1601 (O_1601,N_19998,N_19870);
or UO_1602 (O_1602,N_19979,N_19942);
xnor UO_1603 (O_1603,N_19912,N_19866);
nor UO_1604 (O_1604,N_19859,N_19997);
nand UO_1605 (O_1605,N_19888,N_19860);
or UO_1606 (O_1606,N_19878,N_19990);
nor UO_1607 (O_1607,N_19893,N_19951);
xnor UO_1608 (O_1608,N_19894,N_19973);
or UO_1609 (O_1609,N_19964,N_19879);
nor UO_1610 (O_1610,N_19893,N_19913);
nor UO_1611 (O_1611,N_19892,N_19857);
or UO_1612 (O_1612,N_19998,N_19840);
xnor UO_1613 (O_1613,N_19867,N_19987);
nor UO_1614 (O_1614,N_19860,N_19951);
nand UO_1615 (O_1615,N_19843,N_19951);
nor UO_1616 (O_1616,N_19964,N_19844);
and UO_1617 (O_1617,N_19937,N_19856);
nor UO_1618 (O_1618,N_19981,N_19911);
xnor UO_1619 (O_1619,N_19917,N_19927);
and UO_1620 (O_1620,N_19908,N_19995);
nand UO_1621 (O_1621,N_19844,N_19938);
nand UO_1622 (O_1622,N_19855,N_19920);
or UO_1623 (O_1623,N_19877,N_19925);
and UO_1624 (O_1624,N_19892,N_19956);
nor UO_1625 (O_1625,N_19993,N_19886);
or UO_1626 (O_1626,N_19879,N_19843);
or UO_1627 (O_1627,N_19945,N_19922);
or UO_1628 (O_1628,N_19866,N_19859);
nor UO_1629 (O_1629,N_19898,N_19937);
xor UO_1630 (O_1630,N_19857,N_19845);
or UO_1631 (O_1631,N_19998,N_19908);
nor UO_1632 (O_1632,N_19945,N_19992);
or UO_1633 (O_1633,N_19916,N_19870);
nor UO_1634 (O_1634,N_19998,N_19901);
xor UO_1635 (O_1635,N_19869,N_19887);
nand UO_1636 (O_1636,N_19869,N_19915);
xnor UO_1637 (O_1637,N_19979,N_19960);
and UO_1638 (O_1638,N_19988,N_19866);
or UO_1639 (O_1639,N_19955,N_19863);
or UO_1640 (O_1640,N_19990,N_19961);
xnor UO_1641 (O_1641,N_19980,N_19862);
or UO_1642 (O_1642,N_19987,N_19985);
xnor UO_1643 (O_1643,N_19850,N_19955);
xnor UO_1644 (O_1644,N_19946,N_19940);
nor UO_1645 (O_1645,N_19846,N_19967);
or UO_1646 (O_1646,N_19916,N_19978);
and UO_1647 (O_1647,N_19856,N_19914);
and UO_1648 (O_1648,N_19942,N_19996);
or UO_1649 (O_1649,N_19841,N_19914);
nor UO_1650 (O_1650,N_19961,N_19985);
and UO_1651 (O_1651,N_19955,N_19852);
and UO_1652 (O_1652,N_19863,N_19894);
xor UO_1653 (O_1653,N_19875,N_19937);
xnor UO_1654 (O_1654,N_19950,N_19975);
nand UO_1655 (O_1655,N_19863,N_19976);
and UO_1656 (O_1656,N_19890,N_19914);
nand UO_1657 (O_1657,N_19903,N_19939);
xor UO_1658 (O_1658,N_19866,N_19980);
and UO_1659 (O_1659,N_19841,N_19893);
nor UO_1660 (O_1660,N_19922,N_19969);
xor UO_1661 (O_1661,N_19976,N_19853);
nor UO_1662 (O_1662,N_19874,N_19954);
and UO_1663 (O_1663,N_19991,N_19843);
nor UO_1664 (O_1664,N_19891,N_19959);
and UO_1665 (O_1665,N_19856,N_19954);
nand UO_1666 (O_1666,N_19927,N_19949);
and UO_1667 (O_1667,N_19997,N_19954);
or UO_1668 (O_1668,N_19966,N_19991);
xnor UO_1669 (O_1669,N_19883,N_19880);
nor UO_1670 (O_1670,N_19990,N_19841);
or UO_1671 (O_1671,N_19942,N_19884);
or UO_1672 (O_1672,N_19848,N_19921);
nor UO_1673 (O_1673,N_19860,N_19998);
and UO_1674 (O_1674,N_19870,N_19896);
xnor UO_1675 (O_1675,N_19990,N_19881);
or UO_1676 (O_1676,N_19879,N_19918);
nand UO_1677 (O_1677,N_19941,N_19907);
xor UO_1678 (O_1678,N_19885,N_19991);
or UO_1679 (O_1679,N_19928,N_19875);
nand UO_1680 (O_1680,N_19895,N_19938);
or UO_1681 (O_1681,N_19983,N_19994);
or UO_1682 (O_1682,N_19951,N_19942);
xor UO_1683 (O_1683,N_19990,N_19970);
and UO_1684 (O_1684,N_19928,N_19922);
nand UO_1685 (O_1685,N_19944,N_19867);
xor UO_1686 (O_1686,N_19868,N_19872);
xor UO_1687 (O_1687,N_19954,N_19976);
nand UO_1688 (O_1688,N_19972,N_19859);
nand UO_1689 (O_1689,N_19898,N_19902);
or UO_1690 (O_1690,N_19977,N_19859);
xor UO_1691 (O_1691,N_19842,N_19983);
xor UO_1692 (O_1692,N_19948,N_19861);
xnor UO_1693 (O_1693,N_19993,N_19960);
nor UO_1694 (O_1694,N_19877,N_19844);
xor UO_1695 (O_1695,N_19937,N_19978);
nor UO_1696 (O_1696,N_19995,N_19985);
and UO_1697 (O_1697,N_19977,N_19917);
or UO_1698 (O_1698,N_19869,N_19896);
nor UO_1699 (O_1699,N_19949,N_19851);
xnor UO_1700 (O_1700,N_19883,N_19993);
nor UO_1701 (O_1701,N_19938,N_19919);
nand UO_1702 (O_1702,N_19969,N_19989);
nand UO_1703 (O_1703,N_19877,N_19889);
nand UO_1704 (O_1704,N_19845,N_19854);
or UO_1705 (O_1705,N_19890,N_19957);
nand UO_1706 (O_1706,N_19972,N_19875);
xor UO_1707 (O_1707,N_19942,N_19865);
and UO_1708 (O_1708,N_19963,N_19971);
and UO_1709 (O_1709,N_19912,N_19949);
nor UO_1710 (O_1710,N_19912,N_19923);
xor UO_1711 (O_1711,N_19994,N_19883);
and UO_1712 (O_1712,N_19948,N_19843);
xnor UO_1713 (O_1713,N_19867,N_19923);
nand UO_1714 (O_1714,N_19881,N_19910);
nor UO_1715 (O_1715,N_19899,N_19999);
or UO_1716 (O_1716,N_19967,N_19901);
and UO_1717 (O_1717,N_19966,N_19968);
xnor UO_1718 (O_1718,N_19841,N_19984);
and UO_1719 (O_1719,N_19944,N_19853);
nor UO_1720 (O_1720,N_19869,N_19920);
nand UO_1721 (O_1721,N_19984,N_19991);
and UO_1722 (O_1722,N_19900,N_19844);
nand UO_1723 (O_1723,N_19903,N_19976);
and UO_1724 (O_1724,N_19873,N_19938);
or UO_1725 (O_1725,N_19901,N_19963);
xnor UO_1726 (O_1726,N_19898,N_19960);
and UO_1727 (O_1727,N_19983,N_19861);
or UO_1728 (O_1728,N_19867,N_19940);
or UO_1729 (O_1729,N_19892,N_19955);
nor UO_1730 (O_1730,N_19899,N_19893);
or UO_1731 (O_1731,N_19983,N_19990);
xor UO_1732 (O_1732,N_19905,N_19891);
xnor UO_1733 (O_1733,N_19893,N_19966);
nand UO_1734 (O_1734,N_19914,N_19870);
nand UO_1735 (O_1735,N_19864,N_19987);
and UO_1736 (O_1736,N_19891,N_19841);
nor UO_1737 (O_1737,N_19987,N_19850);
xnor UO_1738 (O_1738,N_19933,N_19885);
nand UO_1739 (O_1739,N_19974,N_19944);
xnor UO_1740 (O_1740,N_19915,N_19937);
or UO_1741 (O_1741,N_19963,N_19926);
nand UO_1742 (O_1742,N_19963,N_19934);
nand UO_1743 (O_1743,N_19943,N_19955);
nand UO_1744 (O_1744,N_19895,N_19992);
and UO_1745 (O_1745,N_19863,N_19860);
and UO_1746 (O_1746,N_19865,N_19940);
nand UO_1747 (O_1747,N_19891,N_19976);
nand UO_1748 (O_1748,N_19955,N_19952);
nand UO_1749 (O_1749,N_19843,N_19953);
and UO_1750 (O_1750,N_19927,N_19877);
or UO_1751 (O_1751,N_19883,N_19911);
or UO_1752 (O_1752,N_19859,N_19939);
xnor UO_1753 (O_1753,N_19990,N_19875);
xnor UO_1754 (O_1754,N_19892,N_19900);
and UO_1755 (O_1755,N_19987,N_19895);
and UO_1756 (O_1756,N_19937,N_19897);
nand UO_1757 (O_1757,N_19938,N_19993);
or UO_1758 (O_1758,N_19988,N_19899);
nor UO_1759 (O_1759,N_19963,N_19990);
nor UO_1760 (O_1760,N_19934,N_19888);
and UO_1761 (O_1761,N_19842,N_19973);
nand UO_1762 (O_1762,N_19874,N_19955);
xnor UO_1763 (O_1763,N_19881,N_19922);
nand UO_1764 (O_1764,N_19905,N_19944);
nand UO_1765 (O_1765,N_19876,N_19912);
or UO_1766 (O_1766,N_19981,N_19907);
nor UO_1767 (O_1767,N_19843,N_19954);
xor UO_1768 (O_1768,N_19943,N_19849);
or UO_1769 (O_1769,N_19914,N_19977);
nor UO_1770 (O_1770,N_19905,N_19924);
nand UO_1771 (O_1771,N_19940,N_19994);
nor UO_1772 (O_1772,N_19958,N_19843);
and UO_1773 (O_1773,N_19897,N_19933);
and UO_1774 (O_1774,N_19970,N_19982);
or UO_1775 (O_1775,N_19867,N_19869);
xor UO_1776 (O_1776,N_19910,N_19921);
nor UO_1777 (O_1777,N_19897,N_19982);
nor UO_1778 (O_1778,N_19841,N_19938);
and UO_1779 (O_1779,N_19974,N_19890);
nor UO_1780 (O_1780,N_19975,N_19926);
or UO_1781 (O_1781,N_19985,N_19860);
and UO_1782 (O_1782,N_19901,N_19876);
or UO_1783 (O_1783,N_19995,N_19905);
xor UO_1784 (O_1784,N_19968,N_19862);
nor UO_1785 (O_1785,N_19967,N_19876);
nor UO_1786 (O_1786,N_19915,N_19905);
and UO_1787 (O_1787,N_19888,N_19957);
nand UO_1788 (O_1788,N_19932,N_19926);
xnor UO_1789 (O_1789,N_19951,N_19873);
and UO_1790 (O_1790,N_19911,N_19936);
nand UO_1791 (O_1791,N_19870,N_19941);
and UO_1792 (O_1792,N_19994,N_19921);
nor UO_1793 (O_1793,N_19860,N_19921);
nor UO_1794 (O_1794,N_19841,N_19986);
and UO_1795 (O_1795,N_19970,N_19946);
or UO_1796 (O_1796,N_19870,N_19986);
nor UO_1797 (O_1797,N_19991,N_19916);
or UO_1798 (O_1798,N_19925,N_19856);
xnor UO_1799 (O_1799,N_19955,N_19982);
xnor UO_1800 (O_1800,N_19968,N_19885);
nor UO_1801 (O_1801,N_19926,N_19990);
nand UO_1802 (O_1802,N_19854,N_19938);
nor UO_1803 (O_1803,N_19986,N_19918);
or UO_1804 (O_1804,N_19951,N_19973);
nand UO_1805 (O_1805,N_19845,N_19920);
and UO_1806 (O_1806,N_19881,N_19933);
xor UO_1807 (O_1807,N_19928,N_19958);
nor UO_1808 (O_1808,N_19871,N_19988);
nand UO_1809 (O_1809,N_19989,N_19932);
or UO_1810 (O_1810,N_19992,N_19846);
xnor UO_1811 (O_1811,N_19959,N_19888);
or UO_1812 (O_1812,N_19964,N_19886);
xnor UO_1813 (O_1813,N_19901,N_19931);
xor UO_1814 (O_1814,N_19937,N_19859);
or UO_1815 (O_1815,N_19926,N_19965);
and UO_1816 (O_1816,N_19897,N_19973);
xor UO_1817 (O_1817,N_19854,N_19927);
or UO_1818 (O_1818,N_19875,N_19959);
nand UO_1819 (O_1819,N_19909,N_19870);
or UO_1820 (O_1820,N_19891,N_19926);
and UO_1821 (O_1821,N_19962,N_19951);
nand UO_1822 (O_1822,N_19973,N_19921);
or UO_1823 (O_1823,N_19999,N_19914);
or UO_1824 (O_1824,N_19927,N_19860);
nand UO_1825 (O_1825,N_19896,N_19980);
and UO_1826 (O_1826,N_19904,N_19852);
nor UO_1827 (O_1827,N_19962,N_19897);
and UO_1828 (O_1828,N_19892,N_19845);
or UO_1829 (O_1829,N_19895,N_19919);
and UO_1830 (O_1830,N_19843,N_19867);
nand UO_1831 (O_1831,N_19909,N_19851);
nor UO_1832 (O_1832,N_19888,N_19840);
nor UO_1833 (O_1833,N_19950,N_19856);
xnor UO_1834 (O_1834,N_19860,N_19876);
xor UO_1835 (O_1835,N_19914,N_19899);
or UO_1836 (O_1836,N_19986,N_19888);
nand UO_1837 (O_1837,N_19889,N_19884);
and UO_1838 (O_1838,N_19909,N_19922);
and UO_1839 (O_1839,N_19937,N_19881);
or UO_1840 (O_1840,N_19946,N_19920);
and UO_1841 (O_1841,N_19888,N_19985);
or UO_1842 (O_1842,N_19995,N_19875);
nand UO_1843 (O_1843,N_19979,N_19854);
or UO_1844 (O_1844,N_19991,N_19986);
nor UO_1845 (O_1845,N_19920,N_19917);
and UO_1846 (O_1846,N_19907,N_19972);
nand UO_1847 (O_1847,N_19974,N_19887);
and UO_1848 (O_1848,N_19870,N_19923);
and UO_1849 (O_1849,N_19948,N_19899);
or UO_1850 (O_1850,N_19922,N_19852);
nand UO_1851 (O_1851,N_19849,N_19954);
or UO_1852 (O_1852,N_19880,N_19961);
nand UO_1853 (O_1853,N_19870,N_19982);
xnor UO_1854 (O_1854,N_19852,N_19921);
nand UO_1855 (O_1855,N_19855,N_19947);
nor UO_1856 (O_1856,N_19971,N_19841);
xor UO_1857 (O_1857,N_19845,N_19997);
nor UO_1858 (O_1858,N_19854,N_19947);
xor UO_1859 (O_1859,N_19860,N_19939);
or UO_1860 (O_1860,N_19851,N_19850);
or UO_1861 (O_1861,N_19903,N_19997);
xor UO_1862 (O_1862,N_19906,N_19846);
and UO_1863 (O_1863,N_19899,N_19973);
nand UO_1864 (O_1864,N_19954,N_19890);
and UO_1865 (O_1865,N_19854,N_19975);
nor UO_1866 (O_1866,N_19902,N_19889);
and UO_1867 (O_1867,N_19968,N_19915);
xor UO_1868 (O_1868,N_19875,N_19964);
xnor UO_1869 (O_1869,N_19911,N_19858);
nor UO_1870 (O_1870,N_19942,N_19940);
nor UO_1871 (O_1871,N_19862,N_19913);
or UO_1872 (O_1872,N_19992,N_19918);
nor UO_1873 (O_1873,N_19935,N_19840);
and UO_1874 (O_1874,N_19850,N_19840);
and UO_1875 (O_1875,N_19899,N_19884);
and UO_1876 (O_1876,N_19861,N_19998);
nand UO_1877 (O_1877,N_19978,N_19992);
nand UO_1878 (O_1878,N_19912,N_19846);
and UO_1879 (O_1879,N_19953,N_19930);
xnor UO_1880 (O_1880,N_19971,N_19974);
and UO_1881 (O_1881,N_19886,N_19885);
and UO_1882 (O_1882,N_19843,N_19979);
nand UO_1883 (O_1883,N_19851,N_19843);
and UO_1884 (O_1884,N_19941,N_19855);
or UO_1885 (O_1885,N_19862,N_19996);
nand UO_1886 (O_1886,N_19966,N_19890);
nor UO_1887 (O_1887,N_19844,N_19895);
nor UO_1888 (O_1888,N_19843,N_19840);
and UO_1889 (O_1889,N_19990,N_19870);
and UO_1890 (O_1890,N_19958,N_19879);
and UO_1891 (O_1891,N_19906,N_19979);
nor UO_1892 (O_1892,N_19993,N_19951);
and UO_1893 (O_1893,N_19933,N_19961);
or UO_1894 (O_1894,N_19932,N_19861);
nand UO_1895 (O_1895,N_19989,N_19946);
nand UO_1896 (O_1896,N_19948,N_19987);
or UO_1897 (O_1897,N_19987,N_19904);
and UO_1898 (O_1898,N_19984,N_19925);
and UO_1899 (O_1899,N_19988,N_19908);
nand UO_1900 (O_1900,N_19916,N_19937);
or UO_1901 (O_1901,N_19878,N_19984);
and UO_1902 (O_1902,N_19918,N_19940);
nand UO_1903 (O_1903,N_19974,N_19957);
xnor UO_1904 (O_1904,N_19844,N_19940);
xnor UO_1905 (O_1905,N_19986,N_19988);
or UO_1906 (O_1906,N_19955,N_19947);
xnor UO_1907 (O_1907,N_19961,N_19969);
nor UO_1908 (O_1908,N_19860,N_19992);
or UO_1909 (O_1909,N_19998,N_19952);
or UO_1910 (O_1910,N_19909,N_19953);
and UO_1911 (O_1911,N_19974,N_19925);
or UO_1912 (O_1912,N_19965,N_19937);
and UO_1913 (O_1913,N_19943,N_19985);
xor UO_1914 (O_1914,N_19924,N_19915);
and UO_1915 (O_1915,N_19857,N_19867);
xnor UO_1916 (O_1916,N_19899,N_19962);
nand UO_1917 (O_1917,N_19955,N_19964);
and UO_1918 (O_1918,N_19959,N_19910);
xor UO_1919 (O_1919,N_19892,N_19989);
or UO_1920 (O_1920,N_19929,N_19884);
or UO_1921 (O_1921,N_19895,N_19980);
and UO_1922 (O_1922,N_19890,N_19984);
nand UO_1923 (O_1923,N_19871,N_19958);
xnor UO_1924 (O_1924,N_19865,N_19895);
xnor UO_1925 (O_1925,N_19966,N_19916);
or UO_1926 (O_1926,N_19885,N_19876);
or UO_1927 (O_1927,N_19932,N_19899);
and UO_1928 (O_1928,N_19939,N_19963);
nor UO_1929 (O_1929,N_19971,N_19901);
nand UO_1930 (O_1930,N_19980,N_19904);
nand UO_1931 (O_1931,N_19983,N_19979);
nor UO_1932 (O_1932,N_19992,N_19855);
and UO_1933 (O_1933,N_19882,N_19840);
xnor UO_1934 (O_1934,N_19968,N_19919);
or UO_1935 (O_1935,N_19998,N_19963);
nand UO_1936 (O_1936,N_19844,N_19951);
xnor UO_1937 (O_1937,N_19973,N_19925);
nand UO_1938 (O_1938,N_19850,N_19979);
xor UO_1939 (O_1939,N_19901,N_19968);
nand UO_1940 (O_1940,N_19988,N_19922);
xnor UO_1941 (O_1941,N_19914,N_19893);
and UO_1942 (O_1942,N_19963,N_19906);
and UO_1943 (O_1943,N_19961,N_19991);
or UO_1944 (O_1944,N_19871,N_19984);
nor UO_1945 (O_1945,N_19849,N_19931);
nand UO_1946 (O_1946,N_19926,N_19946);
nand UO_1947 (O_1947,N_19917,N_19896);
nor UO_1948 (O_1948,N_19930,N_19856);
xnor UO_1949 (O_1949,N_19924,N_19987);
or UO_1950 (O_1950,N_19999,N_19966);
nor UO_1951 (O_1951,N_19868,N_19926);
nand UO_1952 (O_1952,N_19857,N_19949);
nor UO_1953 (O_1953,N_19937,N_19977);
and UO_1954 (O_1954,N_19943,N_19939);
and UO_1955 (O_1955,N_19973,N_19964);
or UO_1956 (O_1956,N_19920,N_19944);
and UO_1957 (O_1957,N_19977,N_19982);
nand UO_1958 (O_1958,N_19993,N_19911);
nor UO_1959 (O_1959,N_19988,N_19848);
xor UO_1960 (O_1960,N_19994,N_19863);
and UO_1961 (O_1961,N_19863,N_19895);
or UO_1962 (O_1962,N_19853,N_19983);
or UO_1963 (O_1963,N_19970,N_19846);
nor UO_1964 (O_1964,N_19923,N_19847);
or UO_1965 (O_1965,N_19979,N_19931);
xnor UO_1966 (O_1966,N_19933,N_19921);
nor UO_1967 (O_1967,N_19899,N_19916);
nand UO_1968 (O_1968,N_19958,N_19968);
or UO_1969 (O_1969,N_19964,N_19978);
and UO_1970 (O_1970,N_19981,N_19958);
nand UO_1971 (O_1971,N_19917,N_19859);
or UO_1972 (O_1972,N_19928,N_19946);
nand UO_1973 (O_1973,N_19945,N_19842);
xor UO_1974 (O_1974,N_19909,N_19955);
or UO_1975 (O_1975,N_19938,N_19961);
nor UO_1976 (O_1976,N_19929,N_19868);
nor UO_1977 (O_1977,N_19954,N_19857);
xnor UO_1978 (O_1978,N_19859,N_19982);
xnor UO_1979 (O_1979,N_19972,N_19992);
nor UO_1980 (O_1980,N_19850,N_19854);
xor UO_1981 (O_1981,N_19955,N_19916);
nand UO_1982 (O_1982,N_19948,N_19984);
nand UO_1983 (O_1983,N_19986,N_19875);
xnor UO_1984 (O_1984,N_19946,N_19875);
xnor UO_1985 (O_1985,N_19885,N_19874);
nor UO_1986 (O_1986,N_19984,N_19939);
xor UO_1987 (O_1987,N_19847,N_19935);
and UO_1988 (O_1988,N_19877,N_19926);
nand UO_1989 (O_1989,N_19970,N_19916);
nand UO_1990 (O_1990,N_19966,N_19937);
nor UO_1991 (O_1991,N_19992,N_19866);
nor UO_1992 (O_1992,N_19959,N_19878);
nand UO_1993 (O_1993,N_19849,N_19955);
nor UO_1994 (O_1994,N_19866,N_19984);
or UO_1995 (O_1995,N_19857,N_19858);
and UO_1996 (O_1996,N_19924,N_19860);
and UO_1997 (O_1997,N_19877,N_19935);
nor UO_1998 (O_1998,N_19873,N_19879);
and UO_1999 (O_1999,N_19919,N_19985);
xor UO_2000 (O_2000,N_19906,N_19952);
nor UO_2001 (O_2001,N_19964,N_19876);
and UO_2002 (O_2002,N_19893,N_19843);
or UO_2003 (O_2003,N_19956,N_19904);
nor UO_2004 (O_2004,N_19983,N_19970);
or UO_2005 (O_2005,N_19856,N_19927);
or UO_2006 (O_2006,N_19909,N_19854);
nand UO_2007 (O_2007,N_19975,N_19961);
and UO_2008 (O_2008,N_19874,N_19934);
nor UO_2009 (O_2009,N_19898,N_19949);
and UO_2010 (O_2010,N_19970,N_19968);
nand UO_2011 (O_2011,N_19940,N_19909);
xnor UO_2012 (O_2012,N_19958,N_19915);
nor UO_2013 (O_2013,N_19973,N_19871);
nor UO_2014 (O_2014,N_19918,N_19870);
nand UO_2015 (O_2015,N_19867,N_19888);
and UO_2016 (O_2016,N_19876,N_19970);
xnor UO_2017 (O_2017,N_19914,N_19885);
and UO_2018 (O_2018,N_19994,N_19946);
xnor UO_2019 (O_2019,N_19857,N_19901);
nand UO_2020 (O_2020,N_19886,N_19985);
or UO_2021 (O_2021,N_19973,N_19889);
or UO_2022 (O_2022,N_19906,N_19934);
nand UO_2023 (O_2023,N_19889,N_19967);
nor UO_2024 (O_2024,N_19896,N_19945);
or UO_2025 (O_2025,N_19846,N_19928);
xnor UO_2026 (O_2026,N_19875,N_19916);
nor UO_2027 (O_2027,N_19858,N_19979);
nor UO_2028 (O_2028,N_19858,N_19951);
xnor UO_2029 (O_2029,N_19871,N_19860);
nand UO_2030 (O_2030,N_19899,N_19844);
xor UO_2031 (O_2031,N_19943,N_19915);
nor UO_2032 (O_2032,N_19968,N_19939);
xnor UO_2033 (O_2033,N_19953,N_19993);
and UO_2034 (O_2034,N_19858,N_19850);
nor UO_2035 (O_2035,N_19945,N_19888);
nor UO_2036 (O_2036,N_19879,N_19951);
nor UO_2037 (O_2037,N_19867,N_19845);
and UO_2038 (O_2038,N_19992,N_19930);
xor UO_2039 (O_2039,N_19887,N_19883);
nor UO_2040 (O_2040,N_19967,N_19989);
nor UO_2041 (O_2041,N_19928,N_19988);
nand UO_2042 (O_2042,N_19944,N_19861);
and UO_2043 (O_2043,N_19847,N_19894);
and UO_2044 (O_2044,N_19854,N_19870);
nand UO_2045 (O_2045,N_19929,N_19952);
xnor UO_2046 (O_2046,N_19912,N_19960);
or UO_2047 (O_2047,N_19880,N_19876);
xnor UO_2048 (O_2048,N_19979,N_19974);
xor UO_2049 (O_2049,N_19922,N_19951);
nor UO_2050 (O_2050,N_19992,N_19999);
and UO_2051 (O_2051,N_19929,N_19869);
or UO_2052 (O_2052,N_19923,N_19891);
nand UO_2053 (O_2053,N_19889,N_19953);
nand UO_2054 (O_2054,N_19906,N_19940);
xor UO_2055 (O_2055,N_19857,N_19933);
nand UO_2056 (O_2056,N_19933,N_19882);
or UO_2057 (O_2057,N_19914,N_19877);
or UO_2058 (O_2058,N_19878,N_19869);
nand UO_2059 (O_2059,N_19999,N_19865);
nand UO_2060 (O_2060,N_19893,N_19944);
nand UO_2061 (O_2061,N_19978,N_19868);
or UO_2062 (O_2062,N_19997,N_19914);
and UO_2063 (O_2063,N_19966,N_19887);
xnor UO_2064 (O_2064,N_19863,N_19911);
nor UO_2065 (O_2065,N_19860,N_19872);
or UO_2066 (O_2066,N_19952,N_19935);
or UO_2067 (O_2067,N_19942,N_19986);
nand UO_2068 (O_2068,N_19949,N_19886);
nand UO_2069 (O_2069,N_19994,N_19970);
and UO_2070 (O_2070,N_19913,N_19867);
nor UO_2071 (O_2071,N_19935,N_19966);
nand UO_2072 (O_2072,N_19976,N_19914);
nand UO_2073 (O_2073,N_19885,N_19963);
and UO_2074 (O_2074,N_19991,N_19952);
xor UO_2075 (O_2075,N_19902,N_19846);
xor UO_2076 (O_2076,N_19881,N_19846);
nor UO_2077 (O_2077,N_19964,N_19999);
nor UO_2078 (O_2078,N_19929,N_19919);
and UO_2079 (O_2079,N_19984,N_19962);
and UO_2080 (O_2080,N_19949,N_19850);
nand UO_2081 (O_2081,N_19843,N_19994);
and UO_2082 (O_2082,N_19983,N_19908);
nor UO_2083 (O_2083,N_19921,N_19964);
nor UO_2084 (O_2084,N_19991,N_19866);
nor UO_2085 (O_2085,N_19980,N_19856);
xnor UO_2086 (O_2086,N_19947,N_19915);
nand UO_2087 (O_2087,N_19881,N_19928);
nor UO_2088 (O_2088,N_19981,N_19977);
and UO_2089 (O_2089,N_19948,N_19866);
nand UO_2090 (O_2090,N_19978,N_19997);
xor UO_2091 (O_2091,N_19962,N_19928);
nor UO_2092 (O_2092,N_19893,N_19869);
xor UO_2093 (O_2093,N_19906,N_19993);
nor UO_2094 (O_2094,N_19865,N_19920);
nand UO_2095 (O_2095,N_19934,N_19945);
xor UO_2096 (O_2096,N_19894,N_19945);
or UO_2097 (O_2097,N_19852,N_19893);
and UO_2098 (O_2098,N_19982,N_19865);
or UO_2099 (O_2099,N_19915,N_19926);
nand UO_2100 (O_2100,N_19871,N_19898);
nor UO_2101 (O_2101,N_19946,N_19960);
or UO_2102 (O_2102,N_19982,N_19915);
nor UO_2103 (O_2103,N_19913,N_19882);
xnor UO_2104 (O_2104,N_19850,N_19904);
and UO_2105 (O_2105,N_19905,N_19938);
or UO_2106 (O_2106,N_19944,N_19863);
or UO_2107 (O_2107,N_19929,N_19896);
or UO_2108 (O_2108,N_19946,N_19869);
nand UO_2109 (O_2109,N_19995,N_19997);
or UO_2110 (O_2110,N_19916,N_19871);
xnor UO_2111 (O_2111,N_19934,N_19974);
and UO_2112 (O_2112,N_19948,N_19944);
nand UO_2113 (O_2113,N_19862,N_19878);
or UO_2114 (O_2114,N_19864,N_19931);
and UO_2115 (O_2115,N_19977,N_19952);
nand UO_2116 (O_2116,N_19941,N_19849);
or UO_2117 (O_2117,N_19939,N_19849);
and UO_2118 (O_2118,N_19936,N_19875);
or UO_2119 (O_2119,N_19879,N_19874);
or UO_2120 (O_2120,N_19849,N_19897);
xor UO_2121 (O_2121,N_19944,N_19915);
nand UO_2122 (O_2122,N_19983,N_19965);
nand UO_2123 (O_2123,N_19868,N_19870);
and UO_2124 (O_2124,N_19876,N_19867);
or UO_2125 (O_2125,N_19995,N_19993);
xor UO_2126 (O_2126,N_19861,N_19889);
nor UO_2127 (O_2127,N_19892,N_19918);
nor UO_2128 (O_2128,N_19913,N_19912);
or UO_2129 (O_2129,N_19927,N_19926);
xnor UO_2130 (O_2130,N_19871,N_19897);
xor UO_2131 (O_2131,N_19937,N_19945);
or UO_2132 (O_2132,N_19965,N_19859);
xnor UO_2133 (O_2133,N_19877,N_19937);
and UO_2134 (O_2134,N_19999,N_19995);
nand UO_2135 (O_2135,N_19863,N_19943);
nor UO_2136 (O_2136,N_19881,N_19964);
and UO_2137 (O_2137,N_19864,N_19903);
xor UO_2138 (O_2138,N_19967,N_19922);
or UO_2139 (O_2139,N_19846,N_19841);
xor UO_2140 (O_2140,N_19945,N_19914);
or UO_2141 (O_2141,N_19885,N_19944);
and UO_2142 (O_2142,N_19941,N_19888);
nand UO_2143 (O_2143,N_19924,N_19880);
or UO_2144 (O_2144,N_19913,N_19859);
or UO_2145 (O_2145,N_19899,N_19935);
xnor UO_2146 (O_2146,N_19857,N_19939);
and UO_2147 (O_2147,N_19860,N_19899);
nor UO_2148 (O_2148,N_19977,N_19878);
nand UO_2149 (O_2149,N_19930,N_19882);
and UO_2150 (O_2150,N_19851,N_19940);
and UO_2151 (O_2151,N_19861,N_19884);
xor UO_2152 (O_2152,N_19972,N_19998);
nor UO_2153 (O_2153,N_19938,N_19870);
or UO_2154 (O_2154,N_19956,N_19910);
or UO_2155 (O_2155,N_19881,N_19900);
xnor UO_2156 (O_2156,N_19920,N_19906);
or UO_2157 (O_2157,N_19934,N_19960);
and UO_2158 (O_2158,N_19929,N_19900);
nand UO_2159 (O_2159,N_19888,N_19954);
nand UO_2160 (O_2160,N_19976,N_19992);
xnor UO_2161 (O_2161,N_19924,N_19865);
and UO_2162 (O_2162,N_19968,N_19891);
and UO_2163 (O_2163,N_19906,N_19996);
nor UO_2164 (O_2164,N_19985,N_19993);
and UO_2165 (O_2165,N_19850,N_19984);
or UO_2166 (O_2166,N_19857,N_19923);
xor UO_2167 (O_2167,N_19885,N_19932);
xnor UO_2168 (O_2168,N_19926,N_19897);
nand UO_2169 (O_2169,N_19985,N_19949);
xnor UO_2170 (O_2170,N_19901,N_19896);
xor UO_2171 (O_2171,N_19898,N_19987);
nand UO_2172 (O_2172,N_19848,N_19879);
xnor UO_2173 (O_2173,N_19934,N_19857);
or UO_2174 (O_2174,N_19901,N_19970);
and UO_2175 (O_2175,N_19924,N_19990);
and UO_2176 (O_2176,N_19841,N_19917);
or UO_2177 (O_2177,N_19949,N_19902);
and UO_2178 (O_2178,N_19988,N_19878);
nand UO_2179 (O_2179,N_19878,N_19921);
xor UO_2180 (O_2180,N_19927,N_19961);
or UO_2181 (O_2181,N_19897,N_19966);
nor UO_2182 (O_2182,N_19869,N_19881);
nor UO_2183 (O_2183,N_19889,N_19928);
xnor UO_2184 (O_2184,N_19919,N_19852);
or UO_2185 (O_2185,N_19955,N_19862);
nand UO_2186 (O_2186,N_19970,N_19969);
xor UO_2187 (O_2187,N_19940,N_19873);
nand UO_2188 (O_2188,N_19874,N_19899);
or UO_2189 (O_2189,N_19972,N_19917);
nand UO_2190 (O_2190,N_19878,N_19860);
nor UO_2191 (O_2191,N_19951,N_19932);
or UO_2192 (O_2192,N_19950,N_19941);
xor UO_2193 (O_2193,N_19935,N_19931);
or UO_2194 (O_2194,N_19859,N_19956);
xnor UO_2195 (O_2195,N_19969,N_19892);
and UO_2196 (O_2196,N_19877,N_19905);
nor UO_2197 (O_2197,N_19949,N_19972);
and UO_2198 (O_2198,N_19859,N_19858);
and UO_2199 (O_2199,N_19992,N_19934);
xor UO_2200 (O_2200,N_19949,N_19947);
and UO_2201 (O_2201,N_19996,N_19921);
and UO_2202 (O_2202,N_19866,N_19894);
nand UO_2203 (O_2203,N_19918,N_19859);
or UO_2204 (O_2204,N_19964,N_19983);
xnor UO_2205 (O_2205,N_19954,N_19877);
and UO_2206 (O_2206,N_19886,N_19980);
xnor UO_2207 (O_2207,N_19917,N_19875);
or UO_2208 (O_2208,N_19880,N_19916);
nor UO_2209 (O_2209,N_19907,N_19947);
nand UO_2210 (O_2210,N_19971,N_19942);
nor UO_2211 (O_2211,N_19957,N_19950);
xnor UO_2212 (O_2212,N_19899,N_19864);
or UO_2213 (O_2213,N_19845,N_19922);
nand UO_2214 (O_2214,N_19987,N_19876);
xnor UO_2215 (O_2215,N_19879,N_19974);
and UO_2216 (O_2216,N_19893,N_19862);
or UO_2217 (O_2217,N_19924,N_19892);
xor UO_2218 (O_2218,N_19938,N_19880);
xnor UO_2219 (O_2219,N_19847,N_19946);
nand UO_2220 (O_2220,N_19862,N_19866);
or UO_2221 (O_2221,N_19993,N_19909);
and UO_2222 (O_2222,N_19910,N_19982);
nand UO_2223 (O_2223,N_19989,N_19944);
nand UO_2224 (O_2224,N_19855,N_19912);
xor UO_2225 (O_2225,N_19932,N_19888);
and UO_2226 (O_2226,N_19883,N_19850);
nand UO_2227 (O_2227,N_19975,N_19995);
and UO_2228 (O_2228,N_19981,N_19928);
nand UO_2229 (O_2229,N_19894,N_19935);
nor UO_2230 (O_2230,N_19906,N_19851);
xor UO_2231 (O_2231,N_19968,N_19903);
or UO_2232 (O_2232,N_19929,N_19921);
xnor UO_2233 (O_2233,N_19854,N_19948);
and UO_2234 (O_2234,N_19873,N_19852);
xnor UO_2235 (O_2235,N_19895,N_19886);
and UO_2236 (O_2236,N_19940,N_19969);
nand UO_2237 (O_2237,N_19938,N_19990);
nor UO_2238 (O_2238,N_19848,N_19914);
xor UO_2239 (O_2239,N_19987,N_19974);
nand UO_2240 (O_2240,N_19989,N_19959);
nand UO_2241 (O_2241,N_19979,N_19912);
and UO_2242 (O_2242,N_19898,N_19923);
nor UO_2243 (O_2243,N_19930,N_19996);
xnor UO_2244 (O_2244,N_19954,N_19940);
and UO_2245 (O_2245,N_19913,N_19887);
nand UO_2246 (O_2246,N_19911,N_19990);
and UO_2247 (O_2247,N_19867,N_19966);
nor UO_2248 (O_2248,N_19850,N_19962);
nand UO_2249 (O_2249,N_19941,N_19881);
or UO_2250 (O_2250,N_19926,N_19976);
nand UO_2251 (O_2251,N_19953,N_19869);
xnor UO_2252 (O_2252,N_19843,N_19907);
and UO_2253 (O_2253,N_19981,N_19931);
and UO_2254 (O_2254,N_19937,N_19917);
or UO_2255 (O_2255,N_19876,N_19909);
xor UO_2256 (O_2256,N_19909,N_19883);
nand UO_2257 (O_2257,N_19883,N_19957);
or UO_2258 (O_2258,N_19863,N_19930);
or UO_2259 (O_2259,N_19962,N_19841);
or UO_2260 (O_2260,N_19931,N_19874);
or UO_2261 (O_2261,N_19948,N_19879);
and UO_2262 (O_2262,N_19938,N_19967);
xor UO_2263 (O_2263,N_19907,N_19970);
or UO_2264 (O_2264,N_19981,N_19859);
nor UO_2265 (O_2265,N_19960,N_19871);
nand UO_2266 (O_2266,N_19983,N_19871);
or UO_2267 (O_2267,N_19843,N_19912);
and UO_2268 (O_2268,N_19943,N_19895);
and UO_2269 (O_2269,N_19848,N_19980);
nand UO_2270 (O_2270,N_19916,N_19887);
nand UO_2271 (O_2271,N_19900,N_19886);
nor UO_2272 (O_2272,N_19942,N_19969);
and UO_2273 (O_2273,N_19982,N_19978);
and UO_2274 (O_2274,N_19863,N_19960);
or UO_2275 (O_2275,N_19910,N_19905);
and UO_2276 (O_2276,N_19848,N_19846);
or UO_2277 (O_2277,N_19872,N_19980);
and UO_2278 (O_2278,N_19950,N_19913);
xor UO_2279 (O_2279,N_19972,N_19879);
and UO_2280 (O_2280,N_19982,N_19894);
and UO_2281 (O_2281,N_19947,N_19948);
or UO_2282 (O_2282,N_19977,N_19990);
nand UO_2283 (O_2283,N_19973,N_19986);
nand UO_2284 (O_2284,N_19920,N_19992);
or UO_2285 (O_2285,N_19846,N_19973);
nor UO_2286 (O_2286,N_19909,N_19910);
nor UO_2287 (O_2287,N_19873,N_19913);
and UO_2288 (O_2288,N_19992,N_19897);
nand UO_2289 (O_2289,N_19924,N_19954);
nand UO_2290 (O_2290,N_19843,N_19939);
or UO_2291 (O_2291,N_19938,N_19859);
or UO_2292 (O_2292,N_19899,N_19875);
nor UO_2293 (O_2293,N_19996,N_19885);
and UO_2294 (O_2294,N_19999,N_19906);
xor UO_2295 (O_2295,N_19946,N_19876);
xor UO_2296 (O_2296,N_19864,N_19856);
nor UO_2297 (O_2297,N_19867,N_19852);
or UO_2298 (O_2298,N_19974,N_19885);
or UO_2299 (O_2299,N_19970,N_19951);
or UO_2300 (O_2300,N_19975,N_19922);
xor UO_2301 (O_2301,N_19898,N_19988);
xor UO_2302 (O_2302,N_19999,N_19919);
or UO_2303 (O_2303,N_19896,N_19881);
xnor UO_2304 (O_2304,N_19929,N_19959);
nand UO_2305 (O_2305,N_19908,N_19855);
nor UO_2306 (O_2306,N_19893,N_19985);
or UO_2307 (O_2307,N_19930,N_19936);
nor UO_2308 (O_2308,N_19909,N_19931);
and UO_2309 (O_2309,N_19915,N_19989);
or UO_2310 (O_2310,N_19847,N_19992);
xor UO_2311 (O_2311,N_19855,N_19999);
and UO_2312 (O_2312,N_19869,N_19974);
nor UO_2313 (O_2313,N_19901,N_19860);
or UO_2314 (O_2314,N_19959,N_19871);
nand UO_2315 (O_2315,N_19842,N_19866);
xnor UO_2316 (O_2316,N_19957,N_19918);
nand UO_2317 (O_2317,N_19927,N_19935);
nand UO_2318 (O_2318,N_19936,N_19891);
nand UO_2319 (O_2319,N_19968,N_19859);
or UO_2320 (O_2320,N_19882,N_19928);
nand UO_2321 (O_2321,N_19925,N_19962);
nor UO_2322 (O_2322,N_19962,N_19881);
xnor UO_2323 (O_2323,N_19977,N_19877);
xnor UO_2324 (O_2324,N_19944,N_19860);
nor UO_2325 (O_2325,N_19914,N_19922);
nor UO_2326 (O_2326,N_19847,N_19863);
or UO_2327 (O_2327,N_19937,N_19866);
nor UO_2328 (O_2328,N_19939,N_19978);
and UO_2329 (O_2329,N_19967,N_19893);
or UO_2330 (O_2330,N_19943,N_19881);
nand UO_2331 (O_2331,N_19997,N_19965);
nand UO_2332 (O_2332,N_19950,N_19841);
or UO_2333 (O_2333,N_19922,N_19985);
nand UO_2334 (O_2334,N_19889,N_19860);
and UO_2335 (O_2335,N_19960,N_19938);
nand UO_2336 (O_2336,N_19842,N_19996);
nor UO_2337 (O_2337,N_19914,N_19918);
or UO_2338 (O_2338,N_19846,N_19885);
nor UO_2339 (O_2339,N_19844,N_19998);
and UO_2340 (O_2340,N_19918,N_19954);
or UO_2341 (O_2341,N_19981,N_19953);
nor UO_2342 (O_2342,N_19939,N_19856);
and UO_2343 (O_2343,N_19927,N_19975);
xnor UO_2344 (O_2344,N_19971,N_19851);
or UO_2345 (O_2345,N_19947,N_19898);
xnor UO_2346 (O_2346,N_19993,N_19854);
or UO_2347 (O_2347,N_19903,N_19882);
and UO_2348 (O_2348,N_19875,N_19983);
nor UO_2349 (O_2349,N_19899,N_19944);
and UO_2350 (O_2350,N_19959,N_19864);
and UO_2351 (O_2351,N_19892,N_19876);
nor UO_2352 (O_2352,N_19938,N_19879);
or UO_2353 (O_2353,N_19966,N_19841);
xnor UO_2354 (O_2354,N_19907,N_19990);
and UO_2355 (O_2355,N_19877,N_19840);
xor UO_2356 (O_2356,N_19989,N_19963);
or UO_2357 (O_2357,N_19954,N_19860);
or UO_2358 (O_2358,N_19851,N_19948);
nor UO_2359 (O_2359,N_19993,N_19984);
xor UO_2360 (O_2360,N_19866,N_19989);
and UO_2361 (O_2361,N_19960,N_19942);
and UO_2362 (O_2362,N_19957,N_19988);
xor UO_2363 (O_2363,N_19970,N_19899);
and UO_2364 (O_2364,N_19993,N_19923);
xnor UO_2365 (O_2365,N_19959,N_19847);
or UO_2366 (O_2366,N_19997,N_19877);
or UO_2367 (O_2367,N_19993,N_19885);
nor UO_2368 (O_2368,N_19981,N_19898);
xnor UO_2369 (O_2369,N_19919,N_19936);
nor UO_2370 (O_2370,N_19917,N_19946);
nand UO_2371 (O_2371,N_19998,N_19948);
and UO_2372 (O_2372,N_19984,N_19955);
nor UO_2373 (O_2373,N_19957,N_19977);
nor UO_2374 (O_2374,N_19861,N_19921);
and UO_2375 (O_2375,N_19887,N_19857);
and UO_2376 (O_2376,N_19932,N_19927);
nor UO_2377 (O_2377,N_19968,N_19962);
nand UO_2378 (O_2378,N_19964,N_19992);
xnor UO_2379 (O_2379,N_19851,N_19916);
xor UO_2380 (O_2380,N_19977,N_19955);
or UO_2381 (O_2381,N_19849,N_19865);
xor UO_2382 (O_2382,N_19860,N_19963);
and UO_2383 (O_2383,N_19992,N_19916);
nand UO_2384 (O_2384,N_19969,N_19851);
xor UO_2385 (O_2385,N_19863,N_19861);
nor UO_2386 (O_2386,N_19919,N_19911);
nand UO_2387 (O_2387,N_19870,N_19935);
or UO_2388 (O_2388,N_19997,N_19968);
and UO_2389 (O_2389,N_19991,N_19877);
nand UO_2390 (O_2390,N_19960,N_19903);
and UO_2391 (O_2391,N_19897,N_19885);
xor UO_2392 (O_2392,N_19932,N_19934);
or UO_2393 (O_2393,N_19997,N_19935);
nor UO_2394 (O_2394,N_19995,N_19966);
and UO_2395 (O_2395,N_19885,N_19864);
and UO_2396 (O_2396,N_19927,N_19858);
nand UO_2397 (O_2397,N_19988,N_19930);
or UO_2398 (O_2398,N_19931,N_19945);
nor UO_2399 (O_2399,N_19928,N_19912);
xnor UO_2400 (O_2400,N_19967,N_19933);
and UO_2401 (O_2401,N_19885,N_19937);
nor UO_2402 (O_2402,N_19995,N_19861);
nand UO_2403 (O_2403,N_19867,N_19958);
or UO_2404 (O_2404,N_19949,N_19967);
or UO_2405 (O_2405,N_19883,N_19854);
or UO_2406 (O_2406,N_19932,N_19984);
nor UO_2407 (O_2407,N_19950,N_19852);
xor UO_2408 (O_2408,N_19915,N_19878);
or UO_2409 (O_2409,N_19964,N_19995);
nor UO_2410 (O_2410,N_19851,N_19888);
and UO_2411 (O_2411,N_19901,N_19999);
and UO_2412 (O_2412,N_19972,N_19916);
xor UO_2413 (O_2413,N_19993,N_19954);
nand UO_2414 (O_2414,N_19842,N_19840);
nand UO_2415 (O_2415,N_19955,N_19842);
xnor UO_2416 (O_2416,N_19884,N_19910);
nand UO_2417 (O_2417,N_19980,N_19990);
and UO_2418 (O_2418,N_19840,N_19957);
nor UO_2419 (O_2419,N_19987,N_19986);
xor UO_2420 (O_2420,N_19928,N_19951);
and UO_2421 (O_2421,N_19920,N_19864);
xnor UO_2422 (O_2422,N_19870,N_19971);
nand UO_2423 (O_2423,N_19943,N_19954);
nand UO_2424 (O_2424,N_19890,N_19996);
nand UO_2425 (O_2425,N_19880,N_19915);
nor UO_2426 (O_2426,N_19844,N_19870);
or UO_2427 (O_2427,N_19880,N_19955);
nor UO_2428 (O_2428,N_19982,N_19840);
xnor UO_2429 (O_2429,N_19939,N_19958);
or UO_2430 (O_2430,N_19894,N_19994);
nand UO_2431 (O_2431,N_19941,N_19973);
and UO_2432 (O_2432,N_19863,N_19853);
nand UO_2433 (O_2433,N_19977,N_19951);
nor UO_2434 (O_2434,N_19877,N_19975);
nor UO_2435 (O_2435,N_19850,N_19973);
xnor UO_2436 (O_2436,N_19966,N_19969);
xor UO_2437 (O_2437,N_19934,N_19965);
xor UO_2438 (O_2438,N_19995,N_19854);
nand UO_2439 (O_2439,N_19969,N_19938);
or UO_2440 (O_2440,N_19903,N_19880);
and UO_2441 (O_2441,N_19840,N_19896);
or UO_2442 (O_2442,N_19888,N_19933);
nand UO_2443 (O_2443,N_19949,N_19854);
xor UO_2444 (O_2444,N_19936,N_19877);
xor UO_2445 (O_2445,N_19938,N_19842);
nor UO_2446 (O_2446,N_19842,N_19961);
nand UO_2447 (O_2447,N_19895,N_19847);
nand UO_2448 (O_2448,N_19966,N_19977);
nand UO_2449 (O_2449,N_19935,N_19874);
xor UO_2450 (O_2450,N_19900,N_19937);
nor UO_2451 (O_2451,N_19878,N_19951);
or UO_2452 (O_2452,N_19961,N_19944);
or UO_2453 (O_2453,N_19852,N_19986);
xnor UO_2454 (O_2454,N_19944,N_19880);
and UO_2455 (O_2455,N_19893,N_19925);
or UO_2456 (O_2456,N_19988,N_19907);
or UO_2457 (O_2457,N_19900,N_19879);
or UO_2458 (O_2458,N_19873,N_19925);
and UO_2459 (O_2459,N_19872,N_19954);
nand UO_2460 (O_2460,N_19926,N_19969);
nor UO_2461 (O_2461,N_19927,N_19982);
and UO_2462 (O_2462,N_19964,N_19892);
or UO_2463 (O_2463,N_19990,N_19876);
xor UO_2464 (O_2464,N_19977,N_19934);
nor UO_2465 (O_2465,N_19988,N_19847);
nor UO_2466 (O_2466,N_19853,N_19845);
or UO_2467 (O_2467,N_19982,N_19841);
and UO_2468 (O_2468,N_19928,N_19878);
nand UO_2469 (O_2469,N_19964,N_19974);
or UO_2470 (O_2470,N_19922,N_19944);
nand UO_2471 (O_2471,N_19942,N_19864);
or UO_2472 (O_2472,N_19885,N_19860);
nor UO_2473 (O_2473,N_19872,N_19920);
or UO_2474 (O_2474,N_19906,N_19946);
and UO_2475 (O_2475,N_19931,N_19951);
nand UO_2476 (O_2476,N_19961,N_19946);
nand UO_2477 (O_2477,N_19998,N_19977);
xor UO_2478 (O_2478,N_19855,N_19882);
nand UO_2479 (O_2479,N_19871,N_19986);
nor UO_2480 (O_2480,N_19934,N_19966);
or UO_2481 (O_2481,N_19872,N_19910);
or UO_2482 (O_2482,N_19851,N_19842);
nor UO_2483 (O_2483,N_19928,N_19968);
nor UO_2484 (O_2484,N_19842,N_19853);
xnor UO_2485 (O_2485,N_19919,N_19890);
and UO_2486 (O_2486,N_19914,N_19946);
or UO_2487 (O_2487,N_19862,N_19956);
nor UO_2488 (O_2488,N_19873,N_19968);
or UO_2489 (O_2489,N_19857,N_19938);
and UO_2490 (O_2490,N_19914,N_19896);
and UO_2491 (O_2491,N_19903,N_19874);
nand UO_2492 (O_2492,N_19925,N_19965);
and UO_2493 (O_2493,N_19990,N_19982);
nand UO_2494 (O_2494,N_19933,N_19951);
nor UO_2495 (O_2495,N_19984,N_19895);
nand UO_2496 (O_2496,N_19879,N_19967);
or UO_2497 (O_2497,N_19996,N_19951);
xor UO_2498 (O_2498,N_19842,N_19893);
and UO_2499 (O_2499,N_19997,N_19950);
endmodule