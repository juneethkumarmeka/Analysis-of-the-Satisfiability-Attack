module basic_1500_15000_2000_50_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
xor U0 (N_0,In_165,In_1143);
and U1 (N_1,In_1061,In_864);
and U2 (N_2,In_842,In_147);
or U3 (N_3,In_710,In_252);
nand U4 (N_4,In_398,In_42);
nor U5 (N_5,In_778,In_622);
or U6 (N_6,In_1039,In_579);
xor U7 (N_7,In_907,In_784);
and U8 (N_8,In_951,In_739);
nor U9 (N_9,In_586,In_930);
and U10 (N_10,In_1194,In_1110);
nor U11 (N_11,In_585,In_146);
nor U12 (N_12,In_599,In_509);
nor U13 (N_13,In_1254,In_94);
and U14 (N_14,In_1083,In_416);
nand U15 (N_15,In_435,In_1414);
or U16 (N_16,In_1478,In_23);
or U17 (N_17,In_724,In_988);
xnor U18 (N_18,In_1227,In_625);
and U19 (N_19,In_333,In_1242);
xnor U20 (N_20,In_313,In_1412);
nand U21 (N_21,In_823,In_872);
and U22 (N_22,In_1329,In_565);
xnor U23 (N_23,In_1308,In_88);
nand U24 (N_24,In_1002,In_795);
nand U25 (N_25,In_689,In_1098);
xnor U26 (N_26,In_47,In_1131);
and U27 (N_27,In_1344,In_853);
and U28 (N_28,In_664,In_63);
and U29 (N_29,In_471,In_1080);
and U30 (N_30,In_1427,In_1332);
nand U31 (N_31,In_745,In_1374);
xnor U32 (N_32,In_366,In_556);
nand U33 (N_33,In_377,In_33);
xor U34 (N_34,In_1073,In_1237);
nor U35 (N_35,In_1186,In_1221);
nand U36 (N_36,In_756,In_187);
nand U37 (N_37,In_250,In_1345);
or U38 (N_38,In_1157,In_300);
nor U39 (N_39,In_1063,In_67);
nand U40 (N_40,In_198,In_761);
xor U41 (N_41,In_125,In_72);
nor U42 (N_42,In_1303,In_32);
or U43 (N_43,In_1159,In_84);
xnor U44 (N_44,In_727,In_518);
or U45 (N_45,In_1078,In_192);
and U46 (N_46,In_1177,In_260);
and U47 (N_47,In_877,In_666);
nor U48 (N_48,In_726,In_145);
nand U49 (N_49,In_623,In_259);
nor U50 (N_50,In_673,In_52);
and U51 (N_51,In_1342,In_858);
and U52 (N_52,In_913,In_845);
nand U53 (N_53,In_48,In_323);
or U54 (N_54,In_31,In_261);
nor U55 (N_55,In_854,In_19);
xnor U56 (N_56,In_1385,In_127);
xnor U57 (N_57,In_244,In_8);
or U58 (N_58,In_640,In_232);
nor U59 (N_59,In_642,In_199);
nand U60 (N_60,In_57,In_1466);
or U61 (N_61,In_144,In_849);
xor U62 (N_62,In_831,In_46);
and U63 (N_63,In_593,In_765);
xor U64 (N_64,In_286,In_275);
or U65 (N_65,In_967,In_97);
and U66 (N_66,In_1264,In_178);
nand U67 (N_67,In_1093,In_278);
xnor U68 (N_68,In_975,In_1053);
and U69 (N_69,In_9,In_119);
or U70 (N_70,In_321,In_177);
and U71 (N_71,In_966,In_457);
and U72 (N_72,In_1323,In_963);
nand U73 (N_73,In_701,In_385);
or U74 (N_74,In_444,In_965);
xnor U75 (N_75,In_357,In_1268);
nand U76 (N_76,In_277,In_1386);
or U77 (N_77,In_671,In_1023);
nor U78 (N_78,In_1096,In_11);
or U79 (N_79,In_825,In_785);
nor U80 (N_80,In_1284,In_1260);
nand U81 (N_81,In_284,In_208);
and U82 (N_82,In_972,In_847);
nor U83 (N_83,In_304,In_424);
or U84 (N_84,In_1309,In_1119);
xor U85 (N_85,In_1072,In_605);
xnor U86 (N_86,In_1442,In_179);
nand U87 (N_87,In_2,In_396);
and U88 (N_88,In_306,In_86);
xor U89 (N_89,In_356,In_1265);
or U90 (N_90,In_1141,In_746);
and U91 (N_91,In_1140,In_279);
and U92 (N_92,In_962,In_1108);
nor U93 (N_93,In_743,In_757);
and U94 (N_94,In_753,In_1241);
and U95 (N_95,In_76,In_941);
or U96 (N_96,In_1132,In_1448);
nand U97 (N_97,In_1364,In_737);
or U98 (N_98,In_866,In_412);
nor U99 (N_99,In_793,In_994);
or U100 (N_100,In_1162,In_769);
and U101 (N_101,In_694,In_821);
xnor U102 (N_102,In_291,In_536);
and U103 (N_103,In_944,In_862);
nor U104 (N_104,In_417,In_1250);
xnor U105 (N_105,In_607,In_855);
nor U106 (N_106,In_740,In_1409);
nor U107 (N_107,In_503,In_632);
nand U108 (N_108,In_368,In_1188);
and U109 (N_109,In_1319,In_129);
nor U110 (N_110,In_58,In_1278);
and U111 (N_111,In_355,In_1213);
and U112 (N_112,In_229,In_686);
xnor U113 (N_113,In_181,In_820);
nand U114 (N_114,In_810,In_519);
and U115 (N_115,In_1088,In_915);
nor U116 (N_116,In_113,In_26);
nor U117 (N_117,In_197,In_834);
xor U118 (N_118,In_557,In_904);
and U119 (N_119,In_1315,In_830);
and U120 (N_120,In_1102,In_383);
xor U121 (N_121,In_505,In_719);
nor U122 (N_122,In_819,In_818);
or U123 (N_123,In_1210,In_1279);
nor U124 (N_124,In_413,In_345);
nand U125 (N_125,In_263,In_1335);
nand U126 (N_126,In_1033,In_652);
and U127 (N_127,In_814,In_438);
xor U128 (N_128,In_79,In_779);
and U129 (N_129,In_875,In_1152);
or U130 (N_130,In_932,In_816);
nand U131 (N_131,In_73,In_215);
nand U132 (N_132,In_1321,In_530);
or U133 (N_133,In_859,In_560);
nand U134 (N_134,In_1195,In_777);
or U135 (N_135,In_93,In_61);
or U136 (N_136,In_400,In_1014);
nor U137 (N_137,In_885,In_1113);
and U138 (N_138,In_461,In_337);
nor U139 (N_139,In_449,In_527);
xor U140 (N_140,In_334,In_812);
or U141 (N_141,In_324,In_910);
and U142 (N_142,In_683,In_470);
xor U143 (N_143,In_307,In_587);
nor U144 (N_144,In_415,In_1300);
xor U145 (N_145,In_718,In_1231);
or U146 (N_146,In_836,In_1355);
nor U147 (N_147,In_191,In_308);
nor U148 (N_148,In_631,In_50);
or U149 (N_149,In_608,In_1290);
nand U150 (N_150,In_1367,In_218);
or U151 (N_151,In_1037,In_603);
nor U152 (N_152,In_1144,In_1469);
nand U153 (N_153,In_639,In_832);
and U154 (N_154,In_1079,In_645);
xnor U155 (N_155,In_564,In_616);
or U156 (N_156,In_302,In_132);
or U157 (N_157,In_708,In_1354);
or U158 (N_158,In_1410,In_1187);
nand U159 (N_159,In_99,In_1200);
xnor U160 (N_160,In_1097,In_950);
or U161 (N_161,In_817,In_1408);
or U162 (N_162,In_574,In_713);
nor U163 (N_163,In_1310,In_647);
or U164 (N_164,In_791,In_706);
or U165 (N_165,In_251,In_1261);
or U166 (N_166,In_936,In_1050);
or U167 (N_167,In_728,In_636);
nand U168 (N_168,In_418,In_576);
nor U169 (N_169,In_696,In_946);
nand U170 (N_170,In_1196,In_531);
nor U171 (N_171,In_421,In_613);
nor U172 (N_172,In_38,In_839);
nor U173 (N_173,In_1293,In_1361);
or U174 (N_174,In_206,In_1009);
or U175 (N_175,In_1433,In_943);
nor U176 (N_176,In_365,In_811);
and U177 (N_177,In_265,In_594);
and U178 (N_178,In_1042,In_1225);
and U179 (N_179,In_285,In_1358);
xnor U180 (N_180,In_399,In_1123);
nor U181 (N_181,In_241,In_1327);
xnor U182 (N_182,In_1435,In_1223);
and U183 (N_183,In_34,In_908);
xnor U184 (N_184,In_1005,In_155);
and U185 (N_185,In_17,In_550);
xor U186 (N_186,In_1467,In_826);
nor U187 (N_187,In_217,In_234);
xor U188 (N_188,In_1322,In_1107);
and U189 (N_189,In_469,In_749);
xor U190 (N_190,In_1135,In_873);
and U191 (N_191,In_380,In_236);
nand U192 (N_192,In_295,In_18);
nor U193 (N_193,In_1205,In_592);
nor U194 (N_194,In_629,In_868);
or U195 (N_195,In_1154,In_1359);
xnor U196 (N_196,In_140,In_1022);
nand U197 (N_197,In_269,In_750);
and U198 (N_198,In_1394,In_1199);
nand U199 (N_199,In_239,In_1288);
or U200 (N_200,In_29,In_233);
nand U201 (N_201,In_1054,In_36);
or U202 (N_202,In_1473,In_1112);
nor U203 (N_203,In_219,In_1100);
and U204 (N_204,In_1198,In_1276);
nor U205 (N_205,In_1007,In_56);
xor U206 (N_206,In_1301,In_95);
or U207 (N_207,In_487,In_397);
or U208 (N_208,In_691,In_997);
and U209 (N_209,In_1437,In_101);
xor U210 (N_210,In_815,In_1403);
xor U211 (N_211,In_867,In_747);
nor U212 (N_212,In_1420,In_153);
and U213 (N_213,In_865,In_1145);
xnor U214 (N_214,In_1189,In_1398);
nand U215 (N_215,In_247,In_1299);
and U216 (N_216,In_894,In_1451);
nand U217 (N_217,In_175,In_1249);
xor U218 (N_218,In_1158,In_1090);
xnor U219 (N_219,In_288,In_433);
nor U220 (N_220,In_1226,In_797);
nand U221 (N_221,In_387,In_89);
or U222 (N_222,In_389,In_827);
xnor U223 (N_223,In_1428,In_524);
nor U224 (N_224,In_445,In_1027);
nand U225 (N_225,In_391,In_1269);
nand U226 (N_226,In_266,In_974);
and U227 (N_227,In_1092,In_1010);
and U228 (N_228,In_262,In_476);
xnor U229 (N_229,In_310,In_346);
nand U230 (N_230,In_508,In_362);
nand U231 (N_231,In_1085,In_102);
and U232 (N_232,In_1470,In_1047);
or U233 (N_233,In_1058,In_870);
xor U234 (N_234,In_453,In_981);
nand U235 (N_235,In_428,In_624);
xnor U236 (N_236,In_431,In_672);
or U237 (N_237,In_567,In_137);
and U238 (N_238,In_43,In_1401);
nand U239 (N_239,In_895,In_927);
and U240 (N_240,In_690,In_712);
and U241 (N_241,In_989,In_643);
xnor U242 (N_242,In_637,In_552);
or U243 (N_243,In_1233,In_69);
or U244 (N_244,In_1230,In_379);
xnor U245 (N_245,In_840,In_744);
nand U246 (N_246,In_361,In_714);
or U247 (N_247,In_1148,In_0);
xnor U248 (N_248,In_730,In_1404);
nand U249 (N_249,In_610,In_1128);
xnor U250 (N_250,In_674,In_316);
or U251 (N_251,In_1064,In_1498);
nor U252 (N_252,In_114,In_837);
or U253 (N_253,In_243,In_1051);
and U254 (N_254,In_376,In_602);
and U255 (N_255,In_841,In_1118);
and U256 (N_256,In_1314,In_1219);
or U257 (N_257,In_343,In_371);
and U258 (N_258,In_452,In_955);
and U259 (N_259,In_1103,In_798);
nand U260 (N_260,In_675,In_276);
or U261 (N_261,In_1173,In_722);
nand U262 (N_262,In_1417,In_41);
xnor U263 (N_263,In_486,In_937);
nand U264 (N_264,In_693,In_4);
xnor U265 (N_265,In_543,In_976);
nand U266 (N_266,In_960,In_615);
nand U267 (N_267,In_143,In_1266);
and U268 (N_268,In_878,In_511);
nor U269 (N_269,In_314,In_1245);
xnor U270 (N_270,In_548,In_157);
xor U271 (N_271,In_1275,In_896);
xor U272 (N_272,In_1235,In_500);
and U273 (N_273,In_1087,In_256);
nand U274 (N_274,In_1295,In_583);
or U275 (N_275,In_949,In_212);
xor U276 (N_276,In_935,In_271);
xor U277 (N_277,In_1445,In_663);
xnor U278 (N_278,In_1418,In_83);
xnor U279 (N_279,In_386,In_1487);
nand U280 (N_280,In_919,In_350);
xnor U281 (N_281,In_479,In_62);
nand U282 (N_282,In_1244,In_169);
and U283 (N_283,In_703,In_451);
nand U284 (N_284,In_403,In_685);
xnor U285 (N_285,In_939,In_495);
nor U286 (N_286,In_1400,In_248);
nor U287 (N_287,In_1311,In_1238);
and U288 (N_288,In_627,In_538);
or U289 (N_289,In_1454,In_786);
nand U290 (N_290,In_709,In_352);
nand U291 (N_291,In_301,In_1164);
nor U292 (N_292,In_1146,In_351);
or U293 (N_293,In_1413,In_534);
nor U294 (N_294,In_922,In_655);
nor U295 (N_295,In_1201,In_733);
xnor U296 (N_296,In_741,In_325);
nor U297 (N_297,In_553,In_402);
or U298 (N_298,In_978,In_755);
or U299 (N_299,In_948,In_1147);
nor U300 (N_300,In_661,In_20);
nor U301 (N_301,In_504,In_237);
nand U302 (N_302,In_360,In_540);
nand U303 (N_303,In_51,N_178);
nand U304 (N_304,In_1362,N_276);
nand U305 (N_305,In_427,In_609);
nor U306 (N_306,In_498,In_973);
or U307 (N_307,N_14,N_125);
and U308 (N_308,In_1056,In_596);
or U309 (N_309,In_1369,In_473);
or U310 (N_310,In_517,In_338);
nor U311 (N_311,In_992,In_228);
xor U312 (N_312,In_98,In_1366);
or U313 (N_313,N_71,N_288);
and U314 (N_314,In_971,In_614);
nor U315 (N_315,In_871,In_419);
and U316 (N_316,N_118,N_290);
or U317 (N_317,In_384,In_1353);
xor U318 (N_318,N_124,In_10);
nand U319 (N_319,In_573,N_11);
nand U320 (N_320,In_335,In_423);
and U321 (N_321,In_200,In_214);
nor U322 (N_322,N_271,In_789);
and U323 (N_323,N_291,N_130);
or U324 (N_324,In_920,In_224);
nor U325 (N_325,N_293,N_216);
nor U326 (N_326,In_1004,N_141);
xor U327 (N_327,In_707,N_281);
and U328 (N_328,In_1181,In_901);
or U329 (N_329,In_898,N_250);
xor U330 (N_330,In_1138,N_51);
or U331 (N_331,In_760,In_1486);
xnor U332 (N_332,In_848,In_670);
or U333 (N_333,In_598,In_1455);
nor U334 (N_334,In_392,In_82);
or U335 (N_335,N_5,N_227);
or U336 (N_336,In_268,In_1191);
nand U337 (N_337,In_1,In_1294);
or U338 (N_338,N_48,N_238);
and U339 (N_339,In_662,In_606);
or U340 (N_340,In_542,In_539);
nor U341 (N_341,In_582,N_136);
nor U342 (N_342,In_1491,In_410);
nor U343 (N_343,In_188,N_12);
and U344 (N_344,N_286,In_60);
xor U345 (N_345,In_688,In_1440);
or U346 (N_346,In_803,In_1378);
or U347 (N_347,In_363,In_202);
nor U348 (N_348,In_804,In_957);
nand U349 (N_349,N_80,In_242);
nand U350 (N_350,In_1423,N_93);
and U351 (N_351,N_228,In_154);
nor U352 (N_352,In_230,In_852);
nor U353 (N_353,N_195,N_129);
or U354 (N_354,In_1318,In_1415);
nand U355 (N_355,In_572,N_230);
and U356 (N_356,In_1352,In_1034);
nor U357 (N_357,In_176,In_465);
nor U358 (N_358,In_1104,In_221);
nor U359 (N_359,In_347,In_1479);
xnor U360 (N_360,In_454,N_89);
and U361 (N_361,In_488,In_1125);
and U362 (N_362,In_796,N_100);
or U363 (N_363,In_577,N_188);
or U364 (N_364,In_523,In_580);
and U365 (N_365,In_1282,In_1267);
and U366 (N_366,In_514,In_717);
nand U367 (N_367,In_692,In_776);
nor U368 (N_368,In_1160,N_32);
xor U369 (N_369,N_215,In_546);
nor U370 (N_370,In_1443,In_604);
or U371 (N_371,In_1336,N_10);
or U372 (N_372,In_1340,N_255);
nor U373 (N_373,N_69,In_1089);
and U374 (N_374,In_1126,In_1124);
and U375 (N_375,In_705,In_494);
nand U376 (N_376,In_533,In_990);
nand U377 (N_377,In_468,In_775);
and U378 (N_378,In_695,In_1043);
xor U379 (N_379,In_59,In_425);
and U380 (N_380,N_8,In_1330);
nand U381 (N_381,In_27,In_492);
nor U382 (N_382,In_267,In_597);
or U383 (N_383,In_861,In_911);
nand U384 (N_384,In_138,In_892);
xor U385 (N_385,In_111,N_233);
and U386 (N_386,N_161,In_1475);
nor U387 (N_387,In_535,In_1020);
xor U388 (N_388,N_277,N_85);
xor U389 (N_389,In_763,In_846);
and U390 (N_390,N_191,N_76);
and U391 (N_391,N_19,In_222);
or U392 (N_392,In_1193,In_1350);
nor U393 (N_393,N_177,N_119);
xnor U394 (N_394,In_118,N_122);
xor U395 (N_395,In_1021,In_253);
or U396 (N_396,N_23,In_12);
nor U397 (N_397,In_501,N_61);
nor U398 (N_398,N_194,In_459);
and U399 (N_399,N_131,In_151);
nor U400 (N_400,In_1496,In_879);
xor U401 (N_401,In_1149,In_1105);
and U402 (N_402,In_886,In_1472);
nor U403 (N_403,N_169,In_982);
xnor U404 (N_404,In_1490,In_408);
or U405 (N_405,In_874,In_1075);
and U406 (N_406,In_771,In_1136);
nor U407 (N_407,In_1477,N_183);
or U408 (N_408,In_891,In_985);
or U409 (N_409,N_289,In_64);
nand U410 (N_410,In_1281,In_303);
and U411 (N_411,In_297,In_1292);
or U412 (N_412,In_437,In_1202);
nand U413 (N_413,In_562,In_1206);
xnor U414 (N_414,In_116,In_748);
nor U415 (N_415,In_1450,N_59);
or U416 (N_416,In_235,In_296);
nand U417 (N_417,In_933,In_293);
nand U418 (N_418,In_496,In_529);
xnor U419 (N_419,In_668,N_202);
and U420 (N_420,N_236,In_13);
nand U421 (N_421,In_1062,In_1019);
xor U422 (N_422,N_180,In_1094);
or U423 (N_423,N_214,In_1182);
nand U424 (N_424,In_1040,In_1036);
and U425 (N_425,In_485,In_829);
nand U426 (N_426,N_207,In_570);
nand U427 (N_427,In_1289,In_1084);
or U428 (N_428,In_824,N_152);
xnor U429 (N_429,In_166,In_1255);
or U430 (N_430,In_554,In_612);
xor U431 (N_431,N_273,In_1424);
nor U432 (N_432,In_467,In_16);
and U433 (N_433,In_758,In_835);
and U434 (N_434,N_81,In_1351);
nand U435 (N_435,In_1493,In_1106);
nand U436 (N_436,N_105,N_234);
and U437 (N_437,In_651,N_231);
and U438 (N_438,In_968,In_945);
and U439 (N_439,In_282,In_1390);
or U440 (N_440,In_39,In_499);
nor U441 (N_441,In_172,In_182);
nand U442 (N_442,In_507,In_136);
and U443 (N_443,In_122,In_270);
nand U444 (N_444,N_40,In_1391);
nor U445 (N_445,In_330,In_958);
nand U446 (N_446,In_1247,In_541);
or U447 (N_447,In_401,In_1407);
and U448 (N_448,In_3,In_1224);
or U449 (N_449,In_1426,N_137);
nand U450 (N_450,N_212,In_1306);
xnor U451 (N_451,N_13,In_738);
and U452 (N_452,In_432,N_21);
and U453 (N_453,N_116,In_545);
and U454 (N_454,In_863,N_218);
nand U455 (N_455,In_1291,In_794);
or U456 (N_456,In_884,In_1368);
and U457 (N_457,In_164,In_1499);
or U458 (N_458,In_1190,In_537);
and U459 (N_459,N_78,In_319);
xor U460 (N_460,In_1025,In_1372);
nand U461 (N_461,In_1253,In_1207);
xor U462 (N_462,N_172,In_938);
xnor U463 (N_463,In_851,In_1494);
and U464 (N_464,N_206,In_676);
and U465 (N_465,In_808,In_1243);
or U466 (N_466,In_1334,In_620);
or U467 (N_467,In_980,In_770);
nor U468 (N_468,N_242,N_166);
nand U469 (N_469,In_1457,N_251);
xor U470 (N_470,In_677,In_81);
xor U471 (N_471,In_790,In_792);
xnor U472 (N_472,In_1001,In_1488);
xnor U473 (N_473,In_1184,N_33);
nand U474 (N_474,In_532,In_1236);
nor U475 (N_475,N_140,In_1307);
xor U476 (N_476,In_226,In_1429);
xor U477 (N_477,In_204,N_237);
nor U478 (N_478,In_1271,In_287);
nand U479 (N_479,In_513,In_152);
xnor U480 (N_480,N_147,In_905);
nand U481 (N_481,N_65,In_1035);
and U482 (N_482,N_88,In_344);
nor U483 (N_483,In_203,In_420);
nor U484 (N_484,N_60,In_1405);
and U485 (N_485,In_90,In_977);
or U486 (N_486,In_1492,In_1167);
nand U487 (N_487,N_107,In_149);
nor U488 (N_488,N_246,In_120);
xor U489 (N_489,In_1048,In_1392);
nand U490 (N_490,In_601,In_626);
nand U491 (N_491,In_566,In_1028);
nand U492 (N_492,N_224,In_160);
nand U493 (N_493,N_150,In_768);
xnor U494 (N_494,In_947,N_75);
nand U495 (N_495,In_578,In_1339);
nor U496 (N_496,In_53,In_887);
nand U497 (N_497,In_80,In_1151);
or U498 (N_498,In_897,In_551);
or U499 (N_499,N_144,In_1076);
xnor U500 (N_500,In_1248,In_1296);
or U501 (N_501,In_942,In_1270);
nor U502 (N_502,N_175,In_1142);
nand U503 (N_503,In_1130,In_1099);
or U504 (N_504,In_921,N_187);
nand U505 (N_505,In_411,In_483);
xnor U506 (N_506,N_46,In_889);
xnor U507 (N_507,In_104,In_1262);
and U508 (N_508,N_92,In_1172);
nor U509 (N_509,In_561,N_52);
and U510 (N_510,In_1333,In_781);
or U511 (N_511,In_1176,In_96);
and U512 (N_512,N_36,In_762);
or U513 (N_513,N_163,In_1463);
xnor U514 (N_514,In_373,In_961);
or U515 (N_515,In_1003,In_774);
nand U516 (N_516,In_342,In_1497);
xor U517 (N_517,N_261,In_780);
xor U518 (N_518,N_278,N_197);
xor U519 (N_519,N_44,In_1439);
nand U520 (N_520,In_274,In_899);
nor U521 (N_521,In_986,In_563);
nor U522 (N_522,In_646,In_161);
and U523 (N_523,N_205,N_196);
and U524 (N_524,In_1425,N_292);
or U525 (N_525,In_341,In_290);
or U526 (N_526,In_1067,In_979);
nor U527 (N_527,In_475,In_174);
xor U528 (N_528,N_26,N_297);
and U529 (N_529,In_489,N_258);
xnor U530 (N_530,In_1285,In_223);
and U531 (N_531,N_174,In_240);
and U532 (N_532,N_274,In_923);
nand U533 (N_533,In_716,N_192);
nand U534 (N_534,N_22,N_156);
nand U535 (N_535,N_20,In_1464);
xnor U536 (N_536,N_86,In_349);
nor U537 (N_537,N_266,In_1380);
and U538 (N_538,In_568,In_751);
or U539 (N_539,In_447,N_115);
and U540 (N_540,N_82,In_305);
nor U541 (N_541,In_216,In_159);
or U542 (N_542,N_24,N_28);
nor U543 (N_543,In_660,In_1397);
or U544 (N_544,In_600,In_103);
nor U545 (N_545,N_138,N_17);
nand U546 (N_546,N_6,In_1222);
nand U547 (N_547,In_1030,N_134);
and U548 (N_548,In_1459,N_295);
xor U549 (N_549,In_156,In_687);
nor U550 (N_550,In_903,In_107);
or U551 (N_551,In_1038,N_133);
or U552 (N_552,In_6,In_124);
and U553 (N_553,In_44,In_953);
nand U554 (N_554,In_1212,In_482);
xor U555 (N_555,In_1008,In_1304);
xor U556 (N_556,In_1326,In_502);
and U557 (N_557,N_185,N_248);
nor U558 (N_558,In_434,In_723);
nand U559 (N_559,In_441,N_126);
xnor U560 (N_560,In_123,In_309);
or U561 (N_561,In_1460,In_571);
nor U562 (N_562,In_439,N_182);
or U563 (N_563,N_111,In_171);
xnor U564 (N_564,In_78,In_37);
nor U565 (N_565,In_348,N_58);
and U566 (N_566,In_336,N_57);
nand U567 (N_567,In_1422,N_222);
or U568 (N_568,In_1077,In_1134);
nand U569 (N_569,In_370,In_30);
nand U570 (N_570,N_123,N_135);
or U571 (N_571,In_246,In_472);
or U572 (N_572,In_1482,In_1183);
nand U573 (N_573,In_1024,In_1447);
nor U574 (N_574,In_1127,In_735);
nor U575 (N_575,In_510,N_148);
and U576 (N_576,In_25,In_1209);
or U577 (N_577,In_184,In_969);
and U578 (N_578,In_1017,In_358);
or U579 (N_579,N_56,In_860);
or U580 (N_580,In_1297,In_1382);
or U581 (N_581,N_62,In_729);
and U582 (N_582,In_654,In_311);
and U583 (N_583,In_1302,In_1495);
nor U584 (N_584,In_1328,N_171);
nand U585 (N_585,N_9,In_254);
or U586 (N_586,In_1109,In_611);
or U587 (N_587,In_1483,In_1341);
or U588 (N_588,In_1438,In_1431);
and U589 (N_589,N_299,In_35);
xor U590 (N_590,In_327,In_764);
and U591 (N_591,In_788,In_1468);
or U592 (N_592,In_249,In_934);
nand U593 (N_593,In_890,In_959);
nor U594 (N_594,In_809,In_914);
nor U595 (N_595,In_312,In_996);
nor U596 (N_596,In_1283,In_956);
xor U597 (N_597,In_1000,In_800);
or U598 (N_598,In_1252,In_100);
xnor U599 (N_599,In_478,In_1485);
nand U600 (N_600,In_1256,N_265);
nand U601 (N_601,N_260,N_0);
or U602 (N_602,N_524,N_326);
or U603 (N_603,N_302,N_419);
xnor U604 (N_604,N_181,N_508);
xor U605 (N_605,N_492,N_318);
or U606 (N_606,N_547,N_439);
or U607 (N_607,In_1046,N_72);
nor U608 (N_608,In_68,N_155);
or U609 (N_609,In_294,N_256);
and U610 (N_610,In_381,In_436);
xor U611 (N_611,In_49,In_443);
nand U612 (N_612,In_388,In_40);
xor U613 (N_613,In_213,In_1192);
or U614 (N_614,N_429,N_262);
or U615 (N_615,N_298,N_398);
and U616 (N_616,In_1060,N_572);
xnor U617 (N_617,In_711,In_1406);
xnor U618 (N_618,In_1052,N_414);
or U619 (N_619,N_168,In_422);
nand U620 (N_620,In_1363,N_356);
nor U621 (N_621,In_1388,N_153);
nand U622 (N_622,In_669,In_1171);
xor U623 (N_623,N_505,N_406);
or U624 (N_624,N_219,In_283);
xnor U625 (N_625,In_66,N_384);
xor U626 (N_626,N_580,N_388);
and U627 (N_627,In_1419,In_455);
nor U628 (N_628,In_1452,N_353);
or U629 (N_629,N_327,In_170);
nor U630 (N_630,N_461,N_385);
or U631 (N_631,N_25,In_258);
xnor U632 (N_632,In_1441,In_998);
and U633 (N_633,N_294,In_1114);
and U634 (N_634,In_430,In_633);
and U635 (N_635,In_555,N_403);
nand U636 (N_636,N_370,In_1257);
nor U637 (N_637,N_466,N_583);
nor U638 (N_638,In_559,In_850);
nor U639 (N_639,N_300,In_617);
or U640 (N_640,In_131,In_1066);
nand U641 (N_641,N_362,N_335);
nor U642 (N_642,N_373,N_452);
or U643 (N_643,In_14,In_1343);
or U644 (N_644,In_569,N_139);
nor U645 (N_645,In_881,In_1139);
and U646 (N_646,In_1331,N_142);
nand U647 (N_647,In_516,N_106);
nand U648 (N_648,N_500,In_665);
or U649 (N_649,In_210,N_267);
xor U650 (N_650,N_90,N_512);
nand U651 (N_651,In_1320,N_533);
or U652 (N_652,In_806,N_441);
or U653 (N_653,N_368,In_772);
and U654 (N_654,In_1137,In_799);
and U655 (N_655,N_18,N_426);
or U656 (N_656,N_425,In_619);
or U657 (N_657,In_1384,In_906);
nand U658 (N_658,In_354,In_117);
or U659 (N_659,N_597,In_481);
nand U660 (N_660,N_390,N_573);
or U661 (N_661,In_1416,N_471);
or U662 (N_662,N_540,In_991);
and U663 (N_663,In_1220,N_74);
xor U664 (N_664,N_45,N_495);
and U665 (N_665,N_574,In_464);
nand U666 (N_666,In_225,In_856);
and U667 (N_667,In_448,N_363);
nand U668 (N_668,In_650,In_189);
xor U669 (N_669,In_121,In_1122);
nand U670 (N_670,N_201,N_176);
nor U671 (N_671,N_469,N_316);
xnor U672 (N_672,In_395,N_436);
nor U673 (N_673,N_528,In_917);
nor U674 (N_674,N_167,N_558);
nand U675 (N_675,In_731,N_438);
nor U676 (N_676,N_313,N_254);
nand U677 (N_677,N_321,In_289);
xnor U678 (N_678,In_318,In_359);
xor U679 (N_679,In_209,In_185);
and U680 (N_680,N_341,In_767);
or U681 (N_681,N_275,N_428);
xor U682 (N_682,N_504,In_1461);
xnor U683 (N_683,N_454,N_585);
nor U684 (N_684,In_742,In_1121);
and U685 (N_685,In_458,In_281);
nor U686 (N_686,In_1462,In_238);
or U687 (N_687,In_801,N_98);
xor U688 (N_688,In_1153,N_520);
nor U689 (N_689,In_382,In_1203);
xor U690 (N_690,N_322,In_1013);
or U691 (N_691,N_15,N_1);
nand U692 (N_692,N_104,N_151);
xor U693 (N_693,In_406,In_1031);
and U694 (N_694,In_802,In_462);
and U695 (N_695,In_644,N_479);
nand U696 (N_696,N_411,In_1474);
nand U697 (N_697,In_699,N_445);
xor U698 (N_698,In_1006,N_483);
or U699 (N_699,In_704,N_494);
nor U700 (N_700,N_349,N_184);
or U701 (N_701,In_659,N_41);
nor U702 (N_702,N_367,In_115);
xor U703 (N_703,N_448,In_1395);
or U704 (N_704,In_477,In_1165);
nand U705 (N_705,N_355,In_679);
nand U706 (N_706,In_782,In_133);
nor U707 (N_707,N_463,In_522);
or U708 (N_708,N_446,N_225);
or U709 (N_709,In_1015,N_412);
and U710 (N_710,N_314,N_350);
and U711 (N_711,In_987,In_367);
nand U712 (N_712,In_497,N_4);
nand U713 (N_713,N_323,N_268);
nor U714 (N_714,N_339,N_331);
nand U715 (N_715,In_721,In_591);
or U716 (N_716,N_239,N_259);
nor U717 (N_717,N_121,N_164);
and U718 (N_718,N_29,N_507);
and U719 (N_719,In_1393,In_528);
nor U720 (N_720,N_409,In_584);
or U721 (N_721,N_444,N_592);
nand U722 (N_722,N_241,In_1273);
or U723 (N_723,In_680,N_455);
nand U724 (N_724,In_183,In_1229);
and U725 (N_725,N_543,N_484);
xor U726 (N_726,In_1430,In_581);
nand U727 (N_727,N_513,In_678);
nor U728 (N_728,In_1133,N_465);
nor U729 (N_729,N_47,In_1251);
nand U730 (N_730,In_190,In_28);
xor U731 (N_731,N_37,In_92);
or U732 (N_732,N_159,In_1258);
or U733 (N_733,In_7,N_537);
nand U734 (N_734,In_1387,N_591);
nand U735 (N_735,In_332,In_1055);
or U736 (N_736,N_488,N_158);
xor U737 (N_737,N_73,N_407);
and U738 (N_738,N_145,N_491);
nand U739 (N_739,In_833,N_599);
or U740 (N_740,In_1120,In_1175);
or U741 (N_741,N_359,In_1305);
xnor U742 (N_742,N_79,N_306);
or U743 (N_743,N_381,N_401);
xor U744 (N_744,In_1347,In_928);
and U745 (N_745,N_343,N_315);
and U746 (N_746,In_1232,In_1095);
xnor U747 (N_747,In_1383,In_292);
xnor U748 (N_748,In_24,In_193);
or U749 (N_749,In_766,N_522);
and U750 (N_750,In_1068,In_196);
or U751 (N_751,N_514,N_393);
and U752 (N_752,N_154,N_269);
nor U753 (N_753,In_1411,N_394);
and U754 (N_754,In_1371,In_1178);
and U755 (N_755,N_336,N_581);
or U756 (N_756,N_475,In_1259);
nor U757 (N_757,N_397,In_575);
and U758 (N_758,In_838,In_1287);
xor U759 (N_759,In_1370,N_35);
nor U760 (N_760,In_460,N_542);
xor U761 (N_761,N_351,In_484);
xnor U762 (N_762,In_1074,In_1338);
xor U763 (N_763,In_1179,In_1129);
xnor U764 (N_764,N_480,In_1166);
nor U765 (N_765,N_348,In_339);
nor U766 (N_766,In_394,N_563);
nor U767 (N_767,N_304,N_213);
or U768 (N_768,N_595,N_54);
nor U769 (N_769,N_173,In_883);
nor U770 (N_770,In_1239,N_517);
nand U771 (N_771,N_527,N_186);
nand U772 (N_772,N_413,N_422);
and U773 (N_773,In_298,N_460);
or U774 (N_774,N_282,N_423);
or U775 (N_775,In_918,N_375);
or U776 (N_776,N_30,In_929);
and U777 (N_777,In_926,N_301);
nor U778 (N_778,In_549,In_167);
or U779 (N_779,In_1082,In_844);
nor U780 (N_780,In_1346,In_1458);
and U781 (N_781,N_204,In_628);
and U782 (N_782,N_519,N_538);
and U783 (N_783,In_162,In_1432);
xor U784 (N_784,In_1044,In_1379);
or U785 (N_785,N_270,N_328);
nand U786 (N_786,N_498,In_364);
nor U787 (N_787,In_805,N_165);
nand U788 (N_788,N_473,In_1170);
nand U789 (N_789,N_143,N_424);
nor U790 (N_790,In_326,In_924);
nand U791 (N_791,N_437,In_173);
nor U792 (N_792,In_1402,N_497);
xor U793 (N_793,N_550,N_99);
nand U794 (N_794,N_420,N_506);
nand U795 (N_795,In_493,In_317);
nor U796 (N_796,N_489,In_621);
or U797 (N_797,N_374,N_312);
or U798 (N_798,In_331,N_561);
nand U799 (N_799,N_55,In_995);
xor U800 (N_800,In_544,N_101);
xnor U801 (N_801,N_50,In_474);
nor U802 (N_802,In_1263,In_1101);
xnor U803 (N_803,In_322,N_244);
nand U804 (N_804,In_128,In_506);
and U805 (N_805,In_450,N_579);
and U806 (N_806,N_120,In_1086);
nor U807 (N_807,N_53,N_94);
or U808 (N_808,In_211,N_383);
nor U809 (N_809,N_544,N_557);
xnor U810 (N_810,In_1357,In_207);
or U811 (N_811,N_576,N_346);
xor U812 (N_812,N_459,In_1032);
or U813 (N_813,N_366,N_462);
nand U814 (N_814,N_577,In_393);
and U815 (N_815,In_525,N_203);
and U816 (N_816,N_582,In_1436);
nand U817 (N_817,N_70,N_354);
or U818 (N_818,In_139,In_463);
xor U819 (N_819,In_5,N_545);
nand U820 (N_820,In_512,In_85);
or U821 (N_821,N_486,In_135);
xnor U822 (N_822,N_376,In_1216);
or U823 (N_823,In_1026,In_925);
or U824 (N_824,In_110,In_1174);
nand U825 (N_825,N_127,N_249);
nand U826 (N_826,N_496,N_96);
nor U827 (N_827,In_163,In_257);
nor U828 (N_828,In_931,In_1049);
nor U829 (N_829,N_31,N_307);
nand U830 (N_830,In_1169,N_369);
and U831 (N_831,In_1228,In_1214);
or U832 (N_832,In_595,N_467);
or U833 (N_833,In_1317,N_208);
xor U834 (N_834,In_1377,N_539);
nand U835 (N_835,N_95,N_458);
or U836 (N_836,N_232,N_554);
or U837 (N_837,N_361,N_332);
and U838 (N_838,In_1356,N_320);
nor U839 (N_839,N_481,In_876);
and U840 (N_840,In_1360,N_211);
or U841 (N_841,N_108,N_113);
xor U842 (N_842,In_734,N_552);
and U843 (N_843,In_888,In_1111);
and U844 (N_844,N_503,In_1312);
and U845 (N_845,In_658,N_499);
nand U846 (N_846,In_1465,N_487);
and U847 (N_847,In_405,In_1218);
and U848 (N_848,In_134,N_477);
xor U849 (N_849,In_1240,N_310);
and U850 (N_850,N_38,N_146);
xor U851 (N_851,In_490,N_372);
or U852 (N_852,N_3,In_1444);
nand U853 (N_853,In_752,In_684);
xnor U854 (N_854,N_400,In_813);
nor U855 (N_855,In_869,N_179);
nand U856 (N_856,N_360,N_296);
nor U857 (N_857,N_365,In_1313);
or U858 (N_858,N_114,In_916);
nand U859 (N_859,N_226,N_405);
nor U860 (N_860,In_857,N_590);
xor U861 (N_861,In_1471,In_902);
and U862 (N_862,N_567,In_1349);
and U863 (N_863,N_162,In_1211);
and U864 (N_864,In_1116,N_170);
xor U865 (N_865,N_117,In_75);
and U866 (N_866,N_396,In_783);
nor U867 (N_867,N_556,N_91);
xor U868 (N_868,In_195,N_565);
nor U869 (N_869,N_243,N_570);
xnor U870 (N_870,In_65,In_375);
nand U871 (N_871,N_272,In_940);
or U872 (N_872,N_209,In_105);
nor U873 (N_873,In_1208,In_588);
nand U874 (N_874,In_1069,In_882);
xnor U875 (N_875,N_518,In_649);
or U876 (N_876,In_589,In_409);
xor U877 (N_877,N_482,N_235);
and U878 (N_878,In_900,In_558);
and U879 (N_879,N_402,N_253);
nand U880 (N_880,N_2,N_283);
nand U881 (N_881,N_377,In_822);
nor U882 (N_882,In_1059,N_378);
xnor U883 (N_883,N_569,In_142);
or U884 (N_884,N_279,In_150);
nor U885 (N_885,N_472,N_523);
nor U886 (N_886,In_54,In_407);
and U887 (N_887,In_618,N_575);
and U888 (N_888,In_328,N_66);
xor U889 (N_889,N_280,In_520);
and U890 (N_890,In_954,In_634);
xor U891 (N_891,N_352,In_630);
xor U892 (N_892,In_1373,In_1274);
and U893 (N_893,N_77,N_220);
xor U894 (N_894,In_667,In_255);
nor U895 (N_895,N_84,N_546);
and U896 (N_896,N_303,In_515);
xor U897 (N_897,In_1246,N_526);
xnor U898 (N_898,N_223,N_109);
or U899 (N_899,In_732,In_456);
nor U900 (N_900,N_864,N_535);
nor U901 (N_901,N_868,N_662);
or U902 (N_902,N_898,N_347);
nor U903 (N_903,N_609,In_414);
nand U904 (N_904,N_638,N_653);
and U905 (N_905,N_594,N_417);
and U906 (N_906,N_719,N_680);
xnor U907 (N_907,N_760,In_547);
nor U908 (N_908,N_284,N_193);
or U909 (N_909,N_391,N_689);
nor U910 (N_910,N_845,In_993);
nor U911 (N_911,N_872,N_765);
nor U912 (N_912,N_836,N_835);
xnor U913 (N_913,N_604,In_1161);
or U914 (N_914,N_309,In_205);
and U915 (N_915,N_705,N_773);
or U916 (N_916,N_571,N_726);
and U917 (N_917,N_668,In_1449);
nand U918 (N_918,N_834,In_773);
nand U919 (N_919,N_800,N_785);
or U920 (N_920,N_735,N_431);
xor U921 (N_921,N_641,In_653);
nor U922 (N_922,N_839,N_379);
xor U923 (N_923,N_64,N_852);
nand U924 (N_924,In_1481,In_109);
xnor U925 (N_925,N_549,N_882);
nor U926 (N_926,N_617,N_763);
or U927 (N_927,N_470,N_799);
nor U928 (N_928,N_588,N_796);
nand U929 (N_929,N_600,N_686);
and U930 (N_930,In_74,N_718);
nor U931 (N_931,N_623,In_1280);
or U932 (N_932,N_564,In_1117);
or U933 (N_933,N_762,N_697);
nor U934 (N_934,N_704,N_530);
and U935 (N_935,N_871,N_826);
xor U936 (N_936,N_478,In_372);
or U937 (N_937,In_657,N_817);
nand U938 (N_938,N_245,N_677);
or U939 (N_939,N_587,N_622);
or U940 (N_940,In_759,N_649);
xnor U941 (N_941,In_446,N_319);
nand U942 (N_942,N_430,N_639);
xnor U943 (N_943,N_778,N_642);
nor U944 (N_944,N_707,N_324);
and U945 (N_945,In_1163,N_859);
nor U946 (N_946,In_148,N_770);
xor U947 (N_947,N_456,N_692);
nor U948 (N_948,N_627,N_700);
nand U949 (N_949,N_750,In_1065);
or U950 (N_950,N_476,N_781);
nand U951 (N_951,N_666,In_1286);
or U952 (N_952,In_55,N_759);
nor U953 (N_953,In_1476,In_1197);
and U954 (N_954,In_1041,N_775);
nor U955 (N_955,N_645,N_801);
nor U956 (N_956,In_1446,N_317);
nor U957 (N_957,N_855,N_43);
and U958 (N_958,N_337,N_618);
nor U959 (N_959,In_1081,N_364);
nor U960 (N_960,N_338,N_667);
and U961 (N_961,N_710,In_45);
nand U962 (N_962,N_749,N_815);
nor U963 (N_963,In_390,N_721);
nand U964 (N_964,N_34,N_634);
and U965 (N_965,In_1484,N_883);
and U966 (N_966,N_730,N_633);
or U967 (N_967,N_240,N_416);
xor U968 (N_968,N_779,N_709);
nand U969 (N_969,N_657,N_695);
nor U970 (N_970,N_637,N_804);
nor U971 (N_971,N_305,N_867);
nor U972 (N_972,N_701,In_638);
xor U973 (N_973,N_808,N_646);
nand U974 (N_974,N_688,N_440);
xnor U975 (N_975,N_399,N_786);
nor U976 (N_976,N_807,In_1156);
xor U977 (N_977,N_83,N_578);
xnor U978 (N_978,N_596,N_714);
nor U979 (N_979,N_584,N_899);
nand U980 (N_980,In_1272,N_189);
nor U981 (N_981,N_757,In_1434);
and U982 (N_982,N_862,N_768);
nand U983 (N_983,N_717,N_607);
xor U984 (N_984,In_1277,In_1375);
and U985 (N_985,N_602,N_102);
xnor U986 (N_986,N_389,N_553);
xor U987 (N_987,N_650,In_641);
nor U988 (N_988,N_837,N_708);
or U989 (N_989,In_1234,In_1150);
or U990 (N_990,N_683,N_515);
nor U991 (N_991,N_751,N_678);
nand U992 (N_992,In_1389,In_843);
and U993 (N_993,In_521,In_378);
xnor U994 (N_994,In_1204,N_342);
xnor U995 (N_995,N_865,N_856);
nand U996 (N_996,In_970,N_629);
nor U997 (N_997,N_157,In_280);
or U998 (N_998,N_731,N_534);
xor U999 (N_999,N_725,N_611);
nand U1000 (N_1000,N_656,N_453);
nor U1001 (N_1001,In_648,In_828);
nand U1002 (N_1002,N_247,N_742);
or U1003 (N_1003,In_1325,N_605);
xor U1004 (N_1004,N_783,N_769);
xnor U1005 (N_1005,N_880,In_112);
nor U1006 (N_1006,N_386,In_909);
and U1007 (N_1007,N_715,N_380);
nand U1008 (N_1008,N_712,In_426);
or U1009 (N_1009,In_1399,N_747);
or U1010 (N_1010,N_614,N_874);
xnor U1011 (N_1011,N_792,N_263);
and U1012 (N_1012,N_788,N_805);
or U1013 (N_1013,N_652,N_635);
xnor U1014 (N_1014,N_674,N_879);
nand U1015 (N_1015,N_625,N_711);
and U1016 (N_1016,In_429,N_198);
or U1017 (N_1017,N_501,N_696);
nand U1018 (N_1018,N_675,N_643);
and U1019 (N_1019,N_408,N_511);
xor U1020 (N_1020,N_598,N_851);
or U1021 (N_1021,N_693,In_1348);
or U1022 (N_1022,N_777,N_744);
or U1023 (N_1023,N_387,N_825);
nor U1024 (N_1024,N_824,In_682);
nor U1025 (N_1025,In_1018,N_340);
xnor U1026 (N_1026,N_87,In_491);
xnor U1027 (N_1027,N_264,N_525);
and U1028 (N_1028,In_1180,In_702);
or U1029 (N_1029,N_887,N_229);
or U1030 (N_1030,N_418,N_764);
nand U1031 (N_1031,N_885,In_273);
nand U1032 (N_1032,N_610,In_1489);
nand U1033 (N_1033,N_654,N_648);
xor U1034 (N_1034,N_630,N_149);
nand U1035 (N_1035,N_766,N_325);
nor U1036 (N_1036,N_427,N_217);
and U1037 (N_1037,In_1396,In_299);
or U1038 (N_1038,N_128,N_897);
or U1039 (N_1039,N_702,N_626);
xor U1040 (N_1040,In_912,N_866);
or U1041 (N_1041,N_628,N_811);
nand U1042 (N_1042,N_754,N_42);
xnor U1043 (N_1043,In_700,N_892);
or U1044 (N_1044,N_63,In_320);
and U1045 (N_1045,N_694,N_823);
nor U1046 (N_1046,N_432,In_21);
xnor U1047 (N_1047,N_698,N_644);
and U1048 (N_1048,In_964,N_822);
and U1049 (N_1049,N_690,In_201);
or U1050 (N_1050,In_725,N_809);
nor U1051 (N_1051,In_754,N_740);
nand U1052 (N_1052,N_112,N_464);
or U1053 (N_1053,In_442,N_849);
nor U1054 (N_1054,N_457,N_451);
or U1055 (N_1055,N_311,N_110);
xor U1056 (N_1056,N_661,N_782);
xnor U1057 (N_1057,In_590,N_371);
nor U1058 (N_1058,In_698,N_889);
xor U1059 (N_1059,In_1480,In_245);
or U1060 (N_1060,N_850,N_392);
or U1061 (N_1061,N_329,N_531);
xnor U1062 (N_1062,N_404,N_741);
and U1063 (N_1063,N_593,N_847);
or U1064 (N_1064,N_893,N_676);
nand U1065 (N_1065,N_703,N_612);
nor U1066 (N_1066,N_555,In_1337);
nor U1067 (N_1067,N_738,In_1011);
nand U1068 (N_1068,N_97,N_842);
and U1069 (N_1069,N_877,In_715);
xor U1070 (N_1070,In_126,In_340);
nor U1071 (N_1071,In_71,In_1324);
nor U1072 (N_1072,N_210,In_526);
xnor U1073 (N_1073,In_1016,N_447);
or U1074 (N_1074,N_797,N_344);
nor U1075 (N_1075,N_357,N_664);
xor U1076 (N_1076,N_761,N_257);
nand U1077 (N_1077,N_831,N_789);
nor U1078 (N_1078,N_636,In_404);
nand U1079 (N_1079,In_681,N_443);
nand U1080 (N_1080,N_891,N_673);
xnor U1081 (N_1081,N_806,N_886);
xor U1082 (N_1082,In_1185,In_141);
xor U1083 (N_1083,N_888,In_158);
nand U1084 (N_1084,In_272,N_621);
nand U1085 (N_1085,N_658,N_562);
nor U1086 (N_1086,N_651,N_795);
and U1087 (N_1087,N_631,In_315);
or U1088 (N_1088,N_632,N_521);
xnor U1089 (N_1089,In_194,In_983);
xnor U1090 (N_1090,N_780,N_529);
nor U1091 (N_1091,N_39,N_890);
nor U1092 (N_1092,N_616,N_827);
and U1093 (N_1093,N_532,N_723);
nor U1094 (N_1094,N_873,N_728);
xnor U1095 (N_1095,N_881,N_624);
nand U1096 (N_1096,N_619,N_790);
nor U1097 (N_1097,N_821,In_108);
or U1098 (N_1098,N_669,N_568);
or U1099 (N_1099,N_132,In_1045);
nor U1100 (N_1100,N_49,N_833);
or U1101 (N_1101,N_510,N_857);
nor U1102 (N_1102,N_358,In_1381);
nand U1103 (N_1103,N_659,N_793);
nand U1104 (N_1104,N_415,N_794);
nor U1105 (N_1105,In_893,N_287);
or U1106 (N_1106,N_840,In_1215);
and U1107 (N_1107,N_813,N_103);
nand U1108 (N_1108,N_832,In_1456);
or U1109 (N_1109,N_671,N_748);
or U1110 (N_1110,N_753,In_1421);
xor U1111 (N_1111,N_767,N_812);
and U1112 (N_1112,N_685,N_308);
and U1113 (N_1113,N_190,N_737);
nor U1114 (N_1114,N_756,N_200);
xor U1115 (N_1115,N_687,N_27);
nor U1116 (N_1116,N_16,N_860);
nor U1117 (N_1117,N_606,In_231);
and U1118 (N_1118,In_180,N_724);
nor U1119 (N_1119,In_22,N_559);
nor U1120 (N_1120,N_752,In_1168);
and U1121 (N_1121,N_199,In_91);
xor U1122 (N_1122,N_672,N_435);
or U1123 (N_1123,In_130,In_952);
xnor U1124 (N_1124,N_803,N_802);
nor U1125 (N_1125,N_876,N_691);
nand U1126 (N_1126,In_787,N_334);
or U1127 (N_1127,N_818,N_665);
or U1128 (N_1128,N_449,In_374);
and U1129 (N_1129,In_440,N_670);
nor U1130 (N_1130,In_1070,N_516);
or U1131 (N_1131,N_679,N_450);
or U1132 (N_1132,N_771,N_828);
or U1133 (N_1133,N_7,N_878);
xor U1134 (N_1134,N_894,N_729);
nor U1135 (N_1135,N_734,N_716);
or U1136 (N_1136,N_589,N_681);
xor U1137 (N_1137,N_682,N_784);
xnor U1138 (N_1138,In_1316,N_746);
xnor U1139 (N_1139,N_442,N_858);
and U1140 (N_1140,N_869,N_838);
xnor U1141 (N_1141,N_896,In_656);
nand U1142 (N_1142,In_70,In_720);
or U1143 (N_1143,In_87,In_999);
and U1144 (N_1144,N_755,N_330);
nand U1145 (N_1145,N_660,N_684);
nand U1146 (N_1146,N_502,N_787);
nand U1147 (N_1147,N_745,In_220);
nand U1148 (N_1148,N_608,N_541);
and U1149 (N_1149,N_791,In_480);
and U1150 (N_1150,In_1115,In_736);
xor U1151 (N_1151,N_382,In_186);
nor U1152 (N_1152,In_1029,N_884);
nor U1153 (N_1153,N_551,N_67);
or U1154 (N_1154,N_841,N_68);
or U1155 (N_1155,In_1298,N_743);
nor U1156 (N_1156,N_816,In_635);
nor U1157 (N_1157,In_466,N_820);
nand U1158 (N_1158,N_814,N_663);
xor U1159 (N_1159,N_720,N_560);
nand U1160 (N_1160,N_733,N_474);
or U1161 (N_1161,In_984,In_77);
nor U1162 (N_1162,N_706,N_221);
nand U1163 (N_1163,N_732,In_1453);
xnor U1164 (N_1164,N_798,N_485);
nor U1165 (N_1165,N_846,In_227);
and U1166 (N_1166,In_1365,N_875);
nand U1167 (N_1167,N_810,N_699);
or U1168 (N_1168,N_434,N_395);
nand U1169 (N_1169,N_421,N_758);
nand U1170 (N_1170,N_655,In_1012);
xor U1171 (N_1171,N_601,N_863);
xor U1172 (N_1172,N_433,N_586);
or U1173 (N_1173,N_829,N_870);
or U1174 (N_1174,N_844,N_603);
and U1175 (N_1175,N_843,N_493);
xnor U1176 (N_1176,In_1155,In_1376);
nor U1177 (N_1177,N_566,N_895);
nor U1178 (N_1178,In_353,In_807);
or U1179 (N_1179,N_615,N_722);
nor U1180 (N_1180,N_739,In_880);
nor U1181 (N_1181,In_1057,N_776);
nor U1182 (N_1182,N_819,N_736);
xnor U1183 (N_1183,N_410,In_697);
nor U1184 (N_1184,N_727,In_264);
xnor U1185 (N_1185,N_160,In_329);
or U1186 (N_1186,N_713,N_345);
or U1187 (N_1187,In_106,N_548);
xor U1188 (N_1188,N_509,N_613);
xnor U1189 (N_1189,N_620,N_468);
nand U1190 (N_1190,N_774,N_854);
nand U1191 (N_1191,N_285,N_647);
nor U1192 (N_1192,N_536,N_333);
and U1193 (N_1193,In_369,In_168);
and U1194 (N_1194,In_15,N_772);
xnor U1195 (N_1195,N_490,N_848);
and U1196 (N_1196,N_861,N_252);
nand U1197 (N_1197,N_640,In_1091);
xor U1198 (N_1198,N_853,N_830);
xor U1199 (N_1199,In_1217,In_1071);
xor U1200 (N_1200,N_998,N_1125);
nand U1201 (N_1201,N_914,N_1002);
or U1202 (N_1202,N_1179,N_935);
and U1203 (N_1203,N_931,N_1094);
xor U1204 (N_1204,N_1180,N_1060);
xnor U1205 (N_1205,N_933,N_909);
nor U1206 (N_1206,N_984,N_1088);
nor U1207 (N_1207,N_1131,N_1159);
nand U1208 (N_1208,N_1175,N_1185);
nand U1209 (N_1209,N_1102,N_1032);
nand U1210 (N_1210,N_1134,N_959);
xor U1211 (N_1211,N_1026,N_1091);
nor U1212 (N_1212,N_1015,N_1072);
xor U1213 (N_1213,N_1056,N_1005);
xnor U1214 (N_1214,N_1043,N_1055);
or U1215 (N_1215,N_1121,N_1151);
nor U1216 (N_1216,N_1053,N_1098);
xor U1217 (N_1217,N_925,N_1143);
xor U1218 (N_1218,N_1158,N_1068);
xor U1219 (N_1219,N_905,N_978);
or U1220 (N_1220,N_1148,N_1074);
nor U1221 (N_1221,N_1090,N_1167);
nor U1222 (N_1222,N_974,N_1122);
or U1223 (N_1223,N_1132,N_927);
nor U1224 (N_1224,N_1100,N_926);
nand U1225 (N_1225,N_901,N_981);
nand U1226 (N_1226,N_979,N_1199);
xor U1227 (N_1227,N_1051,N_1093);
nor U1228 (N_1228,N_928,N_1187);
or U1229 (N_1229,N_919,N_1017);
and U1230 (N_1230,N_1025,N_1110);
and U1231 (N_1231,N_1128,N_1118);
xnor U1232 (N_1232,N_1182,N_1003);
nand U1233 (N_1233,N_910,N_1112);
and U1234 (N_1234,N_1145,N_1194);
or U1235 (N_1235,N_936,N_1044);
and U1236 (N_1236,N_1142,N_1149);
and U1237 (N_1237,N_964,N_1061);
nand U1238 (N_1238,N_1156,N_916);
and U1239 (N_1239,N_947,N_1166);
nor U1240 (N_1240,N_1139,N_943);
and U1241 (N_1241,N_1083,N_983);
xnor U1242 (N_1242,N_1124,N_1073);
xnor U1243 (N_1243,N_1147,N_1186);
and U1244 (N_1244,N_1109,N_975);
and U1245 (N_1245,N_1157,N_1041);
nor U1246 (N_1246,N_1108,N_1107);
xor U1247 (N_1247,N_1009,N_1176);
or U1248 (N_1248,N_1081,N_902);
or U1249 (N_1249,N_1021,N_1066);
xor U1250 (N_1250,N_913,N_1054);
nand U1251 (N_1251,N_904,N_1011);
or U1252 (N_1252,N_934,N_1018);
xor U1253 (N_1253,N_980,N_1184);
or U1254 (N_1254,N_1138,N_973);
or U1255 (N_1255,N_966,N_1019);
nand U1256 (N_1256,N_1195,N_1065);
and U1257 (N_1257,N_1063,N_1155);
xnor U1258 (N_1258,N_906,N_985);
and U1259 (N_1259,N_1196,N_1096);
and U1260 (N_1260,N_956,N_1049);
nand U1261 (N_1261,N_986,N_1169);
nand U1262 (N_1262,N_1150,N_1008);
or U1263 (N_1263,N_1022,N_924);
nor U1264 (N_1264,N_1052,N_903);
xnor U1265 (N_1265,N_997,N_920);
and U1266 (N_1266,N_1127,N_1028);
nor U1267 (N_1267,N_921,N_1178);
or U1268 (N_1268,N_1016,N_1069);
xor U1269 (N_1269,N_1024,N_968);
nand U1270 (N_1270,N_1059,N_1075);
nand U1271 (N_1271,N_976,N_1086);
and U1272 (N_1272,N_945,N_908);
nand U1273 (N_1273,N_1153,N_932);
xor U1274 (N_1274,N_1040,N_922);
or U1275 (N_1275,N_1078,N_1058);
nor U1276 (N_1276,N_1077,N_1190);
and U1277 (N_1277,N_1144,N_1079);
nand U1278 (N_1278,N_1173,N_1038);
or U1279 (N_1279,N_1004,N_1103);
and U1280 (N_1280,N_970,N_1089);
and U1281 (N_1281,N_1029,N_950);
xor U1282 (N_1282,N_990,N_1023);
nor U1283 (N_1283,N_1126,N_941);
xnor U1284 (N_1284,N_1057,N_1120);
and U1285 (N_1285,N_957,N_1039);
xnor U1286 (N_1286,N_988,N_1113);
nand U1287 (N_1287,N_1010,N_1033);
or U1288 (N_1288,N_1042,N_1136);
nor U1289 (N_1289,N_989,N_948);
nor U1290 (N_1290,N_1162,N_1146);
xor U1291 (N_1291,N_949,N_1115);
nand U1292 (N_1292,N_1013,N_1076);
xnor U1293 (N_1293,N_1165,N_1101);
nor U1294 (N_1294,N_911,N_1097);
or U1295 (N_1295,N_1045,N_1172);
nor U1296 (N_1296,N_1007,N_1198);
xnor U1297 (N_1297,N_940,N_1141);
nor U1298 (N_1298,N_1197,N_923);
nand U1299 (N_1299,N_996,N_1030);
nand U1300 (N_1300,N_951,N_1189);
xnor U1301 (N_1301,N_1163,N_930);
xnor U1302 (N_1302,N_937,N_1114);
nand U1303 (N_1303,N_1160,N_939);
nor U1304 (N_1304,N_1048,N_1123);
and U1305 (N_1305,N_907,N_952);
nor U1306 (N_1306,N_992,N_1012);
or U1307 (N_1307,N_953,N_1064);
and U1308 (N_1308,N_1129,N_982);
and U1309 (N_1309,N_1027,N_1000);
nor U1310 (N_1310,N_1119,N_1036);
nand U1311 (N_1311,N_1014,N_1152);
nor U1312 (N_1312,N_1092,N_1117);
and U1313 (N_1313,N_944,N_929);
xor U1314 (N_1314,N_967,N_1104);
xnor U1315 (N_1315,N_938,N_1164);
and U1316 (N_1316,N_971,N_1161);
nor U1317 (N_1317,N_1037,N_999);
xnor U1318 (N_1318,N_1174,N_1192);
or U1319 (N_1319,N_955,N_918);
nor U1320 (N_1320,N_977,N_912);
nand U1321 (N_1321,N_958,N_1031);
nand U1322 (N_1322,N_1062,N_1035);
xor U1323 (N_1323,N_963,N_1168);
and U1324 (N_1324,N_954,N_1170);
xnor U1325 (N_1325,N_960,N_1135);
xnor U1326 (N_1326,N_917,N_1177);
and U1327 (N_1327,N_1034,N_962);
or U1328 (N_1328,N_1183,N_1116);
xnor U1329 (N_1329,N_1087,N_1191);
and U1330 (N_1330,N_915,N_1188);
and U1331 (N_1331,N_1133,N_1099);
or U1332 (N_1332,N_1050,N_961);
xnor U1333 (N_1333,N_987,N_1080);
or U1334 (N_1334,N_995,N_946);
nand U1335 (N_1335,N_991,N_1181);
or U1336 (N_1336,N_972,N_1106);
xnor U1337 (N_1337,N_1084,N_1111);
nand U1338 (N_1338,N_1006,N_993);
nand U1339 (N_1339,N_1137,N_994);
xor U1340 (N_1340,N_1082,N_965);
and U1341 (N_1341,N_969,N_1071);
or U1342 (N_1342,N_1067,N_1140);
xnor U1343 (N_1343,N_1095,N_1047);
nand U1344 (N_1344,N_942,N_1046);
or U1345 (N_1345,N_1105,N_1070);
and U1346 (N_1346,N_1020,N_1001);
nor U1347 (N_1347,N_900,N_1154);
or U1348 (N_1348,N_1085,N_1193);
and U1349 (N_1349,N_1171,N_1130);
nor U1350 (N_1350,N_1002,N_1119);
xnor U1351 (N_1351,N_1163,N_1012);
and U1352 (N_1352,N_973,N_1169);
and U1353 (N_1353,N_1114,N_1187);
or U1354 (N_1354,N_1031,N_1087);
nand U1355 (N_1355,N_1046,N_917);
and U1356 (N_1356,N_1039,N_991);
nor U1357 (N_1357,N_953,N_1160);
and U1358 (N_1358,N_978,N_1157);
xor U1359 (N_1359,N_1126,N_1058);
xor U1360 (N_1360,N_1112,N_1017);
xor U1361 (N_1361,N_1157,N_1026);
xnor U1362 (N_1362,N_1173,N_925);
nor U1363 (N_1363,N_972,N_948);
nor U1364 (N_1364,N_1145,N_919);
or U1365 (N_1365,N_1065,N_1056);
or U1366 (N_1366,N_1155,N_1191);
nor U1367 (N_1367,N_907,N_1049);
xnor U1368 (N_1368,N_1099,N_915);
or U1369 (N_1369,N_974,N_1153);
nor U1370 (N_1370,N_1171,N_1105);
or U1371 (N_1371,N_1038,N_1035);
and U1372 (N_1372,N_932,N_1094);
or U1373 (N_1373,N_912,N_1007);
or U1374 (N_1374,N_1052,N_947);
nor U1375 (N_1375,N_1077,N_924);
or U1376 (N_1376,N_1133,N_976);
nand U1377 (N_1377,N_1031,N_914);
nor U1378 (N_1378,N_957,N_1155);
and U1379 (N_1379,N_976,N_1014);
nand U1380 (N_1380,N_1177,N_1043);
nand U1381 (N_1381,N_945,N_921);
and U1382 (N_1382,N_959,N_1095);
xnor U1383 (N_1383,N_1091,N_958);
xnor U1384 (N_1384,N_1153,N_1120);
xor U1385 (N_1385,N_935,N_1090);
nand U1386 (N_1386,N_1053,N_908);
nor U1387 (N_1387,N_913,N_1110);
or U1388 (N_1388,N_1048,N_973);
xor U1389 (N_1389,N_925,N_976);
xor U1390 (N_1390,N_985,N_1075);
and U1391 (N_1391,N_1038,N_1115);
xnor U1392 (N_1392,N_940,N_1143);
nor U1393 (N_1393,N_1125,N_1193);
nor U1394 (N_1394,N_1196,N_1004);
or U1395 (N_1395,N_1068,N_994);
or U1396 (N_1396,N_1180,N_956);
and U1397 (N_1397,N_1180,N_905);
nand U1398 (N_1398,N_964,N_1162);
nand U1399 (N_1399,N_945,N_1109);
xor U1400 (N_1400,N_1088,N_1197);
xor U1401 (N_1401,N_1136,N_1077);
nor U1402 (N_1402,N_1114,N_953);
and U1403 (N_1403,N_1082,N_998);
or U1404 (N_1404,N_1048,N_1000);
nor U1405 (N_1405,N_1040,N_960);
or U1406 (N_1406,N_1103,N_1025);
xnor U1407 (N_1407,N_969,N_1151);
nand U1408 (N_1408,N_908,N_1125);
nor U1409 (N_1409,N_920,N_1129);
and U1410 (N_1410,N_1129,N_1168);
nand U1411 (N_1411,N_1033,N_938);
nor U1412 (N_1412,N_1183,N_1047);
and U1413 (N_1413,N_1035,N_932);
nor U1414 (N_1414,N_1130,N_1076);
and U1415 (N_1415,N_926,N_1185);
nor U1416 (N_1416,N_955,N_992);
or U1417 (N_1417,N_998,N_901);
or U1418 (N_1418,N_909,N_986);
xnor U1419 (N_1419,N_1038,N_938);
nor U1420 (N_1420,N_1100,N_1011);
xnor U1421 (N_1421,N_921,N_998);
and U1422 (N_1422,N_1084,N_1186);
nor U1423 (N_1423,N_1006,N_1188);
or U1424 (N_1424,N_1108,N_1004);
or U1425 (N_1425,N_976,N_950);
nand U1426 (N_1426,N_1075,N_991);
or U1427 (N_1427,N_1021,N_1128);
nor U1428 (N_1428,N_934,N_1170);
nand U1429 (N_1429,N_910,N_931);
or U1430 (N_1430,N_1047,N_1119);
and U1431 (N_1431,N_1082,N_964);
xnor U1432 (N_1432,N_1021,N_900);
nor U1433 (N_1433,N_1186,N_1145);
nor U1434 (N_1434,N_918,N_1050);
and U1435 (N_1435,N_1003,N_1027);
and U1436 (N_1436,N_1123,N_1176);
or U1437 (N_1437,N_1133,N_1129);
nor U1438 (N_1438,N_1066,N_1116);
nor U1439 (N_1439,N_1182,N_1103);
xnor U1440 (N_1440,N_992,N_1055);
or U1441 (N_1441,N_1053,N_1093);
or U1442 (N_1442,N_1193,N_1025);
nand U1443 (N_1443,N_1080,N_915);
nor U1444 (N_1444,N_1175,N_1160);
and U1445 (N_1445,N_1082,N_1089);
or U1446 (N_1446,N_915,N_992);
nand U1447 (N_1447,N_1034,N_1091);
nand U1448 (N_1448,N_1135,N_1130);
nand U1449 (N_1449,N_1005,N_1009);
xnor U1450 (N_1450,N_1187,N_1066);
nand U1451 (N_1451,N_963,N_1070);
and U1452 (N_1452,N_914,N_961);
and U1453 (N_1453,N_1161,N_902);
nand U1454 (N_1454,N_983,N_916);
or U1455 (N_1455,N_1010,N_1158);
and U1456 (N_1456,N_1086,N_1045);
and U1457 (N_1457,N_1038,N_958);
and U1458 (N_1458,N_903,N_1146);
nor U1459 (N_1459,N_1079,N_1070);
nor U1460 (N_1460,N_1062,N_970);
nor U1461 (N_1461,N_1105,N_1199);
and U1462 (N_1462,N_1034,N_1064);
xor U1463 (N_1463,N_1145,N_1050);
nand U1464 (N_1464,N_1004,N_1055);
nor U1465 (N_1465,N_1145,N_1110);
nand U1466 (N_1466,N_937,N_979);
or U1467 (N_1467,N_1112,N_944);
or U1468 (N_1468,N_934,N_1046);
or U1469 (N_1469,N_1055,N_965);
xnor U1470 (N_1470,N_1166,N_945);
and U1471 (N_1471,N_1031,N_1027);
and U1472 (N_1472,N_1155,N_974);
xor U1473 (N_1473,N_1179,N_1079);
xnor U1474 (N_1474,N_989,N_1040);
nor U1475 (N_1475,N_1173,N_934);
and U1476 (N_1476,N_1188,N_1093);
nor U1477 (N_1477,N_955,N_1115);
or U1478 (N_1478,N_989,N_1147);
xnor U1479 (N_1479,N_1157,N_1141);
nor U1480 (N_1480,N_925,N_1014);
or U1481 (N_1481,N_1016,N_919);
nand U1482 (N_1482,N_1066,N_1047);
nand U1483 (N_1483,N_1034,N_1040);
xor U1484 (N_1484,N_943,N_1106);
xnor U1485 (N_1485,N_1049,N_1124);
nor U1486 (N_1486,N_1056,N_1046);
nand U1487 (N_1487,N_1021,N_972);
nand U1488 (N_1488,N_1145,N_921);
nor U1489 (N_1489,N_986,N_905);
or U1490 (N_1490,N_1173,N_1065);
nor U1491 (N_1491,N_1133,N_1101);
or U1492 (N_1492,N_1156,N_933);
nand U1493 (N_1493,N_1190,N_1003);
xnor U1494 (N_1494,N_941,N_1196);
or U1495 (N_1495,N_965,N_1198);
nor U1496 (N_1496,N_984,N_1186);
xnor U1497 (N_1497,N_1164,N_905);
or U1498 (N_1498,N_987,N_1133);
and U1499 (N_1499,N_1080,N_1024);
and U1500 (N_1500,N_1413,N_1329);
nand U1501 (N_1501,N_1373,N_1448);
xor U1502 (N_1502,N_1435,N_1345);
nand U1503 (N_1503,N_1230,N_1442);
and U1504 (N_1504,N_1419,N_1256);
and U1505 (N_1505,N_1396,N_1222);
and U1506 (N_1506,N_1370,N_1382);
nor U1507 (N_1507,N_1245,N_1441);
xnor U1508 (N_1508,N_1335,N_1307);
nor U1509 (N_1509,N_1494,N_1460);
nand U1510 (N_1510,N_1499,N_1491);
xor U1511 (N_1511,N_1418,N_1263);
or U1512 (N_1512,N_1232,N_1341);
nand U1513 (N_1513,N_1318,N_1259);
nor U1514 (N_1514,N_1313,N_1324);
nor U1515 (N_1515,N_1411,N_1476);
xor U1516 (N_1516,N_1384,N_1445);
and U1517 (N_1517,N_1352,N_1430);
nand U1518 (N_1518,N_1402,N_1268);
or U1519 (N_1519,N_1303,N_1393);
or U1520 (N_1520,N_1200,N_1409);
nor U1521 (N_1521,N_1250,N_1489);
nand U1522 (N_1522,N_1467,N_1277);
nand U1523 (N_1523,N_1255,N_1378);
nor U1524 (N_1524,N_1388,N_1415);
or U1525 (N_1525,N_1210,N_1495);
nor U1526 (N_1526,N_1360,N_1302);
xnor U1527 (N_1527,N_1377,N_1278);
xnor U1528 (N_1528,N_1457,N_1426);
or U1529 (N_1529,N_1219,N_1465);
or U1530 (N_1530,N_1266,N_1216);
and U1531 (N_1531,N_1251,N_1434);
nand U1532 (N_1532,N_1447,N_1408);
or U1533 (N_1533,N_1497,N_1471);
nor U1534 (N_1534,N_1387,N_1272);
nor U1535 (N_1535,N_1308,N_1211);
or U1536 (N_1536,N_1295,N_1486);
nand U1537 (N_1537,N_1473,N_1480);
nor U1538 (N_1538,N_1223,N_1493);
xnor U1539 (N_1539,N_1299,N_1429);
and U1540 (N_1540,N_1414,N_1215);
nand U1541 (N_1541,N_1237,N_1201);
nand U1542 (N_1542,N_1479,N_1338);
and U1543 (N_1543,N_1422,N_1317);
xnor U1544 (N_1544,N_1294,N_1403);
nand U1545 (N_1545,N_1398,N_1264);
xnor U1546 (N_1546,N_1300,N_1433);
nor U1547 (N_1547,N_1217,N_1375);
or U1548 (N_1548,N_1290,N_1391);
nor U1549 (N_1549,N_1466,N_1236);
nand U1550 (N_1550,N_1383,N_1292);
and U1551 (N_1551,N_1253,N_1273);
nor U1552 (N_1552,N_1337,N_1298);
xor U1553 (N_1553,N_1260,N_1349);
and U1554 (N_1554,N_1346,N_1395);
nor U1555 (N_1555,N_1348,N_1356);
nand U1556 (N_1556,N_1463,N_1340);
xnor U1557 (N_1557,N_1364,N_1355);
or U1558 (N_1558,N_1354,N_1453);
and U1559 (N_1559,N_1417,N_1488);
or U1560 (N_1560,N_1496,N_1212);
or U1561 (N_1561,N_1220,N_1311);
xor U1562 (N_1562,N_1362,N_1490);
nand U1563 (N_1563,N_1379,N_1305);
xor U1564 (N_1564,N_1443,N_1416);
nor U1565 (N_1565,N_1241,N_1455);
nor U1566 (N_1566,N_1328,N_1452);
nand U1567 (N_1567,N_1314,N_1454);
xnor U1568 (N_1568,N_1286,N_1380);
or U1569 (N_1569,N_1226,N_1470);
and U1570 (N_1570,N_1254,N_1406);
or U1571 (N_1571,N_1483,N_1249);
xnor U1572 (N_1572,N_1297,N_1291);
nor U1573 (N_1573,N_1482,N_1449);
xnor U1574 (N_1574,N_1353,N_1397);
and U1575 (N_1575,N_1209,N_1390);
nand U1576 (N_1576,N_1410,N_1248);
nand U1577 (N_1577,N_1213,N_1350);
or U1578 (N_1578,N_1316,N_1359);
xor U1579 (N_1579,N_1456,N_1468);
or U1580 (N_1580,N_1431,N_1240);
xnor U1581 (N_1581,N_1386,N_1405);
or U1582 (N_1582,N_1310,N_1458);
nor U1583 (N_1583,N_1381,N_1421);
nor U1584 (N_1584,N_1203,N_1374);
nor U1585 (N_1585,N_1366,N_1440);
and U1586 (N_1586,N_1427,N_1437);
nand U1587 (N_1587,N_1274,N_1235);
nand U1588 (N_1588,N_1309,N_1239);
and U1589 (N_1589,N_1287,N_1214);
nor U1590 (N_1590,N_1306,N_1492);
or U1591 (N_1591,N_1246,N_1400);
or U1592 (N_1592,N_1267,N_1339);
or U1593 (N_1593,N_1234,N_1281);
nor U1594 (N_1594,N_1261,N_1227);
or U1595 (N_1595,N_1385,N_1205);
nand U1596 (N_1596,N_1423,N_1289);
or U1597 (N_1597,N_1464,N_1399);
nor U1598 (N_1598,N_1224,N_1365);
and U1599 (N_1599,N_1438,N_1279);
and U1600 (N_1600,N_1207,N_1444);
nor U1601 (N_1601,N_1342,N_1233);
or U1602 (N_1602,N_1344,N_1367);
nand U1603 (N_1603,N_1280,N_1481);
xor U1604 (N_1604,N_1478,N_1477);
or U1605 (N_1605,N_1484,N_1363);
or U1606 (N_1606,N_1218,N_1229);
nor U1607 (N_1607,N_1371,N_1432);
or U1608 (N_1608,N_1247,N_1336);
xor U1609 (N_1609,N_1242,N_1271);
nand U1610 (N_1610,N_1231,N_1469);
and U1611 (N_1611,N_1320,N_1225);
xnor U1612 (N_1612,N_1228,N_1252);
nand U1613 (N_1613,N_1368,N_1401);
and U1614 (N_1614,N_1351,N_1372);
or U1615 (N_1615,N_1204,N_1420);
xor U1616 (N_1616,N_1221,N_1330);
or U1617 (N_1617,N_1319,N_1282);
or U1618 (N_1618,N_1244,N_1208);
or U1619 (N_1619,N_1276,N_1258);
or U1620 (N_1620,N_1288,N_1474);
nor U1621 (N_1621,N_1322,N_1394);
and U1622 (N_1622,N_1243,N_1475);
and U1623 (N_1623,N_1459,N_1361);
xor U1624 (N_1624,N_1275,N_1301);
nor U1625 (N_1625,N_1315,N_1321);
nor U1626 (N_1626,N_1269,N_1392);
and U1627 (N_1627,N_1334,N_1293);
or U1628 (N_1628,N_1498,N_1326);
or U1629 (N_1629,N_1357,N_1358);
nand U1630 (N_1630,N_1424,N_1327);
xor U1631 (N_1631,N_1404,N_1285);
and U1632 (N_1632,N_1332,N_1257);
or U1633 (N_1633,N_1283,N_1343);
nand U1634 (N_1634,N_1270,N_1284);
nor U1635 (N_1635,N_1376,N_1265);
and U1636 (N_1636,N_1333,N_1262);
or U1637 (N_1637,N_1451,N_1304);
or U1638 (N_1638,N_1436,N_1407);
xnor U1639 (N_1639,N_1461,N_1412);
xnor U1640 (N_1640,N_1331,N_1450);
nand U1641 (N_1641,N_1439,N_1428);
xnor U1642 (N_1642,N_1472,N_1238);
and U1643 (N_1643,N_1446,N_1312);
and U1644 (N_1644,N_1202,N_1296);
or U1645 (N_1645,N_1487,N_1347);
and U1646 (N_1646,N_1325,N_1206);
or U1647 (N_1647,N_1462,N_1389);
nand U1648 (N_1648,N_1485,N_1369);
xor U1649 (N_1649,N_1323,N_1425);
nand U1650 (N_1650,N_1408,N_1349);
or U1651 (N_1651,N_1247,N_1257);
nand U1652 (N_1652,N_1392,N_1256);
xor U1653 (N_1653,N_1403,N_1454);
nand U1654 (N_1654,N_1231,N_1252);
xnor U1655 (N_1655,N_1271,N_1493);
nor U1656 (N_1656,N_1306,N_1431);
or U1657 (N_1657,N_1209,N_1346);
nand U1658 (N_1658,N_1277,N_1229);
nor U1659 (N_1659,N_1304,N_1353);
nand U1660 (N_1660,N_1408,N_1375);
nor U1661 (N_1661,N_1333,N_1470);
and U1662 (N_1662,N_1370,N_1428);
nor U1663 (N_1663,N_1398,N_1351);
nand U1664 (N_1664,N_1471,N_1311);
and U1665 (N_1665,N_1350,N_1435);
nor U1666 (N_1666,N_1268,N_1380);
nand U1667 (N_1667,N_1317,N_1433);
nand U1668 (N_1668,N_1262,N_1404);
or U1669 (N_1669,N_1343,N_1318);
nor U1670 (N_1670,N_1334,N_1217);
nand U1671 (N_1671,N_1216,N_1435);
nor U1672 (N_1672,N_1465,N_1349);
nand U1673 (N_1673,N_1269,N_1384);
nor U1674 (N_1674,N_1371,N_1297);
or U1675 (N_1675,N_1494,N_1451);
xor U1676 (N_1676,N_1375,N_1457);
nand U1677 (N_1677,N_1382,N_1304);
nand U1678 (N_1678,N_1433,N_1272);
and U1679 (N_1679,N_1307,N_1238);
nor U1680 (N_1680,N_1272,N_1206);
nand U1681 (N_1681,N_1316,N_1279);
and U1682 (N_1682,N_1449,N_1461);
nand U1683 (N_1683,N_1360,N_1423);
nor U1684 (N_1684,N_1311,N_1269);
xnor U1685 (N_1685,N_1369,N_1498);
xnor U1686 (N_1686,N_1393,N_1378);
xor U1687 (N_1687,N_1352,N_1438);
xnor U1688 (N_1688,N_1443,N_1357);
xnor U1689 (N_1689,N_1228,N_1476);
nand U1690 (N_1690,N_1330,N_1429);
nand U1691 (N_1691,N_1385,N_1255);
and U1692 (N_1692,N_1465,N_1379);
nand U1693 (N_1693,N_1259,N_1226);
or U1694 (N_1694,N_1302,N_1430);
xnor U1695 (N_1695,N_1355,N_1454);
xnor U1696 (N_1696,N_1429,N_1357);
nand U1697 (N_1697,N_1293,N_1296);
nand U1698 (N_1698,N_1351,N_1488);
nand U1699 (N_1699,N_1216,N_1237);
nor U1700 (N_1700,N_1219,N_1337);
and U1701 (N_1701,N_1383,N_1340);
or U1702 (N_1702,N_1203,N_1484);
nor U1703 (N_1703,N_1304,N_1410);
nor U1704 (N_1704,N_1237,N_1294);
or U1705 (N_1705,N_1462,N_1393);
xor U1706 (N_1706,N_1294,N_1321);
nand U1707 (N_1707,N_1312,N_1481);
nor U1708 (N_1708,N_1346,N_1498);
and U1709 (N_1709,N_1333,N_1396);
nand U1710 (N_1710,N_1311,N_1417);
nor U1711 (N_1711,N_1292,N_1497);
nand U1712 (N_1712,N_1387,N_1429);
nor U1713 (N_1713,N_1430,N_1226);
xor U1714 (N_1714,N_1436,N_1308);
or U1715 (N_1715,N_1269,N_1209);
or U1716 (N_1716,N_1239,N_1401);
or U1717 (N_1717,N_1312,N_1488);
nand U1718 (N_1718,N_1398,N_1299);
and U1719 (N_1719,N_1442,N_1387);
and U1720 (N_1720,N_1440,N_1473);
or U1721 (N_1721,N_1410,N_1380);
and U1722 (N_1722,N_1392,N_1253);
nor U1723 (N_1723,N_1473,N_1224);
xnor U1724 (N_1724,N_1267,N_1381);
or U1725 (N_1725,N_1445,N_1354);
or U1726 (N_1726,N_1210,N_1261);
nor U1727 (N_1727,N_1410,N_1411);
xnor U1728 (N_1728,N_1441,N_1271);
and U1729 (N_1729,N_1481,N_1391);
nor U1730 (N_1730,N_1272,N_1379);
xnor U1731 (N_1731,N_1295,N_1230);
and U1732 (N_1732,N_1241,N_1255);
or U1733 (N_1733,N_1443,N_1303);
or U1734 (N_1734,N_1376,N_1448);
nor U1735 (N_1735,N_1263,N_1211);
nor U1736 (N_1736,N_1334,N_1415);
or U1737 (N_1737,N_1473,N_1246);
nand U1738 (N_1738,N_1356,N_1486);
or U1739 (N_1739,N_1284,N_1362);
nor U1740 (N_1740,N_1475,N_1301);
xor U1741 (N_1741,N_1202,N_1334);
or U1742 (N_1742,N_1367,N_1488);
or U1743 (N_1743,N_1255,N_1459);
nor U1744 (N_1744,N_1422,N_1386);
nand U1745 (N_1745,N_1224,N_1316);
xnor U1746 (N_1746,N_1462,N_1461);
nand U1747 (N_1747,N_1422,N_1497);
and U1748 (N_1748,N_1455,N_1487);
nor U1749 (N_1749,N_1317,N_1432);
xor U1750 (N_1750,N_1396,N_1297);
xnor U1751 (N_1751,N_1236,N_1465);
nor U1752 (N_1752,N_1439,N_1359);
or U1753 (N_1753,N_1452,N_1273);
and U1754 (N_1754,N_1445,N_1250);
xnor U1755 (N_1755,N_1430,N_1497);
nor U1756 (N_1756,N_1270,N_1341);
or U1757 (N_1757,N_1264,N_1493);
or U1758 (N_1758,N_1230,N_1264);
nand U1759 (N_1759,N_1421,N_1454);
xor U1760 (N_1760,N_1384,N_1303);
nand U1761 (N_1761,N_1217,N_1361);
or U1762 (N_1762,N_1306,N_1227);
nor U1763 (N_1763,N_1370,N_1273);
nand U1764 (N_1764,N_1382,N_1492);
xor U1765 (N_1765,N_1466,N_1407);
xor U1766 (N_1766,N_1459,N_1290);
and U1767 (N_1767,N_1449,N_1422);
and U1768 (N_1768,N_1233,N_1293);
or U1769 (N_1769,N_1368,N_1359);
or U1770 (N_1770,N_1237,N_1281);
or U1771 (N_1771,N_1280,N_1409);
and U1772 (N_1772,N_1346,N_1445);
xnor U1773 (N_1773,N_1402,N_1477);
xnor U1774 (N_1774,N_1426,N_1243);
nor U1775 (N_1775,N_1424,N_1208);
and U1776 (N_1776,N_1339,N_1369);
nand U1777 (N_1777,N_1430,N_1291);
nor U1778 (N_1778,N_1465,N_1257);
nor U1779 (N_1779,N_1394,N_1366);
xnor U1780 (N_1780,N_1459,N_1376);
xor U1781 (N_1781,N_1263,N_1430);
and U1782 (N_1782,N_1277,N_1212);
nor U1783 (N_1783,N_1388,N_1463);
and U1784 (N_1784,N_1489,N_1312);
and U1785 (N_1785,N_1496,N_1455);
nand U1786 (N_1786,N_1478,N_1441);
xor U1787 (N_1787,N_1241,N_1274);
nor U1788 (N_1788,N_1480,N_1423);
or U1789 (N_1789,N_1436,N_1332);
and U1790 (N_1790,N_1233,N_1317);
or U1791 (N_1791,N_1386,N_1399);
xor U1792 (N_1792,N_1433,N_1350);
or U1793 (N_1793,N_1319,N_1415);
nand U1794 (N_1794,N_1454,N_1336);
and U1795 (N_1795,N_1468,N_1228);
and U1796 (N_1796,N_1411,N_1345);
xnor U1797 (N_1797,N_1384,N_1485);
and U1798 (N_1798,N_1283,N_1249);
nor U1799 (N_1799,N_1402,N_1396);
or U1800 (N_1800,N_1669,N_1576);
or U1801 (N_1801,N_1717,N_1549);
xor U1802 (N_1802,N_1755,N_1526);
nand U1803 (N_1803,N_1770,N_1541);
or U1804 (N_1804,N_1668,N_1615);
or U1805 (N_1805,N_1546,N_1720);
nand U1806 (N_1806,N_1693,N_1640);
nand U1807 (N_1807,N_1653,N_1609);
and U1808 (N_1808,N_1713,N_1771);
xnor U1809 (N_1809,N_1548,N_1568);
xnor U1810 (N_1810,N_1772,N_1676);
and U1811 (N_1811,N_1697,N_1746);
nor U1812 (N_1812,N_1701,N_1736);
xnor U1813 (N_1813,N_1727,N_1602);
or U1814 (N_1814,N_1675,N_1794);
or U1815 (N_1815,N_1776,N_1501);
and U1816 (N_1816,N_1798,N_1762);
or U1817 (N_1817,N_1633,N_1751);
nand U1818 (N_1818,N_1796,N_1723);
xor U1819 (N_1819,N_1612,N_1559);
nand U1820 (N_1820,N_1705,N_1672);
nor U1821 (N_1821,N_1689,N_1539);
nor U1822 (N_1822,N_1745,N_1550);
nand U1823 (N_1823,N_1587,N_1756);
xor U1824 (N_1824,N_1714,N_1650);
xnor U1825 (N_1825,N_1505,N_1696);
xnor U1826 (N_1826,N_1670,N_1513);
and U1827 (N_1827,N_1608,N_1597);
and U1828 (N_1828,N_1520,N_1622);
nand U1829 (N_1829,N_1715,N_1545);
nand U1830 (N_1830,N_1719,N_1799);
and U1831 (N_1831,N_1542,N_1777);
nand U1832 (N_1832,N_1692,N_1793);
nor U1833 (N_1833,N_1752,N_1765);
nor U1834 (N_1834,N_1632,N_1671);
xnor U1835 (N_1835,N_1710,N_1707);
or U1836 (N_1836,N_1634,N_1786);
nand U1837 (N_1837,N_1682,N_1596);
and U1838 (N_1838,N_1761,N_1709);
and U1839 (N_1839,N_1721,N_1780);
or U1840 (N_1840,N_1698,N_1657);
nand U1841 (N_1841,N_1730,N_1544);
xor U1842 (N_1842,N_1591,N_1665);
xor U1843 (N_1843,N_1699,N_1624);
and U1844 (N_1844,N_1645,N_1528);
nor U1845 (N_1845,N_1789,N_1572);
or U1846 (N_1846,N_1636,N_1625);
nor U1847 (N_1847,N_1790,N_1662);
nor U1848 (N_1848,N_1503,N_1654);
nand U1849 (N_1849,N_1579,N_1763);
or U1850 (N_1850,N_1718,N_1535);
nand U1851 (N_1851,N_1733,N_1614);
nand U1852 (N_1852,N_1511,N_1700);
or U1853 (N_1853,N_1722,N_1651);
and U1854 (N_1854,N_1729,N_1639);
xor U1855 (N_1855,N_1741,N_1647);
nor U1856 (N_1856,N_1641,N_1767);
and U1857 (N_1857,N_1575,N_1571);
xor U1858 (N_1858,N_1522,N_1747);
or U1859 (N_1859,N_1703,N_1795);
nor U1860 (N_1860,N_1552,N_1768);
nor U1861 (N_1861,N_1581,N_1791);
nor U1862 (N_1862,N_1758,N_1578);
or U1863 (N_1863,N_1691,N_1536);
or U1864 (N_1864,N_1557,N_1530);
and U1865 (N_1865,N_1684,N_1616);
or U1866 (N_1866,N_1788,N_1540);
xor U1867 (N_1867,N_1748,N_1617);
or U1868 (N_1868,N_1563,N_1686);
xor U1869 (N_1869,N_1712,N_1588);
xor U1870 (N_1870,N_1594,N_1677);
and U1871 (N_1871,N_1764,N_1562);
and U1872 (N_1872,N_1627,N_1613);
or U1873 (N_1873,N_1585,N_1551);
xnor U1874 (N_1874,N_1678,N_1644);
xor U1875 (N_1875,N_1601,N_1648);
xor U1876 (N_1876,N_1569,N_1655);
nor U1877 (N_1877,N_1754,N_1620);
and U1878 (N_1878,N_1660,N_1740);
nor U1879 (N_1879,N_1659,N_1652);
and U1880 (N_1880,N_1716,N_1739);
nor U1881 (N_1881,N_1529,N_1726);
nand U1882 (N_1882,N_1749,N_1523);
nand U1883 (N_1883,N_1728,N_1792);
nand U1884 (N_1884,N_1553,N_1512);
nand U1885 (N_1885,N_1574,N_1642);
nor U1886 (N_1886,N_1577,N_1628);
nand U1887 (N_1887,N_1610,N_1606);
nand U1888 (N_1888,N_1742,N_1760);
xnor U1889 (N_1889,N_1711,N_1781);
and U1890 (N_1890,N_1573,N_1773);
xor U1891 (N_1891,N_1704,N_1674);
nand U1892 (N_1892,N_1702,N_1527);
xnor U1893 (N_1893,N_1538,N_1524);
or U1894 (N_1894,N_1688,N_1626);
nor U1895 (N_1895,N_1743,N_1533);
nand U1896 (N_1896,N_1566,N_1782);
nor U1897 (N_1897,N_1619,N_1661);
or U1898 (N_1898,N_1507,N_1779);
nand U1899 (N_1899,N_1774,N_1508);
or U1900 (N_1900,N_1695,N_1685);
nor U1901 (N_1901,N_1637,N_1631);
nand U1902 (N_1902,N_1502,N_1738);
xnor U1903 (N_1903,N_1666,N_1744);
nand U1904 (N_1904,N_1680,N_1517);
or U1905 (N_1905,N_1667,N_1778);
nor U1906 (N_1906,N_1732,N_1784);
nor U1907 (N_1907,N_1595,N_1555);
xor U1908 (N_1908,N_1509,N_1621);
xnor U1909 (N_1909,N_1673,N_1554);
nand U1910 (N_1910,N_1506,N_1605);
nand U1911 (N_1911,N_1750,N_1561);
nand U1912 (N_1912,N_1757,N_1769);
xor U1913 (N_1913,N_1504,N_1759);
or U1914 (N_1914,N_1560,N_1656);
and U1915 (N_1915,N_1635,N_1629);
and U1916 (N_1916,N_1516,N_1567);
nand U1917 (N_1917,N_1694,N_1708);
xnor U1918 (N_1918,N_1525,N_1531);
nor U1919 (N_1919,N_1521,N_1681);
xor U1920 (N_1920,N_1593,N_1515);
or U1921 (N_1921,N_1623,N_1664);
nand U1922 (N_1922,N_1663,N_1519);
nand U1923 (N_1923,N_1565,N_1783);
xnor U1924 (N_1924,N_1725,N_1590);
nand U1925 (N_1925,N_1618,N_1510);
nor U1926 (N_1926,N_1586,N_1584);
nand U1927 (N_1927,N_1638,N_1607);
or U1928 (N_1928,N_1731,N_1658);
and U1929 (N_1929,N_1687,N_1690);
and U1930 (N_1930,N_1611,N_1583);
xnor U1931 (N_1931,N_1630,N_1797);
or U1932 (N_1932,N_1604,N_1582);
nor U1933 (N_1933,N_1649,N_1570);
or U1934 (N_1934,N_1558,N_1603);
nor U1935 (N_1935,N_1775,N_1534);
nor U1936 (N_1936,N_1600,N_1766);
nor U1937 (N_1937,N_1500,N_1787);
nand U1938 (N_1938,N_1643,N_1679);
nand U1939 (N_1939,N_1592,N_1532);
and U1940 (N_1940,N_1598,N_1724);
nand U1941 (N_1941,N_1737,N_1564);
and U1942 (N_1942,N_1537,N_1547);
xnor U1943 (N_1943,N_1589,N_1518);
or U1944 (N_1944,N_1753,N_1514);
xor U1945 (N_1945,N_1706,N_1785);
nor U1946 (N_1946,N_1580,N_1735);
xor U1947 (N_1947,N_1599,N_1683);
or U1948 (N_1948,N_1543,N_1734);
and U1949 (N_1949,N_1646,N_1556);
and U1950 (N_1950,N_1539,N_1615);
nand U1951 (N_1951,N_1520,N_1525);
nand U1952 (N_1952,N_1751,N_1779);
and U1953 (N_1953,N_1604,N_1693);
xnor U1954 (N_1954,N_1684,N_1789);
or U1955 (N_1955,N_1711,N_1734);
or U1956 (N_1956,N_1572,N_1606);
and U1957 (N_1957,N_1555,N_1679);
and U1958 (N_1958,N_1555,N_1552);
and U1959 (N_1959,N_1700,N_1764);
and U1960 (N_1960,N_1707,N_1540);
nand U1961 (N_1961,N_1700,N_1556);
and U1962 (N_1962,N_1543,N_1654);
xor U1963 (N_1963,N_1729,N_1517);
and U1964 (N_1964,N_1753,N_1722);
or U1965 (N_1965,N_1528,N_1532);
nor U1966 (N_1966,N_1661,N_1652);
and U1967 (N_1967,N_1640,N_1591);
nand U1968 (N_1968,N_1613,N_1675);
and U1969 (N_1969,N_1780,N_1799);
nor U1970 (N_1970,N_1657,N_1634);
nand U1971 (N_1971,N_1716,N_1766);
or U1972 (N_1972,N_1691,N_1539);
or U1973 (N_1973,N_1748,N_1799);
and U1974 (N_1974,N_1762,N_1550);
nand U1975 (N_1975,N_1582,N_1578);
xor U1976 (N_1976,N_1751,N_1613);
xor U1977 (N_1977,N_1772,N_1571);
or U1978 (N_1978,N_1511,N_1570);
and U1979 (N_1979,N_1581,N_1701);
and U1980 (N_1980,N_1585,N_1776);
nor U1981 (N_1981,N_1755,N_1737);
xor U1982 (N_1982,N_1686,N_1617);
nand U1983 (N_1983,N_1630,N_1525);
nor U1984 (N_1984,N_1582,N_1721);
nand U1985 (N_1985,N_1666,N_1519);
and U1986 (N_1986,N_1579,N_1715);
or U1987 (N_1987,N_1585,N_1661);
nor U1988 (N_1988,N_1517,N_1545);
nor U1989 (N_1989,N_1708,N_1614);
nand U1990 (N_1990,N_1501,N_1724);
nand U1991 (N_1991,N_1704,N_1761);
or U1992 (N_1992,N_1601,N_1552);
or U1993 (N_1993,N_1651,N_1517);
xnor U1994 (N_1994,N_1769,N_1664);
and U1995 (N_1995,N_1728,N_1595);
or U1996 (N_1996,N_1647,N_1603);
xor U1997 (N_1997,N_1628,N_1572);
or U1998 (N_1998,N_1670,N_1514);
and U1999 (N_1999,N_1561,N_1656);
and U2000 (N_2000,N_1691,N_1540);
and U2001 (N_2001,N_1583,N_1738);
nand U2002 (N_2002,N_1670,N_1700);
nor U2003 (N_2003,N_1538,N_1580);
nor U2004 (N_2004,N_1713,N_1760);
xor U2005 (N_2005,N_1755,N_1556);
or U2006 (N_2006,N_1734,N_1692);
nor U2007 (N_2007,N_1714,N_1764);
nor U2008 (N_2008,N_1759,N_1772);
and U2009 (N_2009,N_1631,N_1648);
nand U2010 (N_2010,N_1737,N_1540);
nor U2011 (N_2011,N_1753,N_1660);
nand U2012 (N_2012,N_1652,N_1714);
or U2013 (N_2013,N_1587,N_1744);
nor U2014 (N_2014,N_1766,N_1749);
or U2015 (N_2015,N_1799,N_1674);
and U2016 (N_2016,N_1759,N_1724);
xor U2017 (N_2017,N_1688,N_1527);
and U2018 (N_2018,N_1521,N_1594);
and U2019 (N_2019,N_1764,N_1528);
or U2020 (N_2020,N_1747,N_1599);
or U2021 (N_2021,N_1667,N_1634);
xor U2022 (N_2022,N_1690,N_1635);
nor U2023 (N_2023,N_1662,N_1678);
and U2024 (N_2024,N_1547,N_1795);
xnor U2025 (N_2025,N_1694,N_1703);
nand U2026 (N_2026,N_1546,N_1626);
and U2027 (N_2027,N_1789,N_1587);
xor U2028 (N_2028,N_1796,N_1618);
nor U2029 (N_2029,N_1659,N_1613);
xnor U2030 (N_2030,N_1784,N_1648);
nor U2031 (N_2031,N_1529,N_1599);
or U2032 (N_2032,N_1687,N_1594);
xor U2033 (N_2033,N_1798,N_1608);
nor U2034 (N_2034,N_1694,N_1559);
nand U2035 (N_2035,N_1788,N_1647);
and U2036 (N_2036,N_1611,N_1722);
and U2037 (N_2037,N_1523,N_1789);
or U2038 (N_2038,N_1637,N_1730);
nor U2039 (N_2039,N_1630,N_1756);
nor U2040 (N_2040,N_1563,N_1657);
or U2041 (N_2041,N_1554,N_1732);
or U2042 (N_2042,N_1765,N_1618);
or U2043 (N_2043,N_1556,N_1581);
nor U2044 (N_2044,N_1519,N_1656);
or U2045 (N_2045,N_1508,N_1687);
and U2046 (N_2046,N_1720,N_1616);
nor U2047 (N_2047,N_1719,N_1740);
xnor U2048 (N_2048,N_1645,N_1784);
nand U2049 (N_2049,N_1579,N_1511);
nor U2050 (N_2050,N_1730,N_1584);
or U2051 (N_2051,N_1706,N_1663);
nand U2052 (N_2052,N_1638,N_1636);
nand U2053 (N_2053,N_1623,N_1737);
nand U2054 (N_2054,N_1520,N_1759);
or U2055 (N_2055,N_1591,N_1610);
nand U2056 (N_2056,N_1514,N_1700);
xnor U2057 (N_2057,N_1610,N_1545);
xor U2058 (N_2058,N_1726,N_1700);
or U2059 (N_2059,N_1763,N_1573);
and U2060 (N_2060,N_1675,N_1610);
nor U2061 (N_2061,N_1537,N_1691);
nand U2062 (N_2062,N_1527,N_1551);
nand U2063 (N_2063,N_1541,N_1769);
or U2064 (N_2064,N_1734,N_1544);
xor U2065 (N_2065,N_1721,N_1761);
xnor U2066 (N_2066,N_1506,N_1630);
nor U2067 (N_2067,N_1655,N_1636);
nand U2068 (N_2068,N_1622,N_1721);
or U2069 (N_2069,N_1561,N_1635);
and U2070 (N_2070,N_1657,N_1740);
nand U2071 (N_2071,N_1539,N_1677);
nor U2072 (N_2072,N_1669,N_1746);
nand U2073 (N_2073,N_1719,N_1587);
xnor U2074 (N_2074,N_1623,N_1591);
nor U2075 (N_2075,N_1793,N_1611);
nand U2076 (N_2076,N_1637,N_1787);
nand U2077 (N_2077,N_1557,N_1647);
nor U2078 (N_2078,N_1696,N_1793);
nand U2079 (N_2079,N_1598,N_1571);
and U2080 (N_2080,N_1548,N_1710);
nor U2081 (N_2081,N_1648,N_1567);
nor U2082 (N_2082,N_1621,N_1627);
nand U2083 (N_2083,N_1530,N_1569);
and U2084 (N_2084,N_1793,N_1711);
xnor U2085 (N_2085,N_1754,N_1670);
nand U2086 (N_2086,N_1539,N_1512);
xor U2087 (N_2087,N_1723,N_1642);
and U2088 (N_2088,N_1583,N_1675);
nor U2089 (N_2089,N_1676,N_1782);
or U2090 (N_2090,N_1675,N_1528);
nand U2091 (N_2091,N_1770,N_1542);
and U2092 (N_2092,N_1505,N_1798);
and U2093 (N_2093,N_1569,N_1643);
nor U2094 (N_2094,N_1524,N_1560);
and U2095 (N_2095,N_1590,N_1719);
and U2096 (N_2096,N_1686,N_1656);
or U2097 (N_2097,N_1533,N_1657);
and U2098 (N_2098,N_1527,N_1560);
or U2099 (N_2099,N_1562,N_1785);
nor U2100 (N_2100,N_2008,N_1904);
and U2101 (N_2101,N_1809,N_1872);
xnor U2102 (N_2102,N_1948,N_2017);
nand U2103 (N_2103,N_2065,N_1922);
and U2104 (N_2104,N_2026,N_2032);
or U2105 (N_2105,N_1895,N_2078);
xor U2106 (N_2106,N_2098,N_2072);
xnor U2107 (N_2107,N_2034,N_1881);
nand U2108 (N_2108,N_1868,N_1934);
and U2109 (N_2109,N_2091,N_1827);
and U2110 (N_2110,N_1834,N_2070);
nor U2111 (N_2111,N_2074,N_2093);
xnor U2112 (N_2112,N_2045,N_1919);
xor U2113 (N_2113,N_1929,N_2069);
nand U2114 (N_2114,N_1982,N_1820);
nand U2115 (N_2115,N_2005,N_2052);
or U2116 (N_2116,N_2048,N_1987);
or U2117 (N_2117,N_1915,N_2022);
or U2118 (N_2118,N_1962,N_1873);
and U2119 (N_2119,N_2007,N_1952);
or U2120 (N_2120,N_1983,N_1814);
nand U2121 (N_2121,N_1837,N_1882);
nand U2122 (N_2122,N_1801,N_1829);
and U2123 (N_2123,N_1965,N_2023);
and U2124 (N_2124,N_2024,N_2056);
and U2125 (N_2125,N_1985,N_1889);
nand U2126 (N_2126,N_1943,N_2071);
nor U2127 (N_2127,N_1986,N_1896);
xor U2128 (N_2128,N_1886,N_1863);
and U2129 (N_2129,N_1865,N_1917);
nand U2130 (N_2130,N_1847,N_2049);
nand U2131 (N_2131,N_2054,N_2053);
or U2132 (N_2132,N_2018,N_1926);
xor U2133 (N_2133,N_1930,N_1976);
or U2134 (N_2134,N_2011,N_1979);
or U2135 (N_2135,N_1862,N_1941);
or U2136 (N_2136,N_2058,N_1883);
nand U2137 (N_2137,N_1924,N_1808);
or U2138 (N_2138,N_1902,N_1916);
xnor U2139 (N_2139,N_2006,N_1963);
nor U2140 (N_2140,N_2099,N_1816);
xor U2141 (N_2141,N_1905,N_1844);
xor U2142 (N_2142,N_1861,N_2089);
and U2143 (N_2143,N_1955,N_1860);
xor U2144 (N_2144,N_2087,N_1867);
and U2145 (N_2145,N_2002,N_1984);
nand U2146 (N_2146,N_2079,N_2015);
nand U2147 (N_2147,N_2040,N_1937);
or U2148 (N_2148,N_2035,N_1969);
or U2149 (N_2149,N_1880,N_2025);
or U2150 (N_2150,N_1956,N_1813);
nand U2151 (N_2151,N_1911,N_1804);
nor U2152 (N_2152,N_1836,N_1831);
xnor U2153 (N_2153,N_1996,N_1991);
and U2154 (N_2154,N_1971,N_1980);
xnor U2155 (N_2155,N_1822,N_1953);
nor U2156 (N_2156,N_1977,N_1964);
and U2157 (N_2157,N_2019,N_1933);
and U2158 (N_2158,N_1846,N_1864);
or U2159 (N_2159,N_1879,N_2094);
xnor U2160 (N_2160,N_1841,N_1938);
or U2161 (N_2161,N_1887,N_2021);
nand U2162 (N_2162,N_2095,N_1853);
nand U2163 (N_2163,N_1966,N_1849);
xor U2164 (N_2164,N_1802,N_1954);
and U2165 (N_2165,N_1892,N_1974);
nor U2166 (N_2166,N_1951,N_2047);
xor U2167 (N_2167,N_1852,N_1998);
nand U2168 (N_2168,N_2096,N_2084);
and U2169 (N_2169,N_1894,N_2004);
nor U2170 (N_2170,N_2092,N_2046);
nor U2171 (N_2171,N_2027,N_1840);
or U2172 (N_2172,N_1923,N_1871);
nand U2173 (N_2173,N_1897,N_1859);
nor U2174 (N_2174,N_1970,N_1810);
nand U2175 (N_2175,N_2083,N_2097);
nor U2176 (N_2176,N_2001,N_2010);
and U2177 (N_2177,N_2081,N_1812);
nor U2178 (N_2178,N_2064,N_2041);
xnor U2179 (N_2179,N_1878,N_1913);
xor U2180 (N_2180,N_2061,N_1838);
xnor U2181 (N_2181,N_1939,N_1909);
or U2182 (N_2182,N_2039,N_2051);
and U2183 (N_2183,N_1826,N_1893);
nand U2184 (N_2184,N_1842,N_1817);
xnor U2185 (N_2185,N_2086,N_1990);
nor U2186 (N_2186,N_2014,N_1935);
nor U2187 (N_2187,N_1940,N_2009);
or U2188 (N_2188,N_1805,N_1885);
nor U2189 (N_2189,N_1901,N_1918);
and U2190 (N_2190,N_1988,N_1891);
and U2191 (N_2191,N_2080,N_1931);
or U2192 (N_2192,N_1912,N_2044);
and U2193 (N_2193,N_1855,N_2029);
and U2194 (N_2194,N_1950,N_1925);
xor U2195 (N_2195,N_1958,N_1825);
nor U2196 (N_2196,N_1967,N_1947);
or U2197 (N_2197,N_1907,N_1877);
nand U2198 (N_2198,N_1828,N_1973);
or U2199 (N_2199,N_1876,N_1888);
and U2200 (N_2200,N_1866,N_2085);
nand U2201 (N_2201,N_1830,N_1989);
or U2202 (N_2202,N_2028,N_1936);
nor U2203 (N_2203,N_1803,N_1978);
nor U2204 (N_2204,N_1942,N_2066);
nand U2205 (N_2205,N_2042,N_1884);
nor U2206 (N_2206,N_2075,N_1818);
nor U2207 (N_2207,N_1995,N_1898);
xnor U2208 (N_2208,N_1850,N_1994);
xor U2209 (N_2209,N_1854,N_1839);
and U2210 (N_2210,N_2073,N_1959);
nand U2211 (N_2211,N_1921,N_1960);
xnor U2212 (N_2212,N_2020,N_2037);
nor U2213 (N_2213,N_1957,N_2057);
and U2214 (N_2214,N_1869,N_1928);
and U2215 (N_2215,N_1858,N_1944);
nor U2216 (N_2216,N_1999,N_1832);
nor U2217 (N_2217,N_1833,N_1824);
nor U2218 (N_2218,N_1992,N_1843);
nand U2219 (N_2219,N_1949,N_2067);
or U2220 (N_2220,N_1945,N_2031);
and U2221 (N_2221,N_2000,N_1835);
nand U2222 (N_2222,N_1875,N_1914);
nor U2223 (N_2223,N_1900,N_1903);
and U2224 (N_2224,N_2038,N_2082);
and U2225 (N_2225,N_1806,N_2088);
nand U2226 (N_2226,N_1920,N_1981);
and U2227 (N_2227,N_1927,N_1993);
xnor U2228 (N_2228,N_1968,N_1857);
and U2229 (N_2229,N_1961,N_2016);
xor U2230 (N_2230,N_2013,N_1821);
or U2231 (N_2231,N_1997,N_2077);
and U2232 (N_2232,N_1823,N_1811);
nand U2233 (N_2233,N_2090,N_1851);
nor U2234 (N_2234,N_2030,N_1815);
xnor U2235 (N_2235,N_1906,N_2060);
nand U2236 (N_2236,N_2050,N_1908);
or U2237 (N_2237,N_1890,N_2043);
nand U2238 (N_2238,N_2059,N_2055);
xnor U2239 (N_2239,N_1946,N_1856);
or U2240 (N_2240,N_1848,N_2033);
nand U2241 (N_2241,N_2012,N_2036);
nand U2242 (N_2242,N_2068,N_1845);
xor U2243 (N_2243,N_1975,N_1874);
nand U2244 (N_2244,N_1870,N_1819);
and U2245 (N_2245,N_2062,N_2063);
xor U2246 (N_2246,N_2076,N_1800);
xnor U2247 (N_2247,N_1972,N_1899);
xor U2248 (N_2248,N_1910,N_1932);
xor U2249 (N_2249,N_1807,N_2003);
nand U2250 (N_2250,N_1920,N_1857);
or U2251 (N_2251,N_1976,N_2015);
nor U2252 (N_2252,N_2063,N_2064);
xor U2253 (N_2253,N_1926,N_2003);
and U2254 (N_2254,N_1814,N_1886);
nand U2255 (N_2255,N_1961,N_2009);
xor U2256 (N_2256,N_1867,N_1856);
or U2257 (N_2257,N_1821,N_2028);
nand U2258 (N_2258,N_1892,N_1863);
nand U2259 (N_2259,N_1858,N_1961);
xor U2260 (N_2260,N_1852,N_1829);
xnor U2261 (N_2261,N_1884,N_2083);
nand U2262 (N_2262,N_1819,N_1921);
nand U2263 (N_2263,N_1818,N_1836);
and U2264 (N_2264,N_2077,N_2008);
nand U2265 (N_2265,N_2065,N_1838);
nand U2266 (N_2266,N_2040,N_1896);
nand U2267 (N_2267,N_1968,N_2003);
nand U2268 (N_2268,N_1892,N_1929);
nor U2269 (N_2269,N_2084,N_2010);
xor U2270 (N_2270,N_1971,N_1935);
and U2271 (N_2271,N_1824,N_2086);
xor U2272 (N_2272,N_2090,N_1843);
xor U2273 (N_2273,N_1894,N_1864);
xnor U2274 (N_2274,N_2069,N_1894);
nor U2275 (N_2275,N_2066,N_1975);
xor U2276 (N_2276,N_1937,N_2005);
and U2277 (N_2277,N_1946,N_1901);
xor U2278 (N_2278,N_1987,N_1979);
or U2279 (N_2279,N_2018,N_2045);
nand U2280 (N_2280,N_1838,N_2013);
nand U2281 (N_2281,N_1907,N_1859);
or U2282 (N_2282,N_1956,N_2056);
or U2283 (N_2283,N_2003,N_2090);
xnor U2284 (N_2284,N_2049,N_2007);
xor U2285 (N_2285,N_2007,N_1982);
and U2286 (N_2286,N_1954,N_1879);
nor U2287 (N_2287,N_1918,N_1915);
or U2288 (N_2288,N_1918,N_1825);
nand U2289 (N_2289,N_1900,N_1815);
nor U2290 (N_2290,N_2096,N_1832);
and U2291 (N_2291,N_1941,N_2014);
xor U2292 (N_2292,N_1992,N_2063);
xor U2293 (N_2293,N_1933,N_2062);
xnor U2294 (N_2294,N_1825,N_1805);
or U2295 (N_2295,N_1929,N_1939);
or U2296 (N_2296,N_1853,N_2029);
nand U2297 (N_2297,N_1943,N_1867);
xnor U2298 (N_2298,N_2012,N_2066);
or U2299 (N_2299,N_1845,N_1988);
nand U2300 (N_2300,N_2097,N_1852);
or U2301 (N_2301,N_1950,N_1833);
and U2302 (N_2302,N_1842,N_1921);
and U2303 (N_2303,N_1851,N_2023);
and U2304 (N_2304,N_1979,N_2095);
or U2305 (N_2305,N_2092,N_2004);
nand U2306 (N_2306,N_1870,N_1863);
or U2307 (N_2307,N_1949,N_2086);
nand U2308 (N_2308,N_1926,N_2050);
or U2309 (N_2309,N_1805,N_1853);
nand U2310 (N_2310,N_2012,N_1861);
nand U2311 (N_2311,N_2038,N_1870);
nand U2312 (N_2312,N_1822,N_2082);
nand U2313 (N_2313,N_1862,N_2064);
xor U2314 (N_2314,N_1874,N_2011);
or U2315 (N_2315,N_2064,N_1980);
nand U2316 (N_2316,N_1823,N_1878);
xnor U2317 (N_2317,N_2061,N_1939);
xor U2318 (N_2318,N_2025,N_1854);
or U2319 (N_2319,N_2043,N_1885);
nor U2320 (N_2320,N_1837,N_2034);
or U2321 (N_2321,N_2010,N_1921);
or U2322 (N_2322,N_1981,N_2053);
and U2323 (N_2323,N_1923,N_1827);
nor U2324 (N_2324,N_1828,N_1914);
or U2325 (N_2325,N_1865,N_1804);
and U2326 (N_2326,N_1946,N_1858);
or U2327 (N_2327,N_2030,N_1869);
xor U2328 (N_2328,N_2087,N_1822);
xor U2329 (N_2329,N_2006,N_1832);
nor U2330 (N_2330,N_2006,N_2062);
nand U2331 (N_2331,N_1987,N_2018);
xor U2332 (N_2332,N_2081,N_1982);
nand U2333 (N_2333,N_2089,N_1926);
xnor U2334 (N_2334,N_1888,N_1922);
xnor U2335 (N_2335,N_1928,N_1824);
xor U2336 (N_2336,N_1891,N_1802);
and U2337 (N_2337,N_2061,N_1932);
nand U2338 (N_2338,N_1941,N_1848);
and U2339 (N_2339,N_2015,N_1904);
xnor U2340 (N_2340,N_2047,N_1823);
nand U2341 (N_2341,N_1833,N_1843);
nor U2342 (N_2342,N_2012,N_1862);
and U2343 (N_2343,N_1897,N_2000);
or U2344 (N_2344,N_2065,N_1934);
nor U2345 (N_2345,N_1918,N_1851);
nor U2346 (N_2346,N_1820,N_1948);
xnor U2347 (N_2347,N_2058,N_1817);
xor U2348 (N_2348,N_1815,N_1803);
or U2349 (N_2349,N_1902,N_1828);
and U2350 (N_2350,N_1821,N_1993);
xor U2351 (N_2351,N_1800,N_1815);
and U2352 (N_2352,N_2033,N_1984);
or U2353 (N_2353,N_2092,N_1938);
nand U2354 (N_2354,N_2009,N_2055);
nand U2355 (N_2355,N_2074,N_1848);
nand U2356 (N_2356,N_1880,N_1878);
nor U2357 (N_2357,N_1866,N_1950);
and U2358 (N_2358,N_1892,N_1887);
and U2359 (N_2359,N_2087,N_1897);
nand U2360 (N_2360,N_1934,N_2016);
xor U2361 (N_2361,N_1865,N_1895);
and U2362 (N_2362,N_1923,N_2081);
nor U2363 (N_2363,N_1933,N_1924);
nand U2364 (N_2364,N_2035,N_1861);
nor U2365 (N_2365,N_1803,N_1881);
or U2366 (N_2366,N_1852,N_1889);
or U2367 (N_2367,N_1815,N_2059);
or U2368 (N_2368,N_1976,N_2040);
xor U2369 (N_2369,N_2045,N_1816);
and U2370 (N_2370,N_1912,N_1957);
nor U2371 (N_2371,N_1939,N_1825);
or U2372 (N_2372,N_1997,N_1982);
and U2373 (N_2373,N_2071,N_1891);
nand U2374 (N_2374,N_1804,N_1997);
or U2375 (N_2375,N_1825,N_2068);
nand U2376 (N_2376,N_1854,N_1891);
or U2377 (N_2377,N_2047,N_1995);
nand U2378 (N_2378,N_1995,N_1990);
nand U2379 (N_2379,N_2085,N_1973);
nor U2380 (N_2380,N_1924,N_1809);
or U2381 (N_2381,N_1860,N_1895);
or U2382 (N_2382,N_1978,N_2006);
nand U2383 (N_2383,N_1898,N_1813);
and U2384 (N_2384,N_1949,N_1929);
nand U2385 (N_2385,N_1868,N_1841);
or U2386 (N_2386,N_2052,N_2085);
and U2387 (N_2387,N_1861,N_1835);
xor U2388 (N_2388,N_2059,N_1836);
or U2389 (N_2389,N_1927,N_2097);
or U2390 (N_2390,N_1921,N_1814);
nand U2391 (N_2391,N_1928,N_1976);
and U2392 (N_2392,N_2073,N_1884);
or U2393 (N_2393,N_2038,N_2010);
nand U2394 (N_2394,N_1961,N_1991);
or U2395 (N_2395,N_1936,N_2051);
and U2396 (N_2396,N_2018,N_1852);
nand U2397 (N_2397,N_2089,N_1862);
xor U2398 (N_2398,N_2076,N_1979);
nor U2399 (N_2399,N_1875,N_2085);
nand U2400 (N_2400,N_2167,N_2112);
or U2401 (N_2401,N_2139,N_2352);
xnor U2402 (N_2402,N_2182,N_2135);
nand U2403 (N_2403,N_2117,N_2265);
xor U2404 (N_2404,N_2279,N_2122);
nor U2405 (N_2405,N_2192,N_2118);
and U2406 (N_2406,N_2170,N_2188);
xor U2407 (N_2407,N_2123,N_2399);
nor U2408 (N_2408,N_2321,N_2247);
and U2409 (N_2409,N_2143,N_2371);
or U2410 (N_2410,N_2290,N_2103);
and U2411 (N_2411,N_2193,N_2354);
or U2412 (N_2412,N_2387,N_2238);
xor U2413 (N_2413,N_2115,N_2314);
or U2414 (N_2414,N_2224,N_2319);
nor U2415 (N_2415,N_2308,N_2176);
nand U2416 (N_2416,N_2304,N_2240);
nor U2417 (N_2417,N_2154,N_2160);
and U2418 (N_2418,N_2250,N_2231);
nand U2419 (N_2419,N_2237,N_2328);
nor U2420 (N_2420,N_2269,N_2178);
xor U2421 (N_2421,N_2104,N_2180);
nor U2422 (N_2422,N_2396,N_2125);
nand U2423 (N_2423,N_2145,N_2196);
xnor U2424 (N_2424,N_2305,N_2335);
or U2425 (N_2425,N_2213,N_2191);
or U2426 (N_2426,N_2339,N_2373);
nand U2427 (N_2427,N_2347,N_2174);
nor U2428 (N_2428,N_2183,N_2348);
xnor U2429 (N_2429,N_2368,N_2198);
xor U2430 (N_2430,N_2282,N_2393);
nor U2431 (N_2431,N_2359,N_2260);
nand U2432 (N_2432,N_2206,N_2340);
and U2433 (N_2433,N_2259,N_2173);
nor U2434 (N_2434,N_2380,N_2195);
nand U2435 (N_2435,N_2220,N_2249);
nor U2436 (N_2436,N_2361,N_2200);
nor U2437 (N_2437,N_2254,N_2310);
or U2438 (N_2438,N_2275,N_2293);
or U2439 (N_2439,N_2146,N_2108);
nor U2440 (N_2440,N_2280,N_2201);
or U2441 (N_2441,N_2207,N_2208);
or U2442 (N_2442,N_2150,N_2185);
or U2443 (N_2443,N_2203,N_2360);
and U2444 (N_2444,N_2285,N_2219);
or U2445 (N_2445,N_2131,N_2327);
nor U2446 (N_2446,N_2394,N_2379);
and U2447 (N_2447,N_2107,N_2243);
and U2448 (N_2448,N_2148,N_2391);
nand U2449 (N_2449,N_2311,N_2333);
xnor U2450 (N_2450,N_2168,N_2356);
and U2451 (N_2451,N_2113,N_2245);
or U2452 (N_2452,N_2120,N_2370);
or U2453 (N_2453,N_2345,N_2253);
and U2454 (N_2454,N_2149,N_2133);
or U2455 (N_2455,N_2124,N_2258);
nor U2456 (N_2456,N_2376,N_2332);
nand U2457 (N_2457,N_2251,N_2341);
or U2458 (N_2458,N_2157,N_2186);
nand U2459 (N_2459,N_2129,N_2337);
nor U2460 (N_2460,N_2181,N_2385);
xnor U2461 (N_2461,N_2114,N_2355);
and U2462 (N_2462,N_2302,N_2241);
and U2463 (N_2463,N_2344,N_2246);
and U2464 (N_2464,N_2102,N_2155);
nor U2465 (N_2465,N_2227,N_2236);
or U2466 (N_2466,N_2262,N_2294);
or U2467 (N_2467,N_2144,N_2346);
nand U2468 (N_2468,N_2316,N_2276);
or U2469 (N_2469,N_2357,N_2273);
nand U2470 (N_2470,N_2242,N_2386);
or U2471 (N_2471,N_2306,N_2287);
nand U2472 (N_2472,N_2381,N_2100);
nand U2473 (N_2473,N_2329,N_2256);
and U2474 (N_2474,N_2233,N_2126);
xor U2475 (N_2475,N_2187,N_2334);
or U2476 (N_2476,N_2110,N_2197);
xor U2477 (N_2477,N_2106,N_2392);
and U2478 (N_2478,N_2179,N_2267);
nor U2479 (N_2479,N_2121,N_2277);
or U2480 (N_2480,N_2291,N_2239);
or U2481 (N_2481,N_2172,N_2384);
xnor U2482 (N_2482,N_2209,N_2375);
or U2483 (N_2483,N_2136,N_2390);
or U2484 (N_2484,N_2257,N_2278);
nand U2485 (N_2485,N_2270,N_2169);
nor U2486 (N_2486,N_2322,N_2189);
nor U2487 (N_2487,N_2140,N_2137);
or U2488 (N_2488,N_2217,N_2336);
and U2489 (N_2489,N_2313,N_2252);
xor U2490 (N_2490,N_2138,N_2323);
or U2491 (N_2491,N_2315,N_2266);
nor U2492 (N_2492,N_2382,N_2301);
nand U2493 (N_2493,N_2156,N_2297);
xnor U2494 (N_2494,N_2216,N_2378);
and U2495 (N_2495,N_2397,N_2159);
or U2496 (N_2496,N_2128,N_2369);
nor U2497 (N_2497,N_2289,N_2109);
xor U2498 (N_2498,N_2307,N_2205);
and U2499 (N_2499,N_2184,N_2152);
nor U2500 (N_2500,N_2320,N_2215);
nand U2501 (N_2501,N_2388,N_2210);
nor U2502 (N_2502,N_2300,N_2286);
nor U2503 (N_2503,N_2367,N_2119);
xor U2504 (N_2504,N_2338,N_2325);
nand U2505 (N_2505,N_2317,N_2324);
nand U2506 (N_2506,N_2363,N_2212);
nand U2507 (N_2507,N_2343,N_2350);
nand U2508 (N_2508,N_2202,N_2295);
nor U2509 (N_2509,N_2141,N_2271);
xor U2510 (N_2510,N_2264,N_2312);
and U2511 (N_2511,N_2225,N_2353);
nand U2512 (N_2512,N_2226,N_2101);
xor U2513 (N_2513,N_2134,N_2166);
nor U2514 (N_2514,N_2298,N_2358);
or U2515 (N_2515,N_2248,N_2366);
or U2516 (N_2516,N_2164,N_2362);
nor U2517 (N_2517,N_2281,N_2158);
or U2518 (N_2518,N_2177,N_2309);
and U2519 (N_2519,N_2221,N_2318);
nand U2520 (N_2520,N_2165,N_2283);
xnor U2521 (N_2521,N_2234,N_2364);
and U2522 (N_2522,N_2244,N_2153);
or U2523 (N_2523,N_2171,N_2342);
nand U2524 (N_2524,N_2383,N_2105);
and U2525 (N_2525,N_2398,N_2349);
nor U2526 (N_2526,N_2228,N_2274);
and U2527 (N_2527,N_2142,N_2377);
and U2528 (N_2528,N_2163,N_2351);
nor U2529 (N_2529,N_2284,N_2130);
or U2530 (N_2530,N_2389,N_2223);
and U2531 (N_2531,N_2190,N_2296);
xnor U2532 (N_2532,N_2263,N_2218);
xnor U2533 (N_2533,N_2211,N_2175);
nor U2534 (N_2534,N_2116,N_2214);
nand U2535 (N_2535,N_2374,N_2194);
nand U2536 (N_2536,N_2162,N_2232);
and U2537 (N_2537,N_2365,N_2204);
xor U2538 (N_2538,N_2199,N_2272);
nand U2539 (N_2539,N_2261,N_2132);
nor U2540 (N_2540,N_2255,N_2229);
nand U2541 (N_2541,N_2395,N_2111);
or U2542 (N_2542,N_2127,N_2372);
or U2543 (N_2543,N_2161,N_2230);
xnor U2544 (N_2544,N_2268,N_2235);
or U2545 (N_2545,N_2331,N_2326);
and U2546 (N_2546,N_2330,N_2292);
xnor U2547 (N_2547,N_2147,N_2288);
nor U2548 (N_2548,N_2303,N_2151);
or U2549 (N_2549,N_2299,N_2222);
nor U2550 (N_2550,N_2320,N_2382);
nor U2551 (N_2551,N_2331,N_2157);
xnor U2552 (N_2552,N_2385,N_2394);
nand U2553 (N_2553,N_2196,N_2278);
xnor U2554 (N_2554,N_2119,N_2251);
nor U2555 (N_2555,N_2204,N_2266);
nand U2556 (N_2556,N_2146,N_2180);
xnor U2557 (N_2557,N_2381,N_2129);
and U2558 (N_2558,N_2188,N_2319);
nor U2559 (N_2559,N_2334,N_2259);
nand U2560 (N_2560,N_2383,N_2343);
nand U2561 (N_2561,N_2258,N_2249);
and U2562 (N_2562,N_2302,N_2368);
or U2563 (N_2563,N_2238,N_2379);
nor U2564 (N_2564,N_2278,N_2185);
or U2565 (N_2565,N_2377,N_2145);
nor U2566 (N_2566,N_2221,N_2249);
xor U2567 (N_2567,N_2131,N_2114);
xor U2568 (N_2568,N_2142,N_2295);
nand U2569 (N_2569,N_2214,N_2139);
xor U2570 (N_2570,N_2144,N_2380);
and U2571 (N_2571,N_2388,N_2201);
nor U2572 (N_2572,N_2290,N_2115);
and U2573 (N_2573,N_2171,N_2222);
nor U2574 (N_2574,N_2315,N_2374);
xnor U2575 (N_2575,N_2235,N_2312);
nor U2576 (N_2576,N_2333,N_2270);
nor U2577 (N_2577,N_2319,N_2299);
and U2578 (N_2578,N_2183,N_2329);
or U2579 (N_2579,N_2364,N_2156);
xor U2580 (N_2580,N_2105,N_2266);
nor U2581 (N_2581,N_2345,N_2341);
nand U2582 (N_2582,N_2160,N_2216);
xnor U2583 (N_2583,N_2275,N_2103);
or U2584 (N_2584,N_2336,N_2125);
or U2585 (N_2585,N_2108,N_2133);
nor U2586 (N_2586,N_2163,N_2132);
nand U2587 (N_2587,N_2213,N_2385);
xor U2588 (N_2588,N_2280,N_2227);
nor U2589 (N_2589,N_2325,N_2316);
or U2590 (N_2590,N_2316,N_2252);
nand U2591 (N_2591,N_2284,N_2231);
xnor U2592 (N_2592,N_2163,N_2226);
or U2593 (N_2593,N_2149,N_2146);
or U2594 (N_2594,N_2304,N_2290);
nand U2595 (N_2595,N_2277,N_2199);
and U2596 (N_2596,N_2169,N_2323);
and U2597 (N_2597,N_2380,N_2321);
and U2598 (N_2598,N_2174,N_2337);
or U2599 (N_2599,N_2334,N_2124);
and U2600 (N_2600,N_2284,N_2182);
nand U2601 (N_2601,N_2328,N_2365);
xnor U2602 (N_2602,N_2325,N_2326);
nand U2603 (N_2603,N_2293,N_2372);
xor U2604 (N_2604,N_2258,N_2262);
and U2605 (N_2605,N_2386,N_2124);
or U2606 (N_2606,N_2169,N_2333);
nor U2607 (N_2607,N_2347,N_2109);
nor U2608 (N_2608,N_2221,N_2294);
or U2609 (N_2609,N_2217,N_2165);
nand U2610 (N_2610,N_2227,N_2259);
nand U2611 (N_2611,N_2147,N_2270);
and U2612 (N_2612,N_2100,N_2271);
nor U2613 (N_2613,N_2271,N_2241);
nor U2614 (N_2614,N_2338,N_2300);
nand U2615 (N_2615,N_2141,N_2178);
nand U2616 (N_2616,N_2128,N_2385);
nand U2617 (N_2617,N_2395,N_2275);
and U2618 (N_2618,N_2366,N_2390);
nor U2619 (N_2619,N_2256,N_2226);
or U2620 (N_2620,N_2394,N_2231);
xnor U2621 (N_2621,N_2228,N_2354);
nand U2622 (N_2622,N_2325,N_2252);
nand U2623 (N_2623,N_2250,N_2304);
nor U2624 (N_2624,N_2315,N_2127);
and U2625 (N_2625,N_2362,N_2179);
xnor U2626 (N_2626,N_2369,N_2386);
or U2627 (N_2627,N_2222,N_2373);
or U2628 (N_2628,N_2210,N_2351);
nand U2629 (N_2629,N_2257,N_2274);
xnor U2630 (N_2630,N_2334,N_2172);
and U2631 (N_2631,N_2325,N_2116);
or U2632 (N_2632,N_2329,N_2393);
xnor U2633 (N_2633,N_2380,N_2386);
and U2634 (N_2634,N_2119,N_2266);
nand U2635 (N_2635,N_2217,N_2188);
and U2636 (N_2636,N_2333,N_2204);
xnor U2637 (N_2637,N_2296,N_2269);
and U2638 (N_2638,N_2321,N_2374);
nand U2639 (N_2639,N_2125,N_2267);
and U2640 (N_2640,N_2293,N_2390);
xor U2641 (N_2641,N_2297,N_2143);
and U2642 (N_2642,N_2115,N_2145);
xor U2643 (N_2643,N_2359,N_2210);
or U2644 (N_2644,N_2352,N_2342);
or U2645 (N_2645,N_2298,N_2104);
nor U2646 (N_2646,N_2299,N_2340);
nand U2647 (N_2647,N_2277,N_2141);
nor U2648 (N_2648,N_2200,N_2116);
or U2649 (N_2649,N_2153,N_2339);
xnor U2650 (N_2650,N_2227,N_2211);
or U2651 (N_2651,N_2261,N_2194);
and U2652 (N_2652,N_2135,N_2386);
and U2653 (N_2653,N_2148,N_2242);
and U2654 (N_2654,N_2357,N_2134);
xnor U2655 (N_2655,N_2179,N_2149);
or U2656 (N_2656,N_2140,N_2355);
nand U2657 (N_2657,N_2336,N_2153);
nand U2658 (N_2658,N_2288,N_2282);
and U2659 (N_2659,N_2165,N_2373);
or U2660 (N_2660,N_2199,N_2287);
nand U2661 (N_2661,N_2224,N_2195);
nand U2662 (N_2662,N_2322,N_2106);
or U2663 (N_2663,N_2120,N_2248);
and U2664 (N_2664,N_2331,N_2176);
and U2665 (N_2665,N_2342,N_2324);
nand U2666 (N_2666,N_2368,N_2184);
nand U2667 (N_2667,N_2249,N_2393);
nand U2668 (N_2668,N_2248,N_2140);
nand U2669 (N_2669,N_2398,N_2221);
nand U2670 (N_2670,N_2328,N_2174);
nor U2671 (N_2671,N_2305,N_2272);
nand U2672 (N_2672,N_2312,N_2173);
xor U2673 (N_2673,N_2350,N_2378);
nor U2674 (N_2674,N_2348,N_2125);
or U2675 (N_2675,N_2321,N_2301);
and U2676 (N_2676,N_2336,N_2138);
nor U2677 (N_2677,N_2288,N_2336);
nand U2678 (N_2678,N_2277,N_2395);
and U2679 (N_2679,N_2262,N_2275);
nor U2680 (N_2680,N_2393,N_2213);
xnor U2681 (N_2681,N_2125,N_2328);
or U2682 (N_2682,N_2382,N_2345);
and U2683 (N_2683,N_2231,N_2266);
and U2684 (N_2684,N_2310,N_2226);
nand U2685 (N_2685,N_2390,N_2130);
or U2686 (N_2686,N_2306,N_2245);
nor U2687 (N_2687,N_2365,N_2362);
or U2688 (N_2688,N_2395,N_2113);
or U2689 (N_2689,N_2174,N_2253);
nand U2690 (N_2690,N_2346,N_2393);
nand U2691 (N_2691,N_2164,N_2145);
nor U2692 (N_2692,N_2158,N_2320);
xnor U2693 (N_2693,N_2204,N_2182);
nor U2694 (N_2694,N_2148,N_2236);
or U2695 (N_2695,N_2211,N_2189);
or U2696 (N_2696,N_2231,N_2375);
nand U2697 (N_2697,N_2206,N_2163);
nor U2698 (N_2698,N_2179,N_2333);
nand U2699 (N_2699,N_2166,N_2348);
xor U2700 (N_2700,N_2593,N_2519);
and U2701 (N_2701,N_2464,N_2481);
xor U2702 (N_2702,N_2613,N_2402);
nand U2703 (N_2703,N_2559,N_2618);
and U2704 (N_2704,N_2443,N_2465);
nor U2705 (N_2705,N_2694,N_2672);
and U2706 (N_2706,N_2461,N_2403);
nor U2707 (N_2707,N_2479,N_2596);
xnor U2708 (N_2708,N_2466,N_2420);
nor U2709 (N_2709,N_2523,N_2592);
or U2710 (N_2710,N_2696,N_2631);
and U2711 (N_2711,N_2572,N_2584);
nor U2712 (N_2712,N_2598,N_2690);
nand U2713 (N_2713,N_2543,N_2460);
xnor U2714 (N_2714,N_2676,N_2547);
xnor U2715 (N_2715,N_2662,N_2580);
and U2716 (N_2716,N_2591,N_2432);
or U2717 (N_2717,N_2527,N_2661);
xor U2718 (N_2718,N_2561,N_2655);
nand U2719 (N_2719,N_2495,N_2525);
and U2720 (N_2720,N_2668,N_2484);
xnor U2721 (N_2721,N_2448,N_2638);
and U2722 (N_2722,N_2681,N_2585);
xnor U2723 (N_2723,N_2612,N_2656);
xor U2724 (N_2724,N_2562,N_2490);
and U2725 (N_2725,N_2439,N_2588);
xnor U2726 (N_2726,N_2502,N_2521);
xnor U2727 (N_2727,N_2671,N_2685);
nand U2728 (N_2728,N_2552,N_2548);
or U2729 (N_2729,N_2575,N_2624);
nor U2730 (N_2730,N_2515,N_2440);
and U2731 (N_2731,N_2467,N_2433);
xor U2732 (N_2732,N_2693,N_2601);
nand U2733 (N_2733,N_2582,N_2607);
and U2734 (N_2734,N_2677,N_2493);
and U2735 (N_2735,N_2546,N_2517);
or U2736 (N_2736,N_2608,N_2427);
xnor U2737 (N_2737,N_2435,N_2657);
xnor U2738 (N_2738,N_2497,N_2565);
xnor U2739 (N_2739,N_2508,N_2634);
xnor U2740 (N_2740,N_2578,N_2589);
xor U2741 (N_2741,N_2615,N_2650);
or U2742 (N_2742,N_2472,N_2423);
nand U2743 (N_2743,N_2628,N_2500);
nand U2744 (N_2744,N_2452,N_2666);
xnor U2745 (N_2745,N_2579,N_2529);
nor U2746 (N_2746,N_2573,N_2649);
nor U2747 (N_2747,N_2689,N_2621);
and U2748 (N_2748,N_2444,N_2669);
or U2749 (N_2749,N_2645,N_2471);
xnor U2750 (N_2750,N_2410,N_2533);
xor U2751 (N_2751,N_2453,N_2686);
or U2752 (N_2752,N_2470,N_2475);
nor U2753 (N_2753,N_2688,N_2425);
or U2754 (N_2754,N_2412,N_2658);
nand U2755 (N_2755,N_2407,N_2473);
xnor U2756 (N_2756,N_2447,N_2544);
and U2757 (N_2757,N_2697,N_2554);
or U2758 (N_2758,N_2434,N_2557);
xor U2759 (N_2759,N_2408,N_2503);
or U2760 (N_2760,N_2437,N_2530);
nand U2761 (N_2761,N_2426,N_2587);
and U2762 (N_2762,N_2683,N_2617);
or U2763 (N_2763,N_2455,N_2518);
nor U2764 (N_2764,N_2586,N_2468);
xor U2765 (N_2765,N_2630,N_2698);
or U2766 (N_2766,N_2663,N_2458);
nor U2767 (N_2767,N_2692,N_2441);
nand U2768 (N_2768,N_2651,N_2687);
or U2769 (N_2769,N_2482,N_2405);
and U2770 (N_2770,N_2413,N_2627);
or U2771 (N_2771,N_2513,N_2602);
xnor U2772 (N_2772,N_2563,N_2476);
or U2773 (N_2773,N_2599,N_2480);
and U2774 (N_2774,N_2637,N_2636);
xnor U2775 (N_2775,N_2541,N_2501);
xnor U2776 (N_2776,N_2526,N_2597);
and U2777 (N_2777,N_2577,N_2610);
xor U2778 (N_2778,N_2507,N_2684);
nor U2779 (N_2779,N_2569,N_2556);
xnor U2780 (N_2780,N_2648,N_2635);
nor U2781 (N_2781,N_2675,N_2643);
nand U2782 (N_2782,N_2673,N_2489);
nor U2783 (N_2783,N_2566,N_2600);
xnor U2784 (N_2784,N_2400,N_2477);
nor U2785 (N_2785,N_2505,N_2524);
or U2786 (N_2786,N_2659,N_2616);
nor U2787 (N_2787,N_2611,N_2603);
xnor U2788 (N_2788,N_2539,N_2633);
xnor U2789 (N_2789,N_2504,N_2419);
and U2790 (N_2790,N_2581,N_2674);
or U2791 (N_2791,N_2632,N_2506);
nor U2792 (N_2792,N_2516,N_2654);
or U2793 (N_2793,N_2571,N_2415);
or U2794 (N_2794,N_2535,N_2605);
nor U2795 (N_2795,N_2641,N_2642);
or U2796 (N_2796,N_2457,N_2438);
xnor U2797 (N_2797,N_2646,N_2487);
or U2798 (N_2798,N_2553,N_2644);
nor U2799 (N_2799,N_2512,N_2604);
nor U2800 (N_2800,N_2449,N_2558);
or U2801 (N_2801,N_2492,N_2665);
nand U2802 (N_2802,N_2564,N_2456);
and U2803 (N_2803,N_2478,N_2430);
and U2804 (N_2804,N_2532,N_2670);
nor U2805 (N_2805,N_2647,N_2450);
xnor U2806 (N_2806,N_2560,N_2417);
xnor U2807 (N_2807,N_2620,N_2424);
and U2808 (N_2808,N_2469,N_2451);
nand U2809 (N_2809,N_2680,N_2462);
nor U2810 (N_2810,N_2538,N_2691);
and U2811 (N_2811,N_2446,N_2574);
xor U2812 (N_2812,N_2414,N_2629);
nor U2813 (N_2813,N_2679,N_2428);
and U2814 (N_2814,N_2522,N_2549);
and U2815 (N_2815,N_2609,N_2594);
nor U2816 (N_2816,N_2510,N_2550);
nand U2817 (N_2817,N_2528,N_2422);
and U2818 (N_2818,N_2695,N_2606);
xnor U2819 (N_2819,N_2639,N_2699);
or U2820 (N_2820,N_2653,N_2622);
xor U2821 (N_2821,N_2614,N_2485);
and U2822 (N_2822,N_2595,N_2488);
or U2823 (N_2823,N_2625,N_2498);
nand U2824 (N_2824,N_2551,N_2626);
nor U2825 (N_2825,N_2499,N_2509);
xnor U2826 (N_2826,N_2640,N_2623);
nor U2827 (N_2827,N_2411,N_2496);
nand U2828 (N_2828,N_2442,N_2534);
nand U2829 (N_2829,N_2431,N_2491);
xnor U2830 (N_2830,N_2583,N_2531);
or U2831 (N_2831,N_2483,N_2445);
xor U2832 (N_2832,N_2416,N_2436);
xnor U2833 (N_2833,N_2409,N_2418);
nand U2834 (N_2834,N_2619,N_2664);
and U2835 (N_2835,N_2429,N_2652);
nor U2836 (N_2836,N_2667,N_2421);
or U2837 (N_2837,N_2486,N_2537);
nor U2838 (N_2838,N_2540,N_2545);
xnor U2839 (N_2839,N_2590,N_2520);
and U2840 (N_2840,N_2454,N_2678);
nor U2841 (N_2841,N_2494,N_2555);
nor U2842 (N_2842,N_2542,N_2511);
nor U2843 (N_2843,N_2463,N_2568);
or U2844 (N_2844,N_2459,N_2660);
and U2845 (N_2845,N_2514,N_2406);
nand U2846 (N_2846,N_2401,N_2536);
and U2847 (N_2847,N_2576,N_2682);
nor U2848 (N_2848,N_2570,N_2567);
nand U2849 (N_2849,N_2404,N_2474);
xnor U2850 (N_2850,N_2413,N_2641);
xor U2851 (N_2851,N_2468,N_2521);
or U2852 (N_2852,N_2651,N_2452);
nand U2853 (N_2853,N_2698,N_2671);
and U2854 (N_2854,N_2447,N_2589);
xnor U2855 (N_2855,N_2603,N_2408);
nor U2856 (N_2856,N_2547,N_2488);
nand U2857 (N_2857,N_2599,N_2506);
and U2858 (N_2858,N_2591,N_2636);
and U2859 (N_2859,N_2418,N_2569);
nand U2860 (N_2860,N_2427,N_2691);
or U2861 (N_2861,N_2504,N_2687);
and U2862 (N_2862,N_2430,N_2520);
xor U2863 (N_2863,N_2655,N_2490);
and U2864 (N_2864,N_2598,N_2484);
or U2865 (N_2865,N_2661,N_2563);
nor U2866 (N_2866,N_2595,N_2481);
nor U2867 (N_2867,N_2442,N_2473);
or U2868 (N_2868,N_2584,N_2571);
or U2869 (N_2869,N_2549,N_2424);
or U2870 (N_2870,N_2466,N_2409);
nor U2871 (N_2871,N_2560,N_2539);
xor U2872 (N_2872,N_2566,N_2590);
nand U2873 (N_2873,N_2435,N_2646);
and U2874 (N_2874,N_2576,N_2445);
nor U2875 (N_2875,N_2509,N_2674);
xnor U2876 (N_2876,N_2559,N_2523);
nand U2877 (N_2877,N_2503,N_2626);
nor U2878 (N_2878,N_2613,N_2654);
nand U2879 (N_2879,N_2488,N_2586);
and U2880 (N_2880,N_2459,N_2580);
or U2881 (N_2881,N_2469,N_2642);
and U2882 (N_2882,N_2507,N_2411);
nand U2883 (N_2883,N_2595,N_2564);
nor U2884 (N_2884,N_2428,N_2649);
nor U2885 (N_2885,N_2629,N_2580);
xnor U2886 (N_2886,N_2491,N_2638);
and U2887 (N_2887,N_2401,N_2573);
xnor U2888 (N_2888,N_2631,N_2534);
and U2889 (N_2889,N_2684,N_2514);
nor U2890 (N_2890,N_2527,N_2517);
or U2891 (N_2891,N_2636,N_2629);
nand U2892 (N_2892,N_2445,N_2459);
or U2893 (N_2893,N_2471,N_2654);
nand U2894 (N_2894,N_2443,N_2572);
and U2895 (N_2895,N_2590,N_2668);
or U2896 (N_2896,N_2655,N_2424);
xor U2897 (N_2897,N_2474,N_2553);
and U2898 (N_2898,N_2465,N_2426);
or U2899 (N_2899,N_2656,N_2602);
or U2900 (N_2900,N_2494,N_2576);
or U2901 (N_2901,N_2411,N_2521);
or U2902 (N_2902,N_2465,N_2556);
and U2903 (N_2903,N_2490,N_2560);
nor U2904 (N_2904,N_2432,N_2607);
nand U2905 (N_2905,N_2653,N_2598);
nand U2906 (N_2906,N_2637,N_2404);
or U2907 (N_2907,N_2544,N_2573);
nand U2908 (N_2908,N_2659,N_2569);
and U2909 (N_2909,N_2566,N_2447);
nor U2910 (N_2910,N_2515,N_2512);
or U2911 (N_2911,N_2558,N_2627);
nand U2912 (N_2912,N_2562,N_2686);
and U2913 (N_2913,N_2499,N_2404);
nor U2914 (N_2914,N_2569,N_2681);
nor U2915 (N_2915,N_2643,N_2656);
xor U2916 (N_2916,N_2412,N_2517);
nand U2917 (N_2917,N_2655,N_2640);
nand U2918 (N_2918,N_2657,N_2467);
nor U2919 (N_2919,N_2477,N_2419);
or U2920 (N_2920,N_2650,N_2590);
nor U2921 (N_2921,N_2412,N_2636);
and U2922 (N_2922,N_2484,N_2629);
nand U2923 (N_2923,N_2545,N_2403);
and U2924 (N_2924,N_2645,N_2579);
xnor U2925 (N_2925,N_2435,N_2548);
and U2926 (N_2926,N_2629,N_2430);
nor U2927 (N_2927,N_2620,N_2626);
or U2928 (N_2928,N_2573,N_2528);
or U2929 (N_2929,N_2687,N_2635);
xor U2930 (N_2930,N_2473,N_2692);
and U2931 (N_2931,N_2570,N_2523);
and U2932 (N_2932,N_2590,N_2649);
nor U2933 (N_2933,N_2403,N_2599);
or U2934 (N_2934,N_2495,N_2587);
nand U2935 (N_2935,N_2496,N_2612);
xnor U2936 (N_2936,N_2681,N_2669);
xor U2937 (N_2937,N_2449,N_2600);
nor U2938 (N_2938,N_2558,N_2654);
and U2939 (N_2939,N_2605,N_2516);
nand U2940 (N_2940,N_2491,N_2604);
xnor U2941 (N_2941,N_2662,N_2479);
xnor U2942 (N_2942,N_2652,N_2499);
xnor U2943 (N_2943,N_2439,N_2500);
and U2944 (N_2944,N_2672,N_2683);
nand U2945 (N_2945,N_2408,N_2539);
nor U2946 (N_2946,N_2521,N_2605);
xor U2947 (N_2947,N_2454,N_2598);
or U2948 (N_2948,N_2686,N_2650);
nand U2949 (N_2949,N_2536,N_2453);
or U2950 (N_2950,N_2473,N_2593);
or U2951 (N_2951,N_2408,N_2502);
xor U2952 (N_2952,N_2513,N_2481);
nand U2953 (N_2953,N_2406,N_2553);
xnor U2954 (N_2954,N_2678,N_2582);
nor U2955 (N_2955,N_2610,N_2517);
xnor U2956 (N_2956,N_2604,N_2685);
and U2957 (N_2957,N_2686,N_2475);
nor U2958 (N_2958,N_2469,N_2638);
nor U2959 (N_2959,N_2675,N_2457);
nor U2960 (N_2960,N_2435,N_2672);
or U2961 (N_2961,N_2454,N_2536);
nand U2962 (N_2962,N_2512,N_2521);
nand U2963 (N_2963,N_2508,N_2486);
or U2964 (N_2964,N_2581,N_2417);
and U2965 (N_2965,N_2485,N_2607);
or U2966 (N_2966,N_2412,N_2585);
nand U2967 (N_2967,N_2600,N_2553);
xnor U2968 (N_2968,N_2525,N_2555);
xor U2969 (N_2969,N_2483,N_2435);
nand U2970 (N_2970,N_2471,N_2465);
or U2971 (N_2971,N_2594,N_2572);
and U2972 (N_2972,N_2431,N_2642);
nand U2973 (N_2973,N_2598,N_2657);
nor U2974 (N_2974,N_2452,N_2417);
nand U2975 (N_2975,N_2588,N_2577);
or U2976 (N_2976,N_2438,N_2499);
xor U2977 (N_2977,N_2516,N_2647);
and U2978 (N_2978,N_2662,N_2604);
nand U2979 (N_2979,N_2485,N_2477);
nand U2980 (N_2980,N_2491,N_2522);
and U2981 (N_2981,N_2405,N_2611);
and U2982 (N_2982,N_2476,N_2582);
xor U2983 (N_2983,N_2534,N_2402);
or U2984 (N_2984,N_2402,N_2422);
nand U2985 (N_2985,N_2691,N_2629);
and U2986 (N_2986,N_2429,N_2621);
and U2987 (N_2987,N_2634,N_2507);
and U2988 (N_2988,N_2449,N_2614);
xor U2989 (N_2989,N_2642,N_2453);
nand U2990 (N_2990,N_2605,N_2561);
and U2991 (N_2991,N_2623,N_2665);
or U2992 (N_2992,N_2681,N_2496);
xor U2993 (N_2993,N_2493,N_2678);
and U2994 (N_2994,N_2699,N_2589);
nand U2995 (N_2995,N_2461,N_2411);
and U2996 (N_2996,N_2669,N_2582);
and U2997 (N_2997,N_2533,N_2480);
nand U2998 (N_2998,N_2411,N_2638);
xor U2999 (N_2999,N_2459,N_2629);
nor U3000 (N_3000,N_2911,N_2701);
nor U3001 (N_3001,N_2762,N_2920);
nand U3002 (N_3002,N_2879,N_2909);
xnor U3003 (N_3003,N_2792,N_2732);
nor U3004 (N_3004,N_2825,N_2872);
nand U3005 (N_3005,N_2827,N_2771);
xnor U3006 (N_3006,N_2831,N_2845);
xnor U3007 (N_3007,N_2788,N_2858);
or U3008 (N_3008,N_2961,N_2812);
and U3009 (N_3009,N_2778,N_2970);
nor U3010 (N_3010,N_2804,N_2744);
nor U3011 (N_3011,N_2999,N_2848);
nor U3012 (N_3012,N_2718,N_2763);
and U3013 (N_3013,N_2774,N_2757);
and U3014 (N_3014,N_2838,N_2839);
nor U3015 (N_3015,N_2975,N_2952);
nor U3016 (N_3016,N_2834,N_2708);
xor U3017 (N_3017,N_2795,N_2726);
and U3018 (N_3018,N_2981,N_2809);
or U3019 (N_3019,N_2945,N_2853);
nand U3020 (N_3020,N_2985,N_2968);
xor U3021 (N_3021,N_2821,N_2967);
nor U3022 (N_3022,N_2724,N_2764);
nor U3023 (N_3023,N_2918,N_2852);
and U3024 (N_3024,N_2950,N_2972);
nand U3025 (N_3025,N_2880,N_2815);
nand U3026 (N_3026,N_2801,N_2913);
nor U3027 (N_3027,N_2704,N_2807);
nand U3028 (N_3028,N_2990,N_2980);
xnor U3029 (N_3029,N_2811,N_2751);
or U3030 (N_3030,N_2867,N_2816);
and U3031 (N_3031,N_2758,N_2703);
nand U3032 (N_3032,N_2733,N_2769);
and U3033 (N_3033,N_2844,N_2766);
nor U3034 (N_3034,N_2829,N_2900);
xnor U3035 (N_3035,N_2754,N_2836);
and U3036 (N_3036,N_2780,N_2817);
xor U3037 (N_3037,N_2926,N_2921);
xnor U3038 (N_3038,N_2898,N_2856);
nand U3039 (N_3039,N_2842,N_2720);
xnor U3040 (N_3040,N_2794,N_2702);
or U3041 (N_3041,N_2716,N_2884);
or U3042 (N_3042,N_2934,N_2917);
xnor U3043 (N_3043,N_2925,N_2896);
nand U3044 (N_3044,N_2940,N_2745);
or U3045 (N_3045,N_2765,N_2988);
or U3046 (N_3046,N_2965,N_2916);
or U3047 (N_3047,N_2748,N_2837);
xnor U3048 (N_3048,N_2791,N_2722);
and U3049 (N_3049,N_2796,N_2908);
nor U3050 (N_3050,N_2959,N_2723);
and U3051 (N_3051,N_2759,N_2728);
xnor U3052 (N_3052,N_2750,N_2814);
nor U3053 (N_3053,N_2717,N_2753);
xor U3054 (N_3054,N_2901,N_2871);
nor U3055 (N_3055,N_2855,N_2730);
xnor U3056 (N_3056,N_2863,N_2893);
nor U3057 (N_3057,N_2889,N_2971);
xor U3058 (N_3058,N_2773,N_2857);
xor U3059 (N_3059,N_2713,N_2885);
nand U3060 (N_3060,N_2962,N_2808);
nand U3061 (N_3061,N_2946,N_2873);
nand U3062 (N_3062,N_2897,N_2775);
nand U3063 (N_3063,N_2851,N_2731);
or U3064 (N_3064,N_2986,N_2859);
nand U3065 (N_3065,N_2923,N_2734);
and U3066 (N_3066,N_2951,N_2709);
nand U3067 (N_3067,N_2998,N_2976);
nand U3068 (N_3068,N_2974,N_2942);
xor U3069 (N_3069,N_2785,N_2877);
and U3070 (N_3070,N_2707,N_2932);
and U3071 (N_3071,N_2712,N_2761);
nand U3072 (N_3072,N_2818,N_2833);
or U3073 (N_3073,N_2823,N_2865);
and U3074 (N_3074,N_2755,N_2953);
xor U3075 (N_3075,N_2957,N_2841);
or U3076 (N_3076,N_2881,N_2910);
nor U3077 (N_3077,N_2735,N_2711);
nor U3078 (N_3078,N_2914,N_2805);
or U3079 (N_3079,N_2832,N_2887);
nor U3080 (N_3080,N_2924,N_2937);
or U3081 (N_3081,N_2861,N_2847);
xor U3082 (N_3082,N_2776,N_2800);
nand U3083 (N_3083,N_2928,N_2943);
nor U3084 (N_3084,N_2907,N_2992);
nor U3085 (N_3085,N_2882,N_2875);
and U3086 (N_3086,N_2870,N_2983);
and U3087 (N_3087,N_2888,N_2790);
or U3088 (N_3088,N_2982,N_2949);
nand U3089 (N_3089,N_2860,N_2736);
or U3090 (N_3090,N_2715,N_2803);
xnor U3091 (N_3091,N_2903,N_2770);
and U3092 (N_3092,N_2954,N_2938);
nand U3093 (N_3093,N_2710,N_2714);
xor U3094 (N_3094,N_2793,N_2995);
nand U3095 (N_3095,N_2919,N_2895);
or U3096 (N_3096,N_2705,N_2768);
nor U3097 (N_3097,N_2850,N_2905);
xnor U3098 (N_3098,N_2966,N_2749);
and U3099 (N_3099,N_2941,N_2820);
nand U3100 (N_3100,N_2944,N_2787);
and U3101 (N_3101,N_2984,N_2782);
nand U3102 (N_3102,N_2789,N_2779);
nand U3103 (N_3103,N_2930,N_2947);
xor U3104 (N_3104,N_2799,N_2862);
or U3105 (N_3105,N_2936,N_2892);
nand U3106 (N_3106,N_2840,N_2874);
or U3107 (N_3107,N_2741,N_2899);
or U3108 (N_3108,N_2725,N_2784);
nand U3109 (N_3109,N_2835,N_2721);
or U3110 (N_3110,N_2849,N_2977);
xnor U3111 (N_3111,N_2786,N_2996);
and U3112 (N_3112,N_2846,N_2978);
nor U3113 (N_3113,N_2963,N_2989);
xnor U3114 (N_3114,N_2854,N_2760);
or U3115 (N_3115,N_2706,N_2729);
and U3116 (N_3116,N_2739,N_2819);
nor U3117 (N_3117,N_2783,N_2866);
and U3118 (N_3118,N_2743,N_2902);
and U3119 (N_3119,N_2746,N_2931);
nor U3120 (N_3120,N_2813,N_2890);
nand U3121 (N_3121,N_2935,N_2752);
nor U3122 (N_3122,N_2929,N_2894);
and U3123 (N_3123,N_2876,N_2738);
or U3124 (N_3124,N_2891,N_2843);
nand U3125 (N_3125,N_2830,N_2939);
and U3126 (N_3126,N_2737,N_2824);
xnor U3127 (N_3127,N_2915,N_2991);
xnor U3128 (N_3128,N_2868,N_2927);
and U3129 (N_3129,N_2987,N_2906);
nand U3130 (N_3130,N_2727,N_2781);
or U3131 (N_3131,N_2955,N_2802);
or U3132 (N_3132,N_2973,N_2883);
nand U3133 (N_3133,N_2869,N_2740);
nor U3134 (N_3134,N_2797,N_2767);
or U3135 (N_3135,N_2912,N_2798);
nand U3136 (N_3136,N_2922,N_2826);
and U3137 (N_3137,N_2933,N_2960);
and U3138 (N_3138,N_2878,N_2956);
nor U3139 (N_3139,N_2904,N_2828);
xor U3140 (N_3140,N_2964,N_2864);
nor U3141 (N_3141,N_2979,N_2969);
nor U3142 (N_3142,N_2756,N_2997);
or U3143 (N_3143,N_2948,N_2958);
nor U3144 (N_3144,N_2777,N_2719);
and U3145 (N_3145,N_2742,N_2772);
nor U3146 (N_3146,N_2886,N_2747);
xnor U3147 (N_3147,N_2810,N_2994);
or U3148 (N_3148,N_2993,N_2700);
nand U3149 (N_3149,N_2806,N_2822);
or U3150 (N_3150,N_2992,N_2886);
nor U3151 (N_3151,N_2862,N_2969);
xnor U3152 (N_3152,N_2800,N_2782);
nor U3153 (N_3153,N_2808,N_2830);
and U3154 (N_3154,N_2746,N_2952);
nand U3155 (N_3155,N_2801,N_2713);
nand U3156 (N_3156,N_2703,N_2901);
nor U3157 (N_3157,N_2973,N_2863);
nor U3158 (N_3158,N_2861,N_2888);
nor U3159 (N_3159,N_2784,N_2961);
nand U3160 (N_3160,N_2847,N_2904);
nand U3161 (N_3161,N_2842,N_2950);
nor U3162 (N_3162,N_2885,N_2760);
or U3163 (N_3163,N_2965,N_2810);
and U3164 (N_3164,N_2803,N_2780);
xor U3165 (N_3165,N_2756,N_2911);
xor U3166 (N_3166,N_2732,N_2935);
xnor U3167 (N_3167,N_2994,N_2905);
or U3168 (N_3168,N_2858,N_2900);
or U3169 (N_3169,N_2778,N_2795);
nand U3170 (N_3170,N_2732,N_2793);
and U3171 (N_3171,N_2780,N_2938);
or U3172 (N_3172,N_2906,N_2999);
nand U3173 (N_3173,N_2827,N_2912);
nor U3174 (N_3174,N_2926,N_2905);
nand U3175 (N_3175,N_2743,N_2832);
nand U3176 (N_3176,N_2947,N_2802);
and U3177 (N_3177,N_2950,N_2884);
nor U3178 (N_3178,N_2954,N_2842);
and U3179 (N_3179,N_2866,N_2772);
and U3180 (N_3180,N_2782,N_2767);
and U3181 (N_3181,N_2820,N_2895);
nand U3182 (N_3182,N_2921,N_2875);
or U3183 (N_3183,N_2956,N_2725);
nand U3184 (N_3184,N_2832,N_2898);
nand U3185 (N_3185,N_2824,N_2830);
xnor U3186 (N_3186,N_2731,N_2822);
nor U3187 (N_3187,N_2789,N_2711);
or U3188 (N_3188,N_2716,N_2920);
xnor U3189 (N_3189,N_2808,N_2921);
xnor U3190 (N_3190,N_2714,N_2850);
and U3191 (N_3191,N_2817,N_2827);
nand U3192 (N_3192,N_2998,N_2748);
nor U3193 (N_3193,N_2868,N_2836);
nor U3194 (N_3194,N_2705,N_2796);
xnor U3195 (N_3195,N_2742,N_2785);
and U3196 (N_3196,N_2723,N_2777);
nand U3197 (N_3197,N_2733,N_2779);
and U3198 (N_3198,N_2721,N_2863);
nor U3199 (N_3199,N_2999,N_2948);
xor U3200 (N_3200,N_2872,N_2729);
nand U3201 (N_3201,N_2973,N_2920);
xor U3202 (N_3202,N_2745,N_2944);
xor U3203 (N_3203,N_2743,N_2834);
or U3204 (N_3204,N_2742,N_2751);
and U3205 (N_3205,N_2860,N_2927);
xor U3206 (N_3206,N_2954,N_2963);
and U3207 (N_3207,N_2835,N_2985);
xor U3208 (N_3208,N_2846,N_2827);
and U3209 (N_3209,N_2862,N_2998);
nor U3210 (N_3210,N_2780,N_2869);
nor U3211 (N_3211,N_2942,N_2896);
nand U3212 (N_3212,N_2837,N_2880);
or U3213 (N_3213,N_2768,N_2813);
and U3214 (N_3214,N_2799,N_2778);
and U3215 (N_3215,N_2915,N_2734);
or U3216 (N_3216,N_2924,N_2750);
and U3217 (N_3217,N_2743,N_2772);
nor U3218 (N_3218,N_2791,N_2777);
xor U3219 (N_3219,N_2957,N_2798);
or U3220 (N_3220,N_2921,N_2856);
xnor U3221 (N_3221,N_2917,N_2707);
xor U3222 (N_3222,N_2843,N_2860);
nand U3223 (N_3223,N_2754,N_2909);
nand U3224 (N_3224,N_2892,N_2799);
or U3225 (N_3225,N_2870,N_2923);
nand U3226 (N_3226,N_2815,N_2883);
and U3227 (N_3227,N_2823,N_2798);
nor U3228 (N_3228,N_2857,N_2710);
nor U3229 (N_3229,N_2930,N_2835);
nor U3230 (N_3230,N_2746,N_2758);
or U3231 (N_3231,N_2707,N_2978);
xor U3232 (N_3232,N_2817,N_2788);
or U3233 (N_3233,N_2802,N_2959);
nand U3234 (N_3234,N_2867,N_2719);
nor U3235 (N_3235,N_2742,N_2748);
nand U3236 (N_3236,N_2898,N_2719);
and U3237 (N_3237,N_2918,N_2767);
and U3238 (N_3238,N_2851,N_2970);
and U3239 (N_3239,N_2881,N_2899);
xnor U3240 (N_3240,N_2969,N_2715);
xor U3241 (N_3241,N_2750,N_2974);
nand U3242 (N_3242,N_2916,N_2733);
nand U3243 (N_3243,N_2806,N_2923);
nor U3244 (N_3244,N_2936,N_2768);
xor U3245 (N_3245,N_2754,N_2720);
or U3246 (N_3246,N_2776,N_2866);
nand U3247 (N_3247,N_2965,N_2797);
xor U3248 (N_3248,N_2863,N_2952);
xor U3249 (N_3249,N_2787,N_2838);
nand U3250 (N_3250,N_2956,N_2909);
nor U3251 (N_3251,N_2827,N_2742);
xor U3252 (N_3252,N_2793,N_2974);
xnor U3253 (N_3253,N_2835,N_2879);
xnor U3254 (N_3254,N_2899,N_2986);
nand U3255 (N_3255,N_2936,N_2715);
nand U3256 (N_3256,N_2765,N_2895);
xor U3257 (N_3257,N_2959,N_2773);
nor U3258 (N_3258,N_2976,N_2721);
and U3259 (N_3259,N_2877,N_2727);
and U3260 (N_3260,N_2784,N_2886);
or U3261 (N_3261,N_2877,N_2973);
or U3262 (N_3262,N_2931,N_2754);
and U3263 (N_3263,N_2871,N_2940);
nand U3264 (N_3264,N_2990,N_2777);
nor U3265 (N_3265,N_2725,N_2992);
xnor U3266 (N_3266,N_2745,N_2885);
nand U3267 (N_3267,N_2741,N_2786);
and U3268 (N_3268,N_2922,N_2770);
or U3269 (N_3269,N_2778,N_2803);
and U3270 (N_3270,N_2793,N_2936);
xor U3271 (N_3271,N_2786,N_2888);
nor U3272 (N_3272,N_2851,N_2930);
nor U3273 (N_3273,N_2839,N_2949);
and U3274 (N_3274,N_2748,N_2752);
or U3275 (N_3275,N_2938,N_2877);
or U3276 (N_3276,N_2901,N_2916);
or U3277 (N_3277,N_2927,N_2912);
or U3278 (N_3278,N_2933,N_2964);
or U3279 (N_3279,N_2827,N_2718);
xor U3280 (N_3280,N_2881,N_2901);
xor U3281 (N_3281,N_2844,N_2746);
xor U3282 (N_3282,N_2976,N_2749);
and U3283 (N_3283,N_2888,N_2935);
nor U3284 (N_3284,N_2790,N_2798);
xnor U3285 (N_3285,N_2968,N_2835);
nor U3286 (N_3286,N_2927,N_2782);
xor U3287 (N_3287,N_2766,N_2999);
nor U3288 (N_3288,N_2969,N_2789);
nand U3289 (N_3289,N_2793,N_2780);
nor U3290 (N_3290,N_2825,N_2973);
and U3291 (N_3291,N_2707,N_2923);
and U3292 (N_3292,N_2778,N_2704);
nand U3293 (N_3293,N_2860,N_2986);
or U3294 (N_3294,N_2778,N_2857);
xnor U3295 (N_3295,N_2732,N_2959);
nand U3296 (N_3296,N_2837,N_2791);
or U3297 (N_3297,N_2979,N_2915);
and U3298 (N_3298,N_2705,N_2823);
nand U3299 (N_3299,N_2995,N_2965);
nor U3300 (N_3300,N_3010,N_3159);
or U3301 (N_3301,N_3103,N_3160);
or U3302 (N_3302,N_3209,N_3178);
and U3303 (N_3303,N_3157,N_3239);
xnor U3304 (N_3304,N_3024,N_3051);
or U3305 (N_3305,N_3088,N_3138);
nand U3306 (N_3306,N_3074,N_3216);
nand U3307 (N_3307,N_3210,N_3141);
xnor U3308 (N_3308,N_3270,N_3077);
and U3309 (N_3309,N_3208,N_3238);
nor U3310 (N_3310,N_3104,N_3096);
nand U3311 (N_3311,N_3277,N_3030);
nor U3312 (N_3312,N_3025,N_3260);
xnor U3313 (N_3313,N_3266,N_3023);
nand U3314 (N_3314,N_3139,N_3150);
nand U3315 (N_3315,N_3041,N_3008);
and U3316 (N_3316,N_3113,N_3232);
or U3317 (N_3317,N_3129,N_3043);
nor U3318 (N_3318,N_3197,N_3133);
nand U3319 (N_3319,N_3134,N_3251);
nand U3320 (N_3320,N_3081,N_3156);
nand U3321 (N_3321,N_3070,N_3082);
xnor U3322 (N_3322,N_3241,N_3117);
nor U3323 (N_3323,N_3244,N_3126);
and U3324 (N_3324,N_3035,N_3203);
xnor U3325 (N_3325,N_3089,N_3225);
and U3326 (N_3326,N_3233,N_3111);
nand U3327 (N_3327,N_3254,N_3064);
nand U3328 (N_3328,N_3108,N_3021);
nor U3329 (N_3329,N_3227,N_3243);
and U3330 (N_3330,N_3095,N_3048);
nor U3331 (N_3331,N_3196,N_3223);
nor U3332 (N_3332,N_3242,N_3173);
or U3333 (N_3333,N_3221,N_3107);
xor U3334 (N_3334,N_3115,N_3128);
nand U3335 (N_3335,N_3200,N_3015);
and U3336 (N_3336,N_3259,N_3031);
nand U3337 (N_3337,N_3154,N_3132);
xnor U3338 (N_3338,N_3290,N_3056);
nor U3339 (N_3339,N_3253,N_3009);
nor U3340 (N_3340,N_3072,N_3174);
nand U3341 (N_3341,N_3172,N_3136);
or U3342 (N_3342,N_3257,N_3166);
nor U3343 (N_3343,N_3131,N_3091);
and U3344 (N_3344,N_3247,N_3013);
nand U3345 (N_3345,N_3191,N_3292);
nand U3346 (N_3346,N_3050,N_3019);
and U3347 (N_3347,N_3042,N_3094);
nand U3348 (N_3348,N_3265,N_3256);
nor U3349 (N_3349,N_3175,N_3155);
nand U3350 (N_3350,N_3145,N_3246);
or U3351 (N_3351,N_3059,N_3269);
and U3352 (N_3352,N_3252,N_3002);
nor U3353 (N_3353,N_3230,N_3228);
or U3354 (N_3354,N_3073,N_3274);
nand U3355 (N_3355,N_3123,N_3075);
or U3356 (N_3356,N_3083,N_3135);
xor U3357 (N_3357,N_3118,N_3293);
and U3358 (N_3358,N_3076,N_3218);
nand U3359 (N_3359,N_3183,N_3020);
and U3360 (N_3360,N_3007,N_3215);
xnor U3361 (N_3361,N_3214,N_3177);
or U3362 (N_3362,N_3106,N_3049);
xor U3363 (N_3363,N_3090,N_3144);
nand U3364 (N_3364,N_3057,N_3032);
or U3365 (N_3365,N_3061,N_3190);
xor U3366 (N_3366,N_3109,N_3003);
and U3367 (N_3367,N_3034,N_3182);
nor U3368 (N_3368,N_3261,N_3080);
and U3369 (N_3369,N_3058,N_3069);
nor U3370 (N_3370,N_3062,N_3119);
or U3371 (N_3371,N_3116,N_3276);
or U3372 (N_3372,N_3192,N_3294);
or U3373 (N_3373,N_3263,N_3086);
xor U3374 (N_3374,N_3204,N_3201);
nor U3375 (N_3375,N_3189,N_3176);
or U3376 (N_3376,N_3185,N_3017);
and U3377 (N_3377,N_3219,N_3028);
xnor U3378 (N_3378,N_3255,N_3044);
nor U3379 (N_3379,N_3250,N_3000);
and U3380 (N_3380,N_3281,N_3211);
nor U3381 (N_3381,N_3130,N_3291);
nor U3382 (N_3382,N_3212,N_3120);
and U3383 (N_3383,N_3143,N_3102);
and U3384 (N_3384,N_3137,N_3188);
and U3385 (N_3385,N_3224,N_3187);
nor U3386 (N_3386,N_3078,N_3039);
or U3387 (N_3387,N_3264,N_3026);
or U3388 (N_3388,N_3280,N_3165);
nand U3389 (N_3389,N_3205,N_3275);
nor U3390 (N_3390,N_3033,N_3297);
and U3391 (N_3391,N_3038,N_3198);
nand U3392 (N_3392,N_3164,N_3146);
xnor U3393 (N_3393,N_3283,N_3278);
nand U3394 (N_3394,N_3001,N_3055);
nor U3395 (N_3395,N_3231,N_3045);
and U3396 (N_3396,N_3016,N_3258);
or U3397 (N_3397,N_3124,N_3193);
xnor U3398 (N_3398,N_3063,N_3097);
nor U3399 (N_3399,N_3289,N_3229);
nand U3400 (N_3400,N_3287,N_3158);
xor U3401 (N_3401,N_3112,N_3195);
or U3402 (N_3402,N_3068,N_3127);
and U3403 (N_3403,N_3060,N_3153);
xnor U3404 (N_3404,N_3110,N_3161);
and U3405 (N_3405,N_3168,N_3036);
nand U3406 (N_3406,N_3163,N_3027);
nor U3407 (N_3407,N_3011,N_3226);
or U3408 (N_3408,N_3236,N_3149);
nand U3409 (N_3409,N_3046,N_3213);
and U3410 (N_3410,N_3207,N_3140);
nor U3411 (N_3411,N_3029,N_3184);
nor U3412 (N_3412,N_3288,N_3100);
nand U3413 (N_3413,N_3206,N_3054);
nor U3414 (N_3414,N_3147,N_3114);
and U3415 (N_3415,N_3098,N_3181);
nand U3416 (N_3416,N_3179,N_3167);
nand U3417 (N_3417,N_3240,N_3012);
and U3418 (N_3418,N_3199,N_3125);
and U3419 (N_3419,N_3194,N_3245);
nand U3420 (N_3420,N_3171,N_3202);
and U3421 (N_3421,N_3065,N_3105);
nand U3422 (N_3422,N_3282,N_3170);
xnor U3423 (N_3423,N_3284,N_3249);
nand U3424 (N_3424,N_3222,N_3272);
and U3425 (N_3425,N_3066,N_3295);
or U3426 (N_3426,N_3052,N_3004);
or U3427 (N_3427,N_3273,N_3180);
nand U3428 (N_3428,N_3006,N_3296);
and U3429 (N_3429,N_3084,N_3248);
and U3430 (N_3430,N_3018,N_3014);
nor U3431 (N_3431,N_3101,N_3298);
nor U3432 (N_3432,N_3186,N_3142);
or U3433 (N_3433,N_3148,N_3286);
nand U3434 (N_3434,N_3152,N_3162);
nor U3435 (N_3435,N_3079,N_3093);
nor U3436 (N_3436,N_3087,N_3037);
nand U3437 (N_3437,N_3279,N_3262);
or U3438 (N_3438,N_3047,N_3005);
nor U3439 (N_3439,N_3217,N_3040);
xor U3440 (N_3440,N_3085,N_3237);
xnor U3441 (N_3441,N_3022,N_3121);
or U3442 (N_3442,N_3267,N_3122);
or U3443 (N_3443,N_3285,N_3235);
nor U3444 (N_3444,N_3067,N_3268);
or U3445 (N_3445,N_3099,N_3092);
nor U3446 (N_3446,N_3220,N_3053);
nand U3447 (N_3447,N_3234,N_3299);
or U3448 (N_3448,N_3271,N_3151);
xnor U3449 (N_3449,N_3071,N_3169);
and U3450 (N_3450,N_3117,N_3173);
xnor U3451 (N_3451,N_3012,N_3130);
and U3452 (N_3452,N_3227,N_3240);
or U3453 (N_3453,N_3255,N_3290);
or U3454 (N_3454,N_3287,N_3133);
nand U3455 (N_3455,N_3190,N_3090);
and U3456 (N_3456,N_3089,N_3203);
nand U3457 (N_3457,N_3267,N_3139);
or U3458 (N_3458,N_3154,N_3212);
nor U3459 (N_3459,N_3039,N_3252);
nor U3460 (N_3460,N_3157,N_3205);
nor U3461 (N_3461,N_3016,N_3218);
xor U3462 (N_3462,N_3084,N_3028);
or U3463 (N_3463,N_3107,N_3161);
nor U3464 (N_3464,N_3128,N_3223);
or U3465 (N_3465,N_3026,N_3200);
or U3466 (N_3466,N_3072,N_3018);
or U3467 (N_3467,N_3037,N_3191);
and U3468 (N_3468,N_3125,N_3026);
xnor U3469 (N_3469,N_3183,N_3060);
or U3470 (N_3470,N_3209,N_3220);
xnor U3471 (N_3471,N_3217,N_3152);
and U3472 (N_3472,N_3127,N_3158);
xor U3473 (N_3473,N_3185,N_3088);
nor U3474 (N_3474,N_3242,N_3227);
and U3475 (N_3475,N_3065,N_3195);
and U3476 (N_3476,N_3043,N_3088);
or U3477 (N_3477,N_3128,N_3229);
nor U3478 (N_3478,N_3153,N_3141);
and U3479 (N_3479,N_3082,N_3244);
or U3480 (N_3480,N_3167,N_3042);
nand U3481 (N_3481,N_3252,N_3016);
and U3482 (N_3482,N_3239,N_3184);
xnor U3483 (N_3483,N_3279,N_3039);
or U3484 (N_3484,N_3071,N_3111);
nand U3485 (N_3485,N_3209,N_3238);
xnor U3486 (N_3486,N_3148,N_3130);
or U3487 (N_3487,N_3053,N_3128);
xnor U3488 (N_3488,N_3235,N_3241);
nor U3489 (N_3489,N_3114,N_3083);
nand U3490 (N_3490,N_3229,N_3217);
and U3491 (N_3491,N_3152,N_3044);
and U3492 (N_3492,N_3264,N_3189);
nor U3493 (N_3493,N_3058,N_3003);
xnor U3494 (N_3494,N_3066,N_3145);
and U3495 (N_3495,N_3208,N_3252);
or U3496 (N_3496,N_3201,N_3156);
or U3497 (N_3497,N_3149,N_3259);
xnor U3498 (N_3498,N_3143,N_3089);
nand U3499 (N_3499,N_3215,N_3157);
xor U3500 (N_3500,N_3114,N_3120);
nand U3501 (N_3501,N_3047,N_3009);
or U3502 (N_3502,N_3014,N_3159);
nand U3503 (N_3503,N_3008,N_3240);
or U3504 (N_3504,N_3090,N_3243);
or U3505 (N_3505,N_3103,N_3029);
xor U3506 (N_3506,N_3213,N_3018);
xor U3507 (N_3507,N_3131,N_3272);
nand U3508 (N_3508,N_3291,N_3231);
xor U3509 (N_3509,N_3052,N_3109);
nand U3510 (N_3510,N_3220,N_3195);
and U3511 (N_3511,N_3207,N_3049);
nand U3512 (N_3512,N_3138,N_3218);
nor U3513 (N_3513,N_3251,N_3136);
nand U3514 (N_3514,N_3150,N_3202);
and U3515 (N_3515,N_3166,N_3124);
nand U3516 (N_3516,N_3227,N_3027);
or U3517 (N_3517,N_3098,N_3216);
nand U3518 (N_3518,N_3190,N_3059);
and U3519 (N_3519,N_3166,N_3079);
or U3520 (N_3520,N_3247,N_3175);
and U3521 (N_3521,N_3294,N_3060);
nor U3522 (N_3522,N_3202,N_3291);
xnor U3523 (N_3523,N_3257,N_3049);
nand U3524 (N_3524,N_3213,N_3028);
and U3525 (N_3525,N_3240,N_3254);
xnor U3526 (N_3526,N_3078,N_3164);
nor U3527 (N_3527,N_3137,N_3294);
or U3528 (N_3528,N_3295,N_3017);
xor U3529 (N_3529,N_3031,N_3282);
nand U3530 (N_3530,N_3283,N_3295);
xor U3531 (N_3531,N_3119,N_3149);
nand U3532 (N_3532,N_3206,N_3063);
nand U3533 (N_3533,N_3186,N_3243);
and U3534 (N_3534,N_3153,N_3053);
nor U3535 (N_3535,N_3257,N_3092);
nand U3536 (N_3536,N_3080,N_3128);
nor U3537 (N_3537,N_3218,N_3288);
nor U3538 (N_3538,N_3047,N_3223);
nand U3539 (N_3539,N_3040,N_3253);
and U3540 (N_3540,N_3050,N_3190);
xor U3541 (N_3541,N_3011,N_3151);
xnor U3542 (N_3542,N_3264,N_3127);
or U3543 (N_3543,N_3246,N_3281);
and U3544 (N_3544,N_3077,N_3035);
xnor U3545 (N_3545,N_3181,N_3157);
and U3546 (N_3546,N_3266,N_3117);
nor U3547 (N_3547,N_3113,N_3195);
xor U3548 (N_3548,N_3167,N_3100);
nand U3549 (N_3549,N_3220,N_3130);
xor U3550 (N_3550,N_3003,N_3051);
and U3551 (N_3551,N_3096,N_3041);
and U3552 (N_3552,N_3271,N_3231);
or U3553 (N_3553,N_3281,N_3212);
nor U3554 (N_3554,N_3289,N_3297);
nand U3555 (N_3555,N_3083,N_3163);
or U3556 (N_3556,N_3243,N_3209);
nor U3557 (N_3557,N_3269,N_3285);
xnor U3558 (N_3558,N_3250,N_3152);
nor U3559 (N_3559,N_3039,N_3272);
xnor U3560 (N_3560,N_3077,N_3096);
nand U3561 (N_3561,N_3023,N_3028);
nor U3562 (N_3562,N_3264,N_3247);
xnor U3563 (N_3563,N_3297,N_3240);
and U3564 (N_3564,N_3196,N_3148);
xor U3565 (N_3565,N_3130,N_3098);
nor U3566 (N_3566,N_3247,N_3062);
and U3567 (N_3567,N_3050,N_3254);
nor U3568 (N_3568,N_3030,N_3214);
nor U3569 (N_3569,N_3299,N_3153);
and U3570 (N_3570,N_3129,N_3271);
nor U3571 (N_3571,N_3118,N_3050);
nand U3572 (N_3572,N_3137,N_3037);
nand U3573 (N_3573,N_3290,N_3168);
xor U3574 (N_3574,N_3185,N_3093);
xor U3575 (N_3575,N_3130,N_3172);
nor U3576 (N_3576,N_3267,N_3022);
nor U3577 (N_3577,N_3215,N_3147);
or U3578 (N_3578,N_3008,N_3235);
and U3579 (N_3579,N_3247,N_3016);
xnor U3580 (N_3580,N_3077,N_3141);
xor U3581 (N_3581,N_3211,N_3138);
and U3582 (N_3582,N_3124,N_3234);
or U3583 (N_3583,N_3238,N_3061);
nand U3584 (N_3584,N_3020,N_3129);
xor U3585 (N_3585,N_3031,N_3053);
xor U3586 (N_3586,N_3047,N_3219);
nor U3587 (N_3587,N_3238,N_3170);
and U3588 (N_3588,N_3268,N_3251);
nor U3589 (N_3589,N_3269,N_3198);
or U3590 (N_3590,N_3254,N_3110);
nand U3591 (N_3591,N_3298,N_3266);
nor U3592 (N_3592,N_3242,N_3151);
xnor U3593 (N_3593,N_3015,N_3044);
xor U3594 (N_3594,N_3220,N_3226);
nor U3595 (N_3595,N_3188,N_3237);
or U3596 (N_3596,N_3201,N_3199);
or U3597 (N_3597,N_3061,N_3050);
or U3598 (N_3598,N_3095,N_3243);
nand U3599 (N_3599,N_3291,N_3103);
or U3600 (N_3600,N_3519,N_3453);
nor U3601 (N_3601,N_3376,N_3509);
and U3602 (N_3602,N_3485,N_3531);
nand U3603 (N_3603,N_3366,N_3396);
and U3604 (N_3604,N_3392,N_3550);
nor U3605 (N_3605,N_3539,N_3566);
nor U3606 (N_3606,N_3456,N_3310);
or U3607 (N_3607,N_3560,N_3535);
nor U3608 (N_3608,N_3472,N_3493);
nor U3609 (N_3609,N_3551,N_3348);
nand U3610 (N_3610,N_3542,N_3352);
or U3611 (N_3611,N_3505,N_3431);
nor U3612 (N_3612,N_3450,N_3561);
nand U3613 (N_3613,N_3474,N_3572);
or U3614 (N_3614,N_3395,N_3347);
or U3615 (N_3615,N_3594,N_3574);
xnor U3616 (N_3616,N_3402,N_3552);
and U3617 (N_3617,N_3443,N_3452);
nand U3618 (N_3618,N_3406,N_3300);
nand U3619 (N_3619,N_3436,N_3422);
or U3620 (N_3620,N_3390,N_3559);
xor U3621 (N_3621,N_3394,N_3322);
and U3622 (N_3622,N_3323,N_3384);
nand U3623 (N_3623,N_3454,N_3430);
xnor U3624 (N_3624,N_3547,N_3315);
nor U3625 (N_3625,N_3438,N_3486);
or U3626 (N_3626,N_3584,N_3329);
nor U3627 (N_3627,N_3378,N_3373);
xnor U3628 (N_3628,N_3425,N_3555);
xnor U3629 (N_3629,N_3435,N_3368);
nor U3630 (N_3630,N_3421,N_3525);
xor U3631 (N_3631,N_3313,N_3499);
or U3632 (N_3632,N_3342,N_3344);
xnor U3633 (N_3633,N_3591,N_3416);
nand U3634 (N_3634,N_3334,N_3388);
nand U3635 (N_3635,N_3405,N_3426);
and U3636 (N_3636,N_3418,N_3377);
xnor U3637 (N_3637,N_3432,N_3592);
nor U3638 (N_3638,N_3403,N_3327);
nor U3639 (N_3639,N_3404,N_3595);
nor U3640 (N_3640,N_3512,N_3337);
or U3641 (N_3641,N_3549,N_3570);
nor U3642 (N_3642,N_3502,N_3571);
xor U3643 (N_3643,N_3444,N_3400);
nand U3644 (N_3644,N_3367,N_3320);
xor U3645 (N_3645,N_3356,N_3409);
or U3646 (N_3646,N_3328,N_3381);
nor U3647 (N_3647,N_3309,N_3325);
nand U3648 (N_3648,N_3412,N_3321);
and U3649 (N_3649,N_3354,N_3441);
and U3650 (N_3650,N_3335,N_3599);
or U3651 (N_3651,N_3533,N_3498);
or U3652 (N_3652,N_3480,N_3596);
nor U3653 (N_3653,N_3423,N_3428);
nor U3654 (N_3654,N_3578,N_3511);
xnor U3655 (N_3655,N_3473,N_3590);
and U3656 (N_3656,N_3350,N_3522);
nor U3657 (N_3657,N_3565,N_3410);
xnor U3658 (N_3658,N_3386,N_3538);
nand U3659 (N_3659,N_3380,N_3492);
and U3660 (N_3660,N_3437,N_3548);
nor U3661 (N_3661,N_3371,N_3382);
and U3662 (N_3662,N_3317,N_3387);
or U3663 (N_3663,N_3338,N_3439);
nand U3664 (N_3664,N_3491,N_3339);
nor U3665 (N_3665,N_3460,N_3389);
or U3666 (N_3666,N_3479,N_3484);
nand U3667 (N_3667,N_3359,N_3564);
nor U3668 (N_3668,N_3523,N_3451);
nor U3669 (N_3669,N_3581,N_3307);
and U3670 (N_3670,N_3318,N_3324);
nand U3671 (N_3671,N_3541,N_3459);
xor U3672 (N_3672,N_3407,N_3466);
or U3673 (N_3673,N_3449,N_3467);
nor U3674 (N_3674,N_3483,N_3476);
or U3675 (N_3675,N_3529,N_3575);
nor U3676 (N_3676,N_3587,N_3413);
nand U3677 (N_3677,N_3475,N_3364);
xnor U3678 (N_3678,N_3427,N_3308);
xor U3679 (N_3679,N_3557,N_3496);
xor U3680 (N_3680,N_3362,N_3341);
nand U3681 (N_3681,N_3482,N_3504);
xor U3682 (N_3682,N_3481,N_3556);
nor U3683 (N_3683,N_3363,N_3319);
and U3684 (N_3684,N_3470,N_3517);
and U3685 (N_3685,N_3536,N_3433);
nand U3686 (N_3686,N_3415,N_3417);
or U3687 (N_3687,N_3580,N_3553);
and U3688 (N_3688,N_3489,N_3440);
nor U3689 (N_3689,N_3583,N_3562);
nand U3690 (N_3690,N_3408,N_3464);
nand U3691 (N_3691,N_3497,N_3343);
xor U3692 (N_3692,N_3527,N_3465);
nor U3693 (N_3693,N_3530,N_3537);
xnor U3694 (N_3694,N_3358,N_3503);
nand U3695 (N_3695,N_3369,N_3593);
nand U3696 (N_3696,N_3361,N_3507);
and U3697 (N_3697,N_3494,N_3563);
and U3698 (N_3698,N_3520,N_3304);
nand U3699 (N_3699,N_3314,N_3501);
nand U3700 (N_3700,N_3534,N_3463);
nor U3701 (N_3701,N_3333,N_3316);
nor U3702 (N_3702,N_3442,N_3375);
and U3703 (N_3703,N_3462,N_3558);
xnor U3704 (N_3704,N_3543,N_3568);
nand U3705 (N_3705,N_3585,N_3589);
nor U3706 (N_3706,N_3516,N_3448);
and U3707 (N_3707,N_3305,N_3545);
nand U3708 (N_3708,N_3487,N_3588);
or U3709 (N_3709,N_3379,N_3488);
nand U3710 (N_3710,N_3445,N_3526);
or U3711 (N_3711,N_3420,N_3477);
nand U3712 (N_3712,N_3332,N_3579);
nor U3713 (N_3713,N_3351,N_3302);
xnor U3714 (N_3714,N_3434,N_3429);
nand U3715 (N_3715,N_3508,N_3455);
nor U3716 (N_3716,N_3424,N_3393);
or U3717 (N_3717,N_3521,N_3330);
nand U3718 (N_3718,N_3372,N_3346);
nand U3719 (N_3719,N_3411,N_3357);
nand U3720 (N_3720,N_3345,N_3401);
nand U3721 (N_3721,N_3544,N_3513);
nand U3722 (N_3722,N_3353,N_3515);
nor U3723 (N_3723,N_3471,N_3349);
or U3724 (N_3724,N_3518,N_3500);
xor U3725 (N_3725,N_3567,N_3490);
nor U3726 (N_3726,N_3365,N_3326);
xor U3727 (N_3727,N_3336,N_3554);
nor U3728 (N_3728,N_3331,N_3301);
or U3729 (N_3729,N_3398,N_3355);
nor U3730 (N_3730,N_3478,N_3528);
xor U3731 (N_3731,N_3360,N_3446);
or U3732 (N_3732,N_3370,N_3598);
and U3733 (N_3733,N_3385,N_3506);
nand U3734 (N_3734,N_3312,N_3573);
xnor U3735 (N_3735,N_3397,N_3569);
xnor U3736 (N_3736,N_3514,N_3391);
nand U3737 (N_3737,N_3577,N_3447);
and U3738 (N_3738,N_3461,N_3311);
or U3739 (N_3739,N_3340,N_3532);
nand U3740 (N_3740,N_3540,N_3576);
xnor U3741 (N_3741,N_3597,N_3524);
nand U3742 (N_3742,N_3374,N_3419);
nand U3743 (N_3743,N_3469,N_3495);
nor U3744 (N_3744,N_3582,N_3383);
xnor U3745 (N_3745,N_3546,N_3586);
and U3746 (N_3746,N_3399,N_3468);
nor U3747 (N_3747,N_3303,N_3414);
nand U3748 (N_3748,N_3510,N_3306);
xor U3749 (N_3749,N_3458,N_3457);
nand U3750 (N_3750,N_3354,N_3431);
nor U3751 (N_3751,N_3479,N_3357);
and U3752 (N_3752,N_3389,N_3492);
nand U3753 (N_3753,N_3329,N_3569);
nand U3754 (N_3754,N_3352,N_3446);
and U3755 (N_3755,N_3543,N_3428);
xor U3756 (N_3756,N_3558,N_3520);
nor U3757 (N_3757,N_3501,N_3452);
nor U3758 (N_3758,N_3538,N_3475);
or U3759 (N_3759,N_3495,N_3429);
nor U3760 (N_3760,N_3481,N_3445);
nand U3761 (N_3761,N_3438,N_3310);
and U3762 (N_3762,N_3564,N_3395);
or U3763 (N_3763,N_3340,N_3575);
xnor U3764 (N_3764,N_3470,N_3518);
nor U3765 (N_3765,N_3435,N_3573);
and U3766 (N_3766,N_3381,N_3442);
and U3767 (N_3767,N_3462,N_3514);
nand U3768 (N_3768,N_3433,N_3398);
nand U3769 (N_3769,N_3580,N_3559);
nand U3770 (N_3770,N_3577,N_3347);
or U3771 (N_3771,N_3408,N_3488);
and U3772 (N_3772,N_3347,N_3479);
xnor U3773 (N_3773,N_3413,N_3492);
xnor U3774 (N_3774,N_3511,N_3342);
or U3775 (N_3775,N_3445,N_3310);
or U3776 (N_3776,N_3435,N_3340);
nor U3777 (N_3777,N_3338,N_3464);
nand U3778 (N_3778,N_3374,N_3495);
nand U3779 (N_3779,N_3395,N_3344);
xor U3780 (N_3780,N_3392,N_3596);
nor U3781 (N_3781,N_3366,N_3359);
nor U3782 (N_3782,N_3405,N_3550);
or U3783 (N_3783,N_3548,N_3473);
or U3784 (N_3784,N_3467,N_3409);
or U3785 (N_3785,N_3566,N_3462);
and U3786 (N_3786,N_3436,N_3348);
or U3787 (N_3787,N_3583,N_3357);
nand U3788 (N_3788,N_3539,N_3457);
or U3789 (N_3789,N_3520,N_3478);
and U3790 (N_3790,N_3301,N_3430);
or U3791 (N_3791,N_3394,N_3456);
nor U3792 (N_3792,N_3404,N_3548);
xor U3793 (N_3793,N_3383,N_3453);
and U3794 (N_3794,N_3516,N_3312);
nand U3795 (N_3795,N_3554,N_3322);
nor U3796 (N_3796,N_3374,N_3556);
or U3797 (N_3797,N_3339,N_3569);
and U3798 (N_3798,N_3345,N_3520);
or U3799 (N_3799,N_3313,N_3418);
nand U3800 (N_3800,N_3442,N_3597);
nor U3801 (N_3801,N_3504,N_3562);
nand U3802 (N_3802,N_3337,N_3422);
and U3803 (N_3803,N_3443,N_3590);
and U3804 (N_3804,N_3332,N_3388);
xor U3805 (N_3805,N_3560,N_3518);
or U3806 (N_3806,N_3456,N_3549);
nand U3807 (N_3807,N_3404,N_3422);
nand U3808 (N_3808,N_3302,N_3343);
nor U3809 (N_3809,N_3431,N_3420);
nor U3810 (N_3810,N_3315,N_3539);
xnor U3811 (N_3811,N_3577,N_3410);
nor U3812 (N_3812,N_3480,N_3409);
and U3813 (N_3813,N_3460,N_3564);
and U3814 (N_3814,N_3521,N_3450);
or U3815 (N_3815,N_3413,N_3535);
nand U3816 (N_3816,N_3540,N_3592);
and U3817 (N_3817,N_3384,N_3305);
xnor U3818 (N_3818,N_3546,N_3550);
and U3819 (N_3819,N_3396,N_3463);
nand U3820 (N_3820,N_3466,N_3404);
nor U3821 (N_3821,N_3476,N_3439);
nor U3822 (N_3822,N_3588,N_3371);
nand U3823 (N_3823,N_3512,N_3398);
nand U3824 (N_3824,N_3380,N_3555);
and U3825 (N_3825,N_3574,N_3349);
or U3826 (N_3826,N_3302,N_3422);
or U3827 (N_3827,N_3490,N_3388);
or U3828 (N_3828,N_3560,N_3445);
nor U3829 (N_3829,N_3397,N_3490);
and U3830 (N_3830,N_3321,N_3550);
and U3831 (N_3831,N_3451,N_3401);
xnor U3832 (N_3832,N_3355,N_3500);
nand U3833 (N_3833,N_3574,N_3588);
and U3834 (N_3834,N_3467,N_3465);
nand U3835 (N_3835,N_3417,N_3369);
xnor U3836 (N_3836,N_3364,N_3336);
and U3837 (N_3837,N_3586,N_3344);
nand U3838 (N_3838,N_3332,N_3321);
nor U3839 (N_3839,N_3404,N_3412);
and U3840 (N_3840,N_3344,N_3518);
nand U3841 (N_3841,N_3538,N_3311);
or U3842 (N_3842,N_3383,N_3402);
xnor U3843 (N_3843,N_3587,N_3567);
nor U3844 (N_3844,N_3573,N_3411);
nand U3845 (N_3845,N_3530,N_3352);
xor U3846 (N_3846,N_3364,N_3572);
nand U3847 (N_3847,N_3311,N_3343);
nor U3848 (N_3848,N_3482,N_3354);
or U3849 (N_3849,N_3572,N_3596);
and U3850 (N_3850,N_3332,N_3570);
xnor U3851 (N_3851,N_3320,N_3427);
xnor U3852 (N_3852,N_3509,N_3454);
or U3853 (N_3853,N_3428,N_3337);
nand U3854 (N_3854,N_3583,N_3345);
nor U3855 (N_3855,N_3306,N_3493);
and U3856 (N_3856,N_3439,N_3526);
xor U3857 (N_3857,N_3419,N_3486);
or U3858 (N_3858,N_3559,N_3562);
nor U3859 (N_3859,N_3350,N_3438);
nor U3860 (N_3860,N_3409,N_3512);
nor U3861 (N_3861,N_3518,N_3415);
xnor U3862 (N_3862,N_3551,N_3376);
or U3863 (N_3863,N_3338,N_3340);
and U3864 (N_3864,N_3410,N_3475);
nand U3865 (N_3865,N_3502,N_3409);
or U3866 (N_3866,N_3474,N_3449);
xor U3867 (N_3867,N_3564,N_3327);
xnor U3868 (N_3868,N_3328,N_3395);
nand U3869 (N_3869,N_3521,N_3494);
xor U3870 (N_3870,N_3505,N_3383);
nand U3871 (N_3871,N_3440,N_3573);
and U3872 (N_3872,N_3370,N_3470);
or U3873 (N_3873,N_3597,N_3586);
xnor U3874 (N_3874,N_3594,N_3357);
xor U3875 (N_3875,N_3580,N_3451);
or U3876 (N_3876,N_3301,N_3328);
or U3877 (N_3877,N_3398,N_3389);
nor U3878 (N_3878,N_3505,N_3341);
or U3879 (N_3879,N_3367,N_3526);
nand U3880 (N_3880,N_3372,N_3317);
nor U3881 (N_3881,N_3554,N_3333);
xnor U3882 (N_3882,N_3595,N_3456);
xnor U3883 (N_3883,N_3504,N_3377);
nand U3884 (N_3884,N_3398,N_3338);
nand U3885 (N_3885,N_3512,N_3311);
and U3886 (N_3886,N_3501,N_3531);
nand U3887 (N_3887,N_3355,N_3479);
and U3888 (N_3888,N_3505,N_3443);
or U3889 (N_3889,N_3432,N_3420);
nor U3890 (N_3890,N_3360,N_3409);
nor U3891 (N_3891,N_3323,N_3360);
and U3892 (N_3892,N_3381,N_3534);
and U3893 (N_3893,N_3451,N_3320);
and U3894 (N_3894,N_3528,N_3560);
xor U3895 (N_3895,N_3391,N_3541);
nand U3896 (N_3896,N_3350,N_3314);
and U3897 (N_3897,N_3522,N_3472);
nor U3898 (N_3898,N_3562,N_3405);
and U3899 (N_3899,N_3517,N_3344);
nor U3900 (N_3900,N_3729,N_3817);
nor U3901 (N_3901,N_3809,N_3833);
and U3902 (N_3902,N_3705,N_3764);
and U3903 (N_3903,N_3653,N_3664);
xor U3904 (N_3904,N_3812,N_3709);
xnor U3905 (N_3905,N_3726,N_3756);
nor U3906 (N_3906,N_3630,N_3800);
nand U3907 (N_3907,N_3893,N_3623);
xor U3908 (N_3908,N_3686,N_3641);
and U3909 (N_3909,N_3752,N_3747);
and U3910 (N_3910,N_3811,N_3768);
or U3911 (N_3911,N_3801,N_3652);
xnor U3912 (N_3912,N_3642,N_3829);
nor U3913 (N_3913,N_3616,N_3745);
nor U3914 (N_3914,N_3852,N_3802);
xnor U3915 (N_3915,N_3771,N_3750);
nand U3916 (N_3916,N_3877,N_3883);
xnor U3917 (N_3917,N_3660,N_3763);
nor U3918 (N_3918,N_3897,N_3684);
or U3919 (N_3919,N_3678,N_3673);
or U3920 (N_3920,N_3823,N_3733);
nor U3921 (N_3921,N_3730,N_3867);
and U3922 (N_3922,N_3798,N_3795);
or U3923 (N_3923,N_3741,N_3714);
nor U3924 (N_3924,N_3634,N_3807);
and U3925 (N_3925,N_3813,N_3739);
and U3926 (N_3926,N_3786,N_3721);
xnor U3927 (N_3927,N_3851,N_3853);
and U3928 (N_3928,N_3845,N_3815);
or U3929 (N_3929,N_3693,N_3655);
xnor U3930 (N_3930,N_3870,N_3791);
xnor U3931 (N_3931,N_3844,N_3662);
xor U3932 (N_3932,N_3777,N_3769);
xnor U3933 (N_3933,N_3609,N_3638);
xor U3934 (N_3934,N_3627,N_3842);
or U3935 (N_3935,N_3694,N_3683);
or U3936 (N_3936,N_3849,N_3793);
and U3937 (N_3937,N_3781,N_3792);
and U3938 (N_3938,N_3724,N_3881);
and U3939 (N_3939,N_3799,N_3816);
nor U3940 (N_3940,N_3884,N_3751);
or U3941 (N_3941,N_3888,N_3688);
nor U3942 (N_3942,N_3676,N_3855);
or U3943 (N_3943,N_3667,N_3622);
nand U3944 (N_3944,N_3645,N_3703);
and U3945 (N_3945,N_3766,N_3654);
or U3946 (N_3946,N_3722,N_3889);
or U3947 (N_3947,N_3699,N_3628);
nand U3948 (N_3948,N_3732,N_3675);
and U3949 (N_3949,N_3651,N_3707);
or U3950 (N_3950,N_3615,N_3898);
xor U3951 (N_3951,N_3869,N_3647);
and U3952 (N_3952,N_3697,N_3794);
xor U3953 (N_3953,N_3743,N_3600);
nand U3954 (N_3954,N_3748,N_3740);
or U3955 (N_3955,N_3687,N_3880);
nor U3956 (N_3956,N_3725,N_3830);
and U3957 (N_3957,N_3661,N_3755);
and U3958 (N_3958,N_3831,N_3779);
nand U3959 (N_3959,N_3850,N_3843);
nor U3960 (N_3960,N_3882,N_3737);
nor U3961 (N_3961,N_3734,N_3742);
nor U3962 (N_3962,N_3758,N_3706);
nand U3963 (N_3963,N_3840,N_3787);
nor U3964 (N_3964,N_3859,N_3857);
xor U3965 (N_3965,N_3778,N_3610);
xnor U3966 (N_3966,N_3695,N_3681);
xor U3967 (N_3967,N_3617,N_3670);
nor U3968 (N_3968,N_3605,N_3864);
nand U3969 (N_3969,N_3814,N_3760);
nor U3970 (N_3970,N_3873,N_3780);
xnor U3971 (N_3971,N_3846,N_3735);
nor U3972 (N_3972,N_3784,N_3773);
or U3973 (N_3973,N_3677,N_3818);
and U3974 (N_3974,N_3728,N_3639);
or U3975 (N_3975,N_3736,N_3636);
nor U3976 (N_3976,N_3796,N_3841);
or U3977 (N_3977,N_3650,N_3701);
xor U3978 (N_3978,N_3637,N_3629);
xor U3979 (N_3979,N_3608,N_3828);
xor U3980 (N_3980,N_3607,N_3878);
and U3981 (N_3981,N_3754,N_3723);
nor U3982 (N_3982,N_3863,N_3892);
nor U3983 (N_3983,N_3865,N_3761);
or U3984 (N_3984,N_3682,N_3620);
nand U3985 (N_3985,N_3663,N_3879);
or U3986 (N_3986,N_3614,N_3895);
and U3987 (N_3987,N_3866,N_3790);
or U3988 (N_3988,N_3770,N_3659);
and U3989 (N_3989,N_3890,N_3899);
xnor U3990 (N_3990,N_3718,N_3789);
and U3991 (N_3991,N_3797,N_3804);
nand U3992 (N_3992,N_3753,N_3657);
nand U3993 (N_3993,N_3861,N_3698);
and U3994 (N_3994,N_3679,N_3690);
and U3995 (N_3995,N_3656,N_3826);
nor U3996 (N_3996,N_3819,N_3854);
or U3997 (N_3997,N_3788,N_3765);
nor U3998 (N_3998,N_3702,N_3716);
nor U3999 (N_3999,N_3824,N_3658);
nor U4000 (N_4000,N_3689,N_3624);
and U4001 (N_4001,N_3633,N_3783);
or U4002 (N_4002,N_3820,N_3680);
nand U4003 (N_4003,N_3810,N_3710);
nand U4004 (N_4004,N_3834,N_3875);
and U4005 (N_4005,N_3837,N_3640);
nand U4006 (N_4006,N_3731,N_3772);
xor U4007 (N_4007,N_3625,N_3603);
or U4008 (N_4008,N_3874,N_3708);
nor U4009 (N_4009,N_3757,N_3744);
or U4010 (N_4010,N_3612,N_3775);
xor U4011 (N_4011,N_3604,N_3711);
or U4012 (N_4012,N_3644,N_3871);
or U4013 (N_4013,N_3805,N_3808);
nor U4014 (N_4014,N_3776,N_3782);
xor U4015 (N_4015,N_3832,N_3611);
xnor U4016 (N_4016,N_3719,N_3685);
or U4017 (N_4017,N_3749,N_3692);
nand U4018 (N_4018,N_3891,N_3876);
or U4019 (N_4019,N_3806,N_3602);
or U4020 (N_4020,N_3666,N_3836);
and U4021 (N_4021,N_3606,N_3872);
and U4022 (N_4022,N_3613,N_3648);
xor U4023 (N_4023,N_3886,N_3700);
nand U4024 (N_4024,N_3774,N_3720);
nand U4025 (N_4025,N_3621,N_3860);
nor U4026 (N_4026,N_3618,N_3619);
nor U4027 (N_4027,N_3649,N_3835);
and U4028 (N_4028,N_3767,N_3868);
and U4029 (N_4029,N_3746,N_3759);
or U4030 (N_4030,N_3821,N_3825);
nand U4031 (N_4031,N_3635,N_3738);
or U4032 (N_4032,N_3838,N_3626);
xor U4033 (N_4033,N_3674,N_3727);
nor U4034 (N_4034,N_3856,N_3669);
and U4035 (N_4035,N_3762,N_3712);
xnor U4036 (N_4036,N_3665,N_3785);
nor U4037 (N_4037,N_3803,N_3847);
nand U4038 (N_4038,N_3894,N_3862);
nor U4039 (N_4039,N_3717,N_3646);
nand U4040 (N_4040,N_3672,N_3887);
or U4041 (N_4041,N_3715,N_3696);
nand U4042 (N_4042,N_3713,N_3643);
or U4043 (N_4043,N_3827,N_3896);
or U4044 (N_4044,N_3668,N_3848);
nand U4045 (N_4045,N_3671,N_3885);
and U4046 (N_4046,N_3704,N_3839);
xor U4047 (N_4047,N_3632,N_3822);
or U4048 (N_4048,N_3601,N_3858);
xnor U4049 (N_4049,N_3631,N_3691);
xnor U4050 (N_4050,N_3845,N_3745);
xnor U4051 (N_4051,N_3860,N_3696);
nand U4052 (N_4052,N_3757,N_3827);
and U4053 (N_4053,N_3668,N_3691);
nor U4054 (N_4054,N_3609,N_3830);
nand U4055 (N_4055,N_3872,N_3791);
xnor U4056 (N_4056,N_3739,N_3748);
or U4057 (N_4057,N_3722,N_3779);
nand U4058 (N_4058,N_3642,N_3869);
xnor U4059 (N_4059,N_3852,N_3709);
xnor U4060 (N_4060,N_3647,N_3855);
or U4061 (N_4061,N_3619,N_3716);
xor U4062 (N_4062,N_3883,N_3645);
nand U4063 (N_4063,N_3804,N_3880);
nand U4064 (N_4064,N_3884,N_3732);
xnor U4065 (N_4065,N_3763,N_3779);
and U4066 (N_4066,N_3832,N_3772);
and U4067 (N_4067,N_3849,N_3615);
or U4068 (N_4068,N_3679,N_3817);
nand U4069 (N_4069,N_3884,N_3625);
and U4070 (N_4070,N_3899,N_3700);
nor U4071 (N_4071,N_3753,N_3840);
nand U4072 (N_4072,N_3715,N_3723);
xnor U4073 (N_4073,N_3749,N_3762);
xor U4074 (N_4074,N_3717,N_3607);
nor U4075 (N_4075,N_3705,N_3817);
nand U4076 (N_4076,N_3723,N_3882);
xnor U4077 (N_4077,N_3827,N_3604);
xor U4078 (N_4078,N_3840,N_3644);
xor U4079 (N_4079,N_3859,N_3771);
or U4080 (N_4080,N_3846,N_3758);
nor U4081 (N_4081,N_3641,N_3874);
nand U4082 (N_4082,N_3829,N_3674);
nor U4083 (N_4083,N_3797,N_3853);
and U4084 (N_4084,N_3607,N_3783);
xor U4085 (N_4085,N_3689,N_3641);
xnor U4086 (N_4086,N_3623,N_3711);
xor U4087 (N_4087,N_3841,N_3750);
or U4088 (N_4088,N_3740,N_3724);
xor U4089 (N_4089,N_3796,N_3645);
nand U4090 (N_4090,N_3719,N_3756);
or U4091 (N_4091,N_3736,N_3653);
or U4092 (N_4092,N_3821,N_3672);
xor U4093 (N_4093,N_3848,N_3873);
xor U4094 (N_4094,N_3673,N_3630);
xnor U4095 (N_4095,N_3711,N_3624);
and U4096 (N_4096,N_3744,N_3775);
xnor U4097 (N_4097,N_3897,N_3873);
and U4098 (N_4098,N_3716,N_3638);
nor U4099 (N_4099,N_3619,N_3611);
or U4100 (N_4100,N_3741,N_3655);
nand U4101 (N_4101,N_3899,N_3805);
nand U4102 (N_4102,N_3862,N_3732);
nor U4103 (N_4103,N_3876,N_3633);
nand U4104 (N_4104,N_3646,N_3834);
or U4105 (N_4105,N_3858,N_3869);
nor U4106 (N_4106,N_3885,N_3882);
nor U4107 (N_4107,N_3801,N_3620);
xor U4108 (N_4108,N_3851,N_3620);
and U4109 (N_4109,N_3837,N_3678);
nand U4110 (N_4110,N_3716,N_3632);
and U4111 (N_4111,N_3639,N_3625);
nor U4112 (N_4112,N_3763,N_3635);
nor U4113 (N_4113,N_3762,N_3687);
or U4114 (N_4114,N_3843,N_3648);
nand U4115 (N_4115,N_3659,N_3674);
nand U4116 (N_4116,N_3808,N_3656);
and U4117 (N_4117,N_3729,N_3780);
and U4118 (N_4118,N_3645,N_3862);
nor U4119 (N_4119,N_3885,N_3723);
nand U4120 (N_4120,N_3603,N_3705);
and U4121 (N_4121,N_3684,N_3649);
nor U4122 (N_4122,N_3739,N_3678);
nand U4123 (N_4123,N_3762,N_3624);
and U4124 (N_4124,N_3861,N_3619);
nand U4125 (N_4125,N_3858,N_3849);
or U4126 (N_4126,N_3697,N_3893);
or U4127 (N_4127,N_3776,N_3882);
or U4128 (N_4128,N_3620,N_3657);
xor U4129 (N_4129,N_3835,N_3601);
xnor U4130 (N_4130,N_3635,N_3707);
and U4131 (N_4131,N_3686,N_3608);
and U4132 (N_4132,N_3755,N_3882);
or U4133 (N_4133,N_3804,N_3860);
nand U4134 (N_4134,N_3749,N_3709);
and U4135 (N_4135,N_3736,N_3605);
xor U4136 (N_4136,N_3890,N_3645);
xnor U4137 (N_4137,N_3646,N_3665);
or U4138 (N_4138,N_3871,N_3647);
and U4139 (N_4139,N_3603,N_3897);
or U4140 (N_4140,N_3860,N_3603);
xor U4141 (N_4141,N_3626,N_3705);
nor U4142 (N_4142,N_3757,N_3777);
nand U4143 (N_4143,N_3624,N_3875);
or U4144 (N_4144,N_3651,N_3868);
nand U4145 (N_4145,N_3613,N_3853);
nand U4146 (N_4146,N_3843,N_3894);
and U4147 (N_4147,N_3882,N_3654);
and U4148 (N_4148,N_3758,N_3733);
nand U4149 (N_4149,N_3754,N_3760);
xor U4150 (N_4150,N_3894,N_3779);
xor U4151 (N_4151,N_3764,N_3757);
nor U4152 (N_4152,N_3862,N_3633);
or U4153 (N_4153,N_3650,N_3785);
nor U4154 (N_4154,N_3702,N_3759);
xor U4155 (N_4155,N_3775,N_3780);
xor U4156 (N_4156,N_3833,N_3778);
nor U4157 (N_4157,N_3753,N_3880);
nor U4158 (N_4158,N_3883,N_3713);
or U4159 (N_4159,N_3661,N_3757);
xor U4160 (N_4160,N_3704,N_3794);
nor U4161 (N_4161,N_3608,N_3771);
nand U4162 (N_4162,N_3789,N_3744);
xnor U4163 (N_4163,N_3861,N_3716);
and U4164 (N_4164,N_3613,N_3747);
or U4165 (N_4165,N_3733,N_3855);
and U4166 (N_4166,N_3863,N_3884);
and U4167 (N_4167,N_3705,N_3789);
nor U4168 (N_4168,N_3823,N_3645);
nand U4169 (N_4169,N_3682,N_3697);
xnor U4170 (N_4170,N_3650,N_3853);
and U4171 (N_4171,N_3694,N_3812);
nand U4172 (N_4172,N_3727,N_3603);
or U4173 (N_4173,N_3873,N_3790);
xnor U4174 (N_4174,N_3717,N_3817);
nand U4175 (N_4175,N_3892,N_3781);
and U4176 (N_4176,N_3815,N_3627);
nor U4177 (N_4177,N_3736,N_3754);
xnor U4178 (N_4178,N_3735,N_3882);
nand U4179 (N_4179,N_3631,N_3739);
xor U4180 (N_4180,N_3827,N_3602);
and U4181 (N_4181,N_3875,N_3830);
xor U4182 (N_4182,N_3758,N_3713);
nor U4183 (N_4183,N_3841,N_3623);
or U4184 (N_4184,N_3855,N_3704);
nand U4185 (N_4185,N_3635,N_3625);
nand U4186 (N_4186,N_3717,N_3609);
or U4187 (N_4187,N_3726,N_3669);
and U4188 (N_4188,N_3812,N_3894);
xor U4189 (N_4189,N_3743,N_3726);
or U4190 (N_4190,N_3779,N_3752);
and U4191 (N_4191,N_3655,N_3889);
and U4192 (N_4192,N_3878,N_3714);
or U4193 (N_4193,N_3701,N_3700);
or U4194 (N_4194,N_3876,N_3650);
nand U4195 (N_4195,N_3631,N_3829);
nor U4196 (N_4196,N_3695,N_3867);
nor U4197 (N_4197,N_3700,N_3699);
nor U4198 (N_4198,N_3769,N_3635);
or U4199 (N_4199,N_3846,N_3668);
nor U4200 (N_4200,N_4080,N_3949);
nor U4201 (N_4201,N_3931,N_4098);
nor U4202 (N_4202,N_4094,N_4062);
nor U4203 (N_4203,N_4029,N_4139);
xnor U4204 (N_4204,N_4085,N_4096);
xnor U4205 (N_4205,N_4008,N_4084);
and U4206 (N_4206,N_3942,N_3920);
nor U4207 (N_4207,N_4107,N_4103);
and U4208 (N_4208,N_4081,N_4063);
nor U4209 (N_4209,N_4007,N_4006);
xnor U4210 (N_4210,N_4020,N_4067);
or U4211 (N_4211,N_4071,N_3990);
and U4212 (N_4212,N_4023,N_4050);
xnor U4213 (N_4213,N_3930,N_4091);
and U4214 (N_4214,N_3985,N_4013);
or U4215 (N_4215,N_4053,N_4021);
and U4216 (N_4216,N_4117,N_4001);
nand U4217 (N_4217,N_3991,N_4129);
nor U4218 (N_4218,N_4137,N_3998);
and U4219 (N_4219,N_3923,N_4090);
and U4220 (N_4220,N_4082,N_4069);
or U4221 (N_4221,N_4000,N_3933);
or U4222 (N_4222,N_3962,N_3973);
and U4223 (N_4223,N_3992,N_4189);
xor U4224 (N_4224,N_4036,N_4131);
nand U4225 (N_4225,N_4047,N_4190);
nor U4226 (N_4226,N_3905,N_4054);
xnor U4227 (N_4227,N_3906,N_3925);
and U4228 (N_4228,N_4167,N_3944);
and U4229 (N_4229,N_4128,N_4198);
xor U4230 (N_4230,N_3922,N_4064);
and U4231 (N_4231,N_4015,N_4162);
nand U4232 (N_4232,N_4105,N_3980);
xor U4233 (N_4233,N_4161,N_4159);
or U4234 (N_4234,N_4176,N_3907);
nor U4235 (N_4235,N_3929,N_4175);
nand U4236 (N_4236,N_4030,N_4018);
or U4237 (N_4237,N_3978,N_4123);
nand U4238 (N_4238,N_3952,N_4019);
and U4239 (N_4239,N_3977,N_4075);
or U4240 (N_4240,N_4092,N_4174);
nor U4241 (N_4241,N_4126,N_3921);
nand U4242 (N_4242,N_4114,N_3967);
or U4243 (N_4243,N_4102,N_3986);
nand U4244 (N_4244,N_3916,N_4004);
nand U4245 (N_4245,N_3918,N_4101);
nor U4246 (N_4246,N_4058,N_4164);
and U4247 (N_4247,N_4165,N_3914);
nand U4248 (N_4248,N_3976,N_4150);
nand U4249 (N_4249,N_4099,N_4136);
nor U4250 (N_4250,N_4012,N_3945);
nor U4251 (N_4251,N_3934,N_3951);
nor U4252 (N_4252,N_3956,N_4119);
and U4253 (N_4253,N_4073,N_4017);
and U4254 (N_4254,N_3917,N_4028);
or U4255 (N_4255,N_3983,N_4025);
nor U4256 (N_4256,N_4037,N_3997);
and U4257 (N_4257,N_4118,N_4169);
or U4258 (N_4258,N_4186,N_4056);
nor U4259 (N_4259,N_4158,N_4040);
xnor U4260 (N_4260,N_4193,N_3919);
nand U4261 (N_4261,N_4111,N_4044);
xor U4262 (N_4262,N_4035,N_4183);
xnor U4263 (N_4263,N_3959,N_4177);
or U4264 (N_4264,N_4005,N_3947);
nand U4265 (N_4265,N_4170,N_4066);
xnor U4266 (N_4266,N_4009,N_4187);
nand U4267 (N_4267,N_4196,N_4087);
nor U4268 (N_4268,N_4083,N_3960);
and U4269 (N_4269,N_4145,N_4199);
or U4270 (N_4270,N_4048,N_3910);
xor U4271 (N_4271,N_4022,N_4153);
and U4272 (N_4272,N_3943,N_4110);
nor U4273 (N_4273,N_3989,N_4024);
or U4274 (N_4274,N_4124,N_3957);
or U4275 (N_4275,N_3927,N_4109);
xnor U4276 (N_4276,N_4031,N_3996);
nand U4277 (N_4277,N_3902,N_4016);
nand U4278 (N_4278,N_4144,N_4141);
or U4279 (N_4279,N_4104,N_3950);
xnor U4280 (N_4280,N_4070,N_4149);
nor U4281 (N_4281,N_4130,N_4055);
and U4282 (N_4282,N_4160,N_3994);
nor U4283 (N_4283,N_4045,N_4168);
xor U4284 (N_4284,N_4122,N_4052);
nand U4285 (N_4285,N_4078,N_4138);
xnor U4286 (N_4286,N_4106,N_4039);
nor U4287 (N_4287,N_4059,N_4068);
nand U4288 (N_4288,N_4108,N_4086);
and U4289 (N_4289,N_4076,N_4194);
or U4290 (N_4290,N_3995,N_4157);
nand U4291 (N_4291,N_4182,N_4195);
nand U4292 (N_4292,N_3909,N_3932);
or U4293 (N_4293,N_4046,N_3941);
xor U4294 (N_4294,N_4065,N_4002);
xor U4295 (N_4295,N_3948,N_4115);
nor U4296 (N_4296,N_4155,N_3975);
xnor U4297 (N_4297,N_4188,N_3954);
nor U4298 (N_4298,N_3970,N_4151);
xor U4299 (N_4299,N_3984,N_3913);
xor U4300 (N_4300,N_4043,N_3940);
nor U4301 (N_4301,N_3968,N_4113);
nor U4302 (N_4302,N_4125,N_3955);
and U4303 (N_4303,N_3972,N_4191);
nand U4304 (N_4304,N_3928,N_4032);
nand U4305 (N_4305,N_4135,N_4148);
and U4306 (N_4306,N_4184,N_4163);
nor U4307 (N_4307,N_4171,N_4133);
xor U4308 (N_4308,N_4192,N_4116);
and U4309 (N_4309,N_4180,N_4088);
xnor U4310 (N_4310,N_4112,N_4172);
and U4311 (N_4311,N_3993,N_3988);
nor U4312 (N_4312,N_3982,N_4156);
nor U4313 (N_4313,N_3966,N_3999);
nor U4314 (N_4314,N_4197,N_4097);
or U4315 (N_4315,N_4041,N_3961);
nand U4316 (N_4316,N_4147,N_4079);
nand U4317 (N_4317,N_3912,N_3911);
nand U4318 (N_4318,N_3981,N_3965);
or U4319 (N_4319,N_4034,N_4132);
and U4320 (N_4320,N_4181,N_4185);
nor U4321 (N_4321,N_4003,N_4093);
xnor U4322 (N_4322,N_3903,N_4061);
xor U4323 (N_4323,N_3908,N_4027);
nor U4324 (N_4324,N_4121,N_3926);
nor U4325 (N_4325,N_3974,N_3924);
and U4326 (N_4326,N_3937,N_4152);
xor U4327 (N_4327,N_4077,N_4049);
and U4328 (N_4328,N_4095,N_3953);
nor U4329 (N_4329,N_3987,N_3971);
nand U4330 (N_4330,N_3936,N_4166);
or U4331 (N_4331,N_4146,N_4100);
and U4332 (N_4332,N_4089,N_4173);
nor U4333 (N_4333,N_4010,N_4154);
xnor U4334 (N_4334,N_4051,N_4072);
nor U4335 (N_4335,N_4178,N_3904);
or U4336 (N_4336,N_3900,N_3979);
xnor U4337 (N_4337,N_3963,N_3915);
xnor U4338 (N_4338,N_4026,N_4074);
nor U4339 (N_4339,N_4011,N_3946);
nand U4340 (N_4340,N_4057,N_3901);
and U4341 (N_4341,N_4060,N_3958);
or U4342 (N_4342,N_4038,N_4134);
or U4343 (N_4343,N_4042,N_4120);
and U4344 (N_4344,N_4014,N_3939);
nand U4345 (N_4345,N_4033,N_4179);
xnor U4346 (N_4346,N_3964,N_4142);
xor U4347 (N_4347,N_4127,N_3938);
nand U4348 (N_4348,N_4140,N_4143);
and U4349 (N_4349,N_3969,N_3935);
nand U4350 (N_4350,N_4188,N_4015);
nor U4351 (N_4351,N_4075,N_4195);
xnor U4352 (N_4352,N_3940,N_4056);
nand U4353 (N_4353,N_4049,N_4099);
and U4354 (N_4354,N_4110,N_3911);
nor U4355 (N_4355,N_3933,N_3946);
xor U4356 (N_4356,N_3945,N_4068);
or U4357 (N_4357,N_4147,N_3985);
nand U4358 (N_4358,N_4092,N_4164);
nor U4359 (N_4359,N_4166,N_3991);
and U4360 (N_4360,N_3995,N_3956);
and U4361 (N_4361,N_4126,N_4141);
nand U4362 (N_4362,N_4053,N_3971);
nand U4363 (N_4363,N_4154,N_4049);
nor U4364 (N_4364,N_4048,N_4108);
and U4365 (N_4365,N_4090,N_4147);
nand U4366 (N_4366,N_4061,N_3977);
xnor U4367 (N_4367,N_3957,N_3981);
or U4368 (N_4368,N_4026,N_4040);
xor U4369 (N_4369,N_4122,N_3903);
xor U4370 (N_4370,N_4089,N_3938);
and U4371 (N_4371,N_3987,N_4081);
or U4372 (N_4372,N_3953,N_4169);
or U4373 (N_4373,N_4050,N_3922);
and U4374 (N_4374,N_4045,N_3942);
nor U4375 (N_4375,N_3946,N_4044);
nor U4376 (N_4376,N_4117,N_3913);
xnor U4377 (N_4377,N_4130,N_4160);
and U4378 (N_4378,N_4135,N_4036);
or U4379 (N_4379,N_4082,N_4163);
xor U4380 (N_4380,N_4117,N_4093);
or U4381 (N_4381,N_4036,N_4082);
or U4382 (N_4382,N_4152,N_4113);
or U4383 (N_4383,N_4198,N_4074);
xnor U4384 (N_4384,N_4081,N_3962);
nand U4385 (N_4385,N_4159,N_4042);
or U4386 (N_4386,N_4198,N_4070);
or U4387 (N_4387,N_4170,N_3903);
nor U4388 (N_4388,N_4089,N_3936);
or U4389 (N_4389,N_4001,N_3927);
xor U4390 (N_4390,N_4179,N_3928);
nor U4391 (N_4391,N_4088,N_3949);
xnor U4392 (N_4392,N_4027,N_4029);
nand U4393 (N_4393,N_4182,N_4107);
nand U4394 (N_4394,N_3922,N_4042);
or U4395 (N_4395,N_4042,N_3959);
xnor U4396 (N_4396,N_4068,N_4170);
nor U4397 (N_4397,N_4102,N_4141);
xor U4398 (N_4398,N_4024,N_4067);
and U4399 (N_4399,N_3946,N_4170);
nor U4400 (N_4400,N_4013,N_4037);
nor U4401 (N_4401,N_4152,N_4159);
nor U4402 (N_4402,N_3911,N_4112);
nand U4403 (N_4403,N_4097,N_4137);
nor U4404 (N_4404,N_4111,N_3906);
xnor U4405 (N_4405,N_3960,N_4170);
nor U4406 (N_4406,N_3987,N_3947);
xnor U4407 (N_4407,N_3960,N_3914);
nor U4408 (N_4408,N_4144,N_4086);
nand U4409 (N_4409,N_4030,N_3923);
nor U4410 (N_4410,N_4156,N_4159);
xor U4411 (N_4411,N_3910,N_4159);
and U4412 (N_4412,N_4020,N_4123);
and U4413 (N_4413,N_3993,N_4100);
xnor U4414 (N_4414,N_3966,N_3916);
xnor U4415 (N_4415,N_4199,N_4177);
or U4416 (N_4416,N_4091,N_4018);
xor U4417 (N_4417,N_4121,N_3923);
nand U4418 (N_4418,N_4095,N_4115);
nand U4419 (N_4419,N_4121,N_4052);
xnor U4420 (N_4420,N_4040,N_3951);
xnor U4421 (N_4421,N_3937,N_3962);
xnor U4422 (N_4422,N_3902,N_4030);
or U4423 (N_4423,N_4104,N_4151);
nor U4424 (N_4424,N_4026,N_3968);
and U4425 (N_4425,N_4011,N_4062);
nand U4426 (N_4426,N_3960,N_4122);
and U4427 (N_4427,N_3981,N_3916);
or U4428 (N_4428,N_3945,N_3968);
and U4429 (N_4429,N_3905,N_4091);
or U4430 (N_4430,N_3970,N_3935);
xor U4431 (N_4431,N_3975,N_3971);
and U4432 (N_4432,N_3966,N_4029);
nor U4433 (N_4433,N_3988,N_4072);
nand U4434 (N_4434,N_4103,N_3934);
nor U4435 (N_4435,N_3925,N_4192);
and U4436 (N_4436,N_4140,N_4135);
xnor U4437 (N_4437,N_3984,N_4147);
or U4438 (N_4438,N_3930,N_4182);
and U4439 (N_4439,N_4033,N_4089);
and U4440 (N_4440,N_3962,N_4155);
xnor U4441 (N_4441,N_3927,N_3961);
xor U4442 (N_4442,N_4165,N_4184);
and U4443 (N_4443,N_3962,N_4142);
or U4444 (N_4444,N_4030,N_4174);
xnor U4445 (N_4445,N_4012,N_3980);
or U4446 (N_4446,N_3952,N_4115);
and U4447 (N_4447,N_3950,N_4191);
and U4448 (N_4448,N_4028,N_4022);
nor U4449 (N_4449,N_4159,N_4087);
and U4450 (N_4450,N_3934,N_4079);
and U4451 (N_4451,N_4175,N_4112);
or U4452 (N_4452,N_4159,N_4095);
nand U4453 (N_4453,N_4161,N_4056);
or U4454 (N_4454,N_4020,N_4146);
nor U4455 (N_4455,N_3919,N_4167);
nor U4456 (N_4456,N_3921,N_4035);
and U4457 (N_4457,N_4075,N_4096);
or U4458 (N_4458,N_4165,N_4177);
or U4459 (N_4459,N_3975,N_4072);
nor U4460 (N_4460,N_3910,N_3966);
xor U4461 (N_4461,N_4106,N_4111);
nand U4462 (N_4462,N_3936,N_3931);
nor U4463 (N_4463,N_4071,N_4022);
nor U4464 (N_4464,N_3988,N_3974);
and U4465 (N_4465,N_4163,N_4040);
xnor U4466 (N_4466,N_4132,N_3989);
and U4467 (N_4467,N_3990,N_4193);
nand U4468 (N_4468,N_4179,N_3905);
nor U4469 (N_4469,N_4091,N_4074);
or U4470 (N_4470,N_3969,N_4076);
or U4471 (N_4471,N_4102,N_3980);
and U4472 (N_4472,N_4184,N_3908);
nor U4473 (N_4473,N_4164,N_3913);
xor U4474 (N_4474,N_4089,N_4012);
and U4475 (N_4475,N_4088,N_3915);
and U4476 (N_4476,N_4118,N_4058);
nand U4477 (N_4477,N_4187,N_4087);
xnor U4478 (N_4478,N_3906,N_4008);
xnor U4479 (N_4479,N_3969,N_3938);
nor U4480 (N_4480,N_4022,N_3942);
and U4481 (N_4481,N_4183,N_4057);
nor U4482 (N_4482,N_3974,N_4022);
nand U4483 (N_4483,N_3902,N_4109);
nand U4484 (N_4484,N_4039,N_4011);
nand U4485 (N_4485,N_4105,N_4117);
or U4486 (N_4486,N_4192,N_4169);
and U4487 (N_4487,N_4085,N_4180);
and U4488 (N_4488,N_4091,N_4171);
or U4489 (N_4489,N_3999,N_3926);
or U4490 (N_4490,N_3927,N_4006);
nor U4491 (N_4491,N_4037,N_4121);
and U4492 (N_4492,N_4089,N_4114);
nand U4493 (N_4493,N_4064,N_3965);
xnor U4494 (N_4494,N_3955,N_4046);
xnor U4495 (N_4495,N_3948,N_4150);
xor U4496 (N_4496,N_4177,N_4004);
nand U4497 (N_4497,N_4124,N_4000);
nand U4498 (N_4498,N_3921,N_4032);
or U4499 (N_4499,N_3952,N_3902);
or U4500 (N_4500,N_4356,N_4209);
nor U4501 (N_4501,N_4304,N_4447);
or U4502 (N_4502,N_4492,N_4262);
and U4503 (N_4503,N_4302,N_4458);
xnor U4504 (N_4504,N_4359,N_4497);
nand U4505 (N_4505,N_4316,N_4235);
nor U4506 (N_4506,N_4472,N_4468);
or U4507 (N_4507,N_4210,N_4292);
xnor U4508 (N_4508,N_4330,N_4365);
and U4509 (N_4509,N_4481,N_4342);
nand U4510 (N_4510,N_4445,N_4207);
and U4511 (N_4511,N_4312,N_4275);
and U4512 (N_4512,N_4483,N_4352);
nand U4513 (N_4513,N_4449,N_4269);
xnor U4514 (N_4514,N_4278,N_4396);
nor U4515 (N_4515,N_4250,N_4287);
nand U4516 (N_4516,N_4482,N_4248);
nor U4517 (N_4517,N_4424,N_4421);
nor U4518 (N_4518,N_4344,N_4239);
nand U4519 (N_4519,N_4299,N_4280);
xor U4520 (N_4520,N_4266,N_4470);
nor U4521 (N_4521,N_4383,N_4440);
xnor U4522 (N_4522,N_4335,N_4363);
and U4523 (N_4523,N_4325,N_4347);
and U4524 (N_4524,N_4350,N_4362);
and U4525 (N_4525,N_4341,N_4361);
and U4526 (N_4526,N_4498,N_4446);
nor U4527 (N_4527,N_4283,N_4204);
nand U4528 (N_4528,N_4375,N_4234);
xor U4529 (N_4529,N_4276,N_4442);
nand U4530 (N_4530,N_4386,N_4271);
xor U4531 (N_4531,N_4247,N_4473);
and U4532 (N_4532,N_4268,N_4411);
and U4533 (N_4533,N_4406,N_4264);
nand U4534 (N_4534,N_4286,N_4486);
and U4535 (N_4535,N_4322,N_4318);
or U4536 (N_4536,N_4380,N_4360);
xor U4537 (N_4537,N_4422,N_4461);
nor U4538 (N_4538,N_4412,N_4487);
nand U4539 (N_4539,N_4214,N_4326);
and U4540 (N_4540,N_4374,N_4457);
and U4541 (N_4541,N_4414,N_4246);
or U4542 (N_4542,N_4252,N_4218);
nand U4543 (N_4543,N_4355,N_4391);
nor U4544 (N_4544,N_4290,N_4379);
or U4545 (N_4545,N_4345,N_4272);
xor U4546 (N_4546,N_4392,N_4439);
xor U4547 (N_4547,N_4490,N_4393);
or U4548 (N_4548,N_4381,N_4333);
nand U4549 (N_4549,N_4428,N_4229);
nand U4550 (N_4550,N_4443,N_4479);
xor U4551 (N_4551,N_4223,N_4233);
nor U4552 (N_4552,N_4477,N_4201);
xnor U4553 (N_4553,N_4426,N_4491);
or U4554 (N_4554,N_4225,N_4346);
or U4555 (N_4555,N_4489,N_4314);
and U4556 (N_4556,N_4432,N_4237);
nand U4557 (N_4557,N_4407,N_4433);
or U4558 (N_4558,N_4263,N_4260);
nand U4559 (N_4559,N_4467,N_4436);
nand U4560 (N_4560,N_4448,N_4401);
nand U4561 (N_4561,N_4418,N_4390);
nor U4562 (N_4562,N_4306,N_4296);
or U4563 (N_4563,N_4293,N_4372);
nand U4564 (N_4564,N_4480,N_4308);
xor U4565 (N_4565,N_4315,N_4332);
nor U4566 (N_4566,N_4321,N_4324);
and U4567 (N_4567,N_4434,N_4261);
nand U4568 (N_4568,N_4469,N_4317);
or U4569 (N_4569,N_4227,N_4251);
nand U4570 (N_4570,N_4476,N_4441);
or U4571 (N_4571,N_4409,N_4297);
and U4572 (N_4572,N_4368,N_4205);
or U4573 (N_4573,N_4430,N_4279);
and U4574 (N_4574,N_4213,N_4255);
or U4575 (N_4575,N_4413,N_4242);
nor U4576 (N_4576,N_4222,N_4303);
and U4577 (N_4577,N_4453,N_4257);
or U4578 (N_4578,N_4336,N_4464);
nor U4579 (N_4579,N_4240,N_4385);
nand U4580 (N_4580,N_4456,N_4402);
nor U4581 (N_4581,N_4289,N_4265);
and U4582 (N_4582,N_4284,N_4206);
and U4583 (N_4583,N_4281,N_4202);
and U4584 (N_4584,N_4217,N_4208);
nand U4585 (N_4585,N_4431,N_4323);
and U4586 (N_4586,N_4399,N_4310);
or U4587 (N_4587,N_4277,N_4460);
or U4588 (N_4588,N_4488,N_4273);
and U4589 (N_4589,N_4382,N_4427);
and U4590 (N_4590,N_4267,N_4244);
nor U4591 (N_4591,N_4258,N_4295);
nand U4592 (N_4592,N_4423,N_4466);
nand U4593 (N_4593,N_4337,N_4254);
xor U4594 (N_4594,N_4364,N_4450);
and U4595 (N_4595,N_4400,N_4499);
xor U4596 (N_4596,N_4313,N_4238);
xnor U4597 (N_4597,N_4475,N_4463);
nor U4598 (N_4598,N_4328,N_4340);
and U4599 (N_4599,N_4403,N_4420);
nor U4600 (N_4600,N_4435,N_4241);
nand U4601 (N_4601,N_4465,N_4357);
nand U4602 (N_4602,N_4358,N_4288);
nand U4603 (N_4603,N_4339,N_4455);
xnor U4604 (N_4604,N_4387,N_4496);
nand U4605 (N_4605,N_4212,N_4394);
nand U4606 (N_4606,N_4253,N_4348);
or U4607 (N_4607,N_4395,N_4285);
nor U4608 (N_4608,N_4471,N_4419);
and U4609 (N_4609,N_4373,N_4301);
and U4610 (N_4610,N_4389,N_4397);
or U4611 (N_4611,N_4377,N_4353);
or U4612 (N_4612,N_4416,N_4369);
nand U4613 (N_4613,N_4249,N_4305);
or U4614 (N_4614,N_4216,N_4200);
nand U4615 (N_4615,N_4331,N_4388);
nand U4616 (N_4616,N_4329,N_4495);
nor U4617 (N_4617,N_4298,N_4334);
nand U4618 (N_4618,N_4294,N_4291);
nor U4619 (N_4619,N_4243,N_4384);
and U4620 (N_4620,N_4485,N_4366);
nand U4621 (N_4621,N_4203,N_4454);
nand U4622 (N_4622,N_4319,N_4274);
xnor U4623 (N_4623,N_4343,N_4226);
nor U4624 (N_4624,N_4327,N_4474);
nand U4625 (N_4625,N_4437,N_4478);
nand U4626 (N_4626,N_4230,N_4493);
and U4627 (N_4627,N_4351,N_4404);
or U4628 (N_4628,N_4338,N_4307);
nand U4629 (N_4629,N_4370,N_4245);
or U4630 (N_4630,N_4231,N_4451);
nor U4631 (N_4631,N_4320,N_4349);
and U4632 (N_4632,N_4444,N_4311);
and U4633 (N_4633,N_4354,N_4484);
and U4634 (N_4634,N_4410,N_4256);
and U4635 (N_4635,N_4367,N_4270);
and U4636 (N_4636,N_4425,N_4220);
or U4637 (N_4637,N_4224,N_4232);
or U4638 (N_4638,N_4219,N_4378);
nand U4639 (N_4639,N_4462,N_4429);
xnor U4640 (N_4640,N_4300,N_4211);
nand U4641 (N_4641,N_4376,N_4459);
nand U4642 (N_4642,N_4215,N_4405);
or U4643 (N_4643,N_4398,N_4417);
nand U4644 (N_4644,N_4309,N_4236);
and U4645 (N_4645,N_4371,N_4452);
nand U4646 (N_4646,N_4221,N_4228);
xor U4647 (N_4647,N_4415,N_4282);
or U4648 (N_4648,N_4259,N_4494);
and U4649 (N_4649,N_4408,N_4438);
and U4650 (N_4650,N_4411,N_4397);
and U4651 (N_4651,N_4487,N_4296);
nor U4652 (N_4652,N_4306,N_4236);
nand U4653 (N_4653,N_4214,N_4320);
nor U4654 (N_4654,N_4492,N_4422);
and U4655 (N_4655,N_4407,N_4305);
nor U4656 (N_4656,N_4476,N_4384);
nor U4657 (N_4657,N_4392,N_4200);
nand U4658 (N_4658,N_4450,N_4435);
nor U4659 (N_4659,N_4394,N_4312);
nor U4660 (N_4660,N_4265,N_4232);
nor U4661 (N_4661,N_4474,N_4200);
nand U4662 (N_4662,N_4403,N_4276);
xor U4663 (N_4663,N_4229,N_4455);
or U4664 (N_4664,N_4290,N_4308);
or U4665 (N_4665,N_4397,N_4450);
xnor U4666 (N_4666,N_4431,N_4232);
or U4667 (N_4667,N_4409,N_4271);
or U4668 (N_4668,N_4250,N_4234);
xor U4669 (N_4669,N_4259,N_4264);
nor U4670 (N_4670,N_4368,N_4232);
nand U4671 (N_4671,N_4373,N_4303);
nor U4672 (N_4672,N_4439,N_4322);
nor U4673 (N_4673,N_4401,N_4302);
nand U4674 (N_4674,N_4225,N_4461);
or U4675 (N_4675,N_4432,N_4469);
nor U4676 (N_4676,N_4232,N_4303);
nor U4677 (N_4677,N_4425,N_4446);
or U4678 (N_4678,N_4432,N_4279);
and U4679 (N_4679,N_4415,N_4431);
or U4680 (N_4680,N_4235,N_4482);
and U4681 (N_4681,N_4205,N_4415);
or U4682 (N_4682,N_4426,N_4435);
nor U4683 (N_4683,N_4497,N_4327);
nor U4684 (N_4684,N_4318,N_4244);
or U4685 (N_4685,N_4295,N_4388);
and U4686 (N_4686,N_4473,N_4267);
nor U4687 (N_4687,N_4431,N_4311);
xor U4688 (N_4688,N_4476,N_4424);
or U4689 (N_4689,N_4401,N_4471);
or U4690 (N_4690,N_4271,N_4317);
nor U4691 (N_4691,N_4260,N_4353);
nand U4692 (N_4692,N_4301,N_4310);
and U4693 (N_4693,N_4422,N_4344);
or U4694 (N_4694,N_4268,N_4426);
or U4695 (N_4695,N_4207,N_4428);
and U4696 (N_4696,N_4202,N_4413);
and U4697 (N_4697,N_4320,N_4246);
and U4698 (N_4698,N_4240,N_4344);
xnor U4699 (N_4699,N_4213,N_4405);
and U4700 (N_4700,N_4431,N_4348);
xnor U4701 (N_4701,N_4240,N_4387);
nor U4702 (N_4702,N_4228,N_4354);
nand U4703 (N_4703,N_4286,N_4430);
xor U4704 (N_4704,N_4270,N_4325);
and U4705 (N_4705,N_4455,N_4371);
nor U4706 (N_4706,N_4251,N_4278);
xnor U4707 (N_4707,N_4431,N_4401);
or U4708 (N_4708,N_4330,N_4243);
xor U4709 (N_4709,N_4210,N_4393);
xor U4710 (N_4710,N_4495,N_4478);
nand U4711 (N_4711,N_4486,N_4461);
xnor U4712 (N_4712,N_4326,N_4462);
and U4713 (N_4713,N_4307,N_4228);
nor U4714 (N_4714,N_4247,N_4348);
and U4715 (N_4715,N_4338,N_4410);
or U4716 (N_4716,N_4345,N_4300);
and U4717 (N_4717,N_4272,N_4201);
nand U4718 (N_4718,N_4241,N_4282);
nor U4719 (N_4719,N_4420,N_4230);
or U4720 (N_4720,N_4364,N_4354);
xnor U4721 (N_4721,N_4318,N_4248);
or U4722 (N_4722,N_4318,N_4276);
xnor U4723 (N_4723,N_4273,N_4449);
nor U4724 (N_4724,N_4419,N_4434);
and U4725 (N_4725,N_4371,N_4226);
xnor U4726 (N_4726,N_4387,N_4264);
xnor U4727 (N_4727,N_4211,N_4369);
nor U4728 (N_4728,N_4471,N_4392);
nand U4729 (N_4729,N_4358,N_4316);
xnor U4730 (N_4730,N_4267,N_4443);
or U4731 (N_4731,N_4416,N_4403);
and U4732 (N_4732,N_4368,N_4403);
xnor U4733 (N_4733,N_4405,N_4283);
nor U4734 (N_4734,N_4275,N_4232);
nor U4735 (N_4735,N_4204,N_4251);
or U4736 (N_4736,N_4441,N_4380);
and U4737 (N_4737,N_4210,N_4399);
xnor U4738 (N_4738,N_4367,N_4322);
and U4739 (N_4739,N_4469,N_4232);
and U4740 (N_4740,N_4255,N_4216);
xnor U4741 (N_4741,N_4314,N_4243);
xnor U4742 (N_4742,N_4313,N_4325);
and U4743 (N_4743,N_4355,N_4387);
xnor U4744 (N_4744,N_4326,N_4415);
and U4745 (N_4745,N_4463,N_4222);
nor U4746 (N_4746,N_4341,N_4323);
or U4747 (N_4747,N_4495,N_4355);
and U4748 (N_4748,N_4373,N_4274);
or U4749 (N_4749,N_4480,N_4420);
or U4750 (N_4750,N_4331,N_4311);
or U4751 (N_4751,N_4305,N_4481);
nor U4752 (N_4752,N_4213,N_4229);
or U4753 (N_4753,N_4217,N_4476);
or U4754 (N_4754,N_4478,N_4344);
nor U4755 (N_4755,N_4243,N_4225);
nand U4756 (N_4756,N_4347,N_4245);
and U4757 (N_4757,N_4407,N_4467);
xnor U4758 (N_4758,N_4494,N_4305);
or U4759 (N_4759,N_4225,N_4394);
xnor U4760 (N_4760,N_4337,N_4470);
or U4761 (N_4761,N_4364,N_4391);
or U4762 (N_4762,N_4233,N_4296);
nor U4763 (N_4763,N_4250,N_4296);
or U4764 (N_4764,N_4218,N_4324);
nand U4765 (N_4765,N_4231,N_4422);
or U4766 (N_4766,N_4493,N_4382);
or U4767 (N_4767,N_4407,N_4488);
nand U4768 (N_4768,N_4361,N_4395);
nor U4769 (N_4769,N_4419,N_4265);
nor U4770 (N_4770,N_4473,N_4239);
or U4771 (N_4771,N_4277,N_4267);
nand U4772 (N_4772,N_4274,N_4207);
nor U4773 (N_4773,N_4376,N_4413);
nor U4774 (N_4774,N_4223,N_4335);
nor U4775 (N_4775,N_4396,N_4356);
nor U4776 (N_4776,N_4362,N_4420);
nand U4777 (N_4777,N_4272,N_4489);
and U4778 (N_4778,N_4445,N_4410);
nor U4779 (N_4779,N_4295,N_4458);
or U4780 (N_4780,N_4247,N_4290);
or U4781 (N_4781,N_4385,N_4367);
or U4782 (N_4782,N_4218,N_4468);
nand U4783 (N_4783,N_4320,N_4449);
nor U4784 (N_4784,N_4282,N_4435);
xor U4785 (N_4785,N_4207,N_4291);
and U4786 (N_4786,N_4292,N_4241);
nand U4787 (N_4787,N_4269,N_4403);
nor U4788 (N_4788,N_4230,N_4211);
nand U4789 (N_4789,N_4476,N_4313);
nor U4790 (N_4790,N_4495,N_4308);
or U4791 (N_4791,N_4240,N_4282);
or U4792 (N_4792,N_4441,N_4334);
xnor U4793 (N_4793,N_4449,N_4258);
and U4794 (N_4794,N_4264,N_4407);
nand U4795 (N_4795,N_4315,N_4308);
xor U4796 (N_4796,N_4341,N_4485);
or U4797 (N_4797,N_4246,N_4235);
nor U4798 (N_4798,N_4493,N_4462);
and U4799 (N_4799,N_4340,N_4429);
nor U4800 (N_4800,N_4604,N_4609);
nor U4801 (N_4801,N_4676,N_4788);
xnor U4802 (N_4802,N_4597,N_4738);
xor U4803 (N_4803,N_4530,N_4741);
nand U4804 (N_4804,N_4764,N_4717);
and U4805 (N_4805,N_4590,N_4672);
nand U4806 (N_4806,N_4678,N_4591);
or U4807 (N_4807,N_4752,N_4508);
and U4808 (N_4808,N_4596,N_4760);
or U4809 (N_4809,N_4625,N_4601);
nor U4810 (N_4810,N_4681,N_4722);
nand U4811 (N_4811,N_4538,N_4794);
and U4812 (N_4812,N_4598,N_4734);
xor U4813 (N_4813,N_4773,N_4744);
nand U4814 (N_4814,N_4595,N_4682);
and U4815 (N_4815,N_4616,N_4635);
nand U4816 (N_4816,N_4665,N_4579);
xor U4817 (N_4817,N_4655,N_4535);
nand U4818 (N_4818,N_4661,N_4732);
and U4819 (N_4819,N_4570,N_4526);
nand U4820 (N_4820,N_4748,N_4549);
xnor U4821 (N_4821,N_4627,N_4725);
nand U4822 (N_4822,N_4736,N_4755);
and U4823 (N_4823,N_4565,N_4675);
or U4824 (N_4824,N_4664,N_4726);
xnor U4825 (N_4825,N_4602,N_4552);
and U4826 (N_4826,N_4689,N_4548);
or U4827 (N_4827,N_4782,N_4556);
xor U4828 (N_4828,N_4520,N_4600);
nand U4829 (N_4829,N_4612,N_4550);
xor U4830 (N_4830,N_4668,N_4592);
xnor U4831 (N_4831,N_4614,N_4659);
nor U4832 (N_4832,N_4667,N_4537);
and U4833 (N_4833,N_4685,N_4706);
nand U4834 (N_4834,N_4518,N_4687);
xnor U4835 (N_4835,N_4624,N_4541);
nand U4836 (N_4836,N_4503,N_4674);
xor U4837 (N_4837,N_4688,N_4567);
nor U4838 (N_4838,N_4576,N_4638);
or U4839 (N_4839,N_4683,N_4765);
nand U4840 (N_4840,N_4720,N_4553);
nor U4841 (N_4841,N_4514,N_4581);
nand U4842 (N_4842,N_4573,N_4756);
nand U4843 (N_4843,N_4785,N_4630);
nor U4844 (N_4844,N_4691,N_4619);
nor U4845 (N_4845,N_4733,N_4636);
nand U4846 (N_4846,N_4771,N_4588);
nor U4847 (N_4847,N_4761,N_4634);
xor U4848 (N_4848,N_4730,N_4658);
nand U4849 (N_4849,N_4589,N_4790);
nand U4850 (N_4850,N_4620,N_4737);
xor U4851 (N_4851,N_4613,N_4531);
xnor U4852 (N_4852,N_4580,N_4729);
xnor U4853 (N_4853,N_4714,N_4781);
nand U4854 (N_4854,N_4505,N_4702);
nand U4855 (N_4855,N_4631,N_4750);
xnor U4856 (N_4856,N_4695,N_4787);
xnor U4857 (N_4857,N_4544,N_4608);
and U4858 (N_4858,N_4585,N_4704);
xor U4859 (N_4859,N_4651,N_4605);
xor U4860 (N_4860,N_4677,N_4763);
and U4861 (N_4861,N_4519,N_4746);
nand U4862 (N_4862,N_4504,N_4719);
xnor U4863 (N_4863,N_4663,N_4566);
or U4864 (N_4864,N_4536,N_4522);
and U4865 (N_4865,N_4529,N_4648);
or U4866 (N_4866,N_4618,N_4701);
xor U4867 (N_4867,N_4660,N_4629);
and U4868 (N_4868,N_4769,N_4789);
and U4869 (N_4869,N_4521,N_4586);
or U4870 (N_4870,N_4693,N_4517);
nor U4871 (N_4871,N_4759,N_4735);
and U4872 (N_4872,N_4543,N_4515);
and U4873 (N_4873,N_4742,N_4791);
or U4874 (N_4874,N_4540,N_4584);
nor U4875 (N_4875,N_4692,N_4690);
nand U4876 (N_4876,N_4798,N_4757);
or U4877 (N_4877,N_4745,N_4793);
or U4878 (N_4878,N_4749,N_4780);
nor U4879 (N_4879,N_4545,N_4577);
nor U4880 (N_4880,N_4777,N_4502);
or U4881 (N_4881,N_4709,N_4539);
xor U4882 (N_4882,N_4562,N_4568);
or U4883 (N_4883,N_4778,N_4774);
xor U4884 (N_4884,N_4557,N_4650);
xnor U4885 (N_4885,N_4751,N_4772);
and U4886 (N_4886,N_4571,N_4770);
and U4887 (N_4887,N_4705,N_4640);
nand U4888 (N_4888,N_4569,N_4560);
or U4889 (N_4889,N_4637,N_4776);
or U4890 (N_4890,N_4723,N_4645);
xor U4891 (N_4891,N_4684,N_4786);
and U4892 (N_4892,N_4574,N_4766);
or U4893 (N_4893,N_4647,N_4572);
and U4894 (N_4894,N_4739,N_4662);
xnor U4895 (N_4895,N_4554,N_4657);
and U4896 (N_4896,N_4641,N_4680);
xnor U4897 (N_4897,N_4784,N_4547);
xnor U4898 (N_4898,N_4783,N_4628);
and U4899 (N_4899,N_4673,N_4740);
and U4900 (N_4900,N_4666,N_4697);
and U4901 (N_4901,N_4716,N_4599);
and U4902 (N_4902,N_4626,N_4564);
xnor U4903 (N_4903,N_4587,N_4563);
and U4904 (N_4904,N_4575,N_4699);
nor U4905 (N_4905,N_4644,N_4525);
or U4906 (N_4906,N_4533,N_4649);
nand U4907 (N_4907,N_4527,N_4617);
or U4908 (N_4908,N_4747,N_4679);
nand U4909 (N_4909,N_4712,N_4606);
nor U4910 (N_4910,N_4724,N_4524);
nor U4911 (N_4911,N_4696,N_4561);
and U4912 (N_4912,N_4646,N_4713);
or U4913 (N_4913,N_4583,N_4642);
nor U4914 (N_4914,N_4795,N_4743);
nor U4915 (N_4915,N_4500,N_4758);
xnor U4916 (N_4916,N_4727,N_4779);
and U4917 (N_4917,N_4669,N_4506);
nand U4918 (N_4918,N_4753,N_4542);
nor U4919 (N_4919,N_4728,N_4534);
or U4920 (N_4920,N_4797,N_4710);
and U4921 (N_4921,N_4513,N_4512);
or U4922 (N_4922,N_4754,N_4721);
and U4923 (N_4923,N_4551,N_4523);
nor U4924 (N_4924,N_4643,N_4528);
or U4925 (N_4925,N_4703,N_4593);
or U4926 (N_4926,N_4615,N_4610);
and U4927 (N_4927,N_4623,N_4656);
xor U4928 (N_4928,N_4698,N_4559);
nand U4929 (N_4929,N_4510,N_4555);
nor U4930 (N_4930,N_4731,N_4509);
or U4931 (N_4931,N_4532,N_4670);
xor U4932 (N_4932,N_4546,N_4708);
and U4933 (N_4933,N_4632,N_4767);
nor U4934 (N_4934,N_4622,N_4653);
nand U4935 (N_4935,N_4582,N_4711);
nand U4936 (N_4936,N_4511,N_4700);
and U4937 (N_4937,N_4611,N_4792);
nand U4938 (N_4938,N_4715,N_4558);
and U4939 (N_4939,N_4707,N_4594);
xnor U4940 (N_4940,N_4507,N_4768);
and U4941 (N_4941,N_4686,N_4799);
nor U4942 (N_4942,N_4578,N_4652);
xor U4943 (N_4943,N_4796,N_4516);
and U4944 (N_4944,N_4654,N_4603);
xor U4945 (N_4945,N_4501,N_4775);
and U4946 (N_4946,N_4633,N_4621);
nor U4947 (N_4947,N_4671,N_4607);
nor U4948 (N_4948,N_4718,N_4762);
and U4949 (N_4949,N_4694,N_4639);
nor U4950 (N_4950,N_4540,N_4521);
and U4951 (N_4951,N_4644,N_4778);
nand U4952 (N_4952,N_4675,N_4635);
xnor U4953 (N_4953,N_4598,N_4585);
nand U4954 (N_4954,N_4765,N_4546);
or U4955 (N_4955,N_4729,N_4523);
nand U4956 (N_4956,N_4596,N_4609);
or U4957 (N_4957,N_4692,N_4605);
and U4958 (N_4958,N_4541,N_4792);
nand U4959 (N_4959,N_4550,N_4703);
or U4960 (N_4960,N_4583,N_4664);
xor U4961 (N_4961,N_4584,N_4598);
nor U4962 (N_4962,N_4680,N_4619);
xnor U4963 (N_4963,N_4678,N_4550);
nand U4964 (N_4964,N_4526,N_4562);
nor U4965 (N_4965,N_4587,N_4659);
nand U4966 (N_4966,N_4742,N_4653);
nor U4967 (N_4967,N_4613,N_4748);
and U4968 (N_4968,N_4662,N_4632);
xnor U4969 (N_4969,N_4766,N_4657);
or U4970 (N_4970,N_4774,N_4568);
or U4971 (N_4971,N_4660,N_4608);
nand U4972 (N_4972,N_4566,N_4657);
or U4973 (N_4973,N_4625,N_4741);
or U4974 (N_4974,N_4615,N_4589);
nor U4975 (N_4975,N_4668,N_4646);
or U4976 (N_4976,N_4741,N_4560);
nand U4977 (N_4977,N_4514,N_4717);
and U4978 (N_4978,N_4564,N_4701);
xor U4979 (N_4979,N_4663,N_4767);
and U4980 (N_4980,N_4500,N_4511);
xnor U4981 (N_4981,N_4635,N_4582);
and U4982 (N_4982,N_4680,N_4546);
or U4983 (N_4983,N_4679,N_4507);
or U4984 (N_4984,N_4707,N_4564);
xor U4985 (N_4985,N_4795,N_4684);
nand U4986 (N_4986,N_4660,N_4757);
nor U4987 (N_4987,N_4777,N_4539);
or U4988 (N_4988,N_4620,N_4669);
and U4989 (N_4989,N_4717,N_4796);
nand U4990 (N_4990,N_4762,N_4501);
and U4991 (N_4991,N_4593,N_4717);
xnor U4992 (N_4992,N_4529,N_4551);
or U4993 (N_4993,N_4752,N_4551);
nand U4994 (N_4994,N_4773,N_4511);
nor U4995 (N_4995,N_4701,N_4608);
nand U4996 (N_4996,N_4645,N_4602);
xor U4997 (N_4997,N_4724,N_4695);
and U4998 (N_4998,N_4631,N_4625);
and U4999 (N_4999,N_4568,N_4782);
nand U5000 (N_5000,N_4728,N_4783);
and U5001 (N_5001,N_4745,N_4587);
nor U5002 (N_5002,N_4748,N_4633);
xnor U5003 (N_5003,N_4501,N_4693);
or U5004 (N_5004,N_4745,N_4705);
xnor U5005 (N_5005,N_4721,N_4620);
or U5006 (N_5006,N_4706,N_4767);
or U5007 (N_5007,N_4605,N_4762);
nand U5008 (N_5008,N_4614,N_4549);
and U5009 (N_5009,N_4515,N_4722);
xnor U5010 (N_5010,N_4537,N_4621);
xor U5011 (N_5011,N_4790,N_4516);
xor U5012 (N_5012,N_4517,N_4726);
xnor U5013 (N_5013,N_4667,N_4601);
and U5014 (N_5014,N_4770,N_4747);
nand U5015 (N_5015,N_4507,N_4589);
and U5016 (N_5016,N_4500,N_4705);
nand U5017 (N_5017,N_4675,N_4711);
and U5018 (N_5018,N_4602,N_4615);
xor U5019 (N_5019,N_4777,N_4697);
nor U5020 (N_5020,N_4751,N_4501);
xnor U5021 (N_5021,N_4707,N_4516);
nand U5022 (N_5022,N_4770,N_4638);
and U5023 (N_5023,N_4683,N_4637);
nand U5024 (N_5024,N_4772,N_4585);
and U5025 (N_5025,N_4584,N_4697);
nand U5026 (N_5026,N_4748,N_4664);
and U5027 (N_5027,N_4684,N_4747);
or U5028 (N_5028,N_4609,N_4689);
or U5029 (N_5029,N_4563,N_4626);
or U5030 (N_5030,N_4706,N_4728);
or U5031 (N_5031,N_4593,N_4701);
xor U5032 (N_5032,N_4547,N_4551);
nor U5033 (N_5033,N_4506,N_4794);
or U5034 (N_5034,N_4626,N_4733);
xor U5035 (N_5035,N_4589,N_4799);
and U5036 (N_5036,N_4713,N_4635);
nand U5037 (N_5037,N_4772,N_4701);
nand U5038 (N_5038,N_4572,N_4775);
or U5039 (N_5039,N_4698,N_4762);
or U5040 (N_5040,N_4646,N_4660);
xnor U5041 (N_5041,N_4625,N_4795);
nor U5042 (N_5042,N_4606,N_4552);
nand U5043 (N_5043,N_4770,N_4705);
nand U5044 (N_5044,N_4764,N_4546);
and U5045 (N_5045,N_4693,N_4557);
or U5046 (N_5046,N_4672,N_4696);
nor U5047 (N_5047,N_4781,N_4661);
and U5048 (N_5048,N_4724,N_4681);
nand U5049 (N_5049,N_4662,N_4581);
and U5050 (N_5050,N_4633,N_4575);
nand U5051 (N_5051,N_4567,N_4618);
or U5052 (N_5052,N_4503,N_4616);
xnor U5053 (N_5053,N_4691,N_4542);
nand U5054 (N_5054,N_4685,N_4650);
or U5055 (N_5055,N_4735,N_4631);
nor U5056 (N_5056,N_4770,N_4550);
xor U5057 (N_5057,N_4508,N_4694);
or U5058 (N_5058,N_4786,N_4655);
nand U5059 (N_5059,N_4668,N_4528);
nand U5060 (N_5060,N_4521,N_4652);
xnor U5061 (N_5061,N_4661,N_4791);
or U5062 (N_5062,N_4574,N_4688);
nor U5063 (N_5063,N_4594,N_4733);
or U5064 (N_5064,N_4777,N_4642);
nand U5065 (N_5065,N_4557,N_4531);
nand U5066 (N_5066,N_4566,N_4775);
and U5067 (N_5067,N_4688,N_4663);
and U5068 (N_5068,N_4508,N_4629);
or U5069 (N_5069,N_4690,N_4590);
nand U5070 (N_5070,N_4728,N_4526);
nand U5071 (N_5071,N_4549,N_4632);
or U5072 (N_5072,N_4577,N_4610);
nand U5073 (N_5073,N_4608,N_4783);
and U5074 (N_5074,N_4755,N_4695);
nor U5075 (N_5075,N_4531,N_4510);
and U5076 (N_5076,N_4785,N_4698);
nand U5077 (N_5077,N_4795,N_4580);
and U5078 (N_5078,N_4525,N_4719);
and U5079 (N_5079,N_4558,N_4681);
nand U5080 (N_5080,N_4642,N_4762);
xnor U5081 (N_5081,N_4663,N_4694);
xor U5082 (N_5082,N_4674,N_4767);
and U5083 (N_5083,N_4793,N_4653);
nor U5084 (N_5084,N_4540,N_4535);
xnor U5085 (N_5085,N_4555,N_4620);
xor U5086 (N_5086,N_4711,N_4551);
nand U5087 (N_5087,N_4694,N_4792);
nand U5088 (N_5088,N_4506,N_4501);
nor U5089 (N_5089,N_4575,N_4766);
nor U5090 (N_5090,N_4556,N_4792);
xnor U5091 (N_5091,N_4680,N_4588);
xnor U5092 (N_5092,N_4682,N_4675);
xor U5093 (N_5093,N_4568,N_4652);
nand U5094 (N_5094,N_4725,N_4746);
or U5095 (N_5095,N_4740,N_4765);
xnor U5096 (N_5096,N_4520,N_4521);
and U5097 (N_5097,N_4588,N_4746);
and U5098 (N_5098,N_4755,N_4562);
and U5099 (N_5099,N_4618,N_4642);
or U5100 (N_5100,N_4913,N_5072);
xnor U5101 (N_5101,N_4817,N_4821);
xnor U5102 (N_5102,N_4865,N_4868);
and U5103 (N_5103,N_5097,N_4867);
nand U5104 (N_5104,N_4833,N_4877);
nand U5105 (N_5105,N_5064,N_4823);
and U5106 (N_5106,N_4925,N_4828);
or U5107 (N_5107,N_4825,N_4826);
nor U5108 (N_5108,N_4858,N_5018);
or U5109 (N_5109,N_5080,N_5050);
xor U5110 (N_5110,N_4895,N_4937);
and U5111 (N_5111,N_5059,N_4830);
or U5112 (N_5112,N_4844,N_4950);
nor U5113 (N_5113,N_4919,N_4939);
or U5114 (N_5114,N_5076,N_5051);
nor U5115 (N_5115,N_4840,N_5061);
or U5116 (N_5116,N_4879,N_4874);
or U5117 (N_5117,N_4882,N_4853);
nand U5118 (N_5118,N_4816,N_5078);
and U5119 (N_5119,N_4995,N_5007);
and U5120 (N_5120,N_4902,N_4850);
nor U5121 (N_5121,N_4878,N_5054);
xnor U5122 (N_5122,N_5005,N_4806);
nand U5123 (N_5123,N_4930,N_5069);
nand U5124 (N_5124,N_5026,N_5092);
xnor U5125 (N_5125,N_4966,N_4888);
or U5126 (N_5126,N_4953,N_4860);
nor U5127 (N_5127,N_5011,N_4904);
nor U5128 (N_5128,N_5058,N_4979);
or U5129 (N_5129,N_4864,N_4936);
and U5130 (N_5130,N_5074,N_4892);
or U5131 (N_5131,N_5006,N_5017);
xor U5132 (N_5132,N_4933,N_5053);
or U5133 (N_5133,N_4987,N_5019);
nor U5134 (N_5134,N_5042,N_4898);
nor U5135 (N_5135,N_4805,N_4845);
nand U5136 (N_5136,N_4851,N_4985);
nor U5137 (N_5137,N_4958,N_4869);
nand U5138 (N_5138,N_5099,N_5056);
or U5139 (N_5139,N_5002,N_4996);
nor U5140 (N_5140,N_4848,N_4899);
xor U5141 (N_5141,N_5000,N_4949);
nand U5142 (N_5142,N_4822,N_5014);
xor U5143 (N_5143,N_5063,N_4908);
xnor U5144 (N_5144,N_4955,N_4992);
nor U5145 (N_5145,N_4970,N_4809);
xor U5146 (N_5146,N_4928,N_5015);
and U5147 (N_5147,N_4810,N_4839);
xor U5148 (N_5148,N_4986,N_4814);
xor U5149 (N_5149,N_4800,N_4991);
xor U5150 (N_5150,N_5062,N_4903);
nor U5151 (N_5151,N_4884,N_4829);
or U5152 (N_5152,N_4808,N_5093);
and U5153 (N_5153,N_5031,N_5020);
nor U5154 (N_5154,N_5044,N_4948);
nand U5155 (N_5155,N_5037,N_4931);
nand U5156 (N_5156,N_5030,N_5048);
or U5157 (N_5157,N_4889,N_4818);
and U5158 (N_5158,N_4857,N_5024);
xor U5159 (N_5159,N_4852,N_4961);
nand U5160 (N_5160,N_5055,N_5088);
and U5161 (N_5161,N_4922,N_5090);
or U5162 (N_5162,N_5089,N_4960);
or U5163 (N_5163,N_4965,N_4956);
or U5164 (N_5164,N_4897,N_5095);
nand U5165 (N_5165,N_4990,N_4849);
nor U5166 (N_5166,N_5032,N_5039);
and U5167 (N_5167,N_4998,N_4976);
and U5168 (N_5168,N_5028,N_5004);
xnor U5169 (N_5169,N_4896,N_5091);
and U5170 (N_5170,N_5035,N_4886);
nand U5171 (N_5171,N_4862,N_4945);
nand U5172 (N_5172,N_4926,N_4876);
or U5173 (N_5173,N_4954,N_5052);
and U5174 (N_5174,N_5013,N_4883);
and U5175 (N_5175,N_4835,N_4807);
or U5176 (N_5176,N_4837,N_5094);
xor U5177 (N_5177,N_4927,N_5084);
and U5178 (N_5178,N_4841,N_5082);
nand U5179 (N_5179,N_4880,N_5077);
and U5180 (N_5180,N_4964,N_4803);
or U5181 (N_5181,N_4951,N_4934);
nor U5182 (N_5182,N_5071,N_4832);
or U5183 (N_5183,N_4804,N_5085);
or U5184 (N_5184,N_4952,N_4866);
or U5185 (N_5185,N_4891,N_4893);
xnor U5186 (N_5186,N_4963,N_5043);
xnor U5187 (N_5187,N_5070,N_4983);
xnor U5188 (N_5188,N_5083,N_4988);
nand U5189 (N_5189,N_4915,N_4859);
or U5190 (N_5190,N_4957,N_5045);
or U5191 (N_5191,N_4982,N_5096);
xnor U5192 (N_5192,N_5047,N_4967);
xor U5193 (N_5193,N_4906,N_4812);
xnor U5194 (N_5194,N_4900,N_5029);
or U5195 (N_5195,N_5023,N_4885);
xnor U5196 (N_5196,N_4855,N_5009);
xor U5197 (N_5197,N_4975,N_4811);
or U5198 (N_5198,N_4997,N_4907);
or U5199 (N_5199,N_4929,N_5016);
nor U5200 (N_5200,N_4834,N_4843);
nand U5201 (N_5201,N_5086,N_4881);
or U5202 (N_5202,N_5060,N_4973);
nor U5203 (N_5203,N_4815,N_4972);
nor U5204 (N_5204,N_4971,N_4871);
and U5205 (N_5205,N_4924,N_4827);
and U5206 (N_5206,N_4872,N_4984);
and U5207 (N_5207,N_4890,N_4916);
xor U5208 (N_5208,N_4905,N_4819);
or U5209 (N_5209,N_5025,N_4935);
nand U5210 (N_5210,N_4912,N_4863);
nor U5211 (N_5211,N_4989,N_5012);
or U5212 (N_5212,N_4846,N_4873);
nor U5213 (N_5213,N_5001,N_4968);
or U5214 (N_5214,N_5087,N_4917);
nand U5215 (N_5215,N_4969,N_4959);
and U5216 (N_5216,N_4831,N_5081);
and U5217 (N_5217,N_4847,N_4801);
xor U5218 (N_5218,N_4894,N_5003);
nor U5219 (N_5219,N_5010,N_4947);
and U5220 (N_5220,N_4910,N_4946);
nand U5221 (N_5221,N_5038,N_4824);
or U5222 (N_5222,N_4836,N_4923);
or U5223 (N_5223,N_4861,N_4820);
and U5224 (N_5224,N_4920,N_4901);
xnor U5225 (N_5225,N_4942,N_4978);
nand U5226 (N_5226,N_5040,N_4842);
and U5227 (N_5227,N_5008,N_4999);
nand U5228 (N_5228,N_4943,N_5098);
nor U5229 (N_5229,N_5066,N_4944);
or U5230 (N_5230,N_4932,N_4856);
xnor U5231 (N_5231,N_5021,N_4918);
nor U5232 (N_5232,N_5046,N_4941);
or U5233 (N_5233,N_4909,N_4981);
nor U5234 (N_5234,N_5034,N_4854);
and U5235 (N_5235,N_4993,N_5075);
nor U5236 (N_5236,N_4887,N_5079);
nand U5237 (N_5237,N_5036,N_5022);
or U5238 (N_5238,N_4938,N_5057);
nand U5239 (N_5239,N_4914,N_5027);
nand U5240 (N_5240,N_4994,N_4875);
and U5241 (N_5241,N_4977,N_4838);
nor U5242 (N_5242,N_5041,N_5065);
xnor U5243 (N_5243,N_5033,N_4921);
nor U5244 (N_5244,N_5073,N_4870);
nand U5245 (N_5245,N_4813,N_4980);
nand U5246 (N_5246,N_5068,N_5067);
xor U5247 (N_5247,N_4911,N_4940);
nor U5248 (N_5248,N_4802,N_4974);
or U5249 (N_5249,N_5049,N_4962);
xor U5250 (N_5250,N_4960,N_4958);
or U5251 (N_5251,N_4864,N_4986);
nor U5252 (N_5252,N_5048,N_4927);
nand U5253 (N_5253,N_5009,N_4965);
nor U5254 (N_5254,N_5046,N_5061);
xnor U5255 (N_5255,N_5090,N_4940);
nor U5256 (N_5256,N_4947,N_4878);
nor U5257 (N_5257,N_5034,N_4893);
nand U5258 (N_5258,N_4906,N_4966);
nand U5259 (N_5259,N_4865,N_5085);
or U5260 (N_5260,N_4877,N_5076);
nand U5261 (N_5261,N_5068,N_4877);
xnor U5262 (N_5262,N_5085,N_4923);
nand U5263 (N_5263,N_5068,N_5007);
nand U5264 (N_5264,N_5038,N_5094);
and U5265 (N_5265,N_5061,N_4829);
or U5266 (N_5266,N_5079,N_4949);
and U5267 (N_5267,N_4962,N_5078);
xor U5268 (N_5268,N_5015,N_4962);
xor U5269 (N_5269,N_4900,N_4848);
or U5270 (N_5270,N_5053,N_4809);
xor U5271 (N_5271,N_4839,N_4963);
xnor U5272 (N_5272,N_4862,N_4896);
xor U5273 (N_5273,N_4994,N_4972);
nand U5274 (N_5274,N_4876,N_5062);
and U5275 (N_5275,N_5000,N_5011);
nor U5276 (N_5276,N_5007,N_4860);
xor U5277 (N_5277,N_5045,N_4993);
nor U5278 (N_5278,N_4984,N_5050);
or U5279 (N_5279,N_5002,N_5069);
and U5280 (N_5280,N_5040,N_4944);
nand U5281 (N_5281,N_4982,N_4839);
nand U5282 (N_5282,N_4808,N_4834);
nand U5283 (N_5283,N_4806,N_4901);
xnor U5284 (N_5284,N_4985,N_5041);
nor U5285 (N_5285,N_5027,N_5094);
nand U5286 (N_5286,N_4844,N_4859);
nand U5287 (N_5287,N_4896,N_4892);
and U5288 (N_5288,N_4933,N_4816);
xor U5289 (N_5289,N_4899,N_4929);
and U5290 (N_5290,N_4851,N_4905);
xnor U5291 (N_5291,N_4964,N_5035);
xnor U5292 (N_5292,N_5062,N_4850);
nor U5293 (N_5293,N_4971,N_4824);
nand U5294 (N_5294,N_5004,N_4989);
nand U5295 (N_5295,N_4918,N_4922);
xor U5296 (N_5296,N_4886,N_4864);
or U5297 (N_5297,N_4828,N_5058);
xnor U5298 (N_5298,N_4850,N_4973);
nand U5299 (N_5299,N_5083,N_4989);
or U5300 (N_5300,N_4976,N_4813);
and U5301 (N_5301,N_5073,N_5007);
and U5302 (N_5302,N_5043,N_4955);
xor U5303 (N_5303,N_4991,N_4972);
and U5304 (N_5304,N_5002,N_4858);
and U5305 (N_5305,N_4915,N_5006);
xnor U5306 (N_5306,N_4855,N_4852);
nand U5307 (N_5307,N_5075,N_4888);
nor U5308 (N_5308,N_5066,N_4978);
or U5309 (N_5309,N_4996,N_4858);
xnor U5310 (N_5310,N_4897,N_5000);
or U5311 (N_5311,N_4934,N_5079);
nand U5312 (N_5312,N_4808,N_5068);
xnor U5313 (N_5313,N_4935,N_4940);
xnor U5314 (N_5314,N_5023,N_4818);
or U5315 (N_5315,N_4913,N_5061);
xnor U5316 (N_5316,N_5053,N_5027);
nand U5317 (N_5317,N_5008,N_4815);
nor U5318 (N_5318,N_5099,N_4829);
nand U5319 (N_5319,N_4914,N_4845);
nand U5320 (N_5320,N_4859,N_5078);
xor U5321 (N_5321,N_4847,N_5003);
xor U5322 (N_5322,N_4998,N_4871);
nor U5323 (N_5323,N_5013,N_4882);
nor U5324 (N_5324,N_5077,N_4937);
and U5325 (N_5325,N_4894,N_4895);
nand U5326 (N_5326,N_4967,N_4947);
nor U5327 (N_5327,N_4892,N_5049);
nor U5328 (N_5328,N_5096,N_4841);
nor U5329 (N_5329,N_4841,N_5020);
or U5330 (N_5330,N_4836,N_4846);
xor U5331 (N_5331,N_4968,N_4880);
nand U5332 (N_5332,N_4925,N_4930);
and U5333 (N_5333,N_4814,N_5020);
or U5334 (N_5334,N_4932,N_4931);
nand U5335 (N_5335,N_5082,N_4921);
or U5336 (N_5336,N_4999,N_4985);
xnor U5337 (N_5337,N_4986,N_4956);
and U5338 (N_5338,N_4852,N_4896);
or U5339 (N_5339,N_5030,N_4934);
nand U5340 (N_5340,N_4901,N_5084);
and U5341 (N_5341,N_5098,N_4897);
nand U5342 (N_5342,N_4982,N_4842);
nand U5343 (N_5343,N_5086,N_5070);
and U5344 (N_5344,N_4926,N_5060);
xor U5345 (N_5345,N_5014,N_4891);
nand U5346 (N_5346,N_5063,N_5019);
and U5347 (N_5347,N_4805,N_4920);
xor U5348 (N_5348,N_4960,N_4892);
nand U5349 (N_5349,N_4879,N_4965);
or U5350 (N_5350,N_5046,N_5057);
nand U5351 (N_5351,N_4967,N_4826);
nand U5352 (N_5352,N_5069,N_4837);
nor U5353 (N_5353,N_4933,N_4898);
and U5354 (N_5354,N_4857,N_4855);
xor U5355 (N_5355,N_4936,N_4803);
nand U5356 (N_5356,N_5002,N_5065);
or U5357 (N_5357,N_4831,N_5051);
xnor U5358 (N_5358,N_4921,N_5004);
xor U5359 (N_5359,N_4857,N_5005);
xnor U5360 (N_5360,N_4945,N_5045);
nand U5361 (N_5361,N_4903,N_4928);
or U5362 (N_5362,N_4882,N_5034);
and U5363 (N_5363,N_4973,N_4982);
nand U5364 (N_5364,N_4842,N_4836);
nor U5365 (N_5365,N_4819,N_5074);
nand U5366 (N_5366,N_5005,N_5051);
xor U5367 (N_5367,N_4824,N_5054);
nand U5368 (N_5368,N_4920,N_4999);
xnor U5369 (N_5369,N_4901,N_4869);
xor U5370 (N_5370,N_4895,N_5071);
nand U5371 (N_5371,N_4851,N_5076);
nor U5372 (N_5372,N_4809,N_5035);
nand U5373 (N_5373,N_4992,N_5082);
nand U5374 (N_5374,N_4902,N_4977);
or U5375 (N_5375,N_4811,N_4900);
xnor U5376 (N_5376,N_4978,N_4859);
and U5377 (N_5377,N_4836,N_4820);
and U5378 (N_5378,N_4994,N_5032);
nor U5379 (N_5379,N_4834,N_4897);
nand U5380 (N_5380,N_4845,N_4864);
nand U5381 (N_5381,N_4895,N_5034);
xnor U5382 (N_5382,N_4935,N_5089);
or U5383 (N_5383,N_4894,N_4972);
or U5384 (N_5384,N_4837,N_4957);
and U5385 (N_5385,N_5048,N_4996);
nand U5386 (N_5386,N_4938,N_4961);
nand U5387 (N_5387,N_5060,N_5083);
or U5388 (N_5388,N_4860,N_4838);
xnor U5389 (N_5389,N_5023,N_4803);
nand U5390 (N_5390,N_5077,N_4889);
and U5391 (N_5391,N_4846,N_4947);
xnor U5392 (N_5392,N_4951,N_4920);
and U5393 (N_5393,N_4967,N_5054);
nor U5394 (N_5394,N_4934,N_4940);
nor U5395 (N_5395,N_4848,N_5080);
and U5396 (N_5396,N_4904,N_5031);
and U5397 (N_5397,N_4875,N_4827);
and U5398 (N_5398,N_4800,N_5097);
nand U5399 (N_5399,N_4845,N_5060);
or U5400 (N_5400,N_5264,N_5222);
nand U5401 (N_5401,N_5331,N_5263);
xor U5402 (N_5402,N_5187,N_5307);
nand U5403 (N_5403,N_5253,N_5346);
and U5404 (N_5404,N_5124,N_5109);
or U5405 (N_5405,N_5230,N_5195);
or U5406 (N_5406,N_5143,N_5317);
or U5407 (N_5407,N_5146,N_5373);
and U5408 (N_5408,N_5265,N_5114);
nor U5409 (N_5409,N_5375,N_5254);
xor U5410 (N_5410,N_5341,N_5304);
nand U5411 (N_5411,N_5178,N_5393);
or U5412 (N_5412,N_5386,N_5241);
nor U5413 (N_5413,N_5173,N_5395);
nor U5414 (N_5414,N_5259,N_5295);
nand U5415 (N_5415,N_5193,N_5340);
nor U5416 (N_5416,N_5299,N_5394);
or U5417 (N_5417,N_5199,N_5358);
or U5418 (N_5418,N_5314,N_5203);
nor U5419 (N_5419,N_5336,N_5140);
or U5420 (N_5420,N_5252,N_5158);
nor U5421 (N_5421,N_5359,N_5343);
nor U5422 (N_5422,N_5248,N_5305);
xor U5423 (N_5423,N_5360,N_5311);
nand U5424 (N_5424,N_5162,N_5169);
nor U5425 (N_5425,N_5213,N_5107);
or U5426 (N_5426,N_5227,N_5272);
nor U5427 (N_5427,N_5185,N_5344);
or U5428 (N_5428,N_5152,N_5354);
and U5429 (N_5429,N_5338,N_5167);
xnor U5430 (N_5430,N_5155,N_5244);
and U5431 (N_5431,N_5112,N_5121);
nor U5432 (N_5432,N_5128,N_5371);
nand U5433 (N_5433,N_5353,N_5151);
and U5434 (N_5434,N_5115,N_5239);
xor U5435 (N_5435,N_5132,N_5113);
nor U5436 (N_5436,N_5216,N_5291);
nor U5437 (N_5437,N_5147,N_5172);
nand U5438 (N_5438,N_5176,N_5306);
or U5439 (N_5439,N_5233,N_5348);
or U5440 (N_5440,N_5110,N_5282);
xnor U5441 (N_5441,N_5149,N_5260);
nand U5442 (N_5442,N_5231,N_5181);
nand U5443 (N_5443,N_5196,N_5315);
or U5444 (N_5444,N_5397,N_5246);
nor U5445 (N_5445,N_5104,N_5283);
or U5446 (N_5446,N_5268,N_5322);
and U5447 (N_5447,N_5335,N_5356);
and U5448 (N_5448,N_5165,N_5330);
and U5449 (N_5449,N_5277,N_5321);
nor U5450 (N_5450,N_5370,N_5301);
nand U5451 (N_5451,N_5191,N_5234);
xor U5452 (N_5452,N_5302,N_5364);
xor U5453 (N_5453,N_5355,N_5214);
nor U5454 (N_5454,N_5163,N_5164);
nor U5455 (N_5455,N_5154,N_5221);
nor U5456 (N_5456,N_5137,N_5200);
nand U5457 (N_5457,N_5292,N_5174);
nor U5458 (N_5458,N_5201,N_5224);
xnor U5459 (N_5459,N_5278,N_5189);
nand U5460 (N_5460,N_5148,N_5261);
or U5461 (N_5461,N_5379,N_5120);
nor U5462 (N_5462,N_5168,N_5150);
nor U5463 (N_5463,N_5286,N_5284);
xnor U5464 (N_5464,N_5103,N_5131);
or U5465 (N_5465,N_5318,N_5220);
nor U5466 (N_5466,N_5288,N_5345);
or U5467 (N_5467,N_5217,N_5285);
xor U5468 (N_5468,N_5387,N_5141);
or U5469 (N_5469,N_5366,N_5390);
nor U5470 (N_5470,N_5209,N_5339);
and U5471 (N_5471,N_5334,N_5328);
and U5472 (N_5472,N_5320,N_5376);
and U5473 (N_5473,N_5352,N_5365);
nor U5474 (N_5474,N_5157,N_5287);
nor U5475 (N_5475,N_5275,N_5122);
or U5476 (N_5476,N_5136,N_5350);
and U5477 (N_5477,N_5229,N_5382);
and U5478 (N_5478,N_5271,N_5197);
and U5479 (N_5479,N_5251,N_5333);
nor U5480 (N_5480,N_5236,N_5215);
and U5481 (N_5481,N_5349,N_5342);
nor U5482 (N_5482,N_5347,N_5367);
and U5483 (N_5483,N_5398,N_5326);
nand U5484 (N_5484,N_5383,N_5374);
or U5485 (N_5485,N_5381,N_5294);
and U5486 (N_5486,N_5255,N_5232);
or U5487 (N_5487,N_5243,N_5257);
and U5488 (N_5488,N_5198,N_5276);
nand U5489 (N_5489,N_5378,N_5184);
or U5490 (N_5490,N_5388,N_5205);
and U5491 (N_5491,N_5361,N_5202);
nand U5492 (N_5492,N_5139,N_5175);
nand U5493 (N_5493,N_5138,N_5281);
xnor U5494 (N_5494,N_5385,N_5130);
and U5495 (N_5495,N_5293,N_5310);
and U5496 (N_5496,N_5377,N_5324);
or U5497 (N_5497,N_5303,N_5300);
nor U5498 (N_5498,N_5270,N_5368);
xnor U5499 (N_5499,N_5240,N_5183);
nand U5500 (N_5500,N_5119,N_5204);
or U5501 (N_5501,N_5237,N_5190);
and U5502 (N_5502,N_5225,N_5123);
or U5503 (N_5503,N_5223,N_5384);
nand U5504 (N_5504,N_5242,N_5127);
xor U5505 (N_5505,N_5289,N_5380);
or U5506 (N_5506,N_5273,N_5134);
nand U5507 (N_5507,N_5266,N_5212);
nor U5508 (N_5508,N_5135,N_5129);
xnor U5509 (N_5509,N_5262,N_5101);
nand U5510 (N_5510,N_5274,N_5156);
xnor U5511 (N_5511,N_5207,N_5177);
and U5512 (N_5512,N_5161,N_5125);
xor U5513 (N_5513,N_5194,N_5111);
or U5514 (N_5514,N_5226,N_5160);
nor U5515 (N_5515,N_5362,N_5267);
xor U5516 (N_5516,N_5313,N_5116);
xnor U5517 (N_5517,N_5323,N_5250);
xor U5518 (N_5518,N_5247,N_5279);
xor U5519 (N_5519,N_5389,N_5392);
or U5520 (N_5520,N_5357,N_5351);
nand U5521 (N_5521,N_5218,N_5297);
or U5522 (N_5522,N_5298,N_5396);
and U5523 (N_5523,N_5308,N_5179);
xnor U5524 (N_5524,N_5186,N_5171);
nand U5525 (N_5525,N_5312,N_5144);
or U5526 (N_5526,N_5249,N_5159);
and U5527 (N_5527,N_5399,N_5327);
nor U5528 (N_5528,N_5296,N_5211);
xor U5529 (N_5529,N_5258,N_5145);
nor U5530 (N_5530,N_5170,N_5108);
nor U5531 (N_5531,N_5238,N_5126);
and U5532 (N_5532,N_5269,N_5208);
or U5533 (N_5533,N_5228,N_5142);
nor U5534 (N_5534,N_5100,N_5309);
or U5535 (N_5535,N_5235,N_5337);
and U5536 (N_5536,N_5369,N_5256);
nor U5537 (N_5537,N_5188,N_5219);
or U5538 (N_5538,N_5118,N_5105);
and U5539 (N_5539,N_5153,N_5329);
nand U5540 (N_5540,N_5182,N_5280);
nand U5541 (N_5541,N_5206,N_5316);
nand U5542 (N_5542,N_5180,N_5245);
and U5543 (N_5543,N_5332,N_5391);
nor U5544 (N_5544,N_5372,N_5166);
xnor U5545 (N_5545,N_5133,N_5325);
nand U5546 (N_5546,N_5106,N_5192);
nor U5547 (N_5547,N_5290,N_5210);
xnor U5548 (N_5548,N_5102,N_5363);
xor U5549 (N_5549,N_5319,N_5117);
xnor U5550 (N_5550,N_5165,N_5393);
xor U5551 (N_5551,N_5375,N_5285);
nor U5552 (N_5552,N_5281,N_5342);
and U5553 (N_5553,N_5346,N_5173);
nand U5554 (N_5554,N_5220,N_5180);
nand U5555 (N_5555,N_5267,N_5205);
or U5556 (N_5556,N_5364,N_5162);
or U5557 (N_5557,N_5180,N_5164);
or U5558 (N_5558,N_5313,N_5336);
and U5559 (N_5559,N_5322,N_5246);
or U5560 (N_5560,N_5119,N_5360);
xor U5561 (N_5561,N_5328,N_5189);
xor U5562 (N_5562,N_5335,N_5296);
nand U5563 (N_5563,N_5303,N_5337);
xnor U5564 (N_5564,N_5377,N_5397);
or U5565 (N_5565,N_5342,N_5242);
and U5566 (N_5566,N_5211,N_5300);
and U5567 (N_5567,N_5132,N_5122);
nor U5568 (N_5568,N_5142,N_5229);
or U5569 (N_5569,N_5335,N_5122);
and U5570 (N_5570,N_5176,N_5224);
xnor U5571 (N_5571,N_5270,N_5308);
or U5572 (N_5572,N_5246,N_5118);
or U5573 (N_5573,N_5263,N_5329);
nand U5574 (N_5574,N_5311,N_5397);
and U5575 (N_5575,N_5273,N_5226);
or U5576 (N_5576,N_5306,N_5267);
nor U5577 (N_5577,N_5277,N_5293);
or U5578 (N_5578,N_5381,N_5326);
nor U5579 (N_5579,N_5233,N_5240);
nor U5580 (N_5580,N_5173,N_5274);
nand U5581 (N_5581,N_5228,N_5319);
xor U5582 (N_5582,N_5230,N_5190);
and U5583 (N_5583,N_5331,N_5252);
xor U5584 (N_5584,N_5155,N_5361);
nor U5585 (N_5585,N_5207,N_5171);
nor U5586 (N_5586,N_5305,N_5167);
nor U5587 (N_5587,N_5292,N_5191);
nor U5588 (N_5588,N_5346,N_5352);
nor U5589 (N_5589,N_5399,N_5342);
nand U5590 (N_5590,N_5337,N_5142);
xnor U5591 (N_5591,N_5268,N_5155);
nand U5592 (N_5592,N_5224,N_5347);
xnor U5593 (N_5593,N_5108,N_5218);
and U5594 (N_5594,N_5123,N_5326);
or U5595 (N_5595,N_5165,N_5120);
nand U5596 (N_5596,N_5209,N_5259);
or U5597 (N_5597,N_5207,N_5120);
xnor U5598 (N_5598,N_5179,N_5238);
and U5599 (N_5599,N_5278,N_5184);
nor U5600 (N_5600,N_5283,N_5164);
and U5601 (N_5601,N_5257,N_5165);
and U5602 (N_5602,N_5323,N_5277);
xnor U5603 (N_5603,N_5255,N_5368);
or U5604 (N_5604,N_5204,N_5222);
xor U5605 (N_5605,N_5284,N_5126);
or U5606 (N_5606,N_5115,N_5117);
nor U5607 (N_5607,N_5348,N_5329);
or U5608 (N_5608,N_5396,N_5336);
nand U5609 (N_5609,N_5342,N_5248);
xor U5610 (N_5610,N_5215,N_5155);
or U5611 (N_5611,N_5302,N_5166);
nor U5612 (N_5612,N_5324,N_5333);
nand U5613 (N_5613,N_5360,N_5138);
or U5614 (N_5614,N_5130,N_5268);
and U5615 (N_5615,N_5231,N_5376);
and U5616 (N_5616,N_5342,N_5204);
and U5617 (N_5617,N_5123,N_5250);
nor U5618 (N_5618,N_5254,N_5341);
or U5619 (N_5619,N_5229,N_5366);
or U5620 (N_5620,N_5232,N_5247);
nand U5621 (N_5621,N_5100,N_5352);
and U5622 (N_5622,N_5290,N_5180);
or U5623 (N_5623,N_5343,N_5147);
and U5624 (N_5624,N_5154,N_5361);
or U5625 (N_5625,N_5341,N_5371);
and U5626 (N_5626,N_5380,N_5165);
xnor U5627 (N_5627,N_5305,N_5125);
or U5628 (N_5628,N_5265,N_5325);
xor U5629 (N_5629,N_5307,N_5184);
and U5630 (N_5630,N_5103,N_5341);
xor U5631 (N_5631,N_5144,N_5191);
xnor U5632 (N_5632,N_5390,N_5198);
or U5633 (N_5633,N_5142,N_5280);
xnor U5634 (N_5634,N_5372,N_5321);
nor U5635 (N_5635,N_5225,N_5281);
and U5636 (N_5636,N_5180,N_5386);
nand U5637 (N_5637,N_5235,N_5372);
or U5638 (N_5638,N_5383,N_5343);
and U5639 (N_5639,N_5182,N_5383);
nor U5640 (N_5640,N_5113,N_5281);
or U5641 (N_5641,N_5291,N_5166);
nand U5642 (N_5642,N_5123,N_5301);
and U5643 (N_5643,N_5294,N_5292);
nor U5644 (N_5644,N_5191,N_5210);
and U5645 (N_5645,N_5105,N_5141);
nor U5646 (N_5646,N_5274,N_5397);
nor U5647 (N_5647,N_5335,N_5281);
and U5648 (N_5648,N_5209,N_5366);
nor U5649 (N_5649,N_5284,N_5399);
nand U5650 (N_5650,N_5367,N_5173);
and U5651 (N_5651,N_5178,N_5191);
or U5652 (N_5652,N_5365,N_5380);
xor U5653 (N_5653,N_5257,N_5353);
and U5654 (N_5654,N_5260,N_5175);
and U5655 (N_5655,N_5252,N_5288);
nand U5656 (N_5656,N_5134,N_5370);
or U5657 (N_5657,N_5149,N_5209);
nor U5658 (N_5658,N_5285,N_5167);
nor U5659 (N_5659,N_5337,N_5271);
xor U5660 (N_5660,N_5199,N_5336);
nor U5661 (N_5661,N_5147,N_5188);
xnor U5662 (N_5662,N_5194,N_5160);
xnor U5663 (N_5663,N_5232,N_5158);
and U5664 (N_5664,N_5156,N_5172);
nand U5665 (N_5665,N_5168,N_5189);
nor U5666 (N_5666,N_5181,N_5127);
nor U5667 (N_5667,N_5399,N_5319);
or U5668 (N_5668,N_5239,N_5103);
or U5669 (N_5669,N_5180,N_5155);
nor U5670 (N_5670,N_5112,N_5357);
and U5671 (N_5671,N_5127,N_5172);
nor U5672 (N_5672,N_5385,N_5398);
and U5673 (N_5673,N_5130,N_5365);
or U5674 (N_5674,N_5313,N_5176);
or U5675 (N_5675,N_5228,N_5371);
or U5676 (N_5676,N_5163,N_5298);
nor U5677 (N_5677,N_5267,N_5229);
and U5678 (N_5678,N_5251,N_5292);
or U5679 (N_5679,N_5216,N_5365);
nand U5680 (N_5680,N_5297,N_5193);
xor U5681 (N_5681,N_5240,N_5104);
nand U5682 (N_5682,N_5376,N_5238);
nand U5683 (N_5683,N_5327,N_5235);
and U5684 (N_5684,N_5273,N_5252);
or U5685 (N_5685,N_5147,N_5165);
or U5686 (N_5686,N_5337,N_5260);
nor U5687 (N_5687,N_5275,N_5308);
xnor U5688 (N_5688,N_5348,N_5307);
xor U5689 (N_5689,N_5257,N_5118);
and U5690 (N_5690,N_5212,N_5278);
and U5691 (N_5691,N_5210,N_5119);
and U5692 (N_5692,N_5315,N_5110);
nor U5693 (N_5693,N_5300,N_5395);
and U5694 (N_5694,N_5135,N_5211);
and U5695 (N_5695,N_5334,N_5245);
and U5696 (N_5696,N_5353,N_5277);
nor U5697 (N_5697,N_5257,N_5308);
nand U5698 (N_5698,N_5246,N_5161);
or U5699 (N_5699,N_5350,N_5369);
xnor U5700 (N_5700,N_5465,N_5581);
or U5701 (N_5701,N_5513,N_5567);
nand U5702 (N_5702,N_5616,N_5437);
and U5703 (N_5703,N_5529,N_5556);
xor U5704 (N_5704,N_5541,N_5420);
or U5705 (N_5705,N_5464,N_5456);
nor U5706 (N_5706,N_5589,N_5532);
nand U5707 (N_5707,N_5565,N_5501);
xor U5708 (N_5708,N_5442,N_5525);
nand U5709 (N_5709,N_5404,N_5463);
or U5710 (N_5710,N_5696,N_5553);
and U5711 (N_5711,N_5461,N_5623);
xnor U5712 (N_5712,N_5425,N_5438);
nand U5713 (N_5713,N_5684,N_5618);
and U5714 (N_5714,N_5524,N_5514);
nor U5715 (N_5715,N_5445,N_5542);
xor U5716 (N_5716,N_5605,N_5620);
nand U5717 (N_5717,N_5680,N_5676);
nand U5718 (N_5718,N_5625,N_5570);
nand U5719 (N_5719,N_5689,N_5466);
xnor U5720 (N_5720,N_5478,N_5564);
xnor U5721 (N_5721,N_5666,N_5652);
or U5722 (N_5722,N_5587,N_5537);
xor U5723 (N_5723,N_5606,N_5672);
or U5724 (N_5724,N_5447,N_5613);
nor U5725 (N_5725,N_5462,N_5667);
nand U5726 (N_5726,N_5495,N_5577);
nor U5727 (N_5727,N_5477,N_5610);
nand U5728 (N_5728,N_5687,N_5450);
or U5729 (N_5729,N_5413,N_5663);
and U5730 (N_5730,N_5576,N_5422);
xnor U5731 (N_5731,N_5431,N_5628);
nor U5732 (N_5732,N_5662,N_5569);
nand U5733 (N_5733,N_5551,N_5458);
or U5734 (N_5734,N_5402,N_5615);
xnor U5735 (N_5735,N_5455,N_5481);
nor U5736 (N_5736,N_5506,N_5448);
xnor U5737 (N_5737,N_5492,N_5600);
or U5738 (N_5738,N_5518,N_5545);
nand U5739 (N_5739,N_5609,N_5428);
or U5740 (N_5740,N_5530,N_5601);
nand U5741 (N_5741,N_5683,N_5490);
and U5742 (N_5742,N_5408,N_5583);
xnor U5743 (N_5743,N_5639,N_5657);
xnor U5744 (N_5744,N_5690,N_5632);
nand U5745 (N_5745,N_5608,N_5472);
nor U5746 (N_5746,N_5627,N_5649);
and U5747 (N_5747,N_5670,N_5441);
and U5748 (N_5748,N_5641,N_5651);
or U5749 (N_5749,N_5512,N_5555);
nand U5750 (N_5750,N_5497,N_5411);
xor U5751 (N_5751,N_5434,N_5642);
nor U5752 (N_5752,N_5538,N_5650);
and U5753 (N_5753,N_5645,N_5526);
or U5754 (N_5754,N_5602,N_5635);
nor U5755 (N_5755,N_5661,N_5559);
nand U5756 (N_5756,N_5451,N_5473);
and U5757 (N_5757,N_5469,N_5500);
and U5758 (N_5758,N_5671,N_5636);
and U5759 (N_5759,N_5579,N_5519);
or U5760 (N_5760,N_5622,N_5659);
nor U5761 (N_5761,N_5479,N_5584);
or U5762 (N_5762,N_5489,N_5691);
xnor U5763 (N_5763,N_5646,N_5417);
or U5764 (N_5764,N_5427,N_5452);
nand U5765 (N_5765,N_5654,N_5669);
xnor U5766 (N_5766,N_5644,N_5440);
or U5767 (N_5767,N_5673,N_5590);
xnor U5768 (N_5768,N_5695,N_5488);
or U5769 (N_5769,N_5603,N_5682);
xnor U5770 (N_5770,N_5423,N_5502);
nor U5771 (N_5771,N_5460,N_5634);
nor U5772 (N_5772,N_5499,N_5629);
nor U5773 (N_5773,N_5648,N_5647);
nand U5774 (N_5774,N_5424,N_5694);
or U5775 (N_5775,N_5543,N_5637);
nand U5776 (N_5776,N_5638,N_5435);
or U5777 (N_5777,N_5444,N_5475);
or U5778 (N_5778,N_5697,N_5561);
xnor U5779 (N_5779,N_5407,N_5494);
nor U5780 (N_5780,N_5505,N_5558);
xnor U5781 (N_5781,N_5621,N_5516);
nand U5782 (N_5782,N_5643,N_5496);
or U5783 (N_5783,N_5548,N_5546);
or U5784 (N_5784,N_5493,N_5515);
and U5785 (N_5785,N_5485,N_5523);
and U5786 (N_5786,N_5547,N_5520);
or U5787 (N_5787,N_5534,N_5582);
xnor U5788 (N_5788,N_5467,N_5550);
nor U5789 (N_5789,N_5585,N_5560);
xnor U5790 (N_5790,N_5409,N_5531);
nor U5791 (N_5791,N_5674,N_5401);
nor U5792 (N_5792,N_5403,N_5656);
nand U5793 (N_5793,N_5658,N_5594);
nor U5794 (N_5794,N_5517,N_5429);
or U5795 (N_5795,N_5535,N_5509);
or U5796 (N_5796,N_5470,N_5592);
and U5797 (N_5797,N_5677,N_5688);
or U5798 (N_5798,N_5498,N_5454);
and U5799 (N_5799,N_5508,N_5595);
nand U5800 (N_5800,N_5624,N_5563);
or U5801 (N_5801,N_5571,N_5686);
and U5802 (N_5802,N_5487,N_5588);
xor U5803 (N_5803,N_5678,N_5491);
nand U5804 (N_5804,N_5416,N_5522);
or U5805 (N_5805,N_5503,N_5544);
nor U5806 (N_5806,N_5459,N_5614);
xnor U5807 (N_5807,N_5471,N_5568);
or U5808 (N_5808,N_5631,N_5527);
nor U5809 (N_5809,N_5685,N_5557);
nand U5810 (N_5810,N_5457,N_5415);
nor U5811 (N_5811,N_5607,N_5449);
xnor U5812 (N_5812,N_5681,N_5655);
and U5813 (N_5813,N_5410,N_5630);
and U5814 (N_5814,N_5679,N_5439);
nor U5815 (N_5815,N_5599,N_5507);
or U5816 (N_5816,N_5528,N_5436);
nand U5817 (N_5817,N_5633,N_5574);
or U5818 (N_5818,N_5675,N_5421);
xor U5819 (N_5819,N_5640,N_5664);
or U5820 (N_5820,N_5693,N_5562);
xor U5821 (N_5821,N_5510,N_5430);
xor U5822 (N_5822,N_5698,N_5486);
or U5823 (N_5823,N_5586,N_5483);
or U5824 (N_5824,N_5626,N_5540);
or U5825 (N_5825,N_5419,N_5412);
nand U5826 (N_5826,N_5554,N_5406);
xor U5827 (N_5827,N_5453,N_5539);
or U5828 (N_5828,N_5414,N_5611);
and U5829 (N_5829,N_5468,N_5699);
xnor U5830 (N_5830,N_5433,N_5432);
nand U5831 (N_5831,N_5580,N_5405);
nor U5832 (N_5832,N_5533,N_5446);
xnor U5833 (N_5833,N_5426,N_5443);
nor U5834 (N_5834,N_5572,N_5480);
nand U5835 (N_5835,N_5549,N_5578);
xnor U5836 (N_5836,N_5474,N_5653);
xor U5837 (N_5837,N_5692,N_5660);
xnor U5838 (N_5838,N_5552,N_5511);
or U5839 (N_5839,N_5619,N_5484);
xnor U5840 (N_5840,N_5575,N_5504);
and U5841 (N_5841,N_5598,N_5617);
nor U5842 (N_5842,N_5597,N_5591);
xor U5843 (N_5843,N_5536,N_5400);
nand U5844 (N_5844,N_5482,N_5596);
and U5845 (N_5845,N_5668,N_5573);
xnor U5846 (N_5846,N_5521,N_5593);
and U5847 (N_5847,N_5418,N_5604);
nor U5848 (N_5848,N_5612,N_5566);
nand U5849 (N_5849,N_5665,N_5476);
and U5850 (N_5850,N_5608,N_5522);
nor U5851 (N_5851,N_5480,N_5656);
nand U5852 (N_5852,N_5636,N_5456);
or U5853 (N_5853,N_5402,N_5577);
or U5854 (N_5854,N_5449,N_5408);
xor U5855 (N_5855,N_5446,N_5648);
xor U5856 (N_5856,N_5663,N_5423);
and U5857 (N_5857,N_5686,N_5612);
nand U5858 (N_5858,N_5529,N_5411);
nand U5859 (N_5859,N_5401,N_5516);
or U5860 (N_5860,N_5581,N_5538);
xor U5861 (N_5861,N_5623,N_5452);
nor U5862 (N_5862,N_5564,N_5645);
nor U5863 (N_5863,N_5544,N_5559);
nand U5864 (N_5864,N_5496,N_5550);
or U5865 (N_5865,N_5438,N_5504);
xnor U5866 (N_5866,N_5666,N_5438);
or U5867 (N_5867,N_5524,N_5490);
nand U5868 (N_5868,N_5679,N_5600);
nand U5869 (N_5869,N_5601,N_5634);
or U5870 (N_5870,N_5688,N_5494);
nand U5871 (N_5871,N_5597,N_5494);
nand U5872 (N_5872,N_5671,N_5622);
xnor U5873 (N_5873,N_5647,N_5592);
nand U5874 (N_5874,N_5405,N_5526);
and U5875 (N_5875,N_5523,N_5554);
and U5876 (N_5876,N_5547,N_5601);
nor U5877 (N_5877,N_5695,N_5688);
nand U5878 (N_5878,N_5576,N_5491);
nand U5879 (N_5879,N_5405,N_5623);
or U5880 (N_5880,N_5443,N_5430);
nor U5881 (N_5881,N_5615,N_5613);
or U5882 (N_5882,N_5696,N_5453);
nor U5883 (N_5883,N_5647,N_5695);
and U5884 (N_5884,N_5422,N_5605);
or U5885 (N_5885,N_5512,N_5493);
xnor U5886 (N_5886,N_5696,N_5502);
nand U5887 (N_5887,N_5650,N_5685);
nand U5888 (N_5888,N_5456,N_5591);
xor U5889 (N_5889,N_5489,N_5459);
and U5890 (N_5890,N_5476,N_5526);
nand U5891 (N_5891,N_5668,N_5583);
nand U5892 (N_5892,N_5428,N_5433);
nand U5893 (N_5893,N_5554,N_5513);
nor U5894 (N_5894,N_5647,N_5604);
nor U5895 (N_5895,N_5419,N_5474);
and U5896 (N_5896,N_5565,N_5416);
and U5897 (N_5897,N_5491,N_5663);
nor U5898 (N_5898,N_5402,N_5654);
and U5899 (N_5899,N_5458,N_5429);
xnor U5900 (N_5900,N_5463,N_5416);
nand U5901 (N_5901,N_5494,N_5498);
or U5902 (N_5902,N_5608,N_5525);
and U5903 (N_5903,N_5569,N_5658);
and U5904 (N_5904,N_5540,N_5543);
nand U5905 (N_5905,N_5405,N_5630);
nand U5906 (N_5906,N_5697,N_5446);
nand U5907 (N_5907,N_5412,N_5437);
nor U5908 (N_5908,N_5686,N_5660);
xnor U5909 (N_5909,N_5532,N_5581);
nor U5910 (N_5910,N_5568,N_5591);
or U5911 (N_5911,N_5566,N_5500);
or U5912 (N_5912,N_5452,N_5669);
and U5913 (N_5913,N_5685,N_5624);
or U5914 (N_5914,N_5616,N_5582);
nor U5915 (N_5915,N_5678,N_5508);
nand U5916 (N_5916,N_5433,N_5572);
or U5917 (N_5917,N_5521,N_5444);
nand U5918 (N_5918,N_5558,N_5431);
nor U5919 (N_5919,N_5655,N_5636);
nor U5920 (N_5920,N_5410,N_5488);
or U5921 (N_5921,N_5486,N_5608);
and U5922 (N_5922,N_5449,N_5578);
and U5923 (N_5923,N_5541,N_5484);
nand U5924 (N_5924,N_5591,N_5608);
and U5925 (N_5925,N_5536,N_5563);
and U5926 (N_5926,N_5411,N_5686);
nor U5927 (N_5927,N_5618,N_5622);
xor U5928 (N_5928,N_5575,N_5464);
nor U5929 (N_5929,N_5681,N_5528);
nor U5930 (N_5930,N_5543,N_5562);
xnor U5931 (N_5931,N_5406,N_5470);
xor U5932 (N_5932,N_5619,N_5687);
xor U5933 (N_5933,N_5568,N_5485);
nor U5934 (N_5934,N_5423,N_5414);
xnor U5935 (N_5935,N_5441,N_5437);
nand U5936 (N_5936,N_5536,N_5585);
xor U5937 (N_5937,N_5656,N_5477);
nand U5938 (N_5938,N_5513,N_5668);
or U5939 (N_5939,N_5678,N_5665);
nor U5940 (N_5940,N_5430,N_5650);
or U5941 (N_5941,N_5530,N_5520);
xnor U5942 (N_5942,N_5403,N_5569);
and U5943 (N_5943,N_5409,N_5556);
nor U5944 (N_5944,N_5539,N_5564);
nor U5945 (N_5945,N_5566,N_5531);
and U5946 (N_5946,N_5626,N_5444);
xnor U5947 (N_5947,N_5562,N_5457);
and U5948 (N_5948,N_5636,N_5496);
xor U5949 (N_5949,N_5623,N_5440);
nor U5950 (N_5950,N_5605,N_5563);
nor U5951 (N_5951,N_5690,N_5571);
or U5952 (N_5952,N_5481,N_5482);
and U5953 (N_5953,N_5435,N_5665);
and U5954 (N_5954,N_5561,N_5531);
xor U5955 (N_5955,N_5493,N_5606);
and U5956 (N_5956,N_5662,N_5673);
xor U5957 (N_5957,N_5549,N_5432);
xor U5958 (N_5958,N_5617,N_5498);
nor U5959 (N_5959,N_5548,N_5597);
or U5960 (N_5960,N_5637,N_5521);
xnor U5961 (N_5961,N_5587,N_5648);
xnor U5962 (N_5962,N_5685,N_5471);
and U5963 (N_5963,N_5610,N_5649);
nor U5964 (N_5964,N_5417,N_5633);
or U5965 (N_5965,N_5581,N_5647);
nor U5966 (N_5966,N_5659,N_5617);
nor U5967 (N_5967,N_5580,N_5619);
nor U5968 (N_5968,N_5644,N_5689);
xnor U5969 (N_5969,N_5459,N_5575);
xor U5970 (N_5970,N_5665,N_5426);
or U5971 (N_5971,N_5479,N_5581);
or U5972 (N_5972,N_5531,N_5417);
xor U5973 (N_5973,N_5598,N_5632);
and U5974 (N_5974,N_5514,N_5602);
nor U5975 (N_5975,N_5667,N_5623);
nor U5976 (N_5976,N_5457,N_5570);
or U5977 (N_5977,N_5499,N_5596);
nor U5978 (N_5978,N_5530,N_5671);
nand U5979 (N_5979,N_5624,N_5688);
xnor U5980 (N_5980,N_5622,N_5572);
nor U5981 (N_5981,N_5660,N_5609);
nand U5982 (N_5982,N_5598,N_5527);
or U5983 (N_5983,N_5493,N_5416);
and U5984 (N_5984,N_5568,N_5400);
or U5985 (N_5985,N_5603,N_5423);
xnor U5986 (N_5986,N_5489,N_5436);
nand U5987 (N_5987,N_5455,N_5484);
and U5988 (N_5988,N_5536,N_5592);
nor U5989 (N_5989,N_5552,N_5632);
nand U5990 (N_5990,N_5495,N_5580);
and U5991 (N_5991,N_5519,N_5447);
nand U5992 (N_5992,N_5468,N_5453);
nor U5993 (N_5993,N_5579,N_5567);
nand U5994 (N_5994,N_5539,N_5443);
xnor U5995 (N_5995,N_5697,N_5695);
nor U5996 (N_5996,N_5547,N_5483);
nor U5997 (N_5997,N_5462,N_5408);
xor U5998 (N_5998,N_5401,N_5437);
or U5999 (N_5999,N_5429,N_5537);
and U6000 (N_6000,N_5806,N_5829);
nor U6001 (N_6001,N_5793,N_5760);
nor U6002 (N_6002,N_5761,N_5933);
nor U6003 (N_6003,N_5876,N_5879);
or U6004 (N_6004,N_5759,N_5832);
or U6005 (N_6005,N_5769,N_5710);
nand U6006 (N_6006,N_5967,N_5947);
xor U6007 (N_6007,N_5797,N_5942);
xnor U6008 (N_6008,N_5800,N_5741);
nand U6009 (N_6009,N_5785,N_5786);
and U6010 (N_6010,N_5982,N_5843);
xnor U6011 (N_6011,N_5957,N_5972);
nor U6012 (N_6012,N_5828,N_5747);
xor U6013 (N_6013,N_5861,N_5929);
nand U6014 (N_6014,N_5787,N_5846);
xor U6015 (N_6015,N_5757,N_5810);
nor U6016 (N_6016,N_5824,N_5968);
nand U6017 (N_6017,N_5944,N_5714);
nor U6018 (N_6018,N_5854,N_5790);
nand U6019 (N_6019,N_5976,N_5808);
or U6020 (N_6020,N_5722,N_5858);
and U6021 (N_6021,N_5836,N_5921);
or U6022 (N_6022,N_5926,N_5880);
and U6023 (N_6023,N_5920,N_5905);
and U6024 (N_6024,N_5821,N_5857);
nor U6025 (N_6025,N_5903,N_5753);
nor U6026 (N_6026,N_5763,N_5937);
or U6027 (N_6027,N_5979,N_5706);
nor U6028 (N_6028,N_5814,N_5994);
xor U6029 (N_6029,N_5888,N_5866);
xor U6030 (N_6030,N_5954,N_5733);
or U6031 (N_6031,N_5740,N_5746);
nand U6032 (N_6032,N_5749,N_5711);
nor U6033 (N_6033,N_5923,N_5909);
nand U6034 (N_6034,N_5713,N_5735);
and U6035 (N_6035,N_5900,N_5889);
or U6036 (N_6036,N_5856,N_5984);
xor U6037 (N_6037,N_5703,N_5912);
xor U6038 (N_6038,N_5913,N_5701);
and U6039 (N_6039,N_5813,N_5772);
and U6040 (N_6040,N_5794,N_5766);
nand U6041 (N_6041,N_5958,N_5948);
and U6042 (N_6042,N_5974,N_5991);
and U6043 (N_6043,N_5989,N_5953);
nor U6044 (N_6044,N_5727,N_5988);
xor U6045 (N_6045,N_5840,N_5971);
and U6046 (N_6046,N_5748,N_5805);
nand U6047 (N_6047,N_5924,N_5744);
or U6048 (N_6048,N_5985,N_5737);
and U6049 (N_6049,N_5812,N_5964);
xor U6050 (N_6050,N_5938,N_5927);
and U6051 (N_6051,N_5844,N_5949);
nand U6052 (N_6052,N_5896,N_5914);
nand U6053 (N_6053,N_5922,N_5940);
and U6054 (N_6054,N_5743,N_5887);
nor U6055 (N_6055,N_5899,N_5742);
or U6056 (N_6056,N_5784,N_5853);
nor U6057 (N_6057,N_5980,N_5973);
xnor U6058 (N_6058,N_5878,N_5819);
or U6059 (N_6059,N_5754,N_5756);
nor U6060 (N_6060,N_5709,N_5762);
xnor U6061 (N_6061,N_5816,N_5868);
nor U6062 (N_6062,N_5702,N_5983);
nand U6063 (N_6063,N_5823,N_5936);
xor U6064 (N_6064,N_5897,N_5745);
or U6065 (N_6065,N_5841,N_5770);
or U6066 (N_6066,N_5849,N_5732);
nor U6067 (N_6067,N_5904,N_5919);
or U6068 (N_6068,N_5961,N_5943);
nor U6069 (N_6069,N_5783,N_5777);
xor U6070 (N_6070,N_5768,N_5998);
and U6071 (N_6071,N_5725,N_5700);
or U6072 (N_6072,N_5718,N_5864);
nor U6073 (N_6073,N_5717,N_5881);
and U6074 (N_6074,N_5867,N_5765);
and U6075 (N_6075,N_5822,N_5932);
xor U6076 (N_6076,N_5781,N_5885);
nor U6077 (N_6077,N_5789,N_5731);
nand U6078 (N_6078,N_5833,N_5811);
nand U6079 (N_6079,N_5815,N_5915);
nand U6080 (N_6080,N_5908,N_5935);
nor U6081 (N_6081,N_5893,N_5719);
and U6082 (N_6082,N_5870,N_5838);
nand U6083 (N_6083,N_5752,N_5995);
xor U6084 (N_6084,N_5736,N_5803);
or U6085 (N_6085,N_5895,N_5860);
xnor U6086 (N_6086,N_5946,N_5906);
or U6087 (N_6087,N_5848,N_5963);
nor U6088 (N_6088,N_5758,N_5898);
nand U6089 (N_6089,N_5877,N_5778);
or U6090 (N_6090,N_5862,N_5873);
xor U6091 (N_6091,N_5738,N_5807);
or U6092 (N_6092,N_5825,N_5891);
and U6093 (N_6093,N_5941,N_5997);
nor U6094 (N_6094,N_5950,N_5981);
nand U6095 (N_6095,N_5715,N_5847);
or U6096 (N_6096,N_5939,N_5990);
or U6097 (N_6097,N_5902,N_5863);
or U6098 (N_6098,N_5779,N_5771);
or U6099 (N_6099,N_5751,N_5916);
or U6100 (N_6100,N_5802,N_5835);
and U6101 (N_6101,N_5775,N_5962);
or U6102 (N_6102,N_5830,N_5872);
and U6103 (N_6103,N_5910,N_5969);
nor U6104 (N_6104,N_5774,N_5755);
or U6105 (N_6105,N_5729,N_5977);
xnor U6106 (N_6106,N_5925,N_5956);
nand U6107 (N_6107,N_5782,N_5795);
and U6108 (N_6108,N_5818,N_5721);
nand U6109 (N_6109,N_5917,N_5874);
nor U6110 (N_6110,N_5780,N_5996);
nor U6111 (N_6111,N_5890,N_5928);
nor U6112 (N_6112,N_5750,N_5845);
nor U6113 (N_6113,N_5883,N_5918);
nor U6114 (N_6114,N_5952,N_5827);
nand U6115 (N_6115,N_5882,N_5739);
nand U6116 (N_6116,N_5987,N_5851);
nand U6117 (N_6117,N_5911,N_5842);
or U6118 (N_6118,N_5723,N_5955);
nor U6119 (N_6119,N_5707,N_5884);
or U6120 (N_6120,N_5978,N_5730);
and U6121 (N_6121,N_5930,N_5776);
or U6122 (N_6122,N_5839,N_5993);
xor U6123 (N_6123,N_5960,N_5986);
and U6124 (N_6124,N_5871,N_5951);
nand U6125 (N_6125,N_5975,N_5788);
xor U6126 (N_6126,N_5720,N_5712);
and U6127 (N_6127,N_5892,N_5798);
xnor U6128 (N_6128,N_5970,N_5999);
and U6129 (N_6129,N_5724,N_5894);
nand U6130 (N_6130,N_5792,N_5831);
or U6131 (N_6131,N_5817,N_5934);
or U6132 (N_6132,N_5801,N_5826);
or U6133 (N_6133,N_5796,N_5734);
and U6134 (N_6134,N_5716,N_5865);
and U6135 (N_6135,N_5992,N_5726);
and U6136 (N_6136,N_5764,N_5855);
nand U6137 (N_6137,N_5804,N_5875);
xnor U6138 (N_6138,N_5767,N_5708);
and U6139 (N_6139,N_5837,N_5966);
nor U6140 (N_6140,N_5799,N_5773);
nand U6141 (N_6141,N_5850,N_5704);
and U6142 (N_6142,N_5859,N_5931);
and U6143 (N_6143,N_5820,N_5959);
nor U6144 (N_6144,N_5852,N_5901);
xor U6145 (N_6145,N_5886,N_5705);
and U6146 (N_6146,N_5834,N_5907);
nand U6147 (N_6147,N_5728,N_5869);
nand U6148 (N_6148,N_5965,N_5791);
or U6149 (N_6149,N_5945,N_5809);
or U6150 (N_6150,N_5845,N_5771);
or U6151 (N_6151,N_5781,N_5868);
xor U6152 (N_6152,N_5841,N_5747);
nor U6153 (N_6153,N_5801,N_5762);
or U6154 (N_6154,N_5707,N_5804);
nand U6155 (N_6155,N_5958,N_5912);
nand U6156 (N_6156,N_5960,N_5830);
and U6157 (N_6157,N_5898,N_5722);
and U6158 (N_6158,N_5765,N_5929);
xnor U6159 (N_6159,N_5877,N_5990);
or U6160 (N_6160,N_5836,N_5761);
and U6161 (N_6161,N_5876,N_5935);
or U6162 (N_6162,N_5879,N_5847);
or U6163 (N_6163,N_5749,N_5919);
or U6164 (N_6164,N_5703,N_5957);
nand U6165 (N_6165,N_5946,N_5831);
nand U6166 (N_6166,N_5732,N_5727);
and U6167 (N_6167,N_5714,N_5949);
and U6168 (N_6168,N_5707,N_5818);
and U6169 (N_6169,N_5962,N_5988);
nor U6170 (N_6170,N_5739,N_5765);
or U6171 (N_6171,N_5745,N_5739);
and U6172 (N_6172,N_5776,N_5968);
and U6173 (N_6173,N_5784,N_5734);
and U6174 (N_6174,N_5909,N_5893);
xnor U6175 (N_6175,N_5754,N_5953);
nand U6176 (N_6176,N_5934,N_5757);
and U6177 (N_6177,N_5901,N_5929);
nand U6178 (N_6178,N_5958,N_5904);
nor U6179 (N_6179,N_5727,N_5722);
nand U6180 (N_6180,N_5874,N_5819);
nor U6181 (N_6181,N_5726,N_5911);
nand U6182 (N_6182,N_5837,N_5785);
xnor U6183 (N_6183,N_5996,N_5914);
or U6184 (N_6184,N_5979,N_5722);
or U6185 (N_6185,N_5904,N_5982);
xor U6186 (N_6186,N_5880,N_5962);
xnor U6187 (N_6187,N_5964,N_5845);
and U6188 (N_6188,N_5862,N_5925);
xor U6189 (N_6189,N_5940,N_5902);
nand U6190 (N_6190,N_5962,N_5755);
nand U6191 (N_6191,N_5918,N_5867);
or U6192 (N_6192,N_5813,N_5810);
nor U6193 (N_6193,N_5946,N_5899);
or U6194 (N_6194,N_5748,N_5810);
nand U6195 (N_6195,N_5996,N_5773);
nor U6196 (N_6196,N_5899,N_5962);
nor U6197 (N_6197,N_5726,N_5766);
nor U6198 (N_6198,N_5793,N_5889);
nand U6199 (N_6199,N_5935,N_5981);
or U6200 (N_6200,N_5791,N_5822);
and U6201 (N_6201,N_5924,N_5997);
nor U6202 (N_6202,N_5703,N_5717);
xor U6203 (N_6203,N_5873,N_5951);
nand U6204 (N_6204,N_5758,N_5902);
or U6205 (N_6205,N_5739,N_5763);
nand U6206 (N_6206,N_5941,N_5744);
xor U6207 (N_6207,N_5810,N_5874);
nor U6208 (N_6208,N_5879,N_5781);
xnor U6209 (N_6209,N_5856,N_5807);
nor U6210 (N_6210,N_5851,N_5707);
nor U6211 (N_6211,N_5777,N_5737);
and U6212 (N_6212,N_5918,N_5713);
xnor U6213 (N_6213,N_5940,N_5919);
xor U6214 (N_6214,N_5886,N_5981);
xor U6215 (N_6215,N_5739,N_5810);
nand U6216 (N_6216,N_5858,N_5975);
and U6217 (N_6217,N_5973,N_5813);
and U6218 (N_6218,N_5728,N_5748);
xor U6219 (N_6219,N_5739,N_5962);
xor U6220 (N_6220,N_5897,N_5817);
nor U6221 (N_6221,N_5864,N_5976);
and U6222 (N_6222,N_5743,N_5787);
nand U6223 (N_6223,N_5886,N_5898);
or U6224 (N_6224,N_5704,N_5966);
or U6225 (N_6225,N_5795,N_5819);
or U6226 (N_6226,N_5767,N_5914);
or U6227 (N_6227,N_5876,N_5768);
nand U6228 (N_6228,N_5737,N_5981);
xor U6229 (N_6229,N_5823,N_5745);
and U6230 (N_6230,N_5920,N_5878);
xor U6231 (N_6231,N_5775,N_5969);
xnor U6232 (N_6232,N_5715,N_5992);
and U6233 (N_6233,N_5856,N_5816);
nand U6234 (N_6234,N_5872,N_5720);
nor U6235 (N_6235,N_5711,N_5866);
or U6236 (N_6236,N_5705,N_5938);
nor U6237 (N_6237,N_5813,N_5998);
nor U6238 (N_6238,N_5999,N_5911);
xor U6239 (N_6239,N_5931,N_5783);
or U6240 (N_6240,N_5833,N_5737);
nor U6241 (N_6241,N_5882,N_5701);
nand U6242 (N_6242,N_5740,N_5889);
and U6243 (N_6243,N_5932,N_5784);
nor U6244 (N_6244,N_5930,N_5841);
nand U6245 (N_6245,N_5790,N_5988);
nor U6246 (N_6246,N_5723,N_5979);
and U6247 (N_6247,N_5743,N_5766);
nor U6248 (N_6248,N_5785,N_5741);
and U6249 (N_6249,N_5834,N_5934);
nand U6250 (N_6250,N_5886,N_5768);
and U6251 (N_6251,N_5805,N_5717);
nand U6252 (N_6252,N_5761,N_5815);
xor U6253 (N_6253,N_5715,N_5767);
or U6254 (N_6254,N_5844,N_5994);
xor U6255 (N_6255,N_5742,N_5823);
xor U6256 (N_6256,N_5934,N_5775);
nand U6257 (N_6257,N_5870,N_5920);
xor U6258 (N_6258,N_5871,N_5753);
nand U6259 (N_6259,N_5987,N_5791);
or U6260 (N_6260,N_5860,N_5783);
and U6261 (N_6261,N_5736,N_5700);
nor U6262 (N_6262,N_5867,N_5828);
xor U6263 (N_6263,N_5932,N_5791);
or U6264 (N_6264,N_5703,N_5771);
xor U6265 (N_6265,N_5987,N_5718);
nor U6266 (N_6266,N_5801,N_5914);
nor U6267 (N_6267,N_5725,N_5807);
xnor U6268 (N_6268,N_5922,N_5795);
or U6269 (N_6269,N_5860,N_5873);
or U6270 (N_6270,N_5922,N_5996);
or U6271 (N_6271,N_5865,N_5730);
nor U6272 (N_6272,N_5990,N_5745);
nor U6273 (N_6273,N_5904,N_5859);
or U6274 (N_6274,N_5980,N_5877);
xnor U6275 (N_6275,N_5999,N_5786);
xnor U6276 (N_6276,N_5873,N_5980);
xor U6277 (N_6277,N_5893,N_5730);
or U6278 (N_6278,N_5700,N_5814);
xor U6279 (N_6279,N_5813,N_5870);
and U6280 (N_6280,N_5777,N_5815);
xor U6281 (N_6281,N_5953,N_5955);
and U6282 (N_6282,N_5995,N_5977);
and U6283 (N_6283,N_5787,N_5866);
and U6284 (N_6284,N_5868,N_5799);
or U6285 (N_6285,N_5863,N_5996);
nand U6286 (N_6286,N_5768,N_5715);
nand U6287 (N_6287,N_5703,N_5719);
nor U6288 (N_6288,N_5938,N_5858);
nand U6289 (N_6289,N_5868,N_5855);
nor U6290 (N_6290,N_5721,N_5923);
nor U6291 (N_6291,N_5924,N_5815);
and U6292 (N_6292,N_5782,N_5946);
or U6293 (N_6293,N_5823,N_5720);
nand U6294 (N_6294,N_5922,N_5846);
nor U6295 (N_6295,N_5860,N_5898);
nor U6296 (N_6296,N_5836,N_5812);
nand U6297 (N_6297,N_5876,N_5723);
nor U6298 (N_6298,N_5866,N_5804);
and U6299 (N_6299,N_5956,N_5889);
nand U6300 (N_6300,N_6189,N_6107);
nor U6301 (N_6301,N_6241,N_6231);
and U6302 (N_6302,N_6153,N_6281);
or U6303 (N_6303,N_6194,N_6266);
nand U6304 (N_6304,N_6036,N_6215);
or U6305 (N_6305,N_6179,N_6233);
and U6306 (N_6306,N_6145,N_6104);
or U6307 (N_6307,N_6103,N_6169);
or U6308 (N_6308,N_6174,N_6030);
or U6309 (N_6309,N_6163,N_6079);
xnor U6310 (N_6310,N_6201,N_6198);
nand U6311 (N_6311,N_6018,N_6001);
or U6312 (N_6312,N_6111,N_6138);
or U6313 (N_6313,N_6095,N_6127);
xnor U6314 (N_6314,N_6149,N_6064);
or U6315 (N_6315,N_6046,N_6056);
nand U6316 (N_6316,N_6044,N_6167);
xnor U6317 (N_6317,N_6272,N_6037);
and U6318 (N_6318,N_6264,N_6066);
and U6319 (N_6319,N_6058,N_6039);
or U6320 (N_6320,N_6236,N_6279);
nand U6321 (N_6321,N_6280,N_6229);
and U6322 (N_6322,N_6200,N_6254);
or U6323 (N_6323,N_6119,N_6223);
and U6324 (N_6324,N_6193,N_6202);
xor U6325 (N_6325,N_6096,N_6188);
or U6326 (N_6326,N_6106,N_6252);
nor U6327 (N_6327,N_6156,N_6112);
nor U6328 (N_6328,N_6147,N_6157);
xnor U6329 (N_6329,N_6092,N_6230);
xnor U6330 (N_6330,N_6070,N_6276);
nand U6331 (N_6331,N_6166,N_6128);
nand U6332 (N_6332,N_6265,N_6115);
nand U6333 (N_6333,N_6097,N_6005);
or U6334 (N_6334,N_6288,N_6297);
nor U6335 (N_6335,N_6244,N_6150);
nor U6336 (N_6336,N_6028,N_6113);
xor U6337 (N_6337,N_6052,N_6226);
nand U6338 (N_6338,N_6178,N_6109);
or U6339 (N_6339,N_6135,N_6181);
or U6340 (N_6340,N_6173,N_6067);
and U6341 (N_6341,N_6218,N_6033);
xor U6342 (N_6342,N_6246,N_6224);
or U6343 (N_6343,N_6094,N_6273);
and U6344 (N_6344,N_6197,N_6195);
xnor U6345 (N_6345,N_6019,N_6069);
nand U6346 (N_6346,N_6294,N_6283);
nand U6347 (N_6347,N_6175,N_6017);
xor U6348 (N_6348,N_6054,N_6216);
nand U6349 (N_6349,N_6075,N_6071);
and U6350 (N_6350,N_6275,N_6220);
nor U6351 (N_6351,N_6255,N_6049);
and U6352 (N_6352,N_6006,N_6148);
nor U6353 (N_6353,N_6131,N_6076);
and U6354 (N_6354,N_6062,N_6289);
nor U6355 (N_6355,N_6022,N_6091);
nor U6356 (N_6356,N_6087,N_6009);
xnor U6357 (N_6357,N_6121,N_6185);
nand U6358 (N_6358,N_6291,N_6081);
xor U6359 (N_6359,N_6152,N_6048);
xor U6360 (N_6360,N_6029,N_6100);
nor U6361 (N_6361,N_6098,N_6032);
and U6362 (N_6362,N_6171,N_6105);
nor U6363 (N_6363,N_6060,N_6180);
and U6364 (N_6364,N_6292,N_6168);
nor U6365 (N_6365,N_6116,N_6011);
xor U6366 (N_6366,N_6008,N_6285);
nand U6367 (N_6367,N_6051,N_6047);
and U6368 (N_6368,N_6007,N_6235);
or U6369 (N_6369,N_6093,N_6159);
xor U6370 (N_6370,N_6065,N_6117);
nand U6371 (N_6371,N_6125,N_6059);
or U6372 (N_6372,N_6222,N_6118);
and U6373 (N_6373,N_6074,N_6211);
nand U6374 (N_6374,N_6146,N_6256);
and U6375 (N_6375,N_6025,N_6089);
xnor U6376 (N_6376,N_6120,N_6261);
nor U6377 (N_6377,N_6110,N_6130);
nor U6378 (N_6378,N_6299,N_6205);
nor U6379 (N_6379,N_6225,N_6249);
and U6380 (N_6380,N_6042,N_6141);
xor U6381 (N_6381,N_6122,N_6014);
nor U6382 (N_6382,N_6088,N_6102);
nand U6383 (N_6383,N_6140,N_6248);
or U6384 (N_6384,N_6270,N_6080);
or U6385 (N_6385,N_6274,N_6034);
and U6386 (N_6386,N_6151,N_6114);
xnor U6387 (N_6387,N_6142,N_6003);
nand U6388 (N_6388,N_6043,N_6251);
or U6389 (N_6389,N_6259,N_6078);
nand U6390 (N_6390,N_6284,N_6026);
xor U6391 (N_6391,N_6160,N_6192);
xor U6392 (N_6392,N_6061,N_6035);
or U6393 (N_6393,N_6257,N_6240);
or U6394 (N_6394,N_6072,N_6186);
xor U6395 (N_6395,N_6023,N_6260);
nor U6396 (N_6396,N_6183,N_6253);
nor U6397 (N_6397,N_6258,N_6132);
or U6398 (N_6398,N_6247,N_6268);
nor U6399 (N_6399,N_6126,N_6184);
nor U6400 (N_6400,N_6158,N_6170);
and U6401 (N_6401,N_6243,N_6155);
nor U6402 (N_6402,N_6084,N_6129);
or U6403 (N_6403,N_6012,N_6000);
nor U6404 (N_6404,N_6177,N_6242);
and U6405 (N_6405,N_6267,N_6083);
nor U6406 (N_6406,N_6282,N_6057);
and U6407 (N_6407,N_6015,N_6154);
nand U6408 (N_6408,N_6027,N_6262);
or U6409 (N_6409,N_6077,N_6024);
nor U6410 (N_6410,N_6295,N_6234);
xor U6411 (N_6411,N_6228,N_6271);
nor U6412 (N_6412,N_6296,N_6085);
or U6413 (N_6413,N_6227,N_6239);
nor U6414 (N_6414,N_6090,N_6203);
nor U6415 (N_6415,N_6108,N_6004);
nor U6416 (N_6416,N_6278,N_6073);
xor U6417 (N_6417,N_6164,N_6063);
nor U6418 (N_6418,N_6206,N_6208);
and U6419 (N_6419,N_6213,N_6101);
or U6420 (N_6420,N_6221,N_6250);
nor U6421 (N_6421,N_6162,N_6207);
xor U6422 (N_6422,N_6269,N_6219);
nand U6423 (N_6423,N_6050,N_6143);
and U6424 (N_6424,N_6068,N_6016);
and U6425 (N_6425,N_6041,N_6191);
and U6426 (N_6426,N_6099,N_6245);
and U6427 (N_6427,N_6040,N_6086);
nor U6428 (N_6428,N_6238,N_6199);
and U6429 (N_6429,N_6204,N_6182);
nor U6430 (N_6430,N_6134,N_6144);
or U6431 (N_6431,N_6293,N_6210);
or U6432 (N_6432,N_6123,N_6286);
or U6433 (N_6433,N_6277,N_6045);
and U6434 (N_6434,N_6165,N_6214);
nor U6435 (N_6435,N_6176,N_6237);
and U6436 (N_6436,N_6031,N_6190);
and U6437 (N_6437,N_6298,N_6161);
and U6438 (N_6438,N_6232,N_6139);
and U6439 (N_6439,N_6133,N_6209);
or U6440 (N_6440,N_6172,N_6020);
xnor U6441 (N_6441,N_6137,N_6038);
nor U6442 (N_6442,N_6021,N_6187);
and U6443 (N_6443,N_6082,N_6263);
or U6444 (N_6444,N_6053,N_6055);
or U6445 (N_6445,N_6290,N_6136);
nand U6446 (N_6446,N_6287,N_6002);
xnor U6447 (N_6447,N_6196,N_6212);
or U6448 (N_6448,N_6010,N_6013);
nor U6449 (N_6449,N_6124,N_6217);
xor U6450 (N_6450,N_6285,N_6260);
and U6451 (N_6451,N_6065,N_6054);
nor U6452 (N_6452,N_6167,N_6000);
or U6453 (N_6453,N_6227,N_6065);
or U6454 (N_6454,N_6262,N_6268);
xor U6455 (N_6455,N_6020,N_6170);
nand U6456 (N_6456,N_6156,N_6272);
and U6457 (N_6457,N_6176,N_6094);
or U6458 (N_6458,N_6053,N_6139);
and U6459 (N_6459,N_6243,N_6147);
nand U6460 (N_6460,N_6166,N_6114);
xor U6461 (N_6461,N_6079,N_6082);
or U6462 (N_6462,N_6031,N_6168);
and U6463 (N_6463,N_6284,N_6162);
nand U6464 (N_6464,N_6064,N_6036);
xor U6465 (N_6465,N_6284,N_6025);
xor U6466 (N_6466,N_6212,N_6006);
nand U6467 (N_6467,N_6003,N_6036);
nor U6468 (N_6468,N_6203,N_6086);
nor U6469 (N_6469,N_6087,N_6179);
or U6470 (N_6470,N_6184,N_6188);
xnor U6471 (N_6471,N_6220,N_6077);
xor U6472 (N_6472,N_6136,N_6163);
and U6473 (N_6473,N_6299,N_6245);
xnor U6474 (N_6474,N_6013,N_6273);
nand U6475 (N_6475,N_6101,N_6026);
or U6476 (N_6476,N_6169,N_6226);
xnor U6477 (N_6477,N_6159,N_6010);
xor U6478 (N_6478,N_6298,N_6114);
or U6479 (N_6479,N_6197,N_6027);
or U6480 (N_6480,N_6204,N_6045);
or U6481 (N_6481,N_6229,N_6071);
xor U6482 (N_6482,N_6074,N_6118);
nor U6483 (N_6483,N_6099,N_6050);
or U6484 (N_6484,N_6006,N_6142);
and U6485 (N_6485,N_6220,N_6168);
or U6486 (N_6486,N_6187,N_6059);
and U6487 (N_6487,N_6195,N_6237);
and U6488 (N_6488,N_6070,N_6052);
and U6489 (N_6489,N_6184,N_6138);
xor U6490 (N_6490,N_6139,N_6029);
nand U6491 (N_6491,N_6058,N_6038);
nand U6492 (N_6492,N_6010,N_6079);
xor U6493 (N_6493,N_6037,N_6133);
xnor U6494 (N_6494,N_6207,N_6108);
and U6495 (N_6495,N_6058,N_6168);
and U6496 (N_6496,N_6031,N_6060);
nor U6497 (N_6497,N_6220,N_6121);
xnor U6498 (N_6498,N_6156,N_6080);
nor U6499 (N_6499,N_6034,N_6181);
nor U6500 (N_6500,N_6185,N_6117);
xnor U6501 (N_6501,N_6025,N_6191);
nand U6502 (N_6502,N_6253,N_6076);
nor U6503 (N_6503,N_6187,N_6154);
nand U6504 (N_6504,N_6083,N_6153);
xnor U6505 (N_6505,N_6160,N_6164);
and U6506 (N_6506,N_6279,N_6149);
nor U6507 (N_6507,N_6260,N_6011);
or U6508 (N_6508,N_6020,N_6290);
xnor U6509 (N_6509,N_6213,N_6072);
xnor U6510 (N_6510,N_6109,N_6194);
nor U6511 (N_6511,N_6124,N_6231);
nor U6512 (N_6512,N_6047,N_6265);
nand U6513 (N_6513,N_6090,N_6160);
and U6514 (N_6514,N_6195,N_6105);
nor U6515 (N_6515,N_6077,N_6025);
nor U6516 (N_6516,N_6283,N_6223);
nor U6517 (N_6517,N_6007,N_6162);
xnor U6518 (N_6518,N_6159,N_6165);
nor U6519 (N_6519,N_6273,N_6209);
or U6520 (N_6520,N_6116,N_6069);
nand U6521 (N_6521,N_6231,N_6244);
xnor U6522 (N_6522,N_6286,N_6024);
or U6523 (N_6523,N_6070,N_6101);
nand U6524 (N_6524,N_6131,N_6027);
and U6525 (N_6525,N_6140,N_6059);
or U6526 (N_6526,N_6269,N_6023);
and U6527 (N_6527,N_6125,N_6237);
and U6528 (N_6528,N_6239,N_6015);
xnor U6529 (N_6529,N_6050,N_6264);
nand U6530 (N_6530,N_6084,N_6018);
xnor U6531 (N_6531,N_6165,N_6135);
or U6532 (N_6532,N_6188,N_6118);
nand U6533 (N_6533,N_6068,N_6154);
xor U6534 (N_6534,N_6224,N_6091);
nand U6535 (N_6535,N_6093,N_6129);
xnor U6536 (N_6536,N_6225,N_6219);
or U6537 (N_6537,N_6210,N_6061);
nand U6538 (N_6538,N_6008,N_6232);
xnor U6539 (N_6539,N_6149,N_6102);
nand U6540 (N_6540,N_6113,N_6173);
nand U6541 (N_6541,N_6114,N_6190);
and U6542 (N_6542,N_6250,N_6257);
and U6543 (N_6543,N_6191,N_6086);
nor U6544 (N_6544,N_6212,N_6075);
or U6545 (N_6545,N_6064,N_6181);
nor U6546 (N_6546,N_6008,N_6293);
xnor U6547 (N_6547,N_6134,N_6229);
nor U6548 (N_6548,N_6141,N_6067);
nor U6549 (N_6549,N_6248,N_6166);
or U6550 (N_6550,N_6123,N_6169);
nand U6551 (N_6551,N_6184,N_6249);
or U6552 (N_6552,N_6075,N_6006);
nor U6553 (N_6553,N_6071,N_6147);
nor U6554 (N_6554,N_6219,N_6139);
xnor U6555 (N_6555,N_6286,N_6136);
or U6556 (N_6556,N_6032,N_6214);
nand U6557 (N_6557,N_6274,N_6277);
nor U6558 (N_6558,N_6039,N_6133);
nand U6559 (N_6559,N_6112,N_6292);
nand U6560 (N_6560,N_6205,N_6240);
nand U6561 (N_6561,N_6227,N_6015);
nor U6562 (N_6562,N_6293,N_6010);
nor U6563 (N_6563,N_6116,N_6202);
nor U6564 (N_6564,N_6233,N_6098);
xnor U6565 (N_6565,N_6297,N_6017);
and U6566 (N_6566,N_6113,N_6036);
or U6567 (N_6567,N_6130,N_6223);
xor U6568 (N_6568,N_6177,N_6297);
nand U6569 (N_6569,N_6179,N_6257);
nor U6570 (N_6570,N_6099,N_6079);
nor U6571 (N_6571,N_6214,N_6087);
nor U6572 (N_6572,N_6135,N_6069);
nor U6573 (N_6573,N_6020,N_6202);
xnor U6574 (N_6574,N_6252,N_6071);
nor U6575 (N_6575,N_6203,N_6204);
or U6576 (N_6576,N_6156,N_6282);
xnor U6577 (N_6577,N_6082,N_6150);
or U6578 (N_6578,N_6245,N_6139);
and U6579 (N_6579,N_6013,N_6109);
nor U6580 (N_6580,N_6060,N_6101);
nand U6581 (N_6581,N_6203,N_6137);
nor U6582 (N_6582,N_6012,N_6213);
and U6583 (N_6583,N_6234,N_6290);
xnor U6584 (N_6584,N_6187,N_6087);
xor U6585 (N_6585,N_6125,N_6065);
nand U6586 (N_6586,N_6122,N_6224);
or U6587 (N_6587,N_6217,N_6070);
xor U6588 (N_6588,N_6217,N_6120);
nand U6589 (N_6589,N_6005,N_6137);
nand U6590 (N_6590,N_6105,N_6114);
nand U6591 (N_6591,N_6009,N_6275);
or U6592 (N_6592,N_6200,N_6250);
xor U6593 (N_6593,N_6219,N_6151);
and U6594 (N_6594,N_6117,N_6101);
nand U6595 (N_6595,N_6152,N_6108);
and U6596 (N_6596,N_6187,N_6102);
xnor U6597 (N_6597,N_6109,N_6154);
xor U6598 (N_6598,N_6288,N_6194);
xnor U6599 (N_6599,N_6257,N_6131);
or U6600 (N_6600,N_6569,N_6595);
nand U6601 (N_6601,N_6350,N_6480);
xnor U6602 (N_6602,N_6384,N_6576);
nand U6603 (N_6603,N_6356,N_6483);
or U6604 (N_6604,N_6415,N_6319);
nor U6605 (N_6605,N_6405,N_6311);
nand U6606 (N_6606,N_6455,N_6430);
xnor U6607 (N_6607,N_6365,N_6476);
and U6608 (N_6608,N_6404,N_6372);
nand U6609 (N_6609,N_6467,N_6532);
nand U6610 (N_6610,N_6582,N_6574);
and U6611 (N_6611,N_6514,N_6570);
and U6612 (N_6612,N_6391,N_6301);
or U6613 (N_6613,N_6414,N_6500);
nand U6614 (N_6614,N_6520,N_6460);
and U6615 (N_6615,N_6482,N_6428);
nor U6616 (N_6616,N_6542,N_6591);
or U6617 (N_6617,N_6472,N_6390);
and U6618 (N_6618,N_6556,N_6388);
and U6619 (N_6619,N_6401,N_6361);
and U6620 (N_6620,N_6515,N_6505);
xnor U6621 (N_6621,N_6522,N_6394);
nor U6622 (N_6622,N_6325,N_6453);
xor U6623 (N_6623,N_6377,N_6433);
nand U6624 (N_6624,N_6594,N_6488);
and U6625 (N_6625,N_6306,N_6529);
and U6626 (N_6626,N_6523,N_6370);
or U6627 (N_6627,N_6445,N_6410);
nor U6628 (N_6628,N_6360,N_6320);
nand U6629 (N_6629,N_6492,N_6411);
and U6630 (N_6630,N_6548,N_6440);
and U6631 (N_6631,N_6392,N_6547);
nor U6632 (N_6632,N_6426,N_6499);
nor U6633 (N_6633,N_6530,N_6322);
and U6634 (N_6634,N_6318,N_6373);
xnor U6635 (N_6635,N_6432,N_6450);
nand U6636 (N_6636,N_6553,N_6321);
nand U6637 (N_6637,N_6544,N_6589);
nor U6638 (N_6638,N_6495,N_6592);
xor U6639 (N_6639,N_6442,N_6314);
nand U6640 (N_6640,N_6380,N_6424);
and U6641 (N_6641,N_6403,N_6407);
and U6642 (N_6642,N_6458,N_6474);
nor U6643 (N_6643,N_6496,N_6333);
and U6644 (N_6644,N_6537,N_6409);
and U6645 (N_6645,N_6359,N_6353);
nor U6646 (N_6646,N_6454,N_6456);
xnor U6647 (N_6647,N_6564,N_6581);
and U6648 (N_6648,N_6446,N_6352);
xnor U6649 (N_6649,N_6434,N_6420);
nand U6650 (N_6650,N_6508,N_6347);
nand U6651 (N_6651,N_6571,N_6302);
nand U6652 (N_6652,N_6381,N_6303);
xnor U6653 (N_6653,N_6389,N_6577);
or U6654 (N_6654,N_6540,N_6503);
nand U6655 (N_6655,N_6315,N_6461);
nor U6656 (N_6656,N_6566,N_6357);
xnor U6657 (N_6657,N_6305,N_6551);
nor U6658 (N_6658,N_6341,N_6338);
nor U6659 (N_6659,N_6310,N_6337);
or U6660 (N_6660,N_6399,N_6451);
or U6661 (N_6661,N_6444,N_6316);
nor U6662 (N_6662,N_6531,N_6408);
xor U6663 (N_6663,N_6528,N_6549);
nand U6664 (N_6664,N_6339,N_6598);
xnor U6665 (N_6665,N_6584,N_6429);
xnor U6666 (N_6666,N_6308,N_6518);
xor U6667 (N_6667,N_6507,N_6493);
and U6668 (N_6668,N_6448,N_6465);
nor U6669 (N_6669,N_6546,N_6578);
or U6670 (N_6670,N_6369,N_6590);
nand U6671 (N_6671,N_6335,N_6368);
nor U6672 (N_6672,N_6447,N_6358);
xor U6673 (N_6673,N_6526,N_6400);
nand U6674 (N_6674,N_6562,N_6466);
or U6675 (N_6675,N_6593,N_6561);
nor U6676 (N_6676,N_6364,N_6575);
xnor U6677 (N_6677,N_6473,N_6417);
nand U6678 (N_6678,N_6557,N_6512);
nand U6679 (N_6679,N_6559,N_6525);
nor U6680 (N_6680,N_6348,N_6469);
nand U6681 (N_6681,N_6504,N_6385);
nor U6682 (N_6682,N_6538,N_6344);
nor U6683 (N_6683,N_6452,N_6382);
nand U6684 (N_6684,N_6478,N_6573);
nand U6685 (N_6685,N_6596,N_6539);
xnor U6686 (N_6686,N_6351,N_6509);
and U6687 (N_6687,N_6489,N_6502);
or U6688 (N_6688,N_6497,N_6587);
nand U6689 (N_6689,N_6545,N_6516);
nor U6690 (N_6690,N_6498,N_6330);
xnor U6691 (N_6691,N_6479,N_6565);
xor U6692 (N_6692,N_6307,N_6402);
xor U6693 (N_6693,N_6580,N_6459);
nor U6694 (N_6694,N_6345,N_6331);
nand U6695 (N_6695,N_6378,N_6519);
nand U6696 (N_6696,N_6386,N_6462);
xor U6697 (N_6697,N_6550,N_6457);
and U6698 (N_6698,N_6543,N_6346);
or U6699 (N_6699,N_6567,N_6463);
nand U6700 (N_6700,N_6572,N_6334);
nor U6701 (N_6701,N_6422,N_6371);
or U6702 (N_6702,N_6486,N_6536);
or U6703 (N_6703,N_6313,N_6541);
nand U6704 (N_6704,N_6328,N_6379);
or U6705 (N_6705,N_6477,N_6355);
nor U6706 (N_6706,N_6324,N_6342);
nor U6707 (N_6707,N_6312,N_6506);
xor U6708 (N_6708,N_6533,N_6332);
nand U6709 (N_6709,N_6362,N_6484);
or U6710 (N_6710,N_6494,N_6363);
or U6711 (N_6711,N_6510,N_6563);
and U6712 (N_6712,N_6406,N_6511);
nor U6713 (N_6713,N_6354,N_6329);
nor U6714 (N_6714,N_6326,N_6586);
nor U6715 (N_6715,N_6376,N_6470);
nor U6716 (N_6716,N_6397,N_6413);
nor U6717 (N_6717,N_6387,N_6513);
or U6718 (N_6718,N_6554,N_6568);
nor U6719 (N_6719,N_6421,N_6588);
nor U6720 (N_6720,N_6437,N_6481);
nor U6721 (N_6721,N_6427,N_6468);
nor U6722 (N_6722,N_6501,N_6396);
nand U6723 (N_6723,N_6579,N_6340);
nand U6724 (N_6724,N_6323,N_6491);
and U6725 (N_6725,N_6534,N_6583);
xor U6726 (N_6726,N_6471,N_6552);
nand U6727 (N_6727,N_6517,N_6419);
nand U6728 (N_6728,N_6597,N_6490);
and U6729 (N_6729,N_6395,N_6412);
nor U6730 (N_6730,N_6304,N_6524);
xor U6731 (N_6731,N_6317,N_6343);
nor U6732 (N_6732,N_6441,N_6367);
or U6733 (N_6733,N_6560,N_6383);
xor U6734 (N_6734,N_6521,N_6464);
nand U6735 (N_6735,N_6475,N_6300);
xnor U6736 (N_6736,N_6443,N_6435);
nand U6737 (N_6737,N_6599,N_6535);
and U6738 (N_6738,N_6418,N_6585);
nand U6739 (N_6739,N_6431,N_6487);
or U6740 (N_6740,N_6416,N_6393);
xor U6741 (N_6741,N_6425,N_6558);
nand U6742 (N_6742,N_6555,N_6374);
or U6743 (N_6743,N_6366,N_6349);
and U6744 (N_6744,N_6438,N_6336);
or U6745 (N_6745,N_6375,N_6449);
and U6746 (N_6746,N_6436,N_6423);
xor U6747 (N_6747,N_6439,N_6309);
nand U6748 (N_6748,N_6485,N_6398);
and U6749 (N_6749,N_6327,N_6527);
or U6750 (N_6750,N_6448,N_6510);
or U6751 (N_6751,N_6489,N_6548);
xnor U6752 (N_6752,N_6507,N_6321);
xor U6753 (N_6753,N_6442,N_6543);
nor U6754 (N_6754,N_6304,N_6463);
xnor U6755 (N_6755,N_6415,N_6312);
nand U6756 (N_6756,N_6494,N_6334);
and U6757 (N_6757,N_6461,N_6345);
nor U6758 (N_6758,N_6487,N_6438);
or U6759 (N_6759,N_6485,N_6444);
nand U6760 (N_6760,N_6441,N_6375);
xnor U6761 (N_6761,N_6575,N_6348);
nor U6762 (N_6762,N_6557,N_6430);
nand U6763 (N_6763,N_6337,N_6485);
or U6764 (N_6764,N_6527,N_6573);
or U6765 (N_6765,N_6495,N_6471);
xor U6766 (N_6766,N_6563,N_6333);
or U6767 (N_6767,N_6369,N_6405);
nor U6768 (N_6768,N_6568,N_6308);
or U6769 (N_6769,N_6507,N_6346);
nor U6770 (N_6770,N_6534,N_6449);
xor U6771 (N_6771,N_6453,N_6462);
xor U6772 (N_6772,N_6407,N_6570);
and U6773 (N_6773,N_6334,N_6305);
nand U6774 (N_6774,N_6369,N_6395);
xnor U6775 (N_6775,N_6430,N_6420);
nand U6776 (N_6776,N_6381,N_6373);
or U6777 (N_6777,N_6470,N_6302);
xnor U6778 (N_6778,N_6442,N_6321);
nand U6779 (N_6779,N_6390,N_6467);
nand U6780 (N_6780,N_6392,N_6569);
and U6781 (N_6781,N_6365,N_6453);
xor U6782 (N_6782,N_6358,N_6582);
nor U6783 (N_6783,N_6468,N_6466);
and U6784 (N_6784,N_6443,N_6562);
xor U6785 (N_6785,N_6549,N_6395);
nor U6786 (N_6786,N_6418,N_6380);
nor U6787 (N_6787,N_6349,N_6457);
nor U6788 (N_6788,N_6328,N_6365);
and U6789 (N_6789,N_6442,N_6372);
xnor U6790 (N_6790,N_6442,N_6387);
nor U6791 (N_6791,N_6440,N_6375);
and U6792 (N_6792,N_6415,N_6478);
and U6793 (N_6793,N_6452,N_6470);
xnor U6794 (N_6794,N_6404,N_6408);
nand U6795 (N_6795,N_6469,N_6322);
xor U6796 (N_6796,N_6591,N_6596);
nor U6797 (N_6797,N_6349,N_6510);
xor U6798 (N_6798,N_6462,N_6532);
xor U6799 (N_6799,N_6487,N_6336);
nor U6800 (N_6800,N_6320,N_6344);
or U6801 (N_6801,N_6359,N_6305);
or U6802 (N_6802,N_6406,N_6348);
and U6803 (N_6803,N_6565,N_6303);
nand U6804 (N_6804,N_6375,N_6356);
xor U6805 (N_6805,N_6392,N_6309);
and U6806 (N_6806,N_6330,N_6546);
or U6807 (N_6807,N_6497,N_6389);
and U6808 (N_6808,N_6535,N_6459);
nor U6809 (N_6809,N_6579,N_6465);
xnor U6810 (N_6810,N_6426,N_6527);
xor U6811 (N_6811,N_6419,N_6580);
nor U6812 (N_6812,N_6382,N_6548);
nand U6813 (N_6813,N_6551,N_6344);
nor U6814 (N_6814,N_6395,N_6426);
nand U6815 (N_6815,N_6528,N_6405);
nand U6816 (N_6816,N_6514,N_6465);
and U6817 (N_6817,N_6392,N_6493);
or U6818 (N_6818,N_6361,N_6328);
or U6819 (N_6819,N_6466,N_6470);
and U6820 (N_6820,N_6414,N_6535);
or U6821 (N_6821,N_6386,N_6328);
xor U6822 (N_6822,N_6429,N_6410);
or U6823 (N_6823,N_6542,N_6576);
or U6824 (N_6824,N_6591,N_6527);
xnor U6825 (N_6825,N_6519,N_6522);
and U6826 (N_6826,N_6408,N_6411);
and U6827 (N_6827,N_6572,N_6403);
xor U6828 (N_6828,N_6543,N_6303);
and U6829 (N_6829,N_6576,N_6351);
xnor U6830 (N_6830,N_6493,N_6378);
nand U6831 (N_6831,N_6388,N_6370);
and U6832 (N_6832,N_6454,N_6382);
nand U6833 (N_6833,N_6421,N_6574);
xor U6834 (N_6834,N_6351,N_6520);
nand U6835 (N_6835,N_6310,N_6540);
or U6836 (N_6836,N_6412,N_6581);
xor U6837 (N_6837,N_6450,N_6562);
nor U6838 (N_6838,N_6587,N_6357);
xnor U6839 (N_6839,N_6513,N_6301);
nor U6840 (N_6840,N_6351,N_6477);
nor U6841 (N_6841,N_6334,N_6449);
nand U6842 (N_6842,N_6563,N_6494);
and U6843 (N_6843,N_6363,N_6400);
nand U6844 (N_6844,N_6446,N_6523);
and U6845 (N_6845,N_6350,N_6428);
xnor U6846 (N_6846,N_6435,N_6352);
nor U6847 (N_6847,N_6384,N_6414);
nand U6848 (N_6848,N_6586,N_6339);
nand U6849 (N_6849,N_6489,N_6583);
or U6850 (N_6850,N_6381,N_6387);
nor U6851 (N_6851,N_6484,N_6385);
nand U6852 (N_6852,N_6419,N_6313);
nor U6853 (N_6853,N_6560,N_6404);
xor U6854 (N_6854,N_6595,N_6490);
nand U6855 (N_6855,N_6494,N_6498);
and U6856 (N_6856,N_6504,N_6564);
nand U6857 (N_6857,N_6438,N_6479);
and U6858 (N_6858,N_6436,N_6462);
nor U6859 (N_6859,N_6411,N_6307);
nand U6860 (N_6860,N_6510,N_6565);
or U6861 (N_6861,N_6306,N_6558);
or U6862 (N_6862,N_6401,N_6587);
or U6863 (N_6863,N_6584,N_6516);
and U6864 (N_6864,N_6549,N_6401);
nor U6865 (N_6865,N_6365,N_6538);
nor U6866 (N_6866,N_6527,N_6350);
nor U6867 (N_6867,N_6316,N_6308);
nand U6868 (N_6868,N_6377,N_6358);
nor U6869 (N_6869,N_6425,N_6394);
or U6870 (N_6870,N_6538,N_6346);
or U6871 (N_6871,N_6488,N_6411);
nor U6872 (N_6872,N_6566,N_6558);
nand U6873 (N_6873,N_6352,N_6577);
and U6874 (N_6874,N_6338,N_6452);
nor U6875 (N_6875,N_6308,N_6517);
xor U6876 (N_6876,N_6429,N_6440);
nor U6877 (N_6877,N_6354,N_6319);
and U6878 (N_6878,N_6457,N_6387);
or U6879 (N_6879,N_6481,N_6585);
nor U6880 (N_6880,N_6379,N_6535);
nand U6881 (N_6881,N_6385,N_6528);
nor U6882 (N_6882,N_6498,N_6320);
nor U6883 (N_6883,N_6438,N_6364);
xnor U6884 (N_6884,N_6373,N_6462);
nor U6885 (N_6885,N_6540,N_6375);
nand U6886 (N_6886,N_6462,N_6510);
nor U6887 (N_6887,N_6504,N_6370);
nand U6888 (N_6888,N_6363,N_6379);
or U6889 (N_6889,N_6579,N_6347);
xnor U6890 (N_6890,N_6526,N_6432);
and U6891 (N_6891,N_6530,N_6391);
and U6892 (N_6892,N_6549,N_6573);
and U6893 (N_6893,N_6316,N_6388);
nand U6894 (N_6894,N_6363,N_6542);
xor U6895 (N_6895,N_6423,N_6369);
and U6896 (N_6896,N_6476,N_6340);
nor U6897 (N_6897,N_6495,N_6587);
nor U6898 (N_6898,N_6542,N_6510);
nand U6899 (N_6899,N_6363,N_6423);
xnor U6900 (N_6900,N_6695,N_6730);
or U6901 (N_6901,N_6692,N_6757);
nand U6902 (N_6902,N_6728,N_6867);
nor U6903 (N_6903,N_6762,N_6741);
nor U6904 (N_6904,N_6897,N_6662);
and U6905 (N_6905,N_6686,N_6638);
and U6906 (N_6906,N_6876,N_6796);
xnor U6907 (N_6907,N_6860,N_6841);
xnor U6908 (N_6908,N_6767,N_6822);
xnor U6909 (N_6909,N_6764,N_6843);
nand U6910 (N_6910,N_6613,N_6681);
xnor U6911 (N_6911,N_6604,N_6862);
xnor U6912 (N_6912,N_6827,N_6808);
nand U6913 (N_6913,N_6632,N_6611);
and U6914 (N_6914,N_6806,N_6794);
xor U6915 (N_6915,N_6785,N_6749);
and U6916 (N_6916,N_6780,N_6651);
nor U6917 (N_6917,N_6755,N_6690);
or U6918 (N_6918,N_6709,N_6784);
xnor U6919 (N_6919,N_6866,N_6696);
and U6920 (N_6920,N_6641,N_6700);
or U6921 (N_6921,N_6664,N_6697);
or U6922 (N_6922,N_6620,N_6873);
nand U6923 (N_6923,N_6868,N_6642);
or U6924 (N_6924,N_6615,N_6707);
nor U6925 (N_6925,N_6846,N_6857);
nor U6926 (N_6926,N_6782,N_6809);
nand U6927 (N_6927,N_6607,N_6723);
nor U6928 (N_6928,N_6833,N_6655);
or U6929 (N_6929,N_6787,N_6609);
xor U6930 (N_6930,N_6701,N_6653);
nand U6931 (N_6931,N_6631,N_6874);
nor U6932 (N_6932,N_6859,N_6858);
or U6933 (N_6933,N_6702,N_6880);
nand U6934 (N_6934,N_6824,N_6849);
and U6935 (N_6935,N_6769,N_6750);
or U6936 (N_6936,N_6842,N_6602);
nor U6937 (N_6937,N_6823,N_6654);
xnor U6938 (N_6938,N_6797,N_6618);
or U6939 (N_6939,N_6899,N_6813);
and U6940 (N_6940,N_6805,N_6889);
nand U6941 (N_6941,N_6839,N_6743);
nand U6942 (N_6942,N_6803,N_6886);
or U6943 (N_6943,N_6622,N_6688);
xor U6944 (N_6944,N_6624,N_6721);
nor U6945 (N_6945,N_6756,N_6885);
nand U6946 (N_6946,N_6704,N_6847);
xor U6947 (N_6947,N_6652,N_6870);
nor U6948 (N_6948,N_6814,N_6689);
and U6949 (N_6949,N_6738,N_6819);
or U6950 (N_6950,N_6773,N_6826);
nand U6951 (N_6951,N_6861,N_6856);
nand U6952 (N_6952,N_6614,N_6636);
nand U6953 (N_6953,N_6804,N_6810);
and U6954 (N_6954,N_6894,N_6678);
and U6955 (N_6955,N_6605,N_6768);
nor U6956 (N_6956,N_6674,N_6603);
nand U6957 (N_6957,N_6657,N_6830);
nand U6958 (N_6958,N_6684,N_6747);
xnor U6959 (N_6959,N_6848,N_6844);
or U6960 (N_6960,N_6727,N_6670);
nand U6961 (N_6961,N_6711,N_6772);
nand U6962 (N_6962,N_6724,N_6647);
nor U6963 (N_6963,N_6891,N_6759);
and U6964 (N_6964,N_6896,N_6640);
or U6965 (N_6965,N_6816,N_6845);
xnor U6966 (N_6966,N_6850,N_6671);
or U6967 (N_6967,N_6837,N_6663);
nor U6968 (N_6968,N_6892,N_6853);
nor U6969 (N_6969,N_6659,N_6685);
nand U6970 (N_6970,N_6673,N_6777);
or U6971 (N_6971,N_6855,N_6682);
xor U6972 (N_6972,N_6739,N_6706);
nor U6973 (N_6973,N_6765,N_6606);
xnor U6974 (N_6974,N_6877,N_6815);
and U6975 (N_6975,N_6881,N_6617);
and U6976 (N_6976,N_6601,N_6717);
and U6977 (N_6977,N_6629,N_6879);
xnor U6978 (N_6978,N_6888,N_6715);
and U6979 (N_6979,N_6616,N_6869);
nor U6980 (N_6980,N_6890,N_6751);
nand U6981 (N_6981,N_6731,N_6795);
nor U6982 (N_6982,N_6828,N_6737);
nor U6983 (N_6983,N_6672,N_6746);
or U6984 (N_6984,N_6722,N_6716);
nor U6985 (N_6985,N_6887,N_6771);
or U6986 (N_6986,N_6761,N_6725);
nand U6987 (N_6987,N_6812,N_6748);
nand U6988 (N_6988,N_6838,N_6625);
or U6989 (N_6989,N_6875,N_6644);
nor U6990 (N_6990,N_6893,N_6650);
xor U6991 (N_6991,N_6781,N_6610);
and U6992 (N_6992,N_6821,N_6884);
xnor U6993 (N_6993,N_6788,N_6628);
nor U6994 (N_6994,N_6753,N_6829);
xnor U6995 (N_6995,N_6608,N_6691);
or U6996 (N_6996,N_6705,N_6871);
nor U6997 (N_6997,N_6831,N_6758);
nand U6998 (N_6998,N_6736,N_6648);
nand U6999 (N_6999,N_6735,N_6898);
and U7000 (N_7000,N_6635,N_6710);
nand U7001 (N_7001,N_6752,N_6600);
xnor U7002 (N_7002,N_6786,N_6683);
and U7003 (N_7003,N_6744,N_6801);
or U7004 (N_7004,N_6779,N_6817);
nor U7005 (N_7005,N_6693,N_6745);
xnor U7006 (N_7006,N_6851,N_6679);
nor U7007 (N_7007,N_6612,N_6740);
xnor U7008 (N_7008,N_6699,N_6793);
and U7009 (N_7009,N_6720,N_6726);
or U7010 (N_7010,N_6763,N_6637);
and U7011 (N_7011,N_6770,N_6626);
nand U7012 (N_7012,N_6719,N_6656);
or U7013 (N_7013,N_6643,N_6776);
nor U7014 (N_7014,N_6698,N_6669);
or U7015 (N_7015,N_6694,N_6807);
xor U7016 (N_7016,N_6760,N_6633);
xnor U7017 (N_7017,N_6811,N_6623);
nand U7018 (N_7018,N_6718,N_6754);
or U7019 (N_7019,N_6832,N_6661);
or U7020 (N_7020,N_6791,N_6825);
nand U7021 (N_7021,N_6621,N_6840);
or U7022 (N_7022,N_6766,N_6639);
xnor U7023 (N_7023,N_6802,N_6783);
xor U7024 (N_7024,N_6864,N_6789);
xnor U7025 (N_7025,N_6677,N_6820);
or U7026 (N_7026,N_6818,N_6792);
or U7027 (N_7027,N_6634,N_6835);
or U7028 (N_7028,N_6666,N_6734);
nor U7029 (N_7029,N_6882,N_6676);
and U7030 (N_7030,N_6798,N_6852);
or U7031 (N_7031,N_6799,N_6742);
or U7032 (N_7032,N_6646,N_6733);
nand U7033 (N_7033,N_6883,N_6778);
nor U7034 (N_7034,N_6667,N_6712);
nand U7035 (N_7035,N_6863,N_6627);
nor U7036 (N_7036,N_6675,N_6680);
nor U7037 (N_7037,N_6834,N_6714);
and U7038 (N_7038,N_6703,N_6729);
or U7039 (N_7039,N_6854,N_6865);
xnor U7040 (N_7040,N_6790,N_6665);
xor U7041 (N_7041,N_6658,N_6895);
nand U7042 (N_7042,N_6732,N_6872);
nor U7043 (N_7043,N_6775,N_6660);
or U7044 (N_7044,N_6800,N_6619);
xnor U7045 (N_7045,N_6713,N_6649);
and U7046 (N_7046,N_6645,N_6687);
and U7047 (N_7047,N_6708,N_6836);
nand U7048 (N_7048,N_6630,N_6774);
nor U7049 (N_7049,N_6878,N_6668);
and U7050 (N_7050,N_6710,N_6617);
and U7051 (N_7051,N_6602,N_6646);
xnor U7052 (N_7052,N_6620,N_6861);
and U7053 (N_7053,N_6670,N_6776);
nand U7054 (N_7054,N_6899,N_6768);
and U7055 (N_7055,N_6625,N_6754);
or U7056 (N_7056,N_6758,N_6887);
or U7057 (N_7057,N_6704,N_6666);
nor U7058 (N_7058,N_6717,N_6866);
xnor U7059 (N_7059,N_6627,N_6742);
nor U7060 (N_7060,N_6660,N_6758);
nand U7061 (N_7061,N_6615,N_6803);
nor U7062 (N_7062,N_6810,N_6833);
xnor U7063 (N_7063,N_6735,N_6835);
nand U7064 (N_7064,N_6680,N_6887);
and U7065 (N_7065,N_6689,N_6659);
nor U7066 (N_7066,N_6742,N_6676);
nor U7067 (N_7067,N_6633,N_6824);
or U7068 (N_7068,N_6702,N_6858);
nand U7069 (N_7069,N_6733,N_6657);
nor U7070 (N_7070,N_6823,N_6737);
xor U7071 (N_7071,N_6727,N_6651);
nand U7072 (N_7072,N_6815,N_6727);
or U7073 (N_7073,N_6879,N_6812);
nand U7074 (N_7074,N_6840,N_6777);
xor U7075 (N_7075,N_6653,N_6788);
or U7076 (N_7076,N_6642,N_6681);
and U7077 (N_7077,N_6614,N_6648);
xnor U7078 (N_7078,N_6874,N_6625);
or U7079 (N_7079,N_6805,N_6742);
nand U7080 (N_7080,N_6817,N_6692);
nor U7081 (N_7081,N_6659,N_6609);
xnor U7082 (N_7082,N_6630,N_6755);
nor U7083 (N_7083,N_6693,N_6821);
xor U7084 (N_7084,N_6619,N_6871);
nor U7085 (N_7085,N_6794,N_6672);
or U7086 (N_7086,N_6689,N_6728);
and U7087 (N_7087,N_6609,N_6694);
nand U7088 (N_7088,N_6644,N_6746);
nand U7089 (N_7089,N_6723,N_6890);
nand U7090 (N_7090,N_6874,N_6628);
or U7091 (N_7091,N_6712,N_6669);
and U7092 (N_7092,N_6638,N_6836);
xnor U7093 (N_7093,N_6660,N_6767);
nand U7094 (N_7094,N_6696,N_6797);
and U7095 (N_7095,N_6630,N_6822);
nand U7096 (N_7096,N_6759,N_6606);
and U7097 (N_7097,N_6884,N_6763);
or U7098 (N_7098,N_6629,N_6857);
xor U7099 (N_7099,N_6705,N_6895);
nand U7100 (N_7100,N_6836,N_6835);
or U7101 (N_7101,N_6816,N_6822);
or U7102 (N_7102,N_6777,N_6687);
xor U7103 (N_7103,N_6814,N_6881);
xor U7104 (N_7104,N_6867,N_6861);
and U7105 (N_7105,N_6789,N_6795);
or U7106 (N_7106,N_6683,N_6714);
nor U7107 (N_7107,N_6679,N_6762);
xor U7108 (N_7108,N_6819,N_6674);
xor U7109 (N_7109,N_6850,N_6769);
or U7110 (N_7110,N_6849,N_6601);
xnor U7111 (N_7111,N_6776,N_6862);
xor U7112 (N_7112,N_6708,N_6744);
xor U7113 (N_7113,N_6796,N_6753);
nand U7114 (N_7114,N_6866,N_6843);
nor U7115 (N_7115,N_6703,N_6624);
xnor U7116 (N_7116,N_6832,N_6851);
or U7117 (N_7117,N_6795,N_6653);
or U7118 (N_7118,N_6835,N_6894);
nor U7119 (N_7119,N_6828,N_6897);
xnor U7120 (N_7120,N_6806,N_6652);
nand U7121 (N_7121,N_6684,N_6631);
nor U7122 (N_7122,N_6820,N_6844);
or U7123 (N_7123,N_6638,N_6795);
xor U7124 (N_7124,N_6730,N_6732);
xor U7125 (N_7125,N_6706,N_6873);
or U7126 (N_7126,N_6750,N_6831);
nand U7127 (N_7127,N_6696,N_6694);
nor U7128 (N_7128,N_6604,N_6622);
xnor U7129 (N_7129,N_6876,N_6782);
or U7130 (N_7130,N_6863,N_6859);
nor U7131 (N_7131,N_6654,N_6888);
nand U7132 (N_7132,N_6830,N_6825);
nand U7133 (N_7133,N_6815,N_6706);
nor U7134 (N_7134,N_6865,N_6673);
and U7135 (N_7135,N_6709,N_6832);
nor U7136 (N_7136,N_6818,N_6822);
xor U7137 (N_7137,N_6896,N_6754);
nor U7138 (N_7138,N_6774,N_6871);
or U7139 (N_7139,N_6701,N_6821);
or U7140 (N_7140,N_6846,N_6795);
xor U7141 (N_7141,N_6753,N_6846);
and U7142 (N_7142,N_6694,N_6743);
and U7143 (N_7143,N_6773,N_6618);
or U7144 (N_7144,N_6758,N_6634);
and U7145 (N_7145,N_6618,N_6628);
nor U7146 (N_7146,N_6661,N_6692);
and U7147 (N_7147,N_6767,N_6858);
nand U7148 (N_7148,N_6807,N_6803);
nand U7149 (N_7149,N_6848,N_6698);
xnor U7150 (N_7150,N_6799,N_6785);
and U7151 (N_7151,N_6761,N_6813);
nand U7152 (N_7152,N_6742,N_6609);
xnor U7153 (N_7153,N_6815,N_6748);
or U7154 (N_7154,N_6769,N_6828);
nand U7155 (N_7155,N_6890,N_6893);
nor U7156 (N_7156,N_6634,N_6784);
xnor U7157 (N_7157,N_6699,N_6776);
or U7158 (N_7158,N_6727,N_6707);
nand U7159 (N_7159,N_6762,N_6778);
and U7160 (N_7160,N_6856,N_6609);
and U7161 (N_7161,N_6838,N_6633);
xnor U7162 (N_7162,N_6803,N_6867);
nor U7163 (N_7163,N_6751,N_6806);
xnor U7164 (N_7164,N_6806,N_6705);
or U7165 (N_7165,N_6716,N_6861);
nand U7166 (N_7166,N_6798,N_6858);
and U7167 (N_7167,N_6690,N_6788);
nor U7168 (N_7168,N_6896,N_6864);
xnor U7169 (N_7169,N_6743,N_6692);
or U7170 (N_7170,N_6618,N_6673);
nand U7171 (N_7171,N_6820,N_6755);
or U7172 (N_7172,N_6804,N_6722);
nand U7173 (N_7173,N_6868,N_6881);
or U7174 (N_7174,N_6803,N_6661);
nand U7175 (N_7175,N_6637,N_6868);
xor U7176 (N_7176,N_6885,N_6832);
nor U7177 (N_7177,N_6601,N_6840);
or U7178 (N_7178,N_6850,N_6894);
nor U7179 (N_7179,N_6776,N_6827);
and U7180 (N_7180,N_6821,N_6695);
xnor U7181 (N_7181,N_6810,N_6625);
nand U7182 (N_7182,N_6618,N_6771);
and U7183 (N_7183,N_6608,N_6677);
nor U7184 (N_7184,N_6864,N_6677);
nand U7185 (N_7185,N_6851,N_6668);
nand U7186 (N_7186,N_6812,N_6663);
nor U7187 (N_7187,N_6791,N_6793);
nor U7188 (N_7188,N_6703,N_6873);
nand U7189 (N_7189,N_6713,N_6689);
or U7190 (N_7190,N_6631,N_6749);
and U7191 (N_7191,N_6704,N_6846);
xnor U7192 (N_7192,N_6772,N_6762);
nor U7193 (N_7193,N_6712,N_6681);
nor U7194 (N_7194,N_6743,N_6792);
and U7195 (N_7195,N_6695,N_6621);
nor U7196 (N_7196,N_6760,N_6713);
or U7197 (N_7197,N_6610,N_6739);
and U7198 (N_7198,N_6696,N_6897);
xnor U7199 (N_7199,N_6712,N_6690);
nor U7200 (N_7200,N_7041,N_7049);
and U7201 (N_7201,N_6905,N_6914);
or U7202 (N_7202,N_7152,N_7000);
and U7203 (N_7203,N_7077,N_6958);
or U7204 (N_7204,N_7020,N_6917);
and U7205 (N_7205,N_6987,N_7151);
nor U7206 (N_7206,N_6955,N_6923);
xor U7207 (N_7207,N_7046,N_7119);
nor U7208 (N_7208,N_7168,N_7076);
xor U7209 (N_7209,N_7080,N_7034);
and U7210 (N_7210,N_7062,N_7117);
or U7211 (N_7211,N_7146,N_7091);
and U7212 (N_7212,N_7142,N_6918);
nand U7213 (N_7213,N_6942,N_7144);
or U7214 (N_7214,N_6907,N_7186);
xnor U7215 (N_7215,N_7145,N_6996);
xor U7216 (N_7216,N_6973,N_7054);
xor U7217 (N_7217,N_7134,N_7095);
and U7218 (N_7218,N_7038,N_7036);
nor U7219 (N_7219,N_7100,N_7016);
nor U7220 (N_7220,N_7101,N_6977);
nand U7221 (N_7221,N_7092,N_7118);
nand U7222 (N_7222,N_7114,N_7013);
nor U7223 (N_7223,N_7008,N_7019);
nand U7224 (N_7224,N_6998,N_7172);
xor U7225 (N_7225,N_7175,N_7025);
xor U7226 (N_7226,N_6948,N_7164);
nor U7227 (N_7227,N_7032,N_7170);
and U7228 (N_7228,N_7198,N_6904);
nor U7229 (N_7229,N_7199,N_7193);
and U7230 (N_7230,N_6952,N_6901);
and U7231 (N_7231,N_7147,N_6926);
xor U7232 (N_7232,N_6900,N_7157);
xnor U7233 (N_7233,N_7061,N_7082);
nand U7234 (N_7234,N_7060,N_7014);
xor U7235 (N_7235,N_7088,N_6972);
nor U7236 (N_7236,N_7166,N_7093);
nand U7237 (N_7237,N_6940,N_7187);
nand U7238 (N_7238,N_6989,N_7174);
and U7239 (N_7239,N_7022,N_7131);
nand U7240 (N_7240,N_7056,N_7139);
or U7241 (N_7241,N_7023,N_7110);
and U7242 (N_7242,N_6946,N_6980);
or U7243 (N_7243,N_7084,N_7192);
or U7244 (N_7244,N_7071,N_6944);
xor U7245 (N_7245,N_7051,N_7171);
and U7246 (N_7246,N_7105,N_7154);
nor U7247 (N_7247,N_7140,N_6978);
or U7248 (N_7248,N_7129,N_7126);
nor U7249 (N_7249,N_7148,N_7015);
or U7250 (N_7250,N_7159,N_6986);
or U7251 (N_7251,N_6967,N_7045);
nor U7252 (N_7252,N_7068,N_7085);
nor U7253 (N_7253,N_7055,N_7184);
and U7254 (N_7254,N_7059,N_7173);
nand U7255 (N_7255,N_6939,N_7039);
or U7256 (N_7256,N_7127,N_7162);
and U7257 (N_7257,N_7149,N_7042);
or U7258 (N_7258,N_6976,N_6930);
xnor U7259 (N_7259,N_7160,N_6994);
or U7260 (N_7260,N_7087,N_6916);
nor U7261 (N_7261,N_7132,N_6934);
nor U7262 (N_7262,N_7112,N_7073);
nor U7263 (N_7263,N_7133,N_6949);
nor U7264 (N_7264,N_7111,N_7012);
or U7265 (N_7265,N_6991,N_6915);
or U7266 (N_7266,N_6965,N_6935);
xnor U7267 (N_7267,N_7004,N_7052);
and U7268 (N_7268,N_7047,N_6988);
and U7269 (N_7269,N_7153,N_7120);
nor U7270 (N_7270,N_7081,N_7155);
nand U7271 (N_7271,N_7074,N_6961);
nor U7272 (N_7272,N_6919,N_7031);
xnor U7273 (N_7273,N_6982,N_7001);
nand U7274 (N_7274,N_7072,N_7169);
nand U7275 (N_7275,N_6945,N_7190);
and U7276 (N_7276,N_6936,N_7075);
and U7277 (N_7277,N_6979,N_7083);
xor U7278 (N_7278,N_7136,N_7125);
nor U7279 (N_7279,N_6941,N_6964);
xnor U7280 (N_7280,N_7048,N_7098);
nand U7281 (N_7281,N_6950,N_6908);
nand U7282 (N_7282,N_6911,N_7130);
nor U7283 (N_7283,N_6959,N_7165);
nor U7284 (N_7284,N_7156,N_7044);
nand U7285 (N_7285,N_7058,N_7137);
nor U7286 (N_7286,N_6990,N_6953);
and U7287 (N_7287,N_6925,N_7094);
nand U7288 (N_7288,N_7010,N_7069);
nor U7289 (N_7289,N_6954,N_6928);
nand U7290 (N_7290,N_7035,N_6974);
nor U7291 (N_7291,N_7115,N_7182);
xnor U7292 (N_7292,N_7177,N_7189);
nand U7293 (N_7293,N_7141,N_7099);
or U7294 (N_7294,N_7089,N_7167);
nor U7295 (N_7295,N_6924,N_7103);
xor U7296 (N_7296,N_7090,N_6943);
or U7297 (N_7297,N_6995,N_7197);
nand U7298 (N_7298,N_7138,N_7070);
and U7299 (N_7299,N_7116,N_7053);
xor U7300 (N_7300,N_7188,N_7106);
xnor U7301 (N_7301,N_7161,N_7064);
xnor U7302 (N_7302,N_7040,N_7135);
or U7303 (N_7303,N_7176,N_7109);
or U7304 (N_7304,N_7123,N_7102);
nor U7305 (N_7305,N_7196,N_7179);
xor U7306 (N_7306,N_7002,N_7033);
and U7307 (N_7307,N_7024,N_6933);
xnor U7308 (N_7308,N_7078,N_7150);
and U7309 (N_7309,N_6906,N_6931);
nand U7310 (N_7310,N_7181,N_7096);
nor U7311 (N_7311,N_7097,N_7009);
nor U7312 (N_7312,N_7191,N_6903);
or U7313 (N_7313,N_7143,N_7183);
nand U7314 (N_7314,N_6983,N_6997);
nor U7315 (N_7315,N_6902,N_7017);
nor U7316 (N_7316,N_6921,N_7065);
xnor U7317 (N_7317,N_7030,N_7108);
xor U7318 (N_7318,N_7107,N_6999);
nand U7319 (N_7319,N_6963,N_7163);
and U7320 (N_7320,N_7194,N_7066);
xnor U7321 (N_7321,N_6938,N_6920);
xor U7322 (N_7322,N_6957,N_7028);
xor U7323 (N_7323,N_6951,N_6984);
xor U7324 (N_7324,N_7003,N_7043);
xor U7325 (N_7325,N_6968,N_7079);
or U7326 (N_7326,N_7122,N_7185);
or U7327 (N_7327,N_7104,N_7178);
nor U7328 (N_7328,N_7121,N_7029);
xnor U7329 (N_7329,N_7021,N_7011);
nand U7330 (N_7330,N_6966,N_6970);
nand U7331 (N_7331,N_7063,N_6962);
and U7332 (N_7332,N_6922,N_6932);
nand U7333 (N_7333,N_6981,N_6969);
nand U7334 (N_7334,N_7005,N_7006);
nor U7335 (N_7335,N_6985,N_6912);
nor U7336 (N_7336,N_6960,N_6909);
xnor U7337 (N_7337,N_7018,N_6910);
and U7338 (N_7338,N_7037,N_6913);
nand U7339 (N_7339,N_6937,N_7086);
and U7340 (N_7340,N_7057,N_7128);
and U7341 (N_7341,N_6927,N_7180);
nor U7342 (N_7342,N_7027,N_7124);
and U7343 (N_7343,N_6956,N_7158);
xor U7344 (N_7344,N_6929,N_7113);
or U7345 (N_7345,N_6971,N_7007);
and U7346 (N_7346,N_7067,N_7026);
and U7347 (N_7347,N_7050,N_7195);
nor U7348 (N_7348,N_6975,N_6947);
nand U7349 (N_7349,N_6993,N_6992);
xor U7350 (N_7350,N_6992,N_6986);
nand U7351 (N_7351,N_7002,N_6947);
nand U7352 (N_7352,N_7096,N_7091);
xnor U7353 (N_7353,N_6976,N_7190);
nand U7354 (N_7354,N_7147,N_7155);
xor U7355 (N_7355,N_7048,N_7072);
or U7356 (N_7356,N_6927,N_6980);
and U7357 (N_7357,N_7106,N_7179);
or U7358 (N_7358,N_7057,N_7035);
or U7359 (N_7359,N_6946,N_7024);
xor U7360 (N_7360,N_7176,N_6990);
nand U7361 (N_7361,N_7171,N_7124);
and U7362 (N_7362,N_6931,N_7061);
nor U7363 (N_7363,N_7086,N_7163);
nand U7364 (N_7364,N_7066,N_7084);
and U7365 (N_7365,N_6936,N_6994);
nand U7366 (N_7366,N_7197,N_7148);
and U7367 (N_7367,N_7182,N_7151);
xnor U7368 (N_7368,N_7136,N_6949);
nor U7369 (N_7369,N_7168,N_7034);
and U7370 (N_7370,N_7001,N_7081);
nor U7371 (N_7371,N_7056,N_7175);
nand U7372 (N_7372,N_7039,N_6925);
nand U7373 (N_7373,N_7047,N_6957);
or U7374 (N_7374,N_7199,N_7047);
nor U7375 (N_7375,N_7009,N_6975);
nor U7376 (N_7376,N_7181,N_7120);
xnor U7377 (N_7377,N_6952,N_7166);
nand U7378 (N_7378,N_6908,N_6982);
nand U7379 (N_7379,N_7087,N_7086);
xor U7380 (N_7380,N_7038,N_6988);
or U7381 (N_7381,N_7132,N_6962);
or U7382 (N_7382,N_7079,N_7173);
or U7383 (N_7383,N_7190,N_7108);
xnor U7384 (N_7384,N_7189,N_7173);
and U7385 (N_7385,N_7173,N_6980);
nor U7386 (N_7386,N_7042,N_6977);
nor U7387 (N_7387,N_7003,N_6952);
and U7388 (N_7388,N_6962,N_6912);
nor U7389 (N_7389,N_7123,N_6954);
nor U7390 (N_7390,N_7011,N_7089);
nand U7391 (N_7391,N_7001,N_7018);
or U7392 (N_7392,N_7150,N_7124);
or U7393 (N_7393,N_6918,N_7064);
or U7394 (N_7394,N_7004,N_7148);
or U7395 (N_7395,N_6911,N_7055);
and U7396 (N_7396,N_6966,N_7032);
nand U7397 (N_7397,N_7150,N_6987);
or U7398 (N_7398,N_6967,N_7006);
and U7399 (N_7399,N_6908,N_7081);
nand U7400 (N_7400,N_7152,N_7077);
xor U7401 (N_7401,N_7000,N_7101);
and U7402 (N_7402,N_6983,N_7061);
xnor U7403 (N_7403,N_7059,N_7020);
nor U7404 (N_7404,N_7070,N_6923);
or U7405 (N_7405,N_7129,N_6906);
nand U7406 (N_7406,N_7086,N_6966);
or U7407 (N_7407,N_7110,N_7092);
and U7408 (N_7408,N_7077,N_6943);
xor U7409 (N_7409,N_7039,N_7029);
nand U7410 (N_7410,N_7069,N_7126);
nor U7411 (N_7411,N_7182,N_7088);
xor U7412 (N_7412,N_7012,N_7134);
and U7413 (N_7413,N_7136,N_7155);
nand U7414 (N_7414,N_7168,N_7153);
nand U7415 (N_7415,N_6963,N_6902);
xnor U7416 (N_7416,N_7088,N_7194);
nor U7417 (N_7417,N_7182,N_7032);
nor U7418 (N_7418,N_6901,N_7152);
nor U7419 (N_7419,N_7059,N_7171);
and U7420 (N_7420,N_6987,N_7148);
xnor U7421 (N_7421,N_6917,N_7033);
xnor U7422 (N_7422,N_6957,N_7172);
or U7423 (N_7423,N_7137,N_7088);
xor U7424 (N_7424,N_7176,N_7057);
xnor U7425 (N_7425,N_7170,N_6999);
and U7426 (N_7426,N_7199,N_7028);
and U7427 (N_7427,N_7018,N_7149);
and U7428 (N_7428,N_6984,N_7005);
nor U7429 (N_7429,N_7087,N_7164);
or U7430 (N_7430,N_6948,N_7125);
nor U7431 (N_7431,N_7140,N_7182);
or U7432 (N_7432,N_7160,N_6935);
and U7433 (N_7433,N_7050,N_7108);
nand U7434 (N_7434,N_6924,N_7146);
and U7435 (N_7435,N_7127,N_7166);
nor U7436 (N_7436,N_6956,N_7177);
nand U7437 (N_7437,N_7157,N_7005);
or U7438 (N_7438,N_7093,N_7016);
xor U7439 (N_7439,N_6946,N_6971);
xnor U7440 (N_7440,N_7045,N_7194);
xnor U7441 (N_7441,N_7029,N_7185);
nand U7442 (N_7442,N_7114,N_6996);
xnor U7443 (N_7443,N_6945,N_7061);
xor U7444 (N_7444,N_7195,N_7182);
and U7445 (N_7445,N_6925,N_7010);
nand U7446 (N_7446,N_6951,N_7034);
nor U7447 (N_7447,N_7143,N_7114);
or U7448 (N_7448,N_6999,N_7182);
nand U7449 (N_7449,N_7005,N_6990);
xor U7450 (N_7450,N_7118,N_6910);
nor U7451 (N_7451,N_6982,N_6967);
nor U7452 (N_7452,N_7089,N_6955);
xor U7453 (N_7453,N_6915,N_6923);
nor U7454 (N_7454,N_6931,N_7007);
or U7455 (N_7455,N_7190,N_6943);
xnor U7456 (N_7456,N_6924,N_7010);
nor U7457 (N_7457,N_7147,N_7041);
and U7458 (N_7458,N_7173,N_7130);
nand U7459 (N_7459,N_7093,N_7190);
and U7460 (N_7460,N_7024,N_7196);
and U7461 (N_7461,N_7152,N_7012);
and U7462 (N_7462,N_7007,N_6994);
nand U7463 (N_7463,N_7186,N_7100);
nor U7464 (N_7464,N_7153,N_6947);
nand U7465 (N_7465,N_7188,N_7069);
xor U7466 (N_7466,N_6904,N_7189);
xnor U7467 (N_7467,N_7030,N_7043);
xnor U7468 (N_7468,N_7135,N_7065);
or U7469 (N_7469,N_6970,N_7187);
xor U7470 (N_7470,N_7153,N_7191);
and U7471 (N_7471,N_7135,N_6909);
xor U7472 (N_7472,N_7162,N_6980);
and U7473 (N_7473,N_7154,N_7134);
xor U7474 (N_7474,N_6940,N_7176);
nand U7475 (N_7475,N_7171,N_7028);
or U7476 (N_7476,N_7068,N_7064);
or U7477 (N_7477,N_6981,N_7154);
nor U7478 (N_7478,N_6951,N_7108);
xor U7479 (N_7479,N_7133,N_7158);
nor U7480 (N_7480,N_7014,N_6958);
nor U7481 (N_7481,N_6980,N_7081);
xor U7482 (N_7482,N_7014,N_7169);
nor U7483 (N_7483,N_6926,N_7180);
nor U7484 (N_7484,N_6972,N_7145);
xor U7485 (N_7485,N_7128,N_6986);
nor U7486 (N_7486,N_6962,N_7111);
or U7487 (N_7487,N_7156,N_7016);
nand U7488 (N_7488,N_6992,N_7106);
xor U7489 (N_7489,N_7104,N_7074);
xnor U7490 (N_7490,N_6919,N_7091);
nand U7491 (N_7491,N_7085,N_7121);
or U7492 (N_7492,N_7053,N_7119);
xnor U7493 (N_7493,N_7149,N_6951);
or U7494 (N_7494,N_6907,N_6986);
and U7495 (N_7495,N_7026,N_7157);
xnor U7496 (N_7496,N_7178,N_7010);
or U7497 (N_7497,N_7102,N_7174);
nand U7498 (N_7498,N_7134,N_6932);
xnor U7499 (N_7499,N_7054,N_7174);
and U7500 (N_7500,N_7390,N_7445);
nor U7501 (N_7501,N_7464,N_7385);
nand U7502 (N_7502,N_7405,N_7299);
or U7503 (N_7503,N_7319,N_7212);
xor U7504 (N_7504,N_7288,N_7267);
nor U7505 (N_7505,N_7304,N_7396);
nor U7506 (N_7506,N_7266,N_7347);
nand U7507 (N_7507,N_7485,N_7250);
xor U7508 (N_7508,N_7362,N_7407);
xor U7509 (N_7509,N_7491,N_7303);
xor U7510 (N_7510,N_7412,N_7322);
nor U7511 (N_7511,N_7400,N_7384);
nor U7512 (N_7512,N_7290,N_7348);
or U7513 (N_7513,N_7406,N_7325);
xor U7514 (N_7514,N_7339,N_7298);
and U7515 (N_7515,N_7242,N_7459);
nand U7516 (N_7516,N_7375,N_7440);
or U7517 (N_7517,N_7338,N_7414);
nand U7518 (N_7518,N_7247,N_7429);
nor U7519 (N_7519,N_7286,N_7311);
and U7520 (N_7520,N_7399,N_7230);
xnor U7521 (N_7521,N_7283,N_7248);
or U7522 (N_7522,N_7425,N_7437);
nor U7523 (N_7523,N_7460,N_7474);
nand U7524 (N_7524,N_7222,N_7486);
and U7525 (N_7525,N_7293,N_7203);
and U7526 (N_7526,N_7418,N_7371);
or U7527 (N_7527,N_7234,N_7350);
and U7528 (N_7528,N_7449,N_7229);
or U7529 (N_7529,N_7481,N_7423);
and U7530 (N_7530,N_7421,N_7470);
or U7531 (N_7531,N_7228,N_7336);
nor U7532 (N_7532,N_7469,N_7422);
nand U7533 (N_7533,N_7209,N_7356);
nor U7534 (N_7534,N_7271,N_7458);
nor U7535 (N_7535,N_7296,N_7368);
nand U7536 (N_7536,N_7301,N_7416);
or U7537 (N_7537,N_7492,N_7258);
xor U7538 (N_7538,N_7237,N_7204);
and U7539 (N_7539,N_7346,N_7243);
nand U7540 (N_7540,N_7233,N_7314);
xor U7541 (N_7541,N_7334,N_7330);
and U7542 (N_7542,N_7211,N_7285);
or U7543 (N_7543,N_7241,N_7223);
or U7544 (N_7544,N_7370,N_7224);
and U7545 (N_7545,N_7324,N_7215);
or U7546 (N_7546,N_7256,N_7484);
nor U7547 (N_7547,N_7395,N_7349);
or U7548 (N_7548,N_7456,N_7238);
nor U7549 (N_7549,N_7376,N_7318);
nand U7550 (N_7550,N_7240,N_7309);
xor U7551 (N_7551,N_7262,N_7333);
nand U7552 (N_7552,N_7292,N_7254);
or U7553 (N_7553,N_7214,N_7327);
nor U7554 (N_7554,N_7315,N_7202);
or U7555 (N_7555,N_7381,N_7265);
nor U7556 (N_7556,N_7363,N_7232);
nor U7557 (N_7557,N_7317,N_7221);
xnor U7558 (N_7558,N_7461,N_7270);
xnor U7559 (N_7559,N_7496,N_7446);
or U7560 (N_7560,N_7306,N_7393);
nand U7561 (N_7561,N_7210,N_7320);
nor U7562 (N_7562,N_7340,N_7435);
or U7563 (N_7563,N_7480,N_7373);
and U7564 (N_7564,N_7417,N_7443);
xnor U7565 (N_7565,N_7361,N_7244);
nor U7566 (N_7566,N_7217,N_7335);
and U7567 (N_7567,N_7201,N_7436);
nand U7568 (N_7568,N_7454,N_7386);
and U7569 (N_7569,N_7379,N_7402);
nor U7570 (N_7570,N_7276,N_7216);
nand U7571 (N_7571,N_7354,N_7207);
or U7572 (N_7572,N_7366,N_7358);
nand U7573 (N_7573,N_7415,N_7409);
or U7574 (N_7574,N_7245,N_7208);
or U7575 (N_7575,N_7394,N_7382);
nand U7576 (N_7576,N_7352,N_7428);
or U7577 (N_7577,N_7226,N_7444);
nand U7578 (N_7578,N_7482,N_7323);
xnor U7579 (N_7579,N_7367,N_7355);
nor U7580 (N_7580,N_7275,N_7404);
nand U7581 (N_7581,N_7453,N_7391);
and U7582 (N_7582,N_7475,N_7377);
or U7583 (N_7583,N_7497,N_7277);
nor U7584 (N_7584,N_7280,N_7472);
and U7585 (N_7585,N_7259,N_7269);
nor U7586 (N_7586,N_7434,N_7380);
and U7587 (N_7587,N_7452,N_7344);
or U7588 (N_7588,N_7438,N_7427);
nand U7589 (N_7589,N_7463,N_7307);
nor U7590 (N_7590,N_7357,N_7420);
nor U7591 (N_7591,N_7246,N_7432);
nand U7592 (N_7592,N_7383,N_7279);
xnor U7593 (N_7593,N_7433,N_7466);
or U7594 (N_7594,N_7291,N_7389);
or U7595 (N_7595,N_7424,N_7441);
nand U7596 (N_7596,N_7353,N_7345);
xor U7597 (N_7597,N_7295,N_7220);
xnor U7598 (N_7598,N_7494,N_7479);
nand U7599 (N_7599,N_7200,N_7448);
and U7600 (N_7600,N_7312,N_7272);
nor U7601 (N_7601,N_7455,N_7257);
xor U7602 (N_7602,N_7251,N_7467);
or U7603 (N_7603,N_7498,N_7305);
nand U7604 (N_7604,N_7289,N_7351);
xnor U7605 (N_7605,N_7342,N_7478);
nand U7606 (N_7606,N_7476,N_7457);
and U7607 (N_7607,N_7468,N_7426);
or U7608 (N_7608,N_7218,N_7489);
nor U7609 (N_7609,N_7249,N_7410);
or U7610 (N_7610,N_7392,N_7235);
or U7611 (N_7611,N_7326,N_7281);
and U7612 (N_7612,N_7236,N_7268);
xor U7613 (N_7613,N_7430,N_7493);
xor U7614 (N_7614,N_7343,N_7450);
xor U7615 (N_7615,N_7419,N_7260);
or U7616 (N_7616,N_7387,N_7231);
nor U7617 (N_7617,N_7364,N_7282);
or U7618 (N_7618,N_7451,N_7499);
nor U7619 (N_7619,N_7321,N_7462);
nand U7620 (N_7620,N_7300,N_7439);
nor U7621 (N_7621,N_7227,N_7365);
nor U7622 (N_7622,N_7471,N_7316);
xor U7623 (N_7623,N_7488,N_7388);
and U7624 (N_7624,N_7255,N_7413);
or U7625 (N_7625,N_7397,N_7369);
nand U7626 (N_7626,N_7297,N_7341);
or U7627 (N_7627,N_7213,N_7329);
and U7628 (N_7628,N_7313,N_7378);
nand U7629 (N_7629,N_7274,N_7225);
nor U7630 (N_7630,N_7447,N_7239);
and U7631 (N_7631,N_7264,N_7442);
or U7632 (N_7632,N_7483,N_7205);
and U7633 (N_7633,N_7261,N_7294);
xor U7634 (N_7634,N_7408,N_7253);
nor U7635 (N_7635,N_7278,N_7331);
or U7636 (N_7636,N_7332,N_7328);
nor U7637 (N_7637,N_7398,N_7273);
nor U7638 (N_7638,N_7495,N_7263);
nand U7639 (N_7639,N_7490,N_7477);
xor U7640 (N_7640,N_7465,N_7487);
nand U7641 (N_7641,N_7473,N_7337);
and U7642 (N_7642,N_7252,N_7287);
xnor U7643 (N_7643,N_7219,N_7360);
xor U7644 (N_7644,N_7374,N_7308);
and U7645 (N_7645,N_7401,N_7302);
xnor U7646 (N_7646,N_7284,N_7411);
nand U7647 (N_7647,N_7310,N_7359);
nand U7648 (N_7648,N_7372,N_7431);
nor U7649 (N_7649,N_7403,N_7206);
nand U7650 (N_7650,N_7218,N_7419);
nand U7651 (N_7651,N_7444,N_7237);
xnor U7652 (N_7652,N_7208,N_7313);
or U7653 (N_7653,N_7236,N_7479);
and U7654 (N_7654,N_7263,N_7406);
and U7655 (N_7655,N_7412,N_7274);
nor U7656 (N_7656,N_7418,N_7248);
or U7657 (N_7657,N_7381,N_7444);
nand U7658 (N_7658,N_7413,N_7313);
xnor U7659 (N_7659,N_7225,N_7476);
nand U7660 (N_7660,N_7448,N_7398);
or U7661 (N_7661,N_7464,N_7301);
or U7662 (N_7662,N_7253,N_7357);
nor U7663 (N_7663,N_7442,N_7209);
nand U7664 (N_7664,N_7437,N_7323);
nand U7665 (N_7665,N_7280,N_7426);
or U7666 (N_7666,N_7277,N_7468);
nor U7667 (N_7667,N_7284,N_7378);
or U7668 (N_7668,N_7222,N_7353);
or U7669 (N_7669,N_7426,N_7425);
and U7670 (N_7670,N_7225,N_7341);
or U7671 (N_7671,N_7417,N_7255);
nor U7672 (N_7672,N_7284,N_7317);
or U7673 (N_7673,N_7228,N_7490);
nor U7674 (N_7674,N_7317,N_7380);
nor U7675 (N_7675,N_7214,N_7279);
or U7676 (N_7676,N_7432,N_7327);
nor U7677 (N_7677,N_7214,N_7446);
xor U7678 (N_7678,N_7203,N_7213);
nor U7679 (N_7679,N_7475,N_7205);
nand U7680 (N_7680,N_7203,N_7404);
and U7681 (N_7681,N_7404,N_7337);
xnor U7682 (N_7682,N_7314,N_7470);
nand U7683 (N_7683,N_7499,N_7493);
xor U7684 (N_7684,N_7412,N_7286);
nand U7685 (N_7685,N_7362,N_7329);
nand U7686 (N_7686,N_7352,N_7404);
or U7687 (N_7687,N_7494,N_7234);
xnor U7688 (N_7688,N_7451,N_7215);
nand U7689 (N_7689,N_7482,N_7205);
and U7690 (N_7690,N_7481,N_7205);
xor U7691 (N_7691,N_7408,N_7334);
or U7692 (N_7692,N_7202,N_7289);
xnor U7693 (N_7693,N_7299,N_7221);
xor U7694 (N_7694,N_7461,N_7462);
nand U7695 (N_7695,N_7417,N_7205);
and U7696 (N_7696,N_7380,N_7397);
and U7697 (N_7697,N_7397,N_7421);
or U7698 (N_7698,N_7297,N_7453);
and U7699 (N_7699,N_7302,N_7264);
and U7700 (N_7700,N_7348,N_7207);
and U7701 (N_7701,N_7425,N_7382);
xnor U7702 (N_7702,N_7252,N_7302);
or U7703 (N_7703,N_7475,N_7254);
or U7704 (N_7704,N_7316,N_7346);
or U7705 (N_7705,N_7444,N_7330);
or U7706 (N_7706,N_7454,N_7447);
and U7707 (N_7707,N_7452,N_7412);
xnor U7708 (N_7708,N_7285,N_7218);
nor U7709 (N_7709,N_7460,N_7252);
xor U7710 (N_7710,N_7401,N_7348);
nor U7711 (N_7711,N_7297,N_7409);
and U7712 (N_7712,N_7439,N_7292);
or U7713 (N_7713,N_7343,N_7344);
or U7714 (N_7714,N_7320,N_7464);
nand U7715 (N_7715,N_7387,N_7407);
nor U7716 (N_7716,N_7235,N_7438);
nand U7717 (N_7717,N_7288,N_7305);
or U7718 (N_7718,N_7439,N_7326);
and U7719 (N_7719,N_7344,N_7253);
nor U7720 (N_7720,N_7301,N_7296);
and U7721 (N_7721,N_7312,N_7445);
nor U7722 (N_7722,N_7404,N_7251);
and U7723 (N_7723,N_7214,N_7321);
nor U7724 (N_7724,N_7231,N_7233);
or U7725 (N_7725,N_7249,N_7387);
nand U7726 (N_7726,N_7404,N_7262);
nand U7727 (N_7727,N_7307,N_7289);
xor U7728 (N_7728,N_7382,N_7489);
nand U7729 (N_7729,N_7226,N_7207);
xnor U7730 (N_7730,N_7382,N_7436);
nor U7731 (N_7731,N_7239,N_7467);
xnor U7732 (N_7732,N_7221,N_7440);
nand U7733 (N_7733,N_7292,N_7296);
xnor U7734 (N_7734,N_7452,N_7399);
nor U7735 (N_7735,N_7315,N_7337);
nand U7736 (N_7736,N_7245,N_7453);
nand U7737 (N_7737,N_7421,N_7231);
nand U7738 (N_7738,N_7468,N_7455);
or U7739 (N_7739,N_7444,N_7249);
nand U7740 (N_7740,N_7402,N_7451);
and U7741 (N_7741,N_7372,N_7305);
or U7742 (N_7742,N_7433,N_7440);
and U7743 (N_7743,N_7477,N_7310);
nor U7744 (N_7744,N_7231,N_7211);
or U7745 (N_7745,N_7497,N_7301);
nor U7746 (N_7746,N_7334,N_7383);
nand U7747 (N_7747,N_7402,N_7382);
nand U7748 (N_7748,N_7200,N_7428);
xnor U7749 (N_7749,N_7485,N_7355);
and U7750 (N_7750,N_7369,N_7311);
xnor U7751 (N_7751,N_7420,N_7261);
xor U7752 (N_7752,N_7229,N_7322);
and U7753 (N_7753,N_7346,N_7217);
and U7754 (N_7754,N_7266,N_7206);
or U7755 (N_7755,N_7264,N_7270);
or U7756 (N_7756,N_7497,N_7219);
nor U7757 (N_7757,N_7329,N_7490);
nand U7758 (N_7758,N_7416,N_7307);
or U7759 (N_7759,N_7467,N_7340);
or U7760 (N_7760,N_7289,N_7426);
nor U7761 (N_7761,N_7203,N_7263);
nor U7762 (N_7762,N_7360,N_7229);
nand U7763 (N_7763,N_7459,N_7310);
nor U7764 (N_7764,N_7379,N_7290);
and U7765 (N_7765,N_7272,N_7247);
nand U7766 (N_7766,N_7396,N_7332);
nor U7767 (N_7767,N_7246,N_7341);
xor U7768 (N_7768,N_7377,N_7293);
and U7769 (N_7769,N_7212,N_7268);
nand U7770 (N_7770,N_7406,N_7327);
or U7771 (N_7771,N_7226,N_7333);
xor U7772 (N_7772,N_7467,N_7356);
xnor U7773 (N_7773,N_7485,N_7282);
or U7774 (N_7774,N_7347,N_7471);
and U7775 (N_7775,N_7418,N_7305);
or U7776 (N_7776,N_7390,N_7404);
nand U7777 (N_7777,N_7322,N_7454);
and U7778 (N_7778,N_7342,N_7385);
nand U7779 (N_7779,N_7253,N_7270);
nand U7780 (N_7780,N_7247,N_7447);
xor U7781 (N_7781,N_7285,N_7368);
or U7782 (N_7782,N_7483,N_7425);
nor U7783 (N_7783,N_7321,N_7375);
nor U7784 (N_7784,N_7329,N_7401);
nor U7785 (N_7785,N_7391,N_7467);
nor U7786 (N_7786,N_7454,N_7286);
or U7787 (N_7787,N_7355,N_7293);
xor U7788 (N_7788,N_7301,N_7282);
xor U7789 (N_7789,N_7304,N_7480);
and U7790 (N_7790,N_7477,N_7352);
or U7791 (N_7791,N_7353,N_7226);
and U7792 (N_7792,N_7393,N_7492);
and U7793 (N_7793,N_7210,N_7206);
or U7794 (N_7794,N_7254,N_7204);
and U7795 (N_7795,N_7280,N_7263);
xnor U7796 (N_7796,N_7250,N_7387);
nand U7797 (N_7797,N_7482,N_7467);
xor U7798 (N_7798,N_7251,N_7267);
nor U7799 (N_7799,N_7404,N_7430);
nand U7800 (N_7800,N_7674,N_7699);
nand U7801 (N_7801,N_7543,N_7647);
or U7802 (N_7802,N_7777,N_7612);
and U7803 (N_7803,N_7741,N_7602);
or U7804 (N_7804,N_7693,N_7770);
nor U7805 (N_7805,N_7512,N_7702);
nor U7806 (N_7806,N_7521,N_7724);
or U7807 (N_7807,N_7610,N_7691);
and U7808 (N_7808,N_7781,N_7719);
xor U7809 (N_7809,N_7522,N_7628);
xnor U7810 (N_7810,N_7577,N_7796);
nand U7811 (N_7811,N_7553,N_7574);
or U7812 (N_7812,N_7626,N_7586);
nand U7813 (N_7813,N_7725,N_7508);
nand U7814 (N_7814,N_7726,N_7785);
nand U7815 (N_7815,N_7797,N_7642);
and U7816 (N_7816,N_7709,N_7619);
xnor U7817 (N_7817,N_7609,N_7551);
and U7818 (N_7818,N_7651,N_7523);
nor U7819 (N_7819,N_7767,N_7664);
xor U7820 (N_7820,N_7539,N_7654);
nand U7821 (N_7821,N_7511,N_7742);
xor U7822 (N_7822,N_7547,N_7650);
or U7823 (N_7823,N_7740,N_7762);
nor U7824 (N_7824,N_7698,N_7746);
xnor U7825 (N_7825,N_7751,N_7617);
xor U7826 (N_7826,N_7795,N_7774);
nand U7827 (N_7827,N_7604,N_7581);
nor U7828 (N_7828,N_7528,N_7570);
xor U7829 (N_7829,N_7745,N_7618);
nand U7830 (N_7830,N_7685,N_7768);
xor U7831 (N_7831,N_7713,N_7576);
nor U7832 (N_7832,N_7683,N_7684);
or U7833 (N_7833,N_7678,N_7787);
nand U7834 (N_7834,N_7501,N_7600);
and U7835 (N_7835,N_7749,N_7747);
xnor U7836 (N_7836,N_7660,N_7799);
or U7837 (N_7837,N_7504,N_7648);
and U7838 (N_7838,N_7598,N_7766);
and U7839 (N_7839,N_7603,N_7616);
nor U7840 (N_7840,N_7730,N_7505);
nand U7841 (N_7841,N_7765,N_7564);
or U7842 (N_7842,N_7588,N_7595);
and U7843 (N_7843,N_7646,N_7593);
and U7844 (N_7844,N_7665,N_7686);
nand U7845 (N_7845,N_7780,N_7771);
and U7846 (N_7846,N_7667,N_7644);
or U7847 (N_7847,N_7591,N_7527);
nand U7848 (N_7848,N_7670,N_7723);
nand U7849 (N_7849,N_7736,N_7546);
nand U7850 (N_7850,N_7769,N_7682);
nor U7851 (N_7851,N_7587,N_7605);
nor U7852 (N_7852,N_7607,N_7530);
nand U7853 (N_7853,N_7657,N_7571);
or U7854 (N_7854,N_7789,N_7714);
nor U7855 (N_7855,N_7500,N_7566);
xnor U7856 (N_7856,N_7542,N_7629);
or U7857 (N_7857,N_7583,N_7668);
nand U7858 (N_7858,N_7623,N_7791);
nand U7859 (N_7859,N_7743,N_7611);
and U7860 (N_7860,N_7703,N_7734);
nand U7861 (N_7861,N_7558,N_7753);
nand U7862 (N_7862,N_7666,N_7545);
nor U7863 (N_7863,N_7639,N_7507);
xor U7864 (N_7864,N_7534,N_7782);
or U7865 (N_7865,N_7536,N_7559);
and U7866 (N_7866,N_7631,N_7625);
xnor U7867 (N_7867,N_7537,N_7705);
nor U7868 (N_7868,N_7589,N_7590);
nand U7869 (N_7869,N_7689,N_7656);
nand U7870 (N_7870,N_7649,N_7790);
nor U7871 (N_7871,N_7722,N_7557);
or U7872 (N_7872,N_7517,N_7707);
or U7873 (N_7873,N_7652,N_7622);
nor U7874 (N_7874,N_7706,N_7638);
nor U7875 (N_7875,N_7541,N_7681);
nor U7876 (N_7876,N_7535,N_7721);
or U7877 (N_7877,N_7750,N_7712);
and U7878 (N_7878,N_7503,N_7786);
or U7879 (N_7879,N_7662,N_7748);
or U7880 (N_7880,N_7716,N_7584);
xnor U7881 (N_7881,N_7636,N_7548);
nor U7882 (N_7882,N_7597,N_7761);
xor U7883 (N_7883,N_7759,N_7510);
nand U7884 (N_7884,N_7717,N_7733);
and U7885 (N_7885,N_7515,N_7737);
nand U7886 (N_7886,N_7538,N_7655);
or U7887 (N_7887,N_7540,N_7502);
nand U7888 (N_7888,N_7727,N_7735);
xor U7889 (N_7889,N_7514,N_7578);
nor U7890 (N_7890,N_7739,N_7690);
or U7891 (N_7891,N_7544,N_7701);
and U7892 (N_7892,N_7579,N_7634);
nand U7893 (N_7893,N_7653,N_7692);
or U7894 (N_7894,N_7568,N_7715);
and U7895 (N_7895,N_7760,N_7732);
nor U7896 (N_7896,N_7758,N_7561);
xor U7897 (N_7897,N_7696,N_7755);
or U7898 (N_7898,N_7718,N_7560);
or U7899 (N_7899,N_7757,N_7720);
nor U7900 (N_7900,N_7531,N_7632);
nor U7901 (N_7901,N_7596,N_7635);
nor U7902 (N_7902,N_7599,N_7792);
and U7903 (N_7903,N_7509,N_7779);
xor U7904 (N_7904,N_7763,N_7524);
nor U7905 (N_7905,N_7645,N_7513);
nor U7906 (N_7906,N_7784,N_7567);
nand U7907 (N_7907,N_7679,N_7669);
and U7908 (N_7908,N_7711,N_7710);
xnor U7909 (N_7909,N_7529,N_7687);
and U7910 (N_7910,N_7633,N_7778);
and U7911 (N_7911,N_7671,N_7694);
nor U7912 (N_7912,N_7794,N_7738);
and U7913 (N_7913,N_7637,N_7752);
or U7914 (N_7914,N_7764,N_7573);
or U7915 (N_7915,N_7756,N_7621);
and U7916 (N_7916,N_7614,N_7673);
and U7917 (N_7917,N_7516,N_7549);
xnor U7918 (N_7918,N_7606,N_7798);
nand U7919 (N_7919,N_7556,N_7641);
or U7920 (N_7920,N_7708,N_7555);
nor U7921 (N_7921,N_7772,N_7554);
nor U7922 (N_7922,N_7562,N_7608);
xnor U7923 (N_7923,N_7601,N_7569);
or U7924 (N_7924,N_7533,N_7615);
or U7925 (N_7925,N_7663,N_7520);
xnor U7926 (N_7926,N_7695,N_7697);
or U7927 (N_7927,N_7580,N_7565);
and U7928 (N_7928,N_7677,N_7518);
and U7929 (N_7929,N_7506,N_7563);
or U7930 (N_7930,N_7675,N_7793);
xor U7931 (N_7931,N_7525,N_7526);
nor U7932 (N_7932,N_7728,N_7630);
and U7933 (N_7933,N_7704,N_7700);
or U7934 (N_7934,N_7744,N_7613);
nand U7935 (N_7935,N_7688,N_7627);
nor U7936 (N_7936,N_7582,N_7572);
nor U7937 (N_7937,N_7773,N_7672);
nor U7938 (N_7938,N_7658,N_7640);
nand U7939 (N_7939,N_7754,N_7532);
nor U7940 (N_7940,N_7592,N_7788);
xnor U7941 (N_7941,N_7550,N_7643);
nor U7942 (N_7942,N_7676,N_7620);
nor U7943 (N_7943,N_7585,N_7659);
nand U7944 (N_7944,N_7783,N_7775);
nand U7945 (N_7945,N_7776,N_7729);
nor U7946 (N_7946,N_7552,N_7594);
nand U7947 (N_7947,N_7731,N_7624);
or U7948 (N_7948,N_7680,N_7575);
nor U7949 (N_7949,N_7661,N_7519);
xor U7950 (N_7950,N_7759,N_7746);
and U7951 (N_7951,N_7674,N_7737);
nor U7952 (N_7952,N_7500,N_7502);
xnor U7953 (N_7953,N_7535,N_7665);
nor U7954 (N_7954,N_7699,N_7579);
nand U7955 (N_7955,N_7505,N_7790);
or U7956 (N_7956,N_7652,N_7547);
xnor U7957 (N_7957,N_7682,N_7520);
nor U7958 (N_7958,N_7558,N_7754);
nor U7959 (N_7959,N_7697,N_7756);
or U7960 (N_7960,N_7547,N_7756);
xnor U7961 (N_7961,N_7672,N_7762);
nand U7962 (N_7962,N_7787,N_7672);
nor U7963 (N_7963,N_7697,N_7712);
xor U7964 (N_7964,N_7610,N_7719);
nand U7965 (N_7965,N_7502,N_7769);
nand U7966 (N_7966,N_7662,N_7592);
nand U7967 (N_7967,N_7634,N_7791);
xnor U7968 (N_7968,N_7646,N_7587);
and U7969 (N_7969,N_7726,N_7513);
and U7970 (N_7970,N_7511,N_7521);
and U7971 (N_7971,N_7604,N_7642);
nor U7972 (N_7972,N_7766,N_7733);
and U7973 (N_7973,N_7778,N_7656);
or U7974 (N_7974,N_7597,N_7620);
nor U7975 (N_7975,N_7658,N_7514);
and U7976 (N_7976,N_7540,N_7723);
xor U7977 (N_7977,N_7780,N_7506);
and U7978 (N_7978,N_7777,N_7537);
or U7979 (N_7979,N_7618,N_7541);
nor U7980 (N_7980,N_7529,N_7713);
and U7981 (N_7981,N_7700,N_7566);
and U7982 (N_7982,N_7725,N_7559);
xnor U7983 (N_7983,N_7757,N_7558);
nand U7984 (N_7984,N_7742,N_7560);
xor U7985 (N_7985,N_7783,N_7590);
nor U7986 (N_7986,N_7646,N_7674);
or U7987 (N_7987,N_7736,N_7579);
or U7988 (N_7988,N_7782,N_7746);
nor U7989 (N_7989,N_7640,N_7730);
nand U7990 (N_7990,N_7702,N_7672);
nor U7991 (N_7991,N_7548,N_7516);
nand U7992 (N_7992,N_7575,N_7749);
nand U7993 (N_7993,N_7527,N_7662);
or U7994 (N_7994,N_7695,N_7785);
nor U7995 (N_7995,N_7746,N_7508);
or U7996 (N_7996,N_7524,N_7770);
nand U7997 (N_7997,N_7581,N_7792);
and U7998 (N_7998,N_7708,N_7719);
nand U7999 (N_7999,N_7588,N_7683);
xnor U8000 (N_8000,N_7580,N_7743);
xor U8001 (N_8001,N_7598,N_7660);
xnor U8002 (N_8002,N_7579,N_7663);
nor U8003 (N_8003,N_7523,N_7703);
or U8004 (N_8004,N_7649,N_7721);
nor U8005 (N_8005,N_7532,N_7684);
nand U8006 (N_8006,N_7595,N_7567);
nor U8007 (N_8007,N_7601,N_7509);
nand U8008 (N_8008,N_7520,N_7522);
xnor U8009 (N_8009,N_7724,N_7645);
nand U8010 (N_8010,N_7627,N_7666);
nor U8011 (N_8011,N_7552,N_7674);
and U8012 (N_8012,N_7583,N_7573);
or U8013 (N_8013,N_7584,N_7759);
nand U8014 (N_8014,N_7553,N_7728);
nand U8015 (N_8015,N_7519,N_7758);
and U8016 (N_8016,N_7553,N_7578);
nor U8017 (N_8017,N_7547,N_7749);
and U8018 (N_8018,N_7666,N_7704);
nor U8019 (N_8019,N_7734,N_7694);
xor U8020 (N_8020,N_7798,N_7698);
and U8021 (N_8021,N_7686,N_7617);
and U8022 (N_8022,N_7611,N_7520);
xor U8023 (N_8023,N_7563,N_7540);
xor U8024 (N_8024,N_7787,N_7737);
nor U8025 (N_8025,N_7637,N_7527);
nand U8026 (N_8026,N_7686,N_7630);
nand U8027 (N_8027,N_7579,N_7571);
nor U8028 (N_8028,N_7656,N_7756);
and U8029 (N_8029,N_7649,N_7525);
nand U8030 (N_8030,N_7711,N_7749);
and U8031 (N_8031,N_7704,N_7791);
xor U8032 (N_8032,N_7725,N_7728);
nor U8033 (N_8033,N_7629,N_7728);
nor U8034 (N_8034,N_7667,N_7786);
nand U8035 (N_8035,N_7550,N_7651);
and U8036 (N_8036,N_7778,N_7713);
nor U8037 (N_8037,N_7755,N_7678);
or U8038 (N_8038,N_7707,N_7606);
or U8039 (N_8039,N_7595,N_7693);
and U8040 (N_8040,N_7550,N_7570);
nor U8041 (N_8041,N_7653,N_7616);
or U8042 (N_8042,N_7764,N_7751);
and U8043 (N_8043,N_7788,N_7766);
nand U8044 (N_8044,N_7614,N_7675);
xnor U8045 (N_8045,N_7575,N_7558);
xor U8046 (N_8046,N_7797,N_7647);
xnor U8047 (N_8047,N_7563,N_7536);
or U8048 (N_8048,N_7563,N_7623);
xnor U8049 (N_8049,N_7513,N_7668);
xnor U8050 (N_8050,N_7738,N_7718);
or U8051 (N_8051,N_7579,N_7761);
nor U8052 (N_8052,N_7535,N_7637);
nor U8053 (N_8053,N_7629,N_7548);
nand U8054 (N_8054,N_7601,N_7759);
and U8055 (N_8055,N_7507,N_7710);
and U8056 (N_8056,N_7540,N_7709);
and U8057 (N_8057,N_7547,N_7546);
or U8058 (N_8058,N_7588,N_7572);
and U8059 (N_8059,N_7736,N_7600);
xnor U8060 (N_8060,N_7758,N_7513);
nand U8061 (N_8061,N_7745,N_7746);
nand U8062 (N_8062,N_7529,N_7609);
nor U8063 (N_8063,N_7570,N_7696);
nor U8064 (N_8064,N_7682,N_7561);
or U8065 (N_8065,N_7632,N_7778);
xnor U8066 (N_8066,N_7507,N_7592);
and U8067 (N_8067,N_7567,N_7726);
nand U8068 (N_8068,N_7543,N_7712);
xnor U8069 (N_8069,N_7556,N_7675);
nand U8070 (N_8070,N_7626,N_7728);
nor U8071 (N_8071,N_7593,N_7621);
and U8072 (N_8072,N_7774,N_7699);
xnor U8073 (N_8073,N_7636,N_7694);
xor U8074 (N_8074,N_7761,N_7580);
nor U8075 (N_8075,N_7726,N_7541);
or U8076 (N_8076,N_7587,N_7595);
nor U8077 (N_8077,N_7755,N_7632);
nand U8078 (N_8078,N_7575,N_7737);
and U8079 (N_8079,N_7526,N_7565);
nor U8080 (N_8080,N_7606,N_7588);
nand U8081 (N_8081,N_7521,N_7764);
nor U8082 (N_8082,N_7744,N_7567);
nand U8083 (N_8083,N_7520,N_7569);
and U8084 (N_8084,N_7681,N_7517);
and U8085 (N_8085,N_7731,N_7560);
and U8086 (N_8086,N_7732,N_7548);
nor U8087 (N_8087,N_7749,N_7792);
nand U8088 (N_8088,N_7794,N_7631);
nand U8089 (N_8089,N_7543,N_7619);
or U8090 (N_8090,N_7746,N_7602);
or U8091 (N_8091,N_7526,N_7600);
and U8092 (N_8092,N_7702,N_7631);
nor U8093 (N_8093,N_7575,N_7630);
and U8094 (N_8094,N_7652,N_7658);
and U8095 (N_8095,N_7559,N_7793);
nand U8096 (N_8096,N_7790,N_7794);
nand U8097 (N_8097,N_7624,N_7642);
nand U8098 (N_8098,N_7721,N_7577);
or U8099 (N_8099,N_7599,N_7737);
or U8100 (N_8100,N_7902,N_7865);
xnor U8101 (N_8101,N_8052,N_8087);
nor U8102 (N_8102,N_7888,N_7962);
and U8103 (N_8103,N_7950,N_8090);
or U8104 (N_8104,N_7956,N_7987);
nor U8105 (N_8105,N_8074,N_7973);
nor U8106 (N_8106,N_7979,N_7804);
or U8107 (N_8107,N_7974,N_8034);
nand U8108 (N_8108,N_7854,N_7822);
nor U8109 (N_8109,N_7935,N_7831);
or U8110 (N_8110,N_7880,N_8007);
nor U8111 (N_8111,N_7845,N_7906);
xor U8112 (N_8112,N_7897,N_8026);
nor U8113 (N_8113,N_8088,N_7910);
xnor U8114 (N_8114,N_7961,N_7801);
or U8115 (N_8115,N_8057,N_7901);
nor U8116 (N_8116,N_8039,N_7819);
and U8117 (N_8117,N_7957,N_7802);
nand U8118 (N_8118,N_7969,N_7967);
nor U8119 (N_8119,N_8059,N_7874);
nand U8120 (N_8120,N_7944,N_8038);
nand U8121 (N_8121,N_8095,N_8075);
or U8122 (N_8122,N_7809,N_7928);
xor U8123 (N_8123,N_7864,N_7986);
nand U8124 (N_8124,N_8033,N_7882);
or U8125 (N_8125,N_7859,N_8093);
or U8126 (N_8126,N_7955,N_8047);
xnor U8127 (N_8127,N_7808,N_7847);
or U8128 (N_8128,N_7826,N_7907);
xnor U8129 (N_8129,N_7964,N_7821);
and U8130 (N_8130,N_7949,N_7998);
or U8131 (N_8131,N_8062,N_7940);
or U8132 (N_8132,N_7927,N_8068);
nand U8133 (N_8133,N_8083,N_7810);
xnor U8134 (N_8134,N_7827,N_7958);
xnor U8135 (N_8135,N_8036,N_7886);
and U8136 (N_8136,N_7913,N_7806);
nand U8137 (N_8137,N_7994,N_7889);
xor U8138 (N_8138,N_8001,N_8050);
or U8139 (N_8139,N_7941,N_7851);
and U8140 (N_8140,N_7938,N_7951);
xor U8141 (N_8141,N_8041,N_7895);
and U8142 (N_8142,N_8015,N_7908);
and U8143 (N_8143,N_7918,N_7936);
nor U8144 (N_8144,N_8053,N_7870);
nor U8145 (N_8145,N_8048,N_7983);
xnor U8146 (N_8146,N_7959,N_8044);
xor U8147 (N_8147,N_7990,N_7834);
and U8148 (N_8148,N_7892,N_7824);
nor U8149 (N_8149,N_8002,N_8076);
xnor U8150 (N_8150,N_7900,N_8079);
and U8151 (N_8151,N_7885,N_7850);
nand U8152 (N_8152,N_8022,N_8085);
or U8153 (N_8153,N_8017,N_7972);
or U8154 (N_8154,N_7853,N_8056);
or U8155 (N_8155,N_7948,N_7988);
and U8156 (N_8156,N_7840,N_7909);
and U8157 (N_8157,N_8054,N_7912);
and U8158 (N_8158,N_7884,N_7861);
or U8159 (N_8159,N_8027,N_7818);
or U8160 (N_8160,N_7820,N_7914);
or U8161 (N_8161,N_8049,N_7849);
nor U8162 (N_8162,N_7862,N_7916);
nor U8163 (N_8163,N_8064,N_7881);
and U8164 (N_8164,N_7937,N_7866);
or U8165 (N_8165,N_8071,N_7970);
xnor U8166 (N_8166,N_7890,N_7878);
or U8167 (N_8167,N_7903,N_8091);
and U8168 (N_8168,N_8003,N_7835);
xnor U8169 (N_8169,N_7975,N_8069);
nor U8170 (N_8170,N_7848,N_7813);
nand U8171 (N_8171,N_7931,N_7904);
xor U8172 (N_8172,N_8005,N_8031);
nor U8173 (N_8173,N_8096,N_8066);
nor U8174 (N_8174,N_7960,N_7981);
and U8175 (N_8175,N_7842,N_7971);
nor U8176 (N_8176,N_7857,N_8018);
nand U8177 (N_8177,N_7980,N_7829);
or U8178 (N_8178,N_8014,N_7920);
nand U8179 (N_8179,N_7896,N_7814);
nand U8180 (N_8180,N_8019,N_7926);
nor U8181 (N_8181,N_7879,N_7965);
nor U8182 (N_8182,N_7929,N_8065);
nand U8183 (N_8183,N_7915,N_7877);
or U8184 (N_8184,N_8067,N_7852);
and U8185 (N_8185,N_7856,N_7828);
xnor U8186 (N_8186,N_7800,N_8084);
nor U8187 (N_8187,N_7841,N_7833);
and U8188 (N_8188,N_7966,N_8098);
and U8189 (N_8189,N_8004,N_8029);
nor U8190 (N_8190,N_8006,N_7844);
or U8191 (N_8191,N_8012,N_8008);
xor U8192 (N_8192,N_8061,N_8063);
nand U8193 (N_8193,N_8035,N_7837);
nor U8194 (N_8194,N_7999,N_8023);
xor U8195 (N_8195,N_7843,N_8046);
nand U8196 (N_8196,N_8097,N_8086);
nor U8197 (N_8197,N_7832,N_7815);
and U8198 (N_8198,N_7934,N_8080);
nand U8199 (N_8199,N_7976,N_7860);
xor U8200 (N_8200,N_7807,N_7947);
nand U8201 (N_8201,N_7977,N_7985);
and U8202 (N_8202,N_8072,N_7989);
nand U8203 (N_8203,N_7875,N_7992);
nor U8204 (N_8204,N_7811,N_7868);
and U8205 (N_8205,N_8016,N_7871);
xnor U8206 (N_8206,N_7963,N_7846);
nand U8207 (N_8207,N_7917,N_7891);
and U8208 (N_8208,N_8092,N_8020);
and U8209 (N_8209,N_8073,N_8078);
or U8210 (N_8210,N_7911,N_7876);
nor U8211 (N_8211,N_8045,N_7919);
and U8212 (N_8212,N_8082,N_7839);
nor U8213 (N_8213,N_7930,N_7996);
and U8214 (N_8214,N_7943,N_8032);
or U8215 (N_8215,N_7869,N_7995);
nand U8216 (N_8216,N_7932,N_7855);
or U8217 (N_8217,N_8040,N_7838);
nand U8218 (N_8218,N_7946,N_7945);
nor U8219 (N_8219,N_7925,N_7921);
nand U8220 (N_8220,N_8013,N_8051);
nand U8221 (N_8221,N_7953,N_7867);
xnor U8222 (N_8222,N_7905,N_8043);
or U8223 (N_8223,N_7823,N_8011);
nor U8224 (N_8224,N_7942,N_7893);
xor U8225 (N_8225,N_7984,N_8010);
nor U8226 (N_8226,N_8081,N_7883);
nor U8227 (N_8227,N_7922,N_7816);
or U8228 (N_8228,N_7872,N_7933);
nor U8229 (N_8229,N_8042,N_7982);
xnor U8230 (N_8230,N_8024,N_8009);
nand U8231 (N_8231,N_8030,N_7812);
xor U8232 (N_8232,N_7997,N_7863);
and U8233 (N_8233,N_8025,N_8028);
and U8234 (N_8234,N_8094,N_7894);
nand U8235 (N_8235,N_8037,N_8021);
or U8236 (N_8236,N_8058,N_7825);
nand U8237 (N_8237,N_7836,N_8055);
nor U8238 (N_8238,N_7968,N_7887);
or U8239 (N_8239,N_7858,N_8000);
nand U8240 (N_8240,N_7924,N_8089);
or U8241 (N_8241,N_8099,N_7991);
and U8242 (N_8242,N_7899,N_8070);
xor U8243 (N_8243,N_7830,N_7873);
or U8244 (N_8244,N_8077,N_7898);
and U8245 (N_8245,N_7952,N_7923);
and U8246 (N_8246,N_8060,N_7939);
nand U8247 (N_8247,N_7803,N_7993);
xor U8248 (N_8248,N_7805,N_7978);
nor U8249 (N_8249,N_7954,N_7817);
xnor U8250 (N_8250,N_8066,N_8076);
xor U8251 (N_8251,N_7823,N_8038);
nor U8252 (N_8252,N_8002,N_8070);
nand U8253 (N_8253,N_8021,N_7810);
or U8254 (N_8254,N_8035,N_7902);
and U8255 (N_8255,N_8060,N_7884);
or U8256 (N_8256,N_7980,N_7992);
nand U8257 (N_8257,N_8002,N_8095);
nor U8258 (N_8258,N_8024,N_7828);
xor U8259 (N_8259,N_8046,N_7822);
or U8260 (N_8260,N_7969,N_7908);
or U8261 (N_8261,N_7867,N_8034);
xnor U8262 (N_8262,N_8046,N_8089);
xnor U8263 (N_8263,N_7958,N_7945);
nand U8264 (N_8264,N_8016,N_8005);
nand U8265 (N_8265,N_8093,N_7989);
or U8266 (N_8266,N_7865,N_7937);
and U8267 (N_8267,N_7951,N_7823);
or U8268 (N_8268,N_7832,N_8053);
nand U8269 (N_8269,N_8059,N_8096);
xnor U8270 (N_8270,N_7819,N_8010);
or U8271 (N_8271,N_7858,N_8096);
and U8272 (N_8272,N_7827,N_7895);
nand U8273 (N_8273,N_8038,N_7814);
nand U8274 (N_8274,N_7986,N_7897);
nor U8275 (N_8275,N_8080,N_7900);
or U8276 (N_8276,N_7813,N_7844);
nor U8277 (N_8277,N_8007,N_7939);
xor U8278 (N_8278,N_7954,N_7903);
and U8279 (N_8279,N_8080,N_8098);
nor U8280 (N_8280,N_7862,N_7948);
nor U8281 (N_8281,N_7803,N_8062);
or U8282 (N_8282,N_8034,N_7976);
and U8283 (N_8283,N_7812,N_7844);
or U8284 (N_8284,N_8044,N_7916);
nand U8285 (N_8285,N_8012,N_7858);
nor U8286 (N_8286,N_7840,N_7836);
nand U8287 (N_8287,N_7900,N_7870);
nor U8288 (N_8288,N_8022,N_7874);
and U8289 (N_8289,N_8030,N_8023);
and U8290 (N_8290,N_8034,N_8068);
nand U8291 (N_8291,N_7884,N_7956);
xor U8292 (N_8292,N_8053,N_7918);
nand U8293 (N_8293,N_7937,N_7859);
and U8294 (N_8294,N_7921,N_7811);
xnor U8295 (N_8295,N_7851,N_7923);
or U8296 (N_8296,N_7958,N_7984);
or U8297 (N_8297,N_8019,N_7917);
or U8298 (N_8298,N_7989,N_7877);
nand U8299 (N_8299,N_7845,N_7929);
nand U8300 (N_8300,N_7840,N_7894);
nor U8301 (N_8301,N_7957,N_7915);
xnor U8302 (N_8302,N_7878,N_7862);
nor U8303 (N_8303,N_7859,N_7834);
nand U8304 (N_8304,N_7979,N_8051);
xnor U8305 (N_8305,N_7826,N_8099);
xnor U8306 (N_8306,N_7894,N_8041);
xor U8307 (N_8307,N_7992,N_8075);
nand U8308 (N_8308,N_7967,N_8099);
xor U8309 (N_8309,N_7962,N_8097);
or U8310 (N_8310,N_7857,N_7881);
xor U8311 (N_8311,N_7859,N_7995);
or U8312 (N_8312,N_7914,N_7969);
and U8313 (N_8313,N_8019,N_8029);
nor U8314 (N_8314,N_7919,N_7812);
and U8315 (N_8315,N_7878,N_8086);
nand U8316 (N_8316,N_8048,N_8038);
and U8317 (N_8317,N_7916,N_8078);
xor U8318 (N_8318,N_8046,N_7990);
nor U8319 (N_8319,N_7924,N_8050);
nor U8320 (N_8320,N_7891,N_7867);
and U8321 (N_8321,N_7898,N_7975);
nand U8322 (N_8322,N_7981,N_7952);
nor U8323 (N_8323,N_8093,N_7999);
or U8324 (N_8324,N_7870,N_7849);
and U8325 (N_8325,N_7951,N_7863);
nand U8326 (N_8326,N_7997,N_7986);
xnor U8327 (N_8327,N_8043,N_7982);
and U8328 (N_8328,N_7926,N_8064);
nand U8329 (N_8329,N_8047,N_7859);
or U8330 (N_8330,N_7892,N_7833);
nand U8331 (N_8331,N_7862,N_7999);
and U8332 (N_8332,N_7963,N_7926);
nand U8333 (N_8333,N_7902,N_7819);
nand U8334 (N_8334,N_7930,N_7839);
nor U8335 (N_8335,N_7886,N_7953);
nand U8336 (N_8336,N_8099,N_8019);
nor U8337 (N_8337,N_7894,N_7899);
nand U8338 (N_8338,N_7848,N_7999);
and U8339 (N_8339,N_7820,N_8043);
and U8340 (N_8340,N_8069,N_7805);
xnor U8341 (N_8341,N_8036,N_7854);
or U8342 (N_8342,N_8045,N_7890);
and U8343 (N_8343,N_8005,N_7919);
xnor U8344 (N_8344,N_7973,N_7891);
xnor U8345 (N_8345,N_8072,N_7880);
and U8346 (N_8346,N_8002,N_7988);
or U8347 (N_8347,N_8004,N_7844);
or U8348 (N_8348,N_8009,N_7905);
xnor U8349 (N_8349,N_7869,N_7887);
nor U8350 (N_8350,N_7934,N_7851);
nor U8351 (N_8351,N_7817,N_7801);
nor U8352 (N_8352,N_7893,N_7876);
xnor U8353 (N_8353,N_8081,N_7981);
nor U8354 (N_8354,N_7863,N_7891);
or U8355 (N_8355,N_8002,N_7936);
xor U8356 (N_8356,N_8011,N_7983);
or U8357 (N_8357,N_7861,N_8089);
nand U8358 (N_8358,N_7920,N_7967);
and U8359 (N_8359,N_7937,N_7888);
xnor U8360 (N_8360,N_7909,N_8013);
nand U8361 (N_8361,N_7943,N_7901);
nor U8362 (N_8362,N_7872,N_7919);
nor U8363 (N_8363,N_7900,N_8040);
or U8364 (N_8364,N_8053,N_7864);
or U8365 (N_8365,N_8005,N_7843);
nand U8366 (N_8366,N_7931,N_7934);
or U8367 (N_8367,N_8065,N_7957);
nor U8368 (N_8368,N_8028,N_7828);
xor U8369 (N_8369,N_7850,N_7905);
nand U8370 (N_8370,N_8083,N_7873);
xnor U8371 (N_8371,N_7908,N_7849);
xor U8372 (N_8372,N_7967,N_7832);
xnor U8373 (N_8373,N_7833,N_7902);
or U8374 (N_8374,N_8041,N_7829);
nand U8375 (N_8375,N_8011,N_7837);
or U8376 (N_8376,N_8044,N_7943);
and U8377 (N_8377,N_7861,N_7915);
xor U8378 (N_8378,N_7990,N_8071);
nand U8379 (N_8379,N_7998,N_8036);
or U8380 (N_8380,N_8039,N_7844);
xnor U8381 (N_8381,N_8013,N_8044);
xor U8382 (N_8382,N_7832,N_7989);
or U8383 (N_8383,N_7829,N_8083);
and U8384 (N_8384,N_7828,N_8051);
nand U8385 (N_8385,N_8048,N_7942);
or U8386 (N_8386,N_8046,N_7913);
xnor U8387 (N_8387,N_8033,N_8036);
and U8388 (N_8388,N_7870,N_7861);
nor U8389 (N_8389,N_7917,N_7869);
nand U8390 (N_8390,N_8059,N_7839);
or U8391 (N_8391,N_7801,N_7998);
nand U8392 (N_8392,N_7837,N_8062);
xnor U8393 (N_8393,N_8028,N_7907);
and U8394 (N_8394,N_7963,N_7865);
nand U8395 (N_8395,N_7962,N_7986);
xnor U8396 (N_8396,N_7890,N_7830);
nor U8397 (N_8397,N_8027,N_8098);
nand U8398 (N_8398,N_7976,N_8095);
xnor U8399 (N_8399,N_8042,N_7861);
and U8400 (N_8400,N_8109,N_8390);
or U8401 (N_8401,N_8260,N_8290);
or U8402 (N_8402,N_8167,N_8226);
nor U8403 (N_8403,N_8168,N_8314);
nand U8404 (N_8404,N_8159,N_8382);
xor U8405 (N_8405,N_8137,N_8172);
nand U8406 (N_8406,N_8101,N_8205);
and U8407 (N_8407,N_8397,N_8294);
nor U8408 (N_8408,N_8125,N_8337);
and U8409 (N_8409,N_8111,N_8350);
nand U8410 (N_8410,N_8333,N_8214);
and U8411 (N_8411,N_8395,N_8152);
nand U8412 (N_8412,N_8153,N_8233);
nand U8413 (N_8413,N_8206,N_8120);
or U8414 (N_8414,N_8182,N_8243);
nor U8415 (N_8415,N_8140,N_8307);
or U8416 (N_8416,N_8339,N_8277);
and U8417 (N_8417,N_8176,N_8129);
and U8418 (N_8418,N_8341,N_8173);
or U8419 (N_8419,N_8132,N_8229);
nor U8420 (N_8420,N_8287,N_8138);
and U8421 (N_8421,N_8385,N_8368);
nand U8422 (N_8422,N_8249,N_8192);
nor U8423 (N_8423,N_8178,N_8275);
xor U8424 (N_8424,N_8263,N_8106);
or U8425 (N_8425,N_8361,N_8216);
xnor U8426 (N_8426,N_8242,N_8388);
and U8427 (N_8427,N_8364,N_8384);
and U8428 (N_8428,N_8255,N_8308);
or U8429 (N_8429,N_8288,N_8117);
and U8430 (N_8430,N_8375,N_8234);
xor U8431 (N_8431,N_8380,N_8261);
nor U8432 (N_8432,N_8210,N_8332);
or U8433 (N_8433,N_8256,N_8164);
nand U8434 (N_8434,N_8200,N_8317);
nand U8435 (N_8435,N_8352,N_8113);
nand U8436 (N_8436,N_8326,N_8188);
nor U8437 (N_8437,N_8363,N_8281);
and U8438 (N_8438,N_8369,N_8244);
nand U8439 (N_8439,N_8126,N_8335);
or U8440 (N_8440,N_8160,N_8128);
xor U8441 (N_8441,N_8238,N_8265);
or U8442 (N_8442,N_8246,N_8280);
nor U8443 (N_8443,N_8141,N_8365);
or U8444 (N_8444,N_8104,N_8377);
or U8445 (N_8445,N_8319,N_8230);
or U8446 (N_8446,N_8186,N_8236);
nand U8447 (N_8447,N_8373,N_8386);
or U8448 (N_8448,N_8348,N_8359);
xor U8449 (N_8449,N_8223,N_8283);
or U8450 (N_8450,N_8391,N_8123);
nor U8451 (N_8451,N_8356,N_8196);
nand U8452 (N_8452,N_8169,N_8122);
xor U8453 (N_8453,N_8181,N_8338);
or U8454 (N_8454,N_8145,N_8313);
and U8455 (N_8455,N_8143,N_8279);
xnor U8456 (N_8456,N_8221,N_8394);
nand U8457 (N_8457,N_8306,N_8144);
and U8458 (N_8458,N_8193,N_8376);
xnor U8459 (N_8459,N_8336,N_8150);
nor U8460 (N_8460,N_8170,N_8184);
nor U8461 (N_8461,N_8222,N_8112);
and U8462 (N_8462,N_8220,N_8180);
and U8463 (N_8463,N_8247,N_8165);
or U8464 (N_8464,N_8166,N_8367);
or U8465 (N_8465,N_8115,N_8268);
nand U8466 (N_8466,N_8118,N_8100);
nand U8467 (N_8467,N_8121,N_8292);
or U8468 (N_8468,N_8107,N_8108);
nor U8469 (N_8469,N_8227,N_8372);
or U8470 (N_8470,N_8362,N_8273);
xor U8471 (N_8471,N_8272,N_8328);
or U8472 (N_8472,N_8371,N_8228);
xnor U8473 (N_8473,N_8217,N_8278);
and U8474 (N_8474,N_8149,N_8312);
nand U8475 (N_8475,N_8235,N_8296);
xor U8476 (N_8476,N_8387,N_8102);
or U8477 (N_8477,N_8199,N_8207);
and U8478 (N_8478,N_8346,N_8389);
and U8479 (N_8479,N_8321,N_8378);
or U8480 (N_8480,N_8293,N_8345);
and U8481 (N_8481,N_8379,N_8171);
or U8482 (N_8482,N_8355,N_8383);
nand U8483 (N_8483,N_8110,N_8330);
or U8484 (N_8484,N_8357,N_8318);
or U8485 (N_8485,N_8301,N_8136);
xor U8486 (N_8486,N_8252,N_8212);
nor U8487 (N_8487,N_8274,N_8237);
nor U8488 (N_8488,N_8157,N_8353);
or U8489 (N_8489,N_8240,N_8399);
or U8490 (N_8490,N_8342,N_8329);
and U8491 (N_8491,N_8340,N_8146);
and U8492 (N_8492,N_8269,N_8135);
or U8493 (N_8493,N_8148,N_8198);
xor U8494 (N_8494,N_8161,N_8158);
or U8495 (N_8495,N_8185,N_8191);
nand U8496 (N_8496,N_8322,N_8224);
nand U8497 (N_8497,N_8177,N_8289);
xnor U8498 (N_8498,N_8209,N_8351);
and U8499 (N_8499,N_8291,N_8300);
nand U8500 (N_8500,N_8162,N_8259);
nor U8501 (N_8501,N_8195,N_8190);
xor U8502 (N_8502,N_8334,N_8213);
or U8503 (N_8503,N_8187,N_8253);
nor U8504 (N_8504,N_8324,N_8124);
nor U8505 (N_8505,N_8215,N_8267);
and U8506 (N_8506,N_8134,N_8323);
nor U8507 (N_8507,N_8358,N_8305);
and U8508 (N_8508,N_8262,N_8114);
or U8509 (N_8509,N_8127,N_8211);
nand U8510 (N_8510,N_8154,N_8298);
xnor U8511 (N_8511,N_8201,N_8103);
nor U8512 (N_8512,N_8151,N_8285);
xor U8513 (N_8513,N_8282,N_8366);
xor U8514 (N_8514,N_8232,N_8208);
or U8515 (N_8515,N_8270,N_8320);
or U8516 (N_8516,N_8284,N_8231);
or U8517 (N_8517,N_8303,N_8315);
xor U8518 (N_8518,N_8225,N_8174);
nand U8519 (N_8519,N_8139,N_8248);
nand U8520 (N_8520,N_8189,N_8271);
xnor U8521 (N_8521,N_8254,N_8374);
xor U8522 (N_8522,N_8203,N_8116);
nor U8523 (N_8523,N_8343,N_8142);
xnor U8524 (N_8524,N_8360,N_8302);
nand U8525 (N_8525,N_8295,N_8381);
xnor U8526 (N_8526,N_8310,N_8264);
xor U8527 (N_8527,N_8325,N_8204);
or U8528 (N_8528,N_8202,N_8392);
or U8529 (N_8529,N_8297,N_8250);
xnor U8530 (N_8530,N_8276,N_8393);
nand U8531 (N_8531,N_8131,N_8398);
and U8532 (N_8532,N_8239,N_8331);
or U8533 (N_8533,N_8299,N_8197);
xor U8534 (N_8534,N_8344,N_8257);
xnor U8535 (N_8535,N_8219,N_8251);
or U8536 (N_8536,N_8218,N_8179);
nand U8537 (N_8537,N_8175,N_8396);
xnor U8538 (N_8538,N_8258,N_8309);
xor U8539 (N_8539,N_8311,N_8316);
and U8540 (N_8540,N_8130,N_8347);
or U8541 (N_8541,N_8156,N_8147);
xor U8542 (N_8542,N_8349,N_8327);
or U8543 (N_8543,N_8370,N_8163);
xor U8544 (N_8544,N_8133,N_8105);
nor U8545 (N_8545,N_8266,N_8119);
or U8546 (N_8546,N_8354,N_8286);
xor U8547 (N_8547,N_8194,N_8183);
nor U8548 (N_8548,N_8245,N_8241);
or U8549 (N_8549,N_8304,N_8155);
nand U8550 (N_8550,N_8295,N_8115);
or U8551 (N_8551,N_8344,N_8134);
nor U8552 (N_8552,N_8324,N_8168);
or U8553 (N_8553,N_8328,N_8384);
nor U8554 (N_8554,N_8255,N_8209);
xnor U8555 (N_8555,N_8223,N_8134);
and U8556 (N_8556,N_8159,N_8265);
and U8557 (N_8557,N_8331,N_8235);
nand U8558 (N_8558,N_8183,N_8350);
and U8559 (N_8559,N_8136,N_8232);
nand U8560 (N_8560,N_8378,N_8302);
or U8561 (N_8561,N_8316,N_8231);
or U8562 (N_8562,N_8399,N_8377);
xor U8563 (N_8563,N_8150,N_8378);
and U8564 (N_8564,N_8288,N_8373);
and U8565 (N_8565,N_8291,N_8133);
or U8566 (N_8566,N_8373,N_8124);
and U8567 (N_8567,N_8108,N_8321);
nor U8568 (N_8568,N_8134,N_8118);
nor U8569 (N_8569,N_8317,N_8165);
and U8570 (N_8570,N_8328,N_8144);
and U8571 (N_8571,N_8181,N_8337);
nor U8572 (N_8572,N_8334,N_8196);
xnor U8573 (N_8573,N_8172,N_8365);
xor U8574 (N_8574,N_8106,N_8274);
and U8575 (N_8575,N_8165,N_8379);
nor U8576 (N_8576,N_8372,N_8389);
or U8577 (N_8577,N_8388,N_8268);
nor U8578 (N_8578,N_8326,N_8155);
nand U8579 (N_8579,N_8324,N_8392);
nor U8580 (N_8580,N_8171,N_8128);
or U8581 (N_8581,N_8201,N_8301);
and U8582 (N_8582,N_8144,N_8275);
nand U8583 (N_8583,N_8215,N_8101);
nor U8584 (N_8584,N_8168,N_8376);
and U8585 (N_8585,N_8298,N_8162);
nor U8586 (N_8586,N_8363,N_8330);
and U8587 (N_8587,N_8385,N_8328);
and U8588 (N_8588,N_8383,N_8331);
xor U8589 (N_8589,N_8278,N_8253);
xor U8590 (N_8590,N_8268,N_8396);
and U8591 (N_8591,N_8134,N_8324);
and U8592 (N_8592,N_8310,N_8290);
or U8593 (N_8593,N_8136,N_8255);
xor U8594 (N_8594,N_8312,N_8163);
xor U8595 (N_8595,N_8261,N_8180);
or U8596 (N_8596,N_8225,N_8210);
and U8597 (N_8597,N_8170,N_8351);
nand U8598 (N_8598,N_8325,N_8114);
xor U8599 (N_8599,N_8294,N_8346);
nand U8600 (N_8600,N_8338,N_8263);
or U8601 (N_8601,N_8275,N_8349);
xor U8602 (N_8602,N_8193,N_8167);
nor U8603 (N_8603,N_8368,N_8356);
and U8604 (N_8604,N_8323,N_8361);
or U8605 (N_8605,N_8234,N_8393);
nor U8606 (N_8606,N_8189,N_8344);
xor U8607 (N_8607,N_8374,N_8107);
and U8608 (N_8608,N_8394,N_8105);
nor U8609 (N_8609,N_8275,N_8227);
or U8610 (N_8610,N_8104,N_8385);
nand U8611 (N_8611,N_8291,N_8383);
xor U8612 (N_8612,N_8386,N_8228);
xnor U8613 (N_8613,N_8383,N_8382);
nor U8614 (N_8614,N_8130,N_8248);
and U8615 (N_8615,N_8326,N_8385);
xnor U8616 (N_8616,N_8258,N_8345);
or U8617 (N_8617,N_8149,N_8246);
and U8618 (N_8618,N_8205,N_8358);
or U8619 (N_8619,N_8307,N_8304);
xor U8620 (N_8620,N_8330,N_8345);
or U8621 (N_8621,N_8196,N_8250);
and U8622 (N_8622,N_8349,N_8175);
xor U8623 (N_8623,N_8258,N_8370);
nand U8624 (N_8624,N_8292,N_8373);
nor U8625 (N_8625,N_8389,N_8345);
xor U8626 (N_8626,N_8118,N_8322);
or U8627 (N_8627,N_8298,N_8178);
nor U8628 (N_8628,N_8122,N_8173);
nand U8629 (N_8629,N_8345,N_8254);
xor U8630 (N_8630,N_8257,N_8353);
and U8631 (N_8631,N_8325,N_8115);
nand U8632 (N_8632,N_8104,N_8264);
or U8633 (N_8633,N_8377,N_8225);
or U8634 (N_8634,N_8385,N_8313);
or U8635 (N_8635,N_8286,N_8393);
nand U8636 (N_8636,N_8305,N_8315);
nor U8637 (N_8637,N_8347,N_8300);
or U8638 (N_8638,N_8162,N_8397);
and U8639 (N_8639,N_8299,N_8376);
or U8640 (N_8640,N_8351,N_8105);
nand U8641 (N_8641,N_8135,N_8232);
and U8642 (N_8642,N_8152,N_8102);
xnor U8643 (N_8643,N_8178,N_8348);
or U8644 (N_8644,N_8187,N_8121);
and U8645 (N_8645,N_8177,N_8336);
or U8646 (N_8646,N_8163,N_8300);
nor U8647 (N_8647,N_8246,N_8302);
nor U8648 (N_8648,N_8329,N_8224);
nand U8649 (N_8649,N_8211,N_8145);
nor U8650 (N_8650,N_8263,N_8108);
or U8651 (N_8651,N_8214,N_8373);
or U8652 (N_8652,N_8368,N_8312);
and U8653 (N_8653,N_8235,N_8233);
or U8654 (N_8654,N_8194,N_8293);
or U8655 (N_8655,N_8384,N_8276);
nor U8656 (N_8656,N_8179,N_8375);
nand U8657 (N_8657,N_8242,N_8321);
and U8658 (N_8658,N_8205,N_8220);
nor U8659 (N_8659,N_8160,N_8107);
or U8660 (N_8660,N_8167,N_8300);
or U8661 (N_8661,N_8370,N_8213);
or U8662 (N_8662,N_8296,N_8126);
and U8663 (N_8663,N_8204,N_8225);
nor U8664 (N_8664,N_8101,N_8106);
nor U8665 (N_8665,N_8335,N_8357);
nor U8666 (N_8666,N_8236,N_8196);
nor U8667 (N_8667,N_8198,N_8381);
nand U8668 (N_8668,N_8329,N_8292);
nor U8669 (N_8669,N_8251,N_8143);
nand U8670 (N_8670,N_8344,N_8183);
nand U8671 (N_8671,N_8296,N_8177);
or U8672 (N_8672,N_8397,N_8105);
nand U8673 (N_8673,N_8376,N_8271);
or U8674 (N_8674,N_8331,N_8318);
nand U8675 (N_8675,N_8175,N_8354);
xor U8676 (N_8676,N_8379,N_8182);
nor U8677 (N_8677,N_8248,N_8260);
or U8678 (N_8678,N_8188,N_8195);
and U8679 (N_8679,N_8373,N_8259);
or U8680 (N_8680,N_8240,N_8182);
nor U8681 (N_8681,N_8252,N_8176);
nand U8682 (N_8682,N_8306,N_8211);
or U8683 (N_8683,N_8331,N_8283);
xor U8684 (N_8684,N_8376,N_8243);
nand U8685 (N_8685,N_8272,N_8264);
nand U8686 (N_8686,N_8345,N_8108);
nor U8687 (N_8687,N_8384,N_8153);
nand U8688 (N_8688,N_8243,N_8103);
xnor U8689 (N_8689,N_8333,N_8210);
xnor U8690 (N_8690,N_8340,N_8289);
nor U8691 (N_8691,N_8334,N_8356);
nor U8692 (N_8692,N_8135,N_8393);
xnor U8693 (N_8693,N_8380,N_8202);
or U8694 (N_8694,N_8107,N_8147);
nor U8695 (N_8695,N_8202,N_8165);
nand U8696 (N_8696,N_8203,N_8244);
or U8697 (N_8697,N_8354,N_8315);
or U8698 (N_8698,N_8347,N_8117);
nor U8699 (N_8699,N_8148,N_8337);
and U8700 (N_8700,N_8670,N_8572);
nand U8701 (N_8701,N_8659,N_8426);
nand U8702 (N_8702,N_8688,N_8591);
xor U8703 (N_8703,N_8541,N_8442);
or U8704 (N_8704,N_8446,N_8519);
nor U8705 (N_8705,N_8536,N_8565);
nand U8706 (N_8706,N_8436,N_8498);
nor U8707 (N_8707,N_8407,N_8470);
nor U8708 (N_8708,N_8653,N_8515);
xnor U8709 (N_8709,N_8404,N_8612);
and U8710 (N_8710,N_8545,N_8444);
nand U8711 (N_8711,N_8566,N_8550);
xnor U8712 (N_8712,N_8613,N_8418);
nor U8713 (N_8713,N_8409,N_8481);
or U8714 (N_8714,N_8627,N_8656);
or U8715 (N_8715,N_8524,N_8680);
nand U8716 (N_8716,N_8563,N_8577);
nor U8717 (N_8717,N_8676,N_8672);
nand U8718 (N_8718,N_8514,N_8505);
nand U8719 (N_8719,N_8522,N_8467);
or U8720 (N_8720,N_8585,N_8685);
xnor U8721 (N_8721,N_8594,N_8606);
and U8722 (N_8722,N_8438,N_8678);
xor U8723 (N_8723,N_8521,N_8421);
nor U8724 (N_8724,N_8491,N_8664);
or U8725 (N_8725,N_8490,N_8555);
xnor U8726 (N_8726,N_8400,N_8580);
or U8727 (N_8727,N_8598,N_8658);
nand U8728 (N_8728,N_8668,N_8624);
nor U8729 (N_8729,N_8619,N_8560);
nor U8730 (N_8730,N_8649,N_8452);
or U8731 (N_8731,N_8574,N_8494);
nand U8732 (N_8732,N_8487,N_8636);
or U8733 (N_8733,N_8584,N_8626);
or U8734 (N_8734,N_8643,N_8699);
xnor U8735 (N_8735,N_8543,N_8607);
or U8736 (N_8736,N_8513,N_8506);
or U8737 (N_8737,N_8639,N_8599);
xnor U8738 (N_8738,N_8504,N_8661);
and U8739 (N_8739,N_8679,N_8611);
and U8740 (N_8740,N_8581,N_8546);
and U8741 (N_8741,N_8439,N_8556);
nand U8742 (N_8742,N_8466,N_8674);
nor U8743 (N_8743,N_8665,N_8440);
and U8744 (N_8744,N_8651,N_8547);
nor U8745 (N_8745,N_8632,N_8488);
nand U8746 (N_8746,N_8542,N_8419);
and U8747 (N_8747,N_8596,N_8635);
and U8748 (N_8748,N_8427,N_8424);
nor U8749 (N_8749,N_8423,N_8475);
nor U8750 (N_8750,N_8468,N_8507);
nor U8751 (N_8751,N_8537,N_8479);
nand U8752 (N_8752,N_8601,N_8402);
nor U8753 (N_8753,N_8549,N_8562);
and U8754 (N_8754,N_8569,N_8633);
nor U8755 (N_8755,N_8590,N_8573);
xnor U8756 (N_8756,N_8425,N_8640);
or U8757 (N_8757,N_8692,N_8631);
nand U8758 (N_8758,N_8533,N_8638);
and U8759 (N_8759,N_8625,N_8422);
xor U8760 (N_8760,N_8518,N_8460);
and U8761 (N_8761,N_8647,N_8579);
and U8762 (N_8762,N_8583,N_8551);
nor U8763 (N_8763,N_8482,N_8684);
nor U8764 (N_8764,N_8673,N_8526);
or U8765 (N_8765,N_8682,N_8403);
nand U8766 (N_8766,N_8464,N_8642);
nand U8767 (N_8767,N_8617,N_8530);
or U8768 (N_8768,N_8695,N_8570);
nor U8769 (N_8769,N_8408,N_8630);
or U8770 (N_8770,N_8534,N_8629);
nor U8771 (N_8771,N_8677,N_8662);
or U8772 (N_8772,N_8645,N_8655);
or U8773 (N_8773,N_8535,N_8401);
xnor U8774 (N_8774,N_8480,N_8447);
or U8775 (N_8775,N_8463,N_8628);
and U8776 (N_8776,N_8508,N_8478);
nor U8777 (N_8777,N_8552,N_8553);
nor U8778 (N_8778,N_8589,N_8689);
nor U8779 (N_8779,N_8693,N_8511);
nor U8780 (N_8780,N_8623,N_8435);
nand U8781 (N_8781,N_8483,N_8527);
or U8782 (N_8782,N_8548,N_8492);
and U8783 (N_8783,N_8586,N_8528);
nor U8784 (N_8784,N_8441,N_8465);
or U8785 (N_8785,N_8644,N_8554);
nand U8786 (N_8786,N_8669,N_8477);
xnor U8787 (N_8787,N_8559,N_8600);
or U8788 (N_8788,N_8576,N_8690);
or U8789 (N_8789,N_8461,N_8431);
or U8790 (N_8790,N_8503,N_8578);
nand U8791 (N_8791,N_8621,N_8592);
nand U8792 (N_8792,N_8540,N_8671);
or U8793 (N_8793,N_8501,N_8429);
nor U8794 (N_8794,N_8648,N_8420);
xor U8795 (N_8795,N_8597,N_8634);
xnor U8796 (N_8796,N_8660,N_8687);
nor U8797 (N_8797,N_8694,N_8489);
nor U8798 (N_8798,N_8496,N_8509);
nor U8799 (N_8799,N_8525,N_8430);
and U8800 (N_8800,N_8493,N_8502);
nand U8801 (N_8801,N_8675,N_8428);
or U8802 (N_8802,N_8575,N_8610);
nor U8803 (N_8803,N_8416,N_8450);
nor U8804 (N_8804,N_8512,N_8456);
nor U8805 (N_8805,N_8538,N_8457);
nand U8806 (N_8806,N_8414,N_8568);
or U8807 (N_8807,N_8471,N_8432);
nand U8808 (N_8808,N_8500,N_8458);
xnor U8809 (N_8809,N_8567,N_8455);
xor U8810 (N_8810,N_8698,N_8615);
nand U8811 (N_8811,N_8417,N_8469);
nand U8812 (N_8812,N_8410,N_8454);
and U8813 (N_8813,N_8415,N_8602);
xor U8814 (N_8814,N_8531,N_8614);
and U8815 (N_8815,N_8652,N_8462);
nor U8816 (N_8816,N_8474,N_8654);
nand U8817 (N_8817,N_8641,N_8472);
and U8818 (N_8818,N_8520,N_8434);
and U8819 (N_8819,N_8604,N_8532);
or U8820 (N_8820,N_8587,N_8405);
nand U8821 (N_8821,N_8433,N_8588);
nand U8822 (N_8822,N_8564,N_8561);
nor U8823 (N_8823,N_8681,N_8620);
and U8824 (N_8824,N_8448,N_8646);
and U8825 (N_8825,N_8486,N_8618);
nand U8826 (N_8826,N_8616,N_8406);
or U8827 (N_8827,N_8557,N_8609);
nor U8828 (N_8828,N_8451,N_8691);
or U8829 (N_8829,N_8571,N_8484);
or U8830 (N_8830,N_8411,N_8622);
nor U8831 (N_8831,N_8495,N_8697);
nand U8832 (N_8832,N_8453,N_8485);
nor U8833 (N_8833,N_8412,N_8666);
and U8834 (N_8834,N_8593,N_8459);
xnor U8835 (N_8835,N_8413,N_8582);
or U8836 (N_8836,N_8529,N_8663);
xnor U8837 (N_8837,N_8449,N_8473);
xor U8838 (N_8838,N_8683,N_8443);
nand U8839 (N_8839,N_8523,N_8539);
nor U8840 (N_8840,N_8497,N_8686);
nor U8841 (N_8841,N_8696,N_8595);
and U8842 (N_8842,N_8516,N_8657);
nand U8843 (N_8843,N_8608,N_8637);
and U8844 (N_8844,N_8437,N_8650);
nor U8845 (N_8845,N_8517,N_8667);
nand U8846 (N_8846,N_8499,N_8445);
and U8847 (N_8847,N_8510,N_8544);
nor U8848 (N_8848,N_8558,N_8603);
or U8849 (N_8849,N_8476,N_8605);
and U8850 (N_8850,N_8577,N_8628);
nand U8851 (N_8851,N_8455,N_8685);
nand U8852 (N_8852,N_8684,N_8678);
or U8853 (N_8853,N_8699,N_8492);
nor U8854 (N_8854,N_8524,N_8631);
and U8855 (N_8855,N_8542,N_8511);
xnor U8856 (N_8856,N_8537,N_8643);
nor U8857 (N_8857,N_8696,N_8581);
nand U8858 (N_8858,N_8483,N_8691);
or U8859 (N_8859,N_8426,N_8546);
or U8860 (N_8860,N_8420,N_8484);
and U8861 (N_8861,N_8614,N_8508);
or U8862 (N_8862,N_8447,N_8432);
nand U8863 (N_8863,N_8585,N_8559);
and U8864 (N_8864,N_8671,N_8417);
and U8865 (N_8865,N_8495,N_8525);
and U8866 (N_8866,N_8677,N_8605);
nand U8867 (N_8867,N_8511,N_8449);
nor U8868 (N_8868,N_8499,N_8634);
and U8869 (N_8869,N_8588,N_8473);
or U8870 (N_8870,N_8448,N_8638);
nor U8871 (N_8871,N_8524,N_8421);
xor U8872 (N_8872,N_8584,N_8460);
xor U8873 (N_8873,N_8438,N_8669);
and U8874 (N_8874,N_8660,N_8488);
nor U8875 (N_8875,N_8579,N_8515);
xor U8876 (N_8876,N_8407,N_8537);
nor U8877 (N_8877,N_8633,N_8582);
nand U8878 (N_8878,N_8439,N_8577);
nand U8879 (N_8879,N_8409,N_8642);
nand U8880 (N_8880,N_8689,N_8557);
nor U8881 (N_8881,N_8616,N_8565);
nor U8882 (N_8882,N_8416,N_8657);
xnor U8883 (N_8883,N_8439,N_8530);
nand U8884 (N_8884,N_8691,N_8552);
nand U8885 (N_8885,N_8620,N_8605);
xnor U8886 (N_8886,N_8660,N_8467);
and U8887 (N_8887,N_8647,N_8493);
xnor U8888 (N_8888,N_8409,N_8521);
or U8889 (N_8889,N_8588,N_8687);
xor U8890 (N_8890,N_8559,N_8501);
nor U8891 (N_8891,N_8566,N_8459);
nor U8892 (N_8892,N_8533,N_8618);
xnor U8893 (N_8893,N_8440,N_8659);
nand U8894 (N_8894,N_8593,N_8445);
xnor U8895 (N_8895,N_8481,N_8521);
nand U8896 (N_8896,N_8513,N_8577);
nor U8897 (N_8897,N_8651,N_8633);
and U8898 (N_8898,N_8525,N_8491);
xnor U8899 (N_8899,N_8678,N_8457);
nor U8900 (N_8900,N_8561,N_8633);
xor U8901 (N_8901,N_8461,N_8487);
nor U8902 (N_8902,N_8421,N_8519);
nor U8903 (N_8903,N_8499,N_8595);
and U8904 (N_8904,N_8435,N_8407);
and U8905 (N_8905,N_8443,N_8437);
or U8906 (N_8906,N_8418,N_8490);
xor U8907 (N_8907,N_8403,N_8451);
nand U8908 (N_8908,N_8628,N_8642);
xor U8909 (N_8909,N_8429,N_8407);
and U8910 (N_8910,N_8604,N_8673);
nand U8911 (N_8911,N_8646,N_8494);
nand U8912 (N_8912,N_8699,N_8679);
and U8913 (N_8913,N_8614,N_8611);
nor U8914 (N_8914,N_8473,N_8522);
or U8915 (N_8915,N_8448,N_8556);
or U8916 (N_8916,N_8404,N_8544);
nor U8917 (N_8917,N_8596,N_8618);
xor U8918 (N_8918,N_8489,N_8486);
and U8919 (N_8919,N_8647,N_8509);
or U8920 (N_8920,N_8619,N_8427);
nand U8921 (N_8921,N_8522,N_8459);
nand U8922 (N_8922,N_8421,N_8601);
nand U8923 (N_8923,N_8446,N_8666);
nor U8924 (N_8924,N_8634,N_8515);
and U8925 (N_8925,N_8689,N_8403);
xnor U8926 (N_8926,N_8585,N_8675);
nand U8927 (N_8927,N_8410,N_8639);
and U8928 (N_8928,N_8519,N_8506);
and U8929 (N_8929,N_8412,N_8452);
xor U8930 (N_8930,N_8590,N_8432);
nand U8931 (N_8931,N_8646,N_8640);
xnor U8932 (N_8932,N_8403,N_8438);
nor U8933 (N_8933,N_8669,N_8439);
xnor U8934 (N_8934,N_8469,N_8632);
or U8935 (N_8935,N_8418,N_8485);
or U8936 (N_8936,N_8613,N_8506);
or U8937 (N_8937,N_8656,N_8454);
or U8938 (N_8938,N_8640,N_8442);
nand U8939 (N_8939,N_8622,N_8432);
or U8940 (N_8940,N_8545,N_8608);
and U8941 (N_8941,N_8685,N_8603);
nand U8942 (N_8942,N_8528,N_8645);
or U8943 (N_8943,N_8476,N_8606);
xor U8944 (N_8944,N_8483,N_8531);
nand U8945 (N_8945,N_8627,N_8536);
or U8946 (N_8946,N_8490,N_8445);
and U8947 (N_8947,N_8514,N_8470);
and U8948 (N_8948,N_8405,N_8459);
or U8949 (N_8949,N_8488,N_8667);
nand U8950 (N_8950,N_8423,N_8416);
or U8951 (N_8951,N_8602,N_8635);
nor U8952 (N_8952,N_8427,N_8431);
xor U8953 (N_8953,N_8486,N_8653);
or U8954 (N_8954,N_8635,N_8617);
and U8955 (N_8955,N_8427,N_8539);
or U8956 (N_8956,N_8570,N_8606);
nor U8957 (N_8957,N_8428,N_8493);
and U8958 (N_8958,N_8642,N_8543);
nand U8959 (N_8959,N_8495,N_8458);
nand U8960 (N_8960,N_8467,N_8509);
nor U8961 (N_8961,N_8533,N_8518);
xor U8962 (N_8962,N_8531,N_8598);
nor U8963 (N_8963,N_8429,N_8534);
nand U8964 (N_8964,N_8608,N_8495);
or U8965 (N_8965,N_8544,N_8432);
xnor U8966 (N_8966,N_8577,N_8639);
nand U8967 (N_8967,N_8547,N_8536);
or U8968 (N_8968,N_8565,N_8462);
or U8969 (N_8969,N_8457,N_8593);
nand U8970 (N_8970,N_8492,N_8634);
or U8971 (N_8971,N_8559,N_8572);
nand U8972 (N_8972,N_8505,N_8510);
nor U8973 (N_8973,N_8663,N_8435);
nor U8974 (N_8974,N_8634,N_8672);
or U8975 (N_8975,N_8598,N_8585);
nand U8976 (N_8976,N_8427,N_8699);
or U8977 (N_8977,N_8462,N_8426);
nand U8978 (N_8978,N_8582,N_8553);
or U8979 (N_8979,N_8598,N_8553);
and U8980 (N_8980,N_8558,N_8683);
nor U8981 (N_8981,N_8438,N_8456);
or U8982 (N_8982,N_8549,N_8553);
nor U8983 (N_8983,N_8666,N_8567);
nand U8984 (N_8984,N_8495,N_8448);
nand U8985 (N_8985,N_8454,N_8695);
xnor U8986 (N_8986,N_8619,N_8544);
xnor U8987 (N_8987,N_8682,N_8529);
or U8988 (N_8988,N_8600,N_8529);
nand U8989 (N_8989,N_8405,N_8462);
nand U8990 (N_8990,N_8615,N_8484);
nor U8991 (N_8991,N_8413,N_8666);
and U8992 (N_8992,N_8609,N_8528);
xor U8993 (N_8993,N_8459,N_8519);
nor U8994 (N_8994,N_8628,N_8435);
xor U8995 (N_8995,N_8490,N_8402);
or U8996 (N_8996,N_8697,N_8453);
nor U8997 (N_8997,N_8450,N_8609);
nor U8998 (N_8998,N_8564,N_8524);
xor U8999 (N_8999,N_8480,N_8635);
xor U9000 (N_9000,N_8848,N_8718);
or U9001 (N_9001,N_8846,N_8915);
nand U9002 (N_9002,N_8958,N_8828);
nand U9003 (N_9003,N_8923,N_8991);
nor U9004 (N_9004,N_8759,N_8939);
nor U9005 (N_9005,N_8932,N_8983);
nand U9006 (N_9006,N_8928,N_8804);
nor U9007 (N_9007,N_8784,N_8965);
nor U9008 (N_9008,N_8900,N_8836);
nor U9009 (N_9009,N_8895,N_8978);
or U9010 (N_9010,N_8856,N_8730);
or U9011 (N_9011,N_8777,N_8801);
xor U9012 (N_9012,N_8998,N_8829);
xor U9013 (N_9013,N_8768,N_8946);
nand U9014 (N_9014,N_8857,N_8742);
xnor U9015 (N_9015,N_8729,N_8847);
nand U9016 (N_9016,N_8894,N_8785);
or U9017 (N_9017,N_8853,N_8766);
or U9018 (N_9018,N_8772,N_8883);
xor U9019 (N_9019,N_8957,N_8840);
and U9020 (N_9020,N_8859,N_8897);
nand U9021 (N_9021,N_8796,N_8728);
or U9022 (N_9022,N_8988,N_8929);
or U9023 (N_9023,N_8714,N_8892);
and U9024 (N_9024,N_8980,N_8758);
and U9025 (N_9025,N_8783,N_8954);
xor U9026 (N_9026,N_8996,N_8935);
xor U9027 (N_9027,N_8750,N_8845);
or U9028 (N_9028,N_8986,N_8921);
and U9029 (N_9029,N_8789,N_8955);
nor U9030 (N_9030,N_8969,N_8820);
xnor U9031 (N_9031,N_8731,N_8990);
or U9032 (N_9032,N_8706,N_8740);
xor U9033 (N_9033,N_8934,N_8858);
or U9034 (N_9034,N_8912,N_8925);
nand U9035 (N_9035,N_8924,N_8821);
xor U9036 (N_9036,N_8888,N_8945);
xor U9037 (N_9037,N_8933,N_8745);
and U9038 (N_9038,N_8974,N_8787);
nand U9039 (N_9039,N_8709,N_8802);
and U9040 (N_9040,N_8819,N_8916);
nand U9041 (N_9041,N_8850,N_8962);
or U9042 (N_9042,N_8989,N_8979);
xor U9043 (N_9043,N_8719,N_8757);
xor U9044 (N_9044,N_8815,N_8755);
nor U9045 (N_9045,N_8947,N_8893);
nor U9046 (N_9046,N_8908,N_8737);
or U9047 (N_9047,N_8807,N_8941);
and U9048 (N_9048,N_8876,N_8736);
nand U9049 (N_9049,N_8762,N_8701);
nand U9050 (N_9050,N_8826,N_8767);
nand U9051 (N_9051,N_8964,N_8746);
or U9052 (N_9052,N_8782,N_8860);
and U9053 (N_9053,N_8995,N_8707);
nor U9054 (N_9054,N_8960,N_8884);
nand U9055 (N_9055,N_8806,N_8812);
nor U9056 (N_9056,N_8744,N_8702);
or U9057 (N_9057,N_8752,N_8887);
nand U9058 (N_9058,N_8833,N_8712);
and U9059 (N_9059,N_8715,N_8727);
and U9060 (N_9060,N_8854,N_8753);
or U9061 (N_9061,N_8798,N_8704);
nand U9062 (N_9062,N_8993,N_8976);
and U9063 (N_9063,N_8961,N_8985);
xor U9064 (N_9064,N_8809,N_8973);
nor U9065 (N_9065,N_8867,N_8920);
or U9066 (N_9066,N_8899,N_8811);
and U9067 (N_9067,N_8902,N_8825);
nor U9068 (N_9068,N_8837,N_8891);
or U9069 (N_9069,N_8841,N_8723);
nor U9070 (N_9070,N_8926,N_8832);
xor U9071 (N_9071,N_8901,N_8756);
xor U9072 (N_9072,N_8968,N_8786);
nor U9073 (N_9073,N_8918,N_8844);
nor U9074 (N_9074,N_8999,N_8710);
and U9075 (N_9075,N_8963,N_8880);
nand U9076 (N_9076,N_8975,N_8748);
or U9077 (N_9077,N_8722,N_8910);
and U9078 (N_9078,N_8919,N_8773);
and U9079 (N_9079,N_8713,N_8834);
nand U9080 (N_9080,N_8776,N_8953);
xor U9081 (N_9081,N_8703,N_8913);
and U9082 (N_9082,N_8869,N_8816);
or U9083 (N_9083,N_8780,N_8863);
nand U9084 (N_9084,N_8808,N_8747);
nand U9085 (N_9085,N_8940,N_8865);
or U9086 (N_9086,N_8831,N_8779);
and U9087 (N_9087,N_8938,N_8874);
nand U9088 (N_9088,N_8734,N_8970);
or U9089 (N_9089,N_8862,N_8971);
and U9090 (N_9090,N_8765,N_8977);
xnor U9091 (N_9091,N_8788,N_8878);
or U9092 (N_9092,N_8984,N_8814);
nand U9093 (N_9093,N_8823,N_8864);
nor U9094 (N_9094,N_8800,N_8726);
nor U9095 (N_9095,N_8851,N_8872);
nor U9096 (N_9096,N_8793,N_8795);
or U9097 (N_9097,N_8944,N_8917);
nor U9098 (N_9098,N_8700,N_8922);
nor U9099 (N_9099,N_8914,N_8931);
nor U9100 (N_9100,N_8763,N_8794);
nor U9101 (N_9101,N_8861,N_8855);
or U9102 (N_9102,N_8966,N_8790);
nor U9103 (N_9103,N_8879,N_8906);
nor U9104 (N_9104,N_8911,N_8875);
xor U9105 (N_9105,N_8799,N_8838);
and U9106 (N_9106,N_8760,N_8972);
or U9107 (N_9107,N_8904,N_8959);
xnor U9108 (N_9108,N_8724,N_8882);
xnor U9109 (N_9109,N_8890,N_8805);
or U9110 (N_9110,N_8774,N_8754);
or U9111 (N_9111,N_8791,N_8871);
xor U9112 (N_9112,N_8739,N_8949);
and U9113 (N_9113,N_8956,N_8927);
or U9114 (N_9114,N_8810,N_8716);
or U9115 (N_9115,N_8951,N_8903);
nand U9116 (N_9116,N_8943,N_8997);
nand U9117 (N_9117,N_8705,N_8721);
nand U9118 (N_9118,N_8849,N_8813);
and U9119 (N_9119,N_8907,N_8898);
nor U9120 (N_9120,N_8896,N_8905);
nand U9121 (N_9121,N_8771,N_8937);
xor U9122 (N_9122,N_8797,N_8761);
or U9123 (N_9123,N_8769,N_8885);
nor U9124 (N_9124,N_8881,N_8822);
or U9125 (N_9125,N_8792,N_8948);
nor U9126 (N_9126,N_8952,N_8738);
or U9127 (N_9127,N_8743,N_8725);
or U9128 (N_9128,N_8839,N_8817);
or U9129 (N_9129,N_8830,N_8868);
nor U9130 (N_9130,N_8775,N_8852);
nand U9131 (N_9131,N_8982,N_8781);
and U9132 (N_9132,N_8987,N_8877);
nor U9133 (N_9133,N_8873,N_8866);
nand U9134 (N_9134,N_8992,N_8741);
nor U9135 (N_9135,N_8870,N_8824);
or U9136 (N_9136,N_8733,N_8717);
and U9137 (N_9137,N_8735,N_8749);
and U9138 (N_9138,N_8843,N_8751);
nor U9139 (N_9139,N_8720,N_8994);
nand U9140 (N_9140,N_8770,N_8842);
and U9141 (N_9141,N_8942,N_8967);
xnor U9142 (N_9142,N_8889,N_8708);
or U9143 (N_9143,N_8886,N_8818);
nand U9144 (N_9144,N_8778,N_8950);
nor U9145 (N_9145,N_8827,N_8764);
nand U9146 (N_9146,N_8981,N_8835);
and U9147 (N_9147,N_8936,N_8711);
and U9148 (N_9148,N_8909,N_8803);
or U9149 (N_9149,N_8930,N_8732);
nand U9150 (N_9150,N_8754,N_8973);
and U9151 (N_9151,N_8786,N_8709);
xor U9152 (N_9152,N_8810,N_8988);
nor U9153 (N_9153,N_8856,N_8861);
and U9154 (N_9154,N_8888,N_8955);
xor U9155 (N_9155,N_8954,N_8727);
xor U9156 (N_9156,N_8946,N_8851);
nor U9157 (N_9157,N_8790,N_8971);
nor U9158 (N_9158,N_8947,N_8763);
xnor U9159 (N_9159,N_8894,N_8813);
or U9160 (N_9160,N_8930,N_8936);
xor U9161 (N_9161,N_8796,N_8984);
nor U9162 (N_9162,N_8764,N_8872);
and U9163 (N_9163,N_8911,N_8780);
nand U9164 (N_9164,N_8942,N_8983);
xor U9165 (N_9165,N_8751,N_8882);
nor U9166 (N_9166,N_8953,N_8764);
and U9167 (N_9167,N_8782,N_8976);
and U9168 (N_9168,N_8700,N_8900);
xnor U9169 (N_9169,N_8741,N_8732);
and U9170 (N_9170,N_8878,N_8949);
xnor U9171 (N_9171,N_8757,N_8834);
or U9172 (N_9172,N_8747,N_8997);
nor U9173 (N_9173,N_8716,N_8836);
or U9174 (N_9174,N_8740,N_8942);
nand U9175 (N_9175,N_8842,N_8826);
and U9176 (N_9176,N_8921,N_8933);
nor U9177 (N_9177,N_8828,N_8938);
or U9178 (N_9178,N_8916,N_8984);
nor U9179 (N_9179,N_8702,N_8953);
and U9180 (N_9180,N_8890,N_8815);
nor U9181 (N_9181,N_8968,N_8932);
and U9182 (N_9182,N_8814,N_8989);
and U9183 (N_9183,N_8933,N_8887);
or U9184 (N_9184,N_8945,N_8752);
and U9185 (N_9185,N_8939,N_8912);
xnor U9186 (N_9186,N_8814,N_8703);
nor U9187 (N_9187,N_8956,N_8972);
nand U9188 (N_9188,N_8809,N_8832);
and U9189 (N_9189,N_8998,N_8847);
and U9190 (N_9190,N_8929,N_8759);
nor U9191 (N_9191,N_8825,N_8780);
nor U9192 (N_9192,N_8842,N_8718);
and U9193 (N_9193,N_8861,N_8768);
nor U9194 (N_9194,N_8845,N_8783);
nor U9195 (N_9195,N_8866,N_8706);
nor U9196 (N_9196,N_8800,N_8829);
or U9197 (N_9197,N_8990,N_8744);
xnor U9198 (N_9198,N_8834,N_8740);
and U9199 (N_9199,N_8893,N_8979);
or U9200 (N_9200,N_8810,N_8787);
xor U9201 (N_9201,N_8982,N_8913);
nor U9202 (N_9202,N_8884,N_8992);
nor U9203 (N_9203,N_8794,N_8971);
and U9204 (N_9204,N_8886,N_8922);
nand U9205 (N_9205,N_8852,N_8827);
xnor U9206 (N_9206,N_8997,N_8716);
nand U9207 (N_9207,N_8710,N_8755);
xnor U9208 (N_9208,N_8844,N_8864);
nand U9209 (N_9209,N_8909,N_8929);
nand U9210 (N_9210,N_8779,N_8700);
nand U9211 (N_9211,N_8990,N_8937);
xor U9212 (N_9212,N_8716,N_8919);
or U9213 (N_9213,N_8821,N_8925);
nand U9214 (N_9214,N_8918,N_8867);
xnor U9215 (N_9215,N_8983,N_8810);
and U9216 (N_9216,N_8805,N_8738);
xnor U9217 (N_9217,N_8704,N_8938);
nor U9218 (N_9218,N_8730,N_8784);
nor U9219 (N_9219,N_8746,N_8808);
or U9220 (N_9220,N_8978,N_8908);
or U9221 (N_9221,N_8783,N_8708);
and U9222 (N_9222,N_8823,N_8857);
nor U9223 (N_9223,N_8942,N_8799);
or U9224 (N_9224,N_8958,N_8771);
or U9225 (N_9225,N_8734,N_8815);
xor U9226 (N_9226,N_8852,N_8876);
and U9227 (N_9227,N_8841,N_8706);
xor U9228 (N_9228,N_8909,N_8709);
or U9229 (N_9229,N_8892,N_8766);
xnor U9230 (N_9230,N_8703,N_8764);
or U9231 (N_9231,N_8960,N_8969);
xnor U9232 (N_9232,N_8781,N_8942);
xor U9233 (N_9233,N_8940,N_8961);
nand U9234 (N_9234,N_8933,N_8723);
nand U9235 (N_9235,N_8845,N_8987);
xor U9236 (N_9236,N_8878,N_8792);
or U9237 (N_9237,N_8937,N_8954);
nor U9238 (N_9238,N_8997,N_8833);
and U9239 (N_9239,N_8740,N_8735);
xnor U9240 (N_9240,N_8740,N_8728);
and U9241 (N_9241,N_8946,N_8837);
nor U9242 (N_9242,N_8999,N_8760);
or U9243 (N_9243,N_8709,N_8787);
and U9244 (N_9244,N_8804,N_8965);
xor U9245 (N_9245,N_8804,N_8973);
and U9246 (N_9246,N_8849,N_8776);
and U9247 (N_9247,N_8951,N_8934);
or U9248 (N_9248,N_8772,N_8793);
xnor U9249 (N_9249,N_8771,N_8880);
xnor U9250 (N_9250,N_8761,N_8728);
xor U9251 (N_9251,N_8706,N_8969);
and U9252 (N_9252,N_8824,N_8907);
nand U9253 (N_9253,N_8902,N_8700);
nor U9254 (N_9254,N_8796,N_8815);
and U9255 (N_9255,N_8870,N_8896);
nand U9256 (N_9256,N_8741,N_8875);
nand U9257 (N_9257,N_8820,N_8889);
or U9258 (N_9258,N_8872,N_8793);
nor U9259 (N_9259,N_8897,N_8878);
or U9260 (N_9260,N_8863,N_8773);
xor U9261 (N_9261,N_8787,N_8737);
nand U9262 (N_9262,N_8797,N_8840);
nor U9263 (N_9263,N_8838,N_8839);
nand U9264 (N_9264,N_8794,N_8743);
xor U9265 (N_9265,N_8945,N_8972);
or U9266 (N_9266,N_8899,N_8966);
nor U9267 (N_9267,N_8947,N_8747);
nor U9268 (N_9268,N_8880,N_8891);
xor U9269 (N_9269,N_8756,N_8861);
nor U9270 (N_9270,N_8926,N_8790);
nand U9271 (N_9271,N_8875,N_8867);
nand U9272 (N_9272,N_8765,N_8924);
xor U9273 (N_9273,N_8802,N_8758);
or U9274 (N_9274,N_8826,N_8847);
nor U9275 (N_9275,N_8760,N_8759);
and U9276 (N_9276,N_8923,N_8801);
or U9277 (N_9277,N_8770,N_8873);
or U9278 (N_9278,N_8790,N_8800);
or U9279 (N_9279,N_8721,N_8877);
nand U9280 (N_9280,N_8757,N_8935);
xnor U9281 (N_9281,N_8776,N_8854);
nand U9282 (N_9282,N_8967,N_8755);
nor U9283 (N_9283,N_8765,N_8820);
and U9284 (N_9284,N_8929,N_8944);
xnor U9285 (N_9285,N_8908,N_8773);
xor U9286 (N_9286,N_8778,N_8998);
xor U9287 (N_9287,N_8859,N_8720);
or U9288 (N_9288,N_8900,N_8728);
nand U9289 (N_9289,N_8749,N_8947);
or U9290 (N_9290,N_8843,N_8743);
and U9291 (N_9291,N_8730,N_8875);
xnor U9292 (N_9292,N_8921,N_8943);
xor U9293 (N_9293,N_8732,N_8885);
xor U9294 (N_9294,N_8854,N_8778);
and U9295 (N_9295,N_8765,N_8960);
and U9296 (N_9296,N_8870,N_8991);
or U9297 (N_9297,N_8787,N_8999);
xor U9298 (N_9298,N_8962,N_8837);
or U9299 (N_9299,N_8831,N_8702);
nand U9300 (N_9300,N_9147,N_9226);
and U9301 (N_9301,N_9084,N_9053);
or U9302 (N_9302,N_9250,N_9006);
or U9303 (N_9303,N_9140,N_9034);
nor U9304 (N_9304,N_9012,N_9054);
nand U9305 (N_9305,N_9260,N_9214);
and U9306 (N_9306,N_9058,N_9121);
nor U9307 (N_9307,N_9025,N_9048);
xor U9308 (N_9308,N_9127,N_9029);
and U9309 (N_9309,N_9021,N_9130);
and U9310 (N_9310,N_9016,N_9107);
xor U9311 (N_9311,N_9114,N_9112);
or U9312 (N_9312,N_9266,N_9262);
xnor U9313 (N_9313,N_9027,N_9254);
nand U9314 (N_9314,N_9145,N_9106);
nor U9315 (N_9315,N_9065,N_9292);
xnor U9316 (N_9316,N_9185,N_9208);
or U9317 (N_9317,N_9216,N_9083);
and U9318 (N_9318,N_9090,N_9150);
or U9319 (N_9319,N_9033,N_9204);
or U9320 (N_9320,N_9222,N_9004);
nor U9321 (N_9321,N_9035,N_9026);
and U9322 (N_9322,N_9077,N_9115);
xnor U9323 (N_9323,N_9142,N_9086);
nand U9324 (N_9324,N_9126,N_9186);
xor U9325 (N_9325,N_9201,N_9218);
and U9326 (N_9326,N_9246,N_9171);
xor U9327 (N_9327,N_9244,N_9211);
and U9328 (N_9328,N_9087,N_9091);
nor U9329 (N_9329,N_9129,N_9265);
nor U9330 (N_9330,N_9093,N_9041);
nand U9331 (N_9331,N_9137,N_9269);
nor U9332 (N_9332,N_9072,N_9098);
xnor U9333 (N_9333,N_9227,N_9187);
nand U9334 (N_9334,N_9078,N_9299);
nand U9335 (N_9335,N_9020,N_9296);
or U9336 (N_9336,N_9135,N_9286);
nand U9337 (N_9337,N_9000,N_9096);
xor U9338 (N_9338,N_9195,N_9095);
nor U9339 (N_9339,N_9118,N_9003);
and U9340 (N_9340,N_9133,N_9298);
nand U9341 (N_9341,N_9148,N_9261);
and U9342 (N_9342,N_9040,N_9253);
and U9343 (N_9343,N_9125,N_9258);
and U9344 (N_9344,N_9276,N_9223);
nand U9345 (N_9345,N_9277,N_9167);
or U9346 (N_9346,N_9024,N_9110);
nor U9347 (N_9347,N_9295,N_9213);
nand U9348 (N_9348,N_9032,N_9113);
nand U9349 (N_9349,N_9022,N_9184);
or U9350 (N_9350,N_9289,N_9071);
xor U9351 (N_9351,N_9255,N_9238);
nor U9352 (N_9352,N_9203,N_9144);
and U9353 (N_9353,N_9281,N_9215);
and U9354 (N_9354,N_9177,N_9220);
or U9355 (N_9355,N_9019,N_9263);
or U9356 (N_9356,N_9179,N_9189);
and U9357 (N_9357,N_9156,N_9256);
nor U9358 (N_9358,N_9120,N_9092);
and U9359 (N_9359,N_9221,N_9068);
xor U9360 (N_9360,N_9094,N_9075);
or U9361 (N_9361,N_9067,N_9271);
xor U9362 (N_9362,N_9108,N_9267);
nor U9363 (N_9363,N_9105,N_9264);
nor U9364 (N_9364,N_9097,N_9057);
nor U9365 (N_9365,N_9206,N_9007);
nand U9366 (N_9366,N_9044,N_9070);
xnor U9367 (N_9367,N_9224,N_9194);
or U9368 (N_9368,N_9005,N_9198);
or U9369 (N_9369,N_9045,N_9039);
nand U9370 (N_9370,N_9212,N_9013);
xnor U9371 (N_9371,N_9297,N_9285);
xor U9372 (N_9372,N_9131,N_9104);
nor U9373 (N_9373,N_9178,N_9017);
xnor U9374 (N_9374,N_9279,N_9011);
nor U9375 (N_9375,N_9200,N_9123);
nor U9376 (N_9376,N_9259,N_9138);
or U9377 (N_9377,N_9089,N_9042);
and U9378 (N_9378,N_9190,N_9152);
xor U9379 (N_9379,N_9225,N_9136);
nor U9380 (N_9380,N_9196,N_9273);
nor U9381 (N_9381,N_9085,N_9073);
and U9382 (N_9382,N_9270,N_9111);
and U9383 (N_9383,N_9088,N_9160);
nand U9384 (N_9384,N_9066,N_9237);
and U9385 (N_9385,N_9280,N_9052);
nand U9386 (N_9386,N_9240,N_9268);
xor U9387 (N_9387,N_9182,N_9243);
nand U9388 (N_9388,N_9294,N_9124);
nor U9389 (N_9389,N_9282,N_9175);
and U9390 (N_9390,N_9063,N_9008);
and U9391 (N_9391,N_9101,N_9217);
or U9392 (N_9392,N_9010,N_9275);
nor U9393 (N_9393,N_9151,N_9274);
xor U9394 (N_9394,N_9193,N_9015);
or U9395 (N_9395,N_9119,N_9134);
nand U9396 (N_9396,N_9023,N_9009);
xnor U9397 (N_9397,N_9031,N_9049);
and U9398 (N_9398,N_9290,N_9231);
or U9399 (N_9399,N_9103,N_9219);
or U9400 (N_9400,N_9199,N_9074);
xor U9401 (N_9401,N_9166,N_9176);
nor U9402 (N_9402,N_9146,N_9191);
nor U9403 (N_9403,N_9149,N_9001);
or U9404 (N_9404,N_9170,N_9228);
xor U9405 (N_9405,N_9233,N_9247);
nand U9406 (N_9406,N_9172,N_9163);
nor U9407 (N_9407,N_9153,N_9230);
nor U9408 (N_9408,N_9205,N_9173);
nor U9409 (N_9409,N_9080,N_9252);
and U9410 (N_9410,N_9037,N_9272);
or U9411 (N_9411,N_9062,N_9002);
or U9412 (N_9412,N_9209,N_9229);
nand U9413 (N_9413,N_9030,N_9291);
and U9414 (N_9414,N_9141,N_9079);
and U9415 (N_9415,N_9159,N_9056);
nor U9416 (N_9416,N_9241,N_9197);
and U9417 (N_9417,N_9038,N_9287);
and U9418 (N_9418,N_9014,N_9249);
nor U9419 (N_9419,N_9180,N_9245);
nor U9420 (N_9420,N_9234,N_9059);
xor U9421 (N_9421,N_9161,N_9102);
xor U9422 (N_9422,N_9082,N_9069);
xor U9423 (N_9423,N_9143,N_9100);
and U9424 (N_9424,N_9181,N_9164);
nor U9425 (N_9425,N_9248,N_9202);
or U9426 (N_9426,N_9018,N_9155);
nand U9427 (N_9427,N_9157,N_9128);
nor U9428 (N_9428,N_9278,N_9081);
nor U9429 (N_9429,N_9242,N_9117);
and U9430 (N_9430,N_9109,N_9165);
and U9431 (N_9431,N_9099,N_9183);
or U9432 (N_9432,N_9064,N_9283);
xor U9433 (N_9433,N_9188,N_9288);
and U9434 (N_9434,N_9116,N_9046);
xor U9435 (N_9435,N_9284,N_9192);
or U9436 (N_9436,N_9061,N_9236);
nand U9437 (N_9437,N_9257,N_9207);
nor U9438 (N_9438,N_9043,N_9139);
and U9439 (N_9439,N_9174,N_9158);
or U9440 (N_9440,N_9239,N_9036);
nor U9441 (N_9441,N_9051,N_9028);
nand U9442 (N_9442,N_9293,N_9122);
nand U9443 (N_9443,N_9232,N_9076);
nand U9444 (N_9444,N_9050,N_9047);
and U9445 (N_9445,N_9251,N_9132);
nand U9446 (N_9446,N_9168,N_9055);
xor U9447 (N_9447,N_9154,N_9162);
nand U9448 (N_9448,N_9235,N_9210);
nor U9449 (N_9449,N_9060,N_9169);
nand U9450 (N_9450,N_9297,N_9092);
nand U9451 (N_9451,N_9171,N_9276);
nand U9452 (N_9452,N_9114,N_9019);
xnor U9453 (N_9453,N_9282,N_9007);
xnor U9454 (N_9454,N_9223,N_9266);
nor U9455 (N_9455,N_9055,N_9262);
and U9456 (N_9456,N_9286,N_9208);
or U9457 (N_9457,N_9220,N_9053);
or U9458 (N_9458,N_9188,N_9276);
xnor U9459 (N_9459,N_9272,N_9005);
nor U9460 (N_9460,N_9155,N_9195);
xnor U9461 (N_9461,N_9192,N_9255);
nand U9462 (N_9462,N_9261,N_9047);
nor U9463 (N_9463,N_9027,N_9046);
and U9464 (N_9464,N_9118,N_9254);
nor U9465 (N_9465,N_9185,N_9068);
nand U9466 (N_9466,N_9227,N_9079);
or U9467 (N_9467,N_9080,N_9009);
and U9468 (N_9468,N_9146,N_9247);
xor U9469 (N_9469,N_9028,N_9001);
or U9470 (N_9470,N_9029,N_9146);
xnor U9471 (N_9471,N_9112,N_9063);
nor U9472 (N_9472,N_9240,N_9261);
nor U9473 (N_9473,N_9092,N_9139);
and U9474 (N_9474,N_9286,N_9253);
nand U9475 (N_9475,N_9208,N_9189);
or U9476 (N_9476,N_9048,N_9059);
nor U9477 (N_9477,N_9281,N_9116);
nor U9478 (N_9478,N_9204,N_9121);
nor U9479 (N_9479,N_9168,N_9029);
nand U9480 (N_9480,N_9177,N_9250);
xor U9481 (N_9481,N_9083,N_9263);
nand U9482 (N_9482,N_9241,N_9262);
xnor U9483 (N_9483,N_9288,N_9017);
nand U9484 (N_9484,N_9232,N_9125);
xnor U9485 (N_9485,N_9197,N_9080);
xor U9486 (N_9486,N_9120,N_9041);
nand U9487 (N_9487,N_9041,N_9284);
and U9488 (N_9488,N_9233,N_9177);
and U9489 (N_9489,N_9246,N_9279);
nor U9490 (N_9490,N_9244,N_9118);
nand U9491 (N_9491,N_9224,N_9153);
nand U9492 (N_9492,N_9039,N_9023);
or U9493 (N_9493,N_9113,N_9292);
nor U9494 (N_9494,N_9293,N_9238);
nand U9495 (N_9495,N_9225,N_9061);
or U9496 (N_9496,N_9004,N_9063);
nand U9497 (N_9497,N_9221,N_9104);
nand U9498 (N_9498,N_9066,N_9000);
or U9499 (N_9499,N_9154,N_9275);
or U9500 (N_9500,N_9157,N_9211);
xor U9501 (N_9501,N_9252,N_9074);
or U9502 (N_9502,N_9264,N_9132);
nor U9503 (N_9503,N_9018,N_9072);
or U9504 (N_9504,N_9076,N_9089);
or U9505 (N_9505,N_9064,N_9062);
or U9506 (N_9506,N_9066,N_9292);
or U9507 (N_9507,N_9111,N_9231);
nand U9508 (N_9508,N_9262,N_9027);
nor U9509 (N_9509,N_9175,N_9010);
nor U9510 (N_9510,N_9220,N_9128);
nand U9511 (N_9511,N_9210,N_9005);
xor U9512 (N_9512,N_9109,N_9255);
or U9513 (N_9513,N_9097,N_9040);
nor U9514 (N_9514,N_9137,N_9258);
xor U9515 (N_9515,N_9294,N_9275);
xnor U9516 (N_9516,N_9258,N_9069);
or U9517 (N_9517,N_9164,N_9016);
nand U9518 (N_9518,N_9111,N_9237);
nor U9519 (N_9519,N_9000,N_9176);
xnor U9520 (N_9520,N_9121,N_9137);
and U9521 (N_9521,N_9034,N_9101);
xor U9522 (N_9522,N_9252,N_9195);
nand U9523 (N_9523,N_9038,N_9153);
or U9524 (N_9524,N_9055,N_9266);
nor U9525 (N_9525,N_9224,N_9028);
xor U9526 (N_9526,N_9276,N_9214);
or U9527 (N_9527,N_9275,N_9183);
and U9528 (N_9528,N_9005,N_9264);
and U9529 (N_9529,N_9245,N_9207);
nor U9530 (N_9530,N_9102,N_9177);
or U9531 (N_9531,N_9220,N_9025);
or U9532 (N_9532,N_9195,N_9048);
nand U9533 (N_9533,N_9154,N_9009);
nor U9534 (N_9534,N_9017,N_9246);
or U9535 (N_9535,N_9218,N_9107);
and U9536 (N_9536,N_9222,N_9207);
xnor U9537 (N_9537,N_9217,N_9293);
nand U9538 (N_9538,N_9218,N_9050);
xor U9539 (N_9539,N_9127,N_9253);
xor U9540 (N_9540,N_9249,N_9139);
xnor U9541 (N_9541,N_9053,N_9234);
nand U9542 (N_9542,N_9225,N_9114);
nand U9543 (N_9543,N_9018,N_9168);
xnor U9544 (N_9544,N_9124,N_9292);
nand U9545 (N_9545,N_9037,N_9111);
or U9546 (N_9546,N_9062,N_9121);
xnor U9547 (N_9547,N_9128,N_9299);
and U9548 (N_9548,N_9271,N_9268);
or U9549 (N_9549,N_9082,N_9029);
nor U9550 (N_9550,N_9157,N_9238);
and U9551 (N_9551,N_9234,N_9102);
nor U9552 (N_9552,N_9069,N_9158);
and U9553 (N_9553,N_9010,N_9063);
nand U9554 (N_9554,N_9290,N_9159);
and U9555 (N_9555,N_9225,N_9084);
nor U9556 (N_9556,N_9212,N_9255);
and U9557 (N_9557,N_9247,N_9123);
and U9558 (N_9558,N_9027,N_9005);
or U9559 (N_9559,N_9125,N_9013);
xnor U9560 (N_9560,N_9172,N_9250);
nor U9561 (N_9561,N_9106,N_9203);
and U9562 (N_9562,N_9023,N_9113);
nor U9563 (N_9563,N_9173,N_9082);
nand U9564 (N_9564,N_9005,N_9010);
nor U9565 (N_9565,N_9123,N_9075);
and U9566 (N_9566,N_9170,N_9039);
xor U9567 (N_9567,N_9176,N_9102);
nand U9568 (N_9568,N_9183,N_9241);
nand U9569 (N_9569,N_9277,N_9273);
and U9570 (N_9570,N_9287,N_9007);
nor U9571 (N_9571,N_9112,N_9098);
nand U9572 (N_9572,N_9105,N_9100);
nor U9573 (N_9573,N_9055,N_9295);
nor U9574 (N_9574,N_9014,N_9090);
or U9575 (N_9575,N_9040,N_9064);
nand U9576 (N_9576,N_9204,N_9064);
nor U9577 (N_9577,N_9031,N_9116);
nor U9578 (N_9578,N_9253,N_9115);
or U9579 (N_9579,N_9121,N_9287);
xor U9580 (N_9580,N_9081,N_9245);
and U9581 (N_9581,N_9007,N_9084);
nand U9582 (N_9582,N_9090,N_9167);
nand U9583 (N_9583,N_9250,N_9058);
or U9584 (N_9584,N_9074,N_9140);
and U9585 (N_9585,N_9150,N_9139);
nor U9586 (N_9586,N_9031,N_9111);
and U9587 (N_9587,N_9281,N_9209);
xor U9588 (N_9588,N_9213,N_9212);
nor U9589 (N_9589,N_9208,N_9247);
nand U9590 (N_9590,N_9172,N_9200);
nand U9591 (N_9591,N_9133,N_9107);
nand U9592 (N_9592,N_9280,N_9041);
nand U9593 (N_9593,N_9077,N_9291);
nand U9594 (N_9594,N_9140,N_9147);
and U9595 (N_9595,N_9100,N_9010);
or U9596 (N_9596,N_9197,N_9253);
or U9597 (N_9597,N_9018,N_9066);
nand U9598 (N_9598,N_9275,N_9142);
xor U9599 (N_9599,N_9221,N_9297);
nand U9600 (N_9600,N_9589,N_9528);
nor U9601 (N_9601,N_9336,N_9433);
and U9602 (N_9602,N_9499,N_9300);
and U9603 (N_9603,N_9363,N_9548);
nand U9604 (N_9604,N_9399,N_9542);
or U9605 (N_9605,N_9532,N_9567);
and U9606 (N_9606,N_9397,N_9440);
xor U9607 (N_9607,N_9379,N_9438);
nor U9608 (N_9608,N_9467,N_9412);
nand U9609 (N_9609,N_9387,N_9478);
nand U9610 (N_9610,N_9541,N_9486);
nand U9611 (N_9611,N_9577,N_9329);
nand U9612 (N_9612,N_9314,N_9385);
and U9613 (N_9613,N_9464,N_9504);
nand U9614 (N_9614,N_9351,N_9380);
nand U9615 (N_9615,N_9592,N_9367);
or U9616 (N_9616,N_9362,N_9318);
or U9617 (N_9617,N_9393,N_9304);
or U9618 (N_9618,N_9518,N_9372);
nor U9619 (N_9619,N_9580,N_9368);
nand U9620 (N_9620,N_9484,N_9461);
and U9621 (N_9621,N_9590,N_9466);
nand U9622 (N_9622,N_9340,N_9494);
or U9623 (N_9623,N_9563,N_9373);
and U9624 (N_9624,N_9509,N_9543);
xnor U9625 (N_9625,N_9396,N_9501);
xnor U9626 (N_9626,N_9417,N_9455);
and U9627 (N_9627,N_9488,N_9306);
or U9628 (N_9628,N_9346,N_9560);
xnor U9629 (N_9629,N_9549,N_9534);
or U9630 (N_9630,N_9526,N_9327);
nor U9631 (N_9631,N_9585,N_9578);
or U9632 (N_9632,N_9576,N_9334);
or U9633 (N_9633,N_9366,N_9521);
and U9634 (N_9634,N_9404,N_9452);
nor U9635 (N_9635,N_9448,N_9422);
xnor U9636 (N_9636,N_9591,N_9342);
nor U9637 (N_9637,N_9432,N_9538);
xor U9638 (N_9638,N_9558,N_9571);
and U9639 (N_9639,N_9505,N_9479);
nand U9640 (N_9640,N_9439,N_9490);
or U9641 (N_9641,N_9500,N_9321);
or U9642 (N_9642,N_9460,N_9398);
nor U9643 (N_9643,N_9594,N_9472);
nor U9644 (N_9644,N_9434,N_9361);
xor U9645 (N_9645,N_9312,N_9520);
nand U9646 (N_9646,N_9511,N_9529);
nand U9647 (N_9647,N_9575,N_9508);
nand U9648 (N_9648,N_9584,N_9454);
nor U9649 (N_9649,N_9553,N_9449);
nand U9650 (N_9650,N_9323,N_9487);
xnor U9651 (N_9651,N_9421,N_9507);
xnor U9652 (N_9652,N_9371,N_9309);
and U9653 (N_9653,N_9395,N_9502);
xor U9654 (N_9654,N_9554,N_9583);
xnor U9655 (N_9655,N_9442,N_9358);
nand U9656 (N_9656,N_9572,N_9311);
xor U9657 (N_9657,N_9330,N_9527);
or U9658 (N_9658,N_9431,N_9565);
nand U9659 (N_9659,N_9463,N_9418);
nor U9660 (N_9660,N_9392,N_9447);
and U9661 (N_9661,N_9485,N_9536);
nand U9662 (N_9662,N_9525,N_9471);
xor U9663 (N_9663,N_9531,N_9459);
nand U9664 (N_9664,N_9493,N_9364);
nand U9665 (N_9665,N_9310,N_9474);
or U9666 (N_9666,N_9561,N_9383);
and U9667 (N_9667,N_9517,N_9374);
xor U9668 (N_9668,N_9595,N_9569);
and U9669 (N_9669,N_9557,N_9353);
or U9670 (N_9670,N_9551,N_9313);
nand U9671 (N_9671,N_9350,N_9339);
and U9672 (N_9672,N_9552,N_9457);
nor U9673 (N_9673,N_9319,N_9437);
nand U9674 (N_9674,N_9445,N_9491);
nor U9675 (N_9675,N_9365,N_9302);
and U9676 (N_9676,N_9419,N_9355);
or U9677 (N_9677,N_9483,N_9430);
or U9678 (N_9678,N_9506,N_9359);
or U9679 (N_9679,N_9545,N_9475);
or U9680 (N_9680,N_9377,N_9382);
xnor U9681 (N_9681,N_9320,N_9405);
nor U9682 (N_9682,N_9559,N_9489);
xnor U9683 (N_9683,N_9523,N_9599);
nand U9684 (N_9684,N_9562,N_9325);
nor U9685 (N_9685,N_9401,N_9436);
or U9686 (N_9686,N_9587,N_9441);
xor U9687 (N_9687,N_9515,N_9435);
and U9688 (N_9688,N_9579,N_9588);
xor U9689 (N_9689,N_9573,N_9316);
or U9690 (N_9690,N_9547,N_9376);
xnor U9691 (N_9691,N_9301,N_9391);
and U9692 (N_9692,N_9451,N_9423);
or U9693 (N_9693,N_9386,N_9369);
nand U9694 (N_9694,N_9513,N_9324);
nor U9695 (N_9695,N_9582,N_9349);
nand U9696 (N_9696,N_9307,N_9408);
or U9697 (N_9697,N_9348,N_9535);
nand U9698 (N_9698,N_9413,N_9544);
and U9699 (N_9699,N_9596,N_9522);
nor U9700 (N_9700,N_9458,N_9469);
or U9701 (N_9701,N_9411,N_9403);
xnor U9702 (N_9702,N_9537,N_9514);
or U9703 (N_9703,N_9406,N_9378);
and U9704 (N_9704,N_9356,N_9428);
xor U9705 (N_9705,N_9556,N_9473);
xnor U9706 (N_9706,N_9429,N_9384);
xor U9707 (N_9707,N_9344,N_9597);
or U9708 (N_9708,N_9328,N_9568);
nand U9709 (N_9709,N_9519,N_9381);
xor U9710 (N_9710,N_9453,N_9414);
and U9711 (N_9711,N_9495,N_9546);
nand U9712 (N_9712,N_9352,N_9477);
and U9713 (N_9713,N_9400,N_9415);
or U9714 (N_9714,N_9416,N_9496);
or U9715 (N_9715,N_9388,N_9354);
xnor U9716 (N_9716,N_9555,N_9390);
xor U9717 (N_9717,N_9394,N_9375);
nor U9718 (N_9718,N_9510,N_9539);
and U9719 (N_9719,N_9443,N_9332);
nor U9720 (N_9720,N_9409,N_9343);
and U9721 (N_9721,N_9424,N_9426);
or U9722 (N_9722,N_9326,N_9512);
nor U9723 (N_9723,N_9516,N_9550);
or U9724 (N_9724,N_9598,N_9462);
xnor U9725 (N_9725,N_9303,N_9465);
xor U9726 (N_9726,N_9315,N_9425);
xnor U9727 (N_9727,N_9533,N_9476);
nand U9728 (N_9728,N_9407,N_9492);
or U9729 (N_9729,N_9389,N_9574);
or U9730 (N_9730,N_9481,N_9333);
or U9731 (N_9731,N_9498,N_9480);
nor U9732 (N_9732,N_9420,N_9570);
nand U9733 (N_9733,N_9450,N_9497);
nand U9734 (N_9734,N_9357,N_9337);
or U9735 (N_9735,N_9593,N_9468);
nor U9736 (N_9736,N_9370,N_9566);
and U9737 (N_9737,N_9410,N_9524);
or U9738 (N_9738,N_9586,N_9345);
or U9739 (N_9739,N_9503,N_9308);
or U9740 (N_9740,N_9470,N_9402);
nor U9741 (N_9741,N_9564,N_9317);
and U9742 (N_9742,N_9540,N_9446);
nor U9743 (N_9743,N_9347,N_9322);
and U9744 (N_9744,N_9581,N_9456);
or U9745 (N_9745,N_9444,N_9305);
and U9746 (N_9746,N_9335,N_9530);
xor U9747 (N_9747,N_9341,N_9360);
or U9748 (N_9748,N_9331,N_9338);
nor U9749 (N_9749,N_9427,N_9482);
xnor U9750 (N_9750,N_9510,N_9400);
or U9751 (N_9751,N_9478,N_9551);
and U9752 (N_9752,N_9379,N_9376);
xor U9753 (N_9753,N_9591,N_9334);
xnor U9754 (N_9754,N_9409,N_9444);
nor U9755 (N_9755,N_9309,N_9342);
and U9756 (N_9756,N_9301,N_9579);
nand U9757 (N_9757,N_9525,N_9440);
nand U9758 (N_9758,N_9490,N_9374);
nand U9759 (N_9759,N_9436,N_9439);
xnor U9760 (N_9760,N_9486,N_9460);
and U9761 (N_9761,N_9350,N_9337);
nand U9762 (N_9762,N_9502,N_9572);
nor U9763 (N_9763,N_9375,N_9515);
or U9764 (N_9764,N_9301,N_9496);
or U9765 (N_9765,N_9455,N_9543);
xor U9766 (N_9766,N_9571,N_9417);
nor U9767 (N_9767,N_9507,N_9524);
or U9768 (N_9768,N_9507,N_9328);
xor U9769 (N_9769,N_9351,N_9596);
nor U9770 (N_9770,N_9520,N_9577);
xnor U9771 (N_9771,N_9423,N_9332);
xor U9772 (N_9772,N_9485,N_9489);
nand U9773 (N_9773,N_9583,N_9547);
xnor U9774 (N_9774,N_9428,N_9403);
or U9775 (N_9775,N_9442,N_9557);
or U9776 (N_9776,N_9391,N_9426);
and U9777 (N_9777,N_9485,N_9483);
or U9778 (N_9778,N_9313,N_9437);
nor U9779 (N_9779,N_9595,N_9352);
nor U9780 (N_9780,N_9333,N_9529);
or U9781 (N_9781,N_9560,N_9543);
xor U9782 (N_9782,N_9387,N_9518);
or U9783 (N_9783,N_9547,N_9543);
nand U9784 (N_9784,N_9430,N_9477);
nor U9785 (N_9785,N_9449,N_9303);
or U9786 (N_9786,N_9583,N_9407);
xor U9787 (N_9787,N_9509,N_9381);
xnor U9788 (N_9788,N_9479,N_9301);
and U9789 (N_9789,N_9352,N_9598);
and U9790 (N_9790,N_9454,N_9350);
nand U9791 (N_9791,N_9410,N_9389);
nand U9792 (N_9792,N_9570,N_9355);
and U9793 (N_9793,N_9536,N_9451);
nand U9794 (N_9794,N_9471,N_9349);
xnor U9795 (N_9795,N_9491,N_9338);
or U9796 (N_9796,N_9399,N_9591);
and U9797 (N_9797,N_9427,N_9435);
nand U9798 (N_9798,N_9321,N_9322);
and U9799 (N_9799,N_9421,N_9560);
nand U9800 (N_9800,N_9408,N_9374);
nand U9801 (N_9801,N_9436,N_9345);
xor U9802 (N_9802,N_9328,N_9334);
xnor U9803 (N_9803,N_9377,N_9535);
xor U9804 (N_9804,N_9356,N_9307);
or U9805 (N_9805,N_9549,N_9506);
or U9806 (N_9806,N_9326,N_9433);
nor U9807 (N_9807,N_9573,N_9486);
and U9808 (N_9808,N_9485,N_9372);
xnor U9809 (N_9809,N_9439,N_9529);
nor U9810 (N_9810,N_9492,N_9547);
xnor U9811 (N_9811,N_9494,N_9496);
nand U9812 (N_9812,N_9467,N_9339);
xor U9813 (N_9813,N_9577,N_9378);
or U9814 (N_9814,N_9394,N_9417);
xnor U9815 (N_9815,N_9475,N_9368);
nand U9816 (N_9816,N_9317,N_9582);
nand U9817 (N_9817,N_9482,N_9458);
xor U9818 (N_9818,N_9411,N_9496);
nor U9819 (N_9819,N_9412,N_9528);
or U9820 (N_9820,N_9531,N_9321);
nand U9821 (N_9821,N_9337,N_9540);
nor U9822 (N_9822,N_9305,N_9566);
xnor U9823 (N_9823,N_9550,N_9467);
and U9824 (N_9824,N_9493,N_9441);
nor U9825 (N_9825,N_9519,N_9563);
xnor U9826 (N_9826,N_9432,N_9565);
nor U9827 (N_9827,N_9334,N_9575);
nor U9828 (N_9828,N_9549,N_9569);
and U9829 (N_9829,N_9414,N_9549);
nor U9830 (N_9830,N_9468,N_9584);
nor U9831 (N_9831,N_9530,N_9458);
or U9832 (N_9832,N_9364,N_9574);
or U9833 (N_9833,N_9419,N_9467);
or U9834 (N_9834,N_9377,N_9315);
xnor U9835 (N_9835,N_9313,N_9552);
nand U9836 (N_9836,N_9502,N_9506);
or U9837 (N_9837,N_9526,N_9511);
and U9838 (N_9838,N_9599,N_9453);
nor U9839 (N_9839,N_9439,N_9401);
or U9840 (N_9840,N_9333,N_9532);
xnor U9841 (N_9841,N_9459,N_9432);
or U9842 (N_9842,N_9577,N_9499);
or U9843 (N_9843,N_9446,N_9583);
or U9844 (N_9844,N_9412,N_9333);
xnor U9845 (N_9845,N_9367,N_9528);
nand U9846 (N_9846,N_9390,N_9563);
nor U9847 (N_9847,N_9364,N_9486);
and U9848 (N_9848,N_9461,N_9338);
nand U9849 (N_9849,N_9501,N_9524);
xnor U9850 (N_9850,N_9469,N_9498);
nand U9851 (N_9851,N_9566,N_9301);
or U9852 (N_9852,N_9411,N_9569);
xor U9853 (N_9853,N_9533,N_9414);
nor U9854 (N_9854,N_9554,N_9366);
or U9855 (N_9855,N_9498,N_9489);
xnor U9856 (N_9856,N_9567,N_9472);
or U9857 (N_9857,N_9408,N_9493);
and U9858 (N_9858,N_9463,N_9401);
xnor U9859 (N_9859,N_9471,N_9338);
or U9860 (N_9860,N_9542,N_9596);
xnor U9861 (N_9861,N_9332,N_9334);
nor U9862 (N_9862,N_9594,N_9459);
nor U9863 (N_9863,N_9447,N_9467);
or U9864 (N_9864,N_9430,N_9563);
or U9865 (N_9865,N_9451,N_9580);
xor U9866 (N_9866,N_9342,N_9404);
or U9867 (N_9867,N_9558,N_9579);
xnor U9868 (N_9868,N_9496,N_9433);
nand U9869 (N_9869,N_9460,N_9525);
xnor U9870 (N_9870,N_9351,N_9498);
or U9871 (N_9871,N_9550,N_9554);
nor U9872 (N_9872,N_9530,N_9422);
nand U9873 (N_9873,N_9331,N_9554);
xnor U9874 (N_9874,N_9581,N_9531);
nand U9875 (N_9875,N_9440,N_9595);
xor U9876 (N_9876,N_9465,N_9364);
xnor U9877 (N_9877,N_9456,N_9476);
xnor U9878 (N_9878,N_9430,N_9468);
xor U9879 (N_9879,N_9458,N_9426);
xor U9880 (N_9880,N_9547,N_9561);
nand U9881 (N_9881,N_9358,N_9514);
or U9882 (N_9882,N_9564,N_9326);
nand U9883 (N_9883,N_9514,N_9480);
xnor U9884 (N_9884,N_9590,N_9492);
and U9885 (N_9885,N_9362,N_9423);
or U9886 (N_9886,N_9466,N_9477);
nand U9887 (N_9887,N_9521,N_9526);
and U9888 (N_9888,N_9458,N_9563);
or U9889 (N_9889,N_9572,N_9351);
or U9890 (N_9890,N_9468,N_9336);
and U9891 (N_9891,N_9415,N_9570);
nor U9892 (N_9892,N_9496,N_9597);
and U9893 (N_9893,N_9549,N_9393);
or U9894 (N_9894,N_9324,N_9353);
nor U9895 (N_9895,N_9574,N_9583);
xnor U9896 (N_9896,N_9363,N_9345);
nor U9897 (N_9897,N_9561,N_9570);
xor U9898 (N_9898,N_9455,N_9537);
nor U9899 (N_9899,N_9490,N_9337);
nor U9900 (N_9900,N_9611,N_9815);
nor U9901 (N_9901,N_9770,N_9736);
nand U9902 (N_9902,N_9795,N_9867);
xnor U9903 (N_9903,N_9699,N_9666);
nand U9904 (N_9904,N_9608,N_9631);
nand U9905 (N_9905,N_9771,N_9723);
or U9906 (N_9906,N_9703,N_9683);
and U9907 (N_9907,N_9711,N_9756);
nand U9908 (N_9908,N_9809,N_9724);
xnor U9909 (N_9909,N_9899,N_9757);
nand U9910 (N_9910,N_9602,N_9646);
and U9911 (N_9911,N_9744,N_9836);
or U9912 (N_9912,N_9876,N_9896);
and U9913 (N_9913,N_9701,N_9743);
nor U9914 (N_9914,N_9676,N_9655);
nor U9915 (N_9915,N_9654,N_9621);
nor U9916 (N_9916,N_9812,N_9847);
and U9917 (N_9917,N_9720,N_9615);
xnor U9918 (N_9918,N_9708,N_9633);
and U9919 (N_9919,N_9816,N_9868);
and U9920 (N_9920,N_9688,N_9763);
xor U9921 (N_9921,N_9609,N_9617);
and U9922 (N_9922,N_9828,N_9789);
and U9923 (N_9923,N_9751,N_9832);
nand U9924 (N_9924,N_9728,N_9883);
nand U9925 (N_9925,N_9840,N_9861);
and U9926 (N_9926,N_9650,N_9833);
nand U9927 (N_9927,N_9811,N_9665);
nor U9928 (N_9928,N_9792,N_9645);
and U9929 (N_9929,N_9680,N_9897);
and U9930 (N_9930,N_9664,N_9801);
xor U9931 (N_9931,N_9613,N_9707);
xor U9932 (N_9932,N_9694,N_9855);
or U9933 (N_9933,N_9852,N_9745);
nor U9934 (N_9934,N_9643,N_9618);
nand U9935 (N_9935,N_9869,N_9777);
nand U9936 (N_9936,N_9865,N_9780);
nand U9937 (N_9937,N_9835,N_9870);
xor U9938 (N_9938,N_9857,N_9704);
or U9939 (N_9939,N_9839,N_9651);
xor U9940 (N_9940,N_9829,N_9748);
nor U9941 (N_9941,N_9796,N_9843);
nand U9942 (N_9942,N_9878,N_9649);
nand U9943 (N_9943,N_9894,N_9798);
nor U9944 (N_9944,N_9671,N_9690);
nor U9945 (N_9945,N_9605,N_9717);
nor U9946 (N_9946,N_9725,N_9722);
nand U9947 (N_9947,N_9766,N_9802);
xor U9948 (N_9948,N_9691,N_9889);
nor U9949 (N_9949,N_9797,N_9612);
nor U9950 (N_9950,N_9682,N_9788);
nand U9951 (N_9951,N_9884,N_9875);
or U9952 (N_9952,N_9679,N_9877);
nor U9953 (N_9953,N_9656,N_9782);
nor U9954 (N_9954,N_9641,N_9854);
xor U9955 (N_9955,N_9686,N_9898);
xnor U9956 (N_9956,N_9652,N_9885);
xnor U9957 (N_9957,N_9698,N_9759);
and U9958 (N_9958,N_9862,N_9838);
xnor U9959 (N_9959,N_9687,N_9604);
xor U9960 (N_9960,N_9719,N_9781);
and U9961 (N_9961,N_9783,N_9726);
or U9962 (N_9962,N_9639,N_9776);
and U9963 (N_9963,N_9733,N_9860);
nor U9964 (N_9964,N_9681,N_9871);
xor U9965 (N_9965,N_9805,N_9662);
or U9966 (N_9966,N_9856,N_9842);
or U9967 (N_9967,N_9647,N_9768);
or U9968 (N_9968,N_9834,N_9706);
and U9969 (N_9969,N_9762,N_9734);
nand U9970 (N_9970,N_9684,N_9859);
and U9971 (N_9971,N_9718,N_9674);
nor U9972 (N_9972,N_9661,N_9879);
or U9973 (N_9973,N_9830,N_9814);
nor U9974 (N_9974,N_9697,N_9845);
nor U9975 (N_9975,N_9755,N_9716);
nor U9976 (N_9976,N_9808,N_9807);
and U9977 (N_9977,N_9863,N_9713);
xor U9978 (N_9978,N_9761,N_9672);
and U9979 (N_9979,N_9626,N_9794);
or U9980 (N_9980,N_9764,N_9689);
and U9981 (N_9981,N_9741,N_9635);
nand U9982 (N_9982,N_9758,N_9872);
nor U9983 (N_9983,N_9750,N_9817);
nor U9984 (N_9984,N_9729,N_9601);
xor U9985 (N_9985,N_9873,N_9810);
or U9986 (N_9986,N_9784,N_9657);
nor U9987 (N_9987,N_9858,N_9790);
or U9988 (N_9988,N_9630,N_9831);
and U9989 (N_9989,N_9658,N_9769);
and U9990 (N_9990,N_9732,N_9846);
xnor U9991 (N_9991,N_9827,N_9880);
xnor U9992 (N_9992,N_9826,N_9774);
and U9993 (N_9993,N_9749,N_9712);
xnor U9994 (N_9994,N_9606,N_9739);
nand U9995 (N_9995,N_9642,N_9803);
and U9996 (N_9996,N_9709,N_9685);
nand U9997 (N_9997,N_9637,N_9648);
nor U9998 (N_9998,N_9632,N_9644);
or U9999 (N_9999,N_9752,N_9622);
nor U10000 (N_10000,N_9848,N_9787);
nor U10001 (N_10001,N_9746,N_9714);
nor U10002 (N_10002,N_9853,N_9786);
nand U10003 (N_10003,N_9735,N_9844);
or U10004 (N_10004,N_9804,N_9895);
and U10005 (N_10005,N_9673,N_9623);
or U10006 (N_10006,N_9821,N_9627);
or U10007 (N_10007,N_9737,N_9820);
nand U10008 (N_10008,N_9819,N_9628);
and U10009 (N_10009,N_9888,N_9603);
nor U10010 (N_10010,N_9669,N_9778);
or U10011 (N_10011,N_9696,N_9775);
and U10012 (N_10012,N_9721,N_9663);
nand U10013 (N_10013,N_9600,N_9710);
xnor U10014 (N_10014,N_9610,N_9753);
nand U10015 (N_10015,N_9629,N_9864);
or U10016 (N_10016,N_9693,N_9779);
xor U10017 (N_10017,N_9727,N_9823);
or U10018 (N_10018,N_9841,N_9675);
nor U10019 (N_10019,N_9791,N_9767);
and U10020 (N_10020,N_9730,N_9837);
nor U10021 (N_10021,N_9731,N_9893);
and U10022 (N_10022,N_9891,N_9634);
and U10023 (N_10023,N_9851,N_9670);
and U10024 (N_10024,N_9740,N_9793);
nand U10025 (N_10025,N_9818,N_9692);
nor U10026 (N_10026,N_9607,N_9659);
nor U10027 (N_10027,N_9695,N_9785);
nand U10028 (N_10028,N_9638,N_9700);
nor U10029 (N_10029,N_9660,N_9892);
xnor U10030 (N_10030,N_9800,N_9620);
nand U10031 (N_10031,N_9747,N_9677);
nand U10032 (N_10032,N_9772,N_9799);
or U10033 (N_10033,N_9619,N_9887);
or U10034 (N_10034,N_9625,N_9813);
or U10035 (N_10035,N_9881,N_9773);
and U10036 (N_10036,N_9653,N_9614);
and U10037 (N_10037,N_9822,N_9715);
and U10038 (N_10038,N_9765,N_9824);
nand U10039 (N_10039,N_9825,N_9742);
or U10040 (N_10040,N_9849,N_9882);
nand U10041 (N_10041,N_9624,N_9640);
nor U10042 (N_10042,N_9667,N_9738);
xor U10043 (N_10043,N_9760,N_9678);
xor U10044 (N_10044,N_9806,N_9866);
xnor U10045 (N_10045,N_9668,N_9874);
nor U10046 (N_10046,N_9616,N_9890);
and U10047 (N_10047,N_9850,N_9754);
and U10048 (N_10048,N_9886,N_9636);
nand U10049 (N_10049,N_9702,N_9705);
nand U10050 (N_10050,N_9889,N_9872);
xnor U10051 (N_10051,N_9858,N_9881);
nand U10052 (N_10052,N_9816,N_9646);
xnor U10053 (N_10053,N_9706,N_9648);
nand U10054 (N_10054,N_9764,N_9636);
nor U10055 (N_10055,N_9651,N_9841);
and U10056 (N_10056,N_9788,N_9884);
or U10057 (N_10057,N_9883,N_9715);
nand U10058 (N_10058,N_9773,N_9849);
xnor U10059 (N_10059,N_9674,N_9891);
nand U10060 (N_10060,N_9782,N_9608);
xor U10061 (N_10061,N_9816,N_9884);
nand U10062 (N_10062,N_9609,N_9678);
nor U10063 (N_10063,N_9659,N_9891);
xnor U10064 (N_10064,N_9796,N_9793);
nand U10065 (N_10065,N_9799,N_9840);
xor U10066 (N_10066,N_9633,N_9610);
nand U10067 (N_10067,N_9844,N_9825);
nor U10068 (N_10068,N_9723,N_9820);
or U10069 (N_10069,N_9812,N_9663);
xor U10070 (N_10070,N_9778,N_9750);
and U10071 (N_10071,N_9726,N_9864);
or U10072 (N_10072,N_9657,N_9816);
or U10073 (N_10073,N_9608,N_9678);
xnor U10074 (N_10074,N_9708,N_9664);
and U10075 (N_10075,N_9641,N_9839);
and U10076 (N_10076,N_9627,N_9793);
and U10077 (N_10077,N_9658,N_9653);
or U10078 (N_10078,N_9854,N_9872);
and U10079 (N_10079,N_9849,N_9790);
nand U10080 (N_10080,N_9839,N_9873);
nor U10081 (N_10081,N_9677,N_9899);
xnor U10082 (N_10082,N_9772,N_9656);
nand U10083 (N_10083,N_9685,N_9887);
xnor U10084 (N_10084,N_9812,N_9690);
or U10085 (N_10085,N_9836,N_9891);
and U10086 (N_10086,N_9764,N_9709);
nand U10087 (N_10087,N_9607,N_9828);
xnor U10088 (N_10088,N_9841,N_9856);
or U10089 (N_10089,N_9700,N_9838);
nor U10090 (N_10090,N_9826,N_9605);
or U10091 (N_10091,N_9615,N_9784);
and U10092 (N_10092,N_9753,N_9643);
and U10093 (N_10093,N_9737,N_9872);
and U10094 (N_10094,N_9872,N_9660);
xnor U10095 (N_10095,N_9796,N_9781);
or U10096 (N_10096,N_9755,N_9791);
or U10097 (N_10097,N_9721,N_9787);
and U10098 (N_10098,N_9693,N_9635);
xnor U10099 (N_10099,N_9822,N_9724);
or U10100 (N_10100,N_9861,N_9608);
nand U10101 (N_10101,N_9691,N_9749);
or U10102 (N_10102,N_9691,N_9617);
and U10103 (N_10103,N_9606,N_9697);
and U10104 (N_10104,N_9804,N_9658);
and U10105 (N_10105,N_9612,N_9878);
and U10106 (N_10106,N_9882,N_9863);
nor U10107 (N_10107,N_9626,N_9685);
or U10108 (N_10108,N_9805,N_9613);
nand U10109 (N_10109,N_9805,N_9626);
xnor U10110 (N_10110,N_9842,N_9769);
and U10111 (N_10111,N_9639,N_9673);
xor U10112 (N_10112,N_9659,N_9643);
and U10113 (N_10113,N_9750,N_9803);
or U10114 (N_10114,N_9700,N_9618);
nand U10115 (N_10115,N_9639,N_9770);
nor U10116 (N_10116,N_9741,N_9769);
xnor U10117 (N_10117,N_9612,N_9821);
or U10118 (N_10118,N_9675,N_9830);
nand U10119 (N_10119,N_9687,N_9843);
and U10120 (N_10120,N_9876,N_9815);
nor U10121 (N_10121,N_9618,N_9732);
nand U10122 (N_10122,N_9624,N_9654);
and U10123 (N_10123,N_9676,N_9835);
nor U10124 (N_10124,N_9864,N_9759);
nor U10125 (N_10125,N_9787,N_9826);
and U10126 (N_10126,N_9762,N_9673);
and U10127 (N_10127,N_9895,N_9885);
and U10128 (N_10128,N_9800,N_9663);
or U10129 (N_10129,N_9687,N_9789);
nand U10130 (N_10130,N_9897,N_9683);
nand U10131 (N_10131,N_9728,N_9821);
and U10132 (N_10132,N_9821,N_9631);
and U10133 (N_10133,N_9869,N_9732);
and U10134 (N_10134,N_9753,N_9692);
or U10135 (N_10135,N_9630,N_9826);
nor U10136 (N_10136,N_9635,N_9875);
and U10137 (N_10137,N_9644,N_9838);
and U10138 (N_10138,N_9738,N_9838);
or U10139 (N_10139,N_9761,N_9783);
or U10140 (N_10140,N_9655,N_9681);
xnor U10141 (N_10141,N_9851,N_9771);
xnor U10142 (N_10142,N_9783,N_9676);
nand U10143 (N_10143,N_9804,N_9747);
or U10144 (N_10144,N_9858,N_9711);
nand U10145 (N_10145,N_9834,N_9882);
and U10146 (N_10146,N_9811,N_9646);
xnor U10147 (N_10147,N_9686,N_9664);
xor U10148 (N_10148,N_9740,N_9698);
or U10149 (N_10149,N_9642,N_9725);
or U10150 (N_10150,N_9745,N_9788);
or U10151 (N_10151,N_9727,N_9724);
nor U10152 (N_10152,N_9881,N_9841);
xor U10153 (N_10153,N_9776,N_9687);
nor U10154 (N_10154,N_9699,N_9691);
nand U10155 (N_10155,N_9681,N_9719);
and U10156 (N_10156,N_9723,N_9702);
xor U10157 (N_10157,N_9764,N_9747);
and U10158 (N_10158,N_9691,N_9871);
nand U10159 (N_10159,N_9707,N_9748);
xnor U10160 (N_10160,N_9667,N_9794);
or U10161 (N_10161,N_9782,N_9871);
nand U10162 (N_10162,N_9635,N_9890);
and U10163 (N_10163,N_9655,N_9724);
xor U10164 (N_10164,N_9807,N_9856);
xor U10165 (N_10165,N_9751,N_9768);
nor U10166 (N_10166,N_9870,N_9799);
xor U10167 (N_10167,N_9679,N_9873);
nand U10168 (N_10168,N_9825,N_9870);
nor U10169 (N_10169,N_9677,N_9721);
nand U10170 (N_10170,N_9654,N_9846);
nand U10171 (N_10171,N_9816,N_9877);
nand U10172 (N_10172,N_9742,N_9781);
and U10173 (N_10173,N_9783,N_9728);
and U10174 (N_10174,N_9805,N_9601);
nor U10175 (N_10175,N_9814,N_9720);
nor U10176 (N_10176,N_9782,N_9834);
and U10177 (N_10177,N_9815,N_9678);
and U10178 (N_10178,N_9808,N_9834);
nand U10179 (N_10179,N_9860,N_9604);
nor U10180 (N_10180,N_9630,N_9815);
nand U10181 (N_10181,N_9627,N_9735);
and U10182 (N_10182,N_9648,N_9783);
and U10183 (N_10183,N_9742,N_9880);
nand U10184 (N_10184,N_9843,N_9849);
nor U10185 (N_10185,N_9744,N_9824);
nand U10186 (N_10186,N_9790,N_9782);
nand U10187 (N_10187,N_9693,N_9703);
xor U10188 (N_10188,N_9708,N_9805);
xnor U10189 (N_10189,N_9859,N_9812);
nor U10190 (N_10190,N_9664,N_9771);
or U10191 (N_10191,N_9743,N_9771);
or U10192 (N_10192,N_9702,N_9644);
or U10193 (N_10193,N_9842,N_9823);
nand U10194 (N_10194,N_9807,N_9829);
nand U10195 (N_10195,N_9604,N_9615);
xor U10196 (N_10196,N_9640,N_9891);
nand U10197 (N_10197,N_9641,N_9704);
nor U10198 (N_10198,N_9743,N_9895);
xor U10199 (N_10199,N_9840,N_9655);
or U10200 (N_10200,N_10020,N_10056);
and U10201 (N_10201,N_9936,N_10154);
nor U10202 (N_10202,N_10034,N_10000);
or U10203 (N_10203,N_9940,N_10062);
xor U10204 (N_10204,N_9954,N_10199);
and U10205 (N_10205,N_10148,N_9981);
xor U10206 (N_10206,N_10065,N_10110);
or U10207 (N_10207,N_10181,N_9929);
nand U10208 (N_10208,N_10045,N_9991);
nand U10209 (N_10209,N_10050,N_10145);
nand U10210 (N_10210,N_9977,N_10125);
xnor U10211 (N_10211,N_10035,N_10104);
and U10212 (N_10212,N_9917,N_10012);
or U10213 (N_10213,N_10132,N_10060);
and U10214 (N_10214,N_10066,N_10109);
or U10215 (N_10215,N_10059,N_10180);
xnor U10216 (N_10216,N_10155,N_10025);
xnor U10217 (N_10217,N_9908,N_10043);
or U10218 (N_10218,N_9921,N_9946);
xnor U10219 (N_10219,N_9934,N_9997);
or U10220 (N_10220,N_9972,N_9920);
and U10221 (N_10221,N_9901,N_10079);
or U10222 (N_10222,N_10005,N_9923);
nor U10223 (N_10223,N_10142,N_10166);
nor U10224 (N_10224,N_10040,N_9978);
or U10225 (N_10225,N_10114,N_9957);
and U10226 (N_10226,N_10198,N_10028);
xnor U10227 (N_10227,N_10077,N_10014);
or U10228 (N_10228,N_10058,N_10115);
xor U10229 (N_10229,N_10138,N_10156);
nor U10230 (N_10230,N_10168,N_10108);
and U10231 (N_10231,N_9941,N_9943);
nand U10232 (N_10232,N_10173,N_9995);
nor U10233 (N_10233,N_10096,N_10019);
and U10234 (N_10234,N_10027,N_10193);
or U10235 (N_10235,N_10092,N_10008);
nor U10236 (N_10236,N_10078,N_9969);
nor U10237 (N_10237,N_9994,N_10123);
or U10238 (N_10238,N_9911,N_9950);
and U10239 (N_10239,N_9960,N_10162);
nand U10240 (N_10240,N_10053,N_10068);
or U10241 (N_10241,N_10083,N_9952);
nand U10242 (N_10242,N_10113,N_10188);
xnor U10243 (N_10243,N_10152,N_9973);
nand U10244 (N_10244,N_10021,N_10037);
xor U10245 (N_10245,N_10073,N_9989);
or U10246 (N_10246,N_10135,N_10195);
xnor U10247 (N_10247,N_9986,N_10116);
nand U10248 (N_10248,N_10042,N_10032);
nand U10249 (N_10249,N_9955,N_9964);
or U10250 (N_10250,N_10017,N_10086);
or U10251 (N_10251,N_9919,N_9902);
nor U10252 (N_10252,N_9925,N_9904);
nand U10253 (N_10253,N_10190,N_10146);
nand U10254 (N_10254,N_10127,N_10139);
nand U10255 (N_10255,N_9970,N_10133);
nand U10256 (N_10256,N_9928,N_10192);
nor U10257 (N_10257,N_10074,N_9927);
nand U10258 (N_10258,N_10149,N_10055);
xor U10259 (N_10259,N_10085,N_10186);
xor U10260 (N_10260,N_9967,N_10121);
nand U10261 (N_10261,N_10161,N_10164);
nand U10262 (N_10262,N_10013,N_10070);
and U10263 (N_10263,N_10160,N_10112);
xor U10264 (N_10264,N_10120,N_10006);
or U10265 (N_10265,N_9939,N_10084);
nand U10266 (N_10266,N_10136,N_9987);
or U10267 (N_10267,N_10187,N_10165);
nor U10268 (N_10268,N_10069,N_10071);
xor U10269 (N_10269,N_9942,N_10182);
xnor U10270 (N_10270,N_10080,N_10026);
nand U10271 (N_10271,N_10015,N_10150);
and U10272 (N_10272,N_10038,N_10011);
nor U10273 (N_10273,N_10122,N_10158);
nand U10274 (N_10274,N_9992,N_10126);
nor U10275 (N_10275,N_10140,N_10016);
or U10276 (N_10276,N_10091,N_10049);
nand U10277 (N_10277,N_10039,N_10033);
nand U10278 (N_10278,N_9998,N_9947);
xor U10279 (N_10279,N_10098,N_9971);
xor U10280 (N_10280,N_9938,N_10010);
xor U10281 (N_10281,N_9951,N_10174);
or U10282 (N_10282,N_10047,N_9979);
nor U10283 (N_10283,N_10082,N_9909);
and U10284 (N_10284,N_10089,N_10167);
or U10285 (N_10285,N_9900,N_10087);
xor U10286 (N_10286,N_9974,N_9948);
or U10287 (N_10287,N_10001,N_10044);
or U10288 (N_10288,N_10097,N_10144);
xnor U10289 (N_10289,N_10157,N_10067);
and U10290 (N_10290,N_9912,N_9983);
nand U10291 (N_10291,N_9930,N_9985);
nor U10292 (N_10292,N_10194,N_9906);
or U10293 (N_10293,N_10003,N_10088);
nand U10294 (N_10294,N_9937,N_9988);
nor U10295 (N_10295,N_10093,N_9915);
nor U10296 (N_10296,N_10175,N_10179);
and U10297 (N_10297,N_10197,N_9932);
or U10298 (N_10298,N_9953,N_10170);
or U10299 (N_10299,N_9949,N_10124);
or U10300 (N_10300,N_10018,N_10185);
nor U10301 (N_10301,N_10106,N_9980);
nand U10302 (N_10302,N_9916,N_9914);
or U10303 (N_10303,N_10100,N_9944);
xor U10304 (N_10304,N_10111,N_10009);
nand U10305 (N_10305,N_10141,N_10081);
and U10306 (N_10306,N_9990,N_9903);
or U10307 (N_10307,N_9966,N_10130);
and U10308 (N_10308,N_9962,N_10099);
xor U10309 (N_10309,N_10007,N_9956);
or U10310 (N_10310,N_9945,N_10063);
and U10311 (N_10311,N_10090,N_10029);
xor U10312 (N_10312,N_10134,N_10105);
nand U10313 (N_10313,N_10031,N_10072);
or U10314 (N_10314,N_9907,N_9905);
and U10315 (N_10315,N_10004,N_9982);
xor U10316 (N_10316,N_10041,N_10177);
nor U10317 (N_10317,N_10057,N_9910);
xor U10318 (N_10318,N_10171,N_9993);
and U10319 (N_10319,N_10147,N_10094);
xor U10320 (N_10320,N_10143,N_10051);
nor U10321 (N_10321,N_10076,N_10117);
nand U10322 (N_10322,N_10151,N_10191);
and U10323 (N_10323,N_9958,N_9968);
nor U10324 (N_10324,N_10137,N_9931);
xor U10325 (N_10325,N_10176,N_9918);
or U10326 (N_10326,N_10189,N_10131);
nand U10327 (N_10327,N_9922,N_9984);
or U10328 (N_10328,N_10023,N_10052);
nand U10329 (N_10329,N_9961,N_10183);
nand U10330 (N_10330,N_10054,N_10048);
xor U10331 (N_10331,N_9975,N_9976);
and U10332 (N_10332,N_10118,N_9926);
nand U10333 (N_10333,N_9996,N_9935);
or U10334 (N_10334,N_10046,N_10002);
nor U10335 (N_10335,N_10030,N_10163);
or U10336 (N_10336,N_10128,N_10153);
nand U10337 (N_10337,N_9959,N_10107);
nor U10338 (N_10338,N_9913,N_10022);
or U10339 (N_10339,N_10129,N_10036);
and U10340 (N_10340,N_10102,N_9965);
nand U10341 (N_10341,N_10159,N_10101);
nand U10342 (N_10342,N_10178,N_10064);
nor U10343 (N_10343,N_10061,N_10075);
nor U10344 (N_10344,N_10103,N_9999);
or U10345 (N_10345,N_10119,N_10169);
nor U10346 (N_10346,N_10172,N_9924);
or U10347 (N_10347,N_9933,N_9963);
xor U10348 (N_10348,N_10196,N_10024);
and U10349 (N_10349,N_10184,N_10095);
xnor U10350 (N_10350,N_10180,N_9954);
nor U10351 (N_10351,N_10178,N_9975);
nor U10352 (N_10352,N_10073,N_10092);
nor U10353 (N_10353,N_10007,N_10108);
and U10354 (N_10354,N_10143,N_10025);
nor U10355 (N_10355,N_9946,N_10081);
or U10356 (N_10356,N_9912,N_10014);
xnor U10357 (N_10357,N_10024,N_10195);
or U10358 (N_10358,N_9921,N_9995);
or U10359 (N_10359,N_10170,N_10011);
xor U10360 (N_10360,N_9917,N_10126);
and U10361 (N_10361,N_9992,N_9951);
xnor U10362 (N_10362,N_9959,N_10126);
xnor U10363 (N_10363,N_10090,N_10111);
nand U10364 (N_10364,N_10012,N_10077);
nor U10365 (N_10365,N_10034,N_9933);
xnor U10366 (N_10366,N_9980,N_9978);
nor U10367 (N_10367,N_10083,N_10153);
xnor U10368 (N_10368,N_10115,N_10114);
nor U10369 (N_10369,N_10099,N_10193);
nand U10370 (N_10370,N_10088,N_10046);
and U10371 (N_10371,N_10118,N_10184);
and U10372 (N_10372,N_9904,N_9976);
xor U10373 (N_10373,N_9927,N_10132);
and U10374 (N_10374,N_10011,N_9923);
xor U10375 (N_10375,N_10093,N_10124);
xor U10376 (N_10376,N_9983,N_9903);
xor U10377 (N_10377,N_9925,N_9939);
xnor U10378 (N_10378,N_10140,N_10093);
and U10379 (N_10379,N_10080,N_9982);
or U10380 (N_10380,N_10038,N_10125);
or U10381 (N_10381,N_10159,N_10110);
nand U10382 (N_10382,N_9918,N_10136);
or U10383 (N_10383,N_10115,N_10045);
nand U10384 (N_10384,N_9940,N_10182);
nor U10385 (N_10385,N_10110,N_10000);
nor U10386 (N_10386,N_9907,N_9909);
and U10387 (N_10387,N_10085,N_10185);
nand U10388 (N_10388,N_10118,N_10068);
nand U10389 (N_10389,N_10142,N_10089);
nor U10390 (N_10390,N_9997,N_10074);
or U10391 (N_10391,N_10044,N_9984);
and U10392 (N_10392,N_9906,N_9945);
and U10393 (N_10393,N_10195,N_10046);
or U10394 (N_10394,N_10187,N_10185);
or U10395 (N_10395,N_9925,N_10178);
and U10396 (N_10396,N_9908,N_9931);
nand U10397 (N_10397,N_9950,N_10182);
or U10398 (N_10398,N_9906,N_10149);
or U10399 (N_10399,N_10163,N_9978);
nand U10400 (N_10400,N_10157,N_10052);
or U10401 (N_10401,N_9910,N_10025);
and U10402 (N_10402,N_10073,N_10017);
and U10403 (N_10403,N_9939,N_10159);
or U10404 (N_10404,N_10042,N_10162);
nor U10405 (N_10405,N_10164,N_10035);
and U10406 (N_10406,N_9948,N_10035);
or U10407 (N_10407,N_10064,N_10189);
nand U10408 (N_10408,N_10193,N_9945);
nand U10409 (N_10409,N_9990,N_9963);
and U10410 (N_10410,N_10032,N_10124);
and U10411 (N_10411,N_10078,N_9947);
and U10412 (N_10412,N_10087,N_9966);
and U10413 (N_10413,N_10045,N_10018);
nand U10414 (N_10414,N_10167,N_10119);
nor U10415 (N_10415,N_10117,N_10090);
or U10416 (N_10416,N_9905,N_10033);
or U10417 (N_10417,N_9999,N_10194);
and U10418 (N_10418,N_10055,N_9919);
xnor U10419 (N_10419,N_10131,N_10071);
or U10420 (N_10420,N_10021,N_10189);
and U10421 (N_10421,N_10064,N_10147);
xor U10422 (N_10422,N_10113,N_10102);
nand U10423 (N_10423,N_10104,N_10170);
and U10424 (N_10424,N_10197,N_10054);
and U10425 (N_10425,N_10010,N_10144);
nor U10426 (N_10426,N_9953,N_9937);
and U10427 (N_10427,N_9960,N_10070);
nor U10428 (N_10428,N_10120,N_10155);
xnor U10429 (N_10429,N_10175,N_10100);
or U10430 (N_10430,N_9996,N_9959);
and U10431 (N_10431,N_10023,N_10028);
and U10432 (N_10432,N_9930,N_9911);
nand U10433 (N_10433,N_10119,N_10106);
or U10434 (N_10434,N_10139,N_10152);
nor U10435 (N_10435,N_9910,N_9983);
xnor U10436 (N_10436,N_9993,N_9992);
nand U10437 (N_10437,N_9940,N_10194);
xnor U10438 (N_10438,N_10164,N_9922);
and U10439 (N_10439,N_10136,N_10058);
xnor U10440 (N_10440,N_10117,N_9941);
and U10441 (N_10441,N_10079,N_10098);
nor U10442 (N_10442,N_10173,N_9924);
or U10443 (N_10443,N_10196,N_9943);
xnor U10444 (N_10444,N_10089,N_10110);
or U10445 (N_10445,N_10084,N_9977);
nor U10446 (N_10446,N_9952,N_10170);
nor U10447 (N_10447,N_10173,N_10014);
or U10448 (N_10448,N_9996,N_10092);
and U10449 (N_10449,N_10027,N_10100);
xor U10450 (N_10450,N_10165,N_10170);
nand U10451 (N_10451,N_10190,N_9999);
xnor U10452 (N_10452,N_10155,N_10154);
nor U10453 (N_10453,N_9978,N_10125);
nand U10454 (N_10454,N_9984,N_9940);
xor U10455 (N_10455,N_10070,N_9918);
nand U10456 (N_10456,N_9901,N_9988);
nand U10457 (N_10457,N_10021,N_9948);
nor U10458 (N_10458,N_10118,N_9979);
nand U10459 (N_10459,N_10065,N_10004);
nor U10460 (N_10460,N_10015,N_10036);
or U10461 (N_10461,N_10013,N_10000);
xnor U10462 (N_10462,N_9993,N_10155);
nand U10463 (N_10463,N_10060,N_9966);
or U10464 (N_10464,N_10066,N_10103);
xor U10465 (N_10465,N_10074,N_9910);
and U10466 (N_10466,N_10108,N_9941);
nor U10467 (N_10467,N_10034,N_9968);
nor U10468 (N_10468,N_10039,N_10073);
xnor U10469 (N_10469,N_10096,N_10067);
nand U10470 (N_10470,N_10121,N_10160);
or U10471 (N_10471,N_10175,N_10177);
nor U10472 (N_10472,N_10191,N_9983);
nand U10473 (N_10473,N_10082,N_10159);
nor U10474 (N_10474,N_9963,N_10192);
xnor U10475 (N_10475,N_10130,N_9958);
xnor U10476 (N_10476,N_10095,N_9967);
xnor U10477 (N_10477,N_10051,N_9950);
or U10478 (N_10478,N_9960,N_10106);
nor U10479 (N_10479,N_9908,N_9994);
nor U10480 (N_10480,N_9927,N_9971);
nand U10481 (N_10481,N_10177,N_10012);
or U10482 (N_10482,N_10006,N_10118);
and U10483 (N_10483,N_9943,N_10199);
nand U10484 (N_10484,N_9904,N_10173);
nand U10485 (N_10485,N_10160,N_10167);
nand U10486 (N_10486,N_9959,N_10173);
nand U10487 (N_10487,N_10031,N_10016);
or U10488 (N_10488,N_10024,N_10125);
or U10489 (N_10489,N_10128,N_9961);
and U10490 (N_10490,N_9985,N_10074);
or U10491 (N_10491,N_9954,N_9983);
xor U10492 (N_10492,N_9933,N_10096);
nor U10493 (N_10493,N_9932,N_10117);
xnor U10494 (N_10494,N_10097,N_10189);
nor U10495 (N_10495,N_9926,N_10014);
or U10496 (N_10496,N_10032,N_10096);
nand U10497 (N_10497,N_10072,N_9918);
or U10498 (N_10498,N_9962,N_9946);
nand U10499 (N_10499,N_9908,N_9911);
nand U10500 (N_10500,N_10480,N_10290);
nor U10501 (N_10501,N_10367,N_10481);
and U10502 (N_10502,N_10311,N_10214);
or U10503 (N_10503,N_10417,N_10438);
nand U10504 (N_10504,N_10499,N_10372);
xnor U10505 (N_10505,N_10272,N_10223);
xor U10506 (N_10506,N_10465,N_10406);
nor U10507 (N_10507,N_10256,N_10228);
nand U10508 (N_10508,N_10255,N_10405);
xor U10509 (N_10509,N_10334,N_10307);
xnor U10510 (N_10510,N_10262,N_10246);
nor U10511 (N_10511,N_10289,N_10497);
nor U10512 (N_10512,N_10387,N_10490);
xor U10513 (N_10513,N_10475,N_10401);
nor U10514 (N_10514,N_10350,N_10291);
and U10515 (N_10515,N_10200,N_10202);
nor U10516 (N_10516,N_10376,N_10313);
xnor U10517 (N_10517,N_10331,N_10349);
xor U10518 (N_10518,N_10282,N_10201);
xnor U10519 (N_10519,N_10474,N_10213);
and U10520 (N_10520,N_10306,N_10479);
xnor U10521 (N_10521,N_10339,N_10495);
xnor U10522 (N_10522,N_10207,N_10205);
nand U10523 (N_10523,N_10469,N_10287);
or U10524 (N_10524,N_10276,N_10275);
xor U10525 (N_10525,N_10408,N_10280);
or U10526 (N_10526,N_10298,N_10463);
nor U10527 (N_10527,N_10379,N_10393);
or U10528 (N_10528,N_10448,N_10324);
xnor U10529 (N_10529,N_10317,N_10428);
nor U10530 (N_10530,N_10208,N_10435);
or U10531 (N_10531,N_10380,N_10454);
or U10532 (N_10532,N_10297,N_10375);
nand U10533 (N_10533,N_10348,N_10314);
and U10534 (N_10534,N_10388,N_10278);
or U10535 (N_10535,N_10437,N_10399);
xor U10536 (N_10536,N_10310,N_10390);
xor U10537 (N_10537,N_10312,N_10343);
nor U10538 (N_10538,N_10274,N_10277);
nor U10539 (N_10539,N_10233,N_10316);
nand U10540 (N_10540,N_10257,N_10263);
nor U10541 (N_10541,N_10320,N_10398);
and U10542 (N_10542,N_10327,N_10484);
xor U10543 (N_10543,N_10241,N_10421);
nand U10544 (N_10544,N_10204,N_10493);
nor U10545 (N_10545,N_10452,N_10416);
and U10546 (N_10546,N_10209,N_10411);
nand U10547 (N_10547,N_10221,N_10333);
nand U10548 (N_10548,N_10305,N_10423);
nor U10549 (N_10549,N_10235,N_10472);
nand U10550 (N_10550,N_10212,N_10366);
or U10551 (N_10551,N_10344,N_10336);
and U10552 (N_10552,N_10301,N_10419);
and U10553 (N_10553,N_10422,N_10457);
and U10554 (N_10554,N_10361,N_10449);
xor U10555 (N_10555,N_10477,N_10337);
or U10556 (N_10556,N_10247,N_10227);
nand U10557 (N_10557,N_10450,N_10385);
xor U10558 (N_10558,N_10459,N_10273);
or U10559 (N_10559,N_10325,N_10412);
nand U10560 (N_10560,N_10299,N_10381);
xor U10561 (N_10561,N_10303,N_10468);
nor U10562 (N_10562,N_10357,N_10363);
and U10563 (N_10563,N_10391,N_10210);
or U10564 (N_10564,N_10295,N_10249);
xnor U10565 (N_10565,N_10486,N_10446);
xnor U10566 (N_10566,N_10460,N_10378);
or U10567 (N_10567,N_10230,N_10487);
xnor U10568 (N_10568,N_10395,N_10237);
nor U10569 (N_10569,N_10365,N_10341);
nor U10570 (N_10570,N_10242,N_10476);
nand U10571 (N_10571,N_10383,N_10461);
nand U10572 (N_10572,N_10220,N_10252);
and U10573 (N_10573,N_10342,N_10354);
and U10574 (N_10574,N_10266,N_10473);
nor U10575 (N_10575,N_10425,N_10482);
xnor U10576 (N_10576,N_10329,N_10283);
nor U10577 (N_10577,N_10347,N_10321);
and U10578 (N_10578,N_10386,N_10315);
nor U10579 (N_10579,N_10360,N_10330);
nand U10580 (N_10580,N_10444,N_10478);
xnor U10581 (N_10581,N_10418,N_10264);
nor U10582 (N_10582,N_10281,N_10420);
or U10583 (N_10583,N_10351,N_10394);
nand U10584 (N_10584,N_10489,N_10218);
nor U10585 (N_10585,N_10245,N_10356);
and U10586 (N_10586,N_10466,N_10397);
nor U10587 (N_10587,N_10483,N_10359);
and U10588 (N_10588,N_10234,N_10413);
or U10589 (N_10589,N_10429,N_10492);
xnor U10590 (N_10590,N_10326,N_10410);
and U10591 (N_10591,N_10253,N_10471);
and U10592 (N_10592,N_10293,N_10240);
or U10593 (N_10593,N_10323,N_10370);
xor U10594 (N_10594,N_10396,N_10358);
nand U10595 (N_10595,N_10424,N_10494);
nand U10596 (N_10596,N_10254,N_10271);
xor U10597 (N_10597,N_10203,N_10355);
or U10598 (N_10598,N_10368,N_10216);
or U10599 (N_10599,N_10407,N_10447);
or U10600 (N_10600,N_10261,N_10338);
or U10601 (N_10601,N_10384,N_10467);
nand U10602 (N_10602,N_10427,N_10340);
xnor U10603 (N_10603,N_10335,N_10488);
nor U10604 (N_10604,N_10439,N_10222);
and U10605 (N_10605,N_10403,N_10258);
nor U10606 (N_10606,N_10269,N_10371);
and U10607 (N_10607,N_10345,N_10302);
nand U10608 (N_10608,N_10485,N_10445);
and U10609 (N_10609,N_10250,N_10309);
xor U10610 (N_10610,N_10491,N_10267);
nor U10611 (N_10611,N_10456,N_10279);
or U10612 (N_10612,N_10415,N_10464);
or U10613 (N_10613,N_10362,N_10294);
or U10614 (N_10614,N_10318,N_10239);
or U10615 (N_10615,N_10248,N_10286);
and U10616 (N_10616,N_10409,N_10453);
nor U10617 (N_10617,N_10440,N_10231);
or U10618 (N_10618,N_10451,N_10364);
or U10619 (N_10619,N_10458,N_10243);
nand U10620 (N_10620,N_10260,N_10400);
xnor U10621 (N_10621,N_10265,N_10224);
nor U10622 (N_10622,N_10462,N_10498);
xnor U10623 (N_10623,N_10211,N_10285);
and U10624 (N_10624,N_10431,N_10288);
or U10625 (N_10625,N_10300,N_10319);
or U10626 (N_10626,N_10251,N_10496);
xor U10627 (N_10627,N_10268,N_10328);
or U10628 (N_10628,N_10292,N_10215);
or U10629 (N_10629,N_10470,N_10382);
nand U10630 (N_10630,N_10284,N_10225);
or U10631 (N_10631,N_10352,N_10244);
nor U10632 (N_10632,N_10322,N_10402);
or U10633 (N_10633,N_10434,N_10346);
nand U10634 (N_10634,N_10374,N_10373);
or U10635 (N_10635,N_10353,N_10226);
nor U10636 (N_10636,N_10442,N_10219);
nor U10637 (N_10637,N_10414,N_10430);
and U10638 (N_10638,N_10270,N_10377);
or U10639 (N_10639,N_10332,N_10206);
xor U10640 (N_10640,N_10229,N_10217);
and U10641 (N_10641,N_10432,N_10296);
nand U10642 (N_10642,N_10238,N_10308);
or U10643 (N_10643,N_10259,N_10392);
nor U10644 (N_10644,N_10441,N_10433);
or U10645 (N_10645,N_10455,N_10369);
nand U10646 (N_10646,N_10389,N_10436);
nor U10647 (N_10647,N_10404,N_10443);
and U10648 (N_10648,N_10236,N_10304);
and U10649 (N_10649,N_10232,N_10426);
xor U10650 (N_10650,N_10405,N_10296);
xnor U10651 (N_10651,N_10470,N_10293);
nor U10652 (N_10652,N_10373,N_10230);
nand U10653 (N_10653,N_10365,N_10333);
nor U10654 (N_10654,N_10277,N_10219);
nor U10655 (N_10655,N_10307,N_10367);
nor U10656 (N_10656,N_10315,N_10442);
nand U10657 (N_10657,N_10397,N_10417);
nand U10658 (N_10658,N_10370,N_10264);
xnor U10659 (N_10659,N_10454,N_10460);
or U10660 (N_10660,N_10496,N_10405);
or U10661 (N_10661,N_10371,N_10344);
or U10662 (N_10662,N_10300,N_10492);
or U10663 (N_10663,N_10248,N_10225);
and U10664 (N_10664,N_10357,N_10440);
or U10665 (N_10665,N_10341,N_10398);
nor U10666 (N_10666,N_10417,N_10323);
nor U10667 (N_10667,N_10236,N_10328);
nor U10668 (N_10668,N_10462,N_10228);
xor U10669 (N_10669,N_10246,N_10422);
nand U10670 (N_10670,N_10335,N_10317);
xor U10671 (N_10671,N_10419,N_10240);
nand U10672 (N_10672,N_10372,N_10273);
and U10673 (N_10673,N_10219,N_10304);
nand U10674 (N_10674,N_10494,N_10236);
nand U10675 (N_10675,N_10317,N_10295);
nand U10676 (N_10676,N_10341,N_10221);
and U10677 (N_10677,N_10213,N_10478);
or U10678 (N_10678,N_10497,N_10212);
nand U10679 (N_10679,N_10233,N_10384);
or U10680 (N_10680,N_10482,N_10424);
or U10681 (N_10681,N_10416,N_10342);
nand U10682 (N_10682,N_10212,N_10268);
nor U10683 (N_10683,N_10223,N_10239);
nand U10684 (N_10684,N_10270,N_10240);
xnor U10685 (N_10685,N_10482,N_10337);
xnor U10686 (N_10686,N_10219,N_10307);
nor U10687 (N_10687,N_10231,N_10291);
xnor U10688 (N_10688,N_10441,N_10218);
xor U10689 (N_10689,N_10244,N_10212);
nand U10690 (N_10690,N_10339,N_10441);
xor U10691 (N_10691,N_10313,N_10243);
xnor U10692 (N_10692,N_10203,N_10356);
xnor U10693 (N_10693,N_10334,N_10257);
and U10694 (N_10694,N_10447,N_10301);
xor U10695 (N_10695,N_10245,N_10289);
nor U10696 (N_10696,N_10411,N_10300);
xnor U10697 (N_10697,N_10335,N_10227);
nand U10698 (N_10698,N_10429,N_10366);
and U10699 (N_10699,N_10346,N_10344);
nor U10700 (N_10700,N_10390,N_10386);
xor U10701 (N_10701,N_10429,N_10457);
nand U10702 (N_10702,N_10213,N_10383);
and U10703 (N_10703,N_10440,N_10460);
xnor U10704 (N_10704,N_10490,N_10408);
xnor U10705 (N_10705,N_10497,N_10209);
nor U10706 (N_10706,N_10362,N_10336);
and U10707 (N_10707,N_10428,N_10237);
nand U10708 (N_10708,N_10434,N_10339);
xnor U10709 (N_10709,N_10330,N_10224);
xnor U10710 (N_10710,N_10277,N_10499);
xnor U10711 (N_10711,N_10285,N_10416);
nand U10712 (N_10712,N_10480,N_10280);
and U10713 (N_10713,N_10203,N_10373);
nand U10714 (N_10714,N_10203,N_10244);
xnor U10715 (N_10715,N_10448,N_10447);
and U10716 (N_10716,N_10458,N_10479);
and U10717 (N_10717,N_10452,N_10287);
or U10718 (N_10718,N_10289,N_10418);
or U10719 (N_10719,N_10299,N_10438);
or U10720 (N_10720,N_10435,N_10310);
nor U10721 (N_10721,N_10498,N_10229);
nand U10722 (N_10722,N_10270,N_10207);
or U10723 (N_10723,N_10332,N_10429);
nor U10724 (N_10724,N_10320,N_10384);
xnor U10725 (N_10725,N_10305,N_10486);
xnor U10726 (N_10726,N_10312,N_10307);
and U10727 (N_10727,N_10494,N_10232);
and U10728 (N_10728,N_10436,N_10319);
or U10729 (N_10729,N_10232,N_10470);
and U10730 (N_10730,N_10414,N_10440);
or U10731 (N_10731,N_10225,N_10292);
nand U10732 (N_10732,N_10489,N_10210);
or U10733 (N_10733,N_10262,N_10264);
nand U10734 (N_10734,N_10334,N_10339);
and U10735 (N_10735,N_10394,N_10377);
nand U10736 (N_10736,N_10335,N_10449);
nor U10737 (N_10737,N_10496,N_10330);
xnor U10738 (N_10738,N_10459,N_10409);
nor U10739 (N_10739,N_10274,N_10385);
or U10740 (N_10740,N_10231,N_10260);
nand U10741 (N_10741,N_10363,N_10371);
nand U10742 (N_10742,N_10272,N_10496);
or U10743 (N_10743,N_10404,N_10276);
and U10744 (N_10744,N_10438,N_10490);
and U10745 (N_10745,N_10397,N_10298);
and U10746 (N_10746,N_10493,N_10260);
xor U10747 (N_10747,N_10380,N_10427);
nor U10748 (N_10748,N_10328,N_10298);
nand U10749 (N_10749,N_10349,N_10354);
or U10750 (N_10750,N_10401,N_10316);
and U10751 (N_10751,N_10209,N_10341);
or U10752 (N_10752,N_10233,N_10209);
nor U10753 (N_10753,N_10418,N_10335);
nand U10754 (N_10754,N_10353,N_10368);
and U10755 (N_10755,N_10203,N_10460);
and U10756 (N_10756,N_10291,N_10445);
or U10757 (N_10757,N_10313,N_10442);
or U10758 (N_10758,N_10355,N_10427);
nor U10759 (N_10759,N_10352,N_10441);
nor U10760 (N_10760,N_10223,N_10313);
and U10761 (N_10761,N_10319,N_10285);
nor U10762 (N_10762,N_10387,N_10324);
nor U10763 (N_10763,N_10395,N_10346);
or U10764 (N_10764,N_10482,N_10306);
or U10765 (N_10765,N_10327,N_10295);
xnor U10766 (N_10766,N_10299,N_10369);
nor U10767 (N_10767,N_10308,N_10266);
nand U10768 (N_10768,N_10217,N_10280);
and U10769 (N_10769,N_10274,N_10405);
nor U10770 (N_10770,N_10486,N_10338);
xor U10771 (N_10771,N_10264,N_10491);
and U10772 (N_10772,N_10201,N_10270);
nor U10773 (N_10773,N_10468,N_10320);
xor U10774 (N_10774,N_10365,N_10447);
and U10775 (N_10775,N_10357,N_10348);
nand U10776 (N_10776,N_10244,N_10267);
xor U10777 (N_10777,N_10478,N_10288);
nor U10778 (N_10778,N_10360,N_10413);
xor U10779 (N_10779,N_10345,N_10376);
and U10780 (N_10780,N_10371,N_10284);
xnor U10781 (N_10781,N_10358,N_10488);
nand U10782 (N_10782,N_10306,N_10263);
nor U10783 (N_10783,N_10438,N_10341);
nor U10784 (N_10784,N_10396,N_10230);
or U10785 (N_10785,N_10456,N_10423);
or U10786 (N_10786,N_10320,N_10474);
nand U10787 (N_10787,N_10236,N_10489);
xnor U10788 (N_10788,N_10322,N_10215);
nor U10789 (N_10789,N_10268,N_10487);
xor U10790 (N_10790,N_10409,N_10480);
and U10791 (N_10791,N_10352,N_10469);
or U10792 (N_10792,N_10452,N_10278);
nand U10793 (N_10793,N_10406,N_10415);
or U10794 (N_10794,N_10407,N_10451);
nor U10795 (N_10795,N_10332,N_10224);
and U10796 (N_10796,N_10246,N_10251);
and U10797 (N_10797,N_10330,N_10373);
nand U10798 (N_10798,N_10489,N_10386);
nand U10799 (N_10799,N_10263,N_10278);
or U10800 (N_10800,N_10666,N_10611);
nand U10801 (N_10801,N_10546,N_10702);
or U10802 (N_10802,N_10650,N_10533);
nand U10803 (N_10803,N_10500,N_10784);
nor U10804 (N_10804,N_10585,N_10715);
and U10805 (N_10805,N_10581,N_10723);
xnor U10806 (N_10806,N_10530,N_10799);
and U10807 (N_10807,N_10783,N_10521);
or U10808 (N_10808,N_10518,N_10719);
or U10809 (N_10809,N_10580,N_10712);
or U10810 (N_10810,N_10596,N_10682);
nand U10811 (N_10811,N_10553,N_10535);
xor U10812 (N_10812,N_10538,N_10543);
nor U10813 (N_10813,N_10558,N_10711);
xor U10814 (N_10814,N_10753,N_10695);
or U10815 (N_10815,N_10793,N_10794);
and U10816 (N_10816,N_10792,N_10778);
or U10817 (N_10817,N_10674,N_10577);
or U10818 (N_10818,N_10601,N_10566);
xnor U10819 (N_10819,N_10503,N_10625);
nand U10820 (N_10820,N_10663,N_10759);
xnor U10821 (N_10821,N_10645,N_10796);
and U10822 (N_10822,N_10504,N_10727);
or U10823 (N_10823,N_10705,N_10642);
xnor U10824 (N_10824,N_10547,N_10773);
nand U10825 (N_10825,N_10579,N_10678);
and U10826 (N_10826,N_10676,N_10647);
and U10827 (N_10827,N_10505,N_10629);
nand U10828 (N_10828,N_10698,N_10770);
and U10829 (N_10829,N_10785,N_10714);
and U10830 (N_10830,N_10507,N_10600);
nor U10831 (N_10831,N_10692,N_10709);
nor U10832 (N_10832,N_10680,N_10704);
and U10833 (N_10833,N_10584,N_10755);
nor U10834 (N_10834,N_10631,N_10758);
and U10835 (N_10835,N_10540,N_10743);
and U10836 (N_10836,N_10578,N_10545);
and U10837 (N_10837,N_10575,N_10693);
nor U10838 (N_10838,N_10549,N_10517);
nand U10839 (N_10839,N_10737,N_10722);
or U10840 (N_10840,N_10605,N_10526);
nor U10841 (N_10841,N_10774,N_10637);
or U10842 (N_10842,N_10655,N_10564);
nor U10843 (N_10843,N_10668,N_10527);
xnor U10844 (N_10844,N_10679,N_10516);
nor U10845 (N_10845,N_10544,N_10552);
or U10846 (N_10846,N_10539,N_10536);
nor U10847 (N_10847,N_10617,N_10738);
or U10848 (N_10848,N_10542,N_10616);
nor U10849 (N_10849,N_10664,N_10673);
xor U10850 (N_10850,N_10761,N_10772);
nor U10851 (N_10851,N_10532,N_10561);
and U10852 (N_10852,N_10634,N_10626);
and U10853 (N_10853,N_10652,N_10582);
nor U10854 (N_10854,N_10555,N_10734);
nor U10855 (N_10855,N_10649,N_10602);
or U10856 (N_10856,N_10775,N_10613);
xor U10857 (N_10857,N_10730,N_10754);
xor U10858 (N_10858,N_10548,N_10610);
or U10859 (N_10859,N_10741,N_10639);
xnor U10860 (N_10860,N_10591,N_10609);
and U10861 (N_10861,N_10568,N_10752);
or U10862 (N_10862,N_10615,N_10573);
xor U10863 (N_10863,N_10751,N_10798);
and U10864 (N_10864,N_10716,N_10620);
and U10865 (N_10865,N_10725,N_10740);
and U10866 (N_10866,N_10586,N_10748);
nor U10867 (N_10867,N_10628,N_10736);
nor U10868 (N_10868,N_10764,N_10660);
and U10869 (N_10869,N_10677,N_10641);
nand U10870 (N_10870,N_10635,N_10572);
or U10871 (N_10871,N_10757,N_10681);
nor U10872 (N_10872,N_10721,N_10720);
nor U10873 (N_10873,N_10576,N_10694);
nor U10874 (N_10874,N_10782,N_10750);
or U10875 (N_10875,N_10509,N_10728);
xor U10876 (N_10876,N_10656,N_10658);
or U10877 (N_10877,N_10537,N_10502);
and U10878 (N_10878,N_10787,N_10648);
xnor U10879 (N_10879,N_10523,N_10588);
xor U10880 (N_10880,N_10618,N_10747);
and U10881 (N_10881,N_10671,N_10607);
nor U10882 (N_10882,N_10510,N_10632);
and U10883 (N_10883,N_10706,N_10501);
nor U10884 (N_10884,N_10640,N_10779);
xor U10885 (N_10885,N_10563,N_10684);
nand U10886 (N_10886,N_10797,N_10571);
xnor U10887 (N_10887,N_10767,N_10554);
xor U10888 (N_10888,N_10651,N_10606);
nor U10889 (N_10889,N_10657,N_10519);
nor U10890 (N_10890,N_10732,N_10745);
xor U10891 (N_10891,N_10569,N_10556);
xnor U10892 (N_10892,N_10780,N_10735);
xor U10893 (N_10893,N_10522,N_10691);
or U10894 (N_10894,N_10623,N_10590);
nand U10895 (N_10895,N_10619,N_10622);
or U10896 (N_10896,N_10756,N_10534);
nor U10897 (N_10897,N_10643,N_10739);
or U10898 (N_10898,N_10688,N_10703);
nor U10899 (N_10899,N_10627,N_10795);
nor U10900 (N_10900,N_10675,N_10560);
and U10901 (N_10901,N_10524,N_10541);
nor U10902 (N_10902,N_10708,N_10724);
nand U10903 (N_10903,N_10570,N_10512);
xnor U10904 (N_10904,N_10696,N_10514);
nand U10905 (N_10905,N_10608,N_10713);
and U10906 (N_10906,N_10768,N_10686);
and U10907 (N_10907,N_10670,N_10742);
xor U10908 (N_10908,N_10525,N_10598);
xnor U10909 (N_10909,N_10515,N_10528);
nor U10910 (N_10910,N_10726,N_10665);
xor U10911 (N_10911,N_10599,N_10733);
and U10912 (N_10912,N_10672,N_10621);
and U10913 (N_10913,N_10789,N_10595);
and U10914 (N_10914,N_10667,N_10746);
or U10915 (N_10915,N_10624,N_10683);
nor U10916 (N_10916,N_10653,N_10687);
nand U10917 (N_10917,N_10531,N_10644);
nor U10918 (N_10918,N_10565,N_10559);
and U10919 (N_10919,N_10593,N_10700);
and U10920 (N_10920,N_10669,N_10506);
or U10921 (N_10921,N_10636,N_10562);
and U10922 (N_10922,N_10788,N_10612);
or U10923 (N_10923,N_10760,N_10699);
nand U10924 (N_10924,N_10731,N_10587);
nand U10925 (N_10925,N_10614,N_10765);
or U10926 (N_10926,N_10520,N_10769);
nor U10927 (N_10927,N_10701,N_10685);
nor U10928 (N_10928,N_10654,N_10529);
or U10929 (N_10929,N_10781,N_10790);
nor U10930 (N_10930,N_10710,N_10646);
nand U10931 (N_10931,N_10592,N_10557);
and U10932 (N_10932,N_10638,N_10513);
and U10933 (N_10933,N_10574,N_10567);
or U10934 (N_10934,N_10762,N_10771);
or U10935 (N_10935,N_10744,N_10763);
and U10936 (N_10936,N_10508,N_10583);
or U10937 (N_10937,N_10786,N_10729);
or U10938 (N_10938,N_10550,N_10630);
and U10939 (N_10939,N_10662,N_10659);
nand U10940 (N_10940,N_10589,N_10690);
nand U10941 (N_10941,N_10749,N_10603);
or U10942 (N_10942,N_10511,N_10717);
nor U10943 (N_10943,N_10689,N_10791);
or U10944 (N_10944,N_10777,N_10551);
nand U10945 (N_10945,N_10776,N_10661);
xnor U10946 (N_10946,N_10766,N_10697);
and U10947 (N_10947,N_10633,N_10604);
nand U10948 (N_10948,N_10707,N_10597);
and U10949 (N_10949,N_10594,N_10718);
or U10950 (N_10950,N_10552,N_10638);
nand U10951 (N_10951,N_10681,N_10765);
nor U10952 (N_10952,N_10676,N_10609);
nor U10953 (N_10953,N_10734,N_10693);
xor U10954 (N_10954,N_10773,N_10592);
or U10955 (N_10955,N_10617,N_10609);
nor U10956 (N_10956,N_10729,N_10747);
nand U10957 (N_10957,N_10522,N_10629);
or U10958 (N_10958,N_10579,N_10576);
nand U10959 (N_10959,N_10577,N_10646);
xnor U10960 (N_10960,N_10632,N_10595);
or U10961 (N_10961,N_10575,N_10514);
and U10962 (N_10962,N_10586,N_10559);
xor U10963 (N_10963,N_10599,N_10682);
or U10964 (N_10964,N_10633,N_10661);
nor U10965 (N_10965,N_10554,N_10646);
nand U10966 (N_10966,N_10549,N_10673);
nor U10967 (N_10967,N_10781,N_10603);
or U10968 (N_10968,N_10782,N_10575);
xor U10969 (N_10969,N_10673,N_10525);
nand U10970 (N_10970,N_10696,N_10526);
nand U10971 (N_10971,N_10633,N_10589);
xnor U10972 (N_10972,N_10607,N_10735);
and U10973 (N_10973,N_10503,N_10670);
or U10974 (N_10974,N_10587,N_10774);
nand U10975 (N_10975,N_10746,N_10703);
xor U10976 (N_10976,N_10504,N_10639);
nand U10977 (N_10977,N_10733,N_10783);
and U10978 (N_10978,N_10546,N_10598);
nor U10979 (N_10979,N_10584,N_10799);
or U10980 (N_10980,N_10574,N_10532);
xor U10981 (N_10981,N_10538,N_10714);
or U10982 (N_10982,N_10541,N_10741);
nand U10983 (N_10983,N_10783,N_10563);
nor U10984 (N_10984,N_10646,N_10757);
and U10985 (N_10985,N_10671,N_10646);
or U10986 (N_10986,N_10533,N_10768);
nor U10987 (N_10987,N_10638,N_10700);
or U10988 (N_10988,N_10704,N_10643);
nor U10989 (N_10989,N_10576,N_10667);
nor U10990 (N_10990,N_10615,N_10766);
nand U10991 (N_10991,N_10776,N_10783);
and U10992 (N_10992,N_10710,N_10759);
nand U10993 (N_10993,N_10666,N_10769);
or U10994 (N_10994,N_10748,N_10773);
nand U10995 (N_10995,N_10784,N_10753);
xnor U10996 (N_10996,N_10604,N_10532);
nor U10997 (N_10997,N_10699,N_10503);
nand U10998 (N_10998,N_10595,N_10673);
or U10999 (N_10999,N_10780,N_10784);
nor U11000 (N_11000,N_10605,N_10601);
nor U11001 (N_11001,N_10577,N_10555);
nand U11002 (N_11002,N_10641,N_10554);
nand U11003 (N_11003,N_10662,N_10670);
nand U11004 (N_11004,N_10799,N_10784);
or U11005 (N_11005,N_10747,N_10676);
or U11006 (N_11006,N_10697,N_10693);
nor U11007 (N_11007,N_10684,N_10570);
nor U11008 (N_11008,N_10741,N_10798);
nand U11009 (N_11009,N_10767,N_10680);
xnor U11010 (N_11010,N_10599,N_10797);
nor U11011 (N_11011,N_10763,N_10553);
and U11012 (N_11012,N_10638,N_10782);
nand U11013 (N_11013,N_10772,N_10645);
and U11014 (N_11014,N_10679,N_10707);
nor U11015 (N_11015,N_10572,N_10634);
and U11016 (N_11016,N_10522,N_10749);
or U11017 (N_11017,N_10759,N_10575);
nor U11018 (N_11018,N_10795,N_10591);
and U11019 (N_11019,N_10546,N_10712);
xnor U11020 (N_11020,N_10507,N_10658);
and U11021 (N_11021,N_10527,N_10685);
nor U11022 (N_11022,N_10651,N_10561);
nor U11023 (N_11023,N_10560,N_10586);
or U11024 (N_11024,N_10672,N_10534);
nor U11025 (N_11025,N_10663,N_10743);
and U11026 (N_11026,N_10787,N_10726);
nor U11027 (N_11027,N_10552,N_10702);
and U11028 (N_11028,N_10743,N_10757);
and U11029 (N_11029,N_10710,N_10549);
and U11030 (N_11030,N_10746,N_10602);
or U11031 (N_11031,N_10635,N_10684);
or U11032 (N_11032,N_10575,N_10645);
or U11033 (N_11033,N_10659,N_10689);
nand U11034 (N_11034,N_10574,N_10667);
nor U11035 (N_11035,N_10551,N_10702);
nor U11036 (N_11036,N_10553,N_10590);
nand U11037 (N_11037,N_10557,N_10623);
xor U11038 (N_11038,N_10710,N_10569);
or U11039 (N_11039,N_10634,N_10501);
and U11040 (N_11040,N_10551,N_10505);
and U11041 (N_11041,N_10540,N_10796);
nor U11042 (N_11042,N_10652,N_10695);
or U11043 (N_11043,N_10519,N_10687);
nor U11044 (N_11044,N_10583,N_10608);
xor U11045 (N_11045,N_10514,N_10759);
nor U11046 (N_11046,N_10620,N_10750);
or U11047 (N_11047,N_10589,N_10747);
nor U11048 (N_11048,N_10603,N_10547);
nand U11049 (N_11049,N_10789,N_10597);
nand U11050 (N_11050,N_10705,N_10687);
nand U11051 (N_11051,N_10523,N_10559);
xnor U11052 (N_11052,N_10762,N_10726);
nand U11053 (N_11053,N_10684,N_10795);
xnor U11054 (N_11054,N_10627,N_10779);
nor U11055 (N_11055,N_10636,N_10691);
nor U11056 (N_11056,N_10669,N_10764);
nor U11057 (N_11057,N_10623,N_10713);
or U11058 (N_11058,N_10719,N_10612);
nand U11059 (N_11059,N_10719,N_10541);
nor U11060 (N_11060,N_10790,N_10792);
and U11061 (N_11061,N_10560,N_10758);
nand U11062 (N_11062,N_10544,N_10738);
nor U11063 (N_11063,N_10507,N_10732);
nand U11064 (N_11064,N_10529,N_10731);
nand U11065 (N_11065,N_10562,N_10737);
and U11066 (N_11066,N_10705,N_10650);
or U11067 (N_11067,N_10776,N_10512);
nor U11068 (N_11068,N_10516,N_10798);
or U11069 (N_11069,N_10581,N_10582);
xor U11070 (N_11070,N_10670,N_10644);
or U11071 (N_11071,N_10628,N_10704);
xor U11072 (N_11072,N_10798,N_10557);
nand U11073 (N_11073,N_10665,N_10756);
and U11074 (N_11074,N_10792,N_10709);
or U11075 (N_11075,N_10746,N_10574);
nor U11076 (N_11076,N_10761,N_10762);
or U11077 (N_11077,N_10633,N_10697);
xnor U11078 (N_11078,N_10643,N_10516);
xnor U11079 (N_11079,N_10619,N_10773);
nand U11080 (N_11080,N_10521,N_10506);
nor U11081 (N_11081,N_10598,N_10783);
nand U11082 (N_11082,N_10525,N_10702);
or U11083 (N_11083,N_10527,N_10705);
nor U11084 (N_11084,N_10570,N_10504);
and U11085 (N_11085,N_10547,N_10526);
nand U11086 (N_11086,N_10689,N_10780);
and U11087 (N_11087,N_10735,N_10708);
nor U11088 (N_11088,N_10775,N_10517);
nor U11089 (N_11089,N_10747,N_10508);
nor U11090 (N_11090,N_10774,N_10775);
xnor U11091 (N_11091,N_10640,N_10618);
and U11092 (N_11092,N_10506,N_10507);
nand U11093 (N_11093,N_10515,N_10789);
or U11094 (N_11094,N_10543,N_10645);
xor U11095 (N_11095,N_10652,N_10728);
xnor U11096 (N_11096,N_10740,N_10708);
nand U11097 (N_11097,N_10526,N_10647);
and U11098 (N_11098,N_10583,N_10501);
xnor U11099 (N_11099,N_10509,N_10501);
nand U11100 (N_11100,N_10896,N_10953);
and U11101 (N_11101,N_11022,N_10913);
nand U11102 (N_11102,N_11044,N_11013);
and U11103 (N_11103,N_11019,N_10975);
or U11104 (N_11104,N_10915,N_11065);
or U11105 (N_11105,N_11058,N_11087);
nor U11106 (N_11106,N_10931,N_10956);
or U11107 (N_11107,N_10862,N_10992);
or U11108 (N_11108,N_10943,N_10853);
and U11109 (N_11109,N_10981,N_11016);
nand U11110 (N_11110,N_11025,N_11020);
and U11111 (N_11111,N_11047,N_10925);
or U11112 (N_11112,N_11011,N_11093);
nand U11113 (N_11113,N_11072,N_11073);
and U11114 (N_11114,N_10959,N_10825);
or U11115 (N_11115,N_11081,N_10946);
and U11116 (N_11116,N_10800,N_10918);
nand U11117 (N_11117,N_10979,N_10818);
and U11118 (N_11118,N_10985,N_10816);
nor U11119 (N_11119,N_10908,N_10916);
xor U11120 (N_11120,N_11027,N_10907);
or U11121 (N_11121,N_11039,N_11015);
xor U11122 (N_11122,N_10855,N_10941);
nand U11123 (N_11123,N_11001,N_10937);
nor U11124 (N_11124,N_10876,N_10938);
xnor U11125 (N_11125,N_10854,N_10973);
and U11126 (N_11126,N_10869,N_11002);
xnor U11127 (N_11127,N_10976,N_10830);
and U11128 (N_11128,N_10801,N_11099);
nand U11129 (N_11129,N_10902,N_10998);
nor U11130 (N_11130,N_11079,N_10927);
xnor U11131 (N_11131,N_10929,N_11036);
xnor U11132 (N_11132,N_10878,N_10965);
nor U11133 (N_11133,N_10993,N_10955);
nor U11134 (N_11134,N_10886,N_10815);
xnor U11135 (N_11135,N_10895,N_10819);
or U11136 (N_11136,N_11006,N_10926);
or U11137 (N_11137,N_11000,N_10906);
and U11138 (N_11138,N_10867,N_10870);
or U11139 (N_11139,N_10852,N_11010);
and U11140 (N_11140,N_10983,N_10813);
or U11141 (N_11141,N_10809,N_11014);
nand U11142 (N_11142,N_10921,N_10837);
and U11143 (N_11143,N_10866,N_10893);
and U11144 (N_11144,N_10849,N_11090);
nor U11145 (N_11145,N_11096,N_10880);
xor U11146 (N_11146,N_10887,N_10898);
nor U11147 (N_11147,N_10879,N_10865);
nor U11148 (N_11148,N_10804,N_10935);
nand U11149 (N_11149,N_11092,N_10835);
nor U11150 (N_11150,N_11028,N_10905);
nand U11151 (N_11151,N_11076,N_10970);
nand U11152 (N_11152,N_10950,N_11026);
nand U11153 (N_11153,N_11083,N_10924);
and U11154 (N_11154,N_10892,N_10997);
nor U11155 (N_11155,N_10874,N_11029);
and U11156 (N_11156,N_10994,N_10928);
and U11157 (N_11157,N_10919,N_10860);
and U11158 (N_11158,N_10971,N_10803);
nor U11159 (N_11159,N_10958,N_10805);
or U11160 (N_11160,N_10909,N_10881);
and U11161 (N_11161,N_11095,N_11082);
or U11162 (N_11162,N_10982,N_10939);
and U11163 (N_11163,N_10885,N_11080);
xnor U11164 (N_11164,N_10863,N_10999);
nor U11165 (N_11165,N_11059,N_11005);
nor U11166 (N_11166,N_10850,N_10996);
nor U11167 (N_11167,N_10872,N_10888);
xnor U11168 (N_11168,N_10920,N_10802);
xor U11169 (N_11169,N_10901,N_10810);
nor U11170 (N_11170,N_10891,N_10817);
nand U11171 (N_11171,N_10812,N_11089);
nand U11172 (N_11172,N_10960,N_10977);
nor U11173 (N_11173,N_10990,N_11038);
or U11174 (N_11174,N_10968,N_10875);
xor U11175 (N_11175,N_11049,N_11041);
nand U11176 (N_11176,N_11069,N_10808);
nand U11177 (N_11177,N_11066,N_11042);
nor U11178 (N_11178,N_11046,N_10814);
nand U11179 (N_11179,N_11060,N_10978);
nor U11180 (N_11180,N_10940,N_10832);
and U11181 (N_11181,N_10934,N_11032);
or U11182 (N_11182,N_10845,N_11030);
nand U11183 (N_11183,N_11062,N_11067);
and U11184 (N_11184,N_10884,N_10831);
nor U11185 (N_11185,N_10948,N_10932);
or U11186 (N_11186,N_10986,N_10889);
nand U11187 (N_11187,N_10848,N_11004);
and U11188 (N_11188,N_10841,N_10859);
or U11189 (N_11189,N_11053,N_10944);
or U11190 (N_11190,N_10840,N_10936);
or U11191 (N_11191,N_10836,N_10963);
nand U11192 (N_11192,N_10861,N_10806);
xnor U11193 (N_11193,N_10871,N_11084);
or U11194 (N_11194,N_11077,N_10822);
and U11195 (N_11195,N_11033,N_11031);
xor U11196 (N_11196,N_10829,N_10910);
xor U11197 (N_11197,N_11057,N_11034);
nor U11198 (N_11198,N_11070,N_11024);
nand U11199 (N_11199,N_10972,N_10966);
or U11200 (N_11200,N_10873,N_10917);
or U11201 (N_11201,N_10904,N_10952);
nor U11202 (N_11202,N_10967,N_10846);
nor U11203 (N_11203,N_10897,N_10995);
or U11204 (N_11204,N_10882,N_10949);
nor U11205 (N_11205,N_10933,N_10942);
nor U11206 (N_11206,N_10843,N_11018);
xnor U11207 (N_11207,N_10842,N_10828);
xor U11208 (N_11208,N_10838,N_10945);
nor U11209 (N_11209,N_11051,N_11045);
and U11210 (N_11210,N_10827,N_10868);
and U11211 (N_11211,N_11048,N_10883);
and U11212 (N_11212,N_10962,N_10844);
nand U11213 (N_11213,N_10847,N_10911);
or U11214 (N_11214,N_10894,N_11097);
xor U11215 (N_11215,N_11035,N_10930);
xor U11216 (N_11216,N_10820,N_10857);
nand U11217 (N_11217,N_10947,N_10961);
or U11218 (N_11218,N_10980,N_10991);
nor U11219 (N_11219,N_11086,N_10954);
or U11220 (N_11220,N_10912,N_10834);
nor U11221 (N_11221,N_10988,N_11075);
nand U11222 (N_11222,N_11050,N_10903);
nand U11223 (N_11223,N_11017,N_11055);
nor U11224 (N_11224,N_11008,N_10851);
xnor U11225 (N_11225,N_10839,N_11037);
nand U11226 (N_11226,N_11085,N_11052);
xor U11227 (N_11227,N_10823,N_11094);
nor U11228 (N_11228,N_10856,N_10957);
xnor U11229 (N_11229,N_11064,N_10900);
and U11230 (N_11230,N_11063,N_11003);
nor U11231 (N_11231,N_10890,N_10858);
and U11232 (N_11232,N_10951,N_10811);
xnor U11233 (N_11233,N_10984,N_11054);
nor U11234 (N_11234,N_11056,N_11021);
xor U11235 (N_11235,N_10833,N_10964);
nand U11236 (N_11236,N_11091,N_11007);
nor U11237 (N_11237,N_10877,N_11098);
nor U11238 (N_11238,N_10969,N_11088);
and U11239 (N_11239,N_11061,N_11009);
or U11240 (N_11240,N_10914,N_11040);
and U11241 (N_11241,N_11012,N_11074);
nand U11242 (N_11242,N_10826,N_10824);
and U11243 (N_11243,N_11068,N_10807);
and U11244 (N_11244,N_11043,N_11078);
or U11245 (N_11245,N_10899,N_10923);
nor U11246 (N_11246,N_10821,N_11023);
xnor U11247 (N_11247,N_11071,N_10922);
or U11248 (N_11248,N_10989,N_10987);
nand U11249 (N_11249,N_10864,N_10974);
nor U11250 (N_11250,N_11058,N_11014);
nor U11251 (N_11251,N_10951,N_11054);
nand U11252 (N_11252,N_10991,N_10933);
nand U11253 (N_11253,N_10922,N_10883);
xor U11254 (N_11254,N_10860,N_10875);
or U11255 (N_11255,N_11011,N_11006);
or U11256 (N_11256,N_11000,N_11064);
nor U11257 (N_11257,N_10871,N_10943);
or U11258 (N_11258,N_11039,N_10832);
nand U11259 (N_11259,N_10928,N_10972);
or U11260 (N_11260,N_11044,N_10954);
and U11261 (N_11261,N_11088,N_11027);
nand U11262 (N_11262,N_11032,N_10824);
nand U11263 (N_11263,N_10990,N_10887);
and U11264 (N_11264,N_10938,N_10940);
or U11265 (N_11265,N_10802,N_10942);
and U11266 (N_11266,N_10975,N_10951);
and U11267 (N_11267,N_10837,N_10932);
nor U11268 (N_11268,N_10949,N_10829);
nor U11269 (N_11269,N_11073,N_10874);
xor U11270 (N_11270,N_10889,N_10970);
nor U11271 (N_11271,N_11088,N_10934);
xor U11272 (N_11272,N_10807,N_10966);
xor U11273 (N_11273,N_11068,N_10942);
nor U11274 (N_11274,N_11036,N_10938);
nand U11275 (N_11275,N_11041,N_10835);
nand U11276 (N_11276,N_11082,N_10921);
xor U11277 (N_11277,N_11075,N_10870);
nand U11278 (N_11278,N_11084,N_10895);
xnor U11279 (N_11279,N_10863,N_11037);
and U11280 (N_11280,N_11088,N_11019);
xor U11281 (N_11281,N_10950,N_11021);
and U11282 (N_11282,N_10927,N_10992);
xnor U11283 (N_11283,N_10916,N_10923);
and U11284 (N_11284,N_11061,N_10842);
or U11285 (N_11285,N_10855,N_10931);
nand U11286 (N_11286,N_10811,N_10853);
nand U11287 (N_11287,N_10833,N_10941);
or U11288 (N_11288,N_10950,N_10874);
and U11289 (N_11289,N_11000,N_11058);
and U11290 (N_11290,N_11077,N_10803);
and U11291 (N_11291,N_10972,N_10924);
and U11292 (N_11292,N_10811,N_10844);
and U11293 (N_11293,N_10968,N_10822);
xor U11294 (N_11294,N_10811,N_11014);
and U11295 (N_11295,N_10980,N_10850);
nand U11296 (N_11296,N_11019,N_11059);
nand U11297 (N_11297,N_10809,N_10926);
and U11298 (N_11298,N_10919,N_11035);
nand U11299 (N_11299,N_10841,N_11002);
xor U11300 (N_11300,N_10875,N_10922);
or U11301 (N_11301,N_11000,N_11009);
nand U11302 (N_11302,N_10831,N_11051);
nor U11303 (N_11303,N_10835,N_10895);
xor U11304 (N_11304,N_11051,N_10958);
nor U11305 (N_11305,N_10843,N_10996);
nor U11306 (N_11306,N_10807,N_11020);
nand U11307 (N_11307,N_10982,N_10961);
nor U11308 (N_11308,N_10827,N_11037);
nor U11309 (N_11309,N_10822,N_10978);
nor U11310 (N_11310,N_11076,N_10983);
nor U11311 (N_11311,N_10985,N_10918);
or U11312 (N_11312,N_10976,N_10915);
xor U11313 (N_11313,N_11078,N_11007);
and U11314 (N_11314,N_11055,N_10978);
and U11315 (N_11315,N_11053,N_10907);
or U11316 (N_11316,N_10818,N_10813);
or U11317 (N_11317,N_11083,N_10960);
and U11318 (N_11318,N_10911,N_10954);
and U11319 (N_11319,N_10936,N_11073);
nor U11320 (N_11320,N_10892,N_10941);
nand U11321 (N_11321,N_10952,N_10887);
or U11322 (N_11322,N_10900,N_10814);
and U11323 (N_11323,N_11044,N_10846);
nor U11324 (N_11324,N_11083,N_10815);
nand U11325 (N_11325,N_11060,N_10916);
and U11326 (N_11326,N_11052,N_10966);
nor U11327 (N_11327,N_10915,N_10941);
or U11328 (N_11328,N_10828,N_10910);
nand U11329 (N_11329,N_10985,N_10942);
nand U11330 (N_11330,N_10837,N_10889);
and U11331 (N_11331,N_10867,N_11063);
xnor U11332 (N_11332,N_11088,N_10823);
and U11333 (N_11333,N_10998,N_10896);
and U11334 (N_11334,N_10961,N_10833);
or U11335 (N_11335,N_10804,N_11004);
nand U11336 (N_11336,N_10987,N_10970);
or U11337 (N_11337,N_10929,N_11098);
nor U11338 (N_11338,N_10937,N_10817);
nand U11339 (N_11339,N_11060,N_10829);
nand U11340 (N_11340,N_11026,N_10929);
xnor U11341 (N_11341,N_10924,N_10957);
nand U11342 (N_11342,N_10865,N_11039);
and U11343 (N_11343,N_10907,N_10975);
nand U11344 (N_11344,N_11038,N_10971);
or U11345 (N_11345,N_10849,N_10882);
and U11346 (N_11346,N_10943,N_11029);
nor U11347 (N_11347,N_10843,N_10805);
and U11348 (N_11348,N_11083,N_10999);
or U11349 (N_11349,N_10844,N_10893);
and U11350 (N_11350,N_11091,N_11064);
nor U11351 (N_11351,N_10955,N_10838);
and U11352 (N_11352,N_10818,N_10960);
xnor U11353 (N_11353,N_11054,N_11009);
xor U11354 (N_11354,N_11012,N_11096);
or U11355 (N_11355,N_10999,N_10907);
nand U11356 (N_11356,N_10866,N_11018);
nand U11357 (N_11357,N_10949,N_10977);
and U11358 (N_11358,N_10889,N_10806);
or U11359 (N_11359,N_10929,N_11037);
or U11360 (N_11360,N_10871,N_10843);
and U11361 (N_11361,N_10979,N_10838);
or U11362 (N_11362,N_10930,N_10836);
and U11363 (N_11363,N_10953,N_10881);
xor U11364 (N_11364,N_11010,N_11029);
nand U11365 (N_11365,N_10943,N_10867);
or U11366 (N_11366,N_10862,N_11007);
xor U11367 (N_11367,N_11049,N_10924);
xor U11368 (N_11368,N_10888,N_10853);
nand U11369 (N_11369,N_10816,N_11059);
nor U11370 (N_11370,N_11069,N_10846);
xnor U11371 (N_11371,N_10822,N_11048);
or U11372 (N_11372,N_10827,N_10925);
or U11373 (N_11373,N_10836,N_11013);
and U11374 (N_11374,N_11042,N_10974);
or U11375 (N_11375,N_10975,N_11014);
or U11376 (N_11376,N_10851,N_10900);
xor U11377 (N_11377,N_10959,N_10984);
xor U11378 (N_11378,N_10835,N_10830);
xor U11379 (N_11379,N_10979,N_11023);
xnor U11380 (N_11380,N_10824,N_10943);
nor U11381 (N_11381,N_10856,N_10914);
nor U11382 (N_11382,N_11004,N_10912);
nor U11383 (N_11383,N_10932,N_10864);
and U11384 (N_11384,N_11000,N_10964);
nor U11385 (N_11385,N_10802,N_10925);
nand U11386 (N_11386,N_10881,N_11080);
or U11387 (N_11387,N_11089,N_10924);
nor U11388 (N_11388,N_11026,N_10968);
nand U11389 (N_11389,N_11039,N_10942);
nor U11390 (N_11390,N_10855,N_11057);
nor U11391 (N_11391,N_11062,N_11038);
and U11392 (N_11392,N_10979,N_10866);
or U11393 (N_11393,N_10963,N_10973);
xor U11394 (N_11394,N_10837,N_10930);
xnor U11395 (N_11395,N_10855,N_11061);
or U11396 (N_11396,N_11015,N_10981);
nand U11397 (N_11397,N_10944,N_10932);
xor U11398 (N_11398,N_10872,N_11093);
and U11399 (N_11399,N_11040,N_10881);
xor U11400 (N_11400,N_11139,N_11233);
xnor U11401 (N_11401,N_11379,N_11200);
and U11402 (N_11402,N_11373,N_11247);
or U11403 (N_11403,N_11235,N_11337);
or U11404 (N_11404,N_11123,N_11274);
and U11405 (N_11405,N_11204,N_11210);
or U11406 (N_11406,N_11276,N_11358);
nand U11407 (N_11407,N_11132,N_11342);
or U11408 (N_11408,N_11107,N_11326);
nand U11409 (N_11409,N_11320,N_11258);
and U11410 (N_11410,N_11231,N_11178);
xnor U11411 (N_11411,N_11382,N_11248);
nor U11412 (N_11412,N_11142,N_11369);
or U11413 (N_11413,N_11191,N_11372);
nor U11414 (N_11414,N_11167,N_11182);
xor U11415 (N_11415,N_11209,N_11227);
or U11416 (N_11416,N_11270,N_11309);
or U11417 (N_11417,N_11376,N_11278);
and U11418 (N_11418,N_11144,N_11251);
or U11419 (N_11419,N_11184,N_11224);
nor U11420 (N_11420,N_11230,N_11229);
xor U11421 (N_11421,N_11194,N_11130);
or U11422 (N_11422,N_11299,N_11305);
xor U11423 (N_11423,N_11237,N_11307);
nand U11424 (N_11424,N_11391,N_11164);
xnor U11425 (N_11425,N_11160,N_11202);
or U11426 (N_11426,N_11253,N_11281);
xnor U11427 (N_11427,N_11198,N_11300);
or U11428 (N_11428,N_11241,N_11315);
nor U11429 (N_11429,N_11216,N_11374);
nand U11430 (N_11430,N_11151,N_11285);
xor U11431 (N_11431,N_11311,N_11279);
xnor U11432 (N_11432,N_11163,N_11124);
nand U11433 (N_11433,N_11322,N_11220);
nor U11434 (N_11434,N_11383,N_11221);
and U11435 (N_11435,N_11357,N_11133);
or U11436 (N_11436,N_11206,N_11117);
and U11437 (N_11437,N_11381,N_11156);
and U11438 (N_11438,N_11174,N_11214);
xnor U11439 (N_11439,N_11218,N_11265);
nor U11440 (N_11440,N_11323,N_11339);
or U11441 (N_11441,N_11330,N_11361);
xnor U11442 (N_11442,N_11336,N_11201);
nand U11443 (N_11443,N_11319,N_11189);
and U11444 (N_11444,N_11101,N_11177);
nor U11445 (N_11445,N_11303,N_11169);
xnor U11446 (N_11446,N_11390,N_11368);
or U11447 (N_11447,N_11143,N_11115);
and U11448 (N_11448,N_11212,N_11145);
xor U11449 (N_11449,N_11287,N_11293);
xor U11450 (N_11450,N_11297,N_11329);
and U11451 (N_11451,N_11304,N_11199);
xor U11452 (N_11452,N_11255,N_11347);
nor U11453 (N_11453,N_11110,N_11364);
and U11454 (N_11454,N_11187,N_11360);
or U11455 (N_11455,N_11354,N_11331);
and U11456 (N_11456,N_11334,N_11207);
nor U11457 (N_11457,N_11134,N_11240);
nand U11458 (N_11458,N_11112,N_11302);
and U11459 (N_11459,N_11106,N_11262);
or U11460 (N_11460,N_11286,N_11263);
nand U11461 (N_11461,N_11128,N_11138);
xor U11462 (N_11462,N_11173,N_11245);
and U11463 (N_11463,N_11321,N_11388);
nand U11464 (N_11464,N_11393,N_11272);
nand U11465 (N_11465,N_11399,N_11346);
nor U11466 (N_11466,N_11103,N_11100);
and U11467 (N_11467,N_11148,N_11215);
and U11468 (N_11468,N_11380,N_11385);
nand U11469 (N_11469,N_11291,N_11183);
and U11470 (N_11470,N_11232,N_11118);
or U11471 (N_11471,N_11186,N_11294);
or U11472 (N_11472,N_11219,N_11111);
xnor U11473 (N_11473,N_11359,N_11153);
nor U11474 (N_11474,N_11197,N_11292);
nand U11475 (N_11475,N_11140,N_11289);
xnor U11476 (N_11476,N_11172,N_11332);
and U11477 (N_11477,N_11158,N_11257);
and U11478 (N_11478,N_11324,N_11367);
or U11479 (N_11479,N_11252,N_11389);
and U11480 (N_11480,N_11377,N_11238);
xor U11481 (N_11481,N_11180,N_11314);
nand U11482 (N_11482,N_11121,N_11290);
or U11483 (N_11483,N_11375,N_11205);
nor U11484 (N_11484,N_11269,N_11341);
nand U11485 (N_11485,N_11275,N_11335);
nor U11486 (N_11486,N_11333,N_11176);
nand U11487 (N_11487,N_11365,N_11308);
xnor U11488 (N_11488,N_11296,N_11366);
nor U11489 (N_11489,N_11259,N_11152);
or U11490 (N_11490,N_11126,N_11317);
nor U11491 (N_11491,N_11120,N_11190);
and U11492 (N_11492,N_11243,N_11394);
or U11493 (N_11493,N_11155,N_11280);
nor U11494 (N_11494,N_11246,N_11351);
nor U11495 (N_11495,N_11223,N_11104);
nor U11496 (N_11496,N_11114,N_11256);
nand U11497 (N_11497,N_11159,N_11325);
nand U11498 (N_11498,N_11306,N_11318);
nor U11499 (N_11499,N_11378,N_11298);
xnor U11500 (N_11500,N_11195,N_11340);
or U11501 (N_11501,N_11203,N_11386);
and U11502 (N_11502,N_11149,N_11397);
and U11503 (N_11503,N_11244,N_11157);
nand U11504 (N_11504,N_11113,N_11168);
and U11505 (N_11505,N_11267,N_11328);
nand U11506 (N_11506,N_11362,N_11208);
xor U11507 (N_11507,N_11225,N_11363);
and U11508 (N_11508,N_11154,N_11355);
xor U11509 (N_11509,N_11119,N_11356);
xnor U11510 (N_11510,N_11193,N_11350);
nor U11511 (N_11511,N_11310,N_11338);
nor U11512 (N_11512,N_11162,N_11185);
nand U11513 (N_11513,N_11316,N_11165);
or U11514 (N_11514,N_11348,N_11109);
xor U11515 (N_11515,N_11129,N_11349);
or U11516 (N_11516,N_11370,N_11228);
and U11517 (N_11517,N_11395,N_11384);
and U11518 (N_11518,N_11261,N_11249);
and U11519 (N_11519,N_11283,N_11282);
nor U11520 (N_11520,N_11313,N_11284);
and U11521 (N_11521,N_11108,N_11226);
or U11522 (N_11522,N_11312,N_11398);
nor U11523 (N_11523,N_11141,N_11327);
nor U11524 (N_11524,N_11268,N_11171);
or U11525 (N_11525,N_11371,N_11136);
and U11526 (N_11526,N_11137,N_11102);
nor U11527 (N_11527,N_11295,N_11217);
and U11528 (N_11528,N_11239,N_11122);
xor U11529 (N_11529,N_11188,N_11196);
nor U11530 (N_11530,N_11135,N_11392);
nor U11531 (N_11531,N_11192,N_11234);
and U11532 (N_11532,N_11211,N_11260);
nand U11533 (N_11533,N_11271,N_11288);
nand U11534 (N_11534,N_11254,N_11146);
and U11535 (N_11535,N_11105,N_11166);
or U11536 (N_11536,N_11161,N_11127);
and U11537 (N_11537,N_11387,N_11236);
nand U11538 (N_11538,N_11175,N_11222);
or U11539 (N_11539,N_11353,N_11125);
or U11540 (N_11540,N_11352,N_11147);
and U11541 (N_11541,N_11301,N_11343);
or U11542 (N_11542,N_11150,N_11213);
nor U11543 (N_11543,N_11264,N_11181);
nor U11544 (N_11544,N_11266,N_11250);
nor U11545 (N_11545,N_11116,N_11170);
or U11546 (N_11546,N_11242,N_11131);
and U11547 (N_11547,N_11277,N_11179);
xnor U11548 (N_11548,N_11344,N_11396);
nor U11549 (N_11549,N_11273,N_11345);
and U11550 (N_11550,N_11202,N_11229);
nor U11551 (N_11551,N_11273,N_11330);
nor U11552 (N_11552,N_11177,N_11140);
nand U11553 (N_11553,N_11181,N_11262);
nor U11554 (N_11554,N_11264,N_11205);
nor U11555 (N_11555,N_11373,N_11128);
nor U11556 (N_11556,N_11117,N_11189);
or U11557 (N_11557,N_11213,N_11384);
xor U11558 (N_11558,N_11399,N_11283);
nor U11559 (N_11559,N_11379,N_11212);
nor U11560 (N_11560,N_11373,N_11205);
nand U11561 (N_11561,N_11303,N_11162);
nand U11562 (N_11562,N_11123,N_11199);
or U11563 (N_11563,N_11298,N_11197);
and U11564 (N_11564,N_11159,N_11192);
xnor U11565 (N_11565,N_11315,N_11224);
xor U11566 (N_11566,N_11233,N_11311);
xnor U11567 (N_11567,N_11357,N_11248);
xnor U11568 (N_11568,N_11118,N_11327);
nor U11569 (N_11569,N_11256,N_11352);
nand U11570 (N_11570,N_11280,N_11153);
or U11571 (N_11571,N_11164,N_11240);
nor U11572 (N_11572,N_11162,N_11362);
xnor U11573 (N_11573,N_11350,N_11288);
xnor U11574 (N_11574,N_11218,N_11354);
or U11575 (N_11575,N_11247,N_11336);
nor U11576 (N_11576,N_11241,N_11116);
nand U11577 (N_11577,N_11337,N_11174);
xnor U11578 (N_11578,N_11387,N_11162);
xnor U11579 (N_11579,N_11198,N_11206);
and U11580 (N_11580,N_11283,N_11144);
or U11581 (N_11581,N_11121,N_11193);
or U11582 (N_11582,N_11279,N_11263);
nand U11583 (N_11583,N_11156,N_11218);
nor U11584 (N_11584,N_11204,N_11386);
nor U11585 (N_11585,N_11375,N_11266);
and U11586 (N_11586,N_11272,N_11260);
nand U11587 (N_11587,N_11107,N_11300);
or U11588 (N_11588,N_11263,N_11225);
xnor U11589 (N_11589,N_11242,N_11285);
nand U11590 (N_11590,N_11256,N_11392);
nor U11591 (N_11591,N_11313,N_11166);
nand U11592 (N_11592,N_11173,N_11323);
xnor U11593 (N_11593,N_11399,N_11306);
nand U11594 (N_11594,N_11245,N_11104);
xnor U11595 (N_11595,N_11296,N_11354);
nor U11596 (N_11596,N_11118,N_11205);
nand U11597 (N_11597,N_11381,N_11110);
nand U11598 (N_11598,N_11288,N_11236);
or U11599 (N_11599,N_11216,N_11372);
nor U11600 (N_11600,N_11152,N_11289);
and U11601 (N_11601,N_11399,N_11246);
xor U11602 (N_11602,N_11261,N_11359);
and U11603 (N_11603,N_11305,N_11123);
nand U11604 (N_11604,N_11102,N_11114);
nand U11605 (N_11605,N_11150,N_11235);
nand U11606 (N_11606,N_11155,N_11381);
and U11607 (N_11607,N_11327,N_11200);
xnor U11608 (N_11608,N_11265,N_11229);
nor U11609 (N_11609,N_11338,N_11346);
xnor U11610 (N_11610,N_11373,N_11243);
nand U11611 (N_11611,N_11141,N_11167);
nand U11612 (N_11612,N_11252,N_11142);
nand U11613 (N_11613,N_11207,N_11127);
or U11614 (N_11614,N_11101,N_11156);
nor U11615 (N_11615,N_11292,N_11324);
and U11616 (N_11616,N_11277,N_11122);
xnor U11617 (N_11617,N_11360,N_11136);
or U11618 (N_11618,N_11297,N_11299);
nand U11619 (N_11619,N_11168,N_11207);
nor U11620 (N_11620,N_11385,N_11342);
nand U11621 (N_11621,N_11212,N_11229);
and U11622 (N_11622,N_11239,N_11249);
nand U11623 (N_11623,N_11150,N_11356);
nand U11624 (N_11624,N_11347,N_11312);
or U11625 (N_11625,N_11110,N_11144);
and U11626 (N_11626,N_11339,N_11139);
nor U11627 (N_11627,N_11327,N_11195);
nand U11628 (N_11628,N_11174,N_11207);
or U11629 (N_11629,N_11187,N_11308);
nand U11630 (N_11630,N_11307,N_11201);
or U11631 (N_11631,N_11365,N_11321);
and U11632 (N_11632,N_11106,N_11344);
or U11633 (N_11633,N_11150,N_11188);
nor U11634 (N_11634,N_11249,N_11399);
or U11635 (N_11635,N_11385,N_11298);
and U11636 (N_11636,N_11212,N_11255);
nor U11637 (N_11637,N_11198,N_11214);
xnor U11638 (N_11638,N_11279,N_11137);
or U11639 (N_11639,N_11242,N_11204);
or U11640 (N_11640,N_11231,N_11286);
xor U11641 (N_11641,N_11387,N_11106);
xnor U11642 (N_11642,N_11159,N_11313);
and U11643 (N_11643,N_11316,N_11307);
or U11644 (N_11644,N_11177,N_11319);
nand U11645 (N_11645,N_11135,N_11134);
nor U11646 (N_11646,N_11389,N_11390);
xnor U11647 (N_11647,N_11259,N_11242);
or U11648 (N_11648,N_11280,N_11187);
and U11649 (N_11649,N_11166,N_11294);
and U11650 (N_11650,N_11169,N_11159);
and U11651 (N_11651,N_11196,N_11342);
xor U11652 (N_11652,N_11149,N_11345);
and U11653 (N_11653,N_11319,N_11179);
and U11654 (N_11654,N_11351,N_11370);
or U11655 (N_11655,N_11295,N_11359);
nor U11656 (N_11656,N_11333,N_11312);
or U11657 (N_11657,N_11363,N_11109);
xnor U11658 (N_11658,N_11176,N_11110);
nand U11659 (N_11659,N_11325,N_11115);
xor U11660 (N_11660,N_11112,N_11393);
nor U11661 (N_11661,N_11255,N_11238);
or U11662 (N_11662,N_11221,N_11244);
or U11663 (N_11663,N_11119,N_11225);
xnor U11664 (N_11664,N_11270,N_11188);
and U11665 (N_11665,N_11287,N_11323);
nand U11666 (N_11666,N_11352,N_11267);
or U11667 (N_11667,N_11342,N_11387);
and U11668 (N_11668,N_11113,N_11118);
nand U11669 (N_11669,N_11306,N_11346);
xnor U11670 (N_11670,N_11145,N_11113);
nor U11671 (N_11671,N_11287,N_11168);
and U11672 (N_11672,N_11298,N_11249);
and U11673 (N_11673,N_11269,N_11213);
and U11674 (N_11674,N_11260,N_11301);
and U11675 (N_11675,N_11107,N_11345);
nor U11676 (N_11676,N_11171,N_11164);
or U11677 (N_11677,N_11252,N_11213);
nand U11678 (N_11678,N_11262,N_11100);
nand U11679 (N_11679,N_11357,N_11123);
and U11680 (N_11680,N_11366,N_11260);
nor U11681 (N_11681,N_11301,N_11119);
and U11682 (N_11682,N_11382,N_11282);
or U11683 (N_11683,N_11108,N_11207);
nand U11684 (N_11684,N_11305,N_11289);
nand U11685 (N_11685,N_11256,N_11101);
or U11686 (N_11686,N_11279,N_11367);
nor U11687 (N_11687,N_11147,N_11215);
and U11688 (N_11688,N_11280,N_11348);
nor U11689 (N_11689,N_11179,N_11377);
nand U11690 (N_11690,N_11298,N_11290);
xnor U11691 (N_11691,N_11176,N_11221);
nor U11692 (N_11692,N_11392,N_11171);
xor U11693 (N_11693,N_11176,N_11278);
or U11694 (N_11694,N_11397,N_11135);
nand U11695 (N_11695,N_11236,N_11212);
nand U11696 (N_11696,N_11347,N_11357);
nand U11697 (N_11697,N_11367,N_11111);
or U11698 (N_11698,N_11100,N_11348);
and U11699 (N_11699,N_11373,N_11397);
xnor U11700 (N_11700,N_11688,N_11456);
nand U11701 (N_11701,N_11408,N_11675);
or U11702 (N_11702,N_11462,N_11435);
nor U11703 (N_11703,N_11460,N_11407);
nand U11704 (N_11704,N_11592,N_11447);
xnor U11705 (N_11705,N_11576,N_11562);
xnor U11706 (N_11706,N_11652,N_11653);
nand U11707 (N_11707,N_11659,N_11611);
xor U11708 (N_11708,N_11628,N_11531);
nor U11709 (N_11709,N_11672,N_11547);
and U11710 (N_11710,N_11481,N_11663);
or U11711 (N_11711,N_11596,N_11535);
and U11712 (N_11712,N_11540,N_11406);
nand U11713 (N_11713,N_11421,N_11486);
or U11714 (N_11714,N_11616,N_11420);
nand U11715 (N_11715,N_11503,N_11433);
nand U11716 (N_11716,N_11482,N_11682);
xor U11717 (N_11717,N_11483,N_11475);
or U11718 (N_11718,N_11464,N_11630);
and U11719 (N_11719,N_11454,N_11664);
and U11720 (N_11720,N_11555,N_11466);
nand U11721 (N_11721,N_11666,N_11614);
or U11722 (N_11722,N_11650,N_11570);
and U11723 (N_11723,N_11455,N_11677);
xor U11724 (N_11724,N_11557,N_11444);
xor U11725 (N_11725,N_11591,N_11595);
nor U11726 (N_11726,N_11631,N_11634);
nand U11727 (N_11727,N_11645,N_11641);
nor U11728 (N_11728,N_11495,N_11498);
nand U11729 (N_11729,N_11654,N_11448);
nand U11730 (N_11730,N_11585,N_11425);
and U11731 (N_11731,N_11522,N_11567);
xnor U11732 (N_11732,N_11623,N_11440);
nor U11733 (N_11733,N_11497,N_11507);
nor U11734 (N_11734,N_11584,N_11568);
and U11735 (N_11735,N_11443,N_11457);
nor U11736 (N_11736,N_11441,N_11476);
or U11737 (N_11737,N_11519,N_11680);
nand U11738 (N_11738,N_11501,N_11661);
nor U11739 (N_11739,N_11619,N_11468);
xnor U11740 (N_11740,N_11606,N_11692);
and U11741 (N_11741,N_11569,N_11473);
xor U11742 (N_11742,N_11400,N_11613);
nor U11743 (N_11743,N_11413,N_11496);
nor U11744 (N_11744,N_11532,N_11494);
or U11745 (N_11745,N_11551,N_11453);
or U11746 (N_11746,N_11626,N_11423);
or U11747 (N_11747,N_11644,N_11512);
xor U11748 (N_11748,N_11499,N_11548);
or U11749 (N_11749,N_11667,N_11635);
nor U11750 (N_11750,N_11602,N_11511);
nor U11751 (N_11751,N_11597,N_11523);
nor U11752 (N_11752,N_11693,N_11546);
and U11753 (N_11753,N_11533,N_11428);
nand U11754 (N_11754,N_11474,N_11579);
xor U11755 (N_11755,N_11651,N_11636);
or U11756 (N_11756,N_11446,N_11638);
or U11757 (N_11757,N_11450,N_11479);
and U11758 (N_11758,N_11480,N_11544);
nor U11759 (N_11759,N_11605,N_11669);
nand U11760 (N_11760,N_11678,N_11615);
nor U11761 (N_11761,N_11655,N_11445);
xnor U11762 (N_11762,N_11612,N_11552);
xor U11763 (N_11763,N_11657,N_11604);
or U11764 (N_11764,N_11403,N_11465);
and U11765 (N_11765,N_11558,N_11639);
and U11766 (N_11766,N_11405,N_11541);
xnor U11767 (N_11767,N_11502,N_11438);
nor U11768 (N_11768,N_11637,N_11416);
or U11769 (N_11769,N_11643,N_11593);
xnor U11770 (N_11770,N_11472,N_11571);
and U11771 (N_11771,N_11572,N_11599);
nor U11772 (N_11772,N_11439,N_11536);
xor U11773 (N_11773,N_11469,N_11418);
or U11774 (N_11774,N_11500,N_11538);
nand U11775 (N_11775,N_11437,N_11573);
nor U11776 (N_11776,N_11426,N_11624);
xnor U11777 (N_11777,N_11696,N_11577);
xnor U11778 (N_11778,N_11566,N_11698);
xnor U11779 (N_11779,N_11539,N_11594);
nor U11780 (N_11780,N_11485,N_11581);
and U11781 (N_11781,N_11560,N_11633);
nor U11782 (N_11782,N_11561,N_11489);
xor U11783 (N_11783,N_11665,N_11687);
nor U11784 (N_11784,N_11411,N_11600);
xor U11785 (N_11785,N_11549,N_11658);
nand U11786 (N_11786,N_11563,N_11580);
xnor U11787 (N_11787,N_11543,N_11598);
nor U11788 (N_11788,N_11424,N_11526);
nand U11789 (N_11789,N_11461,N_11647);
or U11790 (N_11790,N_11554,N_11686);
xnor U11791 (N_11791,N_11574,N_11695);
xnor U11792 (N_11792,N_11509,N_11430);
xnor U11793 (N_11793,N_11458,N_11514);
or U11794 (N_11794,N_11697,N_11559);
nand U11795 (N_11795,N_11451,N_11401);
or U11796 (N_11796,N_11685,N_11510);
xnor U11797 (N_11797,N_11404,N_11625);
nor U11798 (N_11798,N_11436,N_11691);
xor U11799 (N_11799,N_11492,N_11449);
or U11800 (N_11800,N_11518,N_11459);
nor U11801 (N_11801,N_11431,N_11530);
nor U11802 (N_11802,N_11627,N_11505);
and U11803 (N_11803,N_11565,N_11506);
nor U11804 (N_11804,N_11681,N_11684);
nand U11805 (N_11805,N_11412,N_11545);
xnor U11806 (N_11806,N_11521,N_11662);
and U11807 (N_11807,N_11640,N_11402);
xnor U11808 (N_11808,N_11427,N_11542);
and U11809 (N_11809,N_11415,N_11582);
and U11810 (N_11810,N_11478,N_11674);
or U11811 (N_11811,N_11537,N_11620);
and U11812 (N_11812,N_11491,N_11670);
and U11813 (N_11813,N_11578,N_11525);
nand U11814 (N_11814,N_11528,N_11660);
or U11815 (N_11815,N_11527,N_11524);
xor U11816 (N_11816,N_11487,N_11609);
or U11817 (N_11817,N_11699,N_11588);
or U11818 (N_11818,N_11419,N_11434);
or U11819 (N_11819,N_11583,N_11610);
xor U11820 (N_11820,N_11410,N_11417);
xnor U11821 (N_11821,N_11586,N_11467);
nor U11822 (N_11822,N_11587,N_11556);
and U11823 (N_11823,N_11589,N_11490);
xor U11824 (N_11824,N_11508,N_11694);
nor U11825 (N_11825,N_11504,N_11683);
xnor U11826 (N_11826,N_11590,N_11516);
nor U11827 (N_11827,N_11575,N_11515);
or U11828 (N_11828,N_11493,N_11642);
or U11829 (N_11829,N_11632,N_11690);
nor U11830 (N_11830,N_11679,N_11648);
and U11831 (N_11831,N_11409,N_11520);
nand U11832 (N_11832,N_11432,N_11617);
nand U11833 (N_11833,N_11517,N_11470);
or U11834 (N_11834,N_11689,N_11429);
and U11835 (N_11835,N_11603,N_11471);
xor U11836 (N_11836,N_11484,N_11452);
and U11837 (N_11837,N_11422,N_11488);
or U11838 (N_11838,N_11608,N_11477);
and U11839 (N_11839,N_11607,N_11463);
nand U11840 (N_11840,N_11649,N_11629);
xnor U11841 (N_11841,N_11534,N_11553);
nand U11842 (N_11842,N_11622,N_11513);
or U11843 (N_11843,N_11673,N_11529);
or U11844 (N_11844,N_11601,N_11656);
nand U11845 (N_11845,N_11414,N_11646);
or U11846 (N_11846,N_11442,N_11621);
nor U11847 (N_11847,N_11671,N_11564);
xor U11848 (N_11848,N_11668,N_11676);
xor U11849 (N_11849,N_11550,N_11618);
nor U11850 (N_11850,N_11421,N_11595);
xnor U11851 (N_11851,N_11626,N_11655);
nor U11852 (N_11852,N_11436,N_11459);
and U11853 (N_11853,N_11610,N_11595);
or U11854 (N_11854,N_11551,N_11582);
xor U11855 (N_11855,N_11531,N_11430);
nor U11856 (N_11856,N_11650,N_11487);
xnor U11857 (N_11857,N_11547,N_11461);
xnor U11858 (N_11858,N_11626,N_11430);
nor U11859 (N_11859,N_11485,N_11429);
or U11860 (N_11860,N_11656,N_11599);
xor U11861 (N_11861,N_11579,N_11537);
nor U11862 (N_11862,N_11481,N_11431);
xnor U11863 (N_11863,N_11629,N_11479);
nor U11864 (N_11864,N_11414,N_11508);
xor U11865 (N_11865,N_11492,N_11519);
nor U11866 (N_11866,N_11528,N_11461);
nand U11867 (N_11867,N_11577,N_11578);
nand U11868 (N_11868,N_11428,N_11674);
and U11869 (N_11869,N_11545,N_11510);
xor U11870 (N_11870,N_11504,N_11576);
xor U11871 (N_11871,N_11465,N_11616);
nand U11872 (N_11872,N_11644,N_11683);
nand U11873 (N_11873,N_11528,N_11498);
nand U11874 (N_11874,N_11481,N_11658);
nand U11875 (N_11875,N_11567,N_11545);
or U11876 (N_11876,N_11601,N_11434);
nand U11877 (N_11877,N_11420,N_11695);
or U11878 (N_11878,N_11597,N_11445);
or U11879 (N_11879,N_11650,N_11406);
xor U11880 (N_11880,N_11627,N_11644);
and U11881 (N_11881,N_11528,N_11565);
nor U11882 (N_11882,N_11628,N_11667);
xor U11883 (N_11883,N_11667,N_11652);
nand U11884 (N_11884,N_11533,N_11669);
nand U11885 (N_11885,N_11487,N_11416);
nor U11886 (N_11886,N_11468,N_11477);
nand U11887 (N_11887,N_11673,N_11630);
nor U11888 (N_11888,N_11542,N_11447);
or U11889 (N_11889,N_11698,N_11599);
and U11890 (N_11890,N_11611,N_11685);
nor U11891 (N_11891,N_11648,N_11438);
nor U11892 (N_11892,N_11491,N_11629);
xnor U11893 (N_11893,N_11511,N_11653);
nor U11894 (N_11894,N_11699,N_11485);
or U11895 (N_11895,N_11453,N_11522);
nor U11896 (N_11896,N_11430,N_11445);
or U11897 (N_11897,N_11689,N_11563);
xnor U11898 (N_11898,N_11539,N_11495);
nand U11899 (N_11899,N_11665,N_11635);
and U11900 (N_11900,N_11697,N_11647);
nor U11901 (N_11901,N_11541,N_11626);
and U11902 (N_11902,N_11630,N_11512);
xnor U11903 (N_11903,N_11451,N_11602);
and U11904 (N_11904,N_11473,N_11692);
xor U11905 (N_11905,N_11413,N_11417);
and U11906 (N_11906,N_11638,N_11505);
nor U11907 (N_11907,N_11649,N_11567);
and U11908 (N_11908,N_11562,N_11692);
and U11909 (N_11909,N_11454,N_11676);
or U11910 (N_11910,N_11666,N_11583);
nor U11911 (N_11911,N_11555,N_11632);
and U11912 (N_11912,N_11556,N_11563);
xnor U11913 (N_11913,N_11558,N_11553);
xnor U11914 (N_11914,N_11454,N_11613);
nor U11915 (N_11915,N_11510,N_11526);
nand U11916 (N_11916,N_11586,N_11508);
xor U11917 (N_11917,N_11618,N_11477);
or U11918 (N_11918,N_11423,N_11666);
and U11919 (N_11919,N_11422,N_11509);
and U11920 (N_11920,N_11603,N_11475);
xor U11921 (N_11921,N_11499,N_11602);
or U11922 (N_11922,N_11430,N_11691);
xor U11923 (N_11923,N_11434,N_11484);
and U11924 (N_11924,N_11607,N_11495);
nor U11925 (N_11925,N_11651,N_11527);
and U11926 (N_11926,N_11437,N_11608);
nor U11927 (N_11927,N_11513,N_11534);
nand U11928 (N_11928,N_11578,N_11555);
xnor U11929 (N_11929,N_11690,N_11482);
and U11930 (N_11930,N_11660,N_11472);
or U11931 (N_11931,N_11473,N_11490);
and U11932 (N_11932,N_11695,N_11428);
and U11933 (N_11933,N_11463,N_11662);
or U11934 (N_11934,N_11673,N_11622);
and U11935 (N_11935,N_11510,N_11432);
and U11936 (N_11936,N_11447,N_11441);
xnor U11937 (N_11937,N_11655,N_11553);
xnor U11938 (N_11938,N_11537,N_11528);
or U11939 (N_11939,N_11438,N_11511);
nand U11940 (N_11940,N_11459,N_11637);
nor U11941 (N_11941,N_11699,N_11404);
nor U11942 (N_11942,N_11624,N_11438);
nor U11943 (N_11943,N_11427,N_11667);
xnor U11944 (N_11944,N_11621,N_11641);
xnor U11945 (N_11945,N_11656,N_11578);
xnor U11946 (N_11946,N_11652,N_11559);
and U11947 (N_11947,N_11635,N_11680);
nand U11948 (N_11948,N_11632,N_11560);
or U11949 (N_11949,N_11635,N_11575);
or U11950 (N_11950,N_11661,N_11579);
nand U11951 (N_11951,N_11446,N_11523);
nand U11952 (N_11952,N_11636,N_11542);
nor U11953 (N_11953,N_11668,N_11594);
or U11954 (N_11954,N_11607,N_11424);
or U11955 (N_11955,N_11686,N_11462);
nor U11956 (N_11956,N_11524,N_11484);
xnor U11957 (N_11957,N_11408,N_11531);
nand U11958 (N_11958,N_11476,N_11402);
or U11959 (N_11959,N_11607,N_11597);
or U11960 (N_11960,N_11664,N_11458);
xor U11961 (N_11961,N_11527,N_11682);
xor U11962 (N_11962,N_11557,N_11472);
and U11963 (N_11963,N_11615,N_11430);
and U11964 (N_11964,N_11642,N_11658);
nor U11965 (N_11965,N_11628,N_11679);
xnor U11966 (N_11966,N_11411,N_11597);
and U11967 (N_11967,N_11615,N_11654);
or U11968 (N_11968,N_11416,N_11536);
or U11969 (N_11969,N_11632,N_11647);
xnor U11970 (N_11970,N_11628,N_11564);
xnor U11971 (N_11971,N_11457,N_11523);
xor U11972 (N_11972,N_11407,N_11680);
or U11973 (N_11973,N_11471,N_11558);
nand U11974 (N_11974,N_11638,N_11513);
nand U11975 (N_11975,N_11618,N_11487);
and U11976 (N_11976,N_11660,N_11506);
nor U11977 (N_11977,N_11438,N_11608);
and U11978 (N_11978,N_11583,N_11592);
nand U11979 (N_11979,N_11585,N_11487);
or U11980 (N_11980,N_11638,N_11403);
nor U11981 (N_11981,N_11622,N_11670);
nand U11982 (N_11982,N_11670,N_11640);
and U11983 (N_11983,N_11587,N_11488);
nand U11984 (N_11984,N_11513,N_11618);
and U11985 (N_11985,N_11412,N_11698);
and U11986 (N_11986,N_11457,N_11531);
or U11987 (N_11987,N_11597,N_11603);
or U11988 (N_11988,N_11667,N_11497);
nor U11989 (N_11989,N_11482,N_11434);
nor U11990 (N_11990,N_11692,N_11496);
xnor U11991 (N_11991,N_11524,N_11403);
nand U11992 (N_11992,N_11571,N_11532);
or U11993 (N_11993,N_11466,N_11514);
or U11994 (N_11994,N_11487,N_11612);
nor U11995 (N_11995,N_11418,N_11483);
or U11996 (N_11996,N_11500,N_11676);
or U11997 (N_11997,N_11608,N_11520);
and U11998 (N_11998,N_11556,N_11409);
or U11999 (N_11999,N_11624,N_11666);
xnor U12000 (N_12000,N_11726,N_11716);
xnor U12001 (N_12001,N_11825,N_11766);
nor U12002 (N_12002,N_11793,N_11996);
or U12003 (N_12003,N_11924,N_11828);
or U12004 (N_12004,N_11822,N_11772);
nor U12005 (N_12005,N_11783,N_11734);
or U12006 (N_12006,N_11906,N_11775);
or U12007 (N_12007,N_11896,N_11882);
nand U12008 (N_12008,N_11886,N_11839);
or U12009 (N_12009,N_11859,N_11731);
or U12010 (N_12010,N_11984,N_11800);
and U12011 (N_12011,N_11911,N_11959);
nor U12012 (N_12012,N_11894,N_11732);
or U12013 (N_12013,N_11934,N_11874);
and U12014 (N_12014,N_11853,N_11867);
nand U12015 (N_12015,N_11747,N_11788);
nand U12016 (N_12016,N_11933,N_11946);
and U12017 (N_12017,N_11976,N_11918);
or U12018 (N_12018,N_11810,N_11968);
and U12019 (N_12019,N_11965,N_11701);
and U12020 (N_12020,N_11893,N_11851);
or U12021 (N_12021,N_11830,N_11908);
or U12022 (N_12022,N_11870,N_11843);
nor U12023 (N_12023,N_11999,N_11904);
xor U12024 (N_12024,N_11890,N_11944);
or U12025 (N_12025,N_11883,N_11771);
nand U12026 (N_12026,N_11765,N_11948);
and U12027 (N_12027,N_11827,N_11804);
nand U12028 (N_12028,N_11717,N_11989);
and U12029 (N_12029,N_11943,N_11921);
or U12030 (N_12030,N_11888,N_11795);
nor U12031 (N_12031,N_11786,N_11813);
or U12032 (N_12032,N_11901,N_11916);
or U12033 (N_12033,N_11849,N_11834);
xor U12034 (N_12034,N_11977,N_11710);
or U12035 (N_12035,N_11891,N_11768);
nor U12036 (N_12036,N_11983,N_11971);
and U12037 (N_12037,N_11758,N_11845);
or U12038 (N_12038,N_11742,N_11833);
xor U12039 (N_12039,N_11997,N_11872);
or U12040 (N_12040,N_11905,N_11820);
xnor U12041 (N_12041,N_11952,N_11981);
nor U12042 (N_12042,N_11991,N_11869);
xnor U12043 (N_12043,N_11954,N_11803);
or U12044 (N_12044,N_11962,N_11974);
or U12045 (N_12045,N_11955,N_11824);
or U12046 (N_12046,N_11735,N_11702);
or U12047 (N_12047,N_11980,N_11743);
and U12048 (N_12048,N_11727,N_11720);
xnor U12049 (N_12049,N_11718,N_11737);
nand U12050 (N_12050,N_11762,N_11801);
or U12051 (N_12051,N_11829,N_11970);
or U12052 (N_12052,N_11840,N_11945);
nor U12053 (N_12053,N_11812,N_11844);
nand U12054 (N_12054,N_11816,N_11958);
or U12055 (N_12055,N_11887,N_11774);
and U12056 (N_12056,N_11986,N_11837);
and U12057 (N_12057,N_11953,N_11831);
nand U12058 (N_12058,N_11744,N_11846);
xor U12059 (N_12059,N_11998,N_11956);
xor U12060 (N_12060,N_11714,N_11763);
nor U12061 (N_12061,N_11769,N_11926);
or U12062 (N_12062,N_11900,N_11935);
and U12063 (N_12063,N_11794,N_11784);
nand U12064 (N_12064,N_11721,N_11884);
or U12065 (N_12065,N_11733,N_11879);
nand U12066 (N_12066,N_11809,N_11725);
xnor U12067 (N_12067,N_11963,N_11841);
nor U12068 (N_12068,N_11960,N_11730);
or U12069 (N_12069,N_11741,N_11875);
or U12070 (N_12070,N_11988,N_11899);
or U12071 (N_12071,N_11973,N_11876);
or U12072 (N_12072,N_11706,N_11722);
nor U12073 (N_12073,N_11993,N_11947);
nor U12074 (N_12074,N_11920,N_11770);
or U12075 (N_12075,N_11990,N_11847);
and U12076 (N_12076,N_11985,N_11767);
nor U12077 (N_12077,N_11818,N_11740);
and U12078 (N_12078,N_11919,N_11982);
nand U12079 (N_12079,N_11815,N_11719);
xor U12080 (N_12080,N_11950,N_11754);
nor U12081 (N_12081,N_11922,N_11739);
nand U12082 (N_12082,N_11756,N_11755);
or U12083 (N_12083,N_11979,N_11814);
nor U12084 (N_12084,N_11703,N_11909);
xnor U12085 (N_12085,N_11877,N_11798);
or U12086 (N_12086,N_11889,N_11759);
xor U12087 (N_12087,N_11917,N_11892);
xnor U12088 (N_12088,N_11961,N_11778);
nand U12089 (N_12089,N_11995,N_11838);
nand U12090 (N_12090,N_11915,N_11790);
or U12091 (N_12091,N_11942,N_11848);
and U12092 (N_12092,N_11964,N_11861);
xor U12093 (N_12093,N_11880,N_11868);
nor U12094 (N_12094,N_11796,N_11836);
and U12095 (N_12095,N_11802,N_11912);
or U12096 (N_12096,N_11805,N_11826);
nor U12097 (N_12097,N_11745,N_11785);
or U12098 (N_12098,N_11992,N_11808);
xnor U12099 (N_12099,N_11817,N_11819);
nand U12100 (N_12100,N_11797,N_11773);
xor U12101 (N_12101,N_11987,N_11746);
nor U12102 (N_12102,N_11724,N_11878);
nor U12103 (N_12103,N_11782,N_11855);
nor U12104 (N_12104,N_11907,N_11913);
or U12105 (N_12105,N_11707,N_11910);
nand U12106 (N_12106,N_11700,N_11736);
and U12107 (N_12107,N_11821,N_11715);
or U12108 (N_12108,N_11873,N_11871);
nand U12109 (N_12109,N_11711,N_11750);
nor U12110 (N_12110,N_11937,N_11897);
nor U12111 (N_12111,N_11760,N_11856);
or U12112 (N_12112,N_11705,N_11780);
or U12113 (N_12113,N_11864,N_11969);
and U12114 (N_12114,N_11881,N_11748);
and U12115 (N_12115,N_11842,N_11738);
xnor U12116 (N_12116,N_11972,N_11930);
and U12117 (N_12117,N_11753,N_11850);
nor U12118 (N_12118,N_11811,N_11957);
nand U12119 (N_12119,N_11761,N_11923);
xor U12120 (N_12120,N_11975,N_11966);
nor U12121 (N_12121,N_11776,N_11823);
xnor U12122 (N_12122,N_11764,N_11885);
xnor U12123 (N_12123,N_11949,N_11858);
and U12124 (N_12124,N_11863,N_11787);
xor U12125 (N_12125,N_11712,N_11951);
and U12126 (N_12126,N_11807,N_11752);
nand U12127 (N_12127,N_11967,N_11728);
or U12128 (N_12128,N_11940,N_11781);
xnor U12129 (N_12129,N_11854,N_11938);
xor U12130 (N_12130,N_11777,N_11779);
xnor U12131 (N_12131,N_11895,N_11751);
nor U12132 (N_12132,N_11852,N_11925);
nand U12133 (N_12133,N_11931,N_11792);
nand U12134 (N_12134,N_11791,N_11729);
nor U12135 (N_12135,N_11994,N_11723);
or U12136 (N_12136,N_11806,N_11862);
nand U12137 (N_12137,N_11929,N_11939);
and U12138 (N_12138,N_11835,N_11903);
nor U12139 (N_12139,N_11914,N_11941);
and U12140 (N_12140,N_11832,N_11713);
xor U12141 (N_12141,N_11978,N_11866);
nand U12142 (N_12142,N_11865,N_11799);
and U12143 (N_12143,N_11789,N_11932);
or U12144 (N_12144,N_11749,N_11936);
and U12145 (N_12145,N_11927,N_11857);
nand U12146 (N_12146,N_11709,N_11928);
nand U12147 (N_12147,N_11902,N_11708);
nand U12148 (N_12148,N_11704,N_11898);
or U12149 (N_12149,N_11860,N_11757);
nand U12150 (N_12150,N_11774,N_11904);
xnor U12151 (N_12151,N_11904,N_11702);
nand U12152 (N_12152,N_11741,N_11954);
and U12153 (N_12153,N_11949,N_11885);
or U12154 (N_12154,N_11812,N_11840);
and U12155 (N_12155,N_11868,N_11919);
or U12156 (N_12156,N_11835,N_11879);
nand U12157 (N_12157,N_11883,N_11819);
and U12158 (N_12158,N_11735,N_11831);
and U12159 (N_12159,N_11879,N_11823);
and U12160 (N_12160,N_11909,N_11787);
and U12161 (N_12161,N_11882,N_11753);
nand U12162 (N_12162,N_11732,N_11995);
and U12163 (N_12163,N_11761,N_11760);
nor U12164 (N_12164,N_11761,N_11746);
xor U12165 (N_12165,N_11854,N_11742);
and U12166 (N_12166,N_11920,N_11907);
xor U12167 (N_12167,N_11858,N_11954);
or U12168 (N_12168,N_11968,N_11911);
or U12169 (N_12169,N_11883,N_11702);
and U12170 (N_12170,N_11951,N_11718);
or U12171 (N_12171,N_11998,N_11768);
nand U12172 (N_12172,N_11910,N_11825);
nor U12173 (N_12173,N_11907,N_11814);
nor U12174 (N_12174,N_11973,N_11962);
or U12175 (N_12175,N_11966,N_11989);
or U12176 (N_12176,N_11956,N_11794);
nand U12177 (N_12177,N_11877,N_11792);
nand U12178 (N_12178,N_11793,N_11977);
nor U12179 (N_12179,N_11781,N_11812);
or U12180 (N_12180,N_11926,N_11959);
nand U12181 (N_12181,N_11787,N_11886);
and U12182 (N_12182,N_11960,N_11866);
nand U12183 (N_12183,N_11704,N_11908);
nor U12184 (N_12184,N_11701,N_11863);
and U12185 (N_12185,N_11811,N_11788);
or U12186 (N_12186,N_11805,N_11772);
xor U12187 (N_12187,N_11886,N_11749);
or U12188 (N_12188,N_11811,N_11786);
and U12189 (N_12189,N_11973,N_11882);
nor U12190 (N_12190,N_11906,N_11846);
nor U12191 (N_12191,N_11758,N_11715);
nand U12192 (N_12192,N_11734,N_11831);
nand U12193 (N_12193,N_11995,N_11822);
or U12194 (N_12194,N_11843,N_11764);
xor U12195 (N_12195,N_11884,N_11724);
nor U12196 (N_12196,N_11981,N_11960);
xor U12197 (N_12197,N_11802,N_11798);
xnor U12198 (N_12198,N_11730,N_11814);
xor U12199 (N_12199,N_11770,N_11935);
and U12200 (N_12200,N_11964,N_11801);
nand U12201 (N_12201,N_11997,N_11708);
xnor U12202 (N_12202,N_11872,N_11842);
xor U12203 (N_12203,N_11885,N_11977);
nor U12204 (N_12204,N_11760,N_11839);
or U12205 (N_12205,N_11735,N_11749);
or U12206 (N_12206,N_11875,N_11873);
xor U12207 (N_12207,N_11881,N_11795);
nand U12208 (N_12208,N_11719,N_11745);
and U12209 (N_12209,N_11869,N_11875);
nor U12210 (N_12210,N_11978,N_11774);
nand U12211 (N_12211,N_11849,N_11811);
xor U12212 (N_12212,N_11863,N_11947);
nand U12213 (N_12213,N_11889,N_11773);
or U12214 (N_12214,N_11983,N_11774);
or U12215 (N_12215,N_11975,N_11833);
xor U12216 (N_12216,N_11782,N_11734);
and U12217 (N_12217,N_11970,N_11795);
and U12218 (N_12218,N_11829,N_11996);
and U12219 (N_12219,N_11971,N_11942);
nor U12220 (N_12220,N_11804,N_11983);
nand U12221 (N_12221,N_11908,N_11951);
or U12222 (N_12222,N_11874,N_11969);
nor U12223 (N_12223,N_11706,N_11814);
nand U12224 (N_12224,N_11935,N_11918);
xor U12225 (N_12225,N_11751,N_11996);
and U12226 (N_12226,N_11950,N_11919);
and U12227 (N_12227,N_11731,N_11964);
nor U12228 (N_12228,N_11837,N_11940);
or U12229 (N_12229,N_11778,N_11815);
and U12230 (N_12230,N_11823,N_11853);
or U12231 (N_12231,N_11938,N_11817);
and U12232 (N_12232,N_11815,N_11907);
nand U12233 (N_12233,N_11971,N_11956);
xor U12234 (N_12234,N_11815,N_11997);
or U12235 (N_12235,N_11926,N_11965);
nor U12236 (N_12236,N_11727,N_11700);
and U12237 (N_12237,N_11710,N_11805);
nor U12238 (N_12238,N_11987,N_11776);
xnor U12239 (N_12239,N_11799,N_11813);
and U12240 (N_12240,N_11709,N_11734);
or U12241 (N_12241,N_11837,N_11977);
and U12242 (N_12242,N_11864,N_11830);
or U12243 (N_12243,N_11799,N_11887);
nand U12244 (N_12244,N_11779,N_11853);
or U12245 (N_12245,N_11880,N_11902);
xnor U12246 (N_12246,N_11738,N_11824);
nor U12247 (N_12247,N_11703,N_11796);
xnor U12248 (N_12248,N_11767,N_11827);
and U12249 (N_12249,N_11838,N_11991);
xnor U12250 (N_12250,N_11916,N_11928);
nand U12251 (N_12251,N_11836,N_11757);
or U12252 (N_12252,N_11712,N_11763);
and U12253 (N_12253,N_11789,N_11710);
nor U12254 (N_12254,N_11933,N_11899);
and U12255 (N_12255,N_11753,N_11861);
nand U12256 (N_12256,N_11877,N_11701);
nor U12257 (N_12257,N_11851,N_11892);
and U12258 (N_12258,N_11944,N_11963);
or U12259 (N_12259,N_11984,N_11998);
or U12260 (N_12260,N_11812,N_11751);
or U12261 (N_12261,N_11981,N_11950);
xnor U12262 (N_12262,N_11801,N_11884);
nand U12263 (N_12263,N_11983,N_11857);
or U12264 (N_12264,N_11823,N_11726);
nor U12265 (N_12265,N_11767,N_11998);
nor U12266 (N_12266,N_11790,N_11710);
or U12267 (N_12267,N_11720,N_11836);
nand U12268 (N_12268,N_11785,N_11799);
nor U12269 (N_12269,N_11922,N_11988);
or U12270 (N_12270,N_11928,N_11785);
nor U12271 (N_12271,N_11973,N_11927);
and U12272 (N_12272,N_11887,N_11738);
nand U12273 (N_12273,N_11706,N_11784);
or U12274 (N_12274,N_11951,N_11782);
or U12275 (N_12275,N_11844,N_11933);
or U12276 (N_12276,N_11919,N_11803);
xor U12277 (N_12277,N_11747,N_11826);
nand U12278 (N_12278,N_11775,N_11876);
nand U12279 (N_12279,N_11745,N_11784);
and U12280 (N_12280,N_11962,N_11760);
and U12281 (N_12281,N_11711,N_11792);
nand U12282 (N_12282,N_11793,N_11998);
nand U12283 (N_12283,N_11868,N_11872);
or U12284 (N_12284,N_11707,N_11925);
nor U12285 (N_12285,N_11714,N_11995);
and U12286 (N_12286,N_11931,N_11959);
nand U12287 (N_12287,N_11765,N_11855);
or U12288 (N_12288,N_11962,N_11964);
nand U12289 (N_12289,N_11993,N_11844);
nor U12290 (N_12290,N_11708,N_11744);
nand U12291 (N_12291,N_11914,N_11797);
nor U12292 (N_12292,N_11995,N_11992);
nor U12293 (N_12293,N_11824,N_11757);
and U12294 (N_12294,N_11926,N_11885);
xnor U12295 (N_12295,N_11902,N_11933);
nand U12296 (N_12296,N_11834,N_11739);
and U12297 (N_12297,N_11920,N_11761);
xnor U12298 (N_12298,N_11778,N_11998);
and U12299 (N_12299,N_11998,N_11899);
or U12300 (N_12300,N_12269,N_12247);
xor U12301 (N_12301,N_12010,N_12046);
xor U12302 (N_12302,N_12198,N_12196);
and U12303 (N_12303,N_12187,N_12284);
and U12304 (N_12304,N_12185,N_12231);
or U12305 (N_12305,N_12176,N_12076);
nand U12306 (N_12306,N_12286,N_12077);
nor U12307 (N_12307,N_12033,N_12193);
nand U12308 (N_12308,N_12096,N_12294);
nor U12309 (N_12309,N_12028,N_12057);
nand U12310 (N_12310,N_12162,N_12233);
and U12311 (N_12311,N_12019,N_12156);
and U12312 (N_12312,N_12045,N_12293);
nand U12313 (N_12313,N_12047,N_12107);
nand U12314 (N_12314,N_12152,N_12189);
nor U12315 (N_12315,N_12201,N_12038);
or U12316 (N_12316,N_12035,N_12098);
and U12317 (N_12317,N_12005,N_12166);
nand U12318 (N_12318,N_12295,N_12190);
and U12319 (N_12319,N_12216,N_12148);
nand U12320 (N_12320,N_12053,N_12296);
nand U12321 (N_12321,N_12275,N_12072);
nor U12322 (N_12322,N_12195,N_12060);
and U12323 (N_12323,N_12088,N_12089);
and U12324 (N_12324,N_12272,N_12168);
and U12325 (N_12325,N_12288,N_12122);
nand U12326 (N_12326,N_12257,N_12281);
nor U12327 (N_12327,N_12297,N_12174);
and U12328 (N_12328,N_12075,N_12209);
nor U12329 (N_12329,N_12215,N_12058);
xor U12330 (N_12330,N_12299,N_12007);
and U12331 (N_12331,N_12267,N_12291);
or U12332 (N_12332,N_12027,N_12192);
and U12333 (N_12333,N_12066,N_12106);
nor U12334 (N_12334,N_12167,N_12221);
xor U12335 (N_12335,N_12102,N_12108);
nor U12336 (N_12336,N_12163,N_12188);
nand U12337 (N_12337,N_12214,N_12292);
nor U12338 (N_12338,N_12055,N_12043);
nand U12339 (N_12339,N_12243,N_12091);
and U12340 (N_12340,N_12094,N_12262);
nand U12341 (N_12341,N_12130,N_12071);
xnor U12342 (N_12342,N_12219,N_12224);
and U12343 (N_12343,N_12242,N_12186);
and U12344 (N_12344,N_12199,N_12173);
nand U12345 (N_12345,N_12085,N_12001);
nor U12346 (N_12346,N_12223,N_12121);
nor U12347 (N_12347,N_12081,N_12036);
nand U12348 (N_12348,N_12137,N_12184);
xnor U12349 (N_12349,N_12205,N_12273);
nor U12350 (N_12350,N_12064,N_12105);
nand U12351 (N_12351,N_12109,N_12136);
nor U12352 (N_12352,N_12128,N_12025);
and U12353 (N_12353,N_12236,N_12276);
or U12354 (N_12354,N_12070,N_12112);
or U12355 (N_12355,N_12041,N_12030);
nor U12356 (N_12356,N_12145,N_12155);
nand U12357 (N_12357,N_12124,N_12208);
nor U12358 (N_12358,N_12274,N_12238);
nor U12359 (N_12359,N_12023,N_12253);
or U12360 (N_12360,N_12283,N_12012);
and U12361 (N_12361,N_12256,N_12259);
xor U12362 (N_12362,N_12252,N_12159);
or U12363 (N_12363,N_12087,N_12200);
nor U12364 (N_12364,N_12228,N_12029);
nor U12365 (N_12365,N_12034,N_12170);
nor U12366 (N_12366,N_12031,N_12289);
nor U12367 (N_12367,N_12138,N_12080);
nand U12368 (N_12368,N_12153,N_12049);
and U12369 (N_12369,N_12054,N_12132);
xnor U12370 (N_12370,N_12048,N_12181);
or U12371 (N_12371,N_12197,N_12013);
xnor U12372 (N_12372,N_12052,N_12022);
nand U12373 (N_12373,N_12270,N_12002);
and U12374 (N_12374,N_12059,N_12182);
xnor U12375 (N_12375,N_12011,N_12093);
xnor U12376 (N_12376,N_12250,N_12149);
and U12377 (N_12377,N_12282,N_12073);
nand U12378 (N_12378,N_12245,N_12063);
xnor U12379 (N_12379,N_12298,N_12164);
or U12380 (N_12380,N_12069,N_12082);
and U12381 (N_12381,N_12266,N_12241);
nor U12382 (N_12382,N_12175,N_12123);
xor U12383 (N_12383,N_12264,N_12056);
or U12384 (N_12384,N_12101,N_12251);
xnor U12385 (N_12385,N_12024,N_12229);
and U12386 (N_12386,N_12120,N_12183);
nor U12387 (N_12387,N_12204,N_12000);
and U12388 (N_12388,N_12116,N_12239);
nor U12389 (N_12389,N_12006,N_12095);
nand U12390 (N_12390,N_12240,N_12017);
xnor U12391 (N_12391,N_12171,N_12014);
or U12392 (N_12392,N_12249,N_12146);
nor U12393 (N_12393,N_12147,N_12263);
nor U12394 (N_12394,N_12232,N_12004);
and U12395 (N_12395,N_12255,N_12258);
nand U12396 (N_12396,N_12131,N_12268);
and U12397 (N_12397,N_12218,N_12074);
xnor U12398 (N_12398,N_12261,N_12110);
or U12399 (N_12399,N_12018,N_12078);
nor U12400 (N_12400,N_12244,N_12003);
xnor U12401 (N_12401,N_12154,N_12139);
nor U12402 (N_12402,N_12279,N_12026);
and U12403 (N_12403,N_12118,N_12160);
nor U12404 (N_12404,N_12061,N_12037);
nand U12405 (N_12405,N_12203,N_12086);
nand U12406 (N_12406,N_12158,N_12092);
and U12407 (N_12407,N_12117,N_12119);
or U12408 (N_12408,N_12265,N_12206);
or U12409 (N_12409,N_12210,N_12125);
nand U12410 (N_12410,N_12285,N_12126);
nor U12411 (N_12411,N_12039,N_12212);
nand U12412 (N_12412,N_12127,N_12194);
and U12413 (N_12413,N_12235,N_12227);
nand U12414 (N_12414,N_12234,N_12226);
nor U12415 (N_12415,N_12172,N_12178);
xnor U12416 (N_12416,N_12083,N_12062);
nand U12417 (N_12417,N_12044,N_12260);
or U12418 (N_12418,N_12129,N_12015);
or U12419 (N_12419,N_12157,N_12222);
and U12420 (N_12420,N_12230,N_12179);
or U12421 (N_12421,N_12051,N_12050);
nand U12422 (N_12422,N_12220,N_12151);
nor U12423 (N_12423,N_12271,N_12180);
or U12424 (N_12424,N_12020,N_12114);
nand U12425 (N_12425,N_12165,N_12290);
xor U12426 (N_12426,N_12211,N_12090);
or U12427 (N_12427,N_12191,N_12115);
nor U12428 (N_12428,N_12150,N_12142);
xnor U12429 (N_12429,N_12040,N_12237);
nand U12430 (N_12430,N_12287,N_12248);
and U12431 (N_12431,N_12217,N_12097);
nor U12432 (N_12432,N_12104,N_12135);
nor U12433 (N_12433,N_12140,N_12111);
and U12434 (N_12434,N_12068,N_12207);
nor U12435 (N_12435,N_12067,N_12213);
nor U12436 (N_12436,N_12016,N_12009);
and U12437 (N_12437,N_12161,N_12177);
and U12438 (N_12438,N_12277,N_12133);
xor U12439 (N_12439,N_12079,N_12246);
and U12440 (N_12440,N_12278,N_12100);
nand U12441 (N_12441,N_12099,N_12254);
nand U12442 (N_12442,N_12169,N_12202);
xor U12443 (N_12443,N_12113,N_12008);
nor U12444 (N_12444,N_12134,N_12144);
and U12445 (N_12445,N_12103,N_12042);
nor U12446 (N_12446,N_12032,N_12141);
nor U12447 (N_12447,N_12021,N_12084);
or U12448 (N_12448,N_12225,N_12280);
nand U12449 (N_12449,N_12065,N_12143);
nor U12450 (N_12450,N_12230,N_12280);
xor U12451 (N_12451,N_12058,N_12227);
and U12452 (N_12452,N_12290,N_12073);
nand U12453 (N_12453,N_12085,N_12184);
and U12454 (N_12454,N_12008,N_12137);
xor U12455 (N_12455,N_12280,N_12213);
nand U12456 (N_12456,N_12294,N_12265);
nor U12457 (N_12457,N_12275,N_12225);
or U12458 (N_12458,N_12073,N_12208);
xnor U12459 (N_12459,N_12076,N_12217);
nand U12460 (N_12460,N_12190,N_12041);
nand U12461 (N_12461,N_12194,N_12061);
nand U12462 (N_12462,N_12006,N_12179);
nand U12463 (N_12463,N_12208,N_12252);
and U12464 (N_12464,N_12238,N_12000);
nor U12465 (N_12465,N_12035,N_12178);
nand U12466 (N_12466,N_12029,N_12247);
nand U12467 (N_12467,N_12298,N_12203);
nor U12468 (N_12468,N_12297,N_12256);
or U12469 (N_12469,N_12111,N_12282);
xor U12470 (N_12470,N_12033,N_12127);
or U12471 (N_12471,N_12069,N_12269);
or U12472 (N_12472,N_12175,N_12127);
xnor U12473 (N_12473,N_12015,N_12252);
or U12474 (N_12474,N_12230,N_12058);
xnor U12475 (N_12475,N_12290,N_12199);
and U12476 (N_12476,N_12159,N_12099);
nor U12477 (N_12477,N_12064,N_12043);
xnor U12478 (N_12478,N_12200,N_12132);
or U12479 (N_12479,N_12032,N_12207);
nand U12480 (N_12480,N_12033,N_12017);
nand U12481 (N_12481,N_12262,N_12026);
nor U12482 (N_12482,N_12154,N_12013);
and U12483 (N_12483,N_12074,N_12140);
xnor U12484 (N_12484,N_12044,N_12134);
and U12485 (N_12485,N_12114,N_12130);
nand U12486 (N_12486,N_12215,N_12137);
nand U12487 (N_12487,N_12243,N_12147);
or U12488 (N_12488,N_12250,N_12068);
nor U12489 (N_12489,N_12054,N_12150);
or U12490 (N_12490,N_12245,N_12260);
nand U12491 (N_12491,N_12216,N_12049);
nand U12492 (N_12492,N_12118,N_12006);
and U12493 (N_12493,N_12219,N_12129);
nor U12494 (N_12494,N_12022,N_12102);
nor U12495 (N_12495,N_12127,N_12139);
nor U12496 (N_12496,N_12208,N_12111);
xnor U12497 (N_12497,N_12054,N_12196);
nor U12498 (N_12498,N_12055,N_12235);
or U12499 (N_12499,N_12259,N_12029);
xnor U12500 (N_12500,N_12125,N_12002);
nand U12501 (N_12501,N_12000,N_12247);
nand U12502 (N_12502,N_12234,N_12290);
nor U12503 (N_12503,N_12205,N_12298);
and U12504 (N_12504,N_12220,N_12033);
nand U12505 (N_12505,N_12081,N_12064);
or U12506 (N_12506,N_12277,N_12165);
nor U12507 (N_12507,N_12029,N_12025);
nor U12508 (N_12508,N_12051,N_12276);
nand U12509 (N_12509,N_12019,N_12070);
and U12510 (N_12510,N_12192,N_12254);
nor U12511 (N_12511,N_12104,N_12113);
or U12512 (N_12512,N_12043,N_12049);
and U12513 (N_12513,N_12188,N_12003);
or U12514 (N_12514,N_12102,N_12030);
nor U12515 (N_12515,N_12097,N_12285);
nand U12516 (N_12516,N_12165,N_12053);
nand U12517 (N_12517,N_12283,N_12180);
or U12518 (N_12518,N_12226,N_12169);
nand U12519 (N_12519,N_12155,N_12142);
nor U12520 (N_12520,N_12297,N_12000);
or U12521 (N_12521,N_12023,N_12085);
nand U12522 (N_12522,N_12139,N_12193);
or U12523 (N_12523,N_12142,N_12031);
or U12524 (N_12524,N_12146,N_12052);
or U12525 (N_12525,N_12273,N_12036);
xnor U12526 (N_12526,N_12232,N_12211);
and U12527 (N_12527,N_12163,N_12089);
and U12528 (N_12528,N_12025,N_12148);
or U12529 (N_12529,N_12195,N_12014);
nand U12530 (N_12530,N_12185,N_12299);
xnor U12531 (N_12531,N_12069,N_12257);
or U12532 (N_12532,N_12155,N_12191);
and U12533 (N_12533,N_12088,N_12078);
xor U12534 (N_12534,N_12243,N_12157);
and U12535 (N_12535,N_12260,N_12086);
nand U12536 (N_12536,N_12106,N_12017);
nor U12537 (N_12537,N_12127,N_12256);
or U12538 (N_12538,N_12190,N_12081);
nor U12539 (N_12539,N_12234,N_12062);
nor U12540 (N_12540,N_12151,N_12021);
nor U12541 (N_12541,N_12260,N_12232);
or U12542 (N_12542,N_12149,N_12044);
xnor U12543 (N_12543,N_12096,N_12251);
or U12544 (N_12544,N_12001,N_12057);
nor U12545 (N_12545,N_12173,N_12045);
and U12546 (N_12546,N_12140,N_12170);
or U12547 (N_12547,N_12284,N_12209);
nor U12548 (N_12548,N_12283,N_12005);
nor U12549 (N_12549,N_12291,N_12283);
nor U12550 (N_12550,N_12088,N_12017);
xnor U12551 (N_12551,N_12278,N_12272);
xnor U12552 (N_12552,N_12193,N_12223);
nor U12553 (N_12553,N_12087,N_12227);
nor U12554 (N_12554,N_12226,N_12105);
nor U12555 (N_12555,N_12077,N_12140);
or U12556 (N_12556,N_12119,N_12049);
and U12557 (N_12557,N_12034,N_12105);
nor U12558 (N_12558,N_12124,N_12244);
xnor U12559 (N_12559,N_12030,N_12157);
or U12560 (N_12560,N_12248,N_12195);
nor U12561 (N_12561,N_12138,N_12173);
or U12562 (N_12562,N_12017,N_12210);
nand U12563 (N_12563,N_12066,N_12127);
and U12564 (N_12564,N_12077,N_12166);
and U12565 (N_12565,N_12286,N_12248);
xnor U12566 (N_12566,N_12138,N_12090);
nand U12567 (N_12567,N_12016,N_12012);
nor U12568 (N_12568,N_12254,N_12047);
xor U12569 (N_12569,N_12063,N_12285);
xor U12570 (N_12570,N_12207,N_12181);
or U12571 (N_12571,N_12053,N_12275);
or U12572 (N_12572,N_12079,N_12217);
and U12573 (N_12573,N_12142,N_12168);
xnor U12574 (N_12574,N_12168,N_12174);
or U12575 (N_12575,N_12209,N_12119);
nor U12576 (N_12576,N_12015,N_12018);
nand U12577 (N_12577,N_12164,N_12077);
and U12578 (N_12578,N_12139,N_12064);
nand U12579 (N_12579,N_12038,N_12118);
and U12580 (N_12580,N_12011,N_12281);
or U12581 (N_12581,N_12255,N_12058);
and U12582 (N_12582,N_12277,N_12251);
xor U12583 (N_12583,N_12160,N_12121);
xnor U12584 (N_12584,N_12207,N_12249);
or U12585 (N_12585,N_12104,N_12166);
nand U12586 (N_12586,N_12100,N_12010);
xnor U12587 (N_12587,N_12156,N_12119);
nor U12588 (N_12588,N_12208,N_12278);
nor U12589 (N_12589,N_12118,N_12232);
or U12590 (N_12590,N_12296,N_12045);
nor U12591 (N_12591,N_12153,N_12164);
xor U12592 (N_12592,N_12209,N_12226);
nor U12593 (N_12593,N_12034,N_12126);
nand U12594 (N_12594,N_12161,N_12024);
xnor U12595 (N_12595,N_12249,N_12104);
xnor U12596 (N_12596,N_12280,N_12021);
nand U12597 (N_12597,N_12170,N_12158);
xor U12598 (N_12598,N_12113,N_12052);
nand U12599 (N_12599,N_12186,N_12080);
and U12600 (N_12600,N_12312,N_12594);
nor U12601 (N_12601,N_12472,N_12593);
xnor U12602 (N_12602,N_12452,N_12556);
xnor U12603 (N_12603,N_12513,N_12359);
xor U12604 (N_12604,N_12474,N_12326);
or U12605 (N_12605,N_12431,N_12532);
nand U12606 (N_12606,N_12500,N_12381);
xnor U12607 (N_12607,N_12367,N_12342);
or U12608 (N_12608,N_12562,N_12555);
or U12609 (N_12609,N_12416,N_12357);
nor U12610 (N_12610,N_12337,N_12522);
xor U12611 (N_12611,N_12393,N_12305);
xor U12612 (N_12612,N_12458,N_12551);
and U12613 (N_12613,N_12443,N_12535);
nand U12614 (N_12614,N_12315,N_12485);
xnor U12615 (N_12615,N_12384,N_12577);
nor U12616 (N_12616,N_12368,N_12507);
nor U12617 (N_12617,N_12456,N_12449);
or U12618 (N_12618,N_12347,N_12308);
nand U12619 (N_12619,N_12564,N_12586);
and U12620 (N_12620,N_12599,N_12523);
and U12621 (N_12621,N_12461,N_12520);
nor U12622 (N_12622,N_12478,N_12477);
xnor U12623 (N_12623,N_12476,N_12467);
or U12624 (N_12624,N_12543,N_12386);
or U12625 (N_12625,N_12496,N_12493);
nand U12626 (N_12626,N_12366,N_12375);
and U12627 (N_12627,N_12313,N_12530);
nor U12628 (N_12628,N_12329,N_12425);
nand U12629 (N_12629,N_12408,N_12322);
nand U12630 (N_12630,N_12440,N_12480);
xor U12631 (N_12631,N_12350,N_12399);
and U12632 (N_12632,N_12438,N_12587);
xor U12633 (N_12633,N_12544,N_12519);
nor U12634 (N_12634,N_12435,N_12418);
nand U12635 (N_12635,N_12469,N_12388);
nand U12636 (N_12636,N_12572,N_12489);
or U12637 (N_12637,N_12411,N_12539);
or U12638 (N_12638,N_12383,N_12509);
or U12639 (N_12639,N_12592,N_12373);
and U12640 (N_12640,N_12470,N_12573);
nand U12641 (N_12641,N_12571,N_12332);
xnor U12642 (N_12642,N_12482,N_12394);
and U12643 (N_12643,N_12429,N_12508);
and U12644 (N_12644,N_12575,N_12553);
or U12645 (N_12645,N_12494,N_12569);
and U12646 (N_12646,N_12439,N_12389);
nand U12647 (N_12647,N_12473,N_12579);
or U12648 (N_12648,N_12321,N_12475);
and U12649 (N_12649,N_12317,N_12304);
nor U12650 (N_12650,N_12323,N_12406);
xnor U12651 (N_12651,N_12537,N_12340);
nand U12652 (N_12652,N_12549,N_12430);
or U12653 (N_12653,N_12385,N_12465);
nand U12654 (N_12654,N_12392,N_12427);
or U12655 (N_12655,N_12504,N_12395);
or U12656 (N_12656,N_12344,N_12306);
xor U12657 (N_12657,N_12526,N_12397);
nand U12658 (N_12658,N_12525,N_12311);
xnor U12659 (N_12659,N_12349,N_12542);
nand U12660 (N_12660,N_12457,N_12582);
xor U12661 (N_12661,N_12568,N_12314);
xor U12662 (N_12662,N_12303,N_12309);
nor U12663 (N_12663,N_12316,N_12421);
nand U12664 (N_12664,N_12591,N_12341);
or U12665 (N_12665,N_12595,N_12527);
xnor U12666 (N_12666,N_12391,N_12518);
nand U12667 (N_12667,N_12302,N_12414);
nand U12668 (N_12668,N_12514,N_12361);
nand U12669 (N_12669,N_12576,N_12567);
and U12670 (N_12670,N_12371,N_12446);
or U12671 (N_12671,N_12468,N_12370);
or U12672 (N_12672,N_12566,N_12335);
or U12673 (N_12673,N_12528,N_12462);
and U12674 (N_12674,N_12409,N_12426);
nor U12675 (N_12675,N_12331,N_12501);
or U12676 (N_12676,N_12401,N_12464);
nand U12677 (N_12677,N_12454,N_12346);
nand U12678 (N_12678,N_12531,N_12538);
or U12679 (N_12679,N_12505,N_12471);
nor U12680 (N_12680,N_12547,N_12415);
and U12681 (N_12681,N_12506,N_12512);
nand U12682 (N_12682,N_12307,N_12407);
and U12683 (N_12683,N_12517,N_12387);
xnor U12684 (N_12684,N_12445,N_12382);
and U12685 (N_12685,N_12398,N_12453);
or U12686 (N_12686,N_12534,N_12374);
and U12687 (N_12687,N_12590,N_12378);
nand U12688 (N_12688,N_12369,N_12360);
nand U12689 (N_12689,N_12447,N_12495);
nand U12690 (N_12690,N_12460,N_12580);
or U12691 (N_12691,N_12403,N_12348);
nand U12692 (N_12692,N_12405,N_12424);
xnor U12693 (N_12693,N_12301,N_12380);
or U12694 (N_12694,N_12338,N_12583);
or U12695 (N_12695,N_12363,N_12351);
xor U12696 (N_12696,N_12423,N_12432);
xor U12697 (N_12697,N_12428,N_12442);
nand U12698 (N_12698,N_12585,N_12441);
xnor U12699 (N_12699,N_12310,N_12356);
xnor U12700 (N_12700,N_12319,N_12434);
nor U12701 (N_12701,N_12444,N_12487);
nand U12702 (N_12702,N_12481,N_12596);
xor U12703 (N_12703,N_12565,N_12516);
and U12704 (N_12704,N_12362,N_12437);
or U12705 (N_12705,N_12358,N_12546);
and U12706 (N_12706,N_12396,N_12578);
or U12707 (N_12707,N_12490,N_12327);
and U12708 (N_12708,N_12492,N_12379);
and U12709 (N_12709,N_12376,N_12559);
nor U12710 (N_12710,N_12355,N_12339);
and U12711 (N_12711,N_12560,N_12545);
nor U12712 (N_12712,N_12488,N_12497);
nand U12713 (N_12713,N_12536,N_12533);
nor U12714 (N_12714,N_12524,N_12354);
xnor U12715 (N_12715,N_12510,N_12515);
nand U12716 (N_12716,N_12402,N_12330);
nand U12717 (N_12717,N_12541,N_12597);
nand U12718 (N_12718,N_12540,N_12324);
or U12719 (N_12719,N_12436,N_12498);
nor U12720 (N_12720,N_12588,N_12410);
and U12721 (N_12721,N_12413,N_12353);
nor U12722 (N_12722,N_12557,N_12372);
nand U12723 (N_12723,N_12502,N_12420);
or U12724 (N_12724,N_12459,N_12365);
and U12725 (N_12725,N_12364,N_12328);
nor U12726 (N_12726,N_12550,N_12521);
nand U12727 (N_12727,N_12336,N_12334);
and U12728 (N_12728,N_12503,N_12529);
nor U12729 (N_12729,N_12491,N_12552);
xor U12730 (N_12730,N_12352,N_12433);
xor U12731 (N_12731,N_12318,N_12343);
nor U12732 (N_12732,N_12466,N_12511);
xor U12733 (N_12733,N_12450,N_12561);
nor U12734 (N_12734,N_12554,N_12479);
or U12735 (N_12735,N_12448,N_12558);
or U12736 (N_12736,N_12486,N_12417);
xor U12737 (N_12737,N_12570,N_12581);
or U12738 (N_12738,N_12377,N_12484);
xnor U12739 (N_12739,N_12325,N_12404);
xnor U12740 (N_12740,N_12563,N_12574);
nor U12741 (N_12741,N_12584,N_12483);
or U12742 (N_12742,N_12548,N_12455);
nand U12743 (N_12743,N_12463,N_12598);
or U12744 (N_12744,N_12419,N_12589);
or U12745 (N_12745,N_12412,N_12320);
nand U12746 (N_12746,N_12333,N_12400);
and U12747 (N_12747,N_12345,N_12300);
nor U12748 (N_12748,N_12390,N_12499);
or U12749 (N_12749,N_12422,N_12451);
and U12750 (N_12750,N_12469,N_12428);
or U12751 (N_12751,N_12479,N_12541);
nor U12752 (N_12752,N_12330,N_12315);
xnor U12753 (N_12753,N_12582,N_12362);
nor U12754 (N_12754,N_12556,N_12525);
nand U12755 (N_12755,N_12305,N_12445);
xnor U12756 (N_12756,N_12538,N_12342);
nor U12757 (N_12757,N_12310,N_12437);
nor U12758 (N_12758,N_12588,N_12532);
nor U12759 (N_12759,N_12338,N_12429);
and U12760 (N_12760,N_12503,N_12313);
xnor U12761 (N_12761,N_12545,N_12567);
or U12762 (N_12762,N_12456,N_12576);
nor U12763 (N_12763,N_12412,N_12495);
nand U12764 (N_12764,N_12366,N_12565);
xor U12765 (N_12765,N_12345,N_12515);
xnor U12766 (N_12766,N_12368,N_12560);
or U12767 (N_12767,N_12495,N_12549);
or U12768 (N_12768,N_12408,N_12467);
and U12769 (N_12769,N_12401,N_12393);
nand U12770 (N_12770,N_12464,N_12414);
nand U12771 (N_12771,N_12500,N_12397);
xor U12772 (N_12772,N_12375,N_12372);
or U12773 (N_12773,N_12515,N_12383);
nor U12774 (N_12774,N_12332,N_12390);
or U12775 (N_12775,N_12429,N_12348);
and U12776 (N_12776,N_12470,N_12545);
and U12777 (N_12777,N_12476,N_12460);
and U12778 (N_12778,N_12342,N_12505);
and U12779 (N_12779,N_12483,N_12324);
and U12780 (N_12780,N_12549,N_12581);
nor U12781 (N_12781,N_12580,N_12367);
or U12782 (N_12782,N_12382,N_12467);
and U12783 (N_12783,N_12366,N_12339);
nor U12784 (N_12784,N_12576,N_12450);
nand U12785 (N_12785,N_12359,N_12562);
and U12786 (N_12786,N_12316,N_12537);
nand U12787 (N_12787,N_12336,N_12341);
nor U12788 (N_12788,N_12506,N_12398);
and U12789 (N_12789,N_12319,N_12471);
nand U12790 (N_12790,N_12405,N_12406);
and U12791 (N_12791,N_12537,N_12592);
xnor U12792 (N_12792,N_12397,N_12543);
nor U12793 (N_12793,N_12510,N_12409);
xnor U12794 (N_12794,N_12339,N_12526);
nor U12795 (N_12795,N_12546,N_12564);
xnor U12796 (N_12796,N_12472,N_12546);
and U12797 (N_12797,N_12544,N_12330);
or U12798 (N_12798,N_12517,N_12441);
or U12799 (N_12799,N_12376,N_12379);
nand U12800 (N_12800,N_12597,N_12434);
nor U12801 (N_12801,N_12521,N_12398);
nand U12802 (N_12802,N_12398,N_12321);
nand U12803 (N_12803,N_12582,N_12548);
xnor U12804 (N_12804,N_12309,N_12321);
or U12805 (N_12805,N_12563,N_12589);
nor U12806 (N_12806,N_12492,N_12502);
xor U12807 (N_12807,N_12361,N_12500);
and U12808 (N_12808,N_12460,N_12330);
nand U12809 (N_12809,N_12493,N_12427);
nand U12810 (N_12810,N_12401,N_12375);
and U12811 (N_12811,N_12337,N_12472);
nand U12812 (N_12812,N_12578,N_12364);
and U12813 (N_12813,N_12512,N_12494);
nand U12814 (N_12814,N_12533,N_12412);
xnor U12815 (N_12815,N_12361,N_12596);
or U12816 (N_12816,N_12482,N_12441);
nor U12817 (N_12817,N_12442,N_12382);
or U12818 (N_12818,N_12533,N_12383);
xnor U12819 (N_12819,N_12593,N_12328);
nand U12820 (N_12820,N_12372,N_12436);
nor U12821 (N_12821,N_12397,N_12394);
or U12822 (N_12822,N_12480,N_12428);
or U12823 (N_12823,N_12380,N_12389);
nor U12824 (N_12824,N_12599,N_12311);
xor U12825 (N_12825,N_12555,N_12522);
xnor U12826 (N_12826,N_12449,N_12426);
xnor U12827 (N_12827,N_12339,N_12590);
nor U12828 (N_12828,N_12547,N_12476);
nor U12829 (N_12829,N_12352,N_12378);
nor U12830 (N_12830,N_12573,N_12563);
nor U12831 (N_12831,N_12533,N_12508);
and U12832 (N_12832,N_12587,N_12324);
or U12833 (N_12833,N_12498,N_12454);
nor U12834 (N_12834,N_12550,N_12576);
nand U12835 (N_12835,N_12336,N_12464);
or U12836 (N_12836,N_12527,N_12375);
nor U12837 (N_12837,N_12421,N_12512);
xnor U12838 (N_12838,N_12544,N_12443);
xor U12839 (N_12839,N_12405,N_12378);
xor U12840 (N_12840,N_12312,N_12495);
nor U12841 (N_12841,N_12576,N_12414);
and U12842 (N_12842,N_12437,N_12520);
xnor U12843 (N_12843,N_12381,N_12539);
and U12844 (N_12844,N_12540,N_12579);
or U12845 (N_12845,N_12379,N_12338);
nor U12846 (N_12846,N_12381,N_12482);
and U12847 (N_12847,N_12499,N_12431);
or U12848 (N_12848,N_12586,N_12437);
and U12849 (N_12849,N_12386,N_12455);
nand U12850 (N_12850,N_12496,N_12476);
and U12851 (N_12851,N_12486,N_12445);
nand U12852 (N_12852,N_12535,N_12325);
xnor U12853 (N_12853,N_12496,N_12311);
nor U12854 (N_12854,N_12416,N_12454);
and U12855 (N_12855,N_12517,N_12371);
and U12856 (N_12856,N_12381,N_12343);
xor U12857 (N_12857,N_12427,N_12576);
nor U12858 (N_12858,N_12464,N_12303);
nand U12859 (N_12859,N_12420,N_12553);
xnor U12860 (N_12860,N_12484,N_12499);
or U12861 (N_12861,N_12331,N_12570);
and U12862 (N_12862,N_12353,N_12331);
xor U12863 (N_12863,N_12535,N_12314);
nand U12864 (N_12864,N_12385,N_12448);
or U12865 (N_12865,N_12486,N_12437);
nor U12866 (N_12866,N_12342,N_12369);
nor U12867 (N_12867,N_12576,N_12494);
nor U12868 (N_12868,N_12444,N_12415);
nand U12869 (N_12869,N_12583,N_12430);
xnor U12870 (N_12870,N_12365,N_12349);
nor U12871 (N_12871,N_12596,N_12418);
nand U12872 (N_12872,N_12433,N_12310);
and U12873 (N_12873,N_12436,N_12392);
and U12874 (N_12874,N_12349,N_12433);
nor U12875 (N_12875,N_12532,N_12339);
nor U12876 (N_12876,N_12492,N_12315);
and U12877 (N_12877,N_12545,N_12425);
nor U12878 (N_12878,N_12500,N_12591);
or U12879 (N_12879,N_12466,N_12425);
nor U12880 (N_12880,N_12562,N_12490);
and U12881 (N_12881,N_12575,N_12548);
and U12882 (N_12882,N_12405,N_12527);
and U12883 (N_12883,N_12467,N_12478);
xor U12884 (N_12884,N_12524,N_12313);
xnor U12885 (N_12885,N_12440,N_12525);
xnor U12886 (N_12886,N_12353,N_12474);
and U12887 (N_12887,N_12377,N_12326);
xor U12888 (N_12888,N_12377,N_12330);
xnor U12889 (N_12889,N_12446,N_12309);
xor U12890 (N_12890,N_12548,N_12597);
nor U12891 (N_12891,N_12395,N_12383);
nand U12892 (N_12892,N_12559,N_12340);
and U12893 (N_12893,N_12340,N_12510);
or U12894 (N_12894,N_12313,N_12572);
or U12895 (N_12895,N_12415,N_12383);
nand U12896 (N_12896,N_12451,N_12587);
or U12897 (N_12897,N_12455,N_12576);
xor U12898 (N_12898,N_12460,N_12457);
or U12899 (N_12899,N_12446,N_12364);
or U12900 (N_12900,N_12685,N_12871);
nor U12901 (N_12901,N_12804,N_12707);
or U12902 (N_12902,N_12606,N_12805);
nor U12903 (N_12903,N_12786,N_12723);
and U12904 (N_12904,N_12653,N_12852);
nor U12905 (N_12905,N_12674,N_12722);
or U12906 (N_12906,N_12779,N_12890);
xnor U12907 (N_12907,N_12845,N_12781);
xnor U12908 (N_12908,N_12615,N_12818);
or U12909 (N_12909,N_12618,N_12761);
nand U12910 (N_12910,N_12635,N_12894);
nor U12911 (N_12911,N_12687,N_12816);
nand U12912 (N_12912,N_12851,N_12616);
nand U12913 (N_12913,N_12870,N_12646);
xor U12914 (N_12914,N_12600,N_12771);
nand U12915 (N_12915,N_12637,N_12648);
nand U12916 (N_12916,N_12746,N_12613);
and U12917 (N_12917,N_12630,N_12706);
nor U12918 (N_12918,N_12895,N_12623);
and U12919 (N_12919,N_12838,N_12847);
or U12920 (N_12920,N_12881,N_12673);
or U12921 (N_12921,N_12607,N_12828);
or U12922 (N_12922,N_12885,N_12820);
nand U12923 (N_12923,N_12645,N_12874);
or U12924 (N_12924,N_12693,N_12799);
or U12925 (N_12925,N_12656,N_12831);
nand U12926 (N_12926,N_12750,N_12736);
nor U12927 (N_12927,N_12756,N_12832);
xor U12928 (N_12928,N_12833,N_12728);
nor U12929 (N_12929,N_12760,N_12768);
and U12930 (N_12930,N_12751,N_12605);
xor U12931 (N_12931,N_12788,N_12879);
nor U12932 (N_12932,N_12810,N_12720);
nor U12933 (N_12933,N_12749,N_12752);
and U12934 (N_12934,N_12797,N_12603);
xnor U12935 (N_12935,N_12711,N_12865);
xor U12936 (N_12936,N_12780,N_12848);
nand U12937 (N_12937,N_12774,N_12855);
xnor U12938 (N_12938,N_12626,N_12856);
nand U12939 (N_12939,N_12854,N_12725);
and U12940 (N_12940,N_12697,N_12633);
xor U12941 (N_12941,N_12712,N_12665);
or U12942 (N_12942,N_12628,N_12873);
nor U12943 (N_12943,N_12664,N_12688);
and U12944 (N_12944,N_12708,N_12668);
or U12945 (N_12945,N_12709,N_12770);
and U12946 (N_12946,N_12621,N_12614);
nand U12947 (N_12947,N_12620,N_12846);
or U12948 (N_12948,N_12784,N_12671);
and U12949 (N_12949,N_12825,N_12667);
nand U12950 (N_12950,N_12806,N_12631);
nand U12951 (N_12951,N_12801,N_12737);
xnor U12952 (N_12952,N_12822,N_12858);
and U12953 (N_12953,N_12721,N_12713);
nand U12954 (N_12954,N_12649,N_12670);
or U12955 (N_12955,N_12627,N_12644);
or U12956 (N_12956,N_12812,N_12669);
and U12957 (N_12957,N_12658,N_12898);
nor U12958 (N_12958,N_12888,N_12640);
xor U12959 (N_12959,N_12823,N_12853);
nor U12960 (N_12960,N_12641,N_12887);
nor U12961 (N_12961,N_12704,N_12884);
nor U12962 (N_12962,N_12840,N_12660);
nor U12963 (N_12963,N_12663,N_12869);
and U12964 (N_12964,N_12839,N_12726);
nand U12965 (N_12965,N_12686,N_12680);
nor U12966 (N_12966,N_12765,N_12604);
nor U12967 (N_12967,N_12834,N_12809);
or U12968 (N_12968,N_12843,N_12730);
nand U12969 (N_12969,N_12740,N_12694);
or U12970 (N_12970,N_12662,N_12792);
and U12971 (N_12971,N_12611,N_12624);
and U12972 (N_12972,N_12876,N_12701);
nor U12973 (N_12973,N_12601,N_12715);
and U12974 (N_12974,N_12836,N_12675);
xnor U12975 (N_12975,N_12717,N_12755);
nand U12976 (N_12976,N_12841,N_12699);
nor U12977 (N_12977,N_12753,N_12657);
xnor U12978 (N_12978,N_12747,N_12827);
and U12979 (N_12979,N_12678,N_12757);
nor U12980 (N_12980,N_12880,N_12692);
and U12981 (N_12981,N_12727,N_12829);
or U12982 (N_12982,N_12861,N_12643);
or U12983 (N_12983,N_12778,N_12877);
and U12984 (N_12984,N_12622,N_12883);
or U12985 (N_12985,N_12850,N_12703);
or U12986 (N_12986,N_12868,N_12808);
nor U12987 (N_12987,N_12741,N_12735);
xor U12988 (N_12988,N_12634,N_12800);
xor U12989 (N_12989,N_12719,N_12666);
nor U12990 (N_12990,N_12654,N_12835);
and U12991 (N_12991,N_12676,N_12602);
or U12992 (N_12992,N_12710,N_12859);
or U12993 (N_12993,N_12743,N_12864);
and U12994 (N_12994,N_12632,N_12650);
and U12995 (N_12995,N_12700,N_12745);
nor U12996 (N_12996,N_12807,N_12695);
or U12997 (N_12997,N_12724,N_12718);
nor U12998 (N_12998,N_12702,N_12672);
nor U12999 (N_12999,N_12754,N_12897);
xor U13000 (N_13000,N_12617,N_12682);
and U13001 (N_13001,N_12683,N_12638);
or U13002 (N_13002,N_12878,N_12679);
nor U13003 (N_13003,N_12733,N_12738);
xor U13004 (N_13004,N_12837,N_12790);
or U13005 (N_13005,N_12659,N_12619);
xor U13006 (N_13006,N_12639,N_12608);
or U13007 (N_13007,N_12892,N_12732);
nand U13008 (N_13008,N_12625,N_12729);
and U13009 (N_13009,N_12661,N_12681);
xor U13010 (N_13010,N_12849,N_12789);
nor U13011 (N_13011,N_12889,N_12748);
or U13012 (N_13012,N_12891,N_12651);
nand U13013 (N_13013,N_12794,N_12758);
nor U13014 (N_13014,N_12691,N_12819);
and U13015 (N_13015,N_12677,N_12776);
xor U13016 (N_13016,N_12690,N_12795);
or U13017 (N_13017,N_12612,N_12636);
nor U13018 (N_13018,N_12742,N_12652);
nand U13019 (N_13019,N_12817,N_12689);
nand U13020 (N_13020,N_12886,N_12811);
and U13021 (N_13021,N_12762,N_12866);
xor U13022 (N_13022,N_12766,N_12875);
xnor U13023 (N_13023,N_12714,N_12821);
xnor U13024 (N_13024,N_12629,N_12796);
and U13025 (N_13025,N_12696,N_12824);
nand U13026 (N_13026,N_12830,N_12739);
nor U13027 (N_13027,N_12863,N_12734);
or U13028 (N_13028,N_12899,N_12893);
nor U13029 (N_13029,N_12647,N_12793);
nor U13030 (N_13030,N_12782,N_12759);
nand U13031 (N_13031,N_12826,N_12787);
nand U13032 (N_13032,N_12610,N_12842);
or U13033 (N_13033,N_12791,N_12872);
or U13034 (N_13034,N_12857,N_12655);
and U13035 (N_13035,N_12814,N_12684);
nor U13036 (N_13036,N_12882,N_12777);
and U13037 (N_13037,N_12698,N_12813);
nand U13038 (N_13038,N_12769,N_12773);
nand U13039 (N_13039,N_12772,N_12798);
nor U13040 (N_13040,N_12785,N_12731);
xnor U13041 (N_13041,N_12764,N_12744);
or U13042 (N_13042,N_12767,N_12803);
nand U13043 (N_13043,N_12716,N_12705);
or U13044 (N_13044,N_12609,N_12896);
nor U13045 (N_13045,N_12642,N_12867);
or U13046 (N_13046,N_12860,N_12783);
nor U13047 (N_13047,N_12844,N_12815);
and U13048 (N_13048,N_12862,N_12775);
nor U13049 (N_13049,N_12802,N_12763);
xor U13050 (N_13050,N_12647,N_12819);
nand U13051 (N_13051,N_12808,N_12665);
and U13052 (N_13052,N_12600,N_12690);
nor U13053 (N_13053,N_12710,N_12660);
nand U13054 (N_13054,N_12752,N_12628);
nand U13055 (N_13055,N_12662,N_12823);
nand U13056 (N_13056,N_12606,N_12662);
nand U13057 (N_13057,N_12875,N_12751);
or U13058 (N_13058,N_12663,N_12611);
nand U13059 (N_13059,N_12696,N_12756);
nor U13060 (N_13060,N_12831,N_12782);
nand U13061 (N_13061,N_12887,N_12839);
and U13062 (N_13062,N_12888,N_12724);
and U13063 (N_13063,N_12867,N_12843);
xor U13064 (N_13064,N_12801,N_12847);
and U13065 (N_13065,N_12662,N_12795);
nand U13066 (N_13066,N_12668,N_12794);
and U13067 (N_13067,N_12841,N_12681);
and U13068 (N_13068,N_12670,N_12619);
or U13069 (N_13069,N_12654,N_12661);
nor U13070 (N_13070,N_12755,N_12663);
nand U13071 (N_13071,N_12678,N_12702);
or U13072 (N_13072,N_12708,N_12746);
or U13073 (N_13073,N_12892,N_12784);
nand U13074 (N_13074,N_12750,N_12794);
xnor U13075 (N_13075,N_12663,N_12893);
nand U13076 (N_13076,N_12792,N_12681);
and U13077 (N_13077,N_12838,N_12848);
nor U13078 (N_13078,N_12674,N_12821);
or U13079 (N_13079,N_12852,N_12748);
nor U13080 (N_13080,N_12843,N_12691);
and U13081 (N_13081,N_12703,N_12863);
nand U13082 (N_13082,N_12757,N_12847);
and U13083 (N_13083,N_12690,N_12705);
xor U13084 (N_13084,N_12892,N_12730);
nand U13085 (N_13085,N_12775,N_12645);
and U13086 (N_13086,N_12642,N_12750);
xnor U13087 (N_13087,N_12759,N_12837);
xnor U13088 (N_13088,N_12847,N_12763);
or U13089 (N_13089,N_12800,N_12620);
and U13090 (N_13090,N_12897,N_12604);
and U13091 (N_13091,N_12699,N_12840);
or U13092 (N_13092,N_12794,N_12636);
nand U13093 (N_13093,N_12857,N_12717);
nand U13094 (N_13094,N_12618,N_12739);
and U13095 (N_13095,N_12713,N_12615);
and U13096 (N_13096,N_12878,N_12701);
nand U13097 (N_13097,N_12854,N_12836);
or U13098 (N_13098,N_12707,N_12894);
and U13099 (N_13099,N_12666,N_12602);
and U13100 (N_13100,N_12885,N_12613);
nand U13101 (N_13101,N_12652,N_12883);
or U13102 (N_13102,N_12772,N_12736);
or U13103 (N_13103,N_12779,N_12628);
xnor U13104 (N_13104,N_12696,N_12803);
or U13105 (N_13105,N_12764,N_12806);
nor U13106 (N_13106,N_12601,N_12735);
nand U13107 (N_13107,N_12822,N_12615);
xor U13108 (N_13108,N_12897,N_12828);
xor U13109 (N_13109,N_12601,N_12644);
and U13110 (N_13110,N_12724,N_12843);
nor U13111 (N_13111,N_12730,N_12845);
and U13112 (N_13112,N_12882,N_12709);
nand U13113 (N_13113,N_12612,N_12698);
and U13114 (N_13114,N_12601,N_12771);
and U13115 (N_13115,N_12832,N_12688);
or U13116 (N_13116,N_12851,N_12833);
nor U13117 (N_13117,N_12728,N_12831);
nor U13118 (N_13118,N_12700,N_12690);
and U13119 (N_13119,N_12883,N_12872);
and U13120 (N_13120,N_12886,N_12860);
and U13121 (N_13121,N_12884,N_12718);
nor U13122 (N_13122,N_12738,N_12847);
and U13123 (N_13123,N_12876,N_12680);
nor U13124 (N_13124,N_12646,N_12880);
nor U13125 (N_13125,N_12678,N_12606);
nand U13126 (N_13126,N_12749,N_12853);
nor U13127 (N_13127,N_12788,N_12810);
or U13128 (N_13128,N_12691,N_12606);
xnor U13129 (N_13129,N_12858,N_12808);
xor U13130 (N_13130,N_12622,N_12786);
nand U13131 (N_13131,N_12722,N_12745);
or U13132 (N_13132,N_12628,N_12708);
and U13133 (N_13133,N_12876,N_12668);
and U13134 (N_13134,N_12709,N_12847);
nor U13135 (N_13135,N_12633,N_12789);
or U13136 (N_13136,N_12668,N_12838);
nand U13137 (N_13137,N_12751,N_12690);
nand U13138 (N_13138,N_12621,N_12626);
or U13139 (N_13139,N_12874,N_12764);
nand U13140 (N_13140,N_12616,N_12693);
or U13141 (N_13141,N_12783,N_12690);
nand U13142 (N_13142,N_12618,N_12693);
and U13143 (N_13143,N_12888,N_12887);
or U13144 (N_13144,N_12671,N_12746);
nor U13145 (N_13145,N_12646,N_12686);
nand U13146 (N_13146,N_12837,N_12787);
nand U13147 (N_13147,N_12870,N_12703);
or U13148 (N_13148,N_12799,N_12794);
nor U13149 (N_13149,N_12712,N_12758);
and U13150 (N_13150,N_12742,N_12645);
or U13151 (N_13151,N_12661,N_12832);
and U13152 (N_13152,N_12767,N_12794);
nand U13153 (N_13153,N_12608,N_12845);
xnor U13154 (N_13154,N_12670,N_12851);
xor U13155 (N_13155,N_12775,N_12732);
or U13156 (N_13156,N_12762,N_12638);
or U13157 (N_13157,N_12813,N_12774);
nand U13158 (N_13158,N_12833,N_12890);
and U13159 (N_13159,N_12727,N_12646);
and U13160 (N_13160,N_12683,N_12875);
and U13161 (N_13161,N_12744,N_12803);
nor U13162 (N_13162,N_12706,N_12683);
nand U13163 (N_13163,N_12649,N_12751);
xnor U13164 (N_13164,N_12772,N_12636);
and U13165 (N_13165,N_12608,N_12697);
nand U13166 (N_13166,N_12820,N_12767);
and U13167 (N_13167,N_12876,N_12855);
and U13168 (N_13168,N_12684,N_12833);
or U13169 (N_13169,N_12653,N_12721);
or U13170 (N_13170,N_12794,N_12742);
nand U13171 (N_13171,N_12633,N_12824);
and U13172 (N_13172,N_12661,N_12842);
or U13173 (N_13173,N_12605,N_12721);
nor U13174 (N_13174,N_12698,N_12742);
nand U13175 (N_13175,N_12600,N_12712);
nand U13176 (N_13176,N_12831,N_12629);
xor U13177 (N_13177,N_12603,N_12878);
xor U13178 (N_13178,N_12641,N_12611);
nor U13179 (N_13179,N_12742,N_12803);
nand U13180 (N_13180,N_12623,N_12735);
xnor U13181 (N_13181,N_12891,N_12863);
xor U13182 (N_13182,N_12774,N_12605);
nand U13183 (N_13183,N_12687,N_12822);
and U13184 (N_13184,N_12846,N_12841);
nand U13185 (N_13185,N_12718,N_12649);
nor U13186 (N_13186,N_12699,N_12736);
xor U13187 (N_13187,N_12698,N_12672);
nor U13188 (N_13188,N_12693,N_12794);
xor U13189 (N_13189,N_12699,N_12895);
xnor U13190 (N_13190,N_12601,N_12604);
xor U13191 (N_13191,N_12672,N_12637);
xnor U13192 (N_13192,N_12866,N_12650);
nand U13193 (N_13193,N_12627,N_12751);
nor U13194 (N_13194,N_12785,N_12655);
nor U13195 (N_13195,N_12871,N_12891);
xor U13196 (N_13196,N_12870,N_12823);
nor U13197 (N_13197,N_12629,N_12661);
nor U13198 (N_13198,N_12732,N_12607);
and U13199 (N_13199,N_12878,N_12803);
and U13200 (N_13200,N_13027,N_13150);
and U13201 (N_13201,N_12920,N_12932);
xor U13202 (N_13202,N_13084,N_13077);
or U13203 (N_13203,N_13160,N_13170);
or U13204 (N_13204,N_12957,N_13165);
xnor U13205 (N_13205,N_12952,N_13029);
or U13206 (N_13206,N_13009,N_12962);
xnor U13207 (N_13207,N_13078,N_13129);
nand U13208 (N_13208,N_12995,N_13106);
nand U13209 (N_13209,N_12965,N_13101);
nand U13210 (N_13210,N_12946,N_13064);
nor U13211 (N_13211,N_13110,N_12900);
and U13212 (N_13212,N_13072,N_13182);
xor U13213 (N_13213,N_13112,N_12989);
nand U13214 (N_13214,N_13046,N_13004);
nor U13215 (N_13215,N_12935,N_12934);
nor U13216 (N_13216,N_12955,N_12994);
and U13217 (N_13217,N_13074,N_13080);
and U13218 (N_13218,N_12944,N_13087);
and U13219 (N_13219,N_13034,N_13193);
xor U13220 (N_13220,N_13091,N_12980);
nor U13221 (N_13221,N_13070,N_13013);
or U13222 (N_13222,N_12976,N_13048);
nor U13223 (N_13223,N_12907,N_13059);
or U13224 (N_13224,N_13017,N_13179);
nand U13225 (N_13225,N_12982,N_13020);
xnor U13226 (N_13226,N_13126,N_13154);
xnor U13227 (N_13227,N_13146,N_13036);
and U13228 (N_13228,N_13163,N_12922);
nand U13229 (N_13229,N_12974,N_13184);
nor U13230 (N_13230,N_13079,N_13134);
or U13231 (N_13231,N_13192,N_12970);
nor U13232 (N_13232,N_12927,N_13132);
nand U13233 (N_13233,N_12903,N_12928);
nand U13234 (N_13234,N_12918,N_12967);
or U13235 (N_13235,N_13001,N_13109);
xor U13236 (N_13236,N_13195,N_13007);
nor U13237 (N_13237,N_13062,N_13143);
nor U13238 (N_13238,N_12953,N_13066);
xor U13239 (N_13239,N_13194,N_12964);
xnor U13240 (N_13240,N_13090,N_13023);
xor U13241 (N_13241,N_13118,N_12924);
nand U13242 (N_13242,N_12998,N_13016);
nand U13243 (N_13243,N_12908,N_13071);
or U13244 (N_13244,N_13044,N_13128);
nand U13245 (N_13245,N_13014,N_12979);
and U13246 (N_13246,N_12996,N_12960);
and U13247 (N_13247,N_13073,N_13124);
nand U13248 (N_13248,N_13125,N_13075);
and U13249 (N_13249,N_13187,N_13190);
and U13250 (N_13250,N_13120,N_13005);
and U13251 (N_13251,N_13156,N_12941);
nor U13252 (N_13252,N_13127,N_12939);
nand U13253 (N_13253,N_13123,N_13056);
and U13254 (N_13254,N_13041,N_13022);
or U13255 (N_13255,N_13038,N_13099);
and U13256 (N_13256,N_13142,N_12992);
xnor U13257 (N_13257,N_12930,N_12902);
or U13258 (N_13258,N_13122,N_12910);
and U13259 (N_13259,N_12916,N_13057);
xor U13260 (N_13260,N_13051,N_12943);
and U13261 (N_13261,N_12954,N_13003);
nand U13262 (N_13262,N_13133,N_13089);
xor U13263 (N_13263,N_12985,N_13053);
xnor U13264 (N_13264,N_12983,N_13010);
xor U13265 (N_13265,N_13082,N_13006);
nand U13266 (N_13266,N_12906,N_13037);
nand U13267 (N_13267,N_13097,N_13063);
or U13268 (N_13268,N_13111,N_13173);
and U13269 (N_13269,N_13196,N_12926);
xnor U13270 (N_13270,N_13104,N_13054);
or U13271 (N_13271,N_13015,N_13168);
nor U13272 (N_13272,N_13065,N_13076);
nand U13273 (N_13273,N_13145,N_12959);
nand U13274 (N_13274,N_12945,N_13177);
and U13275 (N_13275,N_12971,N_12972);
xnor U13276 (N_13276,N_13000,N_13171);
or U13277 (N_13277,N_13026,N_13052);
xor U13278 (N_13278,N_13121,N_13039);
and U13279 (N_13279,N_13148,N_13093);
or U13280 (N_13280,N_12921,N_12909);
xnor U13281 (N_13281,N_13119,N_13117);
and U13282 (N_13282,N_12968,N_12986);
xor U13283 (N_13283,N_13113,N_13152);
nand U13284 (N_13284,N_13030,N_13167);
nor U13285 (N_13285,N_13050,N_13102);
xnor U13286 (N_13286,N_12938,N_12984);
nor U13287 (N_13287,N_13021,N_13094);
nor U13288 (N_13288,N_12947,N_13067);
nor U13289 (N_13289,N_13183,N_12914);
nand U13290 (N_13290,N_12923,N_12937);
or U13291 (N_13291,N_13019,N_13164);
and U13292 (N_13292,N_12981,N_12929);
nand U13293 (N_13293,N_12956,N_13033);
nand U13294 (N_13294,N_13186,N_12949);
and U13295 (N_13295,N_13086,N_13103);
or U13296 (N_13296,N_13155,N_13159);
xor U13297 (N_13297,N_13096,N_13040);
and U13298 (N_13298,N_13185,N_12997);
xor U13299 (N_13299,N_13138,N_13002);
or U13300 (N_13300,N_13098,N_12940);
xnor U13301 (N_13301,N_12966,N_12951);
and U13302 (N_13302,N_12933,N_13025);
or U13303 (N_13303,N_13197,N_12987);
nand U13304 (N_13304,N_12942,N_12961);
xor U13305 (N_13305,N_13162,N_12991);
or U13306 (N_13306,N_13035,N_13105);
xor U13307 (N_13307,N_12931,N_13068);
or U13308 (N_13308,N_12915,N_13172);
nand U13309 (N_13309,N_13141,N_13139);
xnor U13310 (N_13310,N_13137,N_12978);
and U13311 (N_13311,N_13085,N_13083);
or U13312 (N_13312,N_13191,N_13095);
or U13313 (N_13313,N_13147,N_13045);
or U13314 (N_13314,N_12990,N_13061);
nand U13315 (N_13315,N_13060,N_12917);
nand U13316 (N_13316,N_12948,N_13136);
nand U13317 (N_13317,N_13130,N_13131);
nor U13318 (N_13318,N_12911,N_12936);
nor U13319 (N_13319,N_13049,N_13140);
xnor U13320 (N_13320,N_13178,N_13181);
xor U13321 (N_13321,N_12905,N_13024);
or U13322 (N_13322,N_13161,N_13153);
and U13323 (N_13323,N_13166,N_13135);
xor U13324 (N_13324,N_12950,N_13198);
xor U13325 (N_13325,N_13032,N_13081);
and U13326 (N_13326,N_13175,N_12999);
and U13327 (N_13327,N_13169,N_13012);
xor U13328 (N_13328,N_13042,N_12963);
and U13329 (N_13329,N_13088,N_13028);
and U13330 (N_13330,N_13174,N_13114);
and U13331 (N_13331,N_13158,N_12977);
or U13332 (N_13332,N_13188,N_12904);
or U13333 (N_13333,N_13011,N_13058);
nor U13334 (N_13334,N_13176,N_12912);
xor U13335 (N_13335,N_13043,N_12993);
or U13336 (N_13336,N_13092,N_13069);
and U13337 (N_13337,N_13031,N_12958);
or U13338 (N_13338,N_13055,N_12975);
nor U13339 (N_13339,N_13144,N_13115);
nor U13340 (N_13340,N_13151,N_12901);
and U13341 (N_13341,N_12919,N_13047);
and U13342 (N_13342,N_12913,N_13018);
xnor U13343 (N_13343,N_13107,N_13180);
nor U13344 (N_13344,N_13116,N_13157);
nand U13345 (N_13345,N_12969,N_13108);
nor U13346 (N_13346,N_12988,N_12925);
nand U13347 (N_13347,N_13100,N_13149);
and U13348 (N_13348,N_13199,N_13189);
nand U13349 (N_13349,N_13008,N_12973);
and U13350 (N_13350,N_13014,N_12939);
and U13351 (N_13351,N_12942,N_13183);
xnor U13352 (N_13352,N_12921,N_13082);
nor U13353 (N_13353,N_12913,N_13003);
xor U13354 (N_13354,N_12942,N_13135);
or U13355 (N_13355,N_12933,N_12938);
xnor U13356 (N_13356,N_13176,N_13029);
nand U13357 (N_13357,N_13023,N_13035);
and U13358 (N_13358,N_13098,N_13011);
xor U13359 (N_13359,N_13007,N_13078);
or U13360 (N_13360,N_13095,N_13003);
nand U13361 (N_13361,N_12929,N_13085);
and U13362 (N_13362,N_13137,N_13145);
nand U13363 (N_13363,N_13133,N_12906);
nor U13364 (N_13364,N_13110,N_13068);
or U13365 (N_13365,N_13184,N_12992);
or U13366 (N_13366,N_12975,N_13168);
nor U13367 (N_13367,N_12947,N_12919);
nor U13368 (N_13368,N_13084,N_13072);
nand U13369 (N_13369,N_13138,N_13120);
nor U13370 (N_13370,N_12911,N_13129);
and U13371 (N_13371,N_13187,N_13001);
nand U13372 (N_13372,N_12941,N_13194);
and U13373 (N_13373,N_13005,N_13078);
or U13374 (N_13374,N_13126,N_12992);
nand U13375 (N_13375,N_13035,N_13130);
nand U13376 (N_13376,N_13103,N_13175);
or U13377 (N_13377,N_13133,N_13193);
or U13378 (N_13378,N_13181,N_12932);
xor U13379 (N_13379,N_13167,N_12975);
nand U13380 (N_13380,N_13180,N_13141);
and U13381 (N_13381,N_12977,N_12937);
nand U13382 (N_13382,N_13079,N_13159);
nand U13383 (N_13383,N_13180,N_13194);
and U13384 (N_13384,N_12933,N_12986);
and U13385 (N_13385,N_12991,N_12920);
nor U13386 (N_13386,N_13053,N_12922);
or U13387 (N_13387,N_13175,N_13039);
nor U13388 (N_13388,N_12944,N_13188);
xnor U13389 (N_13389,N_13042,N_13083);
nand U13390 (N_13390,N_13183,N_13181);
nor U13391 (N_13391,N_12976,N_13080);
or U13392 (N_13392,N_13023,N_13128);
nor U13393 (N_13393,N_13088,N_12919);
and U13394 (N_13394,N_13057,N_13150);
xor U13395 (N_13395,N_12926,N_12979);
xor U13396 (N_13396,N_13013,N_13009);
or U13397 (N_13397,N_13002,N_13003);
nand U13398 (N_13398,N_13095,N_13012);
or U13399 (N_13399,N_13126,N_13001);
nand U13400 (N_13400,N_12941,N_13187);
xor U13401 (N_13401,N_12911,N_12997);
or U13402 (N_13402,N_12975,N_13188);
or U13403 (N_13403,N_13053,N_13098);
and U13404 (N_13404,N_13151,N_13027);
nand U13405 (N_13405,N_12991,N_12913);
nor U13406 (N_13406,N_13176,N_12975);
xor U13407 (N_13407,N_13062,N_13047);
or U13408 (N_13408,N_12915,N_13168);
and U13409 (N_13409,N_13186,N_13003);
nand U13410 (N_13410,N_13000,N_13150);
and U13411 (N_13411,N_13163,N_13052);
nor U13412 (N_13412,N_13188,N_12932);
or U13413 (N_13413,N_13181,N_13118);
and U13414 (N_13414,N_12939,N_13171);
and U13415 (N_13415,N_13100,N_13122);
nor U13416 (N_13416,N_12988,N_12998);
or U13417 (N_13417,N_13179,N_13165);
and U13418 (N_13418,N_13086,N_13127);
xor U13419 (N_13419,N_12985,N_13060);
or U13420 (N_13420,N_12978,N_13149);
or U13421 (N_13421,N_13155,N_13000);
xnor U13422 (N_13422,N_12997,N_13016);
xor U13423 (N_13423,N_13110,N_13002);
xnor U13424 (N_13424,N_13010,N_12901);
or U13425 (N_13425,N_12918,N_12990);
nor U13426 (N_13426,N_12948,N_13109);
xnor U13427 (N_13427,N_13188,N_12907);
or U13428 (N_13428,N_13175,N_13090);
or U13429 (N_13429,N_12925,N_13026);
and U13430 (N_13430,N_13095,N_12975);
nor U13431 (N_13431,N_13091,N_13075);
xnor U13432 (N_13432,N_13126,N_13043);
nor U13433 (N_13433,N_13186,N_12925);
or U13434 (N_13434,N_13142,N_12966);
and U13435 (N_13435,N_13081,N_13048);
xnor U13436 (N_13436,N_13177,N_13186);
xor U13437 (N_13437,N_13044,N_13050);
nand U13438 (N_13438,N_12919,N_13079);
xnor U13439 (N_13439,N_12991,N_13147);
nand U13440 (N_13440,N_13052,N_13181);
and U13441 (N_13441,N_13037,N_13171);
nand U13442 (N_13442,N_12909,N_12968);
nand U13443 (N_13443,N_13068,N_13007);
xnor U13444 (N_13444,N_13165,N_12959);
or U13445 (N_13445,N_13180,N_13162);
or U13446 (N_13446,N_13119,N_12971);
and U13447 (N_13447,N_13086,N_13101);
nor U13448 (N_13448,N_13116,N_12987);
nand U13449 (N_13449,N_13101,N_13173);
nor U13450 (N_13450,N_12962,N_13197);
nor U13451 (N_13451,N_12994,N_12968);
xor U13452 (N_13452,N_13176,N_13047);
xnor U13453 (N_13453,N_12973,N_13002);
or U13454 (N_13454,N_13158,N_12919);
xnor U13455 (N_13455,N_13047,N_13152);
or U13456 (N_13456,N_13043,N_13066);
or U13457 (N_13457,N_13161,N_13131);
nand U13458 (N_13458,N_12930,N_13164);
nand U13459 (N_13459,N_13118,N_13028);
and U13460 (N_13460,N_13158,N_12944);
or U13461 (N_13461,N_13049,N_13096);
or U13462 (N_13462,N_12920,N_13087);
nand U13463 (N_13463,N_13118,N_13105);
or U13464 (N_13464,N_13014,N_12942);
xor U13465 (N_13465,N_12924,N_13193);
or U13466 (N_13466,N_13000,N_13100);
nor U13467 (N_13467,N_13086,N_13173);
or U13468 (N_13468,N_12917,N_13137);
nor U13469 (N_13469,N_12984,N_13145);
or U13470 (N_13470,N_13157,N_13098);
or U13471 (N_13471,N_13017,N_13096);
nor U13472 (N_13472,N_12964,N_12918);
nor U13473 (N_13473,N_13052,N_12949);
xor U13474 (N_13474,N_13128,N_13143);
and U13475 (N_13475,N_13001,N_12925);
xnor U13476 (N_13476,N_13126,N_13110);
and U13477 (N_13477,N_12933,N_13033);
xnor U13478 (N_13478,N_13160,N_13018);
nand U13479 (N_13479,N_12958,N_13137);
xor U13480 (N_13480,N_13112,N_13118);
or U13481 (N_13481,N_12949,N_12946);
xor U13482 (N_13482,N_13103,N_13068);
nand U13483 (N_13483,N_13115,N_13152);
xnor U13484 (N_13484,N_12952,N_13005);
and U13485 (N_13485,N_13062,N_13081);
xor U13486 (N_13486,N_13103,N_13066);
nor U13487 (N_13487,N_13181,N_12987);
nor U13488 (N_13488,N_13022,N_13170);
or U13489 (N_13489,N_13078,N_13046);
xnor U13490 (N_13490,N_13175,N_13173);
nand U13491 (N_13491,N_13084,N_12918);
and U13492 (N_13492,N_12949,N_13047);
nand U13493 (N_13493,N_13045,N_13176);
nor U13494 (N_13494,N_13053,N_13034);
xor U13495 (N_13495,N_13017,N_13178);
nand U13496 (N_13496,N_13179,N_12932);
nand U13497 (N_13497,N_13107,N_12950);
nor U13498 (N_13498,N_12937,N_12971);
nor U13499 (N_13499,N_13133,N_12945);
or U13500 (N_13500,N_13269,N_13414);
nand U13501 (N_13501,N_13218,N_13245);
or U13502 (N_13502,N_13205,N_13338);
or U13503 (N_13503,N_13479,N_13342);
nand U13504 (N_13504,N_13200,N_13207);
and U13505 (N_13505,N_13247,N_13419);
xor U13506 (N_13506,N_13458,N_13266);
xnor U13507 (N_13507,N_13295,N_13391);
and U13508 (N_13508,N_13324,N_13372);
nand U13509 (N_13509,N_13322,N_13251);
and U13510 (N_13510,N_13480,N_13422);
nor U13511 (N_13511,N_13477,N_13481);
and U13512 (N_13512,N_13380,N_13339);
xor U13513 (N_13513,N_13283,N_13346);
and U13514 (N_13514,N_13433,N_13341);
nand U13515 (N_13515,N_13278,N_13460);
or U13516 (N_13516,N_13489,N_13212);
and U13517 (N_13517,N_13242,N_13457);
or U13518 (N_13518,N_13332,N_13485);
and U13519 (N_13519,N_13470,N_13469);
or U13520 (N_13520,N_13349,N_13415);
nor U13521 (N_13521,N_13314,N_13467);
nor U13522 (N_13522,N_13383,N_13413);
xnor U13523 (N_13523,N_13401,N_13461);
nor U13524 (N_13524,N_13289,N_13454);
or U13525 (N_13525,N_13351,N_13226);
and U13526 (N_13526,N_13224,N_13325);
nor U13527 (N_13527,N_13464,N_13275);
nand U13528 (N_13528,N_13263,N_13434);
or U13529 (N_13529,N_13265,N_13403);
xor U13530 (N_13530,N_13345,N_13233);
and U13531 (N_13531,N_13462,N_13281);
nand U13532 (N_13532,N_13444,N_13409);
xor U13533 (N_13533,N_13276,N_13300);
xnor U13534 (N_13534,N_13468,N_13273);
xor U13535 (N_13535,N_13363,N_13296);
and U13536 (N_13536,N_13347,N_13394);
and U13537 (N_13537,N_13491,N_13404);
nor U13538 (N_13538,N_13298,N_13297);
and U13539 (N_13539,N_13406,N_13411);
or U13540 (N_13540,N_13309,N_13228);
nand U13541 (N_13541,N_13211,N_13216);
and U13542 (N_13542,N_13340,N_13438);
nand U13543 (N_13543,N_13343,N_13279);
or U13544 (N_13544,N_13356,N_13234);
and U13545 (N_13545,N_13416,N_13282);
nand U13546 (N_13546,N_13405,N_13407);
and U13547 (N_13547,N_13476,N_13376);
or U13548 (N_13548,N_13328,N_13313);
xnor U13549 (N_13549,N_13478,N_13486);
nand U13550 (N_13550,N_13291,N_13379);
and U13551 (N_13551,N_13494,N_13261);
nor U13552 (N_13552,N_13255,N_13429);
and U13553 (N_13553,N_13493,N_13483);
or U13554 (N_13554,N_13204,N_13421);
or U13555 (N_13555,N_13437,N_13412);
nor U13556 (N_13556,N_13285,N_13288);
or U13557 (N_13557,N_13495,N_13369);
nor U13558 (N_13558,N_13243,N_13430);
and U13559 (N_13559,N_13327,N_13417);
xnor U13560 (N_13560,N_13286,N_13439);
nand U13561 (N_13561,N_13397,N_13259);
nand U13562 (N_13562,N_13358,N_13331);
or U13563 (N_13563,N_13498,N_13219);
and U13564 (N_13564,N_13353,N_13487);
and U13565 (N_13565,N_13250,N_13350);
or U13566 (N_13566,N_13293,N_13221);
and U13567 (N_13567,N_13240,N_13371);
and U13568 (N_13568,N_13337,N_13451);
xnor U13569 (N_13569,N_13410,N_13492);
nand U13570 (N_13570,N_13215,N_13284);
nand U13571 (N_13571,N_13248,N_13348);
or U13572 (N_13572,N_13287,N_13446);
or U13573 (N_13573,N_13267,N_13333);
or U13574 (N_13574,N_13424,N_13223);
and U13575 (N_13575,N_13323,N_13236);
nand U13576 (N_13576,N_13299,N_13402);
or U13577 (N_13577,N_13482,N_13329);
nor U13578 (N_13578,N_13209,N_13496);
and U13579 (N_13579,N_13393,N_13326);
nor U13580 (N_13580,N_13423,N_13208);
nand U13581 (N_13581,N_13271,N_13244);
nand U13582 (N_13582,N_13474,N_13431);
nand U13583 (N_13583,N_13443,N_13452);
and U13584 (N_13584,N_13442,N_13378);
or U13585 (N_13585,N_13471,N_13453);
nor U13586 (N_13586,N_13373,N_13315);
and U13587 (N_13587,N_13449,N_13355);
xor U13588 (N_13588,N_13260,N_13303);
xnor U13589 (N_13589,N_13440,N_13395);
nand U13590 (N_13590,N_13365,N_13490);
nand U13591 (N_13591,N_13396,N_13357);
xor U13592 (N_13592,N_13320,N_13305);
nand U13593 (N_13593,N_13203,N_13465);
nand U13594 (N_13594,N_13381,N_13249);
and U13595 (N_13595,N_13210,N_13304);
xnor U13596 (N_13596,N_13385,N_13354);
or U13597 (N_13597,N_13231,N_13336);
nor U13598 (N_13598,N_13316,N_13307);
nor U13599 (N_13599,N_13206,N_13466);
or U13600 (N_13600,N_13280,N_13214);
xor U13601 (N_13601,N_13344,N_13277);
or U13602 (N_13602,N_13398,N_13272);
nor U13603 (N_13603,N_13241,N_13377);
nor U13604 (N_13604,N_13256,N_13426);
and U13605 (N_13605,N_13229,N_13235);
and U13606 (N_13606,N_13238,N_13268);
xnor U13607 (N_13607,N_13435,N_13254);
nor U13608 (N_13608,N_13384,N_13463);
xnor U13609 (N_13609,N_13484,N_13366);
and U13610 (N_13610,N_13253,N_13472);
and U13611 (N_13611,N_13499,N_13319);
and U13612 (N_13612,N_13374,N_13428);
nor U13613 (N_13613,N_13274,N_13232);
nor U13614 (N_13614,N_13213,N_13389);
or U13615 (N_13615,N_13222,N_13441);
and U13616 (N_13616,N_13257,N_13359);
xor U13617 (N_13617,N_13217,N_13392);
nand U13618 (N_13618,N_13450,N_13400);
or U13619 (N_13619,N_13367,N_13201);
and U13620 (N_13620,N_13448,N_13361);
xnor U13621 (N_13621,N_13246,N_13311);
xnor U13622 (N_13622,N_13375,N_13227);
xnor U13623 (N_13623,N_13230,N_13262);
or U13624 (N_13624,N_13264,N_13445);
nand U13625 (N_13625,N_13301,N_13387);
nand U13626 (N_13626,N_13306,N_13447);
nand U13627 (N_13627,N_13290,N_13317);
xnor U13628 (N_13628,N_13459,N_13370);
and U13629 (N_13629,N_13252,N_13488);
and U13630 (N_13630,N_13334,N_13408);
nand U13631 (N_13631,N_13456,N_13399);
or U13632 (N_13632,N_13237,N_13302);
nand U13633 (N_13633,N_13225,N_13418);
xnor U13634 (N_13634,N_13425,N_13388);
or U13635 (N_13635,N_13312,N_13382);
nor U13636 (N_13636,N_13294,N_13335);
xor U13637 (N_13637,N_13202,N_13455);
xnor U13638 (N_13638,N_13436,N_13292);
xnor U13639 (N_13639,N_13364,N_13270);
nand U13640 (N_13640,N_13308,N_13386);
xor U13641 (N_13641,N_13420,N_13473);
nor U13642 (N_13642,N_13318,N_13220);
and U13643 (N_13643,N_13310,N_13321);
nand U13644 (N_13644,N_13497,N_13360);
and U13645 (N_13645,N_13352,N_13330);
nand U13646 (N_13646,N_13427,N_13258);
xnor U13647 (N_13647,N_13368,N_13362);
nand U13648 (N_13648,N_13475,N_13239);
xor U13649 (N_13649,N_13432,N_13390);
and U13650 (N_13650,N_13268,N_13220);
or U13651 (N_13651,N_13257,N_13217);
xor U13652 (N_13652,N_13242,N_13488);
or U13653 (N_13653,N_13419,N_13280);
and U13654 (N_13654,N_13481,N_13252);
xnor U13655 (N_13655,N_13344,N_13372);
and U13656 (N_13656,N_13228,N_13362);
or U13657 (N_13657,N_13334,N_13401);
nor U13658 (N_13658,N_13240,N_13407);
or U13659 (N_13659,N_13393,N_13287);
nor U13660 (N_13660,N_13301,N_13356);
nand U13661 (N_13661,N_13263,N_13242);
nor U13662 (N_13662,N_13326,N_13304);
and U13663 (N_13663,N_13294,N_13428);
nand U13664 (N_13664,N_13233,N_13453);
xor U13665 (N_13665,N_13420,N_13424);
nor U13666 (N_13666,N_13453,N_13386);
nor U13667 (N_13667,N_13420,N_13214);
xor U13668 (N_13668,N_13462,N_13325);
and U13669 (N_13669,N_13327,N_13413);
xor U13670 (N_13670,N_13295,N_13302);
and U13671 (N_13671,N_13409,N_13278);
and U13672 (N_13672,N_13214,N_13499);
xnor U13673 (N_13673,N_13438,N_13219);
nand U13674 (N_13674,N_13384,N_13445);
or U13675 (N_13675,N_13445,N_13341);
and U13676 (N_13676,N_13326,N_13317);
xnor U13677 (N_13677,N_13437,N_13461);
nand U13678 (N_13678,N_13324,N_13412);
and U13679 (N_13679,N_13418,N_13470);
or U13680 (N_13680,N_13475,N_13431);
xnor U13681 (N_13681,N_13415,N_13495);
or U13682 (N_13682,N_13460,N_13468);
nor U13683 (N_13683,N_13249,N_13407);
and U13684 (N_13684,N_13275,N_13494);
or U13685 (N_13685,N_13295,N_13294);
xnor U13686 (N_13686,N_13370,N_13395);
xnor U13687 (N_13687,N_13376,N_13432);
xor U13688 (N_13688,N_13405,N_13424);
xor U13689 (N_13689,N_13439,N_13462);
or U13690 (N_13690,N_13266,N_13254);
or U13691 (N_13691,N_13499,N_13409);
nand U13692 (N_13692,N_13381,N_13485);
nor U13693 (N_13693,N_13394,N_13453);
nand U13694 (N_13694,N_13482,N_13298);
xnor U13695 (N_13695,N_13238,N_13403);
nor U13696 (N_13696,N_13241,N_13496);
nor U13697 (N_13697,N_13335,N_13348);
xnor U13698 (N_13698,N_13235,N_13202);
nand U13699 (N_13699,N_13499,N_13255);
or U13700 (N_13700,N_13264,N_13221);
or U13701 (N_13701,N_13205,N_13267);
xor U13702 (N_13702,N_13362,N_13320);
nor U13703 (N_13703,N_13402,N_13487);
xor U13704 (N_13704,N_13476,N_13332);
nand U13705 (N_13705,N_13497,N_13376);
nor U13706 (N_13706,N_13253,N_13430);
nand U13707 (N_13707,N_13307,N_13211);
nand U13708 (N_13708,N_13389,N_13422);
nand U13709 (N_13709,N_13468,N_13243);
nor U13710 (N_13710,N_13267,N_13305);
nand U13711 (N_13711,N_13352,N_13431);
and U13712 (N_13712,N_13391,N_13482);
xnor U13713 (N_13713,N_13412,N_13339);
nand U13714 (N_13714,N_13227,N_13305);
nand U13715 (N_13715,N_13211,N_13330);
and U13716 (N_13716,N_13475,N_13412);
or U13717 (N_13717,N_13409,N_13495);
nor U13718 (N_13718,N_13474,N_13364);
nand U13719 (N_13719,N_13490,N_13278);
or U13720 (N_13720,N_13409,N_13268);
nand U13721 (N_13721,N_13403,N_13475);
and U13722 (N_13722,N_13334,N_13483);
and U13723 (N_13723,N_13287,N_13327);
or U13724 (N_13724,N_13222,N_13413);
nor U13725 (N_13725,N_13228,N_13245);
and U13726 (N_13726,N_13252,N_13420);
and U13727 (N_13727,N_13310,N_13214);
or U13728 (N_13728,N_13283,N_13237);
or U13729 (N_13729,N_13275,N_13324);
nand U13730 (N_13730,N_13360,N_13340);
nor U13731 (N_13731,N_13373,N_13247);
and U13732 (N_13732,N_13303,N_13375);
nand U13733 (N_13733,N_13414,N_13437);
xor U13734 (N_13734,N_13311,N_13284);
nor U13735 (N_13735,N_13439,N_13300);
nand U13736 (N_13736,N_13408,N_13415);
nand U13737 (N_13737,N_13251,N_13258);
or U13738 (N_13738,N_13361,N_13491);
xnor U13739 (N_13739,N_13412,N_13469);
and U13740 (N_13740,N_13367,N_13478);
and U13741 (N_13741,N_13314,N_13271);
nor U13742 (N_13742,N_13354,N_13236);
and U13743 (N_13743,N_13274,N_13276);
nor U13744 (N_13744,N_13386,N_13226);
or U13745 (N_13745,N_13337,N_13223);
nand U13746 (N_13746,N_13461,N_13378);
and U13747 (N_13747,N_13215,N_13466);
nor U13748 (N_13748,N_13320,N_13353);
nand U13749 (N_13749,N_13328,N_13401);
nand U13750 (N_13750,N_13246,N_13496);
nand U13751 (N_13751,N_13239,N_13388);
or U13752 (N_13752,N_13471,N_13459);
or U13753 (N_13753,N_13360,N_13318);
and U13754 (N_13754,N_13432,N_13350);
nand U13755 (N_13755,N_13268,N_13453);
nand U13756 (N_13756,N_13349,N_13475);
or U13757 (N_13757,N_13415,N_13454);
xnor U13758 (N_13758,N_13313,N_13393);
nand U13759 (N_13759,N_13219,N_13463);
nor U13760 (N_13760,N_13282,N_13216);
xnor U13761 (N_13761,N_13272,N_13453);
nand U13762 (N_13762,N_13302,N_13220);
xor U13763 (N_13763,N_13349,N_13480);
or U13764 (N_13764,N_13298,N_13352);
nand U13765 (N_13765,N_13412,N_13427);
and U13766 (N_13766,N_13376,N_13462);
nor U13767 (N_13767,N_13461,N_13414);
nand U13768 (N_13768,N_13485,N_13356);
or U13769 (N_13769,N_13347,N_13435);
and U13770 (N_13770,N_13222,N_13368);
nand U13771 (N_13771,N_13401,N_13331);
and U13772 (N_13772,N_13403,N_13436);
nor U13773 (N_13773,N_13222,N_13410);
or U13774 (N_13774,N_13345,N_13332);
and U13775 (N_13775,N_13381,N_13231);
xor U13776 (N_13776,N_13328,N_13424);
xor U13777 (N_13777,N_13212,N_13429);
or U13778 (N_13778,N_13388,N_13288);
nor U13779 (N_13779,N_13297,N_13390);
and U13780 (N_13780,N_13408,N_13444);
nor U13781 (N_13781,N_13208,N_13211);
nor U13782 (N_13782,N_13299,N_13418);
xor U13783 (N_13783,N_13240,N_13466);
or U13784 (N_13784,N_13378,N_13455);
xnor U13785 (N_13785,N_13245,N_13439);
or U13786 (N_13786,N_13287,N_13329);
nand U13787 (N_13787,N_13259,N_13213);
and U13788 (N_13788,N_13235,N_13377);
nor U13789 (N_13789,N_13443,N_13229);
nand U13790 (N_13790,N_13260,N_13312);
nor U13791 (N_13791,N_13235,N_13259);
and U13792 (N_13792,N_13328,N_13454);
xor U13793 (N_13793,N_13269,N_13482);
or U13794 (N_13794,N_13343,N_13459);
xnor U13795 (N_13795,N_13385,N_13362);
or U13796 (N_13796,N_13389,N_13272);
or U13797 (N_13797,N_13461,N_13324);
and U13798 (N_13798,N_13246,N_13376);
and U13799 (N_13799,N_13463,N_13437);
nand U13800 (N_13800,N_13672,N_13783);
nand U13801 (N_13801,N_13654,N_13753);
nor U13802 (N_13802,N_13630,N_13511);
and U13803 (N_13803,N_13624,N_13618);
nand U13804 (N_13804,N_13636,N_13755);
nor U13805 (N_13805,N_13554,N_13524);
xor U13806 (N_13806,N_13669,N_13552);
nand U13807 (N_13807,N_13589,N_13586);
or U13808 (N_13808,N_13507,N_13612);
or U13809 (N_13809,N_13769,N_13547);
or U13810 (N_13810,N_13629,N_13601);
nand U13811 (N_13811,N_13757,N_13559);
nand U13812 (N_13812,N_13632,N_13527);
nand U13813 (N_13813,N_13637,N_13519);
xor U13814 (N_13814,N_13709,N_13739);
nand U13815 (N_13815,N_13711,N_13676);
or U13816 (N_13816,N_13797,N_13593);
nand U13817 (N_13817,N_13736,N_13787);
xnor U13818 (N_13818,N_13793,N_13714);
nand U13819 (N_13819,N_13608,N_13657);
or U13820 (N_13820,N_13509,N_13567);
or U13821 (N_13821,N_13515,N_13689);
xor U13822 (N_13822,N_13505,N_13772);
nand U13823 (N_13823,N_13707,N_13627);
or U13824 (N_13824,N_13747,N_13531);
nand U13825 (N_13825,N_13641,N_13616);
nand U13826 (N_13826,N_13546,N_13564);
and U13827 (N_13827,N_13710,N_13727);
xor U13828 (N_13828,N_13721,N_13642);
xnor U13829 (N_13829,N_13648,N_13674);
nor U13830 (N_13830,N_13678,N_13556);
and U13831 (N_13831,N_13786,N_13790);
nand U13832 (N_13832,N_13701,N_13516);
nor U13833 (N_13833,N_13743,N_13571);
or U13834 (N_13834,N_13599,N_13652);
nor U13835 (N_13835,N_13660,N_13502);
nand U13836 (N_13836,N_13538,N_13536);
xnor U13837 (N_13837,N_13759,N_13631);
nand U13838 (N_13838,N_13706,N_13661);
nand U13839 (N_13839,N_13735,N_13520);
xor U13840 (N_13840,N_13741,N_13639);
xnor U13841 (N_13841,N_13550,N_13724);
nand U13842 (N_13842,N_13667,N_13588);
and U13843 (N_13843,N_13795,N_13576);
or U13844 (N_13844,N_13776,N_13596);
xnor U13845 (N_13845,N_13728,N_13695);
nor U13846 (N_13846,N_13666,N_13633);
xnor U13847 (N_13847,N_13656,N_13694);
or U13848 (N_13848,N_13725,N_13553);
or U13849 (N_13849,N_13789,N_13578);
or U13850 (N_13850,N_13668,N_13503);
nor U13851 (N_13851,N_13508,N_13575);
nor U13852 (N_13852,N_13692,N_13771);
nand U13853 (N_13853,N_13574,N_13594);
and U13854 (N_13854,N_13526,N_13673);
nand U13855 (N_13855,N_13682,N_13785);
or U13856 (N_13856,N_13671,N_13796);
or U13857 (N_13857,N_13685,N_13653);
and U13858 (N_13858,N_13530,N_13730);
or U13859 (N_13859,N_13570,N_13767);
nor U13860 (N_13860,N_13592,N_13518);
or U13861 (N_13861,N_13696,N_13681);
or U13862 (N_13862,N_13646,N_13698);
or U13863 (N_13863,N_13609,N_13788);
and U13864 (N_13864,N_13623,N_13595);
and U13865 (N_13865,N_13504,N_13545);
nand U13866 (N_13866,N_13621,N_13640);
nand U13867 (N_13867,N_13742,N_13734);
nor U13868 (N_13868,N_13644,N_13606);
xnor U13869 (N_13869,N_13634,N_13523);
and U13870 (N_13870,N_13784,N_13712);
nor U13871 (N_13871,N_13791,N_13675);
or U13872 (N_13872,N_13602,N_13720);
or U13873 (N_13873,N_13563,N_13765);
or U13874 (N_13874,N_13611,N_13517);
or U13875 (N_13875,N_13568,N_13584);
and U13876 (N_13876,N_13732,N_13687);
nor U13877 (N_13877,N_13718,N_13548);
xnor U13878 (N_13878,N_13686,N_13717);
nand U13879 (N_13879,N_13600,N_13643);
and U13880 (N_13880,N_13778,N_13614);
and U13881 (N_13881,N_13615,N_13746);
or U13882 (N_13882,N_13697,N_13535);
and U13883 (N_13883,N_13770,N_13745);
or U13884 (N_13884,N_13604,N_13514);
and U13885 (N_13885,N_13731,N_13635);
nand U13886 (N_13886,N_13613,N_13645);
xnor U13887 (N_13887,N_13549,N_13617);
or U13888 (N_13888,N_13651,N_13665);
nor U13889 (N_13889,N_13537,N_13598);
or U13890 (N_13890,N_13756,N_13655);
xnor U13891 (N_13891,N_13699,N_13581);
or U13892 (N_13892,N_13569,N_13540);
and U13893 (N_13893,N_13691,N_13775);
nand U13894 (N_13894,N_13506,N_13723);
nand U13895 (N_13895,N_13758,N_13590);
nand U13896 (N_13896,N_13565,N_13542);
or U13897 (N_13897,N_13703,N_13761);
xor U13898 (N_13898,N_13561,N_13573);
nor U13899 (N_13899,N_13558,N_13763);
xnor U13900 (N_13900,N_13528,N_13591);
and U13901 (N_13901,N_13700,N_13662);
nor U13902 (N_13902,N_13610,N_13762);
nand U13903 (N_13903,N_13760,N_13541);
or U13904 (N_13904,N_13693,N_13619);
or U13905 (N_13905,N_13664,N_13792);
nor U13906 (N_13906,N_13626,N_13512);
and U13907 (N_13907,N_13713,N_13522);
nor U13908 (N_13908,N_13705,N_13585);
nand U13909 (N_13909,N_13679,N_13582);
nand U13910 (N_13910,N_13777,N_13715);
nor U13911 (N_13911,N_13620,N_13773);
or U13912 (N_13912,N_13702,N_13625);
and U13913 (N_13913,N_13562,N_13780);
nor U13914 (N_13914,N_13677,N_13557);
or U13915 (N_13915,N_13782,N_13534);
and U13916 (N_13916,N_13799,N_13748);
and U13917 (N_13917,N_13583,N_13766);
xnor U13918 (N_13918,N_13622,N_13543);
and U13919 (N_13919,N_13555,N_13751);
nor U13920 (N_13920,N_13539,N_13737);
or U13921 (N_13921,N_13658,N_13774);
nand U13922 (N_13922,N_13794,N_13533);
and U13923 (N_13923,N_13500,N_13638);
nor U13924 (N_13924,N_13501,N_13781);
xor U13925 (N_13925,N_13587,N_13798);
xnor U13926 (N_13926,N_13597,N_13647);
or U13927 (N_13927,N_13680,N_13752);
or U13928 (N_13928,N_13688,N_13579);
xnor U13929 (N_13929,N_13716,N_13708);
nor U13930 (N_13930,N_13605,N_13544);
nand U13931 (N_13931,N_13580,N_13521);
and U13932 (N_13932,N_13684,N_13628);
xor U13933 (N_13933,N_13551,N_13749);
nor U13934 (N_13934,N_13603,N_13729);
nand U13935 (N_13935,N_13722,N_13740);
or U13936 (N_13936,N_13754,N_13510);
or U13937 (N_13937,N_13525,N_13650);
nand U13938 (N_13938,N_13683,N_13649);
nand U13939 (N_13939,N_13560,N_13577);
nor U13940 (N_13940,N_13764,N_13719);
or U13941 (N_13941,N_13566,N_13529);
nor U13942 (N_13942,N_13663,N_13607);
xor U13943 (N_13943,N_13704,N_13738);
xnor U13944 (N_13944,N_13572,N_13513);
and U13945 (N_13945,N_13532,N_13768);
nor U13946 (N_13946,N_13690,N_13659);
xor U13947 (N_13947,N_13779,N_13670);
or U13948 (N_13948,N_13744,N_13733);
nor U13949 (N_13949,N_13750,N_13726);
nor U13950 (N_13950,N_13686,N_13672);
xnor U13951 (N_13951,N_13534,N_13730);
nor U13952 (N_13952,N_13585,N_13569);
xnor U13953 (N_13953,N_13695,N_13636);
and U13954 (N_13954,N_13677,N_13613);
or U13955 (N_13955,N_13567,N_13737);
nor U13956 (N_13956,N_13737,N_13689);
or U13957 (N_13957,N_13626,N_13514);
and U13958 (N_13958,N_13736,N_13636);
or U13959 (N_13959,N_13642,N_13525);
and U13960 (N_13960,N_13558,N_13716);
xor U13961 (N_13961,N_13650,N_13658);
xor U13962 (N_13962,N_13771,N_13507);
nor U13963 (N_13963,N_13580,N_13622);
and U13964 (N_13964,N_13655,N_13579);
nand U13965 (N_13965,N_13656,N_13799);
xor U13966 (N_13966,N_13787,N_13565);
nand U13967 (N_13967,N_13760,N_13635);
or U13968 (N_13968,N_13524,N_13622);
nor U13969 (N_13969,N_13530,N_13766);
nor U13970 (N_13970,N_13634,N_13591);
nor U13971 (N_13971,N_13558,N_13575);
or U13972 (N_13972,N_13782,N_13590);
and U13973 (N_13973,N_13635,N_13708);
nor U13974 (N_13974,N_13725,N_13683);
or U13975 (N_13975,N_13700,N_13794);
nand U13976 (N_13976,N_13614,N_13555);
nand U13977 (N_13977,N_13681,N_13636);
or U13978 (N_13978,N_13594,N_13569);
and U13979 (N_13979,N_13692,N_13718);
or U13980 (N_13980,N_13514,N_13588);
xor U13981 (N_13981,N_13790,N_13737);
and U13982 (N_13982,N_13595,N_13700);
or U13983 (N_13983,N_13584,N_13531);
or U13984 (N_13984,N_13557,N_13706);
xor U13985 (N_13985,N_13680,N_13740);
xnor U13986 (N_13986,N_13700,N_13504);
xor U13987 (N_13987,N_13574,N_13627);
or U13988 (N_13988,N_13703,N_13671);
nor U13989 (N_13989,N_13711,N_13509);
and U13990 (N_13990,N_13560,N_13642);
xor U13991 (N_13991,N_13647,N_13650);
and U13992 (N_13992,N_13684,N_13511);
xor U13993 (N_13993,N_13705,N_13577);
nand U13994 (N_13994,N_13552,N_13754);
nand U13995 (N_13995,N_13595,N_13566);
and U13996 (N_13996,N_13584,N_13591);
and U13997 (N_13997,N_13624,N_13634);
nor U13998 (N_13998,N_13728,N_13780);
xor U13999 (N_13999,N_13775,N_13507);
nand U14000 (N_14000,N_13501,N_13612);
and U14001 (N_14001,N_13511,N_13555);
xnor U14002 (N_14002,N_13704,N_13703);
and U14003 (N_14003,N_13556,N_13641);
nand U14004 (N_14004,N_13789,N_13590);
xor U14005 (N_14005,N_13564,N_13713);
and U14006 (N_14006,N_13514,N_13786);
and U14007 (N_14007,N_13636,N_13509);
xor U14008 (N_14008,N_13720,N_13505);
nor U14009 (N_14009,N_13760,N_13701);
nand U14010 (N_14010,N_13591,N_13657);
nand U14011 (N_14011,N_13736,N_13575);
or U14012 (N_14012,N_13733,N_13648);
nand U14013 (N_14013,N_13628,N_13626);
nand U14014 (N_14014,N_13669,N_13647);
nor U14015 (N_14015,N_13682,N_13725);
and U14016 (N_14016,N_13524,N_13501);
or U14017 (N_14017,N_13791,N_13582);
nor U14018 (N_14018,N_13796,N_13791);
and U14019 (N_14019,N_13711,N_13550);
xnor U14020 (N_14020,N_13633,N_13650);
nor U14021 (N_14021,N_13778,N_13652);
nor U14022 (N_14022,N_13635,N_13552);
or U14023 (N_14023,N_13500,N_13799);
or U14024 (N_14024,N_13723,N_13599);
and U14025 (N_14025,N_13536,N_13669);
and U14026 (N_14026,N_13596,N_13505);
or U14027 (N_14027,N_13741,N_13708);
nor U14028 (N_14028,N_13723,N_13654);
and U14029 (N_14029,N_13632,N_13574);
xor U14030 (N_14030,N_13753,N_13648);
nor U14031 (N_14031,N_13580,N_13601);
nor U14032 (N_14032,N_13547,N_13741);
nor U14033 (N_14033,N_13601,N_13793);
and U14034 (N_14034,N_13600,N_13697);
xnor U14035 (N_14035,N_13625,N_13674);
nand U14036 (N_14036,N_13685,N_13656);
or U14037 (N_14037,N_13594,N_13652);
xor U14038 (N_14038,N_13618,N_13537);
nor U14039 (N_14039,N_13545,N_13527);
nor U14040 (N_14040,N_13749,N_13784);
and U14041 (N_14041,N_13566,N_13775);
nand U14042 (N_14042,N_13531,N_13503);
or U14043 (N_14043,N_13719,N_13704);
xor U14044 (N_14044,N_13608,N_13618);
nand U14045 (N_14045,N_13512,N_13771);
or U14046 (N_14046,N_13647,N_13626);
and U14047 (N_14047,N_13719,N_13614);
and U14048 (N_14048,N_13747,N_13714);
or U14049 (N_14049,N_13624,N_13543);
nand U14050 (N_14050,N_13655,N_13718);
xor U14051 (N_14051,N_13733,N_13741);
xor U14052 (N_14052,N_13739,N_13680);
xnor U14053 (N_14053,N_13784,N_13709);
nand U14054 (N_14054,N_13631,N_13644);
and U14055 (N_14055,N_13663,N_13700);
nor U14056 (N_14056,N_13572,N_13691);
nand U14057 (N_14057,N_13525,N_13714);
nand U14058 (N_14058,N_13523,N_13542);
nand U14059 (N_14059,N_13698,N_13763);
or U14060 (N_14060,N_13724,N_13694);
nor U14061 (N_14061,N_13519,N_13654);
or U14062 (N_14062,N_13584,N_13665);
and U14063 (N_14063,N_13633,N_13554);
xnor U14064 (N_14064,N_13724,N_13645);
nand U14065 (N_14065,N_13628,N_13748);
and U14066 (N_14066,N_13662,N_13611);
and U14067 (N_14067,N_13639,N_13652);
nand U14068 (N_14068,N_13503,N_13659);
xnor U14069 (N_14069,N_13659,N_13738);
xnor U14070 (N_14070,N_13736,N_13797);
or U14071 (N_14071,N_13670,N_13529);
nor U14072 (N_14072,N_13677,N_13662);
xor U14073 (N_14073,N_13799,N_13571);
xnor U14074 (N_14074,N_13768,N_13573);
and U14075 (N_14075,N_13668,N_13572);
nand U14076 (N_14076,N_13741,N_13512);
nand U14077 (N_14077,N_13516,N_13726);
nor U14078 (N_14078,N_13706,N_13609);
and U14079 (N_14079,N_13501,N_13613);
or U14080 (N_14080,N_13667,N_13761);
nand U14081 (N_14081,N_13587,N_13633);
and U14082 (N_14082,N_13581,N_13529);
nor U14083 (N_14083,N_13731,N_13697);
xnor U14084 (N_14084,N_13658,N_13684);
or U14085 (N_14085,N_13723,N_13519);
and U14086 (N_14086,N_13580,N_13699);
nor U14087 (N_14087,N_13539,N_13561);
nand U14088 (N_14088,N_13721,N_13774);
xor U14089 (N_14089,N_13757,N_13615);
nand U14090 (N_14090,N_13558,N_13519);
xnor U14091 (N_14091,N_13683,N_13563);
and U14092 (N_14092,N_13717,N_13532);
nor U14093 (N_14093,N_13588,N_13512);
xnor U14094 (N_14094,N_13523,N_13688);
nor U14095 (N_14095,N_13795,N_13683);
nor U14096 (N_14096,N_13661,N_13598);
or U14097 (N_14097,N_13540,N_13674);
xor U14098 (N_14098,N_13787,N_13697);
xnor U14099 (N_14099,N_13642,N_13582);
nor U14100 (N_14100,N_13806,N_13977);
nand U14101 (N_14101,N_13884,N_14058);
xor U14102 (N_14102,N_14086,N_13991);
xor U14103 (N_14103,N_13925,N_14061);
or U14104 (N_14104,N_13869,N_13932);
nand U14105 (N_14105,N_13910,N_13909);
or U14106 (N_14106,N_13996,N_13994);
nand U14107 (N_14107,N_13985,N_13947);
or U14108 (N_14108,N_14006,N_13978);
nand U14109 (N_14109,N_13864,N_13907);
nor U14110 (N_14110,N_13923,N_13815);
nor U14111 (N_14111,N_13810,N_13883);
nand U14112 (N_14112,N_14062,N_14011);
and U14113 (N_14113,N_14002,N_14096);
nor U14114 (N_14114,N_14083,N_14097);
nand U14115 (N_14115,N_13847,N_14005);
and U14116 (N_14116,N_13916,N_13971);
nor U14117 (N_14117,N_14081,N_13873);
or U14118 (N_14118,N_13837,N_13899);
nand U14119 (N_14119,N_13999,N_14009);
and U14120 (N_14120,N_14000,N_14048);
and U14121 (N_14121,N_13803,N_13993);
xor U14122 (N_14122,N_13877,N_13868);
and U14123 (N_14123,N_13963,N_13912);
xnor U14124 (N_14124,N_13861,N_14050);
or U14125 (N_14125,N_13872,N_13965);
or U14126 (N_14126,N_13862,N_13974);
nand U14127 (N_14127,N_13855,N_13967);
xor U14128 (N_14128,N_14090,N_13885);
nor U14129 (N_14129,N_13905,N_14026);
xor U14130 (N_14130,N_14051,N_13992);
or U14131 (N_14131,N_14021,N_14037);
nor U14132 (N_14132,N_13843,N_14041);
nand U14133 (N_14133,N_13809,N_13856);
or U14134 (N_14134,N_14091,N_13858);
or U14135 (N_14135,N_13957,N_13964);
and U14136 (N_14136,N_13900,N_14013);
nor U14137 (N_14137,N_13898,N_13857);
xnor U14138 (N_14138,N_13920,N_14035);
and U14139 (N_14139,N_14063,N_13969);
nor U14140 (N_14140,N_13807,N_13878);
nor U14141 (N_14141,N_13943,N_13874);
xor U14142 (N_14142,N_13976,N_14018);
or U14143 (N_14143,N_14049,N_13834);
nor U14144 (N_14144,N_14023,N_14004);
nor U14145 (N_14145,N_14092,N_14071);
and U14146 (N_14146,N_13933,N_13917);
or U14147 (N_14147,N_13921,N_13828);
or U14148 (N_14148,N_13879,N_13995);
and U14149 (N_14149,N_14008,N_13846);
nand U14150 (N_14150,N_13959,N_13998);
or U14151 (N_14151,N_13987,N_14070);
or U14152 (N_14152,N_14019,N_13984);
xor U14153 (N_14153,N_13887,N_13913);
nor U14154 (N_14154,N_13990,N_14066);
xor U14155 (N_14155,N_14068,N_13821);
nand U14156 (N_14156,N_13801,N_14017);
xnor U14157 (N_14157,N_13922,N_14059);
and U14158 (N_14158,N_14082,N_13951);
nand U14159 (N_14159,N_14088,N_14085);
xnor U14160 (N_14160,N_13931,N_13825);
xor U14161 (N_14161,N_13863,N_13918);
nand U14162 (N_14162,N_13940,N_14015);
or U14163 (N_14163,N_13935,N_13818);
xnor U14164 (N_14164,N_13832,N_13948);
and U14165 (N_14165,N_13852,N_14045);
nor U14166 (N_14166,N_13954,N_13934);
nor U14167 (N_14167,N_13839,N_14056);
nand U14168 (N_14168,N_13961,N_14094);
and U14169 (N_14169,N_14042,N_13880);
nand U14170 (N_14170,N_14001,N_13953);
nor U14171 (N_14171,N_13930,N_14076);
or U14172 (N_14172,N_13911,N_13929);
xnor U14173 (N_14173,N_13890,N_13891);
nor U14174 (N_14174,N_13894,N_13928);
and U14175 (N_14175,N_14078,N_13986);
nor U14176 (N_14176,N_13981,N_13804);
xor U14177 (N_14177,N_14034,N_13893);
or U14178 (N_14178,N_13860,N_13886);
xor U14179 (N_14179,N_14089,N_13819);
nand U14180 (N_14180,N_14024,N_14020);
and U14181 (N_14181,N_13897,N_13823);
nor U14182 (N_14182,N_14069,N_13870);
xor U14183 (N_14183,N_13972,N_14079);
xor U14184 (N_14184,N_14014,N_13827);
nand U14185 (N_14185,N_14007,N_14046);
nor U14186 (N_14186,N_13853,N_13975);
and U14187 (N_14187,N_13849,N_13896);
nand U14188 (N_14188,N_14038,N_14003);
or U14189 (N_14189,N_13973,N_13830);
and U14190 (N_14190,N_13835,N_14072);
or U14191 (N_14191,N_14044,N_13808);
nand U14192 (N_14192,N_13939,N_13958);
nor U14193 (N_14193,N_14029,N_13942);
and U14194 (N_14194,N_13966,N_13908);
nand U14195 (N_14195,N_13926,N_14077);
xor U14196 (N_14196,N_13840,N_13914);
or U14197 (N_14197,N_13941,N_14025);
xor U14198 (N_14198,N_13968,N_13902);
nor U14199 (N_14199,N_13842,N_14099);
nor U14200 (N_14200,N_14073,N_13816);
nand U14201 (N_14201,N_13824,N_13871);
and U14202 (N_14202,N_14016,N_13812);
or U14203 (N_14203,N_13983,N_13820);
and U14204 (N_14204,N_13945,N_13875);
nor U14205 (N_14205,N_13892,N_13927);
xor U14206 (N_14206,N_13826,N_13980);
xnor U14207 (N_14207,N_14040,N_14093);
nor U14208 (N_14208,N_13854,N_13850);
nand U14209 (N_14209,N_14039,N_14074);
nand U14210 (N_14210,N_13989,N_13988);
nor U14211 (N_14211,N_13924,N_13829);
xnor U14212 (N_14212,N_14031,N_14036);
nor U14213 (N_14213,N_13936,N_13946);
nand U14214 (N_14214,N_13836,N_13848);
nor U14215 (N_14215,N_14028,N_14054);
xor U14216 (N_14216,N_14012,N_13915);
and U14217 (N_14217,N_13960,N_14065);
or U14218 (N_14218,N_13802,N_14064);
and U14219 (N_14219,N_14057,N_13889);
xnor U14220 (N_14220,N_14087,N_13950);
nor U14221 (N_14221,N_13814,N_13895);
nand U14222 (N_14222,N_13956,N_13805);
and U14223 (N_14223,N_13970,N_13876);
xnor U14224 (N_14224,N_13838,N_13903);
and U14225 (N_14225,N_13952,N_13904);
and U14226 (N_14226,N_13962,N_13882);
xnor U14227 (N_14227,N_13944,N_13949);
xor U14228 (N_14228,N_14030,N_13851);
xnor U14229 (N_14229,N_14053,N_13938);
xnor U14230 (N_14230,N_13844,N_13997);
nor U14231 (N_14231,N_13955,N_14027);
nand U14232 (N_14232,N_14022,N_14075);
nand U14233 (N_14233,N_13901,N_14095);
and U14234 (N_14234,N_13822,N_13865);
xnor U14235 (N_14235,N_13866,N_13831);
xnor U14236 (N_14236,N_14098,N_13979);
xnor U14237 (N_14237,N_13881,N_14060);
nand U14238 (N_14238,N_13906,N_13859);
or U14239 (N_14239,N_13845,N_13867);
and U14240 (N_14240,N_13817,N_14047);
xnor U14241 (N_14241,N_14032,N_13982);
nand U14242 (N_14242,N_13811,N_13813);
and U14243 (N_14243,N_14033,N_13800);
and U14244 (N_14244,N_14010,N_14084);
nand U14245 (N_14245,N_13937,N_13888);
nor U14246 (N_14246,N_13841,N_13833);
xnor U14247 (N_14247,N_14067,N_14055);
nor U14248 (N_14248,N_13919,N_14052);
nand U14249 (N_14249,N_14043,N_14080);
xnor U14250 (N_14250,N_13831,N_13845);
nand U14251 (N_14251,N_13868,N_14051);
nor U14252 (N_14252,N_14067,N_13882);
or U14253 (N_14253,N_13829,N_14066);
nor U14254 (N_14254,N_13961,N_13958);
and U14255 (N_14255,N_14015,N_14053);
nor U14256 (N_14256,N_13823,N_14091);
and U14257 (N_14257,N_13825,N_13878);
nand U14258 (N_14258,N_14015,N_13870);
xnor U14259 (N_14259,N_13976,N_13891);
nand U14260 (N_14260,N_13852,N_14073);
or U14261 (N_14261,N_14098,N_13864);
xnor U14262 (N_14262,N_14082,N_13974);
nor U14263 (N_14263,N_13970,N_14074);
xor U14264 (N_14264,N_13863,N_14021);
and U14265 (N_14265,N_13970,N_13943);
xnor U14266 (N_14266,N_13835,N_14027);
nand U14267 (N_14267,N_13858,N_13880);
xnor U14268 (N_14268,N_13933,N_14036);
nor U14269 (N_14269,N_13825,N_13868);
nand U14270 (N_14270,N_13826,N_14060);
nor U14271 (N_14271,N_13885,N_13969);
and U14272 (N_14272,N_13902,N_14097);
nor U14273 (N_14273,N_13889,N_14016);
and U14274 (N_14274,N_14076,N_14033);
xnor U14275 (N_14275,N_13995,N_13949);
nand U14276 (N_14276,N_13834,N_14035);
and U14277 (N_14277,N_13919,N_13955);
and U14278 (N_14278,N_14062,N_13870);
nand U14279 (N_14279,N_14089,N_13858);
nand U14280 (N_14280,N_13879,N_13910);
and U14281 (N_14281,N_14047,N_14036);
xor U14282 (N_14282,N_13949,N_13828);
and U14283 (N_14283,N_13962,N_13849);
nand U14284 (N_14284,N_13867,N_13954);
xor U14285 (N_14285,N_14011,N_13843);
or U14286 (N_14286,N_13827,N_13900);
xnor U14287 (N_14287,N_13957,N_14062);
nor U14288 (N_14288,N_13999,N_13803);
and U14289 (N_14289,N_13838,N_13973);
or U14290 (N_14290,N_13886,N_14086);
or U14291 (N_14291,N_13854,N_13960);
xnor U14292 (N_14292,N_14052,N_14019);
and U14293 (N_14293,N_14037,N_13959);
or U14294 (N_14294,N_13982,N_13861);
and U14295 (N_14295,N_13807,N_13983);
or U14296 (N_14296,N_13853,N_13885);
xor U14297 (N_14297,N_13858,N_13851);
nor U14298 (N_14298,N_13899,N_13869);
and U14299 (N_14299,N_13808,N_14084);
nand U14300 (N_14300,N_13894,N_14013);
nand U14301 (N_14301,N_13964,N_14003);
xor U14302 (N_14302,N_13846,N_13887);
or U14303 (N_14303,N_13950,N_13866);
or U14304 (N_14304,N_13915,N_13852);
nand U14305 (N_14305,N_14077,N_13933);
xor U14306 (N_14306,N_13962,N_13831);
or U14307 (N_14307,N_13826,N_14079);
xnor U14308 (N_14308,N_14054,N_13917);
nand U14309 (N_14309,N_13939,N_14052);
or U14310 (N_14310,N_13895,N_14026);
xor U14311 (N_14311,N_14033,N_13842);
xnor U14312 (N_14312,N_14071,N_14043);
nand U14313 (N_14313,N_14082,N_13925);
xnor U14314 (N_14314,N_13846,N_14062);
and U14315 (N_14315,N_13972,N_14069);
and U14316 (N_14316,N_13869,N_14053);
or U14317 (N_14317,N_14072,N_13894);
or U14318 (N_14318,N_14006,N_13827);
or U14319 (N_14319,N_14077,N_13972);
nor U14320 (N_14320,N_13953,N_13983);
xor U14321 (N_14321,N_13935,N_13862);
nor U14322 (N_14322,N_14044,N_14094);
and U14323 (N_14323,N_14097,N_14043);
nor U14324 (N_14324,N_14095,N_13953);
and U14325 (N_14325,N_13918,N_14005);
nor U14326 (N_14326,N_13955,N_13862);
or U14327 (N_14327,N_13801,N_13904);
nand U14328 (N_14328,N_13966,N_13853);
and U14329 (N_14329,N_14091,N_13978);
nor U14330 (N_14330,N_13813,N_13953);
nor U14331 (N_14331,N_14042,N_13855);
and U14332 (N_14332,N_13857,N_14042);
xnor U14333 (N_14333,N_13809,N_14067);
or U14334 (N_14334,N_14036,N_14086);
and U14335 (N_14335,N_14094,N_13983);
and U14336 (N_14336,N_13822,N_14054);
nand U14337 (N_14337,N_14087,N_13848);
or U14338 (N_14338,N_13942,N_13804);
xnor U14339 (N_14339,N_13854,N_13979);
nand U14340 (N_14340,N_13894,N_13979);
nor U14341 (N_14341,N_13859,N_13905);
and U14342 (N_14342,N_13888,N_14023);
nor U14343 (N_14343,N_14076,N_14005);
or U14344 (N_14344,N_13899,N_13931);
xor U14345 (N_14345,N_13833,N_14093);
or U14346 (N_14346,N_13973,N_13923);
nand U14347 (N_14347,N_13912,N_14007);
nor U14348 (N_14348,N_13845,N_13932);
and U14349 (N_14349,N_14081,N_14048);
nand U14350 (N_14350,N_13898,N_13931);
nor U14351 (N_14351,N_13852,N_13986);
and U14352 (N_14352,N_14009,N_14072);
nor U14353 (N_14353,N_13909,N_13941);
or U14354 (N_14354,N_13976,N_13861);
nand U14355 (N_14355,N_13956,N_14019);
nor U14356 (N_14356,N_14093,N_13982);
and U14357 (N_14357,N_13988,N_13981);
nor U14358 (N_14358,N_13937,N_13850);
xor U14359 (N_14359,N_14058,N_13971);
xor U14360 (N_14360,N_13820,N_13980);
and U14361 (N_14361,N_14084,N_14025);
and U14362 (N_14362,N_13842,N_14039);
nand U14363 (N_14363,N_14094,N_13838);
nand U14364 (N_14364,N_14080,N_13870);
xnor U14365 (N_14365,N_13918,N_13964);
xnor U14366 (N_14366,N_13967,N_13862);
xnor U14367 (N_14367,N_14029,N_14050);
nand U14368 (N_14368,N_13898,N_13813);
nand U14369 (N_14369,N_14055,N_13980);
nand U14370 (N_14370,N_13803,N_13896);
xnor U14371 (N_14371,N_13935,N_13821);
xor U14372 (N_14372,N_13966,N_13920);
nor U14373 (N_14373,N_14048,N_14008);
and U14374 (N_14374,N_14053,N_13855);
nor U14375 (N_14375,N_13829,N_14014);
xor U14376 (N_14376,N_13962,N_14042);
nor U14377 (N_14377,N_14010,N_13820);
and U14378 (N_14378,N_14004,N_14073);
or U14379 (N_14379,N_13894,N_13934);
nor U14380 (N_14380,N_13836,N_13961);
nor U14381 (N_14381,N_14022,N_13887);
nand U14382 (N_14382,N_13841,N_13984);
nor U14383 (N_14383,N_14030,N_14049);
xor U14384 (N_14384,N_13807,N_13870);
xnor U14385 (N_14385,N_13931,N_14031);
nor U14386 (N_14386,N_13936,N_13928);
nand U14387 (N_14387,N_14094,N_13812);
nor U14388 (N_14388,N_13835,N_13848);
or U14389 (N_14389,N_14089,N_14006);
xor U14390 (N_14390,N_13814,N_13952);
nor U14391 (N_14391,N_14001,N_13883);
nor U14392 (N_14392,N_13922,N_13900);
xnor U14393 (N_14393,N_13830,N_13839);
nor U14394 (N_14394,N_13928,N_13802);
xnor U14395 (N_14395,N_14089,N_13904);
nand U14396 (N_14396,N_13851,N_14074);
or U14397 (N_14397,N_14019,N_13888);
xor U14398 (N_14398,N_13942,N_13833);
nor U14399 (N_14399,N_13963,N_13995);
or U14400 (N_14400,N_14303,N_14201);
and U14401 (N_14401,N_14345,N_14323);
and U14402 (N_14402,N_14300,N_14392);
and U14403 (N_14403,N_14151,N_14289);
or U14404 (N_14404,N_14282,N_14257);
xor U14405 (N_14405,N_14301,N_14391);
xor U14406 (N_14406,N_14179,N_14143);
nor U14407 (N_14407,N_14157,N_14125);
or U14408 (N_14408,N_14173,N_14209);
nand U14409 (N_14409,N_14131,N_14297);
xor U14410 (N_14410,N_14255,N_14163);
and U14411 (N_14411,N_14230,N_14160);
nand U14412 (N_14412,N_14393,N_14336);
or U14413 (N_14413,N_14350,N_14141);
nand U14414 (N_14414,N_14318,N_14217);
nand U14415 (N_14415,N_14295,N_14384);
and U14416 (N_14416,N_14137,N_14315);
nor U14417 (N_14417,N_14377,N_14103);
or U14418 (N_14418,N_14106,N_14104);
nor U14419 (N_14419,N_14369,N_14351);
nand U14420 (N_14420,N_14197,N_14145);
and U14421 (N_14421,N_14365,N_14130);
and U14422 (N_14422,N_14328,N_14200);
xnor U14423 (N_14423,N_14340,N_14321);
nor U14424 (N_14424,N_14308,N_14208);
xnor U14425 (N_14425,N_14198,N_14113);
and U14426 (N_14426,N_14362,N_14235);
and U14427 (N_14427,N_14107,N_14155);
xor U14428 (N_14428,N_14119,N_14266);
xor U14429 (N_14429,N_14372,N_14238);
xnor U14430 (N_14430,N_14140,N_14371);
and U14431 (N_14431,N_14128,N_14100);
and U14432 (N_14432,N_14139,N_14211);
nand U14433 (N_14433,N_14376,N_14383);
or U14434 (N_14434,N_14256,N_14136);
xor U14435 (N_14435,N_14379,N_14178);
or U14436 (N_14436,N_14247,N_14364);
xor U14437 (N_14437,N_14135,N_14373);
and U14438 (N_14438,N_14316,N_14156);
and U14439 (N_14439,N_14150,N_14286);
and U14440 (N_14440,N_14176,N_14356);
nand U14441 (N_14441,N_14284,N_14341);
nand U14442 (N_14442,N_14293,N_14149);
and U14443 (N_14443,N_14306,N_14196);
nand U14444 (N_14444,N_14213,N_14395);
or U14445 (N_14445,N_14382,N_14359);
and U14446 (N_14446,N_14352,N_14326);
xor U14447 (N_14447,N_14348,N_14398);
nand U14448 (N_14448,N_14220,N_14115);
nand U14449 (N_14449,N_14245,N_14342);
and U14450 (N_14450,N_14271,N_14314);
nand U14451 (N_14451,N_14317,N_14357);
nor U14452 (N_14452,N_14162,N_14154);
xnor U14453 (N_14453,N_14127,N_14361);
xor U14454 (N_14454,N_14267,N_14338);
and U14455 (N_14455,N_14210,N_14216);
or U14456 (N_14456,N_14347,N_14223);
nor U14457 (N_14457,N_14294,N_14368);
and U14458 (N_14458,N_14184,N_14299);
xnor U14459 (N_14459,N_14152,N_14388);
nand U14460 (N_14460,N_14132,N_14389);
xor U14461 (N_14461,N_14174,N_14307);
xnor U14462 (N_14462,N_14202,N_14385);
nor U14463 (N_14463,N_14126,N_14269);
nand U14464 (N_14464,N_14262,N_14204);
nand U14465 (N_14465,N_14112,N_14225);
xnor U14466 (N_14466,N_14214,N_14167);
nor U14467 (N_14467,N_14311,N_14146);
nor U14468 (N_14468,N_14329,N_14183);
and U14469 (N_14469,N_14124,N_14142);
nor U14470 (N_14470,N_14190,N_14349);
xor U14471 (N_14471,N_14337,N_14195);
and U14472 (N_14472,N_14310,N_14397);
or U14473 (N_14473,N_14360,N_14122);
nor U14474 (N_14474,N_14370,N_14250);
nor U14475 (N_14475,N_14305,N_14165);
or U14476 (N_14476,N_14153,N_14285);
nor U14477 (N_14477,N_14144,N_14258);
or U14478 (N_14478,N_14275,N_14324);
nor U14479 (N_14479,N_14171,N_14319);
xor U14480 (N_14480,N_14327,N_14380);
and U14481 (N_14481,N_14229,N_14236);
and U14482 (N_14482,N_14191,N_14253);
nor U14483 (N_14483,N_14320,N_14203);
and U14484 (N_14484,N_14386,N_14194);
xnor U14485 (N_14485,N_14313,N_14281);
xor U14486 (N_14486,N_14358,N_14292);
nand U14487 (N_14487,N_14374,N_14298);
or U14488 (N_14488,N_14353,N_14366);
or U14489 (N_14489,N_14123,N_14231);
and U14490 (N_14490,N_14354,N_14312);
and U14491 (N_14491,N_14187,N_14218);
nor U14492 (N_14492,N_14239,N_14287);
nand U14493 (N_14493,N_14120,N_14164);
or U14494 (N_14494,N_14277,N_14181);
nand U14495 (N_14495,N_14261,N_14346);
nand U14496 (N_14496,N_14134,N_14116);
and U14497 (N_14497,N_14108,N_14322);
nand U14498 (N_14498,N_14330,N_14110);
nor U14499 (N_14499,N_14268,N_14182);
and U14500 (N_14500,N_14193,N_14249);
nor U14501 (N_14501,N_14233,N_14159);
or U14502 (N_14502,N_14263,N_14279);
nand U14503 (N_14503,N_14309,N_14188);
and U14504 (N_14504,N_14206,N_14363);
and U14505 (N_14505,N_14222,N_14212);
xnor U14506 (N_14506,N_14207,N_14175);
xnor U14507 (N_14507,N_14215,N_14117);
or U14508 (N_14508,N_14332,N_14280);
nand U14509 (N_14509,N_14274,N_14259);
nand U14510 (N_14510,N_14399,N_14367);
or U14511 (N_14511,N_14335,N_14265);
nand U14512 (N_14512,N_14290,N_14390);
nor U14513 (N_14513,N_14260,N_14224);
nor U14514 (N_14514,N_14227,N_14381);
and U14515 (N_14515,N_14147,N_14180);
nand U14516 (N_14516,N_14304,N_14242);
and U14517 (N_14517,N_14355,N_14270);
and U14518 (N_14518,N_14278,N_14254);
nand U14519 (N_14519,N_14387,N_14221);
nand U14520 (N_14520,N_14378,N_14232);
nand U14521 (N_14521,N_14168,N_14252);
or U14522 (N_14522,N_14189,N_14251);
nand U14523 (N_14523,N_14331,N_14291);
nand U14524 (N_14524,N_14343,N_14283);
xnor U14525 (N_14525,N_14240,N_14186);
or U14526 (N_14526,N_14166,N_14272);
and U14527 (N_14527,N_14264,N_14101);
nand U14528 (N_14528,N_14161,N_14118);
or U14529 (N_14529,N_14333,N_14396);
nor U14530 (N_14530,N_14185,N_14114);
or U14531 (N_14531,N_14339,N_14288);
or U14532 (N_14532,N_14102,N_14158);
xnor U14533 (N_14533,N_14172,N_14244);
xnor U14534 (N_14534,N_14170,N_14138);
nand U14535 (N_14535,N_14296,N_14121);
nor U14536 (N_14536,N_14234,N_14219);
and U14537 (N_14537,N_14109,N_14334);
xor U14538 (N_14538,N_14325,N_14246);
nor U14539 (N_14539,N_14302,N_14241);
or U14540 (N_14540,N_14248,N_14105);
or U14541 (N_14541,N_14192,N_14226);
and U14542 (N_14542,N_14375,N_14199);
or U14543 (N_14543,N_14276,N_14177);
nand U14544 (N_14544,N_14205,N_14169);
or U14545 (N_14545,N_14243,N_14237);
nor U14546 (N_14546,N_14133,N_14344);
nor U14547 (N_14547,N_14394,N_14228);
xor U14548 (N_14548,N_14129,N_14273);
or U14549 (N_14549,N_14111,N_14148);
and U14550 (N_14550,N_14342,N_14322);
nor U14551 (N_14551,N_14113,N_14246);
nor U14552 (N_14552,N_14187,N_14131);
xor U14553 (N_14553,N_14241,N_14184);
xnor U14554 (N_14554,N_14274,N_14104);
nor U14555 (N_14555,N_14212,N_14193);
or U14556 (N_14556,N_14358,N_14222);
xor U14557 (N_14557,N_14242,N_14303);
or U14558 (N_14558,N_14126,N_14227);
nand U14559 (N_14559,N_14205,N_14353);
and U14560 (N_14560,N_14389,N_14322);
or U14561 (N_14561,N_14105,N_14273);
nor U14562 (N_14562,N_14152,N_14216);
xor U14563 (N_14563,N_14211,N_14353);
nand U14564 (N_14564,N_14381,N_14286);
and U14565 (N_14565,N_14230,N_14185);
xor U14566 (N_14566,N_14182,N_14359);
xnor U14567 (N_14567,N_14223,N_14371);
and U14568 (N_14568,N_14140,N_14354);
and U14569 (N_14569,N_14113,N_14295);
nand U14570 (N_14570,N_14275,N_14121);
nor U14571 (N_14571,N_14141,N_14116);
and U14572 (N_14572,N_14316,N_14349);
nand U14573 (N_14573,N_14233,N_14366);
or U14574 (N_14574,N_14295,N_14348);
nor U14575 (N_14575,N_14214,N_14384);
or U14576 (N_14576,N_14148,N_14193);
xnor U14577 (N_14577,N_14333,N_14367);
or U14578 (N_14578,N_14106,N_14318);
xor U14579 (N_14579,N_14299,N_14394);
and U14580 (N_14580,N_14154,N_14260);
nand U14581 (N_14581,N_14239,N_14348);
xor U14582 (N_14582,N_14280,N_14310);
nor U14583 (N_14583,N_14160,N_14154);
xor U14584 (N_14584,N_14296,N_14342);
xor U14585 (N_14585,N_14207,N_14262);
or U14586 (N_14586,N_14378,N_14145);
xor U14587 (N_14587,N_14314,N_14359);
nor U14588 (N_14588,N_14345,N_14396);
xnor U14589 (N_14589,N_14358,N_14207);
or U14590 (N_14590,N_14217,N_14105);
xnor U14591 (N_14591,N_14216,N_14119);
xor U14592 (N_14592,N_14219,N_14252);
nand U14593 (N_14593,N_14280,N_14276);
nor U14594 (N_14594,N_14273,N_14332);
nor U14595 (N_14595,N_14336,N_14157);
and U14596 (N_14596,N_14198,N_14333);
xor U14597 (N_14597,N_14232,N_14191);
nor U14598 (N_14598,N_14198,N_14169);
nor U14599 (N_14599,N_14290,N_14348);
nand U14600 (N_14600,N_14398,N_14313);
xnor U14601 (N_14601,N_14166,N_14243);
nor U14602 (N_14602,N_14245,N_14248);
xnor U14603 (N_14603,N_14288,N_14114);
or U14604 (N_14604,N_14281,N_14243);
nand U14605 (N_14605,N_14284,N_14192);
nand U14606 (N_14606,N_14318,N_14293);
nand U14607 (N_14607,N_14281,N_14181);
nand U14608 (N_14608,N_14132,N_14278);
xor U14609 (N_14609,N_14103,N_14357);
or U14610 (N_14610,N_14260,N_14243);
nand U14611 (N_14611,N_14192,N_14313);
or U14612 (N_14612,N_14230,N_14303);
xor U14613 (N_14613,N_14194,N_14284);
xnor U14614 (N_14614,N_14193,N_14351);
xor U14615 (N_14615,N_14327,N_14108);
and U14616 (N_14616,N_14303,N_14266);
nor U14617 (N_14617,N_14396,N_14227);
and U14618 (N_14618,N_14305,N_14258);
nor U14619 (N_14619,N_14368,N_14394);
xnor U14620 (N_14620,N_14355,N_14289);
nor U14621 (N_14621,N_14134,N_14354);
and U14622 (N_14622,N_14316,N_14343);
nor U14623 (N_14623,N_14146,N_14159);
or U14624 (N_14624,N_14162,N_14275);
nor U14625 (N_14625,N_14118,N_14215);
nor U14626 (N_14626,N_14205,N_14184);
nand U14627 (N_14627,N_14140,N_14138);
nand U14628 (N_14628,N_14173,N_14385);
xnor U14629 (N_14629,N_14264,N_14230);
nand U14630 (N_14630,N_14250,N_14117);
or U14631 (N_14631,N_14126,N_14200);
nand U14632 (N_14632,N_14382,N_14209);
or U14633 (N_14633,N_14344,N_14179);
xnor U14634 (N_14634,N_14382,N_14341);
or U14635 (N_14635,N_14202,N_14118);
or U14636 (N_14636,N_14211,N_14382);
xor U14637 (N_14637,N_14149,N_14127);
nor U14638 (N_14638,N_14302,N_14364);
nand U14639 (N_14639,N_14304,N_14312);
xor U14640 (N_14640,N_14354,N_14125);
xor U14641 (N_14641,N_14375,N_14368);
or U14642 (N_14642,N_14254,N_14326);
and U14643 (N_14643,N_14141,N_14240);
nand U14644 (N_14644,N_14385,N_14392);
xnor U14645 (N_14645,N_14179,N_14199);
xnor U14646 (N_14646,N_14281,N_14299);
and U14647 (N_14647,N_14171,N_14285);
or U14648 (N_14648,N_14343,N_14166);
nand U14649 (N_14649,N_14317,N_14140);
and U14650 (N_14650,N_14287,N_14393);
nor U14651 (N_14651,N_14160,N_14305);
and U14652 (N_14652,N_14278,N_14317);
or U14653 (N_14653,N_14152,N_14235);
xor U14654 (N_14654,N_14301,N_14134);
and U14655 (N_14655,N_14301,N_14378);
nor U14656 (N_14656,N_14381,N_14155);
or U14657 (N_14657,N_14255,N_14136);
nand U14658 (N_14658,N_14188,N_14294);
and U14659 (N_14659,N_14322,N_14134);
nand U14660 (N_14660,N_14303,N_14392);
xnor U14661 (N_14661,N_14285,N_14119);
nand U14662 (N_14662,N_14397,N_14101);
nor U14663 (N_14663,N_14317,N_14109);
xnor U14664 (N_14664,N_14254,N_14101);
nand U14665 (N_14665,N_14258,N_14213);
nand U14666 (N_14666,N_14102,N_14217);
xnor U14667 (N_14667,N_14299,N_14130);
xnor U14668 (N_14668,N_14111,N_14339);
nor U14669 (N_14669,N_14139,N_14275);
or U14670 (N_14670,N_14216,N_14103);
xor U14671 (N_14671,N_14199,N_14268);
or U14672 (N_14672,N_14247,N_14179);
nand U14673 (N_14673,N_14177,N_14118);
xnor U14674 (N_14674,N_14271,N_14122);
nand U14675 (N_14675,N_14189,N_14207);
xor U14676 (N_14676,N_14110,N_14342);
xnor U14677 (N_14677,N_14375,N_14124);
xor U14678 (N_14678,N_14108,N_14398);
xor U14679 (N_14679,N_14132,N_14323);
and U14680 (N_14680,N_14305,N_14156);
xnor U14681 (N_14681,N_14377,N_14352);
nor U14682 (N_14682,N_14332,N_14260);
or U14683 (N_14683,N_14389,N_14145);
and U14684 (N_14684,N_14231,N_14357);
nor U14685 (N_14685,N_14290,N_14272);
and U14686 (N_14686,N_14243,N_14391);
nand U14687 (N_14687,N_14241,N_14263);
xor U14688 (N_14688,N_14245,N_14322);
nand U14689 (N_14689,N_14236,N_14396);
or U14690 (N_14690,N_14372,N_14230);
and U14691 (N_14691,N_14103,N_14281);
or U14692 (N_14692,N_14316,N_14190);
nand U14693 (N_14693,N_14328,N_14284);
nor U14694 (N_14694,N_14366,N_14158);
or U14695 (N_14695,N_14369,N_14262);
and U14696 (N_14696,N_14311,N_14264);
or U14697 (N_14697,N_14116,N_14243);
nor U14698 (N_14698,N_14259,N_14148);
nand U14699 (N_14699,N_14184,N_14216);
xor U14700 (N_14700,N_14610,N_14618);
nand U14701 (N_14701,N_14683,N_14686);
and U14702 (N_14702,N_14501,N_14672);
and U14703 (N_14703,N_14636,N_14569);
nand U14704 (N_14704,N_14478,N_14655);
xnor U14705 (N_14705,N_14679,N_14598);
xor U14706 (N_14706,N_14422,N_14443);
xor U14707 (N_14707,N_14600,N_14646);
nand U14708 (N_14708,N_14473,N_14461);
and U14709 (N_14709,N_14680,N_14625);
nor U14710 (N_14710,N_14475,N_14429);
nand U14711 (N_14711,N_14690,N_14476);
nor U14712 (N_14712,N_14510,N_14420);
and U14713 (N_14713,N_14531,N_14511);
nor U14714 (N_14714,N_14417,N_14620);
and U14715 (N_14715,N_14615,N_14468);
or U14716 (N_14716,N_14412,N_14538);
nor U14717 (N_14717,N_14582,N_14436);
and U14718 (N_14718,N_14589,N_14604);
or U14719 (N_14719,N_14602,N_14612);
nor U14720 (N_14720,N_14479,N_14428);
or U14721 (N_14721,N_14611,N_14606);
and U14722 (N_14722,N_14536,N_14546);
xnor U14723 (N_14723,N_14623,N_14601);
nor U14724 (N_14724,N_14493,N_14544);
nand U14725 (N_14725,N_14669,N_14496);
nor U14726 (N_14726,N_14505,N_14557);
xor U14727 (N_14727,N_14627,N_14539);
nand U14728 (N_14728,N_14547,N_14400);
or U14729 (N_14729,N_14518,N_14577);
xnor U14730 (N_14730,N_14503,N_14421);
xor U14731 (N_14731,N_14540,N_14682);
nor U14732 (N_14732,N_14563,N_14595);
nand U14733 (N_14733,N_14652,N_14519);
xor U14734 (N_14734,N_14537,N_14662);
nand U14735 (N_14735,N_14413,N_14489);
or U14736 (N_14736,N_14437,N_14504);
and U14737 (N_14737,N_14454,N_14653);
nor U14738 (N_14738,N_14564,N_14403);
nand U14739 (N_14739,N_14658,N_14432);
xnor U14740 (N_14740,N_14415,N_14659);
xnor U14741 (N_14741,N_14630,N_14430);
xor U14742 (N_14742,N_14433,N_14483);
or U14743 (N_14743,N_14425,N_14462);
nand U14744 (N_14744,N_14522,N_14688);
or U14745 (N_14745,N_14472,N_14626);
xnor U14746 (N_14746,N_14605,N_14427);
nor U14747 (N_14747,N_14671,N_14527);
xnor U14748 (N_14748,N_14444,N_14456);
and U14749 (N_14749,N_14418,N_14593);
or U14750 (N_14750,N_14494,N_14555);
nor U14751 (N_14751,N_14699,N_14534);
and U14752 (N_14752,N_14556,N_14491);
and U14753 (N_14753,N_14463,N_14543);
and U14754 (N_14754,N_14645,N_14525);
or U14755 (N_14755,N_14666,N_14517);
xnor U14756 (N_14756,N_14471,N_14573);
and U14757 (N_14757,N_14624,N_14550);
or U14758 (N_14758,N_14465,N_14692);
xor U14759 (N_14759,N_14594,N_14558);
nor U14760 (N_14760,N_14668,N_14635);
or U14761 (N_14761,N_14445,N_14661);
xor U14762 (N_14762,N_14617,N_14657);
nand U14763 (N_14763,N_14591,N_14466);
and U14764 (N_14764,N_14584,N_14440);
and U14765 (N_14765,N_14632,N_14435);
and U14766 (N_14766,N_14634,N_14514);
nand U14767 (N_14767,N_14684,N_14404);
nor U14768 (N_14768,N_14580,N_14674);
or U14769 (N_14769,N_14667,N_14631);
nand U14770 (N_14770,N_14481,N_14545);
nor U14771 (N_14771,N_14449,N_14490);
xnor U14772 (N_14772,N_14560,N_14665);
nand U14773 (N_14773,N_14687,N_14597);
xnor U14774 (N_14774,N_14438,N_14551);
or U14775 (N_14775,N_14681,N_14638);
xor U14776 (N_14776,N_14434,N_14694);
or U14777 (N_14777,N_14486,N_14520);
nor U14778 (N_14778,N_14696,N_14664);
or U14779 (N_14779,N_14416,N_14528);
xnor U14780 (N_14780,N_14502,N_14693);
nor U14781 (N_14781,N_14571,N_14458);
xnor U14782 (N_14782,N_14500,N_14526);
nor U14783 (N_14783,N_14512,N_14648);
xnor U14784 (N_14784,N_14575,N_14603);
or U14785 (N_14785,N_14450,N_14419);
nand U14786 (N_14786,N_14565,N_14678);
nor U14787 (N_14787,N_14574,N_14570);
and U14788 (N_14788,N_14513,N_14523);
and U14789 (N_14789,N_14549,N_14487);
and U14790 (N_14790,N_14590,N_14559);
nand U14791 (N_14791,N_14643,N_14407);
nor U14792 (N_14792,N_14497,N_14414);
nand U14793 (N_14793,N_14408,N_14495);
xor U14794 (N_14794,N_14609,N_14698);
or U14795 (N_14795,N_14548,N_14424);
xnor U14796 (N_14796,N_14685,N_14405);
or U14797 (N_14797,N_14562,N_14467);
or U14798 (N_14798,N_14524,N_14689);
or U14799 (N_14799,N_14406,N_14647);
and U14800 (N_14800,N_14637,N_14533);
or U14801 (N_14801,N_14629,N_14515);
or U14802 (N_14802,N_14695,N_14516);
xor U14803 (N_14803,N_14578,N_14459);
and U14804 (N_14804,N_14535,N_14452);
xor U14805 (N_14805,N_14485,N_14423);
nor U14806 (N_14806,N_14585,N_14616);
xor U14807 (N_14807,N_14469,N_14411);
and U14808 (N_14808,N_14673,N_14691);
or U14809 (N_14809,N_14656,N_14470);
nand U14810 (N_14810,N_14460,N_14439);
and U14811 (N_14811,N_14457,N_14447);
and U14812 (N_14812,N_14441,N_14676);
nor U14813 (N_14813,N_14608,N_14426);
xnor U14814 (N_14814,N_14509,N_14508);
or U14815 (N_14815,N_14431,N_14554);
nand U14816 (N_14816,N_14566,N_14663);
or U14817 (N_14817,N_14529,N_14644);
and U14818 (N_14818,N_14583,N_14530);
or U14819 (N_14819,N_14542,N_14650);
xnor U14820 (N_14820,N_14649,N_14567);
nor U14821 (N_14821,N_14521,N_14639);
and U14822 (N_14822,N_14552,N_14464);
xnor U14823 (N_14823,N_14654,N_14622);
or U14824 (N_14824,N_14614,N_14677);
nand U14825 (N_14825,N_14477,N_14532);
nand U14826 (N_14826,N_14572,N_14619);
nand U14827 (N_14827,N_14628,N_14507);
nor U14828 (N_14828,N_14561,N_14488);
nor U14829 (N_14829,N_14596,N_14568);
nand U14830 (N_14830,N_14451,N_14660);
and U14831 (N_14831,N_14402,N_14675);
xor U14832 (N_14832,N_14670,N_14409);
or U14833 (N_14833,N_14499,N_14446);
or U14834 (N_14834,N_14506,N_14581);
and U14835 (N_14835,N_14474,N_14613);
nor U14836 (N_14836,N_14579,N_14587);
and U14837 (N_14837,N_14482,N_14633);
nand U14838 (N_14838,N_14553,N_14410);
or U14839 (N_14839,N_14642,N_14453);
or U14840 (N_14840,N_14651,N_14480);
nand U14841 (N_14841,N_14455,N_14498);
xnor U14842 (N_14842,N_14621,N_14640);
nand U14843 (N_14843,N_14401,N_14442);
nand U14844 (N_14844,N_14697,N_14576);
nor U14845 (N_14845,N_14588,N_14541);
nand U14846 (N_14846,N_14586,N_14448);
and U14847 (N_14847,N_14492,N_14599);
nor U14848 (N_14848,N_14607,N_14484);
nor U14849 (N_14849,N_14592,N_14641);
and U14850 (N_14850,N_14413,N_14515);
xnor U14851 (N_14851,N_14573,N_14596);
xnor U14852 (N_14852,N_14431,N_14600);
xor U14853 (N_14853,N_14422,N_14695);
nand U14854 (N_14854,N_14696,N_14628);
xnor U14855 (N_14855,N_14608,N_14458);
nand U14856 (N_14856,N_14439,N_14502);
nor U14857 (N_14857,N_14514,N_14460);
and U14858 (N_14858,N_14676,N_14654);
nor U14859 (N_14859,N_14499,N_14491);
xor U14860 (N_14860,N_14414,N_14522);
nor U14861 (N_14861,N_14557,N_14407);
nor U14862 (N_14862,N_14629,N_14567);
nand U14863 (N_14863,N_14517,N_14494);
and U14864 (N_14864,N_14532,N_14633);
nand U14865 (N_14865,N_14486,N_14405);
xor U14866 (N_14866,N_14477,N_14660);
and U14867 (N_14867,N_14505,N_14604);
nor U14868 (N_14868,N_14651,N_14573);
xor U14869 (N_14869,N_14471,N_14601);
or U14870 (N_14870,N_14609,N_14410);
xnor U14871 (N_14871,N_14402,N_14645);
xor U14872 (N_14872,N_14492,N_14413);
nand U14873 (N_14873,N_14517,N_14418);
nor U14874 (N_14874,N_14673,N_14616);
nor U14875 (N_14875,N_14572,N_14617);
and U14876 (N_14876,N_14596,N_14653);
nor U14877 (N_14877,N_14452,N_14429);
xnor U14878 (N_14878,N_14602,N_14501);
nor U14879 (N_14879,N_14400,N_14501);
or U14880 (N_14880,N_14607,N_14412);
and U14881 (N_14881,N_14540,N_14465);
nor U14882 (N_14882,N_14670,N_14659);
and U14883 (N_14883,N_14478,N_14405);
or U14884 (N_14884,N_14683,N_14607);
or U14885 (N_14885,N_14678,N_14674);
and U14886 (N_14886,N_14655,N_14673);
or U14887 (N_14887,N_14475,N_14480);
or U14888 (N_14888,N_14424,N_14417);
nand U14889 (N_14889,N_14575,N_14663);
nor U14890 (N_14890,N_14494,N_14445);
nor U14891 (N_14891,N_14463,N_14420);
and U14892 (N_14892,N_14620,N_14458);
nor U14893 (N_14893,N_14643,N_14647);
nand U14894 (N_14894,N_14463,N_14565);
or U14895 (N_14895,N_14557,N_14561);
and U14896 (N_14896,N_14471,N_14507);
and U14897 (N_14897,N_14584,N_14646);
xnor U14898 (N_14898,N_14402,N_14692);
nor U14899 (N_14899,N_14478,N_14639);
nor U14900 (N_14900,N_14481,N_14432);
nor U14901 (N_14901,N_14692,N_14472);
nand U14902 (N_14902,N_14641,N_14440);
nor U14903 (N_14903,N_14559,N_14471);
nand U14904 (N_14904,N_14468,N_14467);
xor U14905 (N_14905,N_14431,N_14592);
or U14906 (N_14906,N_14659,N_14677);
nand U14907 (N_14907,N_14434,N_14492);
and U14908 (N_14908,N_14547,N_14684);
and U14909 (N_14909,N_14507,N_14554);
nand U14910 (N_14910,N_14658,N_14416);
xnor U14911 (N_14911,N_14454,N_14603);
nand U14912 (N_14912,N_14612,N_14630);
nand U14913 (N_14913,N_14583,N_14444);
or U14914 (N_14914,N_14407,N_14577);
nand U14915 (N_14915,N_14538,N_14501);
nor U14916 (N_14916,N_14685,N_14652);
xnor U14917 (N_14917,N_14605,N_14411);
nand U14918 (N_14918,N_14653,N_14572);
or U14919 (N_14919,N_14429,N_14642);
and U14920 (N_14920,N_14654,N_14460);
nand U14921 (N_14921,N_14586,N_14641);
xnor U14922 (N_14922,N_14635,N_14553);
and U14923 (N_14923,N_14621,N_14413);
nand U14924 (N_14924,N_14658,N_14669);
nor U14925 (N_14925,N_14425,N_14558);
or U14926 (N_14926,N_14535,N_14410);
and U14927 (N_14927,N_14469,N_14685);
nand U14928 (N_14928,N_14615,N_14568);
xor U14929 (N_14929,N_14653,N_14466);
and U14930 (N_14930,N_14435,N_14471);
nor U14931 (N_14931,N_14439,N_14485);
and U14932 (N_14932,N_14515,N_14620);
nand U14933 (N_14933,N_14457,N_14480);
xor U14934 (N_14934,N_14438,N_14558);
nand U14935 (N_14935,N_14465,N_14523);
and U14936 (N_14936,N_14533,N_14408);
or U14937 (N_14937,N_14468,N_14609);
nand U14938 (N_14938,N_14667,N_14473);
and U14939 (N_14939,N_14449,N_14505);
nor U14940 (N_14940,N_14430,N_14498);
nor U14941 (N_14941,N_14665,N_14559);
nor U14942 (N_14942,N_14461,N_14614);
and U14943 (N_14943,N_14497,N_14681);
nor U14944 (N_14944,N_14654,N_14416);
or U14945 (N_14945,N_14641,N_14517);
xnor U14946 (N_14946,N_14418,N_14566);
nor U14947 (N_14947,N_14403,N_14510);
xor U14948 (N_14948,N_14587,N_14680);
xor U14949 (N_14949,N_14438,N_14444);
xnor U14950 (N_14950,N_14490,N_14570);
nor U14951 (N_14951,N_14632,N_14427);
nand U14952 (N_14952,N_14632,N_14627);
nand U14953 (N_14953,N_14548,N_14501);
nor U14954 (N_14954,N_14450,N_14550);
or U14955 (N_14955,N_14580,N_14658);
nor U14956 (N_14956,N_14696,N_14671);
and U14957 (N_14957,N_14524,N_14405);
nand U14958 (N_14958,N_14547,N_14585);
xnor U14959 (N_14959,N_14443,N_14466);
xor U14960 (N_14960,N_14463,N_14631);
xor U14961 (N_14961,N_14448,N_14639);
xnor U14962 (N_14962,N_14670,N_14556);
or U14963 (N_14963,N_14459,N_14619);
nor U14964 (N_14964,N_14444,N_14465);
xor U14965 (N_14965,N_14400,N_14410);
or U14966 (N_14966,N_14505,N_14591);
xnor U14967 (N_14967,N_14654,N_14638);
and U14968 (N_14968,N_14459,N_14552);
nand U14969 (N_14969,N_14502,N_14584);
and U14970 (N_14970,N_14521,N_14413);
xor U14971 (N_14971,N_14629,N_14447);
nand U14972 (N_14972,N_14663,N_14657);
and U14973 (N_14973,N_14604,N_14672);
nor U14974 (N_14974,N_14619,N_14608);
nand U14975 (N_14975,N_14570,N_14435);
xor U14976 (N_14976,N_14495,N_14528);
or U14977 (N_14977,N_14682,N_14570);
nor U14978 (N_14978,N_14484,N_14461);
nor U14979 (N_14979,N_14469,N_14499);
xor U14980 (N_14980,N_14514,N_14561);
xor U14981 (N_14981,N_14486,N_14478);
nand U14982 (N_14982,N_14683,N_14560);
xnor U14983 (N_14983,N_14652,N_14464);
nor U14984 (N_14984,N_14676,N_14529);
nand U14985 (N_14985,N_14543,N_14609);
nor U14986 (N_14986,N_14579,N_14575);
nand U14987 (N_14987,N_14616,N_14686);
and U14988 (N_14988,N_14608,N_14554);
or U14989 (N_14989,N_14546,N_14412);
and U14990 (N_14990,N_14587,N_14410);
nand U14991 (N_14991,N_14596,N_14577);
xor U14992 (N_14992,N_14587,N_14626);
and U14993 (N_14993,N_14429,N_14483);
or U14994 (N_14994,N_14446,N_14478);
and U14995 (N_14995,N_14669,N_14450);
or U14996 (N_14996,N_14481,N_14680);
nor U14997 (N_14997,N_14491,N_14446);
or U14998 (N_14998,N_14445,N_14416);
nand U14999 (N_14999,N_14472,N_14529);
nand UO_0 (O_0,N_14774,N_14848);
or UO_1 (O_1,N_14792,N_14985);
xnor UO_2 (O_2,N_14920,N_14751);
xnor UO_3 (O_3,N_14932,N_14767);
nor UO_4 (O_4,N_14967,N_14715);
and UO_5 (O_5,N_14914,N_14736);
xor UO_6 (O_6,N_14880,N_14706);
nand UO_7 (O_7,N_14860,N_14712);
nor UO_8 (O_8,N_14870,N_14950);
or UO_9 (O_9,N_14927,N_14891);
and UO_10 (O_10,N_14817,N_14776);
and UO_11 (O_11,N_14924,N_14784);
xnor UO_12 (O_12,N_14794,N_14994);
nand UO_13 (O_13,N_14990,N_14707);
nor UO_14 (O_14,N_14865,N_14704);
or UO_15 (O_15,N_14943,N_14863);
nand UO_16 (O_16,N_14771,N_14778);
or UO_17 (O_17,N_14905,N_14839);
nand UO_18 (O_18,N_14913,N_14906);
nor UO_19 (O_19,N_14945,N_14747);
and UO_20 (O_20,N_14833,N_14808);
nand UO_21 (O_21,N_14965,N_14903);
xor UO_22 (O_22,N_14749,N_14717);
nand UO_23 (O_23,N_14741,N_14814);
nor UO_24 (O_24,N_14804,N_14899);
or UO_25 (O_25,N_14879,N_14700);
xor UO_26 (O_26,N_14872,N_14782);
or UO_27 (O_27,N_14957,N_14962);
nand UO_28 (O_28,N_14830,N_14881);
or UO_29 (O_29,N_14760,N_14827);
nor UO_30 (O_30,N_14998,N_14757);
nor UO_31 (O_31,N_14840,N_14931);
or UO_32 (O_32,N_14705,N_14721);
nand UO_33 (O_33,N_14734,N_14766);
or UO_34 (O_34,N_14867,N_14810);
xnor UO_35 (O_35,N_14798,N_14912);
xor UO_36 (O_36,N_14878,N_14823);
nor UO_37 (O_37,N_14789,N_14761);
xnor UO_38 (O_38,N_14788,N_14919);
xnor UO_39 (O_39,N_14714,N_14873);
xor UO_40 (O_40,N_14701,N_14902);
nand UO_41 (O_41,N_14801,N_14960);
nand UO_42 (O_42,N_14862,N_14755);
xnor UO_43 (O_43,N_14956,N_14738);
xor UO_44 (O_44,N_14874,N_14775);
xor UO_45 (O_45,N_14948,N_14875);
nor UO_46 (O_46,N_14832,N_14959);
nor UO_47 (O_47,N_14971,N_14897);
and UO_48 (O_48,N_14951,N_14984);
and UO_49 (O_49,N_14882,N_14837);
and UO_50 (O_50,N_14941,N_14785);
nand UO_51 (O_51,N_14972,N_14996);
xor UO_52 (O_52,N_14961,N_14890);
or UO_53 (O_53,N_14917,N_14816);
and UO_54 (O_54,N_14711,N_14783);
or UO_55 (O_55,N_14773,N_14974);
or UO_56 (O_56,N_14796,N_14886);
nand UO_57 (O_57,N_14724,N_14849);
nor UO_58 (O_58,N_14979,N_14940);
or UO_59 (O_59,N_14938,N_14790);
nand UO_60 (O_60,N_14800,N_14892);
nor UO_61 (O_61,N_14807,N_14722);
and UO_62 (O_62,N_14929,N_14716);
or UO_63 (O_63,N_14793,N_14861);
and UO_64 (O_64,N_14825,N_14740);
nand UO_65 (O_65,N_14947,N_14909);
or UO_66 (O_66,N_14908,N_14786);
nand UO_67 (O_67,N_14847,N_14992);
or UO_68 (O_68,N_14826,N_14703);
nor UO_69 (O_69,N_14958,N_14828);
or UO_70 (O_70,N_14859,N_14780);
nand UO_71 (O_71,N_14728,N_14991);
xnor UO_72 (O_72,N_14896,N_14748);
xor UO_73 (O_73,N_14987,N_14883);
nand UO_74 (O_74,N_14744,N_14819);
xor UO_75 (O_75,N_14916,N_14730);
nor UO_76 (O_76,N_14752,N_14895);
and UO_77 (O_77,N_14885,N_14973);
nand UO_78 (O_78,N_14753,N_14777);
xnor UO_79 (O_79,N_14710,N_14713);
and UO_80 (O_80,N_14723,N_14888);
nand UO_81 (O_81,N_14799,N_14708);
and UO_82 (O_82,N_14797,N_14756);
or UO_83 (O_83,N_14871,N_14930);
or UO_84 (O_84,N_14904,N_14846);
xor UO_85 (O_85,N_14968,N_14750);
or UO_86 (O_86,N_14763,N_14813);
nand UO_87 (O_87,N_14925,N_14806);
nor UO_88 (O_88,N_14944,N_14745);
or UO_89 (O_89,N_14762,N_14719);
nor UO_90 (O_90,N_14975,N_14964);
nor UO_91 (O_91,N_14988,N_14970);
nor UO_92 (O_92,N_14765,N_14969);
and UO_93 (O_93,N_14999,N_14854);
and UO_94 (O_94,N_14995,N_14787);
xnor UO_95 (O_95,N_14889,N_14836);
or UO_96 (O_96,N_14853,N_14937);
nand UO_97 (O_97,N_14893,N_14923);
or UO_98 (O_98,N_14898,N_14894);
and UO_99 (O_99,N_14918,N_14737);
or UO_100 (O_100,N_14877,N_14815);
nand UO_101 (O_101,N_14842,N_14791);
nor UO_102 (O_102,N_14869,N_14981);
nand UO_103 (O_103,N_14868,N_14746);
nand UO_104 (O_104,N_14844,N_14866);
or UO_105 (O_105,N_14742,N_14758);
and UO_106 (O_106,N_14936,N_14976);
nand UO_107 (O_107,N_14732,N_14911);
and UO_108 (O_108,N_14768,N_14946);
xnor UO_109 (O_109,N_14820,N_14921);
nand UO_110 (O_110,N_14809,N_14831);
and UO_111 (O_111,N_14986,N_14997);
and UO_112 (O_112,N_14852,N_14834);
nand UO_113 (O_113,N_14841,N_14907);
nor UO_114 (O_114,N_14926,N_14993);
and UO_115 (O_115,N_14939,N_14978);
and UO_116 (O_116,N_14935,N_14983);
nand UO_117 (O_117,N_14915,N_14726);
xor UO_118 (O_118,N_14838,N_14764);
or UO_119 (O_119,N_14900,N_14858);
nor UO_120 (O_120,N_14769,N_14727);
xnor UO_121 (O_121,N_14843,N_14795);
and UO_122 (O_122,N_14901,N_14928);
nand UO_123 (O_123,N_14733,N_14933);
nand UO_124 (O_124,N_14942,N_14910);
or UO_125 (O_125,N_14864,N_14821);
nor UO_126 (O_126,N_14702,N_14954);
xor UO_127 (O_127,N_14812,N_14803);
nand UO_128 (O_128,N_14731,N_14811);
and UO_129 (O_129,N_14735,N_14934);
xnor UO_130 (O_130,N_14743,N_14822);
or UO_131 (O_131,N_14802,N_14779);
xor UO_132 (O_132,N_14739,N_14805);
nand UO_133 (O_133,N_14949,N_14718);
and UO_134 (O_134,N_14982,N_14887);
nor UO_135 (O_135,N_14829,N_14709);
or UO_136 (O_136,N_14922,N_14980);
or UO_137 (O_137,N_14977,N_14850);
nor UO_138 (O_138,N_14851,N_14729);
or UO_139 (O_139,N_14720,N_14818);
nor UO_140 (O_140,N_14989,N_14955);
nand UO_141 (O_141,N_14855,N_14963);
nand UO_142 (O_142,N_14770,N_14876);
nand UO_143 (O_143,N_14952,N_14953);
nor UO_144 (O_144,N_14856,N_14725);
nor UO_145 (O_145,N_14857,N_14759);
and UO_146 (O_146,N_14966,N_14781);
nand UO_147 (O_147,N_14884,N_14772);
and UO_148 (O_148,N_14824,N_14754);
xor UO_149 (O_149,N_14835,N_14845);
or UO_150 (O_150,N_14849,N_14998);
or UO_151 (O_151,N_14793,N_14842);
nor UO_152 (O_152,N_14907,N_14764);
or UO_153 (O_153,N_14849,N_14743);
nand UO_154 (O_154,N_14979,N_14737);
or UO_155 (O_155,N_14706,N_14972);
xnor UO_156 (O_156,N_14815,N_14862);
and UO_157 (O_157,N_14869,N_14786);
or UO_158 (O_158,N_14789,N_14911);
nand UO_159 (O_159,N_14825,N_14810);
or UO_160 (O_160,N_14808,N_14847);
and UO_161 (O_161,N_14806,N_14765);
nand UO_162 (O_162,N_14882,N_14774);
nand UO_163 (O_163,N_14999,N_14963);
xor UO_164 (O_164,N_14783,N_14747);
and UO_165 (O_165,N_14712,N_14932);
nand UO_166 (O_166,N_14951,N_14787);
and UO_167 (O_167,N_14957,N_14976);
and UO_168 (O_168,N_14701,N_14924);
or UO_169 (O_169,N_14734,N_14754);
and UO_170 (O_170,N_14811,N_14853);
or UO_171 (O_171,N_14851,N_14963);
or UO_172 (O_172,N_14770,N_14724);
nand UO_173 (O_173,N_14950,N_14789);
xnor UO_174 (O_174,N_14786,N_14984);
xnor UO_175 (O_175,N_14990,N_14718);
nor UO_176 (O_176,N_14767,N_14729);
and UO_177 (O_177,N_14982,N_14781);
or UO_178 (O_178,N_14799,N_14755);
nor UO_179 (O_179,N_14840,N_14901);
nor UO_180 (O_180,N_14901,N_14738);
nand UO_181 (O_181,N_14792,N_14966);
or UO_182 (O_182,N_14900,N_14860);
and UO_183 (O_183,N_14991,N_14809);
or UO_184 (O_184,N_14716,N_14844);
nor UO_185 (O_185,N_14966,N_14962);
or UO_186 (O_186,N_14969,N_14866);
or UO_187 (O_187,N_14934,N_14812);
nor UO_188 (O_188,N_14890,N_14854);
and UO_189 (O_189,N_14861,N_14794);
xnor UO_190 (O_190,N_14830,N_14891);
and UO_191 (O_191,N_14800,N_14900);
or UO_192 (O_192,N_14704,N_14898);
nor UO_193 (O_193,N_14831,N_14814);
or UO_194 (O_194,N_14785,N_14780);
nand UO_195 (O_195,N_14746,N_14964);
xor UO_196 (O_196,N_14821,N_14714);
and UO_197 (O_197,N_14838,N_14872);
xnor UO_198 (O_198,N_14985,N_14885);
xor UO_199 (O_199,N_14963,N_14842);
and UO_200 (O_200,N_14812,N_14787);
or UO_201 (O_201,N_14752,N_14742);
nor UO_202 (O_202,N_14758,N_14821);
or UO_203 (O_203,N_14810,N_14979);
xor UO_204 (O_204,N_14745,N_14729);
nand UO_205 (O_205,N_14711,N_14709);
nor UO_206 (O_206,N_14953,N_14860);
nand UO_207 (O_207,N_14725,N_14980);
nor UO_208 (O_208,N_14980,N_14840);
xor UO_209 (O_209,N_14707,N_14780);
and UO_210 (O_210,N_14901,N_14804);
nor UO_211 (O_211,N_14753,N_14995);
xor UO_212 (O_212,N_14989,N_14775);
or UO_213 (O_213,N_14743,N_14786);
and UO_214 (O_214,N_14948,N_14730);
and UO_215 (O_215,N_14910,N_14929);
and UO_216 (O_216,N_14804,N_14770);
nor UO_217 (O_217,N_14807,N_14700);
xnor UO_218 (O_218,N_14887,N_14903);
nand UO_219 (O_219,N_14927,N_14907);
nor UO_220 (O_220,N_14949,N_14880);
nor UO_221 (O_221,N_14705,N_14944);
or UO_222 (O_222,N_14910,N_14908);
or UO_223 (O_223,N_14740,N_14848);
nor UO_224 (O_224,N_14777,N_14888);
nand UO_225 (O_225,N_14987,N_14841);
nor UO_226 (O_226,N_14769,N_14900);
or UO_227 (O_227,N_14948,N_14782);
xnor UO_228 (O_228,N_14842,N_14941);
xnor UO_229 (O_229,N_14857,N_14725);
and UO_230 (O_230,N_14922,N_14854);
nand UO_231 (O_231,N_14758,N_14991);
or UO_232 (O_232,N_14941,N_14830);
nand UO_233 (O_233,N_14810,N_14864);
xor UO_234 (O_234,N_14728,N_14712);
and UO_235 (O_235,N_14855,N_14947);
or UO_236 (O_236,N_14702,N_14820);
and UO_237 (O_237,N_14754,N_14758);
nand UO_238 (O_238,N_14823,N_14963);
nor UO_239 (O_239,N_14796,N_14763);
nand UO_240 (O_240,N_14838,N_14824);
nor UO_241 (O_241,N_14852,N_14996);
or UO_242 (O_242,N_14856,N_14924);
and UO_243 (O_243,N_14754,N_14762);
nor UO_244 (O_244,N_14943,N_14893);
and UO_245 (O_245,N_14820,N_14824);
and UO_246 (O_246,N_14822,N_14786);
and UO_247 (O_247,N_14836,N_14848);
nor UO_248 (O_248,N_14740,N_14813);
nand UO_249 (O_249,N_14769,N_14967);
and UO_250 (O_250,N_14749,N_14994);
or UO_251 (O_251,N_14857,N_14858);
and UO_252 (O_252,N_14914,N_14825);
xor UO_253 (O_253,N_14760,N_14817);
xnor UO_254 (O_254,N_14814,N_14821);
nand UO_255 (O_255,N_14819,N_14992);
or UO_256 (O_256,N_14868,N_14917);
nand UO_257 (O_257,N_14826,N_14917);
and UO_258 (O_258,N_14934,N_14874);
xor UO_259 (O_259,N_14968,N_14745);
nor UO_260 (O_260,N_14767,N_14832);
nand UO_261 (O_261,N_14791,N_14837);
nand UO_262 (O_262,N_14907,N_14954);
and UO_263 (O_263,N_14967,N_14833);
and UO_264 (O_264,N_14802,N_14903);
nand UO_265 (O_265,N_14729,N_14712);
and UO_266 (O_266,N_14853,N_14841);
xor UO_267 (O_267,N_14929,N_14706);
or UO_268 (O_268,N_14863,N_14726);
and UO_269 (O_269,N_14742,N_14886);
and UO_270 (O_270,N_14869,N_14807);
and UO_271 (O_271,N_14828,N_14800);
nand UO_272 (O_272,N_14978,N_14892);
nand UO_273 (O_273,N_14844,N_14746);
nor UO_274 (O_274,N_14834,N_14859);
or UO_275 (O_275,N_14722,N_14801);
nor UO_276 (O_276,N_14765,N_14758);
nand UO_277 (O_277,N_14937,N_14923);
nor UO_278 (O_278,N_14996,N_14989);
and UO_279 (O_279,N_14971,N_14810);
and UO_280 (O_280,N_14744,N_14937);
and UO_281 (O_281,N_14821,N_14939);
xnor UO_282 (O_282,N_14857,N_14746);
and UO_283 (O_283,N_14976,N_14801);
xor UO_284 (O_284,N_14802,N_14868);
nor UO_285 (O_285,N_14953,N_14778);
nor UO_286 (O_286,N_14987,N_14702);
nor UO_287 (O_287,N_14715,N_14829);
nand UO_288 (O_288,N_14785,N_14898);
xor UO_289 (O_289,N_14878,N_14990);
nand UO_290 (O_290,N_14773,N_14774);
nand UO_291 (O_291,N_14970,N_14815);
xor UO_292 (O_292,N_14718,N_14706);
and UO_293 (O_293,N_14994,N_14978);
or UO_294 (O_294,N_14988,N_14978);
or UO_295 (O_295,N_14739,N_14924);
nor UO_296 (O_296,N_14814,N_14904);
xor UO_297 (O_297,N_14907,N_14702);
xnor UO_298 (O_298,N_14888,N_14905);
xor UO_299 (O_299,N_14842,N_14763);
and UO_300 (O_300,N_14837,N_14741);
or UO_301 (O_301,N_14852,N_14752);
xnor UO_302 (O_302,N_14878,N_14986);
nor UO_303 (O_303,N_14732,N_14716);
nor UO_304 (O_304,N_14964,N_14740);
and UO_305 (O_305,N_14857,N_14828);
nand UO_306 (O_306,N_14968,N_14865);
nor UO_307 (O_307,N_14884,N_14894);
nand UO_308 (O_308,N_14931,N_14753);
nor UO_309 (O_309,N_14910,N_14835);
and UO_310 (O_310,N_14800,N_14923);
or UO_311 (O_311,N_14792,N_14988);
nor UO_312 (O_312,N_14901,N_14757);
or UO_313 (O_313,N_14714,N_14984);
nand UO_314 (O_314,N_14883,N_14973);
nor UO_315 (O_315,N_14823,N_14999);
nor UO_316 (O_316,N_14804,N_14908);
xnor UO_317 (O_317,N_14835,N_14816);
xor UO_318 (O_318,N_14979,N_14782);
and UO_319 (O_319,N_14865,N_14889);
nor UO_320 (O_320,N_14820,N_14789);
and UO_321 (O_321,N_14828,N_14893);
xnor UO_322 (O_322,N_14945,N_14983);
xor UO_323 (O_323,N_14770,N_14982);
nor UO_324 (O_324,N_14713,N_14911);
and UO_325 (O_325,N_14784,N_14798);
nor UO_326 (O_326,N_14990,N_14888);
and UO_327 (O_327,N_14969,N_14847);
and UO_328 (O_328,N_14914,N_14995);
or UO_329 (O_329,N_14712,N_14703);
nor UO_330 (O_330,N_14969,N_14733);
nand UO_331 (O_331,N_14957,N_14975);
nand UO_332 (O_332,N_14788,N_14994);
or UO_333 (O_333,N_14952,N_14791);
nor UO_334 (O_334,N_14837,N_14877);
nand UO_335 (O_335,N_14762,N_14813);
xnor UO_336 (O_336,N_14942,N_14882);
nor UO_337 (O_337,N_14758,N_14920);
xor UO_338 (O_338,N_14889,N_14734);
or UO_339 (O_339,N_14753,N_14809);
nor UO_340 (O_340,N_14869,N_14906);
nand UO_341 (O_341,N_14761,N_14702);
nand UO_342 (O_342,N_14702,N_14718);
nor UO_343 (O_343,N_14777,N_14801);
nor UO_344 (O_344,N_14723,N_14816);
and UO_345 (O_345,N_14837,N_14865);
xnor UO_346 (O_346,N_14823,N_14968);
nand UO_347 (O_347,N_14832,N_14792);
or UO_348 (O_348,N_14820,N_14909);
xor UO_349 (O_349,N_14882,N_14711);
or UO_350 (O_350,N_14890,N_14914);
nor UO_351 (O_351,N_14974,N_14795);
nor UO_352 (O_352,N_14776,N_14825);
or UO_353 (O_353,N_14840,N_14705);
nand UO_354 (O_354,N_14899,N_14927);
or UO_355 (O_355,N_14840,N_14919);
and UO_356 (O_356,N_14739,N_14758);
or UO_357 (O_357,N_14927,N_14982);
or UO_358 (O_358,N_14826,N_14989);
nor UO_359 (O_359,N_14822,N_14947);
nand UO_360 (O_360,N_14815,N_14768);
xnor UO_361 (O_361,N_14948,N_14937);
or UO_362 (O_362,N_14904,N_14981);
or UO_363 (O_363,N_14773,N_14856);
nand UO_364 (O_364,N_14997,N_14727);
xnor UO_365 (O_365,N_14701,N_14758);
and UO_366 (O_366,N_14992,N_14914);
and UO_367 (O_367,N_14784,N_14882);
nor UO_368 (O_368,N_14720,N_14896);
xor UO_369 (O_369,N_14943,N_14743);
nor UO_370 (O_370,N_14865,N_14871);
nor UO_371 (O_371,N_14809,N_14776);
or UO_372 (O_372,N_14703,N_14746);
xnor UO_373 (O_373,N_14887,N_14951);
nor UO_374 (O_374,N_14940,N_14853);
or UO_375 (O_375,N_14855,N_14815);
or UO_376 (O_376,N_14730,N_14990);
or UO_377 (O_377,N_14764,N_14705);
nand UO_378 (O_378,N_14740,N_14910);
and UO_379 (O_379,N_14829,N_14786);
or UO_380 (O_380,N_14962,N_14710);
nor UO_381 (O_381,N_14998,N_14786);
or UO_382 (O_382,N_14886,N_14985);
nand UO_383 (O_383,N_14966,N_14959);
xor UO_384 (O_384,N_14901,N_14705);
nor UO_385 (O_385,N_14742,N_14957);
and UO_386 (O_386,N_14963,N_14804);
and UO_387 (O_387,N_14770,N_14767);
or UO_388 (O_388,N_14948,N_14897);
and UO_389 (O_389,N_14751,N_14703);
and UO_390 (O_390,N_14895,N_14965);
xor UO_391 (O_391,N_14996,N_14701);
or UO_392 (O_392,N_14897,N_14918);
xor UO_393 (O_393,N_14852,N_14872);
and UO_394 (O_394,N_14831,N_14829);
and UO_395 (O_395,N_14939,N_14715);
and UO_396 (O_396,N_14929,N_14907);
nor UO_397 (O_397,N_14731,N_14971);
nand UO_398 (O_398,N_14731,N_14726);
nand UO_399 (O_399,N_14909,N_14781);
xor UO_400 (O_400,N_14758,N_14787);
nor UO_401 (O_401,N_14739,N_14829);
and UO_402 (O_402,N_14946,N_14915);
and UO_403 (O_403,N_14763,N_14848);
xnor UO_404 (O_404,N_14833,N_14711);
or UO_405 (O_405,N_14734,N_14714);
or UO_406 (O_406,N_14729,N_14752);
and UO_407 (O_407,N_14876,N_14807);
xor UO_408 (O_408,N_14802,N_14861);
and UO_409 (O_409,N_14774,N_14802);
xor UO_410 (O_410,N_14941,N_14961);
or UO_411 (O_411,N_14994,N_14735);
nor UO_412 (O_412,N_14714,N_14930);
and UO_413 (O_413,N_14723,N_14756);
nand UO_414 (O_414,N_14895,N_14732);
nand UO_415 (O_415,N_14921,N_14893);
nand UO_416 (O_416,N_14919,N_14927);
and UO_417 (O_417,N_14924,N_14779);
xnor UO_418 (O_418,N_14771,N_14840);
or UO_419 (O_419,N_14949,N_14953);
and UO_420 (O_420,N_14753,N_14773);
nor UO_421 (O_421,N_14739,N_14717);
and UO_422 (O_422,N_14712,N_14789);
nand UO_423 (O_423,N_14855,N_14996);
or UO_424 (O_424,N_14852,N_14864);
and UO_425 (O_425,N_14914,N_14834);
nor UO_426 (O_426,N_14781,N_14712);
nor UO_427 (O_427,N_14958,N_14976);
and UO_428 (O_428,N_14756,N_14795);
nand UO_429 (O_429,N_14739,N_14830);
or UO_430 (O_430,N_14784,N_14929);
nor UO_431 (O_431,N_14912,N_14831);
nand UO_432 (O_432,N_14973,N_14862);
nand UO_433 (O_433,N_14904,N_14735);
and UO_434 (O_434,N_14985,N_14884);
nand UO_435 (O_435,N_14803,N_14727);
nor UO_436 (O_436,N_14972,N_14875);
xnor UO_437 (O_437,N_14967,N_14905);
nor UO_438 (O_438,N_14823,N_14969);
or UO_439 (O_439,N_14776,N_14855);
or UO_440 (O_440,N_14735,N_14786);
or UO_441 (O_441,N_14748,N_14795);
and UO_442 (O_442,N_14863,N_14896);
and UO_443 (O_443,N_14804,N_14962);
or UO_444 (O_444,N_14861,N_14822);
xnor UO_445 (O_445,N_14850,N_14762);
nand UO_446 (O_446,N_14778,N_14913);
xnor UO_447 (O_447,N_14857,N_14913);
or UO_448 (O_448,N_14977,N_14744);
or UO_449 (O_449,N_14785,N_14711);
nor UO_450 (O_450,N_14948,N_14813);
or UO_451 (O_451,N_14942,N_14965);
nor UO_452 (O_452,N_14782,N_14779);
nor UO_453 (O_453,N_14883,N_14956);
xnor UO_454 (O_454,N_14806,N_14911);
nand UO_455 (O_455,N_14710,N_14826);
xor UO_456 (O_456,N_14721,N_14825);
xnor UO_457 (O_457,N_14932,N_14833);
nor UO_458 (O_458,N_14929,N_14951);
xor UO_459 (O_459,N_14766,N_14717);
and UO_460 (O_460,N_14858,N_14913);
or UO_461 (O_461,N_14825,N_14965);
and UO_462 (O_462,N_14933,N_14791);
xnor UO_463 (O_463,N_14847,N_14931);
and UO_464 (O_464,N_14747,N_14856);
nand UO_465 (O_465,N_14896,N_14962);
and UO_466 (O_466,N_14852,N_14892);
xor UO_467 (O_467,N_14835,N_14887);
nor UO_468 (O_468,N_14736,N_14989);
nor UO_469 (O_469,N_14710,N_14905);
or UO_470 (O_470,N_14809,N_14865);
xor UO_471 (O_471,N_14827,N_14706);
and UO_472 (O_472,N_14945,N_14808);
and UO_473 (O_473,N_14798,N_14740);
nand UO_474 (O_474,N_14752,N_14981);
nand UO_475 (O_475,N_14900,N_14774);
xnor UO_476 (O_476,N_14702,N_14918);
nand UO_477 (O_477,N_14910,N_14739);
xnor UO_478 (O_478,N_14981,N_14787);
nand UO_479 (O_479,N_14940,N_14894);
or UO_480 (O_480,N_14774,N_14885);
nor UO_481 (O_481,N_14820,N_14900);
and UO_482 (O_482,N_14953,N_14881);
nor UO_483 (O_483,N_14997,N_14714);
nor UO_484 (O_484,N_14938,N_14835);
xnor UO_485 (O_485,N_14701,N_14732);
nand UO_486 (O_486,N_14930,N_14865);
nor UO_487 (O_487,N_14972,N_14990);
or UO_488 (O_488,N_14827,N_14857);
or UO_489 (O_489,N_14928,N_14841);
nor UO_490 (O_490,N_14760,N_14729);
nand UO_491 (O_491,N_14886,N_14939);
xnor UO_492 (O_492,N_14863,N_14975);
or UO_493 (O_493,N_14886,N_14708);
and UO_494 (O_494,N_14899,N_14847);
and UO_495 (O_495,N_14891,N_14880);
nor UO_496 (O_496,N_14799,N_14786);
and UO_497 (O_497,N_14959,N_14887);
xnor UO_498 (O_498,N_14828,N_14954);
nand UO_499 (O_499,N_14787,N_14999);
xor UO_500 (O_500,N_14745,N_14933);
nor UO_501 (O_501,N_14923,N_14851);
nor UO_502 (O_502,N_14832,N_14873);
nor UO_503 (O_503,N_14702,N_14721);
or UO_504 (O_504,N_14943,N_14995);
nor UO_505 (O_505,N_14788,N_14997);
xnor UO_506 (O_506,N_14904,N_14710);
or UO_507 (O_507,N_14777,N_14736);
and UO_508 (O_508,N_14750,N_14874);
or UO_509 (O_509,N_14903,N_14715);
nand UO_510 (O_510,N_14970,N_14911);
or UO_511 (O_511,N_14823,N_14926);
nand UO_512 (O_512,N_14774,N_14836);
nor UO_513 (O_513,N_14784,N_14829);
nor UO_514 (O_514,N_14868,N_14929);
and UO_515 (O_515,N_14940,N_14824);
or UO_516 (O_516,N_14784,N_14981);
and UO_517 (O_517,N_14859,N_14964);
xnor UO_518 (O_518,N_14773,N_14714);
nand UO_519 (O_519,N_14977,N_14710);
xor UO_520 (O_520,N_14907,N_14866);
xor UO_521 (O_521,N_14803,N_14723);
xor UO_522 (O_522,N_14838,N_14914);
or UO_523 (O_523,N_14986,N_14838);
or UO_524 (O_524,N_14725,N_14791);
xnor UO_525 (O_525,N_14940,N_14774);
nand UO_526 (O_526,N_14723,N_14812);
nand UO_527 (O_527,N_14796,N_14814);
nor UO_528 (O_528,N_14870,N_14905);
xor UO_529 (O_529,N_14701,N_14936);
nor UO_530 (O_530,N_14809,N_14866);
and UO_531 (O_531,N_14826,N_14931);
nand UO_532 (O_532,N_14917,N_14844);
and UO_533 (O_533,N_14878,N_14817);
nand UO_534 (O_534,N_14814,N_14862);
or UO_535 (O_535,N_14793,N_14870);
and UO_536 (O_536,N_14801,N_14911);
and UO_537 (O_537,N_14959,N_14750);
and UO_538 (O_538,N_14880,N_14794);
xor UO_539 (O_539,N_14923,N_14717);
nor UO_540 (O_540,N_14948,N_14715);
nand UO_541 (O_541,N_14729,N_14791);
or UO_542 (O_542,N_14961,N_14888);
nor UO_543 (O_543,N_14854,N_14865);
or UO_544 (O_544,N_14942,N_14837);
and UO_545 (O_545,N_14948,N_14803);
nor UO_546 (O_546,N_14984,N_14707);
or UO_547 (O_547,N_14713,N_14801);
xor UO_548 (O_548,N_14855,N_14832);
and UO_549 (O_549,N_14863,N_14748);
and UO_550 (O_550,N_14827,N_14822);
nor UO_551 (O_551,N_14730,N_14904);
nand UO_552 (O_552,N_14828,N_14842);
xor UO_553 (O_553,N_14787,N_14851);
nand UO_554 (O_554,N_14985,N_14782);
xnor UO_555 (O_555,N_14875,N_14985);
nor UO_556 (O_556,N_14733,N_14943);
and UO_557 (O_557,N_14892,N_14807);
nand UO_558 (O_558,N_14808,N_14800);
or UO_559 (O_559,N_14948,N_14776);
or UO_560 (O_560,N_14799,N_14769);
nor UO_561 (O_561,N_14799,N_14747);
or UO_562 (O_562,N_14787,N_14974);
and UO_563 (O_563,N_14977,N_14844);
nor UO_564 (O_564,N_14909,N_14774);
nor UO_565 (O_565,N_14832,N_14885);
nor UO_566 (O_566,N_14970,N_14937);
nor UO_567 (O_567,N_14727,N_14874);
nand UO_568 (O_568,N_14953,N_14844);
or UO_569 (O_569,N_14895,N_14958);
or UO_570 (O_570,N_14824,N_14873);
nand UO_571 (O_571,N_14782,N_14784);
nor UO_572 (O_572,N_14947,N_14755);
nand UO_573 (O_573,N_14951,N_14701);
xnor UO_574 (O_574,N_14879,N_14755);
xnor UO_575 (O_575,N_14823,N_14744);
and UO_576 (O_576,N_14896,N_14929);
nor UO_577 (O_577,N_14952,N_14832);
nor UO_578 (O_578,N_14896,N_14925);
nand UO_579 (O_579,N_14778,N_14923);
nand UO_580 (O_580,N_14708,N_14714);
nor UO_581 (O_581,N_14767,N_14823);
nor UO_582 (O_582,N_14851,N_14826);
and UO_583 (O_583,N_14934,N_14846);
nor UO_584 (O_584,N_14961,N_14869);
xor UO_585 (O_585,N_14994,N_14850);
or UO_586 (O_586,N_14784,N_14943);
or UO_587 (O_587,N_14742,N_14832);
nor UO_588 (O_588,N_14929,N_14826);
xnor UO_589 (O_589,N_14791,N_14978);
nor UO_590 (O_590,N_14881,N_14818);
xor UO_591 (O_591,N_14901,N_14922);
and UO_592 (O_592,N_14796,N_14752);
nand UO_593 (O_593,N_14713,N_14765);
or UO_594 (O_594,N_14920,N_14720);
xnor UO_595 (O_595,N_14812,N_14708);
nor UO_596 (O_596,N_14929,N_14725);
and UO_597 (O_597,N_14713,N_14991);
nand UO_598 (O_598,N_14760,N_14734);
or UO_599 (O_599,N_14833,N_14950);
and UO_600 (O_600,N_14712,N_14709);
xor UO_601 (O_601,N_14883,N_14909);
or UO_602 (O_602,N_14788,N_14944);
nand UO_603 (O_603,N_14997,N_14879);
xor UO_604 (O_604,N_14784,N_14850);
xor UO_605 (O_605,N_14709,N_14948);
xnor UO_606 (O_606,N_14833,N_14852);
and UO_607 (O_607,N_14718,N_14986);
xor UO_608 (O_608,N_14901,N_14999);
nand UO_609 (O_609,N_14744,N_14904);
and UO_610 (O_610,N_14978,N_14770);
and UO_611 (O_611,N_14911,N_14754);
xor UO_612 (O_612,N_14806,N_14846);
nand UO_613 (O_613,N_14942,N_14743);
nor UO_614 (O_614,N_14736,N_14854);
nand UO_615 (O_615,N_14712,N_14869);
xor UO_616 (O_616,N_14846,N_14841);
nor UO_617 (O_617,N_14990,N_14831);
nand UO_618 (O_618,N_14976,N_14796);
nor UO_619 (O_619,N_14977,N_14801);
nor UO_620 (O_620,N_14741,N_14937);
or UO_621 (O_621,N_14715,N_14738);
or UO_622 (O_622,N_14826,N_14744);
or UO_623 (O_623,N_14947,N_14895);
and UO_624 (O_624,N_14810,N_14967);
nor UO_625 (O_625,N_14752,N_14836);
and UO_626 (O_626,N_14970,N_14796);
nor UO_627 (O_627,N_14752,N_14827);
nor UO_628 (O_628,N_14971,N_14944);
or UO_629 (O_629,N_14906,N_14871);
or UO_630 (O_630,N_14970,N_14924);
and UO_631 (O_631,N_14993,N_14744);
and UO_632 (O_632,N_14739,N_14761);
nand UO_633 (O_633,N_14859,N_14778);
nor UO_634 (O_634,N_14770,N_14984);
nand UO_635 (O_635,N_14914,N_14826);
xor UO_636 (O_636,N_14812,N_14959);
and UO_637 (O_637,N_14874,N_14997);
xnor UO_638 (O_638,N_14731,N_14866);
and UO_639 (O_639,N_14974,N_14933);
and UO_640 (O_640,N_14888,N_14733);
xnor UO_641 (O_641,N_14831,N_14950);
nand UO_642 (O_642,N_14761,N_14826);
or UO_643 (O_643,N_14979,N_14993);
and UO_644 (O_644,N_14895,N_14882);
xor UO_645 (O_645,N_14829,N_14792);
or UO_646 (O_646,N_14721,N_14839);
nand UO_647 (O_647,N_14830,N_14899);
or UO_648 (O_648,N_14755,N_14977);
and UO_649 (O_649,N_14905,N_14923);
or UO_650 (O_650,N_14995,N_14945);
and UO_651 (O_651,N_14836,N_14862);
and UO_652 (O_652,N_14841,N_14997);
nor UO_653 (O_653,N_14848,N_14704);
and UO_654 (O_654,N_14765,N_14742);
or UO_655 (O_655,N_14896,N_14723);
or UO_656 (O_656,N_14779,N_14718);
or UO_657 (O_657,N_14934,N_14878);
or UO_658 (O_658,N_14734,N_14823);
nand UO_659 (O_659,N_14803,N_14852);
xnor UO_660 (O_660,N_14702,N_14862);
or UO_661 (O_661,N_14928,N_14759);
and UO_662 (O_662,N_14760,N_14946);
and UO_663 (O_663,N_14819,N_14906);
xnor UO_664 (O_664,N_14891,N_14934);
or UO_665 (O_665,N_14975,N_14910);
xor UO_666 (O_666,N_14701,N_14839);
nand UO_667 (O_667,N_14897,N_14745);
xor UO_668 (O_668,N_14701,N_14950);
xor UO_669 (O_669,N_14720,N_14978);
nand UO_670 (O_670,N_14847,N_14894);
nand UO_671 (O_671,N_14807,N_14902);
nand UO_672 (O_672,N_14875,N_14945);
or UO_673 (O_673,N_14956,N_14828);
nor UO_674 (O_674,N_14964,N_14729);
xnor UO_675 (O_675,N_14712,N_14807);
nand UO_676 (O_676,N_14889,N_14875);
xor UO_677 (O_677,N_14880,N_14701);
and UO_678 (O_678,N_14739,N_14879);
and UO_679 (O_679,N_14863,N_14785);
nor UO_680 (O_680,N_14891,N_14971);
and UO_681 (O_681,N_14981,N_14749);
and UO_682 (O_682,N_14789,N_14866);
nand UO_683 (O_683,N_14781,N_14815);
nor UO_684 (O_684,N_14938,N_14864);
nor UO_685 (O_685,N_14799,N_14821);
and UO_686 (O_686,N_14862,N_14975);
nor UO_687 (O_687,N_14978,N_14705);
nand UO_688 (O_688,N_14738,N_14994);
nand UO_689 (O_689,N_14941,N_14918);
or UO_690 (O_690,N_14904,N_14968);
xor UO_691 (O_691,N_14712,N_14734);
xnor UO_692 (O_692,N_14813,N_14814);
and UO_693 (O_693,N_14923,N_14845);
nand UO_694 (O_694,N_14830,N_14826);
and UO_695 (O_695,N_14962,N_14976);
or UO_696 (O_696,N_14839,N_14741);
nand UO_697 (O_697,N_14897,N_14734);
xnor UO_698 (O_698,N_14796,N_14965);
xnor UO_699 (O_699,N_14905,N_14924);
nor UO_700 (O_700,N_14851,N_14859);
xnor UO_701 (O_701,N_14984,N_14726);
xnor UO_702 (O_702,N_14998,N_14743);
and UO_703 (O_703,N_14965,N_14985);
xor UO_704 (O_704,N_14861,N_14738);
nand UO_705 (O_705,N_14998,N_14826);
and UO_706 (O_706,N_14788,N_14811);
xnor UO_707 (O_707,N_14959,N_14739);
nand UO_708 (O_708,N_14710,N_14925);
nor UO_709 (O_709,N_14727,N_14744);
nor UO_710 (O_710,N_14718,N_14973);
xnor UO_711 (O_711,N_14987,N_14968);
nor UO_712 (O_712,N_14990,N_14783);
and UO_713 (O_713,N_14953,N_14712);
xor UO_714 (O_714,N_14975,N_14791);
xor UO_715 (O_715,N_14753,N_14880);
nand UO_716 (O_716,N_14703,N_14714);
xnor UO_717 (O_717,N_14806,N_14713);
and UO_718 (O_718,N_14715,N_14748);
and UO_719 (O_719,N_14785,N_14943);
nor UO_720 (O_720,N_14713,N_14916);
xor UO_721 (O_721,N_14759,N_14984);
or UO_722 (O_722,N_14979,N_14930);
and UO_723 (O_723,N_14817,N_14891);
xor UO_724 (O_724,N_14830,N_14733);
nor UO_725 (O_725,N_14845,N_14780);
nand UO_726 (O_726,N_14948,N_14967);
xnor UO_727 (O_727,N_14902,N_14704);
and UO_728 (O_728,N_14716,N_14858);
xor UO_729 (O_729,N_14725,N_14760);
nor UO_730 (O_730,N_14884,N_14780);
or UO_731 (O_731,N_14837,N_14813);
or UO_732 (O_732,N_14750,N_14804);
and UO_733 (O_733,N_14992,N_14720);
or UO_734 (O_734,N_14757,N_14756);
xnor UO_735 (O_735,N_14865,N_14701);
or UO_736 (O_736,N_14963,N_14740);
nand UO_737 (O_737,N_14923,N_14857);
and UO_738 (O_738,N_14909,N_14969);
nand UO_739 (O_739,N_14712,N_14909);
nor UO_740 (O_740,N_14950,N_14859);
nor UO_741 (O_741,N_14994,N_14998);
or UO_742 (O_742,N_14814,N_14892);
nand UO_743 (O_743,N_14870,N_14939);
nor UO_744 (O_744,N_14984,N_14912);
xnor UO_745 (O_745,N_14890,N_14799);
nor UO_746 (O_746,N_14873,N_14963);
xnor UO_747 (O_747,N_14962,N_14923);
or UO_748 (O_748,N_14726,N_14892);
nor UO_749 (O_749,N_14790,N_14880);
and UO_750 (O_750,N_14899,N_14835);
xor UO_751 (O_751,N_14721,N_14974);
nor UO_752 (O_752,N_14845,N_14893);
or UO_753 (O_753,N_14805,N_14935);
and UO_754 (O_754,N_14918,N_14907);
and UO_755 (O_755,N_14943,N_14854);
nand UO_756 (O_756,N_14794,N_14848);
nand UO_757 (O_757,N_14949,N_14744);
xnor UO_758 (O_758,N_14914,N_14798);
xor UO_759 (O_759,N_14727,N_14717);
nand UO_760 (O_760,N_14905,N_14705);
xor UO_761 (O_761,N_14902,N_14978);
xnor UO_762 (O_762,N_14873,N_14842);
and UO_763 (O_763,N_14998,N_14806);
or UO_764 (O_764,N_14978,N_14871);
nand UO_765 (O_765,N_14879,N_14896);
nor UO_766 (O_766,N_14999,N_14855);
nand UO_767 (O_767,N_14712,N_14950);
nand UO_768 (O_768,N_14714,N_14756);
or UO_769 (O_769,N_14794,N_14713);
nor UO_770 (O_770,N_14999,N_14704);
or UO_771 (O_771,N_14995,N_14971);
nor UO_772 (O_772,N_14965,N_14763);
or UO_773 (O_773,N_14940,N_14854);
or UO_774 (O_774,N_14955,N_14902);
and UO_775 (O_775,N_14923,N_14806);
and UO_776 (O_776,N_14954,N_14854);
nor UO_777 (O_777,N_14748,N_14997);
or UO_778 (O_778,N_14746,N_14864);
nor UO_779 (O_779,N_14713,N_14862);
and UO_780 (O_780,N_14912,N_14892);
xnor UO_781 (O_781,N_14946,N_14778);
or UO_782 (O_782,N_14970,N_14804);
nor UO_783 (O_783,N_14845,N_14735);
nor UO_784 (O_784,N_14796,N_14916);
or UO_785 (O_785,N_14906,N_14787);
nand UO_786 (O_786,N_14716,N_14768);
and UO_787 (O_787,N_14802,N_14765);
nand UO_788 (O_788,N_14851,N_14764);
xor UO_789 (O_789,N_14952,N_14754);
xnor UO_790 (O_790,N_14863,N_14911);
nand UO_791 (O_791,N_14769,N_14784);
and UO_792 (O_792,N_14791,N_14790);
nand UO_793 (O_793,N_14820,N_14718);
nand UO_794 (O_794,N_14932,N_14758);
nor UO_795 (O_795,N_14830,N_14854);
or UO_796 (O_796,N_14999,N_14711);
or UO_797 (O_797,N_14762,N_14747);
nand UO_798 (O_798,N_14847,N_14941);
nor UO_799 (O_799,N_14764,N_14924);
xnor UO_800 (O_800,N_14858,N_14860);
nor UO_801 (O_801,N_14920,N_14802);
nor UO_802 (O_802,N_14770,N_14703);
xnor UO_803 (O_803,N_14959,N_14724);
nor UO_804 (O_804,N_14835,N_14788);
xnor UO_805 (O_805,N_14921,N_14834);
nor UO_806 (O_806,N_14936,N_14901);
xnor UO_807 (O_807,N_14735,N_14959);
or UO_808 (O_808,N_14822,N_14904);
xor UO_809 (O_809,N_14843,N_14811);
nand UO_810 (O_810,N_14755,N_14708);
or UO_811 (O_811,N_14750,N_14857);
or UO_812 (O_812,N_14787,N_14877);
nand UO_813 (O_813,N_14921,N_14803);
xnor UO_814 (O_814,N_14822,N_14888);
and UO_815 (O_815,N_14938,N_14927);
nor UO_816 (O_816,N_14899,N_14890);
or UO_817 (O_817,N_14826,N_14902);
nor UO_818 (O_818,N_14908,N_14985);
and UO_819 (O_819,N_14748,N_14765);
or UO_820 (O_820,N_14762,N_14817);
and UO_821 (O_821,N_14900,N_14849);
and UO_822 (O_822,N_14743,N_14879);
or UO_823 (O_823,N_14980,N_14848);
and UO_824 (O_824,N_14940,N_14974);
and UO_825 (O_825,N_14782,N_14818);
or UO_826 (O_826,N_14888,N_14973);
and UO_827 (O_827,N_14954,N_14942);
nand UO_828 (O_828,N_14764,N_14961);
nand UO_829 (O_829,N_14837,N_14756);
xnor UO_830 (O_830,N_14929,N_14809);
xor UO_831 (O_831,N_14705,N_14718);
nand UO_832 (O_832,N_14935,N_14867);
nor UO_833 (O_833,N_14864,N_14803);
xor UO_834 (O_834,N_14753,N_14702);
or UO_835 (O_835,N_14975,N_14933);
and UO_836 (O_836,N_14898,N_14980);
and UO_837 (O_837,N_14864,N_14988);
and UO_838 (O_838,N_14958,N_14936);
nor UO_839 (O_839,N_14916,N_14913);
nand UO_840 (O_840,N_14836,N_14961);
and UO_841 (O_841,N_14971,N_14706);
and UO_842 (O_842,N_14896,N_14946);
or UO_843 (O_843,N_14703,N_14999);
nand UO_844 (O_844,N_14763,N_14745);
or UO_845 (O_845,N_14916,N_14926);
and UO_846 (O_846,N_14982,N_14875);
nand UO_847 (O_847,N_14898,N_14871);
nor UO_848 (O_848,N_14765,N_14791);
or UO_849 (O_849,N_14810,N_14807);
nor UO_850 (O_850,N_14986,N_14762);
xnor UO_851 (O_851,N_14955,N_14911);
and UO_852 (O_852,N_14885,N_14772);
xnor UO_853 (O_853,N_14901,N_14737);
xnor UO_854 (O_854,N_14977,N_14739);
or UO_855 (O_855,N_14905,N_14876);
xnor UO_856 (O_856,N_14749,N_14789);
nand UO_857 (O_857,N_14958,N_14801);
and UO_858 (O_858,N_14735,N_14724);
xor UO_859 (O_859,N_14962,N_14716);
nor UO_860 (O_860,N_14843,N_14707);
or UO_861 (O_861,N_14778,N_14944);
nand UO_862 (O_862,N_14922,N_14781);
nand UO_863 (O_863,N_14976,N_14850);
or UO_864 (O_864,N_14915,N_14962);
nand UO_865 (O_865,N_14795,N_14724);
or UO_866 (O_866,N_14818,N_14754);
or UO_867 (O_867,N_14924,N_14980);
and UO_868 (O_868,N_14882,N_14783);
xor UO_869 (O_869,N_14726,N_14866);
nand UO_870 (O_870,N_14791,N_14835);
nand UO_871 (O_871,N_14807,N_14990);
nor UO_872 (O_872,N_14716,N_14804);
nand UO_873 (O_873,N_14998,N_14951);
xor UO_874 (O_874,N_14974,N_14903);
or UO_875 (O_875,N_14997,N_14984);
and UO_876 (O_876,N_14739,N_14799);
or UO_877 (O_877,N_14733,N_14805);
xnor UO_878 (O_878,N_14726,N_14790);
nor UO_879 (O_879,N_14818,N_14840);
nand UO_880 (O_880,N_14805,N_14737);
nor UO_881 (O_881,N_14753,N_14898);
nand UO_882 (O_882,N_14958,N_14883);
nand UO_883 (O_883,N_14845,N_14954);
or UO_884 (O_884,N_14885,N_14863);
nor UO_885 (O_885,N_14962,N_14932);
and UO_886 (O_886,N_14975,N_14894);
xor UO_887 (O_887,N_14821,N_14730);
xnor UO_888 (O_888,N_14788,N_14827);
xor UO_889 (O_889,N_14961,N_14765);
and UO_890 (O_890,N_14919,N_14745);
nand UO_891 (O_891,N_14727,N_14831);
nor UO_892 (O_892,N_14840,N_14952);
xor UO_893 (O_893,N_14772,N_14962);
nor UO_894 (O_894,N_14800,N_14979);
and UO_895 (O_895,N_14845,N_14781);
and UO_896 (O_896,N_14955,N_14753);
nor UO_897 (O_897,N_14753,N_14928);
and UO_898 (O_898,N_14907,N_14896);
and UO_899 (O_899,N_14784,N_14724);
nor UO_900 (O_900,N_14814,N_14872);
xor UO_901 (O_901,N_14908,N_14744);
xor UO_902 (O_902,N_14865,N_14944);
nand UO_903 (O_903,N_14853,N_14893);
xnor UO_904 (O_904,N_14996,N_14821);
and UO_905 (O_905,N_14849,N_14756);
nor UO_906 (O_906,N_14746,N_14791);
or UO_907 (O_907,N_14931,N_14838);
xor UO_908 (O_908,N_14956,N_14966);
nand UO_909 (O_909,N_14767,N_14974);
xor UO_910 (O_910,N_14817,N_14748);
nand UO_911 (O_911,N_14800,N_14853);
or UO_912 (O_912,N_14919,N_14757);
nand UO_913 (O_913,N_14920,N_14792);
nor UO_914 (O_914,N_14739,N_14778);
xor UO_915 (O_915,N_14979,N_14769);
nand UO_916 (O_916,N_14721,N_14844);
nor UO_917 (O_917,N_14789,N_14868);
and UO_918 (O_918,N_14952,N_14960);
nor UO_919 (O_919,N_14913,N_14962);
nor UO_920 (O_920,N_14973,N_14974);
xor UO_921 (O_921,N_14905,N_14837);
nor UO_922 (O_922,N_14923,N_14871);
and UO_923 (O_923,N_14915,N_14780);
xnor UO_924 (O_924,N_14752,N_14776);
nand UO_925 (O_925,N_14777,N_14752);
xor UO_926 (O_926,N_14772,N_14820);
xnor UO_927 (O_927,N_14960,N_14838);
and UO_928 (O_928,N_14946,N_14859);
nand UO_929 (O_929,N_14989,N_14975);
or UO_930 (O_930,N_14885,N_14980);
nor UO_931 (O_931,N_14814,N_14957);
xor UO_932 (O_932,N_14849,N_14822);
and UO_933 (O_933,N_14709,N_14988);
nand UO_934 (O_934,N_14810,N_14715);
nor UO_935 (O_935,N_14777,N_14977);
and UO_936 (O_936,N_14967,N_14889);
and UO_937 (O_937,N_14934,N_14919);
and UO_938 (O_938,N_14728,N_14886);
xor UO_939 (O_939,N_14980,N_14772);
or UO_940 (O_940,N_14707,N_14801);
nor UO_941 (O_941,N_14904,N_14865);
xnor UO_942 (O_942,N_14909,N_14889);
or UO_943 (O_943,N_14914,N_14975);
and UO_944 (O_944,N_14738,N_14904);
nand UO_945 (O_945,N_14807,N_14816);
nor UO_946 (O_946,N_14989,N_14959);
nor UO_947 (O_947,N_14977,N_14927);
nor UO_948 (O_948,N_14865,N_14819);
nand UO_949 (O_949,N_14744,N_14729);
nand UO_950 (O_950,N_14921,N_14779);
xnor UO_951 (O_951,N_14898,N_14976);
nand UO_952 (O_952,N_14831,N_14816);
xor UO_953 (O_953,N_14862,N_14775);
nor UO_954 (O_954,N_14832,N_14975);
xnor UO_955 (O_955,N_14797,N_14818);
or UO_956 (O_956,N_14977,N_14815);
or UO_957 (O_957,N_14962,N_14731);
xnor UO_958 (O_958,N_14929,N_14870);
nand UO_959 (O_959,N_14871,N_14885);
nor UO_960 (O_960,N_14778,N_14964);
or UO_961 (O_961,N_14953,N_14926);
or UO_962 (O_962,N_14770,N_14946);
xnor UO_963 (O_963,N_14917,N_14918);
nand UO_964 (O_964,N_14933,N_14987);
nand UO_965 (O_965,N_14992,N_14866);
nand UO_966 (O_966,N_14885,N_14764);
xor UO_967 (O_967,N_14724,N_14793);
nor UO_968 (O_968,N_14774,N_14975);
nand UO_969 (O_969,N_14937,N_14710);
nor UO_970 (O_970,N_14940,N_14768);
nor UO_971 (O_971,N_14824,N_14749);
and UO_972 (O_972,N_14835,N_14807);
or UO_973 (O_973,N_14847,N_14850);
xor UO_974 (O_974,N_14926,N_14740);
nand UO_975 (O_975,N_14908,N_14780);
nor UO_976 (O_976,N_14725,N_14950);
xnor UO_977 (O_977,N_14770,N_14899);
nand UO_978 (O_978,N_14717,N_14792);
and UO_979 (O_979,N_14958,N_14731);
xor UO_980 (O_980,N_14766,N_14724);
xor UO_981 (O_981,N_14992,N_14762);
xnor UO_982 (O_982,N_14738,N_14977);
or UO_983 (O_983,N_14993,N_14803);
nor UO_984 (O_984,N_14975,N_14750);
nand UO_985 (O_985,N_14783,N_14737);
or UO_986 (O_986,N_14733,N_14932);
nor UO_987 (O_987,N_14983,N_14807);
nor UO_988 (O_988,N_14783,N_14971);
xor UO_989 (O_989,N_14727,N_14829);
and UO_990 (O_990,N_14880,N_14711);
and UO_991 (O_991,N_14979,N_14917);
xor UO_992 (O_992,N_14997,N_14790);
or UO_993 (O_993,N_14910,N_14759);
xnor UO_994 (O_994,N_14979,N_14898);
nand UO_995 (O_995,N_14826,N_14701);
xnor UO_996 (O_996,N_14777,N_14967);
xor UO_997 (O_997,N_14701,N_14954);
or UO_998 (O_998,N_14715,N_14759);
nand UO_999 (O_999,N_14784,N_14818);
xnor UO_1000 (O_1000,N_14866,N_14796);
or UO_1001 (O_1001,N_14953,N_14756);
xor UO_1002 (O_1002,N_14977,N_14782);
and UO_1003 (O_1003,N_14810,N_14868);
xnor UO_1004 (O_1004,N_14803,N_14941);
and UO_1005 (O_1005,N_14941,N_14984);
nand UO_1006 (O_1006,N_14855,N_14781);
nand UO_1007 (O_1007,N_14765,N_14777);
and UO_1008 (O_1008,N_14724,N_14883);
nand UO_1009 (O_1009,N_14839,N_14712);
and UO_1010 (O_1010,N_14819,N_14830);
nor UO_1011 (O_1011,N_14902,N_14864);
or UO_1012 (O_1012,N_14814,N_14890);
and UO_1013 (O_1013,N_14733,N_14867);
nand UO_1014 (O_1014,N_14774,N_14864);
xor UO_1015 (O_1015,N_14938,N_14998);
or UO_1016 (O_1016,N_14835,N_14918);
nor UO_1017 (O_1017,N_14993,N_14708);
or UO_1018 (O_1018,N_14895,N_14734);
nand UO_1019 (O_1019,N_14980,N_14709);
nand UO_1020 (O_1020,N_14851,N_14715);
nand UO_1021 (O_1021,N_14853,N_14873);
nand UO_1022 (O_1022,N_14872,N_14795);
nor UO_1023 (O_1023,N_14805,N_14921);
or UO_1024 (O_1024,N_14921,N_14915);
or UO_1025 (O_1025,N_14870,N_14982);
xor UO_1026 (O_1026,N_14975,N_14848);
and UO_1027 (O_1027,N_14889,N_14820);
nor UO_1028 (O_1028,N_14845,N_14947);
nor UO_1029 (O_1029,N_14919,N_14728);
nand UO_1030 (O_1030,N_14899,N_14750);
or UO_1031 (O_1031,N_14759,N_14929);
nand UO_1032 (O_1032,N_14974,N_14745);
nand UO_1033 (O_1033,N_14851,N_14984);
nor UO_1034 (O_1034,N_14973,N_14875);
or UO_1035 (O_1035,N_14828,N_14839);
nor UO_1036 (O_1036,N_14742,N_14793);
nor UO_1037 (O_1037,N_14972,N_14983);
nor UO_1038 (O_1038,N_14953,N_14733);
nor UO_1039 (O_1039,N_14937,N_14721);
nand UO_1040 (O_1040,N_14866,N_14954);
or UO_1041 (O_1041,N_14825,N_14895);
xnor UO_1042 (O_1042,N_14725,N_14966);
or UO_1043 (O_1043,N_14933,N_14957);
nor UO_1044 (O_1044,N_14708,N_14985);
nand UO_1045 (O_1045,N_14708,N_14934);
and UO_1046 (O_1046,N_14708,N_14969);
xnor UO_1047 (O_1047,N_14859,N_14841);
nor UO_1048 (O_1048,N_14989,N_14976);
nand UO_1049 (O_1049,N_14952,N_14760);
nand UO_1050 (O_1050,N_14780,N_14947);
xor UO_1051 (O_1051,N_14976,N_14740);
nor UO_1052 (O_1052,N_14795,N_14928);
and UO_1053 (O_1053,N_14840,N_14856);
or UO_1054 (O_1054,N_14819,N_14800);
xor UO_1055 (O_1055,N_14842,N_14815);
nor UO_1056 (O_1056,N_14878,N_14724);
xnor UO_1057 (O_1057,N_14803,N_14956);
xnor UO_1058 (O_1058,N_14904,N_14940);
nor UO_1059 (O_1059,N_14703,N_14921);
xor UO_1060 (O_1060,N_14708,N_14853);
or UO_1061 (O_1061,N_14875,N_14863);
and UO_1062 (O_1062,N_14863,N_14920);
xor UO_1063 (O_1063,N_14906,N_14794);
nand UO_1064 (O_1064,N_14982,N_14999);
nand UO_1065 (O_1065,N_14976,N_14840);
and UO_1066 (O_1066,N_14925,N_14807);
nor UO_1067 (O_1067,N_14821,N_14707);
nor UO_1068 (O_1068,N_14789,N_14933);
xor UO_1069 (O_1069,N_14834,N_14906);
and UO_1070 (O_1070,N_14828,N_14750);
xor UO_1071 (O_1071,N_14815,N_14735);
and UO_1072 (O_1072,N_14759,N_14814);
xnor UO_1073 (O_1073,N_14933,N_14831);
and UO_1074 (O_1074,N_14884,N_14789);
and UO_1075 (O_1075,N_14937,N_14892);
and UO_1076 (O_1076,N_14747,N_14817);
or UO_1077 (O_1077,N_14946,N_14939);
or UO_1078 (O_1078,N_14979,N_14803);
and UO_1079 (O_1079,N_14996,N_14786);
and UO_1080 (O_1080,N_14901,N_14850);
or UO_1081 (O_1081,N_14965,N_14891);
or UO_1082 (O_1082,N_14844,N_14830);
or UO_1083 (O_1083,N_14854,N_14944);
or UO_1084 (O_1084,N_14780,N_14818);
nor UO_1085 (O_1085,N_14976,N_14951);
nor UO_1086 (O_1086,N_14744,N_14857);
xor UO_1087 (O_1087,N_14715,N_14849);
or UO_1088 (O_1088,N_14708,N_14749);
or UO_1089 (O_1089,N_14864,N_14888);
nand UO_1090 (O_1090,N_14905,N_14928);
nand UO_1091 (O_1091,N_14776,N_14724);
or UO_1092 (O_1092,N_14778,N_14920);
and UO_1093 (O_1093,N_14963,N_14816);
xnor UO_1094 (O_1094,N_14729,N_14842);
nor UO_1095 (O_1095,N_14706,N_14819);
nor UO_1096 (O_1096,N_14847,N_14796);
and UO_1097 (O_1097,N_14874,N_14713);
nor UO_1098 (O_1098,N_14936,N_14755);
and UO_1099 (O_1099,N_14966,N_14708);
or UO_1100 (O_1100,N_14735,N_14805);
nand UO_1101 (O_1101,N_14967,N_14736);
or UO_1102 (O_1102,N_14715,N_14957);
and UO_1103 (O_1103,N_14904,N_14838);
nor UO_1104 (O_1104,N_14991,N_14963);
nor UO_1105 (O_1105,N_14742,N_14777);
nand UO_1106 (O_1106,N_14791,N_14868);
xor UO_1107 (O_1107,N_14987,N_14939);
nor UO_1108 (O_1108,N_14724,N_14777);
nor UO_1109 (O_1109,N_14952,N_14919);
and UO_1110 (O_1110,N_14920,N_14737);
and UO_1111 (O_1111,N_14757,N_14773);
xor UO_1112 (O_1112,N_14878,N_14942);
nor UO_1113 (O_1113,N_14777,N_14889);
or UO_1114 (O_1114,N_14995,N_14769);
nor UO_1115 (O_1115,N_14721,N_14900);
nor UO_1116 (O_1116,N_14930,N_14740);
or UO_1117 (O_1117,N_14774,N_14908);
nor UO_1118 (O_1118,N_14880,N_14887);
nor UO_1119 (O_1119,N_14923,N_14897);
or UO_1120 (O_1120,N_14724,N_14965);
nor UO_1121 (O_1121,N_14879,N_14868);
nor UO_1122 (O_1122,N_14858,N_14722);
nand UO_1123 (O_1123,N_14956,N_14953);
nor UO_1124 (O_1124,N_14855,N_14788);
xor UO_1125 (O_1125,N_14863,N_14893);
or UO_1126 (O_1126,N_14886,N_14752);
nand UO_1127 (O_1127,N_14826,N_14978);
nand UO_1128 (O_1128,N_14829,N_14775);
nand UO_1129 (O_1129,N_14792,N_14974);
nand UO_1130 (O_1130,N_14982,N_14758);
and UO_1131 (O_1131,N_14728,N_14799);
nand UO_1132 (O_1132,N_14801,N_14942);
and UO_1133 (O_1133,N_14925,N_14949);
or UO_1134 (O_1134,N_14826,N_14986);
nand UO_1135 (O_1135,N_14719,N_14865);
xnor UO_1136 (O_1136,N_14926,N_14862);
or UO_1137 (O_1137,N_14821,N_14793);
or UO_1138 (O_1138,N_14917,N_14762);
and UO_1139 (O_1139,N_14822,N_14837);
nand UO_1140 (O_1140,N_14862,N_14965);
and UO_1141 (O_1141,N_14868,N_14836);
nand UO_1142 (O_1142,N_14809,N_14790);
nand UO_1143 (O_1143,N_14747,N_14746);
and UO_1144 (O_1144,N_14744,N_14925);
or UO_1145 (O_1145,N_14883,N_14989);
nor UO_1146 (O_1146,N_14796,N_14927);
nor UO_1147 (O_1147,N_14821,N_14831);
nor UO_1148 (O_1148,N_14977,N_14898);
xor UO_1149 (O_1149,N_14942,N_14811);
or UO_1150 (O_1150,N_14780,N_14724);
xnor UO_1151 (O_1151,N_14802,N_14730);
or UO_1152 (O_1152,N_14951,N_14931);
xor UO_1153 (O_1153,N_14899,N_14714);
xnor UO_1154 (O_1154,N_14700,N_14725);
nand UO_1155 (O_1155,N_14831,N_14862);
and UO_1156 (O_1156,N_14862,N_14754);
nand UO_1157 (O_1157,N_14935,N_14754);
nor UO_1158 (O_1158,N_14925,N_14862);
and UO_1159 (O_1159,N_14873,N_14720);
nand UO_1160 (O_1160,N_14948,N_14901);
nand UO_1161 (O_1161,N_14939,N_14826);
nand UO_1162 (O_1162,N_14773,N_14812);
or UO_1163 (O_1163,N_14956,N_14731);
nand UO_1164 (O_1164,N_14949,N_14717);
nor UO_1165 (O_1165,N_14983,N_14882);
nor UO_1166 (O_1166,N_14726,N_14762);
or UO_1167 (O_1167,N_14784,N_14897);
or UO_1168 (O_1168,N_14918,N_14744);
nand UO_1169 (O_1169,N_14727,N_14701);
xor UO_1170 (O_1170,N_14704,N_14762);
xnor UO_1171 (O_1171,N_14893,N_14889);
nor UO_1172 (O_1172,N_14824,N_14953);
nand UO_1173 (O_1173,N_14749,N_14751);
and UO_1174 (O_1174,N_14890,N_14715);
or UO_1175 (O_1175,N_14962,N_14805);
or UO_1176 (O_1176,N_14736,N_14892);
or UO_1177 (O_1177,N_14949,N_14794);
and UO_1178 (O_1178,N_14998,N_14823);
nand UO_1179 (O_1179,N_14822,N_14809);
or UO_1180 (O_1180,N_14857,N_14726);
and UO_1181 (O_1181,N_14915,N_14828);
and UO_1182 (O_1182,N_14890,N_14989);
nor UO_1183 (O_1183,N_14706,N_14738);
and UO_1184 (O_1184,N_14822,N_14732);
or UO_1185 (O_1185,N_14826,N_14854);
or UO_1186 (O_1186,N_14978,N_14869);
and UO_1187 (O_1187,N_14781,N_14859);
and UO_1188 (O_1188,N_14755,N_14990);
or UO_1189 (O_1189,N_14910,N_14828);
or UO_1190 (O_1190,N_14829,N_14706);
and UO_1191 (O_1191,N_14909,N_14751);
xnor UO_1192 (O_1192,N_14870,N_14815);
and UO_1193 (O_1193,N_14752,N_14757);
and UO_1194 (O_1194,N_14976,N_14703);
nand UO_1195 (O_1195,N_14804,N_14904);
or UO_1196 (O_1196,N_14778,N_14912);
and UO_1197 (O_1197,N_14919,N_14893);
and UO_1198 (O_1198,N_14722,N_14844);
and UO_1199 (O_1199,N_14722,N_14962);
xnor UO_1200 (O_1200,N_14726,N_14811);
xnor UO_1201 (O_1201,N_14784,N_14884);
nor UO_1202 (O_1202,N_14941,N_14870);
and UO_1203 (O_1203,N_14906,N_14839);
nor UO_1204 (O_1204,N_14860,N_14958);
or UO_1205 (O_1205,N_14894,N_14754);
or UO_1206 (O_1206,N_14994,N_14977);
nand UO_1207 (O_1207,N_14721,N_14858);
xnor UO_1208 (O_1208,N_14886,N_14715);
nand UO_1209 (O_1209,N_14704,N_14732);
and UO_1210 (O_1210,N_14755,N_14960);
nand UO_1211 (O_1211,N_14961,N_14843);
nor UO_1212 (O_1212,N_14766,N_14933);
nand UO_1213 (O_1213,N_14952,N_14897);
xor UO_1214 (O_1214,N_14722,N_14728);
nand UO_1215 (O_1215,N_14995,N_14701);
and UO_1216 (O_1216,N_14719,N_14961);
or UO_1217 (O_1217,N_14765,N_14947);
nor UO_1218 (O_1218,N_14860,N_14743);
xnor UO_1219 (O_1219,N_14954,N_14892);
and UO_1220 (O_1220,N_14939,N_14865);
and UO_1221 (O_1221,N_14765,N_14972);
and UO_1222 (O_1222,N_14950,N_14751);
nor UO_1223 (O_1223,N_14971,N_14859);
nand UO_1224 (O_1224,N_14925,N_14882);
nor UO_1225 (O_1225,N_14948,N_14914);
xnor UO_1226 (O_1226,N_14793,N_14702);
or UO_1227 (O_1227,N_14700,N_14793);
nor UO_1228 (O_1228,N_14921,N_14711);
nor UO_1229 (O_1229,N_14747,N_14859);
xnor UO_1230 (O_1230,N_14743,N_14768);
nand UO_1231 (O_1231,N_14887,N_14787);
and UO_1232 (O_1232,N_14729,N_14909);
and UO_1233 (O_1233,N_14939,N_14759);
nor UO_1234 (O_1234,N_14889,N_14957);
nor UO_1235 (O_1235,N_14972,N_14784);
or UO_1236 (O_1236,N_14722,N_14997);
or UO_1237 (O_1237,N_14836,N_14851);
nand UO_1238 (O_1238,N_14972,N_14713);
or UO_1239 (O_1239,N_14838,N_14825);
nor UO_1240 (O_1240,N_14723,N_14703);
or UO_1241 (O_1241,N_14892,N_14865);
nor UO_1242 (O_1242,N_14738,N_14758);
xor UO_1243 (O_1243,N_14793,N_14984);
nor UO_1244 (O_1244,N_14805,N_14818);
nand UO_1245 (O_1245,N_14858,N_14973);
nand UO_1246 (O_1246,N_14772,N_14735);
and UO_1247 (O_1247,N_14837,N_14910);
xor UO_1248 (O_1248,N_14971,N_14873);
nor UO_1249 (O_1249,N_14739,N_14707);
xnor UO_1250 (O_1250,N_14838,N_14715);
and UO_1251 (O_1251,N_14799,N_14899);
and UO_1252 (O_1252,N_14712,N_14855);
and UO_1253 (O_1253,N_14982,N_14730);
and UO_1254 (O_1254,N_14709,N_14743);
and UO_1255 (O_1255,N_14888,N_14911);
nand UO_1256 (O_1256,N_14953,N_14959);
nand UO_1257 (O_1257,N_14821,N_14752);
xnor UO_1258 (O_1258,N_14731,N_14894);
or UO_1259 (O_1259,N_14972,N_14951);
nor UO_1260 (O_1260,N_14703,N_14713);
xnor UO_1261 (O_1261,N_14970,N_14861);
or UO_1262 (O_1262,N_14864,N_14823);
or UO_1263 (O_1263,N_14783,N_14754);
or UO_1264 (O_1264,N_14894,N_14954);
or UO_1265 (O_1265,N_14982,N_14941);
nand UO_1266 (O_1266,N_14997,N_14721);
nor UO_1267 (O_1267,N_14772,N_14811);
and UO_1268 (O_1268,N_14937,N_14730);
nand UO_1269 (O_1269,N_14886,N_14813);
nand UO_1270 (O_1270,N_14887,N_14757);
nor UO_1271 (O_1271,N_14923,N_14732);
or UO_1272 (O_1272,N_14787,N_14748);
or UO_1273 (O_1273,N_14716,N_14955);
nand UO_1274 (O_1274,N_14974,N_14971);
nand UO_1275 (O_1275,N_14740,N_14977);
or UO_1276 (O_1276,N_14954,N_14751);
xor UO_1277 (O_1277,N_14952,N_14959);
or UO_1278 (O_1278,N_14934,N_14887);
or UO_1279 (O_1279,N_14811,N_14834);
and UO_1280 (O_1280,N_14793,N_14956);
and UO_1281 (O_1281,N_14713,N_14971);
or UO_1282 (O_1282,N_14970,N_14862);
xnor UO_1283 (O_1283,N_14782,N_14734);
xor UO_1284 (O_1284,N_14933,N_14919);
nand UO_1285 (O_1285,N_14733,N_14804);
and UO_1286 (O_1286,N_14947,N_14799);
nand UO_1287 (O_1287,N_14889,N_14947);
nor UO_1288 (O_1288,N_14991,N_14853);
nand UO_1289 (O_1289,N_14923,N_14757);
xor UO_1290 (O_1290,N_14829,N_14837);
or UO_1291 (O_1291,N_14973,N_14711);
or UO_1292 (O_1292,N_14724,N_14860);
xnor UO_1293 (O_1293,N_14867,N_14878);
and UO_1294 (O_1294,N_14992,N_14977);
xnor UO_1295 (O_1295,N_14755,N_14999);
xnor UO_1296 (O_1296,N_14860,N_14941);
or UO_1297 (O_1297,N_14886,N_14853);
nor UO_1298 (O_1298,N_14932,N_14969);
and UO_1299 (O_1299,N_14785,N_14793);
or UO_1300 (O_1300,N_14766,N_14849);
or UO_1301 (O_1301,N_14883,N_14726);
and UO_1302 (O_1302,N_14828,N_14854);
and UO_1303 (O_1303,N_14767,N_14896);
or UO_1304 (O_1304,N_14718,N_14708);
nor UO_1305 (O_1305,N_14733,N_14971);
nand UO_1306 (O_1306,N_14836,N_14738);
xor UO_1307 (O_1307,N_14763,N_14754);
nor UO_1308 (O_1308,N_14713,N_14983);
xor UO_1309 (O_1309,N_14894,N_14743);
nor UO_1310 (O_1310,N_14872,N_14839);
xor UO_1311 (O_1311,N_14731,N_14987);
xor UO_1312 (O_1312,N_14776,N_14984);
xnor UO_1313 (O_1313,N_14702,N_14931);
nor UO_1314 (O_1314,N_14708,N_14737);
and UO_1315 (O_1315,N_14984,N_14930);
nand UO_1316 (O_1316,N_14742,N_14700);
nand UO_1317 (O_1317,N_14760,N_14747);
nor UO_1318 (O_1318,N_14906,N_14722);
xor UO_1319 (O_1319,N_14884,N_14733);
and UO_1320 (O_1320,N_14953,N_14752);
and UO_1321 (O_1321,N_14918,N_14931);
and UO_1322 (O_1322,N_14750,N_14759);
nand UO_1323 (O_1323,N_14958,N_14718);
or UO_1324 (O_1324,N_14973,N_14870);
or UO_1325 (O_1325,N_14715,N_14758);
nand UO_1326 (O_1326,N_14745,N_14998);
or UO_1327 (O_1327,N_14934,N_14761);
or UO_1328 (O_1328,N_14964,N_14848);
nand UO_1329 (O_1329,N_14969,N_14812);
and UO_1330 (O_1330,N_14809,N_14813);
and UO_1331 (O_1331,N_14812,N_14748);
and UO_1332 (O_1332,N_14939,N_14783);
or UO_1333 (O_1333,N_14749,N_14863);
nor UO_1334 (O_1334,N_14714,N_14746);
and UO_1335 (O_1335,N_14756,N_14735);
or UO_1336 (O_1336,N_14972,N_14979);
and UO_1337 (O_1337,N_14751,N_14884);
or UO_1338 (O_1338,N_14788,N_14850);
or UO_1339 (O_1339,N_14814,N_14891);
xnor UO_1340 (O_1340,N_14778,N_14702);
and UO_1341 (O_1341,N_14718,N_14807);
nand UO_1342 (O_1342,N_14765,N_14949);
nor UO_1343 (O_1343,N_14793,N_14801);
or UO_1344 (O_1344,N_14850,N_14979);
and UO_1345 (O_1345,N_14740,N_14750);
nor UO_1346 (O_1346,N_14884,N_14995);
nor UO_1347 (O_1347,N_14984,N_14801);
or UO_1348 (O_1348,N_14934,N_14885);
or UO_1349 (O_1349,N_14914,N_14873);
xor UO_1350 (O_1350,N_14819,N_14940);
nor UO_1351 (O_1351,N_14731,N_14717);
nor UO_1352 (O_1352,N_14740,N_14978);
nor UO_1353 (O_1353,N_14845,N_14861);
nor UO_1354 (O_1354,N_14995,N_14967);
and UO_1355 (O_1355,N_14700,N_14766);
and UO_1356 (O_1356,N_14859,N_14874);
xnor UO_1357 (O_1357,N_14808,N_14827);
nor UO_1358 (O_1358,N_14787,N_14750);
xor UO_1359 (O_1359,N_14981,N_14788);
nand UO_1360 (O_1360,N_14899,N_14992);
and UO_1361 (O_1361,N_14753,N_14946);
nor UO_1362 (O_1362,N_14725,N_14865);
nand UO_1363 (O_1363,N_14990,N_14951);
nand UO_1364 (O_1364,N_14956,N_14746);
or UO_1365 (O_1365,N_14902,N_14802);
xnor UO_1366 (O_1366,N_14786,N_14770);
and UO_1367 (O_1367,N_14990,N_14830);
nand UO_1368 (O_1368,N_14947,N_14783);
and UO_1369 (O_1369,N_14717,N_14896);
nand UO_1370 (O_1370,N_14734,N_14972);
xor UO_1371 (O_1371,N_14782,N_14736);
nor UO_1372 (O_1372,N_14853,N_14889);
or UO_1373 (O_1373,N_14846,N_14945);
and UO_1374 (O_1374,N_14887,N_14865);
or UO_1375 (O_1375,N_14914,N_14875);
nor UO_1376 (O_1376,N_14704,N_14861);
nor UO_1377 (O_1377,N_14710,N_14772);
nand UO_1378 (O_1378,N_14779,N_14738);
nand UO_1379 (O_1379,N_14772,N_14782);
xnor UO_1380 (O_1380,N_14946,N_14841);
or UO_1381 (O_1381,N_14796,N_14747);
xor UO_1382 (O_1382,N_14742,N_14776);
and UO_1383 (O_1383,N_14847,N_14813);
xnor UO_1384 (O_1384,N_14966,N_14950);
or UO_1385 (O_1385,N_14761,N_14908);
or UO_1386 (O_1386,N_14737,N_14781);
and UO_1387 (O_1387,N_14795,N_14847);
or UO_1388 (O_1388,N_14996,N_14950);
nand UO_1389 (O_1389,N_14906,N_14806);
or UO_1390 (O_1390,N_14859,N_14873);
nand UO_1391 (O_1391,N_14713,N_14925);
or UO_1392 (O_1392,N_14792,N_14784);
xnor UO_1393 (O_1393,N_14754,N_14778);
and UO_1394 (O_1394,N_14911,N_14914);
xor UO_1395 (O_1395,N_14973,N_14919);
and UO_1396 (O_1396,N_14709,N_14739);
nand UO_1397 (O_1397,N_14990,N_14967);
and UO_1398 (O_1398,N_14802,N_14703);
and UO_1399 (O_1399,N_14928,N_14790);
and UO_1400 (O_1400,N_14843,N_14924);
nor UO_1401 (O_1401,N_14835,N_14864);
nor UO_1402 (O_1402,N_14782,N_14749);
xor UO_1403 (O_1403,N_14937,N_14954);
xor UO_1404 (O_1404,N_14932,N_14728);
and UO_1405 (O_1405,N_14901,N_14944);
and UO_1406 (O_1406,N_14959,N_14975);
nor UO_1407 (O_1407,N_14830,N_14938);
nor UO_1408 (O_1408,N_14813,N_14974);
and UO_1409 (O_1409,N_14720,N_14874);
nand UO_1410 (O_1410,N_14894,N_14751);
nor UO_1411 (O_1411,N_14942,N_14948);
xnor UO_1412 (O_1412,N_14842,N_14863);
or UO_1413 (O_1413,N_14838,N_14760);
nor UO_1414 (O_1414,N_14729,N_14829);
or UO_1415 (O_1415,N_14791,N_14780);
or UO_1416 (O_1416,N_14721,N_14734);
and UO_1417 (O_1417,N_14974,N_14964);
and UO_1418 (O_1418,N_14868,N_14887);
nand UO_1419 (O_1419,N_14782,N_14866);
nor UO_1420 (O_1420,N_14780,N_14867);
nor UO_1421 (O_1421,N_14705,N_14859);
nor UO_1422 (O_1422,N_14710,N_14872);
xor UO_1423 (O_1423,N_14810,N_14955);
and UO_1424 (O_1424,N_14971,N_14702);
nand UO_1425 (O_1425,N_14896,N_14936);
nand UO_1426 (O_1426,N_14897,N_14990);
and UO_1427 (O_1427,N_14810,N_14776);
and UO_1428 (O_1428,N_14796,N_14890);
xnor UO_1429 (O_1429,N_14827,N_14735);
nand UO_1430 (O_1430,N_14998,N_14967);
and UO_1431 (O_1431,N_14731,N_14863);
and UO_1432 (O_1432,N_14836,N_14760);
nand UO_1433 (O_1433,N_14838,N_14965);
xor UO_1434 (O_1434,N_14831,N_14972);
nor UO_1435 (O_1435,N_14868,N_14961);
xnor UO_1436 (O_1436,N_14984,N_14977);
and UO_1437 (O_1437,N_14790,N_14707);
and UO_1438 (O_1438,N_14937,N_14945);
xor UO_1439 (O_1439,N_14757,N_14963);
nand UO_1440 (O_1440,N_14793,N_14875);
nand UO_1441 (O_1441,N_14849,N_14902);
nand UO_1442 (O_1442,N_14802,N_14906);
nand UO_1443 (O_1443,N_14996,N_14839);
and UO_1444 (O_1444,N_14732,N_14797);
xor UO_1445 (O_1445,N_14715,N_14995);
xor UO_1446 (O_1446,N_14963,N_14763);
or UO_1447 (O_1447,N_14791,N_14748);
nor UO_1448 (O_1448,N_14920,N_14961);
nor UO_1449 (O_1449,N_14851,N_14868);
and UO_1450 (O_1450,N_14990,N_14877);
and UO_1451 (O_1451,N_14822,N_14843);
nor UO_1452 (O_1452,N_14815,N_14739);
and UO_1453 (O_1453,N_14805,N_14812);
xnor UO_1454 (O_1454,N_14751,N_14718);
and UO_1455 (O_1455,N_14975,N_14797);
nor UO_1456 (O_1456,N_14756,N_14745);
xnor UO_1457 (O_1457,N_14732,N_14913);
nand UO_1458 (O_1458,N_14722,N_14756);
nor UO_1459 (O_1459,N_14735,N_14902);
or UO_1460 (O_1460,N_14856,N_14744);
or UO_1461 (O_1461,N_14905,N_14841);
nor UO_1462 (O_1462,N_14903,N_14775);
nor UO_1463 (O_1463,N_14862,N_14787);
or UO_1464 (O_1464,N_14879,N_14801);
nand UO_1465 (O_1465,N_14771,N_14722);
and UO_1466 (O_1466,N_14769,N_14917);
nor UO_1467 (O_1467,N_14764,N_14922);
or UO_1468 (O_1468,N_14952,N_14920);
nor UO_1469 (O_1469,N_14833,N_14920);
nor UO_1470 (O_1470,N_14792,N_14902);
xnor UO_1471 (O_1471,N_14902,N_14708);
or UO_1472 (O_1472,N_14910,N_14962);
nor UO_1473 (O_1473,N_14892,N_14873);
or UO_1474 (O_1474,N_14989,N_14916);
and UO_1475 (O_1475,N_14895,N_14981);
xor UO_1476 (O_1476,N_14809,N_14765);
and UO_1477 (O_1477,N_14986,N_14755);
nand UO_1478 (O_1478,N_14773,N_14911);
nand UO_1479 (O_1479,N_14770,N_14882);
or UO_1480 (O_1480,N_14937,N_14837);
nand UO_1481 (O_1481,N_14767,N_14934);
nand UO_1482 (O_1482,N_14776,N_14799);
or UO_1483 (O_1483,N_14714,N_14743);
xor UO_1484 (O_1484,N_14704,N_14922);
and UO_1485 (O_1485,N_14729,N_14911);
and UO_1486 (O_1486,N_14827,N_14783);
or UO_1487 (O_1487,N_14742,N_14797);
and UO_1488 (O_1488,N_14977,N_14858);
nor UO_1489 (O_1489,N_14907,N_14933);
and UO_1490 (O_1490,N_14800,N_14708);
xor UO_1491 (O_1491,N_14726,N_14992);
nor UO_1492 (O_1492,N_14819,N_14891);
and UO_1493 (O_1493,N_14787,N_14963);
nor UO_1494 (O_1494,N_14965,N_14770);
nand UO_1495 (O_1495,N_14793,N_14767);
and UO_1496 (O_1496,N_14828,N_14804);
nor UO_1497 (O_1497,N_14704,N_14863);
nand UO_1498 (O_1498,N_14795,N_14772);
or UO_1499 (O_1499,N_14798,N_14854);
nand UO_1500 (O_1500,N_14852,N_14926);
xor UO_1501 (O_1501,N_14869,N_14955);
and UO_1502 (O_1502,N_14913,N_14796);
and UO_1503 (O_1503,N_14860,N_14710);
nand UO_1504 (O_1504,N_14791,N_14998);
or UO_1505 (O_1505,N_14815,N_14795);
or UO_1506 (O_1506,N_14833,N_14777);
xnor UO_1507 (O_1507,N_14775,N_14828);
nand UO_1508 (O_1508,N_14738,N_14859);
xor UO_1509 (O_1509,N_14962,N_14800);
nor UO_1510 (O_1510,N_14783,N_14881);
nor UO_1511 (O_1511,N_14995,N_14907);
xnor UO_1512 (O_1512,N_14805,N_14774);
nor UO_1513 (O_1513,N_14875,N_14777);
and UO_1514 (O_1514,N_14787,N_14972);
and UO_1515 (O_1515,N_14839,N_14911);
nor UO_1516 (O_1516,N_14981,N_14802);
nor UO_1517 (O_1517,N_14839,N_14757);
or UO_1518 (O_1518,N_14757,N_14896);
nor UO_1519 (O_1519,N_14949,N_14988);
xor UO_1520 (O_1520,N_14783,N_14884);
and UO_1521 (O_1521,N_14885,N_14844);
nor UO_1522 (O_1522,N_14820,N_14701);
nand UO_1523 (O_1523,N_14739,N_14951);
nand UO_1524 (O_1524,N_14764,N_14860);
nand UO_1525 (O_1525,N_14895,N_14833);
xnor UO_1526 (O_1526,N_14995,N_14867);
xor UO_1527 (O_1527,N_14999,N_14997);
nand UO_1528 (O_1528,N_14838,N_14757);
or UO_1529 (O_1529,N_14939,N_14907);
and UO_1530 (O_1530,N_14712,N_14872);
nand UO_1531 (O_1531,N_14708,N_14823);
nor UO_1532 (O_1532,N_14820,N_14757);
xor UO_1533 (O_1533,N_14979,N_14946);
and UO_1534 (O_1534,N_14984,N_14781);
xnor UO_1535 (O_1535,N_14766,N_14923);
xnor UO_1536 (O_1536,N_14848,N_14979);
nand UO_1537 (O_1537,N_14773,N_14806);
and UO_1538 (O_1538,N_14885,N_14730);
nand UO_1539 (O_1539,N_14779,N_14986);
and UO_1540 (O_1540,N_14874,N_14968);
nor UO_1541 (O_1541,N_14843,N_14721);
xnor UO_1542 (O_1542,N_14892,N_14872);
or UO_1543 (O_1543,N_14958,N_14737);
nand UO_1544 (O_1544,N_14843,N_14833);
and UO_1545 (O_1545,N_14850,N_14772);
and UO_1546 (O_1546,N_14706,N_14933);
nand UO_1547 (O_1547,N_14796,N_14974);
xor UO_1548 (O_1548,N_14780,N_14865);
nor UO_1549 (O_1549,N_14783,N_14868);
or UO_1550 (O_1550,N_14778,N_14854);
nand UO_1551 (O_1551,N_14823,N_14866);
nor UO_1552 (O_1552,N_14955,N_14701);
nor UO_1553 (O_1553,N_14985,N_14809);
or UO_1554 (O_1554,N_14755,N_14831);
and UO_1555 (O_1555,N_14747,N_14896);
nor UO_1556 (O_1556,N_14879,N_14780);
nand UO_1557 (O_1557,N_14883,N_14901);
xnor UO_1558 (O_1558,N_14799,N_14794);
and UO_1559 (O_1559,N_14712,N_14731);
or UO_1560 (O_1560,N_14962,N_14832);
xor UO_1561 (O_1561,N_14883,N_14782);
xor UO_1562 (O_1562,N_14920,N_14983);
nand UO_1563 (O_1563,N_14905,N_14916);
xnor UO_1564 (O_1564,N_14759,N_14705);
or UO_1565 (O_1565,N_14740,N_14743);
or UO_1566 (O_1566,N_14922,N_14867);
nor UO_1567 (O_1567,N_14906,N_14715);
and UO_1568 (O_1568,N_14734,N_14847);
and UO_1569 (O_1569,N_14934,N_14774);
xor UO_1570 (O_1570,N_14844,N_14723);
or UO_1571 (O_1571,N_14747,N_14901);
nand UO_1572 (O_1572,N_14756,N_14851);
nand UO_1573 (O_1573,N_14706,N_14808);
nand UO_1574 (O_1574,N_14823,N_14712);
nor UO_1575 (O_1575,N_14955,N_14914);
xnor UO_1576 (O_1576,N_14708,N_14828);
nand UO_1577 (O_1577,N_14715,N_14746);
and UO_1578 (O_1578,N_14772,N_14725);
xnor UO_1579 (O_1579,N_14984,N_14840);
nor UO_1580 (O_1580,N_14739,N_14775);
nand UO_1581 (O_1581,N_14771,N_14829);
xnor UO_1582 (O_1582,N_14928,N_14920);
nor UO_1583 (O_1583,N_14986,N_14952);
or UO_1584 (O_1584,N_14972,N_14828);
nand UO_1585 (O_1585,N_14984,N_14971);
or UO_1586 (O_1586,N_14928,N_14712);
nor UO_1587 (O_1587,N_14954,N_14945);
nor UO_1588 (O_1588,N_14912,N_14800);
and UO_1589 (O_1589,N_14985,N_14883);
nor UO_1590 (O_1590,N_14989,N_14707);
nor UO_1591 (O_1591,N_14888,N_14740);
and UO_1592 (O_1592,N_14901,N_14733);
nand UO_1593 (O_1593,N_14770,N_14713);
and UO_1594 (O_1594,N_14721,N_14865);
or UO_1595 (O_1595,N_14978,N_14886);
and UO_1596 (O_1596,N_14941,N_14724);
xor UO_1597 (O_1597,N_14821,N_14747);
or UO_1598 (O_1598,N_14910,N_14970);
and UO_1599 (O_1599,N_14743,N_14924);
and UO_1600 (O_1600,N_14789,N_14875);
and UO_1601 (O_1601,N_14962,N_14938);
nor UO_1602 (O_1602,N_14870,N_14908);
nor UO_1603 (O_1603,N_14857,N_14898);
and UO_1604 (O_1604,N_14717,N_14829);
and UO_1605 (O_1605,N_14842,N_14966);
xnor UO_1606 (O_1606,N_14861,N_14901);
xnor UO_1607 (O_1607,N_14954,N_14934);
and UO_1608 (O_1608,N_14798,N_14960);
xor UO_1609 (O_1609,N_14762,N_14862);
nand UO_1610 (O_1610,N_14988,N_14993);
nand UO_1611 (O_1611,N_14809,N_14855);
nand UO_1612 (O_1612,N_14951,N_14856);
and UO_1613 (O_1613,N_14924,N_14922);
nor UO_1614 (O_1614,N_14761,N_14713);
and UO_1615 (O_1615,N_14924,N_14747);
nor UO_1616 (O_1616,N_14948,N_14806);
nor UO_1617 (O_1617,N_14895,N_14766);
nor UO_1618 (O_1618,N_14932,N_14872);
nor UO_1619 (O_1619,N_14860,N_14920);
or UO_1620 (O_1620,N_14739,N_14883);
xor UO_1621 (O_1621,N_14978,N_14926);
xnor UO_1622 (O_1622,N_14746,N_14907);
nor UO_1623 (O_1623,N_14993,N_14861);
nand UO_1624 (O_1624,N_14768,N_14702);
nor UO_1625 (O_1625,N_14991,N_14759);
nand UO_1626 (O_1626,N_14973,N_14798);
and UO_1627 (O_1627,N_14747,N_14906);
nand UO_1628 (O_1628,N_14763,N_14701);
nand UO_1629 (O_1629,N_14823,N_14780);
nor UO_1630 (O_1630,N_14823,N_14770);
nand UO_1631 (O_1631,N_14886,N_14822);
and UO_1632 (O_1632,N_14962,N_14837);
xor UO_1633 (O_1633,N_14812,N_14887);
xnor UO_1634 (O_1634,N_14850,N_14954);
nor UO_1635 (O_1635,N_14927,N_14737);
or UO_1636 (O_1636,N_14759,N_14793);
nor UO_1637 (O_1637,N_14990,N_14726);
nor UO_1638 (O_1638,N_14854,N_14981);
xnor UO_1639 (O_1639,N_14880,N_14731);
xnor UO_1640 (O_1640,N_14982,N_14954);
nor UO_1641 (O_1641,N_14800,N_14848);
and UO_1642 (O_1642,N_14722,N_14958);
or UO_1643 (O_1643,N_14846,N_14730);
nand UO_1644 (O_1644,N_14975,N_14842);
and UO_1645 (O_1645,N_14762,N_14975);
and UO_1646 (O_1646,N_14700,N_14759);
nand UO_1647 (O_1647,N_14930,N_14706);
nand UO_1648 (O_1648,N_14861,N_14769);
and UO_1649 (O_1649,N_14805,N_14744);
and UO_1650 (O_1650,N_14911,N_14861);
xnor UO_1651 (O_1651,N_14795,N_14940);
and UO_1652 (O_1652,N_14825,N_14747);
or UO_1653 (O_1653,N_14907,N_14910);
nand UO_1654 (O_1654,N_14890,N_14873);
xor UO_1655 (O_1655,N_14984,N_14891);
and UO_1656 (O_1656,N_14779,N_14870);
nor UO_1657 (O_1657,N_14705,N_14784);
and UO_1658 (O_1658,N_14761,N_14703);
or UO_1659 (O_1659,N_14929,N_14938);
and UO_1660 (O_1660,N_14839,N_14780);
xnor UO_1661 (O_1661,N_14842,N_14844);
and UO_1662 (O_1662,N_14724,N_14830);
nand UO_1663 (O_1663,N_14895,N_14846);
or UO_1664 (O_1664,N_14776,N_14779);
xnor UO_1665 (O_1665,N_14738,N_14802);
and UO_1666 (O_1666,N_14793,N_14755);
nand UO_1667 (O_1667,N_14753,N_14767);
and UO_1668 (O_1668,N_14737,N_14772);
and UO_1669 (O_1669,N_14980,N_14755);
nand UO_1670 (O_1670,N_14983,N_14926);
and UO_1671 (O_1671,N_14738,N_14990);
nor UO_1672 (O_1672,N_14947,N_14999);
nand UO_1673 (O_1673,N_14893,N_14723);
or UO_1674 (O_1674,N_14801,N_14774);
and UO_1675 (O_1675,N_14987,N_14929);
nand UO_1676 (O_1676,N_14852,N_14955);
nand UO_1677 (O_1677,N_14811,N_14792);
or UO_1678 (O_1678,N_14847,N_14784);
nand UO_1679 (O_1679,N_14840,N_14869);
or UO_1680 (O_1680,N_14923,N_14788);
xor UO_1681 (O_1681,N_14826,N_14994);
xor UO_1682 (O_1682,N_14999,N_14702);
xor UO_1683 (O_1683,N_14761,N_14889);
xor UO_1684 (O_1684,N_14993,N_14929);
and UO_1685 (O_1685,N_14748,N_14983);
nor UO_1686 (O_1686,N_14853,N_14849);
or UO_1687 (O_1687,N_14771,N_14930);
nor UO_1688 (O_1688,N_14720,N_14740);
nor UO_1689 (O_1689,N_14804,N_14727);
nand UO_1690 (O_1690,N_14898,N_14741);
nor UO_1691 (O_1691,N_14966,N_14884);
nand UO_1692 (O_1692,N_14856,N_14782);
and UO_1693 (O_1693,N_14878,N_14970);
or UO_1694 (O_1694,N_14703,N_14991);
and UO_1695 (O_1695,N_14840,N_14955);
and UO_1696 (O_1696,N_14732,N_14724);
xnor UO_1697 (O_1697,N_14997,N_14925);
nor UO_1698 (O_1698,N_14994,N_14757);
nand UO_1699 (O_1699,N_14994,N_14866);
nand UO_1700 (O_1700,N_14764,N_14748);
or UO_1701 (O_1701,N_14900,N_14763);
nand UO_1702 (O_1702,N_14744,N_14700);
xor UO_1703 (O_1703,N_14867,N_14823);
and UO_1704 (O_1704,N_14776,N_14959);
xor UO_1705 (O_1705,N_14987,N_14999);
nor UO_1706 (O_1706,N_14797,N_14791);
or UO_1707 (O_1707,N_14959,N_14731);
xor UO_1708 (O_1708,N_14799,N_14843);
nor UO_1709 (O_1709,N_14997,N_14915);
or UO_1710 (O_1710,N_14832,N_14806);
xnor UO_1711 (O_1711,N_14908,N_14823);
and UO_1712 (O_1712,N_14738,N_14889);
nor UO_1713 (O_1713,N_14700,N_14794);
nand UO_1714 (O_1714,N_14843,N_14860);
xnor UO_1715 (O_1715,N_14942,N_14927);
or UO_1716 (O_1716,N_14983,N_14896);
and UO_1717 (O_1717,N_14922,N_14939);
and UO_1718 (O_1718,N_14725,N_14827);
or UO_1719 (O_1719,N_14742,N_14799);
nor UO_1720 (O_1720,N_14926,N_14884);
xnor UO_1721 (O_1721,N_14880,N_14861);
nand UO_1722 (O_1722,N_14706,N_14817);
nand UO_1723 (O_1723,N_14836,N_14816);
xor UO_1724 (O_1724,N_14761,N_14978);
xor UO_1725 (O_1725,N_14718,N_14932);
xnor UO_1726 (O_1726,N_14760,N_14937);
xor UO_1727 (O_1727,N_14932,N_14980);
and UO_1728 (O_1728,N_14847,N_14853);
nor UO_1729 (O_1729,N_14822,N_14748);
and UO_1730 (O_1730,N_14716,N_14998);
xor UO_1731 (O_1731,N_14942,N_14850);
xnor UO_1732 (O_1732,N_14843,N_14940);
and UO_1733 (O_1733,N_14987,N_14740);
xor UO_1734 (O_1734,N_14844,N_14753);
nor UO_1735 (O_1735,N_14865,N_14731);
nand UO_1736 (O_1736,N_14932,N_14864);
or UO_1737 (O_1737,N_14945,N_14750);
nor UO_1738 (O_1738,N_14962,N_14965);
or UO_1739 (O_1739,N_14869,N_14757);
or UO_1740 (O_1740,N_14942,N_14720);
nor UO_1741 (O_1741,N_14895,N_14773);
and UO_1742 (O_1742,N_14890,N_14939);
and UO_1743 (O_1743,N_14917,N_14774);
and UO_1744 (O_1744,N_14944,N_14866);
xnor UO_1745 (O_1745,N_14808,N_14910);
nor UO_1746 (O_1746,N_14732,N_14753);
nand UO_1747 (O_1747,N_14746,N_14831);
nand UO_1748 (O_1748,N_14930,N_14803);
nor UO_1749 (O_1749,N_14785,N_14839);
nand UO_1750 (O_1750,N_14710,N_14858);
or UO_1751 (O_1751,N_14772,N_14912);
xor UO_1752 (O_1752,N_14839,N_14807);
and UO_1753 (O_1753,N_14721,N_14901);
or UO_1754 (O_1754,N_14705,N_14953);
nor UO_1755 (O_1755,N_14723,N_14857);
or UO_1756 (O_1756,N_14712,N_14827);
nand UO_1757 (O_1757,N_14789,N_14780);
nor UO_1758 (O_1758,N_14874,N_14927);
or UO_1759 (O_1759,N_14871,N_14768);
nand UO_1760 (O_1760,N_14830,N_14932);
nor UO_1761 (O_1761,N_14858,N_14776);
xor UO_1762 (O_1762,N_14711,N_14870);
xor UO_1763 (O_1763,N_14768,N_14879);
nor UO_1764 (O_1764,N_14824,N_14755);
nand UO_1765 (O_1765,N_14749,N_14965);
nand UO_1766 (O_1766,N_14715,N_14928);
xor UO_1767 (O_1767,N_14791,N_14859);
xor UO_1768 (O_1768,N_14723,N_14940);
and UO_1769 (O_1769,N_14973,N_14822);
nand UO_1770 (O_1770,N_14863,N_14736);
and UO_1771 (O_1771,N_14909,N_14917);
xnor UO_1772 (O_1772,N_14988,N_14762);
xor UO_1773 (O_1773,N_14775,N_14716);
or UO_1774 (O_1774,N_14826,N_14898);
nand UO_1775 (O_1775,N_14855,N_14748);
nand UO_1776 (O_1776,N_14943,N_14764);
and UO_1777 (O_1777,N_14824,N_14892);
or UO_1778 (O_1778,N_14825,N_14873);
and UO_1779 (O_1779,N_14987,N_14930);
xnor UO_1780 (O_1780,N_14837,N_14733);
or UO_1781 (O_1781,N_14812,N_14806);
nor UO_1782 (O_1782,N_14802,N_14754);
or UO_1783 (O_1783,N_14731,N_14745);
nor UO_1784 (O_1784,N_14986,N_14906);
nand UO_1785 (O_1785,N_14981,N_14746);
or UO_1786 (O_1786,N_14782,N_14814);
xor UO_1787 (O_1787,N_14816,N_14975);
nor UO_1788 (O_1788,N_14813,N_14752);
xnor UO_1789 (O_1789,N_14966,N_14813);
and UO_1790 (O_1790,N_14782,N_14712);
xnor UO_1791 (O_1791,N_14977,N_14721);
nor UO_1792 (O_1792,N_14901,N_14789);
or UO_1793 (O_1793,N_14908,N_14859);
and UO_1794 (O_1794,N_14713,N_14933);
and UO_1795 (O_1795,N_14995,N_14877);
or UO_1796 (O_1796,N_14871,N_14824);
nand UO_1797 (O_1797,N_14968,N_14945);
and UO_1798 (O_1798,N_14849,N_14800);
nor UO_1799 (O_1799,N_14902,N_14861);
and UO_1800 (O_1800,N_14813,N_14852);
nand UO_1801 (O_1801,N_14915,N_14910);
xor UO_1802 (O_1802,N_14910,N_14730);
and UO_1803 (O_1803,N_14760,N_14879);
nand UO_1804 (O_1804,N_14846,N_14896);
nor UO_1805 (O_1805,N_14793,N_14948);
nor UO_1806 (O_1806,N_14941,N_14923);
nand UO_1807 (O_1807,N_14981,N_14725);
or UO_1808 (O_1808,N_14713,N_14989);
xor UO_1809 (O_1809,N_14799,N_14849);
or UO_1810 (O_1810,N_14926,N_14960);
and UO_1811 (O_1811,N_14926,N_14915);
nor UO_1812 (O_1812,N_14791,N_14756);
nor UO_1813 (O_1813,N_14832,N_14780);
nand UO_1814 (O_1814,N_14771,N_14741);
nand UO_1815 (O_1815,N_14705,N_14849);
nand UO_1816 (O_1816,N_14721,N_14951);
xor UO_1817 (O_1817,N_14974,N_14881);
or UO_1818 (O_1818,N_14930,N_14889);
xnor UO_1819 (O_1819,N_14990,N_14886);
nor UO_1820 (O_1820,N_14999,N_14954);
or UO_1821 (O_1821,N_14875,N_14935);
and UO_1822 (O_1822,N_14846,N_14919);
nor UO_1823 (O_1823,N_14871,N_14918);
nor UO_1824 (O_1824,N_14846,N_14907);
nand UO_1825 (O_1825,N_14868,N_14919);
xor UO_1826 (O_1826,N_14973,N_14920);
nor UO_1827 (O_1827,N_14978,N_14990);
nand UO_1828 (O_1828,N_14740,N_14980);
or UO_1829 (O_1829,N_14712,N_14918);
nand UO_1830 (O_1830,N_14781,N_14911);
and UO_1831 (O_1831,N_14717,N_14800);
or UO_1832 (O_1832,N_14874,N_14946);
nor UO_1833 (O_1833,N_14841,N_14951);
nand UO_1834 (O_1834,N_14897,N_14731);
nor UO_1835 (O_1835,N_14715,N_14883);
and UO_1836 (O_1836,N_14976,N_14973);
xor UO_1837 (O_1837,N_14744,N_14954);
nor UO_1838 (O_1838,N_14784,N_14770);
and UO_1839 (O_1839,N_14937,N_14865);
nor UO_1840 (O_1840,N_14900,N_14888);
and UO_1841 (O_1841,N_14946,N_14709);
nand UO_1842 (O_1842,N_14929,N_14795);
xor UO_1843 (O_1843,N_14871,N_14818);
or UO_1844 (O_1844,N_14908,N_14756);
or UO_1845 (O_1845,N_14719,N_14850);
nand UO_1846 (O_1846,N_14963,N_14766);
nand UO_1847 (O_1847,N_14906,N_14729);
nor UO_1848 (O_1848,N_14996,N_14796);
nand UO_1849 (O_1849,N_14940,N_14781);
nor UO_1850 (O_1850,N_14753,N_14929);
nor UO_1851 (O_1851,N_14959,N_14789);
nor UO_1852 (O_1852,N_14759,N_14878);
nand UO_1853 (O_1853,N_14868,N_14990);
nand UO_1854 (O_1854,N_14890,N_14846);
nand UO_1855 (O_1855,N_14713,N_14873);
and UO_1856 (O_1856,N_14728,N_14710);
and UO_1857 (O_1857,N_14813,N_14732);
or UO_1858 (O_1858,N_14743,N_14979);
nor UO_1859 (O_1859,N_14947,N_14749);
xor UO_1860 (O_1860,N_14797,N_14773);
nor UO_1861 (O_1861,N_14987,N_14902);
and UO_1862 (O_1862,N_14821,N_14810);
nand UO_1863 (O_1863,N_14801,N_14731);
and UO_1864 (O_1864,N_14702,N_14717);
nor UO_1865 (O_1865,N_14776,N_14922);
or UO_1866 (O_1866,N_14852,N_14706);
or UO_1867 (O_1867,N_14961,N_14778);
nor UO_1868 (O_1868,N_14788,N_14907);
and UO_1869 (O_1869,N_14719,N_14791);
nor UO_1870 (O_1870,N_14929,N_14888);
nand UO_1871 (O_1871,N_14913,N_14855);
nand UO_1872 (O_1872,N_14720,N_14761);
nor UO_1873 (O_1873,N_14701,N_14762);
or UO_1874 (O_1874,N_14740,N_14954);
nor UO_1875 (O_1875,N_14749,N_14724);
or UO_1876 (O_1876,N_14868,N_14774);
xor UO_1877 (O_1877,N_14963,N_14834);
nand UO_1878 (O_1878,N_14737,N_14995);
nand UO_1879 (O_1879,N_14968,N_14905);
and UO_1880 (O_1880,N_14885,N_14987);
or UO_1881 (O_1881,N_14999,N_14875);
and UO_1882 (O_1882,N_14933,N_14720);
xnor UO_1883 (O_1883,N_14977,N_14787);
nor UO_1884 (O_1884,N_14788,N_14757);
nand UO_1885 (O_1885,N_14722,N_14877);
nand UO_1886 (O_1886,N_14764,N_14840);
and UO_1887 (O_1887,N_14735,N_14973);
nor UO_1888 (O_1888,N_14823,N_14769);
nand UO_1889 (O_1889,N_14763,N_14705);
nor UO_1890 (O_1890,N_14977,N_14754);
or UO_1891 (O_1891,N_14912,N_14958);
nor UO_1892 (O_1892,N_14728,N_14833);
nor UO_1893 (O_1893,N_14777,N_14837);
xor UO_1894 (O_1894,N_14938,N_14705);
nand UO_1895 (O_1895,N_14876,N_14826);
and UO_1896 (O_1896,N_14953,N_14804);
or UO_1897 (O_1897,N_14897,N_14744);
and UO_1898 (O_1898,N_14812,N_14832);
and UO_1899 (O_1899,N_14750,N_14741);
nand UO_1900 (O_1900,N_14956,N_14975);
nand UO_1901 (O_1901,N_14770,N_14873);
nand UO_1902 (O_1902,N_14759,N_14771);
or UO_1903 (O_1903,N_14798,N_14719);
xnor UO_1904 (O_1904,N_14801,N_14719);
xor UO_1905 (O_1905,N_14723,N_14904);
and UO_1906 (O_1906,N_14767,N_14836);
and UO_1907 (O_1907,N_14813,N_14833);
nand UO_1908 (O_1908,N_14885,N_14853);
nor UO_1909 (O_1909,N_14705,N_14822);
nor UO_1910 (O_1910,N_14840,N_14773);
or UO_1911 (O_1911,N_14907,N_14830);
xnor UO_1912 (O_1912,N_14808,N_14868);
nor UO_1913 (O_1913,N_14924,N_14704);
nor UO_1914 (O_1914,N_14712,N_14747);
nand UO_1915 (O_1915,N_14934,N_14744);
nand UO_1916 (O_1916,N_14841,N_14703);
and UO_1917 (O_1917,N_14966,N_14952);
or UO_1918 (O_1918,N_14733,N_14824);
nand UO_1919 (O_1919,N_14804,N_14915);
xor UO_1920 (O_1920,N_14803,N_14724);
xor UO_1921 (O_1921,N_14778,N_14787);
nor UO_1922 (O_1922,N_14781,N_14707);
nor UO_1923 (O_1923,N_14844,N_14969);
nand UO_1924 (O_1924,N_14965,N_14955);
xor UO_1925 (O_1925,N_14872,N_14748);
or UO_1926 (O_1926,N_14753,N_14722);
or UO_1927 (O_1927,N_14811,N_14905);
nand UO_1928 (O_1928,N_14719,N_14884);
and UO_1929 (O_1929,N_14843,N_14874);
nor UO_1930 (O_1930,N_14875,N_14979);
and UO_1931 (O_1931,N_14899,N_14712);
or UO_1932 (O_1932,N_14730,N_14838);
nand UO_1933 (O_1933,N_14857,N_14761);
nand UO_1934 (O_1934,N_14970,N_14857);
nand UO_1935 (O_1935,N_14852,N_14795);
nand UO_1936 (O_1936,N_14850,N_14838);
nor UO_1937 (O_1937,N_14710,N_14993);
nor UO_1938 (O_1938,N_14836,N_14987);
and UO_1939 (O_1939,N_14973,N_14743);
xnor UO_1940 (O_1940,N_14876,N_14961);
or UO_1941 (O_1941,N_14766,N_14939);
xnor UO_1942 (O_1942,N_14994,N_14816);
nand UO_1943 (O_1943,N_14966,N_14978);
nor UO_1944 (O_1944,N_14800,N_14949);
nor UO_1945 (O_1945,N_14862,N_14935);
or UO_1946 (O_1946,N_14928,N_14900);
nand UO_1947 (O_1947,N_14786,N_14899);
xor UO_1948 (O_1948,N_14824,N_14863);
and UO_1949 (O_1949,N_14988,N_14992);
xor UO_1950 (O_1950,N_14999,N_14944);
nand UO_1951 (O_1951,N_14772,N_14824);
or UO_1952 (O_1952,N_14996,N_14961);
nand UO_1953 (O_1953,N_14755,N_14828);
or UO_1954 (O_1954,N_14756,N_14821);
and UO_1955 (O_1955,N_14728,N_14876);
nor UO_1956 (O_1956,N_14761,N_14846);
and UO_1957 (O_1957,N_14705,N_14881);
or UO_1958 (O_1958,N_14891,N_14939);
nand UO_1959 (O_1959,N_14820,N_14980);
xnor UO_1960 (O_1960,N_14744,N_14828);
nor UO_1961 (O_1961,N_14838,N_14911);
nand UO_1962 (O_1962,N_14946,N_14784);
xor UO_1963 (O_1963,N_14743,N_14912);
xor UO_1964 (O_1964,N_14821,N_14912);
and UO_1965 (O_1965,N_14704,N_14994);
and UO_1966 (O_1966,N_14701,N_14731);
nor UO_1967 (O_1967,N_14778,N_14772);
nor UO_1968 (O_1968,N_14937,N_14947);
or UO_1969 (O_1969,N_14940,N_14923);
nand UO_1970 (O_1970,N_14827,N_14839);
or UO_1971 (O_1971,N_14948,N_14840);
and UO_1972 (O_1972,N_14964,N_14949);
or UO_1973 (O_1973,N_14849,N_14809);
nand UO_1974 (O_1974,N_14950,N_14857);
xor UO_1975 (O_1975,N_14814,N_14711);
or UO_1976 (O_1976,N_14735,N_14785);
and UO_1977 (O_1977,N_14980,N_14936);
nand UO_1978 (O_1978,N_14808,N_14733);
nor UO_1979 (O_1979,N_14705,N_14930);
xnor UO_1980 (O_1980,N_14708,N_14882);
and UO_1981 (O_1981,N_14915,N_14976);
or UO_1982 (O_1982,N_14800,N_14719);
xor UO_1983 (O_1983,N_14701,N_14802);
and UO_1984 (O_1984,N_14819,N_14860);
and UO_1985 (O_1985,N_14720,N_14966);
nor UO_1986 (O_1986,N_14722,N_14737);
xor UO_1987 (O_1987,N_14733,N_14887);
nor UO_1988 (O_1988,N_14756,N_14738);
nor UO_1989 (O_1989,N_14957,N_14917);
or UO_1990 (O_1990,N_14829,N_14737);
nand UO_1991 (O_1991,N_14982,N_14737);
xnor UO_1992 (O_1992,N_14734,N_14921);
or UO_1993 (O_1993,N_14754,N_14803);
or UO_1994 (O_1994,N_14950,N_14704);
nor UO_1995 (O_1995,N_14714,N_14801);
or UO_1996 (O_1996,N_14953,N_14964);
or UO_1997 (O_1997,N_14790,N_14919);
or UO_1998 (O_1998,N_14755,N_14795);
or UO_1999 (O_1999,N_14736,N_14984);
endmodule