module basic_1500_15000_2000_75_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
or U0 (N_0,In_438,In_316);
and U1 (N_1,In_1260,In_362);
and U2 (N_2,In_1232,In_586);
or U3 (N_3,In_5,In_75);
xnor U4 (N_4,In_1440,In_1115);
xnor U5 (N_5,In_201,In_498);
nand U6 (N_6,In_703,In_499);
and U7 (N_7,In_734,In_579);
xor U8 (N_8,In_1255,In_95);
and U9 (N_9,In_941,In_690);
nor U10 (N_10,In_994,In_618);
xnor U11 (N_11,In_607,In_574);
nand U12 (N_12,In_1394,In_418);
and U13 (N_13,In_1299,In_205);
nand U14 (N_14,In_1414,In_785);
nand U15 (N_15,In_1141,In_47);
nor U16 (N_16,In_374,In_376);
or U17 (N_17,In_515,In_942);
xor U18 (N_18,In_635,In_107);
nor U19 (N_19,In_1402,In_987);
or U20 (N_20,In_236,In_210);
or U21 (N_21,In_344,In_889);
and U22 (N_22,In_1179,In_332);
xnor U23 (N_23,In_1137,In_1286);
nor U24 (N_24,In_222,In_128);
xnor U25 (N_25,In_164,In_805);
or U26 (N_26,In_440,In_280);
or U27 (N_27,In_291,In_373);
nor U28 (N_28,In_1272,In_117);
xor U29 (N_29,In_0,In_427);
nand U30 (N_30,In_435,In_1046);
and U31 (N_31,In_253,In_1093);
or U32 (N_32,In_434,In_166);
xor U33 (N_33,In_764,In_788);
nand U34 (N_34,In_1020,In_691);
nor U35 (N_35,In_350,In_390);
or U36 (N_36,In_273,In_394);
and U37 (N_37,In_35,In_247);
xnor U38 (N_38,In_591,In_363);
xor U39 (N_39,In_81,In_1122);
xnor U40 (N_40,In_552,In_188);
nand U41 (N_41,In_1083,In_17);
nand U42 (N_42,In_127,In_932);
nor U43 (N_43,In_719,In_365);
and U44 (N_44,In_306,In_246);
xnor U45 (N_45,In_423,In_198);
nor U46 (N_46,In_1395,In_525);
nand U47 (N_47,In_1054,In_1373);
or U48 (N_48,In_554,In_1472);
nand U49 (N_49,In_1019,In_87);
or U50 (N_50,In_313,In_1322);
nor U51 (N_51,In_450,In_1326);
and U52 (N_52,In_962,In_257);
and U53 (N_53,In_1123,In_1024);
nand U54 (N_54,In_1492,In_929);
nor U55 (N_55,In_1366,In_80);
xnor U56 (N_56,In_519,In_832);
or U57 (N_57,In_20,In_1092);
nand U58 (N_58,In_1391,In_272);
nor U59 (N_59,In_359,In_1289);
nand U60 (N_60,In_97,In_1204);
nand U61 (N_61,In_1172,In_720);
nand U62 (N_62,In_142,In_102);
or U63 (N_63,In_592,In_820);
and U64 (N_64,In_567,In_1098);
nor U65 (N_65,In_1025,In_1089);
nand U66 (N_66,In_840,In_1283);
xnor U67 (N_67,In_1355,In_689);
or U68 (N_68,In_138,In_855);
nor U69 (N_69,In_202,In_736);
xnor U70 (N_70,In_837,In_896);
xnor U71 (N_71,In_1426,In_1072);
and U72 (N_72,In_1169,In_41);
xnor U73 (N_73,In_1429,In_1433);
nand U74 (N_74,In_318,In_693);
nor U75 (N_75,In_366,In_1453);
xor U76 (N_76,In_333,In_955);
nor U77 (N_77,In_401,In_296);
xnor U78 (N_78,In_162,In_66);
or U79 (N_79,In_1337,In_336);
or U80 (N_80,In_869,In_251);
or U81 (N_81,In_214,In_626);
nand U82 (N_82,In_326,In_865);
nor U83 (N_83,In_405,In_1369);
nand U84 (N_84,In_1487,In_1220);
nand U85 (N_85,In_106,In_1155);
or U86 (N_86,In_1086,In_449);
xor U87 (N_87,In_90,In_346);
or U88 (N_88,In_239,In_371);
nand U89 (N_89,In_1475,In_426);
or U90 (N_90,In_8,In_1251);
and U91 (N_91,In_1409,In_483);
and U92 (N_92,In_713,In_1221);
and U93 (N_93,In_1482,In_425);
and U94 (N_94,In_460,In_914);
xnor U95 (N_95,In_605,In_375);
and U96 (N_96,In_1403,In_1005);
and U97 (N_97,In_311,In_1125);
and U98 (N_98,In_1007,In_46);
xor U99 (N_99,In_705,In_553);
and U100 (N_100,In_388,In_1009);
xnor U101 (N_101,In_77,In_1269);
xor U102 (N_102,In_1063,In_584);
nand U103 (N_103,In_857,In_185);
nand U104 (N_104,In_1461,In_403);
or U105 (N_105,In_503,In_1143);
nand U106 (N_106,In_868,In_1419);
xor U107 (N_107,In_1154,In_152);
or U108 (N_108,In_282,In_98);
nand U109 (N_109,In_549,In_953);
and U110 (N_110,In_276,In_1401);
nand U111 (N_111,In_1457,In_1361);
or U112 (N_112,In_1231,In_601);
and U113 (N_113,In_1151,In_585);
nor U114 (N_114,In_355,In_886);
xnor U115 (N_115,In_864,In_771);
and U116 (N_116,In_817,In_1273);
or U117 (N_117,In_786,In_1420);
and U118 (N_118,In_168,In_977);
nand U119 (N_119,In_1104,In_140);
nor U120 (N_120,In_1474,In_1271);
nor U121 (N_121,In_1160,In_1217);
nand U122 (N_122,In_685,In_244);
nand U123 (N_123,In_923,In_1287);
or U124 (N_124,In_169,In_1132);
or U125 (N_125,In_768,In_576);
xnor U126 (N_126,In_458,In_1319);
and U127 (N_127,In_1079,In_1118);
and U128 (N_128,In_975,In_821);
or U129 (N_129,In_416,In_876);
or U130 (N_130,In_338,In_1171);
nand U131 (N_131,In_668,In_847);
xor U132 (N_132,In_613,In_1168);
or U133 (N_133,In_878,In_1034);
and U134 (N_134,In_1205,In_1434);
and U135 (N_135,In_965,In_904);
nand U136 (N_136,In_1467,In_660);
and U137 (N_137,In_286,In_721);
xnor U138 (N_138,In_184,In_1292);
or U139 (N_139,In_589,In_407);
nand U140 (N_140,In_297,In_1058);
nand U141 (N_141,In_262,In_396);
nand U142 (N_142,In_1274,In_836);
and U143 (N_143,In_1002,In_212);
nor U144 (N_144,In_1078,In_803);
or U145 (N_145,In_1237,In_1211);
xnor U146 (N_146,In_310,In_113);
xor U147 (N_147,In_640,In_321);
nand U148 (N_148,In_320,In_594);
or U149 (N_149,In_85,In_841);
and U150 (N_150,In_1384,In_735);
xnor U151 (N_151,In_1053,In_1101);
nand U152 (N_152,In_756,In_849);
xnor U153 (N_153,In_543,In_322);
nor U154 (N_154,In_369,In_793);
nand U155 (N_155,In_1186,In_759);
or U156 (N_156,In_370,In_686);
xnor U157 (N_157,In_1064,In_1246);
or U158 (N_158,In_1037,In_187);
or U159 (N_159,In_1317,In_459);
or U160 (N_160,In_1379,In_232);
nor U161 (N_161,In_752,In_599);
or U162 (N_162,In_1250,In_615);
nor U163 (N_163,In_1153,In_389);
and U164 (N_164,In_422,In_64);
xor U165 (N_165,In_380,In_1052);
nor U166 (N_166,In_824,In_708);
and U167 (N_167,In_319,In_497);
or U168 (N_168,In_529,In_298);
nor U169 (N_169,In_704,In_650);
or U170 (N_170,In_1008,In_1175);
and U171 (N_171,In_1439,In_789);
and U172 (N_172,In_219,In_192);
nand U173 (N_173,In_1157,In_1334);
or U174 (N_174,In_546,In_1328);
and U175 (N_175,In_744,In_980);
xor U176 (N_176,In_897,In_415);
nor U177 (N_177,In_1012,In_653);
nand U178 (N_178,In_1233,In_1187);
nand U179 (N_179,In_1464,In_639);
and U180 (N_180,In_315,In_491);
nand U181 (N_181,In_421,In_466);
nand U182 (N_182,In_564,In_538);
nand U183 (N_183,In_1185,In_749);
xor U184 (N_184,In_1183,In_11);
nand U185 (N_185,In_37,In_385);
and U186 (N_186,In_178,In_773);
and U187 (N_187,In_14,In_1026);
and U188 (N_188,In_505,In_702);
nor U189 (N_189,In_1349,In_1312);
xnor U190 (N_190,In_1127,In_1057);
xnor U191 (N_191,In_995,In_946);
nand U192 (N_192,In_270,In_745);
nor U193 (N_193,In_1015,In_1470);
and U194 (N_194,In_3,In_1138);
xnor U195 (N_195,In_255,In_597);
xnor U196 (N_196,In_175,In_135);
xor U197 (N_197,In_149,In_1193);
and U198 (N_198,In_1229,In_216);
or U199 (N_199,In_1463,In_217);
xor U200 (N_200,In_1252,In_70);
nor U201 (N_201,In_487,N_71);
and U202 (N_202,In_905,In_517);
or U203 (N_203,In_948,In_806);
nand U204 (N_204,In_807,In_1288);
nand U205 (N_205,In_748,In_1399);
or U206 (N_206,In_741,In_259);
and U207 (N_207,In_1228,In_112);
nor U208 (N_208,In_1449,In_508);
nor U209 (N_209,In_1082,In_227);
xnor U210 (N_210,In_609,In_765);
nand U211 (N_211,In_1333,In_82);
nand U212 (N_212,In_659,In_1392);
nand U213 (N_213,In_1061,In_1077);
xnor U214 (N_214,In_1131,N_68);
nor U215 (N_215,N_20,In_1297);
nor U216 (N_216,In_1416,In_174);
xor U217 (N_217,In_455,In_21);
and U218 (N_218,In_1385,In_2);
or U219 (N_219,In_62,In_1368);
xnor U220 (N_220,In_384,In_195);
and U221 (N_221,In_500,In_943);
nand U222 (N_222,In_409,In_226);
nor U223 (N_223,In_1084,In_299);
nand U224 (N_224,In_610,In_1133);
nand U225 (N_225,In_924,N_120);
and U226 (N_226,In_1048,N_148);
or U227 (N_227,In_1206,In_544);
nand U228 (N_228,In_746,In_608);
or U229 (N_229,In_1378,In_1107);
nor U230 (N_230,In_358,In_263);
and U231 (N_231,In_1109,N_58);
xor U232 (N_232,N_50,In_769);
nand U233 (N_233,In_939,In_731);
and U234 (N_234,In_619,N_155);
and U235 (N_235,In_133,N_116);
or U236 (N_236,In_930,In_875);
or U237 (N_237,In_859,In_898);
nor U238 (N_238,In_1216,In_1055);
or U239 (N_239,In_1190,In_92);
and U240 (N_240,In_1215,In_51);
or U241 (N_241,In_1170,In_1050);
xnor U242 (N_242,N_43,N_196);
and U243 (N_243,In_1374,In_479);
or U244 (N_244,In_883,In_658);
or U245 (N_245,In_1192,N_180);
nand U246 (N_246,In_1425,In_716);
xnor U247 (N_247,In_1313,In_628);
nor U248 (N_248,In_30,In_688);
nor U249 (N_249,In_536,In_947);
and U250 (N_250,In_674,In_634);
nor U251 (N_251,In_1184,N_4);
nand U252 (N_252,In_155,In_377);
nand U253 (N_253,In_1371,N_94);
nand U254 (N_254,In_1448,In_274);
xnor U255 (N_255,N_49,In_234);
nor U256 (N_256,In_451,In_19);
or U257 (N_257,N_144,In_1111);
nand U258 (N_258,In_952,In_652);
or U259 (N_259,In_115,In_367);
nand U260 (N_260,N_42,In_1365);
nor U261 (N_261,In_854,N_56);
nor U262 (N_262,N_8,N_12);
nor U263 (N_263,In_1478,In_442);
nand U264 (N_264,In_317,N_166);
xnor U265 (N_265,In_625,In_915);
nand U266 (N_266,N_5,In_208);
nand U267 (N_267,In_1267,In_603);
or U268 (N_268,In_6,In_911);
nor U269 (N_269,In_1235,In_888);
nor U270 (N_270,In_1212,In_1496);
and U271 (N_271,In_1338,In_870);
and U272 (N_272,In_679,In_271);
xnor U273 (N_273,In_29,N_102);
xor U274 (N_274,In_410,In_1364);
or U275 (N_275,In_1330,In_356);
nand U276 (N_276,In_815,In_1066);
nor U277 (N_277,In_26,In_488);
nor U278 (N_278,N_55,In_1033);
or U279 (N_279,N_146,In_55);
nand U280 (N_280,N_177,In_1120);
and U281 (N_281,In_1280,In_96);
nand U282 (N_282,In_638,In_750);
and U283 (N_283,In_763,In_902);
xnor U284 (N_284,In_1129,In_325);
xor U285 (N_285,In_1346,In_722);
and U286 (N_286,In_349,In_557);
or U287 (N_287,In_710,In_173);
and U288 (N_288,N_197,In_916);
or U289 (N_289,N_17,In_891);
nand U290 (N_290,In_1126,In_541);
xnor U291 (N_291,In_606,In_533);
nor U292 (N_292,N_39,In_324);
and U293 (N_293,In_862,In_481);
and U294 (N_294,In_880,In_1180);
xnor U295 (N_295,In_1265,In_478);
xnor U296 (N_296,In_830,In_1119);
xor U297 (N_297,In_661,In_1097);
and U298 (N_298,N_93,In_191);
xnor U299 (N_299,In_1114,In_1488);
nor U300 (N_300,In_470,N_7);
or U301 (N_301,In_1076,N_41);
xnor U302 (N_302,N_98,In_24);
xnor U303 (N_303,N_76,N_89);
nor U304 (N_304,In_159,N_170);
nand U305 (N_305,In_738,In_1441);
or U306 (N_306,In_1166,In_707);
and U307 (N_307,In_1124,In_678);
nor U308 (N_308,N_48,In_16);
xor U309 (N_309,In_334,In_118);
nand U310 (N_310,N_194,In_1261);
and U311 (N_311,N_80,In_328);
xnor U312 (N_312,In_1159,In_335);
or U313 (N_313,In_476,In_669);
nor U314 (N_314,In_1428,In_726);
or U315 (N_315,In_1422,In_204);
nor U316 (N_316,In_443,In_853);
nand U317 (N_317,In_1094,In_1435);
nor U318 (N_318,In_284,In_562);
nand U319 (N_319,In_211,In_1090);
or U320 (N_320,In_866,In_521);
and U321 (N_321,In_758,In_144);
nand U322 (N_322,N_183,In_268);
and U323 (N_323,N_141,In_622);
nor U324 (N_324,In_1240,In_261);
or U325 (N_325,N_96,In_663);
and U326 (N_326,In_1222,In_908);
nand U327 (N_327,In_1342,In_91);
or U328 (N_328,In_1156,In_148);
xor U329 (N_329,N_103,In_397);
or U330 (N_330,In_797,In_844);
xor U331 (N_331,In_1423,In_522);
or U332 (N_332,In_68,In_467);
nor U333 (N_333,In_922,In_860);
and U334 (N_334,In_134,N_165);
xor U335 (N_335,N_59,In_1412);
xor U336 (N_336,In_330,In_83);
nor U337 (N_337,In_737,In_1320);
nor U338 (N_338,In_1214,In_918);
nor U339 (N_339,In_570,In_1437);
nor U340 (N_340,In_651,In_25);
or U341 (N_341,In_1305,In_1162);
xor U342 (N_342,In_931,In_54);
or U343 (N_343,In_770,In_780);
nand U344 (N_344,In_809,In_811);
and U345 (N_345,In_648,In_1341);
nand U346 (N_346,In_309,In_1087);
nor U347 (N_347,In_1471,In_1016);
xnor U348 (N_348,In_151,In_383);
and U349 (N_349,In_248,In_666);
xnor U350 (N_350,In_833,In_725);
xor U351 (N_351,In_125,In_43);
or U352 (N_352,In_611,In_819);
and U353 (N_353,In_1158,In_1011);
nor U354 (N_354,In_551,In_733);
or U355 (N_355,In_754,In_534);
and U356 (N_356,N_174,In_141);
nand U357 (N_357,N_34,In_13);
and U358 (N_358,In_368,In_361);
or U359 (N_359,In_468,In_910);
nand U360 (N_360,N_162,N_97);
nor U361 (N_361,N_178,In_555);
nand U362 (N_362,In_258,In_1308);
nor U363 (N_363,In_1195,N_9);
xor U364 (N_364,In_1296,N_95);
or U365 (N_365,In_612,In_917);
nor U366 (N_366,N_14,In_988);
xor U367 (N_367,In_379,In_1410);
or U368 (N_368,In_1121,N_187);
or U369 (N_369,N_11,In_1070);
xnor U370 (N_370,In_921,In_774);
xor U371 (N_371,In_233,In_732);
nor U372 (N_372,In_391,In_1480);
nor U373 (N_373,In_681,In_1146);
nor U374 (N_374,In_493,N_193);
and U375 (N_375,In_1389,N_2);
nand U376 (N_376,In_22,In_954);
nand U377 (N_377,In_156,In_93);
and U378 (N_378,In_108,In_1248);
xnor U379 (N_379,In_1081,In_777);
or U380 (N_380,N_176,In_684);
nor U381 (N_381,In_457,In_49);
nand U382 (N_382,In_945,In_935);
nand U383 (N_383,In_1262,In_1350);
or U384 (N_384,In_1051,In_1181);
xor U385 (N_385,In_1238,In_671);
and U386 (N_386,In_1257,In_267);
or U387 (N_387,N_53,In_150);
and U388 (N_388,In_839,N_70);
xnor U389 (N_389,In_285,In_1022);
or U390 (N_390,In_620,In_1259);
nor U391 (N_391,N_110,In_327);
and U392 (N_392,In_343,N_108);
xor U393 (N_393,In_672,In_506);
and U394 (N_394,In_110,In_348);
nor U395 (N_395,In_456,In_1256);
and U396 (N_396,In_27,In_1310);
nand U397 (N_397,In_834,In_1438);
and U398 (N_398,In_912,N_161);
nor U399 (N_399,In_602,N_54);
nor U400 (N_400,In_67,N_221);
xor U401 (N_401,In_337,In_1149);
nand U402 (N_402,In_596,In_360);
or U403 (N_403,In_957,In_277);
xor U404 (N_404,In_254,In_480);
or U405 (N_405,In_163,In_527);
or U406 (N_406,In_630,In_999);
nor U407 (N_407,N_30,N_241);
xnor U408 (N_408,In_1208,In_964);
nand U409 (N_409,In_59,In_221);
and U410 (N_410,N_217,In_1460);
nand U411 (N_411,In_959,N_318);
and U412 (N_412,In_877,N_184);
or U413 (N_413,N_270,In_119);
and U414 (N_414,In_1469,In_632);
or U415 (N_415,N_206,In_161);
or U416 (N_416,N_395,In_1466);
nand U417 (N_417,N_278,N_245);
nand U418 (N_418,In_243,In_495);
nor U419 (N_419,In_1413,In_469);
xnor U420 (N_420,N_330,In_548);
or U421 (N_421,In_1188,In_984);
or U422 (N_422,In_1110,In_772);
or U423 (N_423,In_484,In_1404);
or U424 (N_424,N_247,N_173);
xor U425 (N_425,In_1230,In_727);
nor U426 (N_426,In_1130,N_224);
xor U427 (N_427,In_431,In_1021);
nand U428 (N_428,In_940,In_1135);
xnor U429 (N_429,In_1103,N_205);
nand U430 (N_430,In_676,N_310);
and U431 (N_431,In_1315,N_192);
nor U432 (N_432,N_126,In_1088);
xnor U433 (N_433,In_1477,In_44);
xnor U434 (N_434,N_243,In_667);
nand U435 (N_435,N_32,In_1234);
xnor U436 (N_436,In_1030,In_242);
and U437 (N_437,In_489,In_983);
or U438 (N_438,In_1400,In_237);
nor U439 (N_439,In_509,In_1145);
or U440 (N_440,In_1321,N_377);
xor U441 (N_441,N_311,N_175);
or U442 (N_442,N_301,N_363);
nand U443 (N_443,In_677,In_1300);
and U444 (N_444,In_176,N_152);
xnor U445 (N_445,In_714,In_1307);
nor U446 (N_446,In_697,N_27);
and U447 (N_447,N_19,In_743);
and U448 (N_448,In_200,N_239);
nor U449 (N_449,In_968,In_879);
or U450 (N_450,In_1035,In_1178);
xnor U451 (N_451,In_623,N_350);
or U452 (N_452,N_259,In_1249);
and U453 (N_453,N_373,In_1398);
and U454 (N_454,N_202,In_706);
and U455 (N_455,In_979,N_91);
or U456 (N_456,In_307,In_1291);
xor U457 (N_457,In_717,N_129);
xor U458 (N_458,In_882,N_65);
and U459 (N_459,N_254,In_991);
xor U460 (N_460,In_1163,N_37);
nor U461 (N_461,In_779,In_981);
nor U462 (N_462,In_129,In_531);
nand U463 (N_463,N_356,In_1468);
nor U464 (N_464,N_360,In_65);
and U465 (N_465,N_303,In_1290);
or U466 (N_466,In_1386,In_153);
xnor U467 (N_467,N_249,In_825);
or U468 (N_468,In_1309,In_1085);
xor U469 (N_469,In_206,In_776);
nand U470 (N_470,In_472,In_913);
xnor U471 (N_471,In_1031,In_516);
or U472 (N_472,N_60,In_1336);
nand U473 (N_473,In_1177,In_132);
and U474 (N_474,In_664,In_1325);
and U475 (N_475,In_196,N_199);
and U476 (N_476,N_28,In_1038);
nand U477 (N_477,In_966,N_160);
nand U478 (N_478,In_631,In_1279);
xnor U479 (N_479,In_1277,In_7);
nand U480 (N_480,In_890,N_284);
and U481 (N_481,In_747,N_38);
and U482 (N_482,N_13,In_1359);
xnor U483 (N_483,In_850,N_319);
and U484 (N_484,In_1303,N_219);
nand U485 (N_485,N_391,In_795);
nand U486 (N_486,In_39,N_328);
or U487 (N_487,In_512,N_313);
or U488 (N_488,In_130,In_718);
nand U489 (N_489,In_1362,N_172);
and U490 (N_490,In_290,In_1356);
or U491 (N_491,In_818,In_218);
and U492 (N_492,In_701,In_1323);
nor U493 (N_493,In_74,In_675);
and U494 (N_494,N_134,In_1406);
nand U495 (N_495,N_320,In_281);
nand U496 (N_496,In_960,N_114);
xnor U497 (N_497,In_465,In_813);
xnor U498 (N_498,N_396,N_132);
nor U499 (N_499,In_79,In_1003);
nor U500 (N_500,In_1000,In_1176);
or U501 (N_501,In_775,In_986);
and U502 (N_502,In_1043,In_1150);
xnor U503 (N_503,In_1294,In_871);
nor U504 (N_504,In_944,N_64);
nor U505 (N_505,N_85,N_45);
or U506 (N_506,In_812,In_1494);
or U507 (N_507,In_934,N_44);
nand U508 (N_508,In_1014,N_213);
nor U509 (N_509,In_289,N_375);
nand U510 (N_510,In_798,In_408);
nand U511 (N_511,In_696,In_1278);
or U512 (N_512,In_1452,N_229);
and U513 (N_513,N_268,In_545);
nor U514 (N_514,N_88,In_1479);
nand U515 (N_515,In_199,In_114);
and U516 (N_516,N_269,In_1293);
and U517 (N_517,In_56,In_997);
nand U518 (N_518,In_429,N_86);
and U519 (N_519,N_248,N_190);
xor U520 (N_520,In_9,In_528);
nand U521 (N_521,In_1128,In_477);
or U522 (N_522,In_1210,In_903);
nor U523 (N_523,In_167,In_189);
nor U524 (N_524,In_1202,N_264);
xnor U525 (N_525,N_81,In_492);
nand U526 (N_526,In_99,In_1096);
xnor U527 (N_527,In_1199,N_203);
and U528 (N_528,In_1484,In_462);
nand U529 (N_529,In_1284,In_105);
nor U530 (N_530,In_4,In_1226);
xnor U531 (N_531,In_1363,In_203);
nor U532 (N_532,In_18,N_35);
nor U533 (N_533,In_1454,In_969);
nand U534 (N_534,N_21,N_256);
nor U535 (N_535,N_378,N_337);
or U536 (N_536,In_973,In_392);
nand U537 (N_537,In_559,In_437);
or U538 (N_538,In_1390,In_52);
xor U539 (N_539,N_371,In_504);
or U540 (N_540,N_361,In_683);
xnor U541 (N_541,N_154,In_1224);
nor U542 (N_542,In_919,In_1071);
nor U543 (N_543,In_1213,N_274);
xor U544 (N_544,In_873,In_73);
xor U545 (N_545,In_874,In_295);
and U546 (N_546,In_220,In_294);
nand U547 (N_547,In_928,N_140);
and U548 (N_548,N_163,In_12);
nor U549 (N_549,In_419,In_1243);
xor U550 (N_550,In_532,In_347);
or U551 (N_551,N_220,N_299);
nor U552 (N_552,In_84,In_1142);
and U553 (N_553,N_40,In_40);
xor U554 (N_554,In_621,In_1462);
nand U555 (N_555,N_195,N_253);
nand U556 (N_556,N_390,In_1383);
xnor U557 (N_557,In_1450,In_1264);
nand U558 (N_558,In_1415,N_340);
nand U559 (N_559,N_362,In_1189);
xnor U560 (N_560,N_357,In_446);
or U561 (N_561,In_45,N_142);
nor U562 (N_562,In_1068,N_290);
nand U563 (N_563,N_232,In_1316);
xor U564 (N_564,In_266,In_646);
and U565 (N_565,N_341,In_474);
nand U566 (N_566,In_542,In_655);
xnor U567 (N_567,In_1045,In_513);
nand U568 (N_568,N_298,N_314);
nor U569 (N_569,N_342,In_1006);
nor U570 (N_570,In_1446,In_453);
xor U571 (N_571,In_1340,N_164);
xnor U572 (N_572,N_246,In_936);
xor U573 (N_573,N_389,In_1147);
xor U574 (N_574,In_473,In_302);
nand U575 (N_575,In_89,In_633);
nand U576 (N_576,In_1444,In_1332);
and U577 (N_577,In_1263,In_1282);
nor U578 (N_578,In_171,N_201);
and U579 (N_579,In_131,N_352);
nand U580 (N_580,N_22,In_101);
nand U581 (N_581,In_1004,In_814);
xor U582 (N_582,In_989,In_1497);
or U583 (N_583,N_119,In_1253);
and U584 (N_584,In_342,In_580);
nand U585 (N_585,N_325,In_1388);
or U586 (N_586,In_395,In_424);
or U587 (N_587,In_1165,N_212);
nor U588 (N_588,In_1295,N_250);
nor U589 (N_589,In_573,In_949);
nand U590 (N_590,In_828,N_275);
xnor U591 (N_591,N_112,In_364);
nor U592 (N_592,N_285,In_1351);
nor U593 (N_593,In_556,In_887);
nor U594 (N_594,In_804,N_78);
or U595 (N_595,N_185,In_933);
nand U596 (N_596,N_265,In_838);
or U597 (N_597,N_151,In_179);
nor U598 (N_598,N_107,In_1112);
nor U599 (N_599,In_1304,In_961);
and U600 (N_600,N_348,N_90);
or U601 (N_601,In_240,N_150);
or U602 (N_602,N_403,N_451);
nor U603 (N_603,N_15,N_331);
or U604 (N_604,In_1357,In_790);
xor U605 (N_605,N_226,In_139);
xor U606 (N_606,N_421,N_435);
nand U607 (N_607,In_1148,In_972);
nor U608 (N_608,In_800,N_560);
and U609 (N_609,In_1059,In_582);
and U610 (N_610,In_100,In_1370);
nand U611 (N_611,N_204,N_283);
nand U612 (N_612,N_564,In_588);
nor U613 (N_613,N_555,N_260);
nor U614 (N_614,In_436,N_503);
and U615 (N_615,In_637,In_402);
nand U616 (N_616,N_516,N_445);
nand U617 (N_617,N_149,In_1100);
xor U618 (N_618,N_476,N_10);
nor U619 (N_619,N_289,N_145);
xor U620 (N_620,In_794,N_211);
or U621 (N_621,In_1,N_137);
and U622 (N_622,N_511,N_433);
xnor U623 (N_623,N_501,In_441);
and U624 (N_624,In_452,In_1490);
nand U625 (N_625,In_822,N_167);
nand U626 (N_626,In_1314,In_146);
nand U627 (N_627,N_427,N_46);
xnor U628 (N_628,In_1161,In_147);
xnor U629 (N_629,N_47,In_345);
nor U630 (N_630,N_575,N_304);
nor U631 (N_631,In_843,In_967);
nor U632 (N_632,In_177,In_951);
and U633 (N_633,In_136,In_894);
and U634 (N_634,N_31,In_406);
nand U635 (N_635,N_135,In_1254);
nor U636 (N_636,N_534,In_293);
or U637 (N_637,In_892,In_124);
xnor U638 (N_638,In_767,N_424);
nand U639 (N_639,In_404,In_996);
and U640 (N_640,N_469,In_1302);
and U641 (N_641,In_523,N_561);
or U642 (N_642,In_575,In_1074);
nor U643 (N_643,N_494,N_251);
nand U644 (N_644,In_1029,In_414);
and U645 (N_645,In_137,In_1270);
or U646 (N_646,N_487,N_430);
nand U647 (N_647,In_762,N_491);
xnor U648 (N_648,N_453,N_321);
xnor U649 (N_649,In_595,In_292);
nor U650 (N_650,N_51,In_34);
or U651 (N_651,N_506,In_1476);
and U652 (N_652,N_481,N_309);
xnor U653 (N_653,N_349,N_411);
nand U654 (N_654,In_561,In_329);
or U655 (N_655,In_799,In_1044);
and U656 (N_656,N_413,In_1223);
and U657 (N_657,In_207,N_29);
xnor U658 (N_658,N_567,In_1027);
nor U659 (N_659,In_160,In_673);
or U660 (N_660,N_440,In_760);
xnor U661 (N_661,N_416,In_300);
nor U662 (N_662,N_235,In_1152);
nand U663 (N_663,In_884,In_539);
or U664 (N_664,N_329,N_588);
or U665 (N_665,In_982,In_715);
or U666 (N_666,In_560,In_907);
or U667 (N_667,In_695,N_18);
xor U668 (N_668,In_180,N_593);
nand U669 (N_669,N_380,N_225);
and U670 (N_670,In_126,In_1458);
nor U671 (N_671,N_286,In_1095);
xnor U672 (N_672,N_553,In_1348);
or U673 (N_673,N_74,In_157);
nor U674 (N_674,In_53,In_122);
and U675 (N_675,In_742,N_312);
nand U676 (N_676,In_1498,In_111);
and U677 (N_677,In_215,In_872);
and U678 (N_678,N_379,In_649);
xnor U679 (N_679,N_591,In_382);
and U680 (N_680,In_642,In_1001);
or U681 (N_681,N_552,N_595);
xor U682 (N_682,N_255,In_976);
or U683 (N_683,In_413,N_470);
nor U684 (N_684,N_536,In_471);
nor U685 (N_685,N_442,N_429);
xnor U686 (N_686,In_448,In_1173);
nor U687 (N_687,N_263,N_580);
or U688 (N_688,In_900,N_169);
or U689 (N_689,In_1358,N_336);
and U690 (N_690,N_62,In_558);
and U691 (N_691,N_530,N_288);
and U692 (N_692,N_147,N_61);
nor U693 (N_693,N_537,In_308);
nor U694 (N_694,In_998,N_252);
nor U695 (N_695,N_316,In_120);
nor U696 (N_696,In_121,In_1099);
nor U697 (N_697,In_566,In_1377);
nand U698 (N_698,In_1459,In_229);
nor U699 (N_699,In_1039,In_1069);
and U700 (N_700,N_410,In_856);
xnor U701 (N_701,In_1481,In_10);
xnor U702 (N_702,In_445,N_258);
xnor U703 (N_703,N_334,N_480);
nor U704 (N_704,In_183,In_1473);
and U705 (N_705,N_234,In_724);
nor U706 (N_706,N_139,N_338);
xor U707 (N_707,In_490,N_428);
nand U708 (N_708,N_381,In_835);
and U709 (N_709,In_1117,N_452);
xor U710 (N_710,In_461,In_1380);
xnor U711 (N_711,In_1405,N_446);
and U712 (N_712,N_408,N_437);
and U713 (N_713,N_109,N_188);
nor U714 (N_714,In_518,N_412);
and U715 (N_715,In_881,N_458);
nor U716 (N_716,In_1418,N_510);
nand U717 (N_717,In_104,N_492);
or U718 (N_718,N_490,In_616);
and U719 (N_719,In_1375,N_417);
and U720 (N_720,N_277,In_1047);
xor U721 (N_721,In_1198,N_448);
xnor U722 (N_722,N_460,In_303);
nand U723 (N_723,N_374,In_48);
and U724 (N_724,In_305,In_1443);
and U725 (N_725,N_209,N_138);
and U726 (N_726,N_597,N_556);
and U727 (N_727,In_71,N_63);
nand U728 (N_728,In_331,N_520);
xor U729 (N_729,N_351,In_1174);
nor U730 (N_730,N_181,In_194);
or U731 (N_731,N_6,N_401);
xor U732 (N_732,In_454,N_585);
or U733 (N_733,In_398,In_1483);
xor U734 (N_734,N_550,In_78);
xnor U735 (N_735,In_581,In_1360);
nand U736 (N_736,In_1430,In_399);
nor U737 (N_737,In_260,In_572);
or U738 (N_738,In_1106,N_528);
and U739 (N_739,N_127,N_223);
xor U740 (N_740,In_1318,N_354);
xor U741 (N_741,N_366,In_751);
or U742 (N_742,In_740,N_384);
xor U743 (N_743,N_157,N_542);
nand U744 (N_744,N_383,In_1065);
nand U745 (N_745,In_172,In_61);
or U746 (N_746,N_158,N_441);
or U747 (N_747,N_300,N_496);
and U748 (N_748,In_829,In_411);
nand U749 (N_749,In_1424,In_958);
or U750 (N_750,N_423,N_287);
and U751 (N_751,In_1331,N_572);
and U752 (N_752,N_153,In_1499);
nor U753 (N_753,In_1144,In_1219);
nand U754 (N_754,In_1080,N_406);
or U755 (N_755,N_121,In_502);
nor U756 (N_756,N_409,N_207);
and U757 (N_757,N_257,In_57);
nor U758 (N_758,N_482,N_508);
nor U759 (N_759,N_493,N_186);
xor U760 (N_760,N_333,N_529);
and U761 (N_761,N_358,In_831);
or U762 (N_762,N_397,In_31);
nor U763 (N_763,N_272,N_365);
and U764 (N_764,In_439,N_295);
nor U765 (N_765,In_1134,In_170);
nor U766 (N_766,N_540,N_323);
nand U767 (N_767,N_370,In_1067);
nand U768 (N_768,N_261,N_488);
nand U769 (N_769,In_1018,N_574);
nand U770 (N_770,In_617,N_473);
nor U771 (N_771,In_312,In_372);
and U772 (N_772,N_486,In_1102);
nor U773 (N_773,N_554,In_88);
nand U774 (N_774,N_198,In_692);
nand U775 (N_775,In_950,In_1455);
or U776 (N_776,In_1372,N_407);
or U777 (N_777,In_1311,In_723);
nand U778 (N_778,In_792,In_197);
and U779 (N_779,N_179,In_250);
nor U780 (N_780,In_158,N_118);
nand U781 (N_781,In_978,In_1049);
nand U782 (N_782,N_386,N_439);
and U783 (N_783,In_23,N_233);
nand U784 (N_784,In_937,In_901);
or U785 (N_785,In_1010,In_1073);
and U786 (N_786,N_502,N_522);
or U787 (N_787,In_287,In_547);
or U788 (N_788,N_507,N_394);
and U789 (N_789,N_77,In_846);
xnor U790 (N_790,N_570,N_236);
nor U791 (N_791,In_699,In_893);
nand U792 (N_792,In_1393,In_238);
and U793 (N_793,In_698,N_551);
or U794 (N_794,In_1167,N_297);
and U795 (N_795,In_909,In_1182);
or U796 (N_796,N_566,In_1247);
and U797 (N_797,In_1196,N_517);
or U798 (N_798,N_583,In_304);
nand U799 (N_799,In_823,N_519);
nand U800 (N_800,N_761,N_635);
nand U801 (N_801,In_378,N_462);
nand U802 (N_802,N_449,In_656);
and U803 (N_803,In_520,N_794);
and U804 (N_804,N_657,N_613);
and U805 (N_805,N_579,N_645);
or U806 (N_806,In_213,N_296);
nand U807 (N_807,N_783,N_438);
nor U808 (N_808,In_657,In_1427);
and U809 (N_809,N_231,In_209);
nand U810 (N_810,In_1266,In_801);
nand U811 (N_811,In_69,N_719);
nand U812 (N_812,In_645,In_654);
xor U813 (N_813,In_1091,In_109);
or U814 (N_814,N_663,N_326);
or U815 (N_815,N_587,In_895);
xnor U816 (N_816,N_686,N_741);
or U817 (N_817,N_772,N_0);
xor U818 (N_818,In_463,N_504);
xnor U819 (N_819,In_583,In_387);
xor U820 (N_820,N_727,N_625);
nor U821 (N_821,N_425,In_1200);
and U822 (N_822,N_607,In_230);
nand U823 (N_823,In_486,N_355);
nand U824 (N_824,N_419,N_688);
and U825 (N_825,N_762,N_652);
and U826 (N_826,N_539,N_716);
and U827 (N_827,In_283,In_1164);
or U828 (N_828,In_784,N_92);
nand U829 (N_829,In_265,In_1451);
and U830 (N_830,N_291,N_79);
xnor U831 (N_831,In_587,In_644);
nand U832 (N_832,In_339,In_600);
nor U833 (N_833,In_501,N_771);
xnor U834 (N_834,N_786,N_280);
xnor U835 (N_835,In_1268,In_535);
nor U836 (N_836,In_475,N_614);
xnor U837 (N_837,N_450,N_782);
or U838 (N_838,In_1382,In_1447);
or U839 (N_839,N_710,N_382);
and U840 (N_840,In_357,In_1495);
and U841 (N_841,N_662,N_513);
and U842 (N_842,In_1335,In_353);
and U843 (N_843,In_927,N_115);
or U844 (N_844,In_970,N_622);
and U845 (N_845,N_25,In_245);
xor U846 (N_846,N_515,N_557);
and U847 (N_847,In_511,In_956);
nand U848 (N_848,In_627,N_483);
xor U849 (N_849,In_32,N_523);
nor U850 (N_850,N_680,In_614);
xnor U851 (N_851,In_1258,In_1042);
and U852 (N_852,In_1381,N_568);
or U853 (N_853,N_498,N_305);
nand U854 (N_854,N_735,N_317);
and U855 (N_855,N_130,In_279);
xor U856 (N_856,N_582,N_455);
or U857 (N_857,In_826,N_793);
nor U858 (N_858,N_227,N_668);
xor U859 (N_859,In_1285,N_732);
nand U860 (N_860,In_38,N_133);
and U861 (N_861,N_708,In_990);
or U862 (N_862,N_644,In_58);
xor U863 (N_863,N_733,N_676);
xnor U864 (N_864,In_1013,In_728);
nor U865 (N_865,In_1281,N_495);
nor U866 (N_866,In_852,In_569);
nor U867 (N_867,N_798,In_103);
nand U868 (N_868,N_665,In_1108);
nand U869 (N_869,N_237,N_306);
and U870 (N_870,In_1062,N_444);
nor U871 (N_871,N_533,N_705);
nand U872 (N_872,N_388,In_787);
or U873 (N_873,N_608,In_223);
nor U874 (N_874,N_262,N_673);
nor U875 (N_875,In_757,In_712);
nor U876 (N_876,N_308,In_143);
xor U877 (N_877,N_69,N_525);
xnor U878 (N_878,N_454,N_279);
or U879 (N_879,In_1227,In_1203);
and U880 (N_880,N_767,In_670);
nor U881 (N_881,N_753,N_535);
or U882 (N_882,N_67,N_577);
or U883 (N_883,N_592,N_646);
and U884 (N_884,N_558,In_808);
xor U885 (N_885,N_712,N_468);
xor U886 (N_886,In_885,N_302);
xnor U887 (N_887,In_165,In_1056);
and U888 (N_888,N_690,N_124);
nor U889 (N_889,N_569,In_906);
xnor U890 (N_890,N_633,In_1493);
and U891 (N_891,N_466,N_293);
or U892 (N_892,N_621,In_249);
nor U893 (N_893,N_604,In_1023);
and U894 (N_894,In_354,N_785);
or U895 (N_895,N_467,In_432);
and U896 (N_896,N_474,N_546);
or U897 (N_897,N_514,In_963);
and U898 (N_898,N_431,N_189);
nor U899 (N_899,In_781,In_1191);
nand U900 (N_900,In_154,N_307);
nand U901 (N_901,In_1244,In_802);
and U902 (N_902,N_75,In_123);
xnor U903 (N_903,In_485,In_851);
nand U904 (N_904,N_434,N_656);
nor U905 (N_905,N_746,In_755);
xor U906 (N_906,N_620,N_526);
nor U907 (N_907,N_531,In_1306);
or U908 (N_908,N_565,N_734);
xor U909 (N_909,N_598,N_82);
xnor U910 (N_910,N_632,N_740);
or U911 (N_911,N_105,In_1225);
or U912 (N_912,N_590,N_66);
and U913 (N_913,N_586,In_1245);
or U914 (N_914,In_1352,N_703);
or U915 (N_915,In_1387,N_420);
or U916 (N_916,N_182,In_753);
or U917 (N_917,In_938,N_600);
xor U918 (N_918,N_228,In_60);
nor U919 (N_919,N_649,In_15);
and U920 (N_920,N_521,N_640);
and U921 (N_921,In_1354,N_617);
or U922 (N_922,In_1236,In_507);
xnor U923 (N_923,In_231,In_433);
and U924 (N_924,N_276,N_436);
and U925 (N_925,N_200,In_1028);
xor U926 (N_926,N_713,N_547);
xor U927 (N_927,N_106,N_722);
or U928 (N_928,In_447,N_748);
nand U929 (N_929,In_28,In_264);
nand U930 (N_930,N_111,N_647);
nand U931 (N_931,N_594,N_742);
nand U932 (N_932,N_789,In_971);
xnor U933 (N_933,N_671,In_193);
xor U934 (N_934,In_1040,N_730);
or U935 (N_935,In_624,N_768);
xor U936 (N_936,In_783,In_1397);
and U937 (N_937,In_729,In_381);
nand U938 (N_938,N_218,N_677);
and U939 (N_939,N_532,In_1445);
nand U940 (N_940,N_770,N_653);
or U941 (N_941,N_57,N_706);
and U942 (N_942,N_459,N_792);
nand U943 (N_943,N_143,N_661);
or U944 (N_944,N_678,N_267);
nor U945 (N_945,N_790,N_799);
xor U946 (N_946,N_505,In_1432);
xnor U947 (N_947,In_845,N_404);
and U948 (N_948,N_364,In_393);
nor U949 (N_949,N_769,N_699);
nand U950 (N_950,In_1367,N_766);
nand U951 (N_951,In_86,In_920);
nor U952 (N_952,N_725,N_527);
nor U953 (N_953,In_182,N_500);
and U954 (N_954,N_584,N_292);
xor U955 (N_955,In_1489,In_269);
nand U956 (N_956,N_589,In_565);
nand U957 (N_957,N_497,N_739);
xnor U958 (N_958,N_368,N_638);
xnor U959 (N_959,N_775,N_773);
or U960 (N_960,In_662,N_392);
xnor U961 (N_961,N_788,N_335);
xor U962 (N_962,In_417,In_694);
nand U963 (N_963,N_543,N_538);
and U964 (N_964,N_282,N_726);
nor U965 (N_965,N_99,N_443);
nor U966 (N_966,N_266,N_675);
xnor U967 (N_967,In_420,N_683);
and U968 (N_968,N_724,N_744);
nor U969 (N_969,In_1417,N_685);
xnor U970 (N_970,In_537,N_707);
nor U971 (N_971,N_737,N_654);
or U972 (N_972,N_651,N_619);
nand U973 (N_973,N_512,In_861);
xor U974 (N_974,N_650,In_1408);
xor U975 (N_975,N_702,N_658);
or U976 (N_976,N_315,In_700);
or U977 (N_977,N_743,N_136);
nor U978 (N_978,N_215,N_774);
nand U979 (N_979,N_581,N_636);
xor U980 (N_980,In_1396,In_430);
xor U981 (N_981,N_692,In_464);
nor U982 (N_982,N_601,N_615);
or U983 (N_983,In_181,N_701);
and U984 (N_984,N_549,N_414);
and U985 (N_985,In_665,In_778);
nand U986 (N_986,N_52,In_985);
xnor U987 (N_987,N_216,In_278);
nand U988 (N_988,N_398,N_627);
nand U989 (N_989,N_332,N_36);
and U990 (N_990,N_698,N_23);
nand U991 (N_991,In_641,In_256);
nand U992 (N_992,In_766,N_655);
xnor U993 (N_993,N_387,N_562);
nand U994 (N_994,N_240,N_475);
xnor U995 (N_995,N_796,N_728);
or U996 (N_996,N_750,In_709);
xnor U997 (N_997,N_367,N_787);
nand U998 (N_998,In_568,N_736);
nor U999 (N_999,In_782,In_36);
or U1000 (N_1000,N_687,N_980);
and U1001 (N_1001,N_908,N_987);
or U1002 (N_1002,N_684,N_827);
nor U1003 (N_1003,N_679,In_1207);
and U1004 (N_1004,N_966,N_624);
nor U1005 (N_1005,In_1241,N_853);
nand U1006 (N_1006,In_1209,N_24);
xnor U1007 (N_1007,N_634,N_917);
xnor U1008 (N_1008,In_400,N_611);
nor U1009 (N_1009,N_855,In_590);
and U1010 (N_1010,In_1060,N_931);
nand U1011 (N_1011,N_369,N_912);
or U1012 (N_1012,N_964,N_795);
or U1013 (N_1013,In_1201,N_610);
nand U1014 (N_1014,In_858,N_911);
or U1015 (N_1015,N_720,N_666);
and U1016 (N_1016,N_875,N_631);
xnor U1017 (N_1017,In_1275,N_894);
and U1018 (N_1018,N_877,N_916);
nor U1019 (N_1019,N_524,N_955);
nand U1020 (N_1020,N_756,N_791);
and U1021 (N_1021,N_937,N_982);
or U1022 (N_1022,In_1431,N_84);
or U1023 (N_1023,N_87,N_672);
xnor U1024 (N_1024,In_1298,N_682);
nand U1025 (N_1025,N_602,In_563);
and U1026 (N_1026,N_889,N_755);
xor U1027 (N_1027,N_806,N_898);
xnor U1028 (N_1028,N_696,N_970);
and U1029 (N_1029,In_593,N_880);
nor U1030 (N_1030,N_191,In_428);
or U1031 (N_1031,N_999,In_341);
and U1032 (N_1032,N_847,N_974);
and U1033 (N_1033,N_405,N_709);
and U1034 (N_1034,N_571,N_499);
or U1035 (N_1035,In_351,N_885);
and U1036 (N_1036,N_893,N_886);
or U1037 (N_1037,In_730,N_909);
xor U1038 (N_1038,N_933,In_235);
nand U1039 (N_1039,N_947,N_758);
or U1040 (N_1040,N_884,In_598);
nand U1041 (N_1041,In_827,N_418);
nand U1042 (N_1042,In_604,N_950);
xor U1043 (N_1043,N_965,N_961);
or U1044 (N_1044,N_346,N_996);
nand U1045 (N_1045,N_890,N_883);
nor U1046 (N_1046,N_952,N_463);
xor U1047 (N_1047,N_828,In_224);
or U1048 (N_1048,N_975,N_778);
xor U1049 (N_1049,In_228,N_956);
xor U1050 (N_1050,N_958,In_1136);
nor U1051 (N_1051,N_729,N_751);
or U1052 (N_1052,In_1075,N_642);
xor U1053 (N_1053,N_393,N_819);
and U1054 (N_1054,N_100,N_954);
nand U1055 (N_1055,N_932,In_687);
or U1056 (N_1056,In_577,N_464);
and U1057 (N_1057,N_372,N_208);
and U1058 (N_1058,N_576,N_72);
xnor U1059 (N_1059,N_997,N_113);
or U1060 (N_1060,N_674,N_988);
or U1061 (N_1061,N_643,N_344);
nand U1062 (N_1062,N_16,N_101);
or U1063 (N_1063,In_899,In_578);
nor U1064 (N_1064,N_816,In_680);
nor U1065 (N_1065,N_835,N_807);
xnor U1066 (N_1066,In_1197,In_1239);
and U1067 (N_1067,N_915,In_524);
and U1068 (N_1068,In_1347,In_761);
nor U1069 (N_1069,N_861,N_628);
xnor U1070 (N_1070,N_479,N_869);
and U1071 (N_1071,N_896,In_252);
and U1072 (N_1072,N_923,N_415);
nand U1073 (N_1073,In_926,N_843);
xnor U1074 (N_1074,N_629,In_1376);
and U1075 (N_1075,In_992,N_422);
xnor U1076 (N_1076,In_190,N_478);
nand U1077 (N_1077,N_948,N_609);
xnor U1078 (N_1078,N_818,In_629);
xor U1079 (N_1079,In_514,N_920);
and U1080 (N_1080,N_944,N_817);
or U1081 (N_1081,In_1032,N_844);
xnor U1082 (N_1082,In_1442,N_242);
and U1083 (N_1083,N_830,N_977);
and U1084 (N_1084,N_852,N_868);
nand U1085 (N_1085,N_992,N_752);
nor U1086 (N_1086,N_518,N_541);
nand U1087 (N_1087,N_951,N_978);
and U1088 (N_1088,N_718,N_942);
nor U1089 (N_1089,N_823,N_881);
xnor U1090 (N_1090,N_929,N_935);
or U1091 (N_1091,In_482,N_171);
nor U1092 (N_1092,N_973,N_664);
or U1093 (N_1093,N_472,N_821);
nand U1094 (N_1094,N_578,N_913);
xnor U1095 (N_1095,N_159,N_829);
nor U1096 (N_1096,N_826,In_571);
xor U1097 (N_1097,N_104,N_969);
and U1098 (N_1098,N_836,N_385);
or U1099 (N_1099,In_1344,N_715);
nor U1100 (N_1100,N_33,N_700);
nor U1101 (N_1101,N_850,N_863);
or U1102 (N_1102,N_156,N_926);
and U1103 (N_1103,In_816,N_848);
or U1104 (N_1104,N_812,In_50);
nand U1105 (N_1105,N_765,In_647);
nand U1106 (N_1106,N_695,N_906);
nor U1107 (N_1107,N_919,N_993);
nand U1108 (N_1108,N_811,N_324);
xor U1109 (N_1109,N_887,N_122);
xnor U1110 (N_1110,N_637,N_757);
nand U1111 (N_1111,In_1486,N_747);
and U1112 (N_1112,N_959,N_559);
nor U1113 (N_1113,N_339,N_83);
or U1114 (N_1114,N_271,In_1327);
or U1115 (N_1115,N_359,In_1242);
or U1116 (N_1116,N_131,In_1353);
nand U1117 (N_1117,N_902,In_1324);
nand U1118 (N_1118,N_477,N_839);
xnor U1119 (N_1119,N_858,In_796);
and U1120 (N_1120,In_496,In_540);
or U1121 (N_1121,In_842,N_489);
nor U1122 (N_1122,N_803,N_281);
or U1123 (N_1123,N_901,N_810);
and U1124 (N_1124,In_1301,N_693);
xor U1125 (N_1125,In_867,N_934);
xnor U1126 (N_1126,In_94,N_777);
or U1127 (N_1127,N_907,N_888);
nor U1128 (N_1128,In_925,N_878);
xor U1129 (N_1129,N_862,N_764);
nand U1130 (N_1130,N_957,N_903);
nor U1131 (N_1131,In_323,N_623);
or U1132 (N_1132,N_872,N_800);
or U1133 (N_1133,N_612,N_831);
xor U1134 (N_1134,N_626,N_618);
nor U1135 (N_1135,N_347,In_1116);
nor U1136 (N_1136,N_936,N_731);
nor U1137 (N_1137,N_605,N_941);
nand U1138 (N_1138,N_924,N_465);
nor U1139 (N_1139,N_548,In_1140);
and U1140 (N_1140,N_986,In_116);
xor U1141 (N_1141,N_984,N_865);
nor U1142 (N_1142,N_400,N_925);
and U1143 (N_1143,In_510,In_76);
and U1144 (N_1144,In_444,In_1491);
and U1145 (N_1145,In_993,N_648);
nor U1146 (N_1146,N_985,N_447);
xor U1147 (N_1147,N_669,N_905);
nand U1148 (N_1148,In_1485,N_849);
nand U1149 (N_1149,N_857,In_386);
nor U1150 (N_1150,N_432,N_873);
nand U1151 (N_1151,N_691,In_352);
xor U1152 (N_1152,In_412,N_953);
nor U1153 (N_1153,N_784,N_837);
and U1154 (N_1154,In_494,N_238);
nand U1155 (N_1155,N_928,N_864);
nor U1156 (N_1156,N_976,In_739);
nand U1157 (N_1157,N_938,N_871);
nand U1158 (N_1158,In_33,N_990);
xnor U1159 (N_1159,In_1041,N_484);
and U1160 (N_1160,N_711,N_641);
xnor U1161 (N_1161,N_979,N_824);
nor U1162 (N_1162,In_1436,N_776);
nor U1163 (N_1163,N_921,N_214);
nor U1164 (N_1164,In_241,N_599);
or U1165 (N_1165,N_763,N_943);
nor U1166 (N_1166,N_667,In_1276);
xnor U1167 (N_1167,N_681,N_704);
xnor U1168 (N_1168,N_842,N_840);
or U1169 (N_1169,In_225,N_128);
or U1170 (N_1170,N_822,In_1407);
xor U1171 (N_1171,N_222,N_343);
nor U1172 (N_1172,In_1218,N_879);
nor U1173 (N_1173,N_399,N_813);
or U1174 (N_1174,N_841,N_991);
and U1175 (N_1175,N_376,N_882);
nor U1176 (N_1176,In_848,N_876);
and U1177 (N_1177,N_760,N_946);
or U1178 (N_1178,In_1036,N_838);
and U1179 (N_1179,In_1329,N_820);
nor U1180 (N_1180,N_714,N_900);
nor U1181 (N_1181,N_989,N_899);
nor U1182 (N_1182,N_854,N_825);
nor U1183 (N_1183,N_603,N_606);
xor U1184 (N_1184,N_244,N_870);
nand U1185 (N_1185,In_550,N_273);
nand U1186 (N_1186,In_643,N_834);
and U1187 (N_1187,N_910,N_780);
or U1188 (N_1188,N_918,N_859);
and U1189 (N_1189,In_1345,N_804);
nor U1190 (N_1190,N_867,In_1113);
nor U1191 (N_1191,N_994,N_851);
or U1192 (N_1192,N_125,N_971);
xnor U1193 (N_1193,N_759,In_1105);
and U1194 (N_1194,N_866,In_1421);
xor U1195 (N_1195,N_967,N_998);
and U1196 (N_1196,N_721,N_168);
nand U1197 (N_1197,In_1017,In_1411);
and U1198 (N_1198,In_1194,N_210);
xnor U1199 (N_1199,N_3,N_802);
nor U1200 (N_1200,N_660,N_1051);
and U1201 (N_1201,N_1161,N_485);
or U1202 (N_1202,N_779,In_810);
xnor U1203 (N_1203,In_63,N_1016);
nor U1204 (N_1204,N_1085,N_781);
xnor U1205 (N_1205,N_1185,N_1110);
xnor U1206 (N_1206,N_1046,N_749);
nand U1207 (N_1207,N_949,In_1456);
nand U1208 (N_1208,N_456,N_1083);
or U1209 (N_1209,N_1058,N_717);
and U1210 (N_1210,N_1167,N_808);
nand U1211 (N_1211,N_1025,N_1176);
and U1212 (N_1212,N_1104,N_1098);
xnor U1213 (N_1213,N_1129,N_1108);
nand U1214 (N_1214,N_1160,N_1030);
nor U1215 (N_1215,N_1139,N_1078);
nand U1216 (N_1216,N_1173,N_983);
nand U1217 (N_1217,N_1124,N_1140);
xor U1218 (N_1218,N_1162,N_1197);
or U1219 (N_1219,N_1152,N_1113);
or U1220 (N_1220,N_1195,N_1024);
and U1221 (N_1221,N_1069,N_1023);
and U1222 (N_1222,N_1116,N_1087);
and U1223 (N_1223,N_1045,N_1182);
nand U1224 (N_1224,N_1050,N_1036);
xnor U1225 (N_1225,N_1155,N_1177);
or U1226 (N_1226,N_1187,In_636);
xnor U1227 (N_1227,N_1114,In_275);
xor U1228 (N_1228,N_1099,N_801);
nand U1229 (N_1229,N_1164,N_1000);
xor U1230 (N_1230,N_1004,N_797);
nand U1231 (N_1231,N_814,N_1014);
xor U1232 (N_1232,In_974,N_1052);
nand U1233 (N_1233,N_1165,N_809);
and U1234 (N_1234,N_1148,N_322);
and U1235 (N_1235,N_345,N_856);
xor U1236 (N_1236,N_1077,N_1035);
nor U1237 (N_1237,N_1076,N_1138);
or U1238 (N_1238,N_73,N_1112);
nor U1239 (N_1239,N_1001,N_1175);
and U1240 (N_1240,N_1181,N_904);
and U1241 (N_1241,N_1169,N_1088);
nor U1242 (N_1242,N_1101,N_1017);
or U1243 (N_1243,In_530,N_897);
or U1244 (N_1244,N_1084,N_1071);
nor U1245 (N_1245,N_1153,N_1082);
or U1246 (N_1246,In_314,N_723);
nor U1247 (N_1247,N_1003,N_1072);
nor U1248 (N_1248,N_1190,N_1193);
xor U1249 (N_1249,N_1102,N_1070);
nor U1250 (N_1250,N_914,N_694);
nor U1251 (N_1251,N_1199,N_1037);
nor U1252 (N_1252,N_1141,N_1020);
or U1253 (N_1253,N_1150,N_922);
nor U1254 (N_1254,N_1127,N_805);
nor U1255 (N_1255,N_573,N_230);
and U1256 (N_1256,N_945,N_1057);
or U1257 (N_1257,N_1128,N_1029);
and U1258 (N_1258,N_1005,N_1130);
nor U1259 (N_1259,N_1147,N_689);
or U1260 (N_1260,N_846,In_791);
nor U1261 (N_1261,N_745,N_940);
nand U1262 (N_1262,N_697,N_1040);
or U1263 (N_1263,N_1094,N_1031);
nand U1264 (N_1264,N_616,N_1043);
or U1265 (N_1265,N_1038,N_1015);
and U1266 (N_1266,N_471,N_1186);
xnor U1267 (N_1267,In_72,N_874);
nor U1268 (N_1268,N_1053,In_340);
xor U1269 (N_1269,N_1068,N_891);
nor U1270 (N_1270,N_939,N_1032);
nand U1271 (N_1271,N_1097,N_1146);
nor U1272 (N_1272,N_1196,N_1066);
nor U1273 (N_1273,N_815,N_1171);
or U1274 (N_1274,N_972,N_1075);
or U1275 (N_1275,N_892,N_1151);
xnor U1276 (N_1276,N_968,N_1158);
and U1277 (N_1277,N_1047,N_1118);
nor U1278 (N_1278,N_1134,In_186);
nand U1279 (N_1279,N_1091,N_1188);
nand U1280 (N_1280,N_1132,N_1);
and U1281 (N_1281,N_1157,N_930);
or U1282 (N_1282,N_1093,In_1339);
or U1283 (N_1283,N_832,N_1149);
or U1284 (N_1284,N_1198,N_1121);
nand U1285 (N_1285,N_545,In_1139);
or U1286 (N_1286,N_1065,N_1009);
xor U1287 (N_1287,In_863,N_1049);
and U1288 (N_1288,N_1095,N_1081);
or U1289 (N_1289,N_544,N_1063);
nor U1290 (N_1290,N_895,N_1067);
and U1291 (N_1291,N_1166,N_1194);
xnor U1292 (N_1292,N_960,N_1089);
or U1293 (N_1293,In_1465,N_1055);
or U1294 (N_1294,N_1191,In_1343);
xnor U1295 (N_1295,N_1021,N_1143);
nand U1296 (N_1296,N_1056,In_682);
and U1297 (N_1297,N_1142,N_294);
nor U1298 (N_1298,N_1117,N_670);
or U1299 (N_1299,N_1096,In_288);
or U1300 (N_1300,N_1180,N_1145);
xnor U1301 (N_1301,N_1044,N_1007);
nor U1302 (N_1302,N_1074,N_1106);
xnor U1303 (N_1303,N_860,N_1136);
nor U1304 (N_1304,N_1135,N_833);
or U1305 (N_1305,N_1183,N_1027);
or U1306 (N_1306,N_1115,In_526);
and U1307 (N_1307,N_596,N_1189);
xor U1308 (N_1308,N_1062,N_1048);
and U1309 (N_1309,N_981,N_1086);
nand U1310 (N_1310,N_1126,N_26);
nor U1311 (N_1311,N_123,N_1008);
nand U1312 (N_1312,N_1111,N_1006);
or U1313 (N_1313,N_457,N_1073);
nand U1314 (N_1314,N_962,N_1107);
nor U1315 (N_1315,N_738,N_1041);
nor U1316 (N_1316,N_1156,N_1172);
xnor U1317 (N_1317,N_1011,N_1174);
nand U1318 (N_1318,N_1154,N_1092);
nand U1319 (N_1319,N_995,N_1179);
nand U1320 (N_1320,N_1059,N_117);
nand U1321 (N_1321,N_327,N_1090);
nand U1322 (N_1322,N_1012,N_1170);
or U1323 (N_1323,N_1060,N_1033);
and U1324 (N_1324,N_659,In_145);
and U1325 (N_1325,N_1054,N_1018);
nand U1326 (N_1326,N_1137,N_1019);
xnor U1327 (N_1327,N_509,N_1105);
nand U1328 (N_1328,N_461,N_1010);
xnor U1329 (N_1329,N_1100,N_1168);
nor U1330 (N_1330,N_1120,N_1163);
nor U1331 (N_1331,In_42,N_1042);
or U1332 (N_1332,N_402,N_1103);
nor U1333 (N_1333,N_1028,N_1109);
nand U1334 (N_1334,N_1026,N_1184);
nand U1335 (N_1335,In_711,N_1122);
nor U1336 (N_1336,N_426,N_1013);
nor U1337 (N_1337,N_845,N_1192);
nand U1338 (N_1338,N_1144,N_353);
nor U1339 (N_1339,N_1002,N_1039);
nand U1340 (N_1340,N_927,N_630);
and U1341 (N_1341,N_1061,In_301);
nand U1342 (N_1342,N_1119,N_1034);
or U1343 (N_1343,N_1022,N_1178);
or U1344 (N_1344,N_1159,N_639);
xnor U1345 (N_1345,N_1125,N_1080);
nand U1346 (N_1346,N_1079,N_1133);
xor U1347 (N_1347,N_1064,N_1131);
nor U1348 (N_1348,N_1123,N_563);
xnor U1349 (N_1349,N_963,N_754);
xnor U1350 (N_1350,N_1135,N_660);
nand U1351 (N_1351,N_1082,N_1007);
nand U1352 (N_1352,N_1163,N_960);
and U1353 (N_1353,N_73,N_1192);
and U1354 (N_1354,N_456,N_117);
xnor U1355 (N_1355,N_697,N_930);
and U1356 (N_1356,N_983,N_639);
nor U1357 (N_1357,N_1130,N_1074);
nand U1358 (N_1358,In_1456,N_1040);
or U1359 (N_1359,N_981,In_530);
or U1360 (N_1360,N_1157,N_1186);
nor U1361 (N_1361,N_1185,N_1111);
nand U1362 (N_1362,N_1143,N_1037);
or U1363 (N_1363,N_327,N_1182);
or U1364 (N_1364,N_1145,N_1032);
xnor U1365 (N_1365,N_1103,N_456);
nand U1366 (N_1366,N_1040,N_1168);
nand U1367 (N_1367,N_738,N_1098);
nand U1368 (N_1368,N_1074,N_1073);
nand U1369 (N_1369,N_895,N_1181);
or U1370 (N_1370,N_963,N_1025);
nor U1371 (N_1371,N_1067,N_294);
nor U1372 (N_1372,N_616,N_1121);
nand U1373 (N_1373,N_1028,N_1141);
nand U1374 (N_1374,N_1089,N_1095);
and U1375 (N_1375,N_1075,N_754);
nand U1376 (N_1376,N_1158,N_1096);
and U1377 (N_1377,N_1013,In_340);
xnor U1378 (N_1378,N_1128,N_1176);
nor U1379 (N_1379,N_1078,N_1019);
nor U1380 (N_1380,N_509,N_717);
or U1381 (N_1381,N_1105,N_1010);
and U1382 (N_1382,N_1070,N_1167);
and U1383 (N_1383,N_1073,N_1141);
or U1384 (N_1384,N_1082,N_1039);
and U1385 (N_1385,N_230,N_1166);
and U1386 (N_1386,N_1121,N_1048);
xnor U1387 (N_1387,N_1072,N_1118);
and U1388 (N_1388,N_1078,N_1077);
and U1389 (N_1389,In_636,In_288);
or U1390 (N_1390,N_801,N_1146);
and U1391 (N_1391,N_1032,N_940);
nand U1392 (N_1392,N_1067,N_1169);
and U1393 (N_1393,N_1194,N_1185);
xnor U1394 (N_1394,N_596,N_968);
xor U1395 (N_1395,N_939,N_1006);
and U1396 (N_1396,N_927,N_717);
and U1397 (N_1397,N_981,N_1057);
nor U1398 (N_1398,N_1029,N_1116);
nand U1399 (N_1399,N_1162,N_1169);
nand U1400 (N_1400,N_1357,N_1262);
xor U1401 (N_1401,N_1393,N_1226);
or U1402 (N_1402,N_1261,N_1290);
nand U1403 (N_1403,N_1379,N_1342);
and U1404 (N_1404,N_1306,N_1370);
or U1405 (N_1405,N_1236,N_1256);
nand U1406 (N_1406,N_1211,N_1221);
nor U1407 (N_1407,N_1229,N_1216);
and U1408 (N_1408,N_1279,N_1314);
and U1409 (N_1409,N_1209,N_1249);
nor U1410 (N_1410,N_1259,N_1277);
nand U1411 (N_1411,N_1337,N_1207);
nor U1412 (N_1412,N_1394,N_1202);
xnor U1413 (N_1413,N_1364,N_1358);
nand U1414 (N_1414,N_1371,N_1372);
xor U1415 (N_1415,N_1285,N_1374);
nand U1416 (N_1416,N_1299,N_1347);
or U1417 (N_1417,N_1389,N_1270);
or U1418 (N_1418,N_1242,N_1341);
nor U1419 (N_1419,N_1344,N_1243);
and U1420 (N_1420,N_1291,N_1377);
nand U1421 (N_1421,N_1296,N_1362);
or U1422 (N_1422,N_1395,N_1361);
xor U1423 (N_1423,N_1302,N_1324);
and U1424 (N_1424,N_1235,N_1293);
xor U1425 (N_1425,N_1227,N_1263);
or U1426 (N_1426,N_1315,N_1303);
or U1427 (N_1427,N_1297,N_1248);
and U1428 (N_1428,N_1334,N_1366);
nor U1429 (N_1429,N_1311,N_1355);
nor U1430 (N_1430,N_1266,N_1320);
nand U1431 (N_1431,N_1304,N_1330);
xnor U1432 (N_1432,N_1203,N_1278);
nand U1433 (N_1433,N_1219,N_1369);
or U1434 (N_1434,N_1222,N_1289);
and U1435 (N_1435,N_1295,N_1252);
and U1436 (N_1436,N_1386,N_1368);
nor U1437 (N_1437,N_1231,N_1367);
nand U1438 (N_1438,N_1391,N_1325);
and U1439 (N_1439,N_1275,N_1359);
xor U1440 (N_1440,N_1392,N_1271);
xor U1441 (N_1441,N_1310,N_1268);
and U1442 (N_1442,N_1354,N_1336);
and U1443 (N_1443,N_1329,N_1380);
nor U1444 (N_1444,N_1382,N_1308);
and U1445 (N_1445,N_1287,N_1399);
and U1446 (N_1446,N_1265,N_1321);
nor U1447 (N_1447,N_1232,N_1381);
or U1448 (N_1448,N_1345,N_1346);
nor U1449 (N_1449,N_1319,N_1230);
or U1450 (N_1450,N_1333,N_1282);
or U1451 (N_1451,N_1356,N_1339);
and U1452 (N_1452,N_1280,N_1388);
or U1453 (N_1453,N_1288,N_1352);
nand U1454 (N_1454,N_1228,N_1241);
xor U1455 (N_1455,N_1326,N_1301);
and U1456 (N_1456,N_1237,N_1281);
nor U1457 (N_1457,N_1384,N_1273);
or U1458 (N_1458,N_1218,N_1349);
and U1459 (N_1459,N_1267,N_1383);
xor U1460 (N_1460,N_1378,N_1213);
nand U1461 (N_1461,N_1307,N_1253);
xnor U1462 (N_1462,N_1343,N_1206);
nor U1463 (N_1463,N_1251,N_1254);
and U1464 (N_1464,N_1269,N_1244);
nor U1465 (N_1465,N_1286,N_1340);
xor U1466 (N_1466,N_1322,N_1257);
xor U1467 (N_1467,N_1387,N_1215);
xor U1468 (N_1468,N_1376,N_1390);
or U1469 (N_1469,N_1375,N_1365);
xor U1470 (N_1470,N_1255,N_1208);
nor U1471 (N_1471,N_1245,N_1283);
or U1472 (N_1472,N_1335,N_1398);
nor U1473 (N_1473,N_1204,N_1348);
nand U1474 (N_1474,N_1328,N_1294);
xnor U1475 (N_1475,N_1247,N_1201);
nor U1476 (N_1476,N_1238,N_1234);
or U1477 (N_1477,N_1309,N_1360);
nor U1478 (N_1478,N_1212,N_1250);
and U1479 (N_1479,N_1317,N_1318);
and U1480 (N_1480,N_1233,N_1385);
and U1481 (N_1481,N_1225,N_1210);
and U1482 (N_1482,N_1260,N_1353);
and U1483 (N_1483,N_1332,N_1305);
xnor U1484 (N_1484,N_1258,N_1300);
nor U1485 (N_1485,N_1351,N_1240);
xnor U1486 (N_1486,N_1292,N_1298);
and U1487 (N_1487,N_1396,N_1338);
xor U1488 (N_1488,N_1363,N_1276);
or U1489 (N_1489,N_1214,N_1264);
nor U1490 (N_1490,N_1373,N_1323);
and U1491 (N_1491,N_1220,N_1239);
or U1492 (N_1492,N_1224,N_1205);
and U1493 (N_1493,N_1350,N_1284);
or U1494 (N_1494,N_1274,N_1397);
xnor U1495 (N_1495,N_1312,N_1313);
or U1496 (N_1496,N_1331,N_1316);
nand U1497 (N_1497,N_1223,N_1272);
xnor U1498 (N_1498,N_1327,N_1246);
or U1499 (N_1499,N_1200,N_1217);
or U1500 (N_1500,N_1237,N_1261);
and U1501 (N_1501,N_1329,N_1307);
and U1502 (N_1502,N_1344,N_1245);
nor U1503 (N_1503,N_1290,N_1276);
xnor U1504 (N_1504,N_1218,N_1265);
and U1505 (N_1505,N_1378,N_1374);
or U1506 (N_1506,N_1283,N_1343);
xnor U1507 (N_1507,N_1383,N_1305);
nor U1508 (N_1508,N_1224,N_1342);
nand U1509 (N_1509,N_1354,N_1319);
nand U1510 (N_1510,N_1361,N_1371);
or U1511 (N_1511,N_1336,N_1369);
xor U1512 (N_1512,N_1340,N_1247);
nor U1513 (N_1513,N_1384,N_1356);
xnor U1514 (N_1514,N_1250,N_1252);
xnor U1515 (N_1515,N_1314,N_1211);
or U1516 (N_1516,N_1303,N_1281);
nand U1517 (N_1517,N_1216,N_1372);
nand U1518 (N_1518,N_1215,N_1293);
nor U1519 (N_1519,N_1351,N_1245);
nor U1520 (N_1520,N_1329,N_1291);
and U1521 (N_1521,N_1379,N_1290);
and U1522 (N_1522,N_1316,N_1247);
nand U1523 (N_1523,N_1323,N_1205);
nor U1524 (N_1524,N_1221,N_1392);
xnor U1525 (N_1525,N_1300,N_1303);
nor U1526 (N_1526,N_1274,N_1222);
nand U1527 (N_1527,N_1219,N_1217);
nand U1528 (N_1528,N_1234,N_1218);
xor U1529 (N_1529,N_1320,N_1270);
or U1530 (N_1530,N_1221,N_1294);
nand U1531 (N_1531,N_1394,N_1205);
nand U1532 (N_1532,N_1315,N_1251);
nand U1533 (N_1533,N_1365,N_1203);
nand U1534 (N_1534,N_1328,N_1273);
nor U1535 (N_1535,N_1228,N_1376);
or U1536 (N_1536,N_1222,N_1215);
xor U1537 (N_1537,N_1357,N_1258);
nand U1538 (N_1538,N_1347,N_1219);
nand U1539 (N_1539,N_1306,N_1290);
xnor U1540 (N_1540,N_1269,N_1298);
nor U1541 (N_1541,N_1217,N_1233);
and U1542 (N_1542,N_1379,N_1209);
nor U1543 (N_1543,N_1279,N_1240);
xor U1544 (N_1544,N_1358,N_1261);
or U1545 (N_1545,N_1338,N_1205);
or U1546 (N_1546,N_1289,N_1312);
nor U1547 (N_1547,N_1361,N_1327);
and U1548 (N_1548,N_1246,N_1298);
nor U1549 (N_1549,N_1373,N_1344);
or U1550 (N_1550,N_1378,N_1295);
xnor U1551 (N_1551,N_1311,N_1372);
xnor U1552 (N_1552,N_1203,N_1236);
or U1553 (N_1553,N_1357,N_1391);
nor U1554 (N_1554,N_1398,N_1355);
xor U1555 (N_1555,N_1266,N_1346);
and U1556 (N_1556,N_1308,N_1235);
nand U1557 (N_1557,N_1362,N_1395);
nand U1558 (N_1558,N_1224,N_1358);
and U1559 (N_1559,N_1317,N_1264);
xor U1560 (N_1560,N_1326,N_1314);
and U1561 (N_1561,N_1304,N_1253);
and U1562 (N_1562,N_1200,N_1242);
xor U1563 (N_1563,N_1364,N_1392);
and U1564 (N_1564,N_1374,N_1297);
nand U1565 (N_1565,N_1302,N_1364);
nand U1566 (N_1566,N_1341,N_1319);
nand U1567 (N_1567,N_1231,N_1387);
and U1568 (N_1568,N_1319,N_1394);
xnor U1569 (N_1569,N_1249,N_1270);
nand U1570 (N_1570,N_1302,N_1338);
and U1571 (N_1571,N_1332,N_1315);
or U1572 (N_1572,N_1230,N_1268);
or U1573 (N_1573,N_1268,N_1206);
and U1574 (N_1574,N_1292,N_1284);
nor U1575 (N_1575,N_1286,N_1386);
and U1576 (N_1576,N_1298,N_1202);
and U1577 (N_1577,N_1373,N_1212);
and U1578 (N_1578,N_1372,N_1251);
nand U1579 (N_1579,N_1211,N_1289);
xor U1580 (N_1580,N_1353,N_1202);
xor U1581 (N_1581,N_1289,N_1261);
and U1582 (N_1582,N_1305,N_1304);
nand U1583 (N_1583,N_1288,N_1299);
xor U1584 (N_1584,N_1279,N_1362);
and U1585 (N_1585,N_1307,N_1366);
and U1586 (N_1586,N_1387,N_1334);
xor U1587 (N_1587,N_1245,N_1234);
xor U1588 (N_1588,N_1350,N_1349);
nand U1589 (N_1589,N_1296,N_1288);
or U1590 (N_1590,N_1327,N_1364);
nand U1591 (N_1591,N_1273,N_1220);
or U1592 (N_1592,N_1287,N_1355);
nand U1593 (N_1593,N_1229,N_1399);
or U1594 (N_1594,N_1373,N_1393);
nand U1595 (N_1595,N_1230,N_1201);
nor U1596 (N_1596,N_1292,N_1234);
xor U1597 (N_1597,N_1358,N_1200);
and U1598 (N_1598,N_1338,N_1375);
xnor U1599 (N_1599,N_1239,N_1297);
nor U1600 (N_1600,N_1503,N_1484);
nand U1601 (N_1601,N_1402,N_1568);
and U1602 (N_1602,N_1467,N_1440);
xnor U1603 (N_1603,N_1526,N_1561);
nor U1604 (N_1604,N_1500,N_1448);
or U1605 (N_1605,N_1567,N_1487);
or U1606 (N_1606,N_1439,N_1590);
and U1607 (N_1607,N_1514,N_1428);
xor U1608 (N_1608,N_1494,N_1471);
xnor U1609 (N_1609,N_1545,N_1447);
or U1610 (N_1610,N_1411,N_1430);
nand U1611 (N_1611,N_1585,N_1466);
nor U1612 (N_1612,N_1596,N_1420);
or U1613 (N_1613,N_1505,N_1453);
and U1614 (N_1614,N_1588,N_1501);
and U1615 (N_1615,N_1455,N_1509);
or U1616 (N_1616,N_1424,N_1523);
and U1617 (N_1617,N_1542,N_1513);
or U1618 (N_1618,N_1525,N_1574);
and U1619 (N_1619,N_1499,N_1597);
and U1620 (N_1620,N_1481,N_1539);
xnor U1621 (N_1621,N_1422,N_1463);
xnor U1622 (N_1622,N_1479,N_1493);
nor U1623 (N_1623,N_1496,N_1524);
xnor U1624 (N_1624,N_1584,N_1409);
xnor U1625 (N_1625,N_1556,N_1446);
nor U1626 (N_1626,N_1470,N_1593);
or U1627 (N_1627,N_1401,N_1461);
and U1628 (N_1628,N_1576,N_1432);
xor U1629 (N_1629,N_1478,N_1450);
nand U1630 (N_1630,N_1480,N_1591);
nor U1631 (N_1631,N_1595,N_1414);
and U1632 (N_1632,N_1594,N_1598);
or U1633 (N_1633,N_1502,N_1537);
nand U1634 (N_1634,N_1551,N_1541);
and U1635 (N_1635,N_1435,N_1511);
nand U1636 (N_1636,N_1578,N_1528);
and U1637 (N_1637,N_1571,N_1452);
nor U1638 (N_1638,N_1538,N_1485);
or U1639 (N_1639,N_1400,N_1498);
or U1640 (N_1640,N_1469,N_1549);
or U1641 (N_1641,N_1504,N_1583);
nor U1642 (N_1642,N_1429,N_1550);
nand U1643 (N_1643,N_1433,N_1460);
nor U1644 (N_1644,N_1415,N_1475);
nor U1645 (N_1645,N_1405,N_1510);
and U1646 (N_1646,N_1572,N_1410);
and U1647 (N_1647,N_1560,N_1554);
nor U1648 (N_1648,N_1407,N_1477);
nand U1649 (N_1649,N_1419,N_1425);
nor U1650 (N_1650,N_1559,N_1497);
or U1651 (N_1651,N_1474,N_1530);
or U1652 (N_1652,N_1412,N_1473);
nand U1653 (N_1653,N_1516,N_1581);
and U1654 (N_1654,N_1490,N_1417);
xor U1655 (N_1655,N_1544,N_1580);
xnor U1656 (N_1656,N_1437,N_1468);
and U1657 (N_1657,N_1427,N_1575);
or U1658 (N_1658,N_1413,N_1406);
and U1659 (N_1659,N_1536,N_1472);
or U1660 (N_1660,N_1529,N_1531);
nor U1661 (N_1661,N_1535,N_1423);
nor U1662 (N_1662,N_1486,N_1518);
and U1663 (N_1663,N_1403,N_1570);
and U1664 (N_1664,N_1586,N_1507);
and U1665 (N_1665,N_1459,N_1519);
xor U1666 (N_1666,N_1443,N_1488);
nand U1667 (N_1667,N_1555,N_1558);
xnor U1668 (N_1668,N_1482,N_1547);
nor U1669 (N_1669,N_1562,N_1442);
and U1670 (N_1670,N_1416,N_1548);
and U1671 (N_1671,N_1457,N_1464);
or U1672 (N_1672,N_1579,N_1589);
and U1673 (N_1673,N_1506,N_1517);
and U1674 (N_1674,N_1564,N_1512);
nand U1675 (N_1675,N_1532,N_1465);
nor U1676 (N_1676,N_1444,N_1404);
xnor U1677 (N_1677,N_1495,N_1492);
and U1678 (N_1678,N_1563,N_1426);
and U1679 (N_1679,N_1599,N_1582);
xor U1680 (N_1680,N_1454,N_1491);
nand U1681 (N_1681,N_1557,N_1587);
xnor U1682 (N_1682,N_1515,N_1436);
xnor U1683 (N_1683,N_1438,N_1458);
and U1684 (N_1684,N_1441,N_1527);
xnor U1685 (N_1685,N_1577,N_1456);
xor U1686 (N_1686,N_1592,N_1565);
nand U1687 (N_1687,N_1483,N_1462);
and U1688 (N_1688,N_1566,N_1543);
nor U1689 (N_1689,N_1408,N_1534);
and U1690 (N_1690,N_1421,N_1489);
nand U1691 (N_1691,N_1546,N_1533);
xor U1692 (N_1692,N_1569,N_1476);
or U1693 (N_1693,N_1553,N_1431);
or U1694 (N_1694,N_1521,N_1445);
nand U1695 (N_1695,N_1520,N_1540);
xnor U1696 (N_1696,N_1451,N_1449);
xnor U1697 (N_1697,N_1508,N_1552);
xnor U1698 (N_1698,N_1573,N_1418);
nand U1699 (N_1699,N_1434,N_1522);
or U1700 (N_1700,N_1574,N_1529);
nand U1701 (N_1701,N_1419,N_1434);
and U1702 (N_1702,N_1456,N_1558);
or U1703 (N_1703,N_1414,N_1596);
nand U1704 (N_1704,N_1420,N_1554);
nor U1705 (N_1705,N_1444,N_1546);
xor U1706 (N_1706,N_1583,N_1560);
or U1707 (N_1707,N_1512,N_1527);
or U1708 (N_1708,N_1455,N_1426);
xor U1709 (N_1709,N_1437,N_1496);
nand U1710 (N_1710,N_1414,N_1538);
nand U1711 (N_1711,N_1426,N_1425);
and U1712 (N_1712,N_1429,N_1599);
and U1713 (N_1713,N_1443,N_1539);
or U1714 (N_1714,N_1536,N_1474);
nand U1715 (N_1715,N_1514,N_1505);
xor U1716 (N_1716,N_1536,N_1529);
and U1717 (N_1717,N_1547,N_1446);
nand U1718 (N_1718,N_1453,N_1497);
and U1719 (N_1719,N_1438,N_1419);
and U1720 (N_1720,N_1457,N_1521);
nand U1721 (N_1721,N_1429,N_1443);
nand U1722 (N_1722,N_1568,N_1460);
nand U1723 (N_1723,N_1472,N_1400);
xor U1724 (N_1724,N_1406,N_1555);
nand U1725 (N_1725,N_1558,N_1491);
and U1726 (N_1726,N_1545,N_1442);
and U1727 (N_1727,N_1470,N_1433);
and U1728 (N_1728,N_1423,N_1443);
and U1729 (N_1729,N_1542,N_1490);
or U1730 (N_1730,N_1543,N_1439);
and U1731 (N_1731,N_1505,N_1534);
or U1732 (N_1732,N_1483,N_1591);
and U1733 (N_1733,N_1449,N_1580);
or U1734 (N_1734,N_1439,N_1517);
and U1735 (N_1735,N_1419,N_1598);
nand U1736 (N_1736,N_1477,N_1582);
xnor U1737 (N_1737,N_1471,N_1551);
nand U1738 (N_1738,N_1566,N_1423);
nand U1739 (N_1739,N_1454,N_1453);
nor U1740 (N_1740,N_1516,N_1502);
xor U1741 (N_1741,N_1478,N_1482);
and U1742 (N_1742,N_1527,N_1477);
nand U1743 (N_1743,N_1579,N_1523);
nand U1744 (N_1744,N_1539,N_1524);
or U1745 (N_1745,N_1401,N_1541);
and U1746 (N_1746,N_1531,N_1407);
nor U1747 (N_1747,N_1513,N_1568);
or U1748 (N_1748,N_1494,N_1452);
nand U1749 (N_1749,N_1523,N_1481);
or U1750 (N_1750,N_1544,N_1446);
xor U1751 (N_1751,N_1597,N_1506);
and U1752 (N_1752,N_1487,N_1471);
and U1753 (N_1753,N_1521,N_1403);
xor U1754 (N_1754,N_1519,N_1510);
or U1755 (N_1755,N_1500,N_1598);
nand U1756 (N_1756,N_1528,N_1533);
and U1757 (N_1757,N_1495,N_1451);
or U1758 (N_1758,N_1579,N_1582);
and U1759 (N_1759,N_1445,N_1498);
or U1760 (N_1760,N_1415,N_1596);
xor U1761 (N_1761,N_1518,N_1547);
nand U1762 (N_1762,N_1514,N_1595);
nor U1763 (N_1763,N_1419,N_1545);
xnor U1764 (N_1764,N_1423,N_1411);
nor U1765 (N_1765,N_1434,N_1520);
xor U1766 (N_1766,N_1525,N_1453);
nand U1767 (N_1767,N_1406,N_1530);
and U1768 (N_1768,N_1435,N_1404);
xor U1769 (N_1769,N_1582,N_1485);
and U1770 (N_1770,N_1435,N_1423);
or U1771 (N_1771,N_1568,N_1522);
and U1772 (N_1772,N_1496,N_1430);
and U1773 (N_1773,N_1570,N_1547);
or U1774 (N_1774,N_1415,N_1478);
and U1775 (N_1775,N_1405,N_1554);
nor U1776 (N_1776,N_1526,N_1494);
xnor U1777 (N_1777,N_1435,N_1460);
or U1778 (N_1778,N_1423,N_1544);
nor U1779 (N_1779,N_1575,N_1565);
xnor U1780 (N_1780,N_1491,N_1435);
or U1781 (N_1781,N_1538,N_1562);
or U1782 (N_1782,N_1565,N_1570);
xnor U1783 (N_1783,N_1486,N_1447);
xor U1784 (N_1784,N_1474,N_1535);
nor U1785 (N_1785,N_1412,N_1552);
and U1786 (N_1786,N_1402,N_1421);
and U1787 (N_1787,N_1583,N_1530);
nor U1788 (N_1788,N_1535,N_1487);
xor U1789 (N_1789,N_1448,N_1470);
and U1790 (N_1790,N_1577,N_1400);
nand U1791 (N_1791,N_1533,N_1423);
nand U1792 (N_1792,N_1591,N_1535);
nand U1793 (N_1793,N_1449,N_1441);
or U1794 (N_1794,N_1525,N_1500);
and U1795 (N_1795,N_1524,N_1519);
nor U1796 (N_1796,N_1536,N_1407);
nor U1797 (N_1797,N_1449,N_1406);
nor U1798 (N_1798,N_1482,N_1534);
or U1799 (N_1799,N_1515,N_1430);
xnor U1800 (N_1800,N_1731,N_1789);
nand U1801 (N_1801,N_1777,N_1654);
xor U1802 (N_1802,N_1771,N_1786);
xor U1803 (N_1803,N_1662,N_1724);
xor U1804 (N_1804,N_1708,N_1773);
nor U1805 (N_1805,N_1603,N_1756);
or U1806 (N_1806,N_1775,N_1764);
xor U1807 (N_1807,N_1798,N_1621);
or U1808 (N_1808,N_1784,N_1683);
xor U1809 (N_1809,N_1672,N_1655);
nor U1810 (N_1810,N_1645,N_1642);
nor U1811 (N_1811,N_1650,N_1766);
nand U1812 (N_1812,N_1791,N_1661);
or U1813 (N_1813,N_1622,N_1684);
nand U1814 (N_1814,N_1617,N_1620);
xor U1815 (N_1815,N_1692,N_1790);
xor U1816 (N_1816,N_1727,N_1643);
and U1817 (N_1817,N_1663,N_1640);
nand U1818 (N_1818,N_1744,N_1701);
or U1819 (N_1819,N_1671,N_1606);
nor U1820 (N_1820,N_1730,N_1610);
nand U1821 (N_1821,N_1689,N_1656);
and U1822 (N_1822,N_1675,N_1740);
xnor U1823 (N_1823,N_1633,N_1696);
or U1824 (N_1824,N_1720,N_1647);
nand U1825 (N_1825,N_1710,N_1649);
and U1826 (N_1826,N_1752,N_1693);
nor U1827 (N_1827,N_1750,N_1676);
or U1828 (N_1828,N_1611,N_1698);
or U1829 (N_1829,N_1729,N_1761);
and U1830 (N_1830,N_1711,N_1637);
or U1831 (N_1831,N_1670,N_1697);
xnor U1832 (N_1832,N_1631,N_1719);
xor U1833 (N_1833,N_1660,N_1691);
or U1834 (N_1834,N_1747,N_1601);
or U1835 (N_1835,N_1688,N_1749);
and U1836 (N_1836,N_1769,N_1703);
xor U1837 (N_1837,N_1799,N_1746);
xnor U1838 (N_1838,N_1751,N_1635);
nand U1839 (N_1839,N_1739,N_1795);
or U1840 (N_1840,N_1624,N_1627);
nand U1841 (N_1841,N_1623,N_1706);
nor U1842 (N_1842,N_1772,N_1794);
nand U1843 (N_1843,N_1788,N_1665);
and U1844 (N_1844,N_1629,N_1634);
and U1845 (N_1845,N_1709,N_1609);
nand U1846 (N_1846,N_1605,N_1664);
nor U1847 (N_1847,N_1613,N_1717);
and U1848 (N_1848,N_1741,N_1638);
xor U1849 (N_1849,N_1715,N_1785);
xnor U1850 (N_1850,N_1705,N_1658);
or U1851 (N_1851,N_1653,N_1699);
nor U1852 (N_1852,N_1694,N_1607);
nor U1853 (N_1853,N_1733,N_1742);
nor U1854 (N_1854,N_1625,N_1755);
nand U1855 (N_1855,N_1792,N_1734);
and U1856 (N_1856,N_1608,N_1753);
nand U1857 (N_1857,N_1781,N_1669);
nand U1858 (N_1858,N_1722,N_1736);
and U1859 (N_1859,N_1723,N_1757);
nor U1860 (N_1860,N_1651,N_1754);
or U1861 (N_1861,N_1721,N_1685);
or U1862 (N_1862,N_1695,N_1718);
or U1863 (N_1863,N_1712,N_1632);
xor U1864 (N_1864,N_1732,N_1686);
and U1865 (N_1865,N_1615,N_1687);
and U1866 (N_1866,N_1770,N_1780);
nor U1867 (N_1867,N_1614,N_1760);
xnor U1868 (N_1868,N_1707,N_1782);
nor U1869 (N_1869,N_1636,N_1767);
and U1870 (N_1870,N_1797,N_1716);
nor U1871 (N_1871,N_1762,N_1783);
and U1872 (N_1872,N_1677,N_1700);
nand U1873 (N_1873,N_1679,N_1674);
or U1874 (N_1874,N_1673,N_1793);
xnor U1875 (N_1875,N_1616,N_1659);
nand U1876 (N_1876,N_1678,N_1743);
nand U1877 (N_1877,N_1745,N_1612);
nand U1878 (N_1878,N_1704,N_1765);
xor U1879 (N_1879,N_1728,N_1667);
xor U1880 (N_1880,N_1618,N_1725);
nand U1881 (N_1881,N_1668,N_1652);
and U1882 (N_1882,N_1657,N_1644);
or U1883 (N_1883,N_1681,N_1630);
nand U1884 (N_1884,N_1759,N_1702);
and U1885 (N_1885,N_1639,N_1726);
xnor U1886 (N_1886,N_1768,N_1776);
and U1887 (N_1887,N_1628,N_1779);
or U1888 (N_1888,N_1682,N_1641);
nand U1889 (N_1889,N_1735,N_1774);
nor U1890 (N_1890,N_1758,N_1778);
or U1891 (N_1891,N_1666,N_1787);
and U1892 (N_1892,N_1748,N_1690);
nor U1893 (N_1893,N_1680,N_1737);
nor U1894 (N_1894,N_1626,N_1648);
and U1895 (N_1895,N_1763,N_1604);
nor U1896 (N_1896,N_1602,N_1646);
nand U1897 (N_1897,N_1796,N_1713);
xor U1898 (N_1898,N_1738,N_1600);
or U1899 (N_1899,N_1714,N_1619);
nor U1900 (N_1900,N_1731,N_1624);
nand U1901 (N_1901,N_1768,N_1608);
nor U1902 (N_1902,N_1638,N_1677);
or U1903 (N_1903,N_1704,N_1613);
and U1904 (N_1904,N_1796,N_1664);
nand U1905 (N_1905,N_1691,N_1668);
or U1906 (N_1906,N_1694,N_1798);
xor U1907 (N_1907,N_1764,N_1750);
nand U1908 (N_1908,N_1672,N_1696);
nor U1909 (N_1909,N_1710,N_1798);
nand U1910 (N_1910,N_1651,N_1730);
nor U1911 (N_1911,N_1616,N_1656);
nand U1912 (N_1912,N_1682,N_1743);
xnor U1913 (N_1913,N_1763,N_1617);
or U1914 (N_1914,N_1661,N_1685);
or U1915 (N_1915,N_1778,N_1773);
and U1916 (N_1916,N_1663,N_1692);
nand U1917 (N_1917,N_1764,N_1600);
or U1918 (N_1918,N_1784,N_1679);
nor U1919 (N_1919,N_1780,N_1610);
or U1920 (N_1920,N_1659,N_1709);
and U1921 (N_1921,N_1656,N_1600);
nor U1922 (N_1922,N_1766,N_1602);
or U1923 (N_1923,N_1792,N_1757);
and U1924 (N_1924,N_1625,N_1799);
and U1925 (N_1925,N_1704,N_1746);
xor U1926 (N_1926,N_1782,N_1748);
and U1927 (N_1927,N_1655,N_1601);
and U1928 (N_1928,N_1700,N_1734);
xnor U1929 (N_1929,N_1721,N_1683);
nor U1930 (N_1930,N_1614,N_1620);
nor U1931 (N_1931,N_1648,N_1658);
xor U1932 (N_1932,N_1632,N_1737);
xor U1933 (N_1933,N_1639,N_1745);
xor U1934 (N_1934,N_1758,N_1646);
or U1935 (N_1935,N_1738,N_1703);
nand U1936 (N_1936,N_1737,N_1657);
nand U1937 (N_1937,N_1648,N_1719);
or U1938 (N_1938,N_1725,N_1757);
or U1939 (N_1939,N_1741,N_1676);
nand U1940 (N_1940,N_1608,N_1680);
and U1941 (N_1941,N_1649,N_1767);
or U1942 (N_1942,N_1680,N_1670);
nor U1943 (N_1943,N_1666,N_1760);
nor U1944 (N_1944,N_1719,N_1703);
xor U1945 (N_1945,N_1608,N_1696);
nand U1946 (N_1946,N_1657,N_1658);
nand U1947 (N_1947,N_1672,N_1746);
nor U1948 (N_1948,N_1715,N_1732);
nor U1949 (N_1949,N_1708,N_1644);
or U1950 (N_1950,N_1683,N_1620);
and U1951 (N_1951,N_1672,N_1712);
and U1952 (N_1952,N_1748,N_1636);
xnor U1953 (N_1953,N_1720,N_1632);
xnor U1954 (N_1954,N_1666,N_1735);
xnor U1955 (N_1955,N_1677,N_1686);
xor U1956 (N_1956,N_1757,N_1795);
nor U1957 (N_1957,N_1785,N_1749);
or U1958 (N_1958,N_1679,N_1666);
nor U1959 (N_1959,N_1674,N_1658);
nand U1960 (N_1960,N_1798,N_1678);
or U1961 (N_1961,N_1658,N_1644);
nor U1962 (N_1962,N_1787,N_1639);
nor U1963 (N_1963,N_1606,N_1652);
or U1964 (N_1964,N_1745,N_1698);
nand U1965 (N_1965,N_1772,N_1773);
and U1966 (N_1966,N_1681,N_1770);
or U1967 (N_1967,N_1751,N_1690);
or U1968 (N_1968,N_1614,N_1638);
nand U1969 (N_1969,N_1608,N_1650);
xor U1970 (N_1970,N_1761,N_1623);
xor U1971 (N_1971,N_1726,N_1675);
nand U1972 (N_1972,N_1643,N_1758);
and U1973 (N_1973,N_1787,N_1741);
xnor U1974 (N_1974,N_1721,N_1617);
nand U1975 (N_1975,N_1620,N_1759);
or U1976 (N_1976,N_1773,N_1661);
nand U1977 (N_1977,N_1650,N_1697);
or U1978 (N_1978,N_1768,N_1695);
xnor U1979 (N_1979,N_1646,N_1665);
or U1980 (N_1980,N_1775,N_1667);
and U1981 (N_1981,N_1780,N_1603);
or U1982 (N_1982,N_1627,N_1620);
nand U1983 (N_1983,N_1695,N_1694);
nor U1984 (N_1984,N_1701,N_1620);
and U1985 (N_1985,N_1737,N_1774);
or U1986 (N_1986,N_1689,N_1741);
xnor U1987 (N_1987,N_1603,N_1651);
or U1988 (N_1988,N_1678,N_1625);
or U1989 (N_1989,N_1751,N_1732);
nor U1990 (N_1990,N_1699,N_1789);
nor U1991 (N_1991,N_1727,N_1699);
or U1992 (N_1992,N_1699,N_1600);
nor U1993 (N_1993,N_1601,N_1614);
xor U1994 (N_1994,N_1613,N_1719);
nand U1995 (N_1995,N_1782,N_1647);
nor U1996 (N_1996,N_1613,N_1755);
or U1997 (N_1997,N_1798,N_1728);
and U1998 (N_1998,N_1694,N_1654);
nor U1999 (N_1999,N_1741,N_1781);
nor U2000 (N_2000,N_1932,N_1848);
xnor U2001 (N_2001,N_1844,N_1805);
nand U2002 (N_2002,N_1900,N_1929);
nand U2003 (N_2003,N_1966,N_1999);
xnor U2004 (N_2004,N_1970,N_1987);
nand U2005 (N_2005,N_1813,N_1975);
xnor U2006 (N_2006,N_1845,N_1892);
and U2007 (N_2007,N_1919,N_1925);
or U2008 (N_2008,N_1901,N_1863);
nand U2009 (N_2009,N_1983,N_1902);
nand U2010 (N_2010,N_1853,N_1953);
xor U2011 (N_2011,N_1904,N_1864);
and U2012 (N_2012,N_1822,N_1920);
or U2013 (N_2013,N_1923,N_1930);
or U2014 (N_2014,N_1912,N_1982);
or U2015 (N_2015,N_1993,N_1927);
or U2016 (N_2016,N_1831,N_1801);
and U2017 (N_2017,N_1865,N_1833);
xnor U2018 (N_2018,N_1977,N_1886);
xor U2019 (N_2019,N_1937,N_1958);
xor U2020 (N_2020,N_1951,N_1944);
and U2021 (N_2021,N_1941,N_1911);
xnor U2022 (N_2022,N_1917,N_1811);
nand U2023 (N_2023,N_1849,N_1964);
and U2024 (N_2024,N_1942,N_1835);
xnor U2025 (N_2025,N_1820,N_1856);
xnor U2026 (N_2026,N_1979,N_1968);
or U2027 (N_2027,N_1910,N_1924);
xnor U2028 (N_2028,N_1928,N_1978);
nor U2029 (N_2029,N_1894,N_1877);
nand U2030 (N_2030,N_1803,N_1967);
and U2031 (N_2031,N_1880,N_1842);
nand U2032 (N_2032,N_1869,N_1893);
xnor U2033 (N_2033,N_1806,N_1949);
and U2034 (N_2034,N_1963,N_1934);
xor U2035 (N_2035,N_1837,N_1843);
nor U2036 (N_2036,N_1821,N_1800);
nand U2037 (N_2037,N_1818,N_1885);
nor U2038 (N_2038,N_1908,N_1828);
and U2039 (N_2039,N_1809,N_1956);
nor U2040 (N_2040,N_1829,N_1860);
nand U2041 (N_2041,N_1873,N_1935);
xor U2042 (N_2042,N_1945,N_1984);
xor U2043 (N_2043,N_1802,N_1887);
nand U2044 (N_2044,N_1827,N_1846);
and U2045 (N_2045,N_1915,N_1896);
xor U2046 (N_2046,N_1936,N_1895);
nor U2047 (N_2047,N_1868,N_1980);
or U2048 (N_2048,N_1916,N_1991);
nor U2049 (N_2049,N_1959,N_1807);
nand U2050 (N_2050,N_1965,N_1976);
nor U2051 (N_2051,N_1897,N_1832);
or U2052 (N_2052,N_1943,N_1998);
nand U2053 (N_2053,N_1955,N_1939);
or U2054 (N_2054,N_1876,N_1819);
nand U2055 (N_2055,N_1992,N_1899);
xnor U2056 (N_2056,N_1817,N_1898);
nand U2057 (N_2057,N_1862,N_1960);
and U2058 (N_2058,N_1883,N_1997);
nor U2059 (N_2059,N_1909,N_1855);
and U2060 (N_2060,N_1867,N_1950);
and U2061 (N_2061,N_1882,N_1861);
nor U2062 (N_2062,N_1812,N_1814);
nand U2063 (N_2063,N_1988,N_1884);
nand U2064 (N_2064,N_1931,N_1808);
and U2065 (N_2065,N_1952,N_1804);
nand U2066 (N_2066,N_1825,N_1826);
xnor U2067 (N_2067,N_1859,N_1954);
nand U2068 (N_2068,N_1836,N_1971);
and U2069 (N_2069,N_1858,N_1841);
and U2070 (N_2070,N_1995,N_1874);
xor U2071 (N_2071,N_1957,N_1926);
xor U2072 (N_2072,N_1921,N_1875);
xor U2073 (N_2073,N_1903,N_1889);
or U2074 (N_2074,N_1879,N_1852);
xor U2075 (N_2075,N_1823,N_1986);
nor U2076 (N_2076,N_1938,N_1871);
xor U2077 (N_2077,N_1946,N_1810);
nor U2078 (N_2078,N_1996,N_1854);
nor U2079 (N_2079,N_1840,N_1989);
and U2080 (N_2080,N_1839,N_1981);
nand U2081 (N_2081,N_1985,N_1857);
nand U2082 (N_2082,N_1913,N_1947);
and U2083 (N_2083,N_1922,N_1890);
and U2084 (N_2084,N_1830,N_1851);
nor U2085 (N_2085,N_1948,N_1834);
or U2086 (N_2086,N_1961,N_1870);
nand U2087 (N_2087,N_1838,N_1850);
nor U2088 (N_2088,N_1891,N_1969);
and U2089 (N_2089,N_1905,N_1907);
nor U2090 (N_2090,N_1973,N_1914);
and U2091 (N_2091,N_1878,N_1962);
xnor U2092 (N_2092,N_1866,N_1918);
nor U2093 (N_2093,N_1994,N_1974);
or U2094 (N_2094,N_1906,N_1847);
nor U2095 (N_2095,N_1824,N_1816);
and U2096 (N_2096,N_1872,N_1972);
xnor U2097 (N_2097,N_1815,N_1888);
xor U2098 (N_2098,N_1990,N_1933);
or U2099 (N_2099,N_1940,N_1881);
or U2100 (N_2100,N_1976,N_1859);
xor U2101 (N_2101,N_1965,N_1989);
nor U2102 (N_2102,N_1979,N_1958);
nor U2103 (N_2103,N_1843,N_1903);
and U2104 (N_2104,N_1990,N_1949);
nand U2105 (N_2105,N_1998,N_1924);
xnor U2106 (N_2106,N_1913,N_1907);
and U2107 (N_2107,N_1974,N_1902);
or U2108 (N_2108,N_1978,N_1879);
xnor U2109 (N_2109,N_1995,N_1878);
nor U2110 (N_2110,N_1990,N_1889);
xor U2111 (N_2111,N_1838,N_1871);
xor U2112 (N_2112,N_1986,N_1909);
nand U2113 (N_2113,N_1894,N_1851);
nor U2114 (N_2114,N_1818,N_1914);
or U2115 (N_2115,N_1901,N_1904);
nand U2116 (N_2116,N_1944,N_1969);
nand U2117 (N_2117,N_1945,N_1813);
nor U2118 (N_2118,N_1813,N_1908);
or U2119 (N_2119,N_1946,N_1877);
and U2120 (N_2120,N_1845,N_1846);
xnor U2121 (N_2121,N_1865,N_1845);
xnor U2122 (N_2122,N_1900,N_1855);
nand U2123 (N_2123,N_1953,N_1899);
and U2124 (N_2124,N_1812,N_1852);
nand U2125 (N_2125,N_1948,N_1928);
and U2126 (N_2126,N_1897,N_1942);
nor U2127 (N_2127,N_1957,N_1857);
or U2128 (N_2128,N_1810,N_1828);
or U2129 (N_2129,N_1827,N_1950);
nor U2130 (N_2130,N_1943,N_1846);
nand U2131 (N_2131,N_1923,N_1906);
nor U2132 (N_2132,N_1870,N_1968);
nor U2133 (N_2133,N_1967,N_1843);
xnor U2134 (N_2134,N_1942,N_1857);
nand U2135 (N_2135,N_1980,N_1957);
and U2136 (N_2136,N_1954,N_1835);
xor U2137 (N_2137,N_1992,N_1852);
and U2138 (N_2138,N_1996,N_1928);
nand U2139 (N_2139,N_1804,N_1810);
or U2140 (N_2140,N_1947,N_1826);
or U2141 (N_2141,N_1865,N_1891);
and U2142 (N_2142,N_1877,N_1830);
nand U2143 (N_2143,N_1987,N_1870);
nand U2144 (N_2144,N_1939,N_1848);
xor U2145 (N_2145,N_1936,N_1913);
and U2146 (N_2146,N_1883,N_1838);
xnor U2147 (N_2147,N_1880,N_1966);
nand U2148 (N_2148,N_1992,N_1942);
nor U2149 (N_2149,N_1849,N_1814);
xnor U2150 (N_2150,N_1950,N_1801);
or U2151 (N_2151,N_1978,N_1905);
nand U2152 (N_2152,N_1917,N_1800);
and U2153 (N_2153,N_1935,N_1897);
nor U2154 (N_2154,N_1910,N_1859);
and U2155 (N_2155,N_1966,N_1948);
and U2156 (N_2156,N_1902,N_1907);
or U2157 (N_2157,N_1803,N_1865);
nor U2158 (N_2158,N_1806,N_1821);
or U2159 (N_2159,N_1834,N_1836);
xor U2160 (N_2160,N_1958,N_1947);
xnor U2161 (N_2161,N_1907,N_1838);
and U2162 (N_2162,N_1848,N_1871);
and U2163 (N_2163,N_1834,N_1835);
xnor U2164 (N_2164,N_1854,N_1891);
xor U2165 (N_2165,N_1952,N_1831);
nor U2166 (N_2166,N_1941,N_1976);
nand U2167 (N_2167,N_1884,N_1847);
or U2168 (N_2168,N_1971,N_1921);
xor U2169 (N_2169,N_1811,N_1907);
nand U2170 (N_2170,N_1824,N_1909);
or U2171 (N_2171,N_1947,N_1888);
nand U2172 (N_2172,N_1994,N_1858);
or U2173 (N_2173,N_1919,N_1818);
nand U2174 (N_2174,N_1854,N_1983);
and U2175 (N_2175,N_1998,N_1954);
xor U2176 (N_2176,N_1896,N_1891);
and U2177 (N_2177,N_1923,N_1937);
or U2178 (N_2178,N_1929,N_1845);
nand U2179 (N_2179,N_1961,N_1902);
or U2180 (N_2180,N_1975,N_1880);
nand U2181 (N_2181,N_1823,N_1852);
or U2182 (N_2182,N_1984,N_1843);
xor U2183 (N_2183,N_1820,N_1989);
or U2184 (N_2184,N_1936,N_1867);
nor U2185 (N_2185,N_1998,N_1827);
or U2186 (N_2186,N_1943,N_1811);
nand U2187 (N_2187,N_1959,N_1889);
nand U2188 (N_2188,N_1807,N_1927);
xnor U2189 (N_2189,N_1855,N_1901);
xnor U2190 (N_2190,N_1803,N_1811);
and U2191 (N_2191,N_1967,N_1804);
or U2192 (N_2192,N_1958,N_1989);
and U2193 (N_2193,N_1891,N_1824);
nor U2194 (N_2194,N_1867,N_1937);
nor U2195 (N_2195,N_1831,N_1998);
or U2196 (N_2196,N_1908,N_1866);
nor U2197 (N_2197,N_1869,N_1846);
or U2198 (N_2198,N_1871,N_1862);
nand U2199 (N_2199,N_1813,N_1886);
nand U2200 (N_2200,N_2086,N_2081);
and U2201 (N_2201,N_2059,N_2052);
or U2202 (N_2202,N_2179,N_2113);
and U2203 (N_2203,N_2132,N_2026);
or U2204 (N_2204,N_2105,N_2054);
xor U2205 (N_2205,N_2111,N_2031);
nor U2206 (N_2206,N_2048,N_2047);
or U2207 (N_2207,N_2187,N_2013);
xnor U2208 (N_2208,N_2064,N_2112);
nand U2209 (N_2209,N_2123,N_2055);
nor U2210 (N_2210,N_2174,N_2165);
or U2211 (N_2211,N_2139,N_2195);
nor U2212 (N_2212,N_2029,N_2061);
nand U2213 (N_2213,N_2040,N_2087);
and U2214 (N_2214,N_2003,N_2154);
or U2215 (N_2215,N_2056,N_2143);
xnor U2216 (N_2216,N_2152,N_2067);
or U2217 (N_2217,N_2011,N_2097);
nor U2218 (N_2218,N_2118,N_2109);
and U2219 (N_2219,N_2153,N_2126);
or U2220 (N_2220,N_2119,N_2102);
and U2221 (N_2221,N_2150,N_2070);
or U2222 (N_2222,N_2117,N_2182);
and U2223 (N_2223,N_2190,N_2115);
or U2224 (N_2224,N_2001,N_2095);
xnor U2225 (N_2225,N_2155,N_2122);
and U2226 (N_2226,N_2058,N_2138);
and U2227 (N_2227,N_2027,N_2144);
or U2228 (N_2228,N_2193,N_2076);
nand U2229 (N_2229,N_2014,N_2158);
nand U2230 (N_2230,N_2141,N_2010);
nor U2231 (N_2231,N_2006,N_2044);
and U2232 (N_2232,N_2041,N_2098);
or U2233 (N_2233,N_2110,N_2194);
and U2234 (N_2234,N_2114,N_2017);
or U2235 (N_2235,N_2121,N_2125);
nand U2236 (N_2236,N_2180,N_2039);
or U2237 (N_2237,N_2079,N_2140);
xor U2238 (N_2238,N_2106,N_2162);
xnor U2239 (N_2239,N_2103,N_2129);
nor U2240 (N_2240,N_2068,N_2025);
nor U2241 (N_2241,N_2099,N_2100);
nand U2242 (N_2242,N_2151,N_2020);
or U2243 (N_2243,N_2177,N_2074);
or U2244 (N_2244,N_2065,N_2082);
xor U2245 (N_2245,N_2198,N_2080);
and U2246 (N_2246,N_2015,N_2042);
nor U2247 (N_2247,N_2089,N_2127);
and U2248 (N_2248,N_2168,N_2175);
xor U2249 (N_2249,N_2009,N_2033);
and U2250 (N_2250,N_2134,N_2057);
nand U2251 (N_2251,N_2131,N_2021);
nor U2252 (N_2252,N_2156,N_2050);
nor U2253 (N_2253,N_2077,N_2191);
nand U2254 (N_2254,N_2000,N_2008);
or U2255 (N_2255,N_2172,N_2049);
xor U2256 (N_2256,N_2116,N_2024);
nand U2257 (N_2257,N_2171,N_2069);
nor U2258 (N_2258,N_2004,N_2007);
or U2259 (N_2259,N_2090,N_2018);
and U2260 (N_2260,N_2169,N_2071);
xor U2261 (N_2261,N_2032,N_2088);
nor U2262 (N_2262,N_2034,N_2160);
nand U2263 (N_2263,N_2188,N_2043);
nor U2264 (N_2264,N_2146,N_2045);
or U2265 (N_2265,N_2094,N_2128);
nand U2266 (N_2266,N_2159,N_2136);
and U2267 (N_2267,N_2030,N_2176);
xnor U2268 (N_2268,N_2173,N_2016);
nand U2269 (N_2269,N_2022,N_2178);
nor U2270 (N_2270,N_2051,N_2183);
and U2271 (N_2271,N_2037,N_2192);
nand U2272 (N_2272,N_2093,N_2101);
and U2273 (N_2273,N_2142,N_2107);
xnor U2274 (N_2274,N_2167,N_2038);
xnor U2275 (N_2275,N_2072,N_2157);
and U2276 (N_2276,N_2137,N_2197);
xor U2277 (N_2277,N_2028,N_2066);
and U2278 (N_2278,N_2083,N_2170);
and U2279 (N_2279,N_2005,N_2163);
nor U2280 (N_2280,N_2185,N_2145);
xnor U2281 (N_2281,N_2196,N_2108);
and U2282 (N_2282,N_2053,N_2075);
xor U2283 (N_2283,N_2085,N_2060);
nor U2284 (N_2284,N_2164,N_2130);
and U2285 (N_2285,N_2161,N_2073);
nand U2286 (N_2286,N_2135,N_2002);
and U2287 (N_2287,N_2084,N_2184);
or U2288 (N_2288,N_2035,N_2078);
or U2289 (N_2289,N_2104,N_2124);
or U2290 (N_2290,N_2019,N_2046);
or U2291 (N_2291,N_2096,N_2091);
or U2292 (N_2292,N_2023,N_2036);
xnor U2293 (N_2293,N_2063,N_2062);
nor U2294 (N_2294,N_2186,N_2147);
and U2295 (N_2295,N_2149,N_2092);
or U2296 (N_2296,N_2181,N_2189);
nor U2297 (N_2297,N_2133,N_2166);
nor U2298 (N_2298,N_2120,N_2148);
and U2299 (N_2299,N_2199,N_2012);
xnor U2300 (N_2300,N_2150,N_2074);
xnor U2301 (N_2301,N_2133,N_2008);
or U2302 (N_2302,N_2184,N_2049);
or U2303 (N_2303,N_2143,N_2198);
and U2304 (N_2304,N_2134,N_2171);
nor U2305 (N_2305,N_2009,N_2173);
xnor U2306 (N_2306,N_2126,N_2147);
or U2307 (N_2307,N_2162,N_2058);
or U2308 (N_2308,N_2116,N_2066);
nand U2309 (N_2309,N_2021,N_2064);
xnor U2310 (N_2310,N_2104,N_2108);
xnor U2311 (N_2311,N_2182,N_2069);
nand U2312 (N_2312,N_2093,N_2194);
xor U2313 (N_2313,N_2122,N_2124);
and U2314 (N_2314,N_2015,N_2018);
xor U2315 (N_2315,N_2026,N_2015);
and U2316 (N_2316,N_2057,N_2128);
or U2317 (N_2317,N_2170,N_2072);
nand U2318 (N_2318,N_2069,N_2149);
or U2319 (N_2319,N_2131,N_2168);
nand U2320 (N_2320,N_2078,N_2020);
nor U2321 (N_2321,N_2128,N_2070);
xor U2322 (N_2322,N_2085,N_2001);
nor U2323 (N_2323,N_2128,N_2025);
or U2324 (N_2324,N_2032,N_2147);
or U2325 (N_2325,N_2097,N_2147);
xor U2326 (N_2326,N_2180,N_2018);
xnor U2327 (N_2327,N_2185,N_2011);
xnor U2328 (N_2328,N_2123,N_2192);
nand U2329 (N_2329,N_2105,N_2063);
or U2330 (N_2330,N_2006,N_2171);
or U2331 (N_2331,N_2146,N_2068);
nand U2332 (N_2332,N_2019,N_2129);
or U2333 (N_2333,N_2170,N_2025);
and U2334 (N_2334,N_2017,N_2101);
xor U2335 (N_2335,N_2001,N_2124);
and U2336 (N_2336,N_2024,N_2011);
nand U2337 (N_2337,N_2196,N_2023);
and U2338 (N_2338,N_2093,N_2164);
nand U2339 (N_2339,N_2056,N_2133);
xor U2340 (N_2340,N_2131,N_2101);
nor U2341 (N_2341,N_2074,N_2016);
or U2342 (N_2342,N_2196,N_2075);
nand U2343 (N_2343,N_2167,N_2069);
nand U2344 (N_2344,N_2164,N_2187);
and U2345 (N_2345,N_2011,N_2160);
and U2346 (N_2346,N_2090,N_2123);
or U2347 (N_2347,N_2170,N_2111);
and U2348 (N_2348,N_2056,N_2029);
nor U2349 (N_2349,N_2040,N_2136);
and U2350 (N_2350,N_2120,N_2026);
nand U2351 (N_2351,N_2112,N_2082);
and U2352 (N_2352,N_2116,N_2067);
xor U2353 (N_2353,N_2076,N_2006);
and U2354 (N_2354,N_2134,N_2074);
and U2355 (N_2355,N_2134,N_2005);
or U2356 (N_2356,N_2177,N_2022);
and U2357 (N_2357,N_2013,N_2115);
or U2358 (N_2358,N_2165,N_2172);
xnor U2359 (N_2359,N_2197,N_2057);
nor U2360 (N_2360,N_2116,N_2168);
nor U2361 (N_2361,N_2189,N_2022);
nor U2362 (N_2362,N_2060,N_2072);
xnor U2363 (N_2363,N_2039,N_2197);
and U2364 (N_2364,N_2152,N_2117);
or U2365 (N_2365,N_2106,N_2085);
and U2366 (N_2366,N_2085,N_2027);
xor U2367 (N_2367,N_2125,N_2046);
xnor U2368 (N_2368,N_2194,N_2188);
or U2369 (N_2369,N_2084,N_2187);
xor U2370 (N_2370,N_2033,N_2067);
nor U2371 (N_2371,N_2093,N_2065);
and U2372 (N_2372,N_2063,N_2190);
or U2373 (N_2373,N_2122,N_2071);
and U2374 (N_2374,N_2022,N_2024);
or U2375 (N_2375,N_2185,N_2199);
and U2376 (N_2376,N_2055,N_2042);
or U2377 (N_2377,N_2124,N_2074);
and U2378 (N_2378,N_2028,N_2151);
or U2379 (N_2379,N_2006,N_2086);
or U2380 (N_2380,N_2109,N_2170);
xor U2381 (N_2381,N_2012,N_2120);
or U2382 (N_2382,N_2150,N_2122);
xnor U2383 (N_2383,N_2123,N_2158);
or U2384 (N_2384,N_2048,N_2189);
or U2385 (N_2385,N_2167,N_2107);
or U2386 (N_2386,N_2004,N_2069);
nor U2387 (N_2387,N_2038,N_2180);
xor U2388 (N_2388,N_2057,N_2100);
or U2389 (N_2389,N_2074,N_2161);
nand U2390 (N_2390,N_2086,N_2119);
xnor U2391 (N_2391,N_2050,N_2199);
or U2392 (N_2392,N_2038,N_2033);
or U2393 (N_2393,N_2168,N_2185);
and U2394 (N_2394,N_2120,N_2168);
nand U2395 (N_2395,N_2192,N_2097);
or U2396 (N_2396,N_2194,N_2197);
nor U2397 (N_2397,N_2040,N_2036);
or U2398 (N_2398,N_2111,N_2090);
and U2399 (N_2399,N_2172,N_2181);
nor U2400 (N_2400,N_2274,N_2302);
nor U2401 (N_2401,N_2356,N_2204);
nor U2402 (N_2402,N_2376,N_2290);
nand U2403 (N_2403,N_2317,N_2222);
nand U2404 (N_2404,N_2381,N_2280);
nor U2405 (N_2405,N_2293,N_2201);
and U2406 (N_2406,N_2285,N_2216);
nand U2407 (N_2407,N_2227,N_2343);
nor U2408 (N_2408,N_2257,N_2329);
nor U2409 (N_2409,N_2273,N_2221);
xnor U2410 (N_2410,N_2377,N_2292);
nor U2411 (N_2411,N_2339,N_2265);
nor U2412 (N_2412,N_2388,N_2312);
and U2413 (N_2413,N_2384,N_2373);
or U2414 (N_2414,N_2305,N_2300);
or U2415 (N_2415,N_2287,N_2237);
nand U2416 (N_2416,N_2207,N_2225);
nand U2417 (N_2417,N_2360,N_2203);
and U2418 (N_2418,N_2233,N_2387);
xor U2419 (N_2419,N_2232,N_2246);
nor U2420 (N_2420,N_2276,N_2362);
or U2421 (N_2421,N_2235,N_2341);
and U2422 (N_2422,N_2398,N_2311);
and U2423 (N_2423,N_2294,N_2289);
and U2424 (N_2424,N_2330,N_2219);
nor U2425 (N_2425,N_2368,N_2314);
xnor U2426 (N_2426,N_2351,N_2363);
and U2427 (N_2427,N_2318,N_2392);
xor U2428 (N_2428,N_2217,N_2279);
and U2429 (N_2429,N_2323,N_2327);
xor U2430 (N_2430,N_2261,N_2281);
or U2431 (N_2431,N_2324,N_2245);
or U2432 (N_2432,N_2242,N_2220);
or U2433 (N_2433,N_2282,N_2306);
nor U2434 (N_2434,N_2364,N_2239);
and U2435 (N_2435,N_2256,N_2248);
and U2436 (N_2436,N_2338,N_2218);
and U2437 (N_2437,N_2321,N_2355);
xnor U2438 (N_2438,N_2230,N_2291);
nand U2439 (N_2439,N_2288,N_2320);
nand U2440 (N_2440,N_2263,N_2268);
xnor U2441 (N_2441,N_2319,N_2266);
xnor U2442 (N_2442,N_2301,N_2352);
nand U2443 (N_2443,N_2342,N_2325);
nor U2444 (N_2444,N_2208,N_2213);
or U2445 (N_2445,N_2357,N_2332);
nand U2446 (N_2446,N_2365,N_2366);
or U2447 (N_2447,N_2299,N_2370);
xor U2448 (N_2448,N_2262,N_2315);
and U2449 (N_2449,N_2260,N_2395);
nand U2450 (N_2450,N_2389,N_2359);
and U2451 (N_2451,N_2250,N_2354);
and U2452 (N_2452,N_2283,N_2252);
nand U2453 (N_2453,N_2361,N_2234);
or U2454 (N_2454,N_2303,N_2277);
or U2455 (N_2455,N_2310,N_2214);
and U2456 (N_2456,N_2334,N_2378);
xor U2457 (N_2457,N_2307,N_2372);
nand U2458 (N_2458,N_2226,N_2215);
nand U2459 (N_2459,N_2333,N_2238);
and U2460 (N_2460,N_2313,N_2296);
nor U2461 (N_2461,N_2336,N_2347);
and U2462 (N_2462,N_2251,N_2259);
nand U2463 (N_2463,N_2371,N_2316);
and U2464 (N_2464,N_2249,N_2255);
nor U2465 (N_2465,N_2247,N_2390);
or U2466 (N_2466,N_2397,N_2304);
and U2467 (N_2467,N_2209,N_2298);
and U2468 (N_2468,N_2326,N_2345);
nor U2469 (N_2469,N_2241,N_2382);
nor U2470 (N_2470,N_2267,N_2297);
and U2471 (N_2471,N_2353,N_2258);
and U2472 (N_2472,N_2391,N_2358);
and U2473 (N_2473,N_2200,N_2253);
xor U2474 (N_2474,N_2272,N_2224);
or U2475 (N_2475,N_2206,N_2205);
xnor U2476 (N_2476,N_2284,N_2394);
or U2477 (N_2477,N_2308,N_2335);
and U2478 (N_2478,N_2270,N_2337);
nand U2479 (N_2479,N_2240,N_2367);
xnor U2480 (N_2480,N_2322,N_2295);
nand U2481 (N_2481,N_2379,N_2211);
nor U2482 (N_2482,N_2286,N_2340);
and U2483 (N_2483,N_2244,N_2228);
nand U2484 (N_2484,N_2396,N_2271);
or U2485 (N_2485,N_2385,N_2383);
xnor U2486 (N_2486,N_2348,N_2386);
nor U2487 (N_2487,N_2243,N_2264);
xor U2488 (N_2488,N_2374,N_2212);
nor U2489 (N_2489,N_2210,N_2393);
or U2490 (N_2490,N_2229,N_2369);
nor U2491 (N_2491,N_2346,N_2309);
and U2492 (N_2492,N_2349,N_2350);
and U2493 (N_2493,N_2380,N_2328);
nand U2494 (N_2494,N_2275,N_2331);
nand U2495 (N_2495,N_2254,N_2231);
nor U2496 (N_2496,N_2236,N_2202);
nand U2497 (N_2497,N_2278,N_2223);
nand U2498 (N_2498,N_2269,N_2344);
nand U2499 (N_2499,N_2399,N_2375);
nand U2500 (N_2500,N_2206,N_2362);
nand U2501 (N_2501,N_2272,N_2214);
nand U2502 (N_2502,N_2396,N_2368);
or U2503 (N_2503,N_2255,N_2301);
nor U2504 (N_2504,N_2224,N_2316);
or U2505 (N_2505,N_2294,N_2238);
nand U2506 (N_2506,N_2255,N_2209);
xnor U2507 (N_2507,N_2283,N_2348);
xor U2508 (N_2508,N_2324,N_2264);
nand U2509 (N_2509,N_2276,N_2242);
nor U2510 (N_2510,N_2360,N_2343);
or U2511 (N_2511,N_2294,N_2242);
nor U2512 (N_2512,N_2382,N_2254);
xnor U2513 (N_2513,N_2394,N_2214);
and U2514 (N_2514,N_2360,N_2370);
xor U2515 (N_2515,N_2289,N_2362);
and U2516 (N_2516,N_2334,N_2396);
nor U2517 (N_2517,N_2263,N_2277);
nand U2518 (N_2518,N_2346,N_2383);
and U2519 (N_2519,N_2320,N_2340);
nand U2520 (N_2520,N_2356,N_2243);
nand U2521 (N_2521,N_2344,N_2310);
or U2522 (N_2522,N_2286,N_2374);
and U2523 (N_2523,N_2248,N_2211);
nor U2524 (N_2524,N_2214,N_2368);
nand U2525 (N_2525,N_2338,N_2221);
or U2526 (N_2526,N_2336,N_2225);
nand U2527 (N_2527,N_2313,N_2311);
nand U2528 (N_2528,N_2207,N_2227);
or U2529 (N_2529,N_2353,N_2321);
nand U2530 (N_2530,N_2379,N_2327);
and U2531 (N_2531,N_2395,N_2261);
and U2532 (N_2532,N_2300,N_2363);
nand U2533 (N_2533,N_2208,N_2232);
nand U2534 (N_2534,N_2236,N_2395);
xnor U2535 (N_2535,N_2263,N_2247);
xnor U2536 (N_2536,N_2399,N_2303);
nand U2537 (N_2537,N_2226,N_2353);
or U2538 (N_2538,N_2221,N_2362);
xor U2539 (N_2539,N_2272,N_2274);
nor U2540 (N_2540,N_2205,N_2360);
nor U2541 (N_2541,N_2376,N_2328);
and U2542 (N_2542,N_2362,N_2234);
nor U2543 (N_2543,N_2226,N_2235);
nor U2544 (N_2544,N_2282,N_2366);
xor U2545 (N_2545,N_2394,N_2368);
xor U2546 (N_2546,N_2302,N_2286);
nor U2547 (N_2547,N_2261,N_2262);
or U2548 (N_2548,N_2254,N_2233);
or U2549 (N_2549,N_2267,N_2273);
nand U2550 (N_2550,N_2282,N_2201);
xnor U2551 (N_2551,N_2242,N_2336);
nor U2552 (N_2552,N_2389,N_2387);
nand U2553 (N_2553,N_2220,N_2372);
nand U2554 (N_2554,N_2364,N_2283);
nand U2555 (N_2555,N_2363,N_2308);
nor U2556 (N_2556,N_2276,N_2325);
nor U2557 (N_2557,N_2217,N_2204);
nor U2558 (N_2558,N_2374,N_2232);
xor U2559 (N_2559,N_2391,N_2300);
xor U2560 (N_2560,N_2219,N_2251);
and U2561 (N_2561,N_2305,N_2297);
nor U2562 (N_2562,N_2341,N_2259);
nor U2563 (N_2563,N_2348,N_2249);
or U2564 (N_2564,N_2219,N_2331);
or U2565 (N_2565,N_2225,N_2214);
nand U2566 (N_2566,N_2294,N_2333);
or U2567 (N_2567,N_2312,N_2330);
or U2568 (N_2568,N_2376,N_2395);
nand U2569 (N_2569,N_2219,N_2335);
nor U2570 (N_2570,N_2293,N_2387);
or U2571 (N_2571,N_2314,N_2290);
nand U2572 (N_2572,N_2290,N_2303);
nor U2573 (N_2573,N_2287,N_2231);
nor U2574 (N_2574,N_2200,N_2339);
xor U2575 (N_2575,N_2346,N_2395);
or U2576 (N_2576,N_2211,N_2352);
or U2577 (N_2577,N_2371,N_2225);
xor U2578 (N_2578,N_2325,N_2327);
nor U2579 (N_2579,N_2295,N_2384);
or U2580 (N_2580,N_2281,N_2202);
and U2581 (N_2581,N_2244,N_2249);
xnor U2582 (N_2582,N_2266,N_2309);
and U2583 (N_2583,N_2303,N_2229);
nand U2584 (N_2584,N_2203,N_2258);
and U2585 (N_2585,N_2215,N_2286);
and U2586 (N_2586,N_2289,N_2361);
xor U2587 (N_2587,N_2230,N_2278);
xor U2588 (N_2588,N_2284,N_2298);
and U2589 (N_2589,N_2371,N_2385);
and U2590 (N_2590,N_2218,N_2372);
or U2591 (N_2591,N_2273,N_2389);
or U2592 (N_2592,N_2381,N_2243);
or U2593 (N_2593,N_2287,N_2374);
xnor U2594 (N_2594,N_2394,N_2213);
nand U2595 (N_2595,N_2250,N_2263);
nor U2596 (N_2596,N_2214,N_2349);
nand U2597 (N_2597,N_2348,N_2262);
nand U2598 (N_2598,N_2229,N_2373);
and U2599 (N_2599,N_2305,N_2232);
and U2600 (N_2600,N_2453,N_2560);
xor U2601 (N_2601,N_2414,N_2462);
or U2602 (N_2602,N_2484,N_2490);
and U2603 (N_2603,N_2538,N_2501);
nand U2604 (N_2604,N_2423,N_2421);
and U2605 (N_2605,N_2449,N_2563);
and U2606 (N_2606,N_2406,N_2474);
and U2607 (N_2607,N_2596,N_2509);
and U2608 (N_2608,N_2562,N_2457);
or U2609 (N_2609,N_2524,N_2499);
and U2610 (N_2610,N_2544,N_2419);
xnor U2611 (N_2611,N_2520,N_2577);
and U2612 (N_2612,N_2543,N_2554);
xnor U2613 (N_2613,N_2489,N_2441);
and U2614 (N_2614,N_2506,N_2442);
and U2615 (N_2615,N_2545,N_2440);
or U2616 (N_2616,N_2576,N_2472);
xor U2617 (N_2617,N_2519,N_2460);
nand U2618 (N_2618,N_2542,N_2429);
nand U2619 (N_2619,N_2592,N_2425);
nor U2620 (N_2620,N_2480,N_2424);
or U2621 (N_2621,N_2412,N_2467);
or U2622 (N_2622,N_2475,N_2485);
nor U2623 (N_2623,N_2468,N_2402);
xnor U2624 (N_2624,N_2535,N_2452);
nor U2625 (N_2625,N_2479,N_2586);
xor U2626 (N_2626,N_2444,N_2428);
or U2627 (N_2627,N_2583,N_2436);
nor U2628 (N_2628,N_2439,N_2558);
xor U2629 (N_2629,N_2529,N_2450);
xor U2630 (N_2630,N_2448,N_2420);
xor U2631 (N_2631,N_2486,N_2415);
nor U2632 (N_2632,N_2456,N_2500);
xor U2633 (N_2633,N_2568,N_2553);
or U2634 (N_2634,N_2401,N_2571);
xor U2635 (N_2635,N_2505,N_2591);
xor U2636 (N_2636,N_2559,N_2422);
and U2637 (N_2637,N_2516,N_2471);
xor U2638 (N_2638,N_2585,N_2557);
and U2639 (N_2639,N_2455,N_2464);
nor U2640 (N_2640,N_2527,N_2407);
nand U2641 (N_2641,N_2416,N_2589);
nor U2642 (N_2642,N_2426,N_2552);
xor U2643 (N_2643,N_2496,N_2555);
or U2644 (N_2644,N_2598,N_2463);
and U2645 (N_2645,N_2447,N_2532);
or U2646 (N_2646,N_2581,N_2473);
nand U2647 (N_2647,N_2478,N_2564);
nand U2648 (N_2648,N_2408,N_2570);
xnor U2649 (N_2649,N_2430,N_2572);
or U2650 (N_2650,N_2493,N_2481);
or U2651 (N_2651,N_2411,N_2461);
or U2652 (N_2652,N_2502,N_2561);
nand U2653 (N_2653,N_2512,N_2491);
xnor U2654 (N_2654,N_2587,N_2522);
xor U2655 (N_2655,N_2579,N_2497);
nor U2656 (N_2656,N_2580,N_2599);
nor U2657 (N_2657,N_2418,N_2569);
nor U2658 (N_2658,N_2488,N_2518);
and U2659 (N_2659,N_2417,N_2515);
and U2660 (N_2660,N_2517,N_2409);
nor U2661 (N_2661,N_2556,N_2458);
or U2662 (N_2662,N_2437,N_2593);
xnor U2663 (N_2663,N_2400,N_2597);
xnor U2664 (N_2664,N_2483,N_2494);
or U2665 (N_2665,N_2413,N_2405);
xnor U2666 (N_2666,N_2547,N_2536);
xor U2667 (N_2667,N_2525,N_2504);
and U2668 (N_2668,N_2438,N_2445);
nand U2669 (N_2669,N_2548,N_2528);
nand U2670 (N_2670,N_2521,N_2451);
nand U2671 (N_2671,N_2541,N_2503);
nand U2672 (N_2672,N_2495,N_2530);
nand U2673 (N_2673,N_2523,N_2550);
or U2674 (N_2674,N_2574,N_2573);
nor U2675 (N_2675,N_2578,N_2537);
nand U2676 (N_2676,N_2469,N_2477);
xnor U2677 (N_2677,N_2531,N_2540);
and U2678 (N_2678,N_2443,N_2526);
nor U2679 (N_2679,N_2487,N_2410);
nor U2680 (N_2680,N_2434,N_2565);
nand U2681 (N_2681,N_2575,N_2466);
and U2682 (N_2682,N_2594,N_2546);
xnor U2683 (N_2683,N_2539,N_2482);
xnor U2684 (N_2684,N_2492,N_2590);
and U2685 (N_2685,N_2508,N_2534);
nor U2686 (N_2686,N_2567,N_2403);
nand U2687 (N_2687,N_2566,N_2432);
nand U2688 (N_2688,N_2476,N_2507);
nor U2689 (N_2689,N_2454,N_2584);
nor U2690 (N_2690,N_2595,N_2551);
xnor U2691 (N_2691,N_2514,N_2435);
nand U2692 (N_2692,N_2465,N_2588);
nand U2693 (N_2693,N_2459,N_2446);
or U2694 (N_2694,N_2533,N_2431);
xnor U2695 (N_2695,N_2510,N_2511);
xor U2696 (N_2696,N_2498,N_2470);
xor U2697 (N_2697,N_2404,N_2433);
or U2698 (N_2698,N_2549,N_2427);
or U2699 (N_2699,N_2513,N_2582);
and U2700 (N_2700,N_2482,N_2556);
xnor U2701 (N_2701,N_2409,N_2586);
and U2702 (N_2702,N_2453,N_2557);
xnor U2703 (N_2703,N_2455,N_2582);
nand U2704 (N_2704,N_2553,N_2595);
or U2705 (N_2705,N_2588,N_2418);
xor U2706 (N_2706,N_2462,N_2514);
and U2707 (N_2707,N_2440,N_2563);
or U2708 (N_2708,N_2543,N_2470);
nand U2709 (N_2709,N_2583,N_2479);
or U2710 (N_2710,N_2490,N_2573);
and U2711 (N_2711,N_2458,N_2477);
nand U2712 (N_2712,N_2545,N_2513);
or U2713 (N_2713,N_2523,N_2547);
xnor U2714 (N_2714,N_2494,N_2577);
or U2715 (N_2715,N_2475,N_2470);
or U2716 (N_2716,N_2409,N_2450);
and U2717 (N_2717,N_2475,N_2494);
xor U2718 (N_2718,N_2517,N_2435);
xnor U2719 (N_2719,N_2428,N_2420);
and U2720 (N_2720,N_2560,N_2404);
or U2721 (N_2721,N_2574,N_2404);
xnor U2722 (N_2722,N_2490,N_2589);
or U2723 (N_2723,N_2508,N_2548);
xnor U2724 (N_2724,N_2464,N_2471);
or U2725 (N_2725,N_2407,N_2503);
or U2726 (N_2726,N_2492,N_2435);
nand U2727 (N_2727,N_2528,N_2564);
nor U2728 (N_2728,N_2515,N_2582);
or U2729 (N_2729,N_2431,N_2480);
xor U2730 (N_2730,N_2491,N_2566);
nor U2731 (N_2731,N_2414,N_2501);
or U2732 (N_2732,N_2527,N_2436);
nand U2733 (N_2733,N_2591,N_2475);
or U2734 (N_2734,N_2457,N_2471);
nor U2735 (N_2735,N_2419,N_2444);
nor U2736 (N_2736,N_2546,N_2458);
or U2737 (N_2737,N_2451,N_2471);
xor U2738 (N_2738,N_2452,N_2568);
and U2739 (N_2739,N_2574,N_2539);
nor U2740 (N_2740,N_2402,N_2467);
nor U2741 (N_2741,N_2473,N_2439);
and U2742 (N_2742,N_2451,N_2533);
xnor U2743 (N_2743,N_2539,N_2486);
nand U2744 (N_2744,N_2520,N_2495);
or U2745 (N_2745,N_2484,N_2428);
nor U2746 (N_2746,N_2482,N_2559);
or U2747 (N_2747,N_2418,N_2438);
and U2748 (N_2748,N_2574,N_2409);
nand U2749 (N_2749,N_2549,N_2475);
and U2750 (N_2750,N_2473,N_2565);
nor U2751 (N_2751,N_2529,N_2453);
nor U2752 (N_2752,N_2519,N_2472);
xor U2753 (N_2753,N_2505,N_2449);
nor U2754 (N_2754,N_2598,N_2557);
or U2755 (N_2755,N_2462,N_2405);
xor U2756 (N_2756,N_2522,N_2415);
or U2757 (N_2757,N_2431,N_2421);
and U2758 (N_2758,N_2490,N_2447);
nor U2759 (N_2759,N_2512,N_2534);
or U2760 (N_2760,N_2518,N_2511);
nand U2761 (N_2761,N_2558,N_2476);
xnor U2762 (N_2762,N_2569,N_2584);
xnor U2763 (N_2763,N_2561,N_2473);
nor U2764 (N_2764,N_2443,N_2593);
and U2765 (N_2765,N_2427,N_2457);
xor U2766 (N_2766,N_2420,N_2486);
or U2767 (N_2767,N_2587,N_2583);
xor U2768 (N_2768,N_2527,N_2590);
or U2769 (N_2769,N_2514,N_2570);
xor U2770 (N_2770,N_2438,N_2572);
nor U2771 (N_2771,N_2589,N_2450);
xor U2772 (N_2772,N_2420,N_2496);
nand U2773 (N_2773,N_2539,N_2559);
xor U2774 (N_2774,N_2434,N_2427);
or U2775 (N_2775,N_2439,N_2533);
nor U2776 (N_2776,N_2466,N_2461);
xnor U2777 (N_2777,N_2534,N_2498);
and U2778 (N_2778,N_2549,N_2489);
nor U2779 (N_2779,N_2552,N_2457);
xnor U2780 (N_2780,N_2478,N_2568);
nor U2781 (N_2781,N_2500,N_2593);
nor U2782 (N_2782,N_2593,N_2552);
and U2783 (N_2783,N_2512,N_2412);
or U2784 (N_2784,N_2569,N_2511);
nand U2785 (N_2785,N_2572,N_2588);
or U2786 (N_2786,N_2574,N_2468);
xnor U2787 (N_2787,N_2402,N_2418);
nand U2788 (N_2788,N_2537,N_2591);
nor U2789 (N_2789,N_2508,N_2462);
nand U2790 (N_2790,N_2569,N_2557);
nand U2791 (N_2791,N_2572,N_2510);
nor U2792 (N_2792,N_2435,N_2536);
nand U2793 (N_2793,N_2504,N_2425);
or U2794 (N_2794,N_2580,N_2493);
and U2795 (N_2795,N_2549,N_2452);
xnor U2796 (N_2796,N_2573,N_2463);
or U2797 (N_2797,N_2562,N_2409);
xnor U2798 (N_2798,N_2525,N_2461);
nor U2799 (N_2799,N_2596,N_2489);
xnor U2800 (N_2800,N_2639,N_2672);
nand U2801 (N_2801,N_2635,N_2686);
nand U2802 (N_2802,N_2612,N_2630);
and U2803 (N_2803,N_2775,N_2749);
and U2804 (N_2804,N_2627,N_2696);
nor U2805 (N_2805,N_2680,N_2764);
nor U2806 (N_2806,N_2768,N_2713);
nand U2807 (N_2807,N_2670,N_2755);
nor U2808 (N_2808,N_2602,N_2700);
or U2809 (N_2809,N_2750,N_2788);
or U2810 (N_2810,N_2625,N_2721);
or U2811 (N_2811,N_2714,N_2632);
or U2812 (N_2812,N_2648,N_2781);
nand U2813 (N_2813,N_2640,N_2608);
xnor U2814 (N_2814,N_2615,N_2616);
nand U2815 (N_2815,N_2682,N_2646);
nand U2816 (N_2816,N_2609,N_2786);
and U2817 (N_2817,N_2666,N_2614);
xor U2818 (N_2818,N_2730,N_2641);
or U2819 (N_2819,N_2743,N_2758);
nand U2820 (N_2820,N_2643,N_2657);
nor U2821 (N_2821,N_2791,N_2711);
xnor U2822 (N_2822,N_2681,N_2606);
or U2823 (N_2823,N_2604,N_2620);
nand U2824 (N_2824,N_2633,N_2738);
nand U2825 (N_2825,N_2601,N_2794);
nor U2826 (N_2826,N_2645,N_2770);
or U2827 (N_2827,N_2676,N_2732);
nor U2828 (N_2828,N_2787,N_2754);
nand U2829 (N_2829,N_2647,N_2663);
or U2830 (N_2830,N_2626,N_2741);
and U2831 (N_2831,N_2629,N_2780);
and U2832 (N_2832,N_2740,N_2623);
nor U2833 (N_2833,N_2603,N_2733);
and U2834 (N_2834,N_2659,N_2656);
nand U2835 (N_2835,N_2783,N_2644);
or U2836 (N_2836,N_2724,N_2655);
and U2837 (N_2837,N_2708,N_2600);
xor U2838 (N_2838,N_2718,N_2756);
nand U2839 (N_2839,N_2717,N_2747);
xor U2840 (N_2840,N_2766,N_2729);
xnor U2841 (N_2841,N_2765,N_2723);
xnor U2842 (N_2842,N_2618,N_2772);
nand U2843 (N_2843,N_2660,N_2607);
nor U2844 (N_2844,N_2795,N_2690);
or U2845 (N_2845,N_2720,N_2748);
nor U2846 (N_2846,N_2716,N_2691);
or U2847 (N_2847,N_2683,N_2636);
nand U2848 (N_2848,N_2761,N_2796);
nor U2849 (N_2849,N_2726,N_2688);
nor U2850 (N_2850,N_2728,N_2605);
nor U2851 (N_2851,N_2699,N_2777);
or U2852 (N_2852,N_2611,N_2739);
and U2853 (N_2853,N_2722,N_2707);
and U2854 (N_2854,N_2752,N_2649);
or U2855 (N_2855,N_2727,N_2624);
nor U2856 (N_2856,N_2631,N_2694);
xor U2857 (N_2857,N_2785,N_2712);
nor U2858 (N_2858,N_2746,N_2689);
or U2859 (N_2859,N_2737,N_2684);
or U2860 (N_2860,N_2710,N_2767);
or U2861 (N_2861,N_2703,N_2734);
or U2862 (N_2862,N_2651,N_2669);
and U2863 (N_2863,N_2695,N_2658);
nor U2864 (N_2864,N_2742,N_2705);
nand U2865 (N_2865,N_2771,N_2665);
nand U2866 (N_2866,N_2773,N_2673);
and U2867 (N_2867,N_2634,N_2709);
nand U2868 (N_2868,N_2745,N_2675);
and U2869 (N_2869,N_2744,N_2790);
nand U2870 (N_2870,N_2719,N_2693);
or U2871 (N_2871,N_2613,N_2753);
and U2872 (N_2872,N_2704,N_2619);
and U2873 (N_2873,N_2692,N_2760);
nor U2874 (N_2874,N_2735,N_2664);
xor U2875 (N_2875,N_2774,N_2685);
or U2876 (N_2876,N_2650,N_2642);
nor U2877 (N_2877,N_2662,N_2679);
or U2878 (N_2878,N_2671,N_2799);
or U2879 (N_2879,N_2698,N_2702);
nor U2880 (N_2880,N_2653,N_2674);
xor U2881 (N_2881,N_2762,N_2797);
nor U2882 (N_2882,N_2792,N_2652);
and U2883 (N_2883,N_2731,N_2798);
xnor U2884 (N_2884,N_2677,N_2654);
or U2885 (N_2885,N_2769,N_2793);
or U2886 (N_2886,N_2776,N_2667);
nand U2887 (N_2887,N_2736,N_2610);
nand U2888 (N_2888,N_2622,N_2621);
and U2889 (N_2889,N_2789,N_2687);
or U2890 (N_2890,N_2617,N_2759);
and U2891 (N_2891,N_2697,N_2725);
nand U2892 (N_2892,N_2706,N_2637);
and U2893 (N_2893,N_2757,N_2778);
or U2894 (N_2894,N_2779,N_2784);
nor U2895 (N_2895,N_2668,N_2715);
and U2896 (N_2896,N_2701,N_2678);
xnor U2897 (N_2897,N_2782,N_2638);
xnor U2898 (N_2898,N_2628,N_2751);
xor U2899 (N_2899,N_2661,N_2763);
and U2900 (N_2900,N_2779,N_2649);
and U2901 (N_2901,N_2741,N_2656);
nand U2902 (N_2902,N_2672,N_2649);
xnor U2903 (N_2903,N_2682,N_2774);
and U2904 (N_2904,N_2626,N_2795);
nor U2905 (N_2905,N_2730,N_2658);
or U2906 (N_2906,N_2744,N_2773);
nand U2907 (N_2907,N_2771,N_2716);
nor U2908 (N_2908,N_2726,N_2706);
xnor U2909 (N_2909,N_2610,N_2600);
nand U2910 (N_2910,N_2665,N_2706);
nor U2911 (N_2911,N_2602,N_2608);
nand U2912 (N_2912,N_2789,N_2761);
or U2913 (N_2913,N_2778,N_2700);
or U2914 (N_2914,N_2684,N_2715);
nand U2915 (N_2915,N_2646,N_2657);
nor U2916 (N_2916,N_2750,N_2602);
or U2917 (N_2917,N_2613,N_2751);
and U2918 (N_2918,N_2618,N_2625);
nand U2919 (N_2919,N_2678,N_2605);
or U2920 (N_2920,N_2695,N_2607);
or U2921 (N_2921,N_2613,N_2763);
and U2922 (N_2922,N_2781,N_2626);
nand U2923 (N_2923,N_2606,N_2743);
or U2924 (N_2924,N_2639,N_2760);
nor U2925 (N_2925,N_2653,N_2769);
and U2926 (N_2926,N_2687,N_2741);
nand U2927 (N_2927,N_2690,N_2617);
nand U2928 (N_2928,N_2703,N_2650);
nor U2929 (N_2929,N_2609,N_2689);
nor U2930 (N_2930,N_2738,N_2795);
xnor U2931 (N_2931,N_2701,N_2683);
nand U2932 (N_2932,N_2647,N_2734);
nor U2933 (N_2933,N_2610,N_2659);
xor U2934 (N_2934,N_2687,N_2792);
nand U2935 (N_2935,N_2773,N_2632);
xor U2936 (N_2936,N_2787,N_2617);
nand U2937 (N_2937,N_2684,N_2685);
and U2938 (N_2938,N_2631,N_2779);
and U2939 (N_2939,N_2738,N_2619);
and U2940 (N_2940,N_2724,N_2638);
and U2941 (N_2941,N_2606,N_2702);
nor U2942 (N_2942,N_2618,N_2730);
nand U2943 (N_2943,N_2702,N_2630);
or U2944 (N_2944,N_2688,N_2787);
and U2945 (N_2945,N_2719,N_2619);
and U2946 (N_2946,N_2615,N_2603);
nand U2947 (N_2947,N_2756,N_2791);
nor U2948 (N_2948,N_2663,N_2725);
and U2949 (N_2949,N_2630,N_2723);
xor U2950 (N_2950,N_2705,N_2726);
nor U2951 (N_2951,N_2795,N_2652);
or U2952 (N_2952,N_2701,N_2750);
xor U2953 (N_2953,N_2635,N_2673);
xor U2954 (N_2954,N_2796,N_2789);
nor U2955 (N_2955,N_2762,N_2654);
or U2956 (N_2956,N_2698,N_2757);
nand U2957 (N_2957,N_2752,N_2781);
xnor U2958 (N_2958,N_2730,N_2601);
and U2959 (N_2959,N_2610,N_2656);
xnor U2960 (N_2960,N_2694,N_2619);
and U2961 (N_2961,N_2748,N_2783);
xnor U2962 (N_2962,N_2625,N_2780);
xor U2963 (N_2963,N_2799,N_2697);
nand U2964 (N_2964,N_2691,N_2644);
and U2965 (N_2965,N_2704,N_2751);
and U2966 (N_2966,N_2726,N_2659);
xor U2967 (N_2967,N_2733,N_2796);
nor U2968 (N_2968,N_2739,N_2719);
xnor U2969 (N_2969,N_2664,N_2639);
and U2970 (N_2970,N_2744,N_2648);
nor U2971 (N_2971,N_2679,N_2640);
and U2972 (N_2972,N_2655,N_2699);
nor U2973 (N_2973,N_2708,N_2692);
or U2974 (N_2974,N_2631,N_2605);
nand U2975 (N_2975,N_2685,N_2687);
xor U2976 (N_2976,N_2634,N_2731);
xnor U2977 (N_2977,N_2687,N_2761);
and U2978 (N_2978,N_2753,N_2706);
nor U2979 (N_2979,N_2657,N_2605);
or U2980 (N_2980,N_2711,N_2653);
nor U2981 (N_2981,N_2688,N_2621);
nand U2982 (N_2982,N_2627,N_2625);
nor U2983 (N_2983,N_2613,N_2650);
and U2984 (N_2984,N_2781,N_2691);
nor U2985 (N_2985,N_2714,N_2604);
and U2986 (N_2986,N_2722,N_2725);
nand U2987 (N_2987,N_2762,N_2782);
xnor U2988 (N_2988,N_2682,N_2728);
nor U2989 (N_2989,N_2672,N_2650);
nor U2990 (N_2990,N_2613,N_2737);
xor U2991 (N_2991,N_2621,N_2638);
or U2992 (N_2992,N_2698,N_2634);
and U2993 (N_2993,N_2746,N_2612);
and U2994 (N_2994,N_2656,N_2674);
or U2995 (N_2995,N_2691,N_2614);
nand U2996 (N_2996,N_2748,N_2781);
or U2997 (N_2997,N_2750,N_2713);
nand U2998 (N_2998,N_2656,N_2782);
nor U2999 (N_2999,N_2787,N_2624);
and U3000 (N_3000,N_2924,N_2991);
xnor U3001 (N_3001,N_2853,N_2810);
xor U3002 (N_3002,N_2899,N_2851);
xnor U3003 (N_3003,N_2848,N_2831);
nor U3004 (N_3004,N_2852,N_2840);
nand U3005 (N_3005,N_2963,N_2844);
nand U3006 (N_3006,N_2898,N_2947);
nand U3007 (N_3007,N_2895,N_2864);
nand U3008 (N_3008,N_2925,N_2922);
or U3009 (N_3009,N_2964,N_2861);
xnor U3010 (N_3010,N_2958,N_2849);
or U3011 (N_3011,N_2982,N_2882);
xor U3012 (N_3012,N_2827,N_2870);
nand U3013 (N_3013,N_2955,N_2920);
nor U3014 (N_3014,N_2886,N_2806);
nand U3015 (N_3015,N_2868,N_2866);
and U3016 (N_3016,N_2966,N_2874);
nand U3017 (N_3017,N_2934,N_2807);
nand U3018 (N_3018,N_2915,N_2994);
and U3019 (N_3019,N_2904,N_2959);
and U3020 (N_3020,N_2987,N_2812);
nor U3021 (N_3021,N_2952,N_2903);
and U3022 (N_3022,N_2859,N_2912);
nand U3023 (N_3023,N_2818,N_2819);
and U3024 (N_3024,N_2967,N_2956);
xor U3025 (N_3025,N_2927,N_2858);
nor U3026 (N_3026,N_2824,N_2873);
nor U3027 (N_3027,N_2916,N_2829);
nor U3028 (N_3028,N_2802,N_2901);
xor U3029 (N_3029,N_2847,N_2826);
and U3030 (N_3030,N_2835,N_2932);
nand U3031 (N_3031,N_2983,N_2862);
xnor U3032 (N_3032,N_2816,N_2945);
and U3033 (N_3033,N_2979,N_2817);
and U3034 (N_3034,N_2871,N_2821);
and U3035 (N_3035,N_2875,N_2972);
nor U3036 (N_3036,N_2803,N_2970);
and U3037 (N_3037,N_2978,N_2909);
nand U3038 (N_3038,N_2804,N_2814);
or U3039 (N_3039,N_2973,N_2949);
nand U3040 (N_3040,N_2845,N_2836);
xor U3041 (N_3041,N_2855,N_2939);
or U3042 (N_3042,N_2943,N_2995);
or U3043 (N_3043,N_2885,N_2883);
or U3044 (N_3044,N_2998,N_2989);
xnor U3045 (N_3045,N_2999,N_2977);
or U3046 (N_3046,N_2888,N_2857);
nand U3047 (N_3047,N_2820,N_2974);
nor U3048 (N_3048,N_2872,N_2921);
nor U3049 (N_3049,N_2919,N_2877);
nand U3050 (N_3050,N_2842,N_2856);
xnor U3051 (N_3051,N_2910,N_2954);
or U3052 (N_3052,N_2838,N_2908);
nand U3053 (N_3053,N_2823,N_2962);
or U3054 (N_3054,N_2892,N_2928);
nor U3055 (N_3055,N_2992,N_2902);
nand U3056 (N_3056,N_2944,N_2953);
nor U3057 (N_3057,N_2834,N_2846);
or U3058 (N_3058,N_2897,N_2906);
and U3059 (N_3059,N_2905,N_2941);
nor U3060 (N_3060,N_2980,N_2907);
and U3061 (N_3061,N_2811,N_2911);
nor U3062 (N_3062,N_2996,N_2997);
nor U3063 (N_3063,N_2930,N_2984);
and U3064 (N_3064,N_2957,N_2813);
or U3065 (N_3065,N_2809,N_2931);
nor U3066 (N_3066,N_2976,N_2933);
or U3067 (N_3067,N_2950,N_2815);
and U3068 (N_3068,N_2938,N_2879);
xnor U3069 (N_3069,N_2854,N_2843);
nor U3070 (N_3070,N_2929,N_2968);
xnor U3071 (N_3071,N_2993,N_2960);
and U3072 (N_3072,N_2865,N_2981);
or U3073 (N_3073,N_2884,N_2841);
nor U3074 (N_3074,N_2832,N_2918);
nand U3075 (N_3075,N_2917,N_2990);
xor U3076 (N_3076,N_2869,N_2975);
or U3077 (N_3077,N_2881,N_2837);
xnor U3078 (N_3078,N_2808,N_2863);
nor U3079 (N_3079,N_2926,N_2914);
nor U3080 (N_3080,N_2860,N_2887);
xor U3081 (N_3081,N_2894,N_2900);
xor U3082 (N_3082,N_2890,N_2825);
xor U3083 (N_3083,N_2805,N_2801);
and U3084 (N_3084,N_2951,N_2850);
nor U3085 (N_3085,N_2896,N_2830);
nor U3086 (N_3086,N_2828,N_2889);
nand U3087 (N_3087,N_2822,N_2833);
nand U3088 (N_3088,N_2891,N_2935);
nor U3089 (N_3089,N_2867,N_2876);
and U3090 (N_3090,N_2988,N_2985);
and U3091 (N_3091,N_2878,N_2986);
nand U3092 (N_3092,N_2942,N_2800);
nor U3093 (N_3093,N_2923,N_2937);
or U3094 (N_3094,N_2948,N_2969);
xnor U3095 (N_3095,N_2961,N_2965);
or U3096 (N_3096,N_2913,N_2936);
nor U3097 (N_3097,N_2971,N_2940);
and U3098 (N_3098,N_2893,N_2839);
and U3099 (N_3099,N_2946,N_2880);
xnor U3100 (N_3100,N_2894,N_2906);
nor U3101 (N_3101,N_2824,N_2998);
nand U3102 (N_3102,N_2849,N_2950);
and U3103 (N_3103,N_2954,N_2881);
nor U3104 (N_3104,N_2983,N_2996);
nand U3105 (N_3105,N_2967,N_2965);
nand U3106 (N_3106,N_2983,N_2898);
nand U3107 (N_3107,N_2872,N_2905);
nand U3108 (N_3108,N_2941,N_2807);
or U3109 (N_3109,N_2826,N_2896);
and U3110 (N_3110,N_2819,N_2830);
xnor U3111 (N_3111,N_2991,N_2825);
or U3112 (N_3112,N_2834,N_2878);
nor U3113 (N_3113,N_2926,N_2878);
and U3114 (N_3114,N_2815,N_2933);
xor U3115 (N_3115,N_2885,N_2818);
nand U3116 (N_3116,N_2833,N_2816);
xnor U3117 (N_3117,N_2904,N_2935);
xnor U3118 (N_3118,N_2972,N_2963);
xor U3119 (N_3119,N_2974,N_2947);
or U3120 (N_3120,N_2904,N_2908);
and U3121 (N_3121,N_2898,N_2954);
nand U3122 (N_3122,N_2801,N_2871);
nor U3123 (N_3123,N_2804,N_2992);
and U3124 (N_3124,N_2889,N_2920);
nand U3125 (N_3125,N_2942,N_2805);
or U3126 (N_3126,N_2901,N_2993);
nor U3127 (N_3127,N_2918,N_2855);
and U3128 (N_3128,N_2878,N_2854);
xor U3129 (N_3129,N_2850,N_2986);
nand U3130 (N_3130,N_2961,N_2975);
or U3131 (N_3131,N_2953,N_2946);
xor U3132 (N_3132,N_2846,N_2955);
nor U3133 (N_3133,N_2804,N_2865);
and U3134 (N_3134,N_2932,N_2836);
nor U3135 (N_3135,N_2940,N_2961);
nand U3136 (N_3136,N_2987,N_2901);
or U3137 (N_3137,N_2986,N_2886);
xnor U3138 (N_3138,N_2968,N_2949);
nor U3139 (N_3139,N_2980,N_2833);
nor U3140 (N_3140,N_2861,N_2939);
xnor U3141 (N_3141,N_2921,N_2866);
xor U3142 (N_3142,N_2924,N_2963);
and U3143 (N_3143,N_2894,N_2978);
and U3144 (N_3144,N_2884,N_2886);
nor U3145 (N_3145,N_2873,N_2986);
nand U3146 (N_3146,N_2904,N_2897);
xor U3147 (N_3147,N_2911,N_2855);
or U3148 (N_3148,N_2862,N_2802);
nor U3149 (N_3149,N_2985,N_2860);
xor U3150 (N_3150,N_2998,N_2904);
and U3151 (N_3151,N_2988,N_2834);
or U3152 (N_3152,N_2902,N_2925);
or U3153 (N_3153,N_2925,N_2894);
xor U3154 (N_3154,N_2985,N_2856);
or U3155 (N_3155,N_2871,N_2951);
xor U3156 (N_3156,N_2978,N_2981);
nor U3157 (N_3157,N_2815,N_2873);
or U3158 (N_3158,N_2813,N_2873);
nor U3159 (N_3159,N_2893,N_2809);
xor U3160 (N_3160,N_2965,N_2934);
xor U3161 (N_3161,N_2899,N_2871);
xnor U3162 (N_3162,N_2962,N_2862);
nand U3163 (N_3163,N_2841,N_2970);
nand U3164 (N_3164,N_2887,N_2926);
xnor U3165 (N_3165,N_2901,N_2919);
or U3166 (N_3166,N_2926,N_2814);
nand U3167 (N_3167,N_2851,N_2924);
nor U3168 (N_3168,N_2828,N_2817);
and U3169 (N_3169,N_2968,N_2915);
xnor U3170 (N_3170,N_2862,N_2845);
or U3171 (N_3171,N_2949,N_2928);
xor U3172 (N_3172,N_2967,N_2959);
or U3173 (N_3173,N_2978,N_2979);
xor U3174 (N_3174,N_2972,N_2895);
xor U3175 (N_3175,N_2925,N_2821);
nor U3176 (N_3176,N_2959,N_2841);
xor U3177 (N_3177,N_2847,N_2831);
nor U3178 (N_3178,N_2922,N_2911);
nand U3179 (N_3179,N_2933,N_2893);
and U3180 (N_3180,N_2879,N_2969);
nor U3181 (N_3181,N_2842,N_2912);
nor U3182 (N_3182,N_2908,N_2996);
xnor U3183 (N_3183,N_2948,N_2863);
xnor U3184 (N_3184,N_2976,N_2931);
and U3185 (N_3185,N_2812,N_2927);
or U3186 (N_3186,N_2893,N_2801);
xor U3187 (N_3187,N_2915,N_2843);
nand U3188 (N_3188,N_2996,N_2963);
xor U3189 (N_3189,N_2976,N_2980);
nand U3190 (N_3190,N_2920,N_2928);
xnor U3191 (N_3191,N_2935,N_2842);
or U3192 (N_3192,N_2898,N_2879);
nand U3193 (N_3193,N_2905,N_2837);
nor U3194 (N_3194,N_2907,N_2960);
nand U3195 (N_3195,N_2871,N_2864);
or U3196 (N_3196,N_2852,N_2863);
nor U3197 (N_3197,N_2994,N_2899);
and U3198 (N_3198,N_2943,N_2866);
or U3199 (N_3199,N_2837,N_2824);
xor U3200 (N_3200,N_3141,N_3116);
and U3201 (N_3201,N_3075,N_3064);
xor U3202 (N_3202,N_3019,N_3040);
xor U3203 (N_3203,N_3129,N_3083);
xnor U3204 (N_3204,N_3059,N_3166);
nor U3205 (N_3205,N_3155,N_3099);
nor U3206 (N_3206,N_3048,N_3024);
and U3207 (N_3207,N_3118,N_3168);
nor U3208 (N_3208,N_3011,N_3085);
nor U3209 (N_3209,N_3001,N_3189);
or U3210 (N_3210,N_3126,N_3162);
nor U3211 (N_3211,N_3097,N_3098);
or U3212 (N_3212,N_3092,N_3136);
nand U3213 (N_3213,N_3114,N_3177);
nor U3214 (N_3214,N_3113,N_3121);
or U3215 (N_3215,N_3005,N_3123);
nor U3216 (N_3216,N_3181,N_3161);
nand U3217 (N_3217,N_3179,N_3138);
and U3218 (N_3218,N_3086,N_3038);
xor U3219 (N_3219,N_3062,N_3016);
nand U3220 (N_3220,N_3159,N_3056);
xor U3221 (N_3221,N_3147,N_3195);
nor U3222 (N_3222,N_3151,N_3190);
nor U3223 (N_3223,N_3088,N_3046);
or U3224 (N_3224,N_3192,N_3144);
nor U3225 (N_3225,N_3057,N_3007);
nand U3226 (N_3226,N_3132,N_3013);
xnor U3227 (N_3227,N_3125,N_3087);
xor U3228 (N_3228,N_3010,N_3119);
or U3229 (N_3229,N_3146,N_3145);
nand U3230 (N_3230,N_3060,N_3030);
xor U3231 (N_3231,N_3026,N_3015);
and U3232 (N_3232,N_3152,N_3133);
nor U3233 (N_3233,N_3149,N_3041);
nand U3234 (N_3234,N_3020,N_3176);
nor U3235 (N_3235,N_3081,N_3187);
and U3236 (N_3236,N_3096,N_3182);
nand U3237 (N_3237,N_3003,N_3094);
nand U3238 (N_3238,N_3130,N_3006);
and U3239 (N_3239,N_3042,N_3063);
or U3240 (N_3240,N_3186,N_3037);
nand U3241 (N_3241,N_3029,N_3091);
nor U3242 (N_3242,N_3128,N_3169);
and U3243 (N_3243,N_3106,N_3143);
nand U3244 (N_3244,N_3110,N_3089);
xor U3245 (N_3245,N_3032,N_3178);
nand U3246 (N_3246,N_3154,N_3095);
or U3247 (N_3247,N_3072,N_3171);
nand U3248 (N_3248,N_3058,N_3153);
xor U3249 (N_3249,N_3053,N_3196);
or U3250 (N_3250,N_3012,N_3023);
xor U3251 (N_3251,N_3165,N_3148);
or U3252 (N_3252,N_3055,N_3080);
or U3253 (N_3253,N_3028,N_3049);
nor U3254 (N_3254,N_3185,N_3076);
nor U3255 (N_3255,N_3142,N_3051);
or U3256 (N_3256,N_3120,N_3140);
nor U3257 (N_3257,N_3111,N_3107);
and U3258 (N_3258,N_3043,N_3014);
nand U3259 (N_3259,N_3071,N_3199);
and U3260 (N_3260,N_3157,N_3082);
nand U3261 (N_3261,N_3115,N_3184);
nor U3262 (N_3262,N_3077,N_3137);
nand U3263 (N_3263,N_3090,N_3172);
nand U3264 (N_3264,N_3193,N_3194);
or U3265 (N_3265,N_3078,N_3052);
nor U3266 (N_3266,N_3069,N_3002);
or U3267 (N_3267,N_3039,N_3124);
xnor U3268 (N_3268,N_3070,N_3067);
nor U3269 (N_3269,N_3104,N_3008);
nor U3270 (N_3270,N_3197,N_3021);
and U3271 (N_3271,N_3093,N_3050);
or U3272 (N_3272,N_3073,N_3173);
nand U3273 (N_3273,N_3027,N_3164);
or U3274 (N_3274,N_3112,N_3127);
nand U3275 (N_3275,N_3108,N_3101);
or U3276 (N_3276,N_3160,N_3061);
and U3277 (N_3277,N_3035,N_3031);
or U3278 (N_3278,N_3188,N_3066);
xor U3279 (N_3279,N_3004,N_3009);
or U3280 (N_3280,N_3175,N_3174);
nand U3281 (N_3281,N_3084,N_3100);
xnor U3282 (N_3282,N_3131,N_3135);
xnor U3283 (N_3283,N_3167,N_3109);
or U3284 (N_3284,N_3183,N_3045);
nor U3285 (N_3285,N_3163,N_3134);
or U3286 (N_3286,N_3122,N_3102);
or U3287 (N_3287,N_3025,N_3033);
nor U3288 (N_3288,N_3017,N_3156);
nor U3289 (N_3289,N_3158,N_3044);
and U3290 (N_3290,N_3065,N_3198);
nor U3291 (N_3291,N_3191,N_3105);
nor U3292 (N_3292,N_3117,N_3054);
xnor U3293 (N_3293,N_3047,N_3103);
or U3294 (N_3294,N_3000,N_3180);
or U3295 (N_3295,N_3018,N_3139);
or U3296 (N_3296,N_3034,N_3150);
and U3297 (N_3297,N_3068,N_3170);
nor U3298 (N_3298,N_3079,N_3074);
nor U3299 (N_3299,N_3022,N_3036);
nand U3300 (N_3300,N_3101,N_3123);
nor U3301 (N_3301,N_3003,N_3180);
and U3302 (N_3302,N_3146,N_3045);
nand U3303 (N_3303,N_3149,N_3014);
and U3304 (N_3304,N_3017,N_3029);
and U3305 (N_3305,N_3131,N_3106);
xor U3306 (N_3306,N_3164,N_3102);
nor U3307 (N_3307,N_3150,N_3044);
nor U3308 (N_3308,N_3161,N_3083);
nand U3309 (N_3309,N_3191,N_3030);
nand U3310 (N_3310,N_3001,N_3013);
nor U3311 (N_3311,N_3023,N_3191);
xor U3312 (N_3312,N_3075,N_3091);
or U3313 (N_3313,N_3165,N_3003);
nand U3314 (N_3314,N_3114,N_3072);
or U3315 (N_3315,N_3070,N_3097);
xnor U3316 (N_3316,N_3163,N_3027);
and U3317 (N_3317,N_3120,N_3040);
nor U3318 (N_3318,N_3128,N_3179);
xnor U3319 (N_3319,N_3099,N_3103);
nand U3320 (N_3320,N_3023,N_3053);
or U3321 (N_3321,N_3095,N_3086);
nor U3322 (N_3322,N_3059,N_3094);
or U3323 (N_3323,N_3000,N_3114);
xor U3324 (N_3324,N_3039,N_3189);
nand U3325 (N_3325,N_3140,N_3166);
and U3326 (N_3326,N_3192,N_3019);
or U3327 (N_3327,N_3138,N_3005);
nand U3328 (N_3328,N_3078,N_3019);
xor U3329 (N_3329,N_3196,N_3033);
or U3330 (N_3330,N_3074,N_3095);
nand U3331 (N_3331,N_3092,N_3179);
nand U3332 (N_3332,N_3070,N_3041);
nor U3333 (N_3333,N_3192,N_3182);
nand U3334 (N_3334,N_3020,N_3179);
nor U3335 (N_3335,N_3006,N_3080);
nor U3336 (N_3336,N_3104,N_3036);
and U3337 (N_3337,N_3167,N_3054);
and U3338 (N_3338,N_3058,N_3161);
nor U3339 (N_3339,N_3033,N_3061);
and U3340 (N_3340,N_3026,N_3172);
nor U3341 (N_3341,N_3017,N_3166);
nand U3342 (N_3342,N_3045,N_3092);
nor U3343 (N_3343,N_3069,N_3198);
xnor U3344 (N_3344,N_3096,N_3108);
or U3345 (N_3345,N_3100,N_3065);
nand U3346 (N_3346,N_3069,N_3071);
and U3347 (N_3347,N_3028,N_3004);
and U3348 (N_3348,N_3145,N_3182);
nand U3349 (N_3349,N_3008,N_3099);
and U3350 (N_3350,N_3115,N_3123);
nor U3351 (N_3351,N_3044,N_3060);
nor U3352 (N_3352,N_3116,N_3010);
xor U3353 (N_3353,N_3056,N_3092);
nand U3354 (N_3354,N_3031,N_3106);
and U3355 (N_3355,N_3164,N_3160);
or U3356 (N_3356,N_3160,N_3171);
nor U3357 (N_3357,N_3101,N_3188);
xor U3358 (N_3358,N_3086,N_3005);
xnor U3359 (N_3359,N_3010,N_3095);
nor U3360 (N_3360,N_3180,N_3069);
xnor U3361 (N_3361,N_3042,N_3160);
xor U3362 (N_3362,N_3000,N_3068);
and U3363 (N_3363,N_3186,N_3039);
xor U3364 (N_3364,N_3137,N_3058);
and U3365 (N_3365,N_3085,N_3190);
nor U3366 (N_3366,N_3010,N_3157);
xor U3367 (N_3367,N_3172,N_3069);
nor U3368 (N_3368,N_3168,N_3035);
nand U3369 (N_3369,N_3023,N_3122);
nor U3370 (N_3370,N_3122,N_3077);
and U3371 (N_3371,N_3071,N_3141);
xnor U3372 (N_3372,N_3047,N_3161);
or U3373 (N_3373,N_3190,N_3100);
or U3374 (N_3374,N_3199,N_3039);
nor U3375 (N_3375,N_3151,N_3143);
xor U3376 (N_3376,N_3126,N_3190);
xor U3377 (N_3377,N_3040,N_3154);
and U3378 (N_3378,N_3147,N_3033);
and U3379 (N_3379,N_3096,N_3106);
xnor U3380 (N_3380,N_3157,N_3174);
or U3381 (N_3381,N_3159,N_3106);
or U3382 (N_3382,N_3072,N_3100);
or U3383 (N_3383,N_3031,N_3113);
and U3384 (N_3384,N_3164,N_3000);
nor U3385 (N_3385,N_3063,N_3077);
nand U3386 (N_3386,N_3108,N_3030);
xor U3387 (N_3387,N_3051,N_3171);
nand U3388 (N_3388,N_3047,N_3165);
xor U3389 (N_3389,N_3003,N_3007);
or U3390 (N_3390,N_3117,N_3013);
or U3391 (N_3391,N_3113,N_3103);
nand U3392 (N_3392,N_3028,N_3080);
xnor U3393 (N_3393,N_3136,N_3063);
or U3394 (N_3394,N_3161,N_3176);
and U3395 (N_3395,N_3091,N_3099);
xnor U3396 (N_3396,N_3143,N_3181);
nand U3397 (N_3397,N_3021,N_3064);
and U3398 (N_3398,N_3005,N_3025);
and U3399 (N_3399,N_3058,N_3009);
xor U3400 (N_3400,N_3359,N_3206);
or U3401 (N_3401,N_3235,N_3306);
or U3402 (N_3402,N_3335,N_3288);
and U3403 (N_3403,N_3212,N_3222);
xnor U3404 (N_3404,N_3389,N_3386);
xnor U3405 (N_3405,N_3279,N_3218);
nor U3406 (N_3406,N_3375,N_3347);
xor U3407 (N_3407,N_3376,N_3275);
and U3408 (N_3408,N_3249,N_3358);
nand U3409 (N_3409,N_3327,N_3228);
and U3410 (N_3410,N_3242,N_3263);
or U3411 (N_3411,N_3302,N_3274);
nand U3412 (N_3412,N_3293,N_3282);
or U3413 (N_3413,N_3277,N_3292);
xnor U3414 (N_3414,N_3334,N_3333);
xor U3415 (N_3415,N_3332,N_3337);
nand U3416 (N_3416,N_3202,N_3200);
and U3417 (N_3417,N_3244,N_3285);
or U3418 (N_3418,N_3323,N_3201);
nand U3419 (N_3419,N_3330,N_3252);
nand U3420 (N_3420,N_3314,N_3294);
nor U3421 (N_3421,N_3287,N_3384);
or U3422 (N_3422,N_3296,N_3204);
nand U3423 (N_3423,N_3239,N_3388);
nor U3424 (N_3424,N_3216,N_3398);
xor U3425 (N_3425,N_3355,N_3313);
and U3426 (N_3426,N_3234,N_3365);
nor U3427 (N_3427,N_3262,N_3341);
or U3428 (N_3428,N_3353,N_3290);
nor U3429 (N_3429,N_3383,N_3338);
and U3430 (N_3430,N_3297,N_3203);
or U3431 (N_3431,N_3309,N_3268);
nor U3432 (N_3432,N_3267,N_3369);
nand U3433 (N_3433,N_3397,N_3246);
nand U3434 (N_3434,N_3352,N_3344);
or U3435 (N_3435,N_3247,N_3390);
nand U3436 (N_3436,N_3250,N_3266);
and U3437 (N_3437,N_3303,N_3231);
nand U3438 (N_3438,N_3240,N_3260);
nand U3439 (N_3439,N_3245,N_3304);
or U3440 (N_3440,N_3393,N_3286);
nor U3441 (N_3441,N_3380,N_3326);
nor U3442 (N_3442,N_3350,N_3301);
nor U3443 (N_3443,N_3280,N_3254);
and U3444 (N_3444,N_3354,N_3382);
xnor U3445 (N_3445,N_3318,N_3232);
xor U3446 (N_3446,N_3394,N_3317);
or U3447 (N_3447,N_3362,N_3361);
nand U3448 (N_3448,N_3328,N_3300);
nor U3449 (N_3449,N_3289,N_3238);
or U3450 (N_3450,N_3230,N_3364);
nor U3451 (N_3451,N_3316,N_3272);
and U3452 (N_3452,N_3209,N_3366);
nand U3453 (N_3453,N_3324,N_3339);
and U3454 (N_3454,N_3224,N_3258);
nor U3455 (N_3455,N_3223,N_3295);
and U3456 (N_3456,N_3319,N_3342);
or U3457 (N_3457,N_3322,N_3227);
and U3458 (N_3458,N_3377,N_3284);
or U3459 (N_3459,N_3255,N_3367);
xor U3460 (N_3460,N_3276,N_3378);
and U3461 (N_3461,N_3311,N_3373);
xnor U3462 (N_3462,N_3357,N_3379);
nand U3463 (N_3463,N_3256,N_3221);
and U3464 (N_3464,N_3320,N_3281);
xnor U3465 (N_3465,N_3243,N_3237);
or U3466 (N_3466,N_3351,N_3208);
and U3467 (N_3467,N_3264,N_3315);
nor U3468 (N_3468,N_3211,N_3269);
and U3469 (N_3469,N_3372,N_3213);
nor U3470 (N_3470,N_3299,N_3370);
nor U3471 (N_3471,N_3205,N_3368);
xnor U3472 (N_3472,N_3253,N_3298);
xnor U3473 (N_3473,N_3374,N_3321);
nor U3474 (N_3474,N_3265,N_3336);
and U3475 (N_3475,N_3214,N_3312);
and U3476 (N_3476,N_3207,N_3226);
nor U3477 (N_3477,N_3259,N_3283);
or U3478 (N_3478,N_3308,N_3229);
nor U3479 (N_3479,N_3340,N_3251);
or U3480 (N_3480,N_3331,N_3307);
nor U3481 (N_3481,N_3310,N_3305);
or U3482 (N_3482,N_3391,N_3325);
nor U3483 (N_3483,N_3387,N_3360);
nor U3484 (N_3484,N_3248,N_3396);
or U3485 (N_3485,N_3257,N_3329);
or U3486 (N_3486,N_3225,N_3385);
or U3487 (N_3487,N_3343,N_3395);
xor U3488 (N_3488,N_3363,N_3291);
or U3489 (N_3489,N_3349,N_3371);
or U3490 (N_3490,N_3215,N_3348);
nand U3491 (N_3491,N_3233,N_3273);
and U3492 (N_3492,N_3345,N_3236);
and U3493 (N_3493,N_3210,N_3346);
xor U3494 (N_3494,N_3261,N_3271);
and U3495 (N_3495,N_3278,N_3241);
or U3496 (N_3496,N_3392,N_3220);
nand U3497 (N_3497,N_3270,N_3217);
and U3498 (N_3498,N_3399,N_3219);
xnor U3499 (N_3499,N_3381,N_3356);
nand U3500 (N_3500,N_3244,N_3234);
xor U3501 (N_3501,N_3215,N_3373);
nand U3502 (N_3502,N_3212,N_3256);
and U3503 (N_3503,N_3239,N_3340);
xnor U3504 (N_3504,N_3375,N_3363);
nor U3505 (N_3505,N_3202,N_3374);
xnor U3506 (N_3506,N_3374,N_3227);
or U3507 (N_3507,N_3283,N_3261);
or U3508 (N_3508,N_3272,N_3374);
nor U3509 (N_3509,N_3387,N_3329);
or U3510 (N_3510,N_3324,N_3290);
or U3511 (N_3511,N_3310,N_3396);
nand U3512 (N_3512,N_3308,N_3258);
nand U3513 (N_3513,N_3229,N_3233);
xnor U3514 (N_3514,N_3246,N_3261);
nor U3515 (N_3515,N_3229,N_3375);
xor U3516 (N_3516,N_3381,N_3330);
nand U3517 (N_3517,N_3235,N_3316);
or U3518 (N_3518,N_3281,N_3207);
xor U3519 (N_3519,N_3245,N_3356);
nor U3520 (N_3520,N_3236,N_3287);
nor U3521 (N_3521,N_3339,N_3383);
nor U3522 (N_3522,N_3260,N_3327);
or U3523 (N_3523,N_3372,N_3360);
and U3524 (N_3524,N_3267,N_3338);
nor U3525 (N_3525,N_3369,N_3304);
and U3526 (N_3526,N_3227,N_3305);
nand U3527 (N_3527,N_3207,N_3271);
xnor U3528 (N_3528,N_3319,N_3361);
and U3529 (N_3529,N_3213,N_3361);
and U3530 (N_3530,N_3312,N_3242);
xor U3531 (N_3531,N_3282,N_3252);
and U3532 (N_3532,N_3207,N_3255);
and U3533 (N_3533,N_3389,N_3205);
nand U3534 (N_3534,N_3336,N_3312);
or U3535 (N_3535,N_3281,N_3377);
nor U3536 (N_3536,N_3315,N_3371);
or U3537 (N_3537,N_3220,N_3207);
nand U3538 (N_3538,N_3212,N_3377);
nor U3539 (N_3539,N_3366,N_3394);
and U3540 (N_3540,N_3219,N_3246);
xnor U3541 (N_3541,N_3276,N_3300);
xor U3542 (N_3542,N_3397,N_3383);
or U3543 (N_3543,N_3212,N_3263);
and U3544 (N_3544,N_3358,N_3231);
nand U3545 (N_3545,N_3251,N_3201);
nor U3546 (N_3546,N_3308,N_3376);
nor U3547 (N_3547,N_3305,N_3337);
or U3548 (N_3548,N_3321,N_3286);
nand U3549 (N_3549,N_3246,N_3356);
or U3550 (N_3550,N_3207,N_3217);
nand U3551 (N_3551,N_3215,N_3399);
nand U3552 (N_3552,N_3299,N_3329);
nor U3553 (N_3553,N_3257,N_3316);
nand U3554 (N_3554,N_3347,N_3208);
nand U3555 (N_3555,N_3382,N_3315);
and U3556 (N_3556,N_3205,N_3263);
nand U3557 (N_3557,N_3311,N_3289);
and U3558 (N_3558,N_3354,N_3337);
or U3559 (N_3559,N_3206,N_3369);
or U3560 (N_3560,N_3363,N_3260);
nand U3561 (N_3561,N_3258,N_3372);
nor U3562 (N_3562,N_3242,N_3231);
or U3563 (N_3563,N_3301,N_3296);
and U3564 (N_3564,N_3214,N_3278);
and U3565 (N_3565,N_3334,N_3319);
and U3566 (N_3566,N_3331,N_3310);
and U3567 (N_3567,N_3271,N_3231);
xnor U3568 (N_3568,N_3279,N_3270);
xor U3569 (N_3569,N_3288,N_3268);
nand U3570 (N_3570,N_3243,N_3343);
or U3571 (N_3571,N_3212,N_3214);
nand U3572 (N_3572,N_3389,N_3395);
xnor U3573 (N_3573,N_3201,N_3278);
and U3574 (N_3574,N_3241,N_3368);
nand U3575 (N_3575,N_3211,N_3289);
xnor U3576 (N_3576,N_3202,N_3352);
or U3577 (N_3577,N_3378,N_3343);
nor U3578 (N_3578,N_3374,N_3301);
nor U3579 (N_3579,N_3286,N_3212);
xor U3580 (N_3580,N_3346,N_3329);
and U3581 (N_3581,N_3303,N_3398);
nand U3582 (N_3582,N_3333,N_3323);
nand U3583 (N_3583,N_3367,N_3233);
nand U3584 (N_3584,N_3317,N_3300);
nor U3585 (N_3585,N_3250,N_3323);
nand U3586 (N_3586,N_3243,N_3379);
xnor U3587 (N_3587,N_3252,N_3306);
and U3588 (N_3588,N_3395,N_3235);
xnor U3589 (N_3589,N_3302,N_3346);
or U3590 (N_3590,N_3201,N_3392);
xor U3591 (N_3591,N_3228,N_3292);
nand U3592 (N_3592,N_3395,N_3396);
and U3593 (N_3593,N_3244,N_3363);
xor U3594 (N_3594,N_3298,N_3284);
and U3595 (N_3595,N_3219,N_3216);
or U3596 (N_3596,N_3231,N_3262);
nand U3597 (N_3597,N_3349,N_3226);
xor U3598 (N_3598,N_3344,N_3250);
xnor U3599 (N_3599,N_3367,N_3218);
or U3600 (N_3600,N_3584,N_3409);
or U3601 (N_3601,N_3460,N_3585);
or U3602 (N_3602,N_3527,N_3405);
nor U3603 (N_3603,N_3446,N_3440);
xnor U3604 (N_3604,N_3562,N_3500);
nand U3605 (N_3605,N_3422,N_3519);
and U3606 (N_3606,N_3563,N_3525);
or U3607 (N_3607,N_3407,N_3454);
nor U3608 (N_3608,N_3566,N_3415);
xor U3609 (N_3609,N_3553,N_3521);
xnor U3610 (N_3610,N_3499,N_3464);
nand U3611 (N_3611,N_3469,N_3512);
xor U3612 (N_3612,N_3557,N_3581);
nand U3613 (N_3613,N_3477,N_3474);
and U3614 (N_3614,N_3449,N_3536);
or U3615 (N_3615,N_3551,N_3411);
nand U3616 (N_3616,N_3430,N_3567);
and U3617 (N_3617,N_3442,N_3421);
nand U3618 (N_3618,N_3548,N_3495);
nand U3619 (N_3619,N_3423,N_3559);
xnor U3620 (N_3620,N_3485,N_3540);
xnor U3621 (N_3621,N_3556,N_3510);
or U3622 (N_3622,N_3480,N_3537);
xor U3623 (N_3623,N_3457,N_3478);
and U3624 (N_3624,N_3497,N_3417);
nor U3625 (N_3625,N_3573,N_3441);
nand U3626 (N_3626,N_3578,N_3513);
or U3627 (N_3627,N_3443,N_3444);
nor U3628 (N_3628,N_3429,N_3428);
nand U3629 (N_3629,N_3574,N_3471);
and U3630 (N_3630,N_3436,N_3598);
xor U3631 (N_3631,N_3432,N_3597);
nand U3632 (N_3632,N_3491,N_3552);
xnor U3633 (N_3633,N_3522,N_3487);
nor U3634 (N_3634,N_3472,N_3586);
nand U3635 (N_3635,N_3410,N_3418);
xnor U3636 (N_3636,N_3402,N_3572);
nand U3637 (N_3637,N_3504,N_3403);
or U3638 (N_3638,N_3558,N_3517);
and U3639 (N_3639,N_3550,N_3484);
nand U3640 (N_3640,N_3535,N_3467);
and U3641 (N_3641,N_3524,N_3544);
nand U3642 (N_3642,N_3425,N_3515);
xnor U3643 (N_3643,N_3420,N_3528);
and U3644 (N_3644,N_3486,N_3530);
nand U3645 (N_3645,N_3571,N_3577);
nand U3646 (N_3646,N_3498,N_3489);
xnor U3647 (N_3647,N_3419,N_3564);
or U3648 (N_3648,N_3408,N_3455);
nand U3649 (N_3649,N_3549,N_3523);
nand U3650 (N_3650,N_3416,N_3545);
and U3651 (N_3651,N_3599,N_3511);
nor U3652 (N_3652,N_3518,N_3539);
nor U3653 (N_3653,N_3505,N_3452);
and U3654 (N_3654,N_3435,N_3470);
or U3655 (N_3655,N_3414,N_3588);
or U3656 (N_3656,N_3493,N_3488);
nor U3657 (N_3657,N_3547,N_3501);
and U3658 (N_3658,N_3568,N_3592);
nor U3659 (N_3659,N_3502,N_3582);
nor U3660 (N_3660,N_3575,N_3426);
and U3661 (N_3661,N_3579,N_3533);
nand U3662 (N_3662,N_3561,N_3476);
nor U3663 (N_3663,N_3459,N_3438);
and U3664 (N_3664,N_3496,N_3412);
nor U3665 (N_3665,N_3424,N_3433);
nor U3666 (N_3666,N_3570,N_3531);
nand U3667 (N_3667,N_3596,N_3481);
or U3668 (N_3668,N_3445,N_3437);
nand U3669 (N_3669,N_3590,N_3509);
and U3670 (N_3670,N_3462,N_3401);
or U3671 (N_3671,N_3434,N_3580);
nand U3672 (N_3672,N_3456,N_3514);
nor U3673 (N_3673,N_3516,N_3542);
or U3674 (N_3674,N_3587,N_3555);
and U3675 (N_3675,N_3560,N_3482);
nand U3676 (N_3676,N_3554,N_3526);
nor U3677 (N_3677,N_3413,N_3507);
or U3678 (N_3678,N_3494,N_3594);
and U3679 (N_3679,N_3439,N_3534);
xnor U3680 (N_3680,N_3538,N_3453);
nand U3681 (N_3681,N_3520,N_3479);
nand U3682 (N_3682,N_3503,N_3569);
nand U3683 (N_3683,N_3475,N_3506);
and U3684 (N_3684,N_3591,N_3593);
and U3685 (N_3685,N_3431,N_3595);
or U3686 (N_3686,N_3543,N_3400);
nand U3687 (N_3687,N_3450,N_3546);
and U3688 (N_3688,N_3465,N_3473);
or U3689 (N_3689,N_3448,N_3427);
and U3690 (N_3690,N_3583,N_3466);
and U3691 (N_3691,N_3508,N_3490);
nand U3692 (N_3692,N_3461,N_3492);
xnor U3693 (N_3693,N_3532,N_3463);
nand U3694 (N_3694,N_3483,N_3447);
nor U3695 (N_3695,N_3541,N_3565);
nor U3696 (N_3696,N_3451,N_3589);
and U3697 (N_3697,N_3458,N_3529);
nand U3698 (N_3698,N_3468,N_3576);
nand U3699 (N_3699,N_3404,N_3406);
nand U3700 (N_3700,N_3549,N_3413);
and U3701 (N_3701,N_3549,N_3434);
and U3702 (N_3702,N_3491,N_3407);
or U3703 (N_3703,N_3420,N_3410);
and U3704 (N_3704,N_3402,N_3407);
or U3705 (N_3705,N_3579,N_3515);
and U3706 (N_3706,N_3523,N_3417);
xor U3707 (N_3707,N_3434,N_3589);
and U3708 (N_3708,N_3581,N_3401);
nand U3709 (N_3709,N_3490,N_3486);
and U3710 (N_3710,N_3538,N_3489);
nor U3711 (N_3711,N_3564,N_3422);
xnor U3712 (N_3712,N_3456,N_3441);
nand U3713 (N_3713,N_3552,N_3425);
xor U3714 (N_3714,N_3582,N_3564);
nand U3715 (N_3715,N_3533,N_3452);
xnor U3716 (N_3716,N_3540,N_3441);
nand U3717 (N_3717,N_3418,N_3551);
nor U3718 (N_3718,N_3528,N_3539);
nor U3719 (N_3719,N_3537,N_3402);
or U3720 (N_3720,N_3447,N_3468);
xnor U3721 (N_3721,N_3595,N_3439);
xor U3722 (N_3722,N_3598,N_3440);
nand U3723 (N_3723,N_3508,N_3523);
xnor U3724 (N_3724,N_3563,N_3540);
xor U3725 (N_3725,N_3495,N_3479);
and U3726 (N_3726,N_3533,N_3460);
nor U3727 (N_3727,N_3576,N_3563);
or U3728 (N_3728,N_3559,N_3471);
xnor U3729 (N_3729,N_3438,N_3502);
xnor U3730 (N_3730,N_3557,N_3465);
and U3731 (N_3731,N_3519,N_3454);
nor U3732 (N_3732,N_3435,N_3542);
nor U3733 (N_3733,N_3454,N_3594);
or U3734 (N_3734,N_3453,N_3578);
nand U3735 (N_3735,N_3532,N_3423);
nand U3736 (N_3736,N_3485,N_3541);
and U3737 (N_3737,N_3436,N_3501);
nor U3738 (N_3738,N_3541,N_3460);
nor U3739 (N_3739,N_3547,N_3577);
nor U3740 (N_3740,N_3505,N_3448);
or U3741 (N_3741,N_3442,N_3450);
xnor U3742 (N_3742,N_3565,N_3526);
nor U3743 (N_3743,N_3598,N_3447);
nor U3744 (N_3744,N_3553,N_3528);
nand U3745 (N_3745,N_3538,N_3448);
nand U3746 (N_3746,N_3573,N_3517);
or U3747 (N_3747,N_3403,N_3467);
xor U3748 (N_3748,N_3538,N_3422);
nand U3749 (N_3749,N_3587,N_3488);
nand U3750 (N_3750,N_3571,N_3512);
nand U3751 (N_3751,N_3506,N_3431);
and U3752 (N_3752,N_3598,N_3421);
nand U3753 (N_3753,N_3468,N_3579);
or U3754 (N_3754,N_3568,N_3493);
nor U3755 (N_3755,N_3488,N_3536);
and U3756 (N_3756,N_3430,N_3440);
and U3757 (N_3757,N_3540,N_3436);
nor U3758 (N_3758,N_3443,N_3507);
xor U3759 (N_3759,N_3515,N_3446);
nor U3760 (N_3760,N_3523,N_3452);
nand U3761 (N_3761,N_3449,N_3480);
xnor U3762 (N_3762,N_3578,N_3529);
nand U3763 (N_3763,N_3442,N_3568);
and U3764 (N_3764,N_3542,N_3537);
nand U3765 (N_3765,N_3438,N_3441);
and U3766 (N_3766,N_3409,N_3502);
or U3767 (N_3767,N_3515,N_3469);
nor U3768 (N_3768,N_3583,N_3407);
nor U3769 (N_3769,N_3470,N_3527);
xor U3770 (N_3770,N_3403,N_3583);
and U3771 (N_3771,N_3400,N_3453);
or U3772 (N_3772,N_3530,N_3494);
nor U3773 (N_3773,N_3479,N_3564);
xnor U3774 (N_3774,N_3486,N_3532);
or U3775 (N_3775,N_3415,N_3423);
nor U3776 (N_3776,N_3596,N_3430);
and U3777 (N_3777,N_3434,N_3570);
nand U3778 (N_3778,N_3595,N_3569);
or U3779 (N_3779,N_3521,N_3590);
xnor U3780 (N_3780,N_3557,N_3542);
or U3781 (N_3781,N_3548,N_3416);
xnor U3782 (N_3782,N_3462,N_3589);
or U3783 (N_3783,N_3425,N_3531);
nand U3784 (N_3784,N_3430,N_3400);
or U3785 (N_3785,N_3598,N_3498);
nand U3786 (N_3786,N_3406,N_3408);
xor U3787 (N_3787,N_3558,N_3568);
xor U3788 (N_3788,N_3546,N_3453);
nor U3789 (N_3789,N_3436,N_3468);
and U3790 (N_3790,N_3430,N_3402);
nor U3791 (N_3791,N_3510,N_3580);
and U3792 (N_3792,N_3445,N_3456);
or U3793 (N_3793,N_3521,N_3435);
or U3794 (N_3794,N_3517,N_3461);
nor U3795 (N_3795,N_3426,N_3586);
xor U3796 (N_3796,N_3505,N_3500);
and U3797 (N_3797,N_3488,N_3462);
or U3798 (N_3798,N_3437,N_3584);
nand U3799 (N_3799,N_3551,N_3575);
nand U3800 (N_3800,N_3718,N_3647);
nor U3801 (N_3801,N_3711,N_3683);
and U3802 (N_3802,N_3777,N_3754);
or U3803 (N_3803,N_3785,N_3692);
xor U3804 (N_3804,N_3731,N_3627);
nor U3805 (N_3805,N_3618,N_3600);
and U3806 (N_3806,N_3659,N_3727);
and U3807 (N_3807,N_3742,N_3697);
nand U3808 (N_3808,N_3679,N_3724);
nor U3809 (N_3809,N_3781,N_3721);
or U3810 (N_3810,N_3734,N_3793);
nor U3811 (N_3811,N_3716,N_3786);
xnor U3812 (N_3812,N_3706,N_3748);
and U3813 (N_3813,N_3769,N_3732);
nor U3814 (N_3814,N_3637,N_3617);
nor U3815 (N_3815,N_3606,N_3789);
or U3816 (N_3816,N_3794,N_3714);
or U3817 (N_3817,N_3788,N_3642);
nor U3818 (N_3818,N_3750,N_3644);
and U3819 (N_3819,N_3796,N_3755);
or U3820 (N_3820,N_3779,N_3611);
and U3821 (N_3821,N_3656,N_3751);
xor U3822 (N_3822,N_3763,N_3704);
or U3823 (N_3823,N_3649,N_3638);
or U3824 (N_3824,N_3625,N_3792);
and U3825 (N_3825,N_3621,N_3672);
or U3826 (N_3826,N_3626,N_3631);
and U3827 (N_3827,N_3613,N_3798);
or U3828 (N_3828,N_3743,N_3673);
or U3829 (N_3829,N_3761,N_3620);
nand U3830 (N_3830,N_3665,N_3605);
and U3831 (N_3831,N_3681,N_3765);
nor U3832 (N_3832,N_3680,N_3653);
xor U3833 (N_3833,N_3787,N_3738);
nand U3834 (N_3834,N_3699,N_3780);
or U3835 (N_3835,N_3753,N_3703);
or U3836 (N_3836,N_3614,N_3691);
nand U3837 (N_3837,N_3773,N_3641);
or U3838 (N_3838,N_3624,N_3776);
nor U3839 (N_3839,N_3764,N_3768);
xor U3840 (N_3840,N_3607,N_3729);
xor U3841 (N_3841,N_3602,N_3640);
and U3842 (N_3842,N_3636,N_3762);
nor U3843 (N_3843,N_3689,N_3759);
nor U3844 (N_3844,N_3654,N_3630);
nand U3845 (N_3845,N_3662,N_3799);
nand U3846 (N_3846,N_3682,N_3639);
nor U3847 (N_3847,N_3666,N_3717);
xor U3848 (N_3848,N_3609,N_3733);
or U3849 (N_3849,N_3752,N_3702);
and U3850 (N_3850,N_3745,N_3661);
and U3851 (N_3851,N_3628,N_3726);
xor U3852 (N_3852,N_3728,N_3712);
and U3853 (N_3853,N_3686,N_3629);
and U3854 (N_3854,N_3667,N_3645);
xor U3855 (N_3855,N_3676,N_3736);
xor U3856 (N_3856,N_3719,N_3713);
and U3857 (N_3857,N_3778,N_3670);
or U3858 (N_3858,N_3635,N_3693);
or U3859 (N_3859,N_3674,N_3690);
xor U3860 (N_3860,N_3700,N_3657);
or U3861 (N_3861,N_3797,N_3756);
and U3862 (N_3862,N_3610,N_3705);
nor U3863 (N_3863,N_3740,N_3650);
nand U3864 (N_3864,N_3677,N_3723);
nand U3865 (N_3865,N_3744,N_3646);
nor U3866 (N_3866,N_3766,N_3771);
xnor U3867 (N_3867,N_3668,N_3678);
and U3868 (N_3868,N_3725,N_3648);
nor U3869 (N_3869,N_3695,N_3601);
xor U3870 (N_3870,N_3660,N_3772);
xnor U3871 (N_3871,N_3782,N_3634);
nor U3872 (N_3872,N_3767,N_3612);
nor U3873 (N_3873,N_3757,N_3669);
and U3874 (N_3874,N_3608,N_3758);
nand U3875 (N_3875,N_3675,N_3619);
or U3876 (N_3876,N_3749,N_3791);
nor U3877 (N_3877,N_3663,N_3687);
xor U3878 (N_3878,N_3658,N_3715);
nand U3879 (N_3879,N_3710,N_3688);
nor U3880 (N_3880,N_3664,N_3655);
xor U3881 (N_3881,N_3746,N_3615);
or U3882 (N_3882,N_3739,N_3790);
and U3883 (N_3883,N_3623,N_3694);
nand U3884 (N_3884,N_3671,N_3747);
xnor U3885 (N_3885,N_3616,N_3603);
or U3886 (N_3886,N_3775,N_3722);
xor U3887 (N_3887,N_3698,N_3701);
xnor U3888 (N_3888,N_3760,N_3709);
xor U3889 (N_3889,N_3784,N_3652);
nor U3890 (N_3890,N_3737,N_3684);
xor U3891 (N_3891,N_3795,N_3622);
and U3892 (N_3892,N_3696,N_3730);
nor U3893 (N_3893,N_3774,N_3770);
nand U3894 (N_3894,N_3685,N_3735);
nor U3895 (N_3895,N_3651,N_3604);
nand U3896 (N_3896,N_3741,N_3708);
xnor U3897 (N_3897,N_3720,N_3633);
and U3898 (N_3898,N_3783,N_3707);
nand U3899 (N_3899,N_3632,N_3643);
and U3900 (N_3900,N_3709,N_3630);
or U3901 (N_3901,N_3744,N_3737);
nor U3902 (N_3902,N_3620,N_3720);
or U3903 (N_3903,N_3764,N_3638);
nand U3904 (N_3904,N_3687,N_3757);
xor U3905 (N_3905,N_3729,N_3600);
xnor U3906 (N_3906,N_3737,N_3680);
xor U3907 (N_3907,N_3639,N_3637);
xnor U3908 (N_3908,N_3664,N_3769);
nor U3909 (N_3909,N_3762,N_3607);
nor U3910 (N_3910,N_3654,N_3740);
or U3911 (N_3911,N_3695,N_3702);
xor U3912 (N_3912,N_3613,N_3692);
and U3913 (N_3913,N_3695,N_3635);
and U3914 (N_3914,N_3679,N_3688);
nand U3915 (N_3915,N_3762,N_3655);
xor U3916 (N_3916,N_3756,N_3631);
or U3917 (N_3917,N_3622,N_3648);
nand U3918 (N_3918,N_3670,N_3624);
xnor U3919 (N_3919,N_3600,N_3662);
nor U3920 (N_3920,N_3796,N_3653);
nor U3921 (N_3921,N_3762,N_3657);
or U3922 (N_3922,N_3767,N_3626);
nand U3923 (N_3923,N_3763,N_3785);
and U3924 (N_3924,N_3725,N_3730);
and U3925 (N_3925,N_3620,N_3652);
nand U3926 (N_3926,N_3605,N_3774);
and U3927 (N_3927,N_3785,N_3708);
or U3928 (N_3928,N_3796,N_3616);
nand U3929 (N_3929,N_3705,N_3715);
nor U3930 (N_3930,N_3605,N_3696);
xor U3931 (N_3931,N_3794,N_3653);
xor U3932 (N_3932,N_3617,N_3760);
nor U3933 (N_3933,N_3601,N_3787);
and U3934 (N_3934,N_3761,N_3640);
or U3935 (N_3935,N_3638,N_3681);
xnor U3936 (N_3936,N_3763,N_3712);
and U3937 (N_3937,N_3635,N_3703);
nor U3938 (N_3938,N_3705,N_3731);
or U3939 (N_3939,N_3713,N_3601);
nand U3940 (N_3940,N_3705,N_3627);
and U3941 (N_3941,N_3791,N_3740);
nand U3942 (N_3942,N_3678,N_3642);
or U3943 (N_3943,N_3760,N_3708);
nand U3944 (N_3944,N_3719,N_3779);
nor U3945 (N_3945,N_3675,N_3660);
nor U3946 (N_3946,N_3735,N_3606);
or U3947 (N_3947,N_3610,N_3730);
nand U3948 (N_3948,N_3682,N_3752);
nor U3949 (N_3949,N_3661,N_3644);
nor U3950 (N_3950,N_3758,N_3796);
nand U3951 (N_3951,N_3714,N_3745);
xnor U3952 (N_3952,N_3781,N_3752);
nor U3953 (N_3953,N_3771,N_3673);
xor U3954 (N_3954,N_3663,N_3694);
xor U3955 (N_3955,N_3632,N_3691);
nor U3956 (N_3956,N_3633,N_3653);
nand U3957 (N_3957,N_3693,N_3645);
or U3958 (N_3958,N_3765,N_3745);
or U3959 (N_3959,N_3734,N_3654);
nand U3960 (N_3960,N_3639,N_3629);
xor U3961 (N_3961,N_3623,N_3754);
and U3962 (N_3962,N_3756,N_3678);
or U3963 (N_3963,N_3703,N_3781);
or U3964 (N_3964,N_3647,N_3745);
xnor U3965 (N_3965,N_3758,N_3792);
nand U3966 (N_3966,N_3743,N_3675);
or U3967 (N_3967,N_3760,N_3650);
nor U3968 (N_3968,N_3785,N_3720);
or U3969 (N_3969,N_3680,N_3714);
and U3970 (N_3970,N_3612,N_3715);
and U3971 (N_3971,N_3790,N_3772);
and U3972 (N_3972,N_3662,N_3689);
and U3973 (N_3973,N_3649,N_3635);
nor U3974 (N_3974,N_3617,N_3702);
xor U3975 (N_3975,N_3739,N_3675);
and U3976 (N_3976,N_3606,N_3624);
nand U3977 (N_3977,N_3662,N_3677);
nor U3978 (N_3978,N_3763,N_3710);
xor U3979 (N_3979,N_3709,N_3656);
or U3980 (N_3980,N_3703,N_3617);
xnor U3981 (N_3981,N_3781,N_3642);
nor U3982 (N_3982,N_3775,N_3659);
nor U3983 (N_3983,N_3774,N_3789);
or U3984 (N_3984,N_3636,N_3747);
or U3985 (N_3985,N_3619,N_3736);
xnor U3986 (N_3986,N_3660,N_3622);
nor U3987 (N_3987,N_3683,N_3714);
nor U3988 (N_3988,N_3670,N_3777);
nand U3989 (N_3989,N_3699,N_3773);
or U3990 (N_3990,N_3777,N_3792);
nor U3991 (N_3991,N_3745,N_3766);
or U3992 (N_3992,N_3696,N_3705);
nor U3993 (N_3993,N_3670,N_3642);
and U3994 (N_3994,N_3666,N_3748);
and U3995 (N_3995,N_3650,N_3624);
nand U3996 (N_3996,N_3755,N_3786);
xnor U3997 (N_3997,N_3628,N_3725);
nor U3998 (N_3998,N_3625,N_3635);
nor U3999 (N_3999,N_3744,N_3620);
nor U4000 (N_4000,N_3960,N_3934);
or U4001 (N_4001,N_3923,N_3889);
nand U4002 (N_4002,N_3875,N_3984);
nand U4003 (N_4003,N_3991,N_3822);
nand U4004 (N_4004,N_3814,N_3932);
and U4005 (N_4005,N_3989,N_3954);
xnor U4006 (N_4006,N_3827,N_3918);
xor U4007 (N_4007,N_3801,N_3941);
nand U4008 (N_4008,N_3919,N_3845);
nor U4009 (N_4009,N_3821,N_3961);
and U4010 (N_4010,N_3888,N_3841);
nand U4011 (N_4011,N_3800,N_3808);
or U4012 (N_4012,N_3933,N_3967);
nor U4013 (N_4013,N_3907,N_3832);
nor U4014 (N_4014,N_3839,N_3897);
nor U4015 (N_4015,N_3955,N_3892);
xnor U4016 (N_4016,N_3810,N_3980);
or U4017 (N_4017,N_3838,N_3862);
nor U4018 (N_4018,N_3968,N_3931);
nand U4019 (N_4019,N_3804,N_3886);
or U4020 (N_4020,N_3953,N_3908);
and U4021 (N_4021,N_3803,N_3971);
nor U4022 (N_4022,N_3902,N_3912);
xor U4023 (N_4023,N_3866,N_3915);
nor U4024 (N_4024,N_3950,N_3929);
xnor U4025 (N_4025,N_3859,N_3811);
nor U4026 (N_4026,N_3853,N_3986);
xor U4027 (N_4027,N_3865,N_3816);
or U4028 (N_4028,N_3863,N_3935);
and U4029 (N_4029,N_3812,N_3911);
or U4030 (N_4030,N_3946,N_3854);
nand U4031 (N_4031,N_3997,N_3921);
or U4032 (N_4032,N_3927,N_3834);
xnor U4033 (N_4033,N_3844,N_3995);
or U4034 (N_4034,N_3856,N_3940);
nor U4035 (N_4035,N_3881,N_3894);
or U4036 (N_4036,N_3817,N_3823);
and U4037 (N_4037,N_3899,N_3849);
nor U4038 (N_4038,N_3962,N_3824);
or U4039 (N_4039,N_3880,N_3998);
or U4040 (N_4040,N_3906,N_3951);
nand U4041 (N_4041,N_3871,N_3999);
nand U4042 (N_4042,N_3876,N_3973);
or U4043 (N_4043,N_3884,N_3861);
and U4044 (N_4044,N_3873,N_3891);
nor U4045 (N_4045,N_3835,N_3958);
xnor U4046 (N_4046,N_3868,N_3818);
xnor U4047 (N_4047,N_3837,N_3842);
or U4048 (N_4048,N_3936,N_3938);
xnor U4049 (N_4049,N_3969,N_3901);
or U4050 (N_4050,N_3981,N_3852);
and U4051 (N_4051,N_3964,N_3959);
and U4052 (N_4052,N_3952,N_3872);
xor U4053 (N_4053,N_3848,N_3963);
and U4054 (N_4054,N_3982,N_3975);
nand U4055 (N_4055,N_3949,N_3820);
and U4056 (N_4056,N_3979,N_3855);
xnor U4057 (N_4057,N_3885,N_3860);
xnor U4058 (N_4058,N_3813,N_3976);
or U4059 (N_4059,N_3833,N_3831);
nor U4060 (N_4060,N_3957,N_3994);
nor U4061 (N_4061,N_3992,N_3937);
nor U4062 (N_4062,N_3809,N_3978);
nor U4063 (N_4063,N_3914,N_3930);
xor U4064 (N_4064,N_3945,N_3883);
and U4065 (N_4065,N_3879,N_3895);
and U4066 (N_4066,N_3829,N_3864);
or U4067 (N_4067,N_3970,N_3898);
xnor U4068 (N_4068,N_3920,N_3926);
nand U4069 (N_4069,N_3836,N_3922);
nand U4070 (N_4070,N_3944,N_3987);
nor U4071 (N_4071,N_3806,N_3948);
and U4072 (N_4072,N_3828,N_3878);
nand U4073 (N_4073,N_3877,N_3928);
and U4074 (N_4074,N_3900,N_3887);
and U4075 (N_4075,N_3925,N_3867);
xnor U4076 (N_4076,N_3974,N_3947);
nor U4077 (N_4077,N_3857,N_3904);
nand U4078 (N_4078,N_3990,N_3802);
or U4079 (N_4079,N_3996,N_3896);
xnor U4080 (N_4080,N_3869,N_3826);
nand U4081 (N_4081,N_3850,N_3890);
nor U4082 (N_4082,N_3903,N_3966);
xnor U4083 (N_4083,N_3988,N_3870);
nor U4084 (N_4084,N_3913,N_3905);
xor U4085 (N_4085,N_3983,N_3893);
nand U4086 (N_4086,N_3943,N_3847);
xnor U4087 (N_4087,N_3874,N_3916);
nand U4088 (N_4088,N_3993,N_3843);
nand U4089 (N_4089,N_3819,N_3977);
or U4090 (N_4090,N_3924,N_3882);
or U4091 (N_4091,N_3917,N_3985);
nor U4092 (N_4092,N_3965,N_3956);
and U4093 (N_4093,N_3942,N_3939);
and U4094 (N_4094,N_3805,N_3858);
nor U4095 (N_4095,N_3909,N_3846);
and U4096 (N_4096,N_3807,N_3825);
and U4097 (N_4097,N_3815,N_3830);
xor U4098 (N_4098,N_3851,N_3840);
nor U4099 (N_4099,N_3972,N_3910);
xnor U4100 (N_4100,N_3932,N_3863);
nor U4101 (N_4101,N_3892,N_3941);
nor U4102 (N_4102,N_3973,N_3831);
and U4103 (N_4103,N_3864,N_3994);
xor U4104 (N_4104,N_3965,N_3859);
or U4105 (N_4105,N_3852,N_3811);
and U4106 (N_4106,N_3859,N_3899);
xnor U4107 (N_4107,N_3857,N_3957);
nand U4108 (N_4108,N_3852,N_3868);
or U4109 (N_4109,N_3934,N_3965);
nor U4110 (N_4110,N_3932,N_3995);
nor U4111 (N_4111,N_3808,N_3948);
nor U4112 (N_4112,N_3868,N_3923);
or U4113 (N_4113,N_3973,N_3857);
nand U4114 (N_4114,N_3988,N_3953);
nor U4115 (N_4115,N_3955,N_3808);
xnor U4116 (N_4116,N_3981,N_3938);
or U4117 (N_4117,N_3867,N_3946);
nor U4118 (N_4118,N_3987,N_3965);
nand U4119 (N_4119,N_3815,N_3967);
nor U4120 (N_4120,N_3826,N_3993);
and U4121 (N_4121,N_3944,N_3990);
nor U4122 (N_4122,N_3969,N_3902);
and U4123 (N_4123,N_3886,N_3856);
xor U4124 (N_4124,N_3914,N_3869);
nor U4125 (N_4125,N_3973,N_3894);
xnor U4126 (N_4126,N_3878,N_3837);
nand U4127 (N_4127,N_3876,N_3868);
or U4128 (N_4128,N_3884,N_3900);
and U4129 (N_4129,N_3946,N_3873);
xnor U4130 (N_4130,N_3941,N_3945);
nand U4131 (N_4131,N_3853,N_3968);
nor U4132 (N_4132,N_3859,N_3820);
nor U4133 (N_4133,N_3823,N_3952);
xor U4134 (N_4134,N_3999,N_3904);
nand U4135 (N_4135,N_3885,N_3986);
and U4136 (N_4136,N_3973,N_3860);
nand U4137 (N_4137,N_3961,N_3959);
or U4138 (N_4138,N_3933,N_3877);
xor U4139 (N_4139,N_3889,N_3885);
and U4140 (N_4140,N_3955,N_3801);
nor U4141 (N_4141,N_3894,N_3955);
and U4142 (N_4142,N_3942,N_3836);
xnor U4143 (N_4143,N_3859,N_3968);
nor U4144 (N_4144,N_3876,N_3829);
nand U4145 (N_4145,N_3984,N_3972);
nand U4146 (N_4146,N_3830,N_3992);
or U4147 (N_4147,N_3967,N_3931);
or U4148 (N_4148,N_3982,N_3855);
xnor U4149 (N_4149,N_3911,N_3829);
xor U4150 (N_4150,N_3863,N_3986);
nand U4151 (N_4151,N_3966,N_3859);
xor U4152 (N_4152,N_3989,N_3836);
nand U4153 (N_4153,N_3835,N_3979);
nand U4154 (N_4154,N_3953,N_3950);
xor U4155 (N_4155,N_3933,N_3845);
xnor U4156 (N_4156,N_3810,N_3975);
nand U4157 (N_4157,N_3915,N_3819);
nor U4158 (N_4158,N_3945,N_3919);
nor U4159 (N_4159,N_3832,N_3869);
nand U4160 (N_4160,N_3948,N_3940);
and U4161 (N_4161,N_3862,N_3854);
nor U4162 (N_4162,N_3875,N_3867);
xor U4163 (N_4163,N_3880,N_3855);
nor U4164 (N_4164,N_3930,N_3980);
nand U4165 (N_4165,N_3816,N_3925);
and U4166 (N_4166,N_3849,N_3979);
or U4167 (N_4167,N_3981,N_3890);
and U4168 (N_4168,N_3908,N_3944);
and U4169 (N_4169,N_3839,N_3830);
and U4170 (N_4170,N_3974,N_3822);
and U4171 (N_4171,N_3805,N_3904);
nor U4172 (N_4172,N_3864,N_3975);
and U4173 (N_4173,N_3990,N_3884);
xor U4174 (N_4174,N_3982,N_3858);
nor U4175 (N_4175,N_3908,N_3842);
and U4176 (N_4176,N_3856,N_3956);
and U4177 (N_4177,N_3909,N_3845);
nand U4178 (N_4178,N_3970,N_3909);
or U4179 (N_4179,N_3845,N_3903);
xnor U4180 (N_4180,N_3984,N_3891);
and U4181 (N_4181,N_3843,N_3937);
nand U4182 (N_4182,N_3818,N_3847);
or U4183 (N_4183,N_3891,N_3921);
and U4184 (N_4184,N_3913,N_3912);
and U4185 (N_4185,N_3966,N_3934);
and U4186 (N_4186,N_3924,N_3926);
nand U4187 (N_4187,N_3911,N_3943);
nor U4188 (N_4188,N_3952,N_3896);
and U4189 (N_4189,N_3960,N_3975);
nand U4190 (N_4190,N_3830,N_3807);
nor U4191 (N_4191,N_3974,N_3990);
or U4192 (N_4192,N_3901,N_3858);
nand U4193 (N_4193,N_3927,N_3825);
xor U4194 (N_4194,N_3915,N_3947);
nor U4195 (N_4195,N_3861,N_3845);
or U4196 (N_4196,N_3911,N_3915);
xnor U4197 (N_4197,N_3854,N_3905);
or U4198 (N_4198,N_3804,N_3914);
xnor U4199 (N_4199,N_3956,N_3868);
nor U4200 (N_4200,N_4159,N_4108);
and U4201 (N_4201,N_4043,N_4035);
nand U4202 (N_4202,N_4120,N_4123);
nand U4203 (N_4203,N_4110,N_4117);
and U4204 (N_4204,N_4080,N_4021);
nor U4205 (N_4205,N_4148,N_4175);
xnor U4206 (N_4206,N_4024,N_4011);
or U4207 (N_4207,N_4033,N_4121);
or U4208 (N_4208,N_4018,N_4126);
nor U4209 (N_4209,N_4057,N_4105);
nor U4210 (N_4210,N_4193,N_4194);
xnor U4211 (N_4211,N_4041,N_4083);
or U4212 (N_4212,N_4113,N_4149);
xnor U4213 (N_4213,N_4002,N_4009);
or U4214 (N_4214,N_4056,N_4196);
nand U4215 (N_4215,N_4107,N_4199);
nor U4216 (N_4216,N_4000,N_4156);
xor U4217 (N_4217,N_4114,N_4138);
nor U4218 (N_4218,N_4190,N_4029);
or U4219 (N_4219,N_4037,N_4042);
and U4220 (N_4220,N_4005,N_4028);
nor U4221 (N_4221,N_4001,N_4169);
nand U4222 (N_4222,N_4151,N_4177);
nand U4223 (N_4223,N_4004,N_4010);
nand U4224 (N_4224,N_4012,N_4109);
xnor U4225 (N_4225,N_4128,N_4170);
and U4226 (N_4226,N_4143,N_4058);
and U4227 (N_4227,N_4103,N_4036);
or U4228 (N_4228,N_4191,N_4136);
xnor U4229 (N_4229,N_4008,N_4066);
xor U4230 (N_4230,N_4118,N_4049);
nor U4231 (N_4231,N_4053,N_4071);
and U4232 (N_4232,N_4168,N_4050);
nand U4233 (N_4233,N_4052,N_4155);
and U4234 (N_4234,N_4074,N_4184);
nand U4235 (N_4235,N_4088,N_4097);
or U4236 (N_4236,N_4059,N_4069);
xnor U4237 (N_4237,N_4163,N_4179);
nor U4238 (N_4238,N_4051,N_4197);
and U4239 (N_4239,N_4189,N_4176);
nor U4240 (N_4240,N_4178,N_4072);
or U4241 (N_4241,N_4183,N_4137);
xor U4242 (N_4242,N_4104,N_4026);
nor U4243 (N_4243,N_4091,N_4034);
nand U4244 (N_4244,N_4082,N_4124);
and U4245 (N_4245,N_4016,N_4084);
xor U4246 (N_4246,N_4116,N_4048);
nor U4247 (N_4247,N_4046,N_4003);
xnor U4248 (N_4248,N_4192,N_4047);
nand U4249 (N_4249,N_4160,N_4065);
xor U4250 (N_4250,N_4164,N_4150);
or U4251 (N_4251,N_4073,N_4064);
or U4252 (N_4252,N_4135,N_4131);
or U4253 (N_4253,N_4078,N_4173);
or U4254 (N_4254,N_4022,N_4070);
xor U4255 (N_4255,N_4077,N_4141);
xor U4256 (N_4256,N_4076,N_4198);
nor U4257 (N_4257,N_4154,N_4090);
or U4258 (N_4258,N_4174,N_4133);
and U4259 (N_4259,N_4157,N_4032);
xnor U4260 (N_4260,N_4092,N_4039);
nand U4261 (N_4261,N_4098,N_4086);
and U4262 (N_4262,N_4172,N_4101);
xnor U4263 (N_4263,N_4015,N_4181);
and U4264 (N_4264,N_4106,N_4067);
nor U4265 (N_4265,N_4093,N_4099);
and U4266 (N_4266,N_4068,N_4102);
nor U4267 (N_4267,N_4115,N_4095);
nor U4268 (N_4268,N_4167,N_4013);
xor U4269 (N_4269,N_4038,N_4100);
xnor U4270 (N_4270,N_4014,N_4161);
or U4271 (N_4271,N_4125,N_4006);
xor U4272 (N_4272,N_4187,N_4055);
nor U4273 (N_4273,N_4030,N_4185);
and U4274 (N_4274,N_4119,N_4027);
and U4275 (N_4275,N_4122,N_4096);
and U4276 (N_4276,N_4165,N_4075);
nand U4277 (N_4277,N_4085,N_4060);
nand U4278 (N_4278,N_4017,N_4158);
xnor U4279 (N_4279,N_4171,N_4146);
and U4280 (N_4280,N_4061,N_4182);
and U4281 (N_4281,N_4019,N_4089);
nor U4282 (N_4282,N_4081,N_4153);
and U4283 (N_4283,N_4147,N_4139);
nand U4284 (N_4284,N_4144,N_4111);
nand U4285 (N_4285,N_4063,N_4087);
nor U4286 (N_4286,N_4044,N_4180);
or U4287 (N_4287,N_4142,N_4162);
and U4288 (N_4288,N_4040,N_4025);
xnor U4289 (N_4289,N_4020,N_4140);
xnor U4290 (N_4290,N_4145,N_4152);
nand U4291 (N_4291,N_4186,N_4127);
xor U4292 (N_4292,N_4045,N_4054);
nand U4293 (N_4293,N_4007,N_4023);
nor U4294 (N_4294,N_4132,N_4031);
xnor U4295 (N_4295,N_4195,N_4130);
nand U4296 (N_4296,N_4129,N_4094);
nor U4297 (N_4297,N_4062,N_4134);
and U4298 (N_4298,N_4112,N_4166);
and U4299 (N_4299,N_4188,N_4079);
xnor U4300 (N_4300,N_4190,N_4119);
or U4301 (N_4301,N_4162,N_4176);
or U4302 (N_4302,N_4176,N_4109);
nor U4303 (N_4303,N_4030,N_4176);
nand U4304 (N_4304,N_4128,N_4081);
or U4305 (N_4305,N_4037,N_4024);
and U4306 (N_4306,N_4169,N_4197);
xor U4307 (N_4307,N_4162,N_4145);
and U4308 (N_4308,N_4126,N_4144);
nand U4309 (N_4309,N_4043,N_4108);
or U4310 (N_4310,N_4117,N_4034);
nand U4311 (N_4311,N_4185,N_4147);
nor U4312 (N_4312,N_4030,N_4135);
xnor U4313 (N_4313,N_4032,N_4104);
and U4314 (N_4314,N_4058,N_4072);
xor U4315 (N_4315,N_4144,N_4159);
and U4316 (N_4316,N_4125,N_4059);
or U4317 (N_4317,N_4053,N_4170);
xnor U4318 (N_4318,N_4185,N_4084);
or U4319 (N_4319,N_4070,N_4014);
and U4320 (N_4320,N_4173,N_4133);
nor U4321 (N_4321,N_4171,N_4102);
nor U4322 (N_4322,N_4000,N_4049);
nand U4323 (N_4323,N_4085,N_4044);
xor U4324 (N_4324,N_4013,N_4177);
and U4325 (N_4325,N_4082,N_4072);
xor U4326 (N_4326,N_4003,N_4078);
nand U4327 (N_4327,N_4024,N_4142);
and U4328 (N_4328,N_4177,N_4144);
nor U4329 (N_4329,N_4033,N_4002);
or U4330 (N_4330,N_4188,N_4075);
nand U4331 (N_4331,N_4178,N_4137);
and U4332 (N_4332,N_4100,N_4179);
nor U4333 (N_4333,N_4178,N_4186);
xnor U4334 (N_4334,N_4126,N_4010);
nand U4335 (N_4335,N_4098,N_4145);
and U4336 (N_4336,N_4083,N_4183);
nor U4337 (N_4337,N_4094,N_4074);
xnor U4338 (N_4338,N_4068,N_4049);
and U4339 (N_4339,N_4157,N_4080);
or U4340 (N_4340,N_4047,N_4052);
nand U4341 (N_4341,N_4085,N_4181);
or U4342 (N_4342,N_4147,N_4003);
xnor U4343 (N_4343,N_4030,N_4192);
xor U4344 (N_4344,N_4099,N_4139);
or U4345 (N_4345,N_4086,N_4131);
xnor U4346 (N_4346,N_4151,N_4103);
or U4347 (N_4347,N_4164,N_4079);
or U4348 (N_4348,N_4089,N_4031);
nand U4349 (N_4349,N_4155,N_4109);
nand U4350 (N_4350,N_4076,N_4160);
nand U4351 (N_4351,N_4012,N_4142);
nand U4352 (N_4352,N_4160,N_4043);
nand U4353 (N_4353,N_4182,N_4172);
xor U4354 (N_4354,N_4111,N_4022);
nor U4355 (N_4355,N_4012,N_4033);
nor U4356 (N_4356,N_4169,N_4149);
xnor U4357 (N_4357,N_4114,N_4023);
nor U4358 (N_4358,N_4191,N_4098);
xnor U4359 (N_4359,N_4131,N_4004);
and U4360 (N_4360,N_4193,N_4190);
and U4361 (N_4361,N_4012,N_4139);
nor U4362 (N_4362,N_4177,N_4044);
or U4363 (N_4363,N_4142,N_4095);
and U4364 (N_4364,N_4028,N_4041);
and U4365 (N_4365,N_4162,N_4069);
nor U4366 (N_4366,N_4023,N_4195);
nand U4367 (N_4367,N_4137,N_4194);
or U4368 (N_4368,N_4104,N_4057);
and U4369 (N_4369,N_4014,N_4029);
or U4370 (N_4370,N_4006,N_4146);
nor U4371 (N_4371,N_4080,N_4065);
xor U4372 (N_4372,N_4154,N_4156);
nor U4373 (N_4373,N_4180,N_4096);
xor U4374 (N_4374,N_4012,N_4169);
or U4375 (N_4375,N_4020,N_4132);
nor U4376 (N_4376,N_4114,N_4004);
or U4377 (N_4377,N_4050,N_4176);
nand U4378 (N_4378,N_4161,N_4036);
and U4379 (N_4379,N_4021,N_4028);
nor U4380 (N_4380,N_4109,N_4158);
nand U4381 (N_4381,N_4133,N_4197);
nor U4382 (N_4382,N_4048,N_4176);
nand U4383 (N_4383,N_4001,N_4055);
or U4384 (N_4384,N_4035,N_4055);
nand U4385 (N_4385,N_4022,N_4038);
or U4386 (N_4386,N_4042,N_4157);
and U4387 (N_4387,N_4126,N_4131);
xor U4388 (N_4388,N_4112,N_4016);
nor U4389 (N_4389,N_4025,N_4143);
and U4390 (N_4390,N_4115,N_4164);
and U4391 (N_4391,N_4199,N_4181);
and U4392 (N_4392,N_4020,N_4017);
xnor U4393 (N_4393,N_4173,N_4064);
xnor U4394 (N_4394,N_4035,N_4175);
nor U4395 (N_4395,N_4099,N_4009);
xor U4396 (N_4396,N_4191,N_4052);
xor U4397 (N_4397,N_4026,N_4131);
or U4398 (N_4398,N_4120,N_4020);
or U4399 (N_4399,N_4015,N_4001);
and U4400 (N_4400,N_4341,N_4316);
and U4401 (N_4401,N_4270,N_4246);
and U4402 (N_4402,N_4299,N_4282);
nand U4403 (N_4403,N_4313,N_4204);
or U4404 (N_4404,N_4315,N_4274);
or U4405 (N_4405,N_4391,N_4321);
or U4406 (N_4406,N_4354,N_4245);
nor U4407 (N_4407,N_4214,N_4235);
and U4408 (N_4408,N_4343,N_4281);
nand U4409 (N_4409,N_4257,N_4250);
nand U4410 (N_4410,N_4320,N_4225);
nand U4411 (N_4411,N_4284,N_4350);
and U4412 (N_4412,N_4337,N_4330);
and U4413 (N_4413,N_4290,N_4241);
xnor U4414 (N_4414,N_4385,N_4226);
xor U4415 (N_4415,N_4348,N_4342);
or U4416 (N_4416,N_4353,N_4355);
or U4417 (N_4417,N_4389,N_4302);
nor U4418 (N_4418,N_4288,N_4307);
and U4419 (N_4419,N_4292,N_4278);
or U4420 (N_4420,N_4206,N_4397);
nand U4421 (N_4421,N_4242,N_4224);
nor U4422 (N_4422,N_4393,N_4314);
and U4423 (N_4423,N_4269,N_4279);
xnor U4424 (N_4424,N_4373,N_4251);
nand U4425 (N_4425,N_4211,N_4253);
nand U4426 (N_4426,N_4255,N_4243);
xor U4427 (N_4427,N_4358,N_4240);
nand U4428 (N_4428,N_4227,N_4249);
xnor U4429 (N_4429,N_4297,N_4212);
or U4430 (N_4430,N_4230,N_4305);
nor U4431 (N_4431,N_4306,N_4380);
nand U4432 (N_4432,N_4232,N_4247);
and U4433 (N_4433,N_4272,N_4362);
xor U4434 (N_4434,N_4387,N_4287);
and U4435 (N_4435,N_4339,N_4392);
nor U4436 (N_4436,N_4293,N_4333);
and U4437 (N_4437,N_4361,N_4219);
nand U4438 (N_4438,N_4216,N_4218);
and U4439 (N_4439,N_4283,N_4369);
nand U4440 (N_4440,N_4220,N_4398);
nand U4441 (N_4441,N_4329,N_4202);
nand U4442 (N_4442,N_4357,N_4322);
xnor U4443 (N_4443,N_4261,N_4285);
nand U4444 (N_4444,N_4208,N_4396);
and U4445 (N_4445,N_4395,N_4324);
nor U4446 (N_4446,N_4221,N_4296);
nor U4447 (N_4447,N_4325,N_4205);
xor U4448 (N_4448,N_4256,N_4248);
or U4449 (N_4449,N_4377,N_4271);
xnor U4450 (N_4450,N_4335,N_4338);
nand U4451 (N_4451,N_4258,N_4229);
and U4452 (N_4452,N_4310,N_4349);
or U4453 (N_4453,N_4375,N_4363);
and U4454 (N_4454,N_4352,N_4323);
xnor U4455 (N_4455,N_4317,N_4301);
or U4456 (N_4456,N_4328,N_4234);
and U4457 (N_4457,N_4201,N_4351);
nand U4458 (N_4458,N_4200,N_4259);
nor U4459 (N_4459,N_4318,N_4376);
nand U4460 (N_4460,N_4346,N_4370);
nand U4461 (N_4461,N_4267,N_4347);
nand U4462 (N_4462,N_4217,N_4238);
nand U4463 (N_4463,N_4304,N_4336);
or U4464 (N_4464,N_4378,N_4244);
and U4465 (N_4465,N_4366,N_4308);
or U4466 (N_4466,N_4311,N_4231);
or U4467 (N_4467,N_4309,N_4289);
and U4468 (N_4468,N_4359,N_4332);
or U4469 (N_4469,N_4237,N_4294);
xor U4470 (N_4470,N_4273,N_4327);
or U4471 (N_4471,N_4312,N_4295);
xnor U4472 (N_4472,N_4254,N_4364);
xor U4473 (N_4473,N_4233,N_4239);
or U4474 (N_4474,N_4210,N_4344);
and U4475 (N_4475,N_4207,N_4213);
and U4476 (N_4476,N_4326,N_4381);
or U4477 (N_4477,N_4264,N_4223);
and U4478 (N_4478,N_4286,N_4372);
nand U4479 (N_4479,N_4368,N_4356);
and U4480 (N_4480,N_4334,N_4331);
nor U4481 (N_4481,N_4300,N_4371);
nand U4482 (N_4482,N_4236,N_4263);
and U4483 (N_4483,N_4276,N_4374);
nand U4484 (N_4484,N_4298,N_4367);
or U4485 (N_4485,N_4291,N_4386);
nand U4486 (N_4486,N_4388,N_4303);
or U4487 (N_4487,N_4275,N_4382);
nor U4488 (N_4488,N_4215,N_4394);
and U4489 (N_4489,N_4262,N_4379);
or U4490 (N_4490,N_4319,N_4384);
and U4491 (N_4491,N_4266,N_4222);
xnor U4492 (N_4492,N_4265,N_4390);
or U4493 (N_4493,N_4252,N_4399);
or U4494 (N_4494,N_4365,N_4209);
xor U4495 (N_4495,N_4203,N_4268);
nor U4496 (N_4496,N_4277,N_4340);
or U4497 (N_4497,N_4280,N_4360);
or U4498 (N_4498,N_4383,N_4228);
nor U4499 (N_4499,N_4345,N_4260);
nor U4500 (N_4500,N_4200,N_4231);
xor U4501 (N_4501,N_4389,N_4258);
nand U4502 (N_4502,N_4263,N_4217);
xor U4503 (N_4503,N_4333,N_4281);
nand U4504 (N_4504,N_4265,N_4369);
nand U4505 (N_4505,N_4215,N_4278);
or U4506 (N_4506,N_4204,N_4328);
nand U4507 (N_4507,N_4329,N_4272);
nor U4508 (N_4508,N_4367,N_4221);
and U4509 (N_4509,N_4234,N_4240);
nand U4510 (N_4510,N_4242,N_4395);
nor U4511 (N_4511,N_4334,N_4200);
or U4512 (N_4512,N_4220,N_4291);
nor U4513 (N_4513,N_4302,N_4354);
or U4514 (N_4514,N_4370,N_4309);
and U4515 (N_4515,N_4232,N_4255);
nor U4516 (N_4516,N_4319,N_4275);
xor U4517 (N_4517,N_4222,N_4277);
or U4518 (N_4518,N_4326,N_4214);
xor U4519 (N_4519,N_4226,N_4399);
nor U4520 (N_4520,N_4287,N_4252);
xnor U4521 (N_4521,N_4388,N_4217);
or U4522 (N_4522,N_4311,N_4393);
or U4523 (N_4523,N_4363,N_4297);
nand U4524 (N_4524,N_4259,N_4333);
xor U4525 (N_4525,N_4275,N_4301);
xor U4526 (N_4526,N_4217,N_4360);
and U4527 (N_4527,N_4346,N_4390);
and U4528 (N_4528,N_4209,N_4223);
nand U4529 (N_4529,N_4250,N_4354);
xor U4530 (N_4530,N_4281,N_4325);
nand U4531 (N_4531,N_4256,N_4249);
nor U4532 (N_4532,N_4282,N_4356);
nand U4533 (N_4533,N_4306,N_4333);
or U4534 (N_4534,N_4247,N_4212);
xor U4535 (N_4535,N_4201,N_4368);
nor U4536 (N_4536,N_4280,N_4289);
or U4537 (N_4537,N_4225,N_4355);
nand U4538 (N_4538,N_4208,N_4339);
nor U4539 (N_4539,N_4272,N_4269);
and U4540 (N_4540,N_4282,N_4236);
and U4541 (N_4541,N_4330,N_4338);
nor U4542 (N_4542,N_4323,N_4328);
or U4543 (N_4543,N_4298,N_4365);
nor U4544 (N_4544,N_4280,N_4226);
nand U4545 (N_4545,N_4340,N_4314);
nand U4546 (N_4546,N_4244,N_4230);
nor U4547 (N_4547,N_4271,N_4204);
nand U4548 (N_4548,N_4337,N_4242);
or U4549 (N_4549,N_4209,N_4299);
xor U4550 (N_4550,N_4258,N_4356);
and U4551 (N_4551,N_4285,N_4343);
nand U4552 (N_4552,N_4365,N_4255);
xnor U4553 (N_4553,N_4339,N_4299);
nor U4554 (N_4554,N_4300,N_4327);
nor U4555 (N_4555,N_4229,N_4374);
or U4556 (N_4556,N_4305,N_4285);
nand U4557 (N_4557,N_4300,N_4324);
or U4558 (N_4558,N_4248,N_4295);
or U4559 (N_4559,N_4280,N_4208);
and U4560 (N_4560,N_4351,N_4258);
or U4561 (N_4561,N_4289,N_4285);
nor U4562 (N_4562,N_4219,N_4342);
and U4563 (N_4563,N_4389,N_4230);
xor U4564 (N_4564,N_4273,N_4320);
and U4565 (N_4565,N_4362,N_4342);
nor U4566 (N_4566,N_4271,N_4292);
and U4567 (N_4567,N_4337,N_4237);
and U4568 (N_4568,N_4226,N_4225);
nor U4569 (N_4569,N_4289,N_4206);
or U4570 (N_4570,N_4239,N_4305);
xnor U4571 (N_4571,N_4234,N_4363);
nand U4572 (N_4572,N_4300,N_4345);
or U4573 (N_4573,N_4227,N_4210);
and U4574 (N_4574,N_4273,N_4333);
nand U4575 (N_4575,N_4284,N_4269);
and U4576 (N_4576,N_4218,N_4367);
nor U4577 (N_4577,N_4367,N_4232);
xor U4578 (N_4578,N_4360,N_4283);
nand U4579 (N_4579,N_4380,N_4254);
nand U4580 (N_4580,N_4286,N_4316);
xnor U4581 (N_4581,N_4253,N_4378);
nor U4582 (N_4582,N_4218,N_4206);
xnor U4583 (N_4583,N_4239,N_4329);
xnor U4584 (N_4584,N_4363,N_4373);
xor U4585 (N_4585,N_4238,N_4391);
nand U4586 (N_4586,N_4207,N_4272);
nor U4587 (N_4587,N_4290,N_4302);
nor U4588 (N_4588,N_4334,N_4381);
or U4589 (N_4589,N_4389,N_4375);
nor U4590 (N_4590,N_4368,N_4390);
and U4591 (N_4591,N_4320,N_4242);
and U4592 (N_4592,N_4287,N_4212);
nand U4593 (N_4593,N_4273,N_4233);
and U4594 (N_4594,N_4259,N_4215);
xor U4595 (N_4595,N_4337,N_4384);
nor U4596 (N_4596,N_4339,N_4330);
nor U4597 (N_4597,N_4200,N_4387);
or U4598 (N_4598,N_4357,N_4293);
and U4599 (N_4599,N_4342,N_4202);
and U4600 (N_4600,N_4583,N_4525);
or U4601 (N_4601,N_4575,N_4424);
nor U4602 (N_4602,N_4568,N_4482);
and U4603 (N_4603,N_4426,N_4570);
xor U4604 (N_4604,N_4534,N_4449);
nand U4605 (N_4605,N_4517,N_4579);
nor U4606 (N_4606,N_4454,N_4413);
xnor U4607 (N_4607,N_4436,N_4523);
nor U4608 (N_4608,N_4421,N_4505);
nor U4609 (N_4609,N_4492,N_4455);
or U4610 (N_4610,N_4567,N_4537);
xor U4611 (N_4611,N_4539,N_4582);
nand U4612 (N_4612,N_4440,N_4469);
xor U4613 (N_4613,N_4559,N_4589);
xor U4614 (N_4614,N_4437,N_4414);
nor U4615 (N_4615,N_4562,N_4401);
or U4616 (N_4616,N_4466,N_4553);
xor U4617 (N_4617,N_4485,N_4410);
nand U4618 (N_4618,N_4576,N_4544);
and U4619 (N_4619,N_4591,N_4462);
or U4620 (N_4620,N_4503,N_4425);
xor U4621 (N_4621,N_4404,N_4422);
and U4622 (N_4622,N_4402,N_4484);
and U4623 (N_4623,N_4555,N_4581);
xor U4624 (N_4624,N_4416,N_4545);
xor U4625 (N_4625,N_4486,N_4442);
xor U4626 (N_4626,N_4467,N_4471);
or U4627 (N_4627,N_4557,N_4594);
and U4628 (N_4628,N_4536,N_4490);
xnor U4629 (N_4629,N_4580,N_4513);
and U4630 (N_4630,N_4558,N_4461);
nand U4631 (N_4631,N_4538,N_4499);
nand U4632 (N_4632,N_4574,N_4596);
nand U4633 (N_4633,N_4542,N_4412);
xnor U4634 (N_4634,N_4464,N_4566);
or U4635 (N_4635,N_4527,N_4405);
xnor U4636 (N_4636,N_4551,N_4514);
or U4637 (N_4637,N_4474,N_4428);
nand U4638 (N_4638,N_4586,N_4500);
nand U4639 (N_4639,N_4494,N_4451);
or U4640 (N_4640,N_4577,N_4479);
nor U4641 (N_4641,N_4434,N_4445);
xnor U4642 (N_4642,N_4460,N_4560);
and U4643 (N_4643,N_4430,N_4590);
nor U4644 (N_4644,N_4521,N_4403);
or U4645 (N_4645,N_4483,N_4417);
or U4646 (N_4646,N_4497,N_4443);
nor U4647 (N_4647,N_4592,N_4532);
nand U4648 (N_4648,N_4510,N_4515);
xor U4649 (N_4649,N_4447,N_4495);
or U4650 (N_4650,N_4456,N_4465);
xor U4651 (N_4651,N_4524,N_4535);
and U4652 (N_4652,N_4491,N_4473);
nor U4653 (N_4653,N_4530,N_4593);
and U4654 (N_4654,N_4458,N_4477);
nand U4655 (N_4655,N_4438,N_4439);
and U4656 (N_4656,N_4498,N_4502);
nand U4657 (N_4657,N_4441,N_4541);
nor U4658 (N_4658,N_4506,N_4470);
or U4659 (N_4659,N_4533,N_4457);
nor U4660 (N_4660,N_4420,N_4585);
xnor U4661 (N_4661,N_4411,N_4598);
xor U4662 (N_4662,N_4432,N_4406);
and U4663 (N_4663,N_4597,N_4540);
or U4664 (N_4664,N_4529,N_4407);
nor U4665 (N_4665,N_4400,N_4468);
nand U4666 (N_4666,N_4507,N_4423);
xnor U4667 (N_4667,N_4599,N_4409);
xor U4668 (N_4668,N_4552,N_4475);
or U4669 (N_4669,N_4584,N_4565);
nand U4670 (N_4670,N_4526,N_4549);
or U4671 (N_4671,N_4450,N_4446);
and U4672 (N_4672,N_4516,N_4550);
xnor U4673 (N_4673,N_4543,N_4419);
xnor U4674 (N_4674,N_4427,N_4587);
nor U4675 (N_4675,N_4429,N_4472);
or U4676 (N_4676,N_4573,N_4488);
or U4677 (N_4677,N_4481,N_4548);
nor U4678 (N_4678,N_4556,N_4435);
nor U4679 (N_4679,N_4563,N_4431);
or U4680 (N_4680,N_4519,N_4588);
nor U4681 (N_4681,N_4453,N_4554);
and U4682 (N_4682,N_4578,N_4511);
or U4683 (N_4683,N_4408,N_4520);
nand U4684 (N_4684,N_4569,N_4509);
nor U4685 (N_4685,N_4433,N_4489);
and U4686 (N_4686,N_4463,N_4487);
nor U4687 (N_4687,N_4459,N_4528);
xnor U4688 (N_4688,N_4448,N_4415);
nor U4689 (N_4689,N_4444,N_4418);
xor U4690 (N_4690,N_4518,N_4476);
and U4691 (N_4691,N_4504,N_4522);
nand U4692 (N_4692,N_4547,N_4452);
nor U4693 (N_4693,N_4478,N_4531);
nand U4694 (N_4694,N_4496,N_4571);
or U4695 (N_4695,N_4595,N_4564);
nor U4696 (N_4696,N_4546,N_4512);
nand U4697 (N_4697,N_4572,N_4508);
or U4698 (N_4698,N_4480,N_4501);
nor U4699 (N_4699,N_4493,N_4561);
nor U4700 (N_4700,N_4525,N_4523);
nand U4701 (N_4701,N_4560,N_4489);
and U4702 (N_4702,N_4595,N_4438);
and U4703 (N_4703,N_4427,N_4578);
xor U4704 (N_4704,N_4485,N_4518);
and U4705 (N_4705,N_4428,N_4439);
and U4706 (N_4706,N_4416,N_4490);
or U4707 (N_4707,N_4507,N_4464);
or U4708 (N_4708,N_4510,N_4406);
xnor U4709 (N_4709,N_4466,N_4519);
and U4710 (N_4710,N_4529,N_4421);
nor U4711 (N_4711,N_4483,N_4471);
and U4712 (N_4712,N_4445,N_4484);
xnor U4713 (N_4713,N_4438,N_4521);
nand U4714 (N_4714,N_4464,N_4527);
and U4715 (N_4715,N_4532,N_4499);
xnor U4716 (N_4716,N_4543,N_4526);
nand U4717 (N_4717,N_4419,N_4533);
or U4718 (N_4718,N_4479,N_4444);
and U4719 (N_4719,N_4499,N_4588);
nand U4720 (N_4720,N_4456,N_4458);
or U4721 (N_4721,N_4544,N_4593);
or U4722 (N_4722,N_4595,N_4597);
nor U4723 (N_4723,N_4597,N_4523);
xnor U4724 (N_4724,N_4523,N_4537);
and U4725 (N_4725,N_4593,N_4466);
xnor U4726 (N_4726,N_4450,N_4456);
and U4727 (N_4727,N_4543,N_4570);
nor U4728 (N_4728,N_4562,N_4532);
nor U4729 (N_4729,N_4483,N_4459);
nor U4730 (N_4730,N_4402,N_4529);
and U4731 (N_4731,N_4401,N_4523);
and U4732 (N_4732,N_4413,N_4557);
or U4733 (N_4733,N_4518,N_4498);
xor U4734 (N_4734,N_4542,N_4467);
nand U4735 (N_4735,N_4468,N_4552);
nor U4736 (N_4736,N_4433,N_4586);
xor U4737 (N_4737,N_4543,N_4584);
nor U4738 (N_4738,N_4476,N_4462);
xnor U4739 (N_4739,N_4459,N_4553);
nand U4740 (N_4740,N_4423,N_4471);
nor U4741 (N_4741,N_4518,N_4488);
nand U4742 (N_4742,N_4497,N_4466);
nand U4743 (N_4743,N_4439,N_4492);
nor U4744 (N_4744,N_4506,N_4405);
or U4745 (N_4745,N_4435,N_4495);
and U4746 (N_4746,N_4467,N_4421);
and U4747 (N_4747,N_4491,N_4472);
nand U4748 (N_4748,N_4413,N_4499);
nor U4749 (N_4749,N_4521,N_4542);
and U4750 (N_4750,N_4409,N_4426);
nor U4751 (N_4751,N_4569,N_4536);
nand U4752 (N_4752,N_4560,N_4459);
nand U4753 (N_4753,N_4470,N_4474);
xor U4754 (N_4754,N_4472,N_4496);
or U4755 (N_4755,N_4577,N_4419);
xor U4756 (N_4756,N_4514,N_4588);
nand U4757 (N_4757,N_4498,N_4411);
or U4758 (N_4758,N_4413,N_4417);
xor U4759 (N_4759,N_4504,N_4590);
nand U4760 (N_4760,N_4584,N_4476);
nor U4761 (N_4761,N_4468,N_4466);
and U4762 (N_4762,N_4508,N_4434);
xor U4763 (N_4763,N_4449,N_4554);
nor U4764 (N_4764,N_4421,N_4587);
or U4765 (N_4765,N_4575,N_4550);
or U4766 (N_4766,N_4446,N_4547);
nor U4767 (N_4767,N_4452,N_4473);
nand U4768 (N_4768,N_4457,N_4407);
and U4769 (N_4769,N_4567,N_4594);
nand U4770 (N_4770,N_4447,N_4511);
or U4771 (N_4771,N_4502,N_4552);
or U4772 (N_4772,N_4595,N_4462);
nor U4773 (N_4773,N_4486,N_4449);
nand U4774 (N_4774,N_4584,N_4448);
nand U4775 (N_4775,N_4431,N_4547);
or U4776 (N_4776,N_4536,N_4542);
or U4777 (N_4777,N_4429,N_4496);
nand U4778 (N_4778,N_4598,N_4506);
xnor U4779 (N_4779,N_4428,N_4497);
xor U4780 (N_4780,N_4509,N_4480);
nor U4781 (N_4781,N_4516,N_4565);
or U4782 (N_4782,N_4594,N_4463);
nor U4783 (N_4783,N_4477,N_4506);
or U4784 (N_4784,N_4531,N_4445);
nor U4785 (N_4785,N_4449,N_4445);
nand U4786 (N_4786,N_4402,N_4403);
and U4787 (N_4787,N_4437,N_4586);
and U4788 (N_4788,N_4597,N_4485);
or U4789 (N_4789,N_4496,N_4503);
nand U4790 (N_4790,N_4418,N_4516);
nand U4791 (N_4791,N_4582,N_4543);
nor U4792 (N_4792,N_4583,N_4593);
nand U4793 (N_4793,N_4482,N_4486);
nor U4794 (N_4794,N_4465,N_4571);
and U4795 (N_4795,N_4567,N_4441);
or U4796 (N_4796,N_4467,N_4509);
xor U4797 (N_4797,N_4487,N_4446);
or U4798 (N_4798,N_4577,N_4593);
nand U4799 (N_4799,N_4438,N_4483);
xor U4800 (N_4800,N_4622,N_4621);
nand U4801 (N_4801,N_4674,N_4708);
nor U4802 (N_4802,N_4721,N_4773);
and U4803 (N_4803,N_4660,N_4691);
nand U4804 (N_4804,N_4764,N_4612);
xor U4805 (N_4805,N_4702,N_4781);
nor U4806 (N_4806,N_4700,N_4745);
xnor U4807 (N_4807,N_4690,N_4620);
xor U4808 (N_4808,N_4667,N_4775);
nor U4809 (N_4809,N_4607,N_4625);
xor U4810 (N_4810,N_4614,N_4705);
and U4811 (N_4811,N_4756,N_4635);
and U4812 (N_4812,N_4684,N_4780);
nand U4813 (N_4813,N_4662,N_4728);
xor U4814 (N_4814,N_4740,N_4623);
and U4815 (N_4815,N_4743,N_4730);
nor U4816 (N_4816,N_4799,N_4676);
xor U4817 (N_4817,N_4718,N_4641);
or U4818 (N_4818,N_4712,N_4693);
xnor U4819 (N_4819,N_4634,N_4654);
or U4820 (N_4820,N_4703,N_4771);
xnor U4821 (N_4821,N_4772,N_4608);
xor U4822 (N_4822,N_4639,N_4670);
xor U4823 (N_4823,N_4637,N_4646);
xor U4824 (N_4824,N_4661,N_4701);
or U4825 (N_4825,N_4733,N_4704);
or U4826 (N_4826,N_4784,N_4659);
nand U4827 (N_4827,N_4707,N_4752);
and U4828 (N_4828,N_4663,N_4672);
and U4829 (N_4829,N_4600,N_4717);
or U4830 (N_4830,N_4782,N_4619);
nand U4831 (N_4831,N_4658,N_4769);
xor U4832 (N_4832,N_4793,N_4795);
and U4833 (N_4833,N_4748,N_4741);
or U4834 (N_4834,N_4631,N_4759);
or U4835 (N_4835,N_4651,N_4636);
or U4836 (N_4836,N_4779,N_4706);
nand U4837 (N_4837,N_4618,N_4605);
nor U4838 (N_4838,N_4650,N_4649);
and U4839 (N_4839,N_4739,N_4669);
nor U4840 (N_4840,N_4736,N_4754);
nand U4841 (N_4841,N_4794,N_4768);
nand U4842 (N_4842,N_4760,N_4688);
nand U4843 (N_4843,N_4642,N_4766);
nor U4844 (N_4844,N_4626,N_4722);
or U4845 (N_4845,N_4729,N_4763);
or U4846 (N_4846,N_4778,N_4777);
xnor U4847 (N_4847,N_4624,N_4603);
or U4848 (N_4848,N_4644,N_4652);
nand U4849 (N_4849,N_4696,N_4668);
xnor U4850 (N_4850,N_4720,N_4665);
nor U4851 (N_4851,N_4744,N_4711);
nand U4852 (N_4852,N_4742,N_4755);
or U4853 (N_4853,N_4750,N_4798);
nor U4854 (N_4854,N_4695,N_4689);
or U4855 (N_4855,N_4627,N_4757);
or U4856 (N_4856,N_4666,N_4792);
xor U4857 (N_4857,N_4762,N_4789);
or U4858 (N_4858,N_4685,N_4602);
xor U4859 (N_4859,N_4783,N_4664);
or U4860 (N_4860,N_4682,N_4675);
or U4861 (N_4861,N_4606,N_4788);
and U4862 (N_4862,N_4692,N_4681);
xnor U4863 (N_4863,N_4648,N_4785);
nor U4864 (N_4864,N_4796,N_4791);
nand U4865 (N_4865,N_4677,N_4776);
and U4866 (N_4866,N_4610,N_4719);
nor U4867 (N_4867,N_4679,N_4671);
nor U4868 (N_4868,N_4632,N_4633);
nand U4869 (N_4869,N_4687,N_4656);
nand U4870 (N_4870,N_4774,N_4604);
xnor U4871 (N_4871,N_4797,N_4725);
or U4872 (N_4872,N_4727,N_4724);
and U4873 (N_4873,N_4761,N_4680);
nand U4874 (N_4874,N_4735,N_4749);
or U4875 (N_4875,N_4616,N_4787);
or U4876 (N_4876,N_4726,N_4697);
nand U4877 (N_4877,N_4638,N_4790);
xor U4878 (N_4878,N_4732,N_4655);
and U4879 (N_4879,N_4628,N_4715);
nor U4880 (N_4880,N_4734,N_4710);
or U4881 (N_4881,N_4678,N_4694);
nand U4882 (N_4882,N_4673,N_4731);
xor U4883 (N_4883,N_4640,N_4786);
or U4884 (N_4884,N_4758,N_4629);
nor U4885 (N_4885,N_4683,N_4686);
or U4886 (N_4886,N_4747,N_4601);
nor U4887 (N_4887,N_4765,N_4653);
nand U4888 (N_4888,N_4709,N_4738);
and U4889 (N_4889,N_4716,N_4645);
or U4890 (N_4890,N_4737,N_4698);
nand U4891 (N_4891,N_4723,N_4643);
nor U4892 (N_4892,N_4753,N_4699);
and U4893 (N_4893,N_4751,N_4609);
or U4894 (N_4894,N_4746,N_4615);
nor U4895 (N_4895,N_4713,N_4770);
or U4896 (N_4896,N_4617,N_4767);
and U4897 (N_4897,N_4714,N_4613);
nand U4898 (N_4898,N_4647,N_4630);
nand U4899 (N_4899,N_4611,N_4657);
nor U4900 (N_4900,N_4782,N_4715);
xnor U4901 (N_4901,N_4728,N_4775);
or U4902 (N_4902,N_4602,N_4711);
or U4903 (N_4903,N_4736,N_4695);
nand U4904 (N_4904,N_4704,N_4622);
or U4905 (N_4905,N_4775,N_4740);
or U4906 (N_4906,N_4781,N_4771);
xor U4907 (N_4907,N_4694,N_4746);
nand U4908 (N_4908,N_4726,N_4647);
nand U4909 (N_4909,N_4628,N_4658);
nor U4910 (N_4910,N_4780,N_4781);
nor U4911 (N_4911,N_4671,N_4613);
or U4912 (N_4912,N_4780,N_4635);
or U4913 (N_4913,N_4719,N_4725);
nor U4914 (N_4914,N_4742,N_4658);
nor U4915 (N_4915,N_4776,N_4780);
nor U4916 (N_4916,N_4767,N_4786);
nand U4917 (N_4917,N_4701,N_4662);
xor U4918 (N_4918,N_4677,N_4658);
or U4919 (N_4919,N_4624,N_4611);
or U4920 (N_4920,N_4703,N_4770);
xnor U4921 (N_4921,N_4785,N_4759);
nor U4922 (N_4922,N_4776,N_4603);
nand U4923 (N_4923,N_4691,N_4724);
or U4924 (N_4924,N_4664,N_4729);
nand U4925 (N_4925,N_4686,N_4690);
and U4926 (N_4926,N_4640,N_4675);
and U4927 (N_4927,N_4610,N_4770);
xor U4928 (N_4928,N_4641,N_4792);
nand U4929 (N_4929,N_4722,N_4783);
and U4930 (N_4930,N_4691,N_4612);
and U4931 (N_4931,N_4714,N_4650);
or U4932 (N_4932,N_4720,N_4693);
xor U4933 (N_4933,N_4723,N_4703);
nor U4934 (N_4934,N_4670,N_4680);
and U4935 (N_4935,N_4685,N_4625);
or U4936 (N_4936,N_4612,N_4700);
or U4937 (N_4937,N_4789,N_4628);
and U4938 (N_4938,N_4693,N_4715);
xor U4939 (N_4939,N_4720,N_4664);
and U4940 (N_4940,N_4608,N_4719);
xnor U4941 (N_4941,N_4767,N_4687);
nand U4942 (N_4942,N_4753,N_4713);
nor U4943 (N_4943,N_4741,N_4732);
or U4944 (N_4944,N_4713,N_4701);
or U4945 (N_4945,N_4755,N_4734);
or U4946 (N_4946,N_4718,N_4790);
and U4947 (N_4947,N_4786,N_4673);
nand U4948 (N_4948,N_4694,N_4757);
and U4949 (N_4949,N_4629,N_4709);
or U4950 (N_4950,N_4654,N_4675);
or U4951 (N_4951,N_4643,N_4781);
nor U4952 (N_4952,N_4699,N_4654);
nor U4953 (N_4953,N_4610,N_4686);
and U4954 (N_4954,N_4789,N_4761);
nor U4955 (N_4955,N_4699,N_4705);
or U4956 (N_4956,N_4651,N_4630);
nand U4957 (N_4957,N_4657,N_4798);
nand U4958 (N_4958,N_4648,N_4712);
or U4959 (N_4959,N_4793,N_4707);
and U4960 (N_4960,N_4625,N_4774);
nor U4961 (N_4961,N_4690,N_4661);
and U4962 (N_4962,N_4786,N_4717);
and U4963 (N_4963,N_4646,N_4614);
and U4964 (N_4964,N_4788,N_4725);
and U4965 (N_4965,N_4658,N_4770);
and U4966 (N_4966,N_4678,N_4761);
or U4967 (N_4967,N_4782,N_4607);
and U4968 (N_4968,N_4654,N_4624);
and U4969 (N_4969,N_4652,N_4645);
xor U4970 (N_4970,N_4726,N_4721);
nand U4971 (N_4971,N_4642,N_4651);
or U4972 (N_4972,N_4624,N_4695);
nor U4973 (N_4973,N_4741,N_4698);
xnor U4974 (N_4974,N_4651,N_4633);
nor U4975 (N_4975,N_4724,N_4614);
and U4976 (N_4976,N_4678,N_4681);
or U4977 (N_4977,N_4672,N_4760);
or U4978 (N_4978,N_4755,N_4662);
or U4979 (N_4979,N_4681,N_4630);
or U4980 (N_4980,N_4677,N_4720);
nand U4981 (N_4981,N_4749,N_4782);
xor U4982 (N_4982,N_4723,N_4688);
or U4983 (N_4983,N_4704,N_4786);
or U4984 (N_4984,N_4715,N_4732);
xor U4985 (N_4985,N_4666,N_4721);
or U4986 (N_4986,N_4713,N_4724);
nand U4987 (N_4987,N_4737,N_4661);
xor U4988 (N_4988,N_4620,N_4664);
nand U4989 (N_4989,N_4793,N_4666);
nor U4990 (N_4990,N_4715,N_4614);
and U4991 (N_4991,N_4643,N_4691);
nor U4992 (N_4992,N_4636,N_4749);
nor U4993 (N_4993,N_4762,N_4693);
xnor U4994 (N_4994,N_4693,N_4713);
and U4995 (N_4995,N_4756,N_4651);
or U4996 (N_4996,N_4618,N_4798);
nor U4997 (N_4997,N_4649,N_4678);
nand U4998 (N_4998,N_4667,N_4762);
and U4999 (N_4999,N_4757,N_4735);
or U5000 (N_5000,N_4944,N_4813);
nor U5001 (N_5001,N_4865,N_4851);
nand U5002 (N_5002,N_4933,N_4889);
and U5003 (N_5003,N_4970,N_4885);
xnor U5004 (N_5004,N_4913,N_4935);
xor U5005 (N_5005,N_4923,N_4937);
nand U5006 (N_5006,N_4906,N_4819);
or U5007 (N_5007,N_4956,N_4907);
nor U5008 (N_5008,N_4957,N_4862);
nand U5009 (N_5009,N_4940,N_4841);
xor U5010 (N_5010,N_4836,N_4946);
or U5011 (N_5011,N_4883,N_4809);
nand U5012 (N_5012,N_4893,N_4854);
and U5013 (N_5013,N_4942,N_4999);
or U5014 (N_5014,N_4870,N_4860);
or U5015 (N_5015,N_4949,N_4989);
xor U5016 (N_5016,N_4815,N_4924);
or U5017 (N_5017,N_4886,N_4995);
nor U5018 (N_5018,N_4996,N_4805);
nor U5019 (N_5019,N_4961,N_4838);
nand U5020 (N_5020,N_4983,N_4842);
nand U5021 (N_5021,N_4839,N_4824);
and U5022 (N_5022,N_4863,N_4919);
nand U5023 (N_5023,N_4878,N_4954);
xor U5024 (N_5024,N_4834,N_4958);
nor U5025 (N_5025,N_4847,N_4803);
and U5026 (N_5026,N_4908,N_4914);
xor U5027 (N_5027,N_4807,N_4828);
nor U5028 (N_5028,N_4821,N_4825);
or U5029 (N_5029,N_4800,N_4922);
and U5030 (N_5030,N_4855,N_4894);
xnor U5031 (N_5031,N_4829,N_4912);
xnor U5032 (N_5032,N_4977,N_4896);
xor U5033 (N_5033,N_4822,N_4965);
nor U5034 (N_5034,N_4897,N_4837);
nand U5035 (N_5035,N_4917,N_4968);
nand U5036 (N_5036,N_4874,N_4918);
nor U5037 (N_5037,N_4945,N_4895);
nand U5038 (N_5038,N_4812,N_4816);
and U5039 (N_5039,N_4856,N_4926);
and U5040 (N_5040,N_4846,N_4871);
nor U5041 (N_5041,N_4960,N_4869);
nor U5042 (N_5042,N_4879,N_4848);
xnor U5043 (N_5043,N_4963,N_4985);
or U5044 (N_5044,N_4966,N_4941);
or U5045 (N_5045,N_4982,N_4911);
and U5046 (N_5046,N_4801,N_4984);
xnor U5047 (N_5047,N_4810,N_4990);
or U5048 (N_5048,N_4998,N_4868);
nand U5049 (N_5049,N_4902,N_4950);
nand U5050 (N_5050,N_4814,N_4927);
and U5051 (N_5051,N_4844,N_4861);
nand U5052 (N_5052,N_4997,N_4974);
xor U5053 (N_5053,N_4853,N_4887);
nand U5054 (N_5054,N_4951,N_4978);
nand U5055 (N_5055,N_4929,N_4909);
or U5056 (N_5056,N_4811,N_4915);
or U5057 (N_5057,N_4988,N_4955);
or U5058 (N_5058,N_4964,N_4875);
xor U5059 (N_5059,N_4943,N_4882);
xor U5060 (N_5060,N_4872,N_4938);
xor U5061 (N_5061,N_4804,N_4934);
xnor U5062 (N_5062,N_4817,N_4930);
and U5063 (N_5063,N_4858,N_4877);
nand U5064 (N_5064,N_4873,N_4852);
xor U5065 (N_5065,N_4901,N_4962);
and U5066 (N_5066,N_4820,N_4979);
nor U5067 (N_5067,N_4973,N_4802);
nor U5068 (N_5068,N_4859,N_4928);
xor U5069 (N_5069,N_4831,N_4976);
or U5070 (N_5070,N_4864,N_4903);
nand U5071 (N_5071,N_4857,N_4932);
xnor U5072 (N_5072,N_4959,N_4975);
nor U5073 (N_5073,N_4981,N_4818);
nand U5074 (N_5074,N_4840,N_4888);
xnor U5075 (N_5075,N_4920,N_4850);
nand U5076 (N_5076,N_4830,N_4925);
xor U5077 (N_5077,N_4823,N_4884);
or U5078 (N_5078,N_4953,N_4931);
or U5079 (N_5079,N_4904,N_4835);
nor U5080 (N_5080,N_4971,N_4881);
nand U5081 (N_5081,N_4827,N_4900);
and U5082 (N_5082,N_4826,N_4972);
and U5083 (N_5083,N_4892,N_4987);
and U5084 (N_5084,N_4986,N_4980);
nand U5085 (N_5085,N_4994,N_4947);
xor U5086 (N_5086,N_4898,N_4910);
and U5087 (N_5087,N_4866,N_4832);
or U5088 (N_5088,N_4992,N_4921);
xnor U5089 (N_5089,N_4991,N_4891);
or U5090 (N_5090,N_4952,N_4890);
or U5091 (N_5091,N_4833,N_4969);
or U5092 (N_5092,N_4867,N_4936);
xor U5093 (N_5093,N_4808,N_4849);
and U5094 (N_5094,N_4905,N_4876);
xnor U5095 (N_5095,N_4880,N_4845);
or U5096 (N_5096,N_4916,N_4899);
nand U5097 (N_5097,N_4948,N_4967);
nor U5098 (N_5098,N_4843,N_4993);
or U5099 (N_5099,N_4939,N_4806);
nand U5100 (N_5100,N_4845,N_4992);
nor U5101 (N_5101,N_4827,N_4938);
xnor U5102 (N_5102,N_4961,N_4867);
nor U5103 (N_5103,N_4800,N_4872);
xor U5104 (N_5104,N_4972,N_4987);
nor U5105 (N_5105,N_4841,N_4857);
and U5106 (N_5106,N_4840,N_4812);
or U5107 (N_5107,N_4949,N_4937);
xnor U5108 (N_5108,N_4906,N_4957);
and U5109 (N_5109,N_4974,N_4827);
nand U5110 (N_5110,N_4893,N_4957);
or U5111 (N_5111,N_4881,N_4832);
xor U5112 (N_5112,N_4933,N_4915);
and U5113 (N_5113,N_4822,N_4896);
or U5114 (N_5114,N_4916,N_4969);
nand U5115 (N_5115,N_4826,N_4938);
nor U5116 (N_5116,N_4890,N_4958);
and U5117 (N_5117,N_4989,N_4883);
nor U5118 (N_5118,N_4814,N_4884);
nand U5119 (N_5119,N_4974,N_4958);
xor U5120 (N_5120,N_4854,N_4992);
xor U5121 (N_5121,N_4879,N_4916);
nand U5122 (N_5122,N_4819,N_4832);
or U5123 (N_5123,N_4800,N_4828);
and U5124 (N_5124,N_4998,N_4924);
nand U5125 (N_5125,N_4941,N_4965);
nor U5126 (N_5126,N_4840,N_4989);
nor U5127 (N_5127,N_4910,N_4846);
or U5128 (N_5128,N_4910,N_4912);
and U5129 (N_5129,N_4937,N_4830);
or U5130 (N_5130,N_4881,N_4906);
xnor U5131 (N_5131,N_4997,N_4874);
nand U5132 (N_5132,N_4945,N_4956);
xor U5133 (N_5133,N_4997,N_4989);
nand U5134 (N_5134,N_4820,N_4814);
or U5135 (N_5135,N_4878,N_4896);
nor U5136 (N_5136,N_4910,N_4845);
and U5137 (N_5137,N_4846,N_4819);
xor U5138 (N_5138,N_4890,N_4830);
xor U5139 (N_5139,N_4814,N_4980);
xor U5140 (N_5140,N_4925,N_4949);
or U5141 (N_5141,N_4961,N_4898);
and U5142 (N_5142,N_4834,N_4904);
and U5143 (N_5143,N_4955,N_4857);
nand U5144 (N_5144,N_4961,N_4872);
or U5145 (N_5145,N_4897,N_4904);
xnor U5146 (N_5146,N_4978,N_4855);
nand U5147 (N_5147,N_4873,N_4993);
nor U5148 (N_5148,N_4991,N_4841);
xnor U5149 (N_5149,N_4868,N_4838);
or U5150 (N_5150,N_4983,N_4890);
nand U5151 (N_5151,N_4815,N_4958);
and U5152 (N_5152,N_4887,N_4905);
or U5153 (N_5153,N_4916,N_4860);
xnor U5154 (N_5154,N_4942,N_4967);
nor U5155 (N_5155,N_4892,N_4959);
or U5156 (N_5156,N_4904,N_4845);
nand U5157 (N_5157,N_4877,N_4888);
nand U5158 (N_5158,N_4906,N_4965);
xnor U5159 (N_5159,N_4969,N_4876);
or U5160 (N_5160,N_4837,N_4831);
nand U5161 (N_5161,N_4965,N_4902);
and U5162 (N_5162,N_4905,N_4881);
or U5163 (N_5163,N_4954,N_4850);
or U5164 (N_5164,N_4986,N_4935);
nor U5165 (N_5165,N_4942,N_4915);
nor U5166 (N_5166,N_4945,N_4977);
xnor U5167 (N_5167,N_4955,N_4908);
nand U5168 (N_5168,N_4886,N_4820);
nor U5169 (N_5169,N_4843,N_4805);
nand U5170 (N_5170,N_4837,N_4968);
xnor U5171 (N_5171,N_4816,N_4862);
nand U5172 (N_5172,N_4882,N_4803);
nor U5173 (N_5173,N_4991,N_4949);
xnor U5174 (N_5174,N_4844,N_4853);
xor U5175 (N_5175,N_4876,N_4898);
or U5176 (N_5176,N_4979,N_4935);
and U5177 (N_5177,N_4872,N_4815);
nor U5178 (N_5178,N_4926,N_4904);
nor U5179 (N_5179,N_4800,N_4983);
nor U5180 (N_5180,N_4835,N_4939);
and U5181 (N_5181,N_4834,N_4866);
nand U5182 (N_5182,N_4821,N_4845);
nor U5183 (N_5183,N_4937,N_4876);
nand U5184 (N_5184,N_4987,N_4913);
nor U5185 (N_5185,N_4978,N_4986);
nor U5186 (N_5186,N_4962,N_4876);
xnor U5187 (N_5187,N_4892,N_4881);
and U5188 (N_5188,N_4815,N_4921);
xnor U5189 (N_5189,N_4929,N_4891);
nor U5190 (N_5190,N_4944,N_4866);
xnor U5191 (N_5191,N_4885,N_4865);
or U5192 (N_5192,N_4978,N_4980);
or U5193 (N_5193,N_4963,N_4941);
nor U5194 (N_5194,N_4867,N_4999);
xor U5195 (N_5195,N_4889,N_4959);
or U5196 (N_5196,N_4868,N_4804);
or U5197 (N_5197,N_4914,N_4990);
and U5198 (N_5198,N_4972,N_4989);
nand U5199 (N_5199,N_4996,N_4955);
nor U5200 (N_5200,N_5089,N_5103);
or U5201 (N_5201,N_5131,N_5167);
nor U5202 (N_5202,N_5032,N_5122);
nand U5203 (N_5203,N_5008,N_5106);
and U5204 (N_5204,N_5001,N_5196);
nor U5205 (N_5205,N_5178,N_5197);
xor U5206 (N_5206,N_5066,N_5194);
or U5207 (N_5207,N_5003,N_5043);
or U5208 (N_5208,N_5145,N_5171);
xor U5209 (N_5209,N_5024,N_5095);
and U5210 (N_5210,N_5058,N_5198);
and U5211 (N_5211,N_5130,N_5144);
nand U5212 (N_5212,N_5085,N_5162);
or U5213 (N_5213,N_5030,N_5132);
nor U5214 (N_5214,N_5012,N_5160);
xnor U5215 (N_5215,N_5015,N_5137);
nor U5216 (N_5216,N_5011,N_5175);
and U5217 (N_5217,N_5177,N_5061);
nand U5218 (N_5218,N_5000,N_5064);
or U5219 (N_5219,N_5185,N_5101);
nand U5220 (N_5220,N_5051,N_5017);
nor U5221 (N_5221,N_5082,N_5086);
or U5222 (N_5222,N_5195,N_5170);
or U5223 (N_5223,N_5142,N_5045);
nand U5224 (N_5224,N_5046,N_5152);
and U5225 (N_5225,N_5020,N_5121);
or U5226 (N_5226,N_5147,N_5149);
nand U5227 (N_5227,N_5134,N_5191);
and U5228 (N_5228,N_5031,N_5010);
nor U5229 (N_5229,N_5063,N_5146);
nor U5230 (N_5230,N_5019,N_5021);
nand U5231 (N_5231,N_5027,N_5151);
nand U5232 (N_5232,N_5189,N_5156);
and U5233 (N_5233,N_5055,N_5005);
nor U5234 (N_5234,N_5108,N_5068);
or U5235 (N_5235,N_5013,N_5075);
nor U5236 (N_5236,N_5009,N_5093);
xor U5237 (N_5237,N_5157,N_5141);
and U5238 (N_5238,N_5150,N_5173);
nor U5239 (N_5239,N_5098,N_5136);
or U5240 (N_5240,N_5129,N_5067);
nor U5241 (N_5241,N_5099,N_5091);
xor U5242 (N_5242,N_5034,N_5087);
or U5243 (N_5243,N_5125,N_5153);
or U5244 (N_5244,N_5080,N_5081);
xnor U5245 (N_5245,N_5181,N_5065);
nor U5246 (N_5246,N_5036,N_5053);
or U5247 (N_5247,N_5190,N_5154);
nor U5248 (N_5248,N_5140,N_5118);
and U5249 (N_5249,N_5041,N_5114);
and U5250 (N_5250,N_5047,N_5018);
xor U5251 (N_5251,N_5007,N_5022);
nand U5252 (N_5252,N_5113,N_5105);
xor U5253 (N_5253,N_5104,N_5168);
nand U5254 (N_5254,N_5148,N_5123);
xnor U5255 (N_5255,N_5138,N_5038);
or U5256 (N_5256,N_5078,N_5016);
and U5257 (N_5257,N_5143,N_5096);
nand U5258 (N_5258,N_5042,N_5110);
and U5259 (N_5259,N_5112,N_5002);
or U5260 (N_5260,N_5026,N_5193);
xor U5261 (N_5261,N_5062,N_5165);
xor U5262 (N_5262,N_5073,N_5052);
nor U5263 (N_5263,N_5035,N_5180);
or U5264 (N_5264,N_5023,N_5079);
nor U5265 (N_5265,N_5172,N_5128);
or U5266 (N_5266,N_5074,N_5083);
and U5267 (N_5267,N_5159,N_5166);
nand U5268 (N_5268,N_5037,N_5183);
xnor U5269 (N_5269,N_5109,N_5169);
xnor U5270 (N_5270,N_5164,N_5076);
nor U5271 (N_5271,N_5158,N_5033);
or U5272 (N_5272,N_5116,N_5126);
nand U5273 (N_5273,N_5176,N_5072);
nand U5274 (N_5274,N_5025,N_5120);
xnor U5275 (N_5275,N_5028,N_5192);
or U5276 (N_5276,N_5094,N_5100);
and U5277 (N_5277,N_5060,N_5139);
xor U5278 (N_5278,N_5182,N_5050);
and U5279 (N_5279,N_5044,N_5059);
and U5280 (N_5280,N_5187,N_5054);
nor U5281 (N_5281,N_5090,N_5006);
nand U5282 (N_5282,N_5004,N_5039);
or U5283 (N_5283,N_5070,N_5155);
nor U5284 (N_5284,N_5119,N_5014);
or U5285 (N_5285,N_5188,N_5057);
and U5286 (N_5286,N_5029,N_5049);
nand U5287 (N_5287,N_5088,N_5069);
nand U5288 (N_5288,N_5127,N_5117);
nor U5289 (N_5289,N_5071,N_5077);
or U5290 (N_5290,N_5133,N_5097);
xor U5291 (N_5291,N_5048,N_5084);
xor U5292 (N_5292,N_5135,N_5111);
xor U5293 (N_5293,N_5184,N_5199);
nand U5294 (N_5294,N_5179,N_5161);
and U5295 (N_5295,N_5163,N_5107);
nand U5296 (N_5296,N_5092,N_5056);
or U5297 (N_5297,N_5186,N_5174);
nor U5298 (N_5298,N_5124,N_5115);
nor U5299 (N_5299,N_5040,N_5102);
nand U5300 (N_5300,N_5049,N_5195);
or U5301 (N_5301,N_5120,N_5103);
or U5302 (N_5302,N_5152,N_5075);
xnor U5303 (N_5303,N_5124,N_5030);
and U5304 (N_5304,N_5050,N_5179);
nor U5305 (N_5305,N_5136,N_5086);
or U5306 (N_5306,N_5125,N_5136);
xor U5307 (N_5307,N_5091,N_5016);
nand U5308 (N_5308,N_5106,N_5018);
nor U5309 (N_5309,N_5039,N_5178);
nor U5310 (N_5310,N_5126,N_5024);
xor U5311 (N_5311,N_5064,N_5010);
and U5312 (N_5312,N_5187,N_5012);
and U5313 (N_5313,N_5000,N_5105);
or U5314 (N_5314,N_5040,N_5001);
xor U5315 (N_5315,N_5065,N_5093);
nand U5316 (N_5316,N_5121,N_5177);
and U5317 (N_5317,N_5008,N_5074);
and U5318 (N_5318,N_5088,N_5123);
nand U5319 (N_5319,N_5050,N_5133);
nand U5320 (N_5320,N_5137,N_5195);
or U5321 (N_5321,N_5060,N_5128);
xor U5322 (N_5322,N_5037,N_5051);
nand U5323 (N_5323,N_5155,N_5053);
and U5324 (N_5324,N_5100,N_5076);
or U5325 (N_5325,N_5027,N_5141);
or U5326 (N_5326,N_5146,N_5144);
nor U5327 (N_5327,N_5151,N_5078);
and U5328 (N_5328,N_5111,N_5148);
or U5329 (N_5329,N_5192,N_5093);
xor U5330 (N_5330,N_5173,N_5085);
and U5331 (N_5331,N_5122,N_5040);
nor U5332 (N_5332,N_5083,N_5046);
xor U5333 (N_5333,N_5060,N_5002);
xor U5334 (N_5334,N_5085,N_5098);
or U5335 (N_5335,N_5026,N_5188);
nor U5336 (N_5336,N_5164,N_5079);
and U5337 (N_5337,N_5025,N_5075);
and U5338 (N_5338,N_5093,N_5031);
and U5339 (N_5339,N_5045,N_5036);
xor U5340 (N_5340,N_5024,N_5140);
nor U5341 (N_5341,N_5076,N_5002);
xor U5342 (N_5342,N_5070,N_5172);
nor U5343 (N_5343,N_5190,N_5079);
nand U5344 (N_5344,N_5098,N_5084);
or U5345 (N_5345,N_5128,N_5147);
or U5346 (N_5346,N_5040,N_5147);
nor U5347 (N_5347,N_5017,N_5021);
nor U5348 (N_5348,N_5089,N_5191);
nand U5349 (N_5349,N_5099,N_5177);
xnor U5350 (N_5350,N_5072,N_5103);
and U5351 (N_5351,N_5071,N_5156);
nor U5352 (N_5352,N_5160,N_5105);
and U5353 (N_5353,N_5000,N_5189);
xnor U5354 (N_5354,N_5022,N_5087);
xnor U5355 (N_5355,N_5114,N_5190);
xnor U5356 (N_5356,N_5049,N_5165);
nor U5357 (N_5357,N_5146,N_5005);
nor U5358 (N_5358,N_5050,N_5156);
or U5359 (N_5359,N_5077,N_5182);
nand U5360 (N_5360,N_5169,N_5173);
xor U5361 (N_5361,N_5184,N_5051);
nand U5362 (N_5362,N_5089,N_5059);
or U5363 (N_5363,N_5122,N_5022);
or U5364 (N_5364,N_5059,N_5134);
or U5365 (N_5365,N_5012,N_5010);
nand U5366 (N_5366,N_5141,N_5002);
and U5367 (N_5367,N_5197,N_5018);
or U5368 (N_5368,N_5126,N_5101);
and U5369 (N_5369,N_5183,N_5018);
xnor U5370 (N_5370,N_5015,N_5172);
nand U5371 (N_5371,N_5134,N_5142);
or U5372 (N_5372,N_5180,N_5097);
xor U5373 (N_5373,N_5005,N_5188);
and U5374 (N_5374,N_5025,N_5029);
nor U5375 (N_5375,N_5146,N_5168);
nand U5376 (N_5376,N_5151,N_5016);
nand U5377 (N_5377,N_5059,N_5194);
nand U5378 (N_5378,N_5012,N_5150);
or U5379 (N_5379,N_5097,N_5111);
and U5380 (N_5380,N_5003,N_5167);
or U5381 (N_5381,N_5081,N_5084);
nand U5382 (N_5382,N_5175,N_5153);
nor U5383 (N_5383,N_5004,N_5061);
nand U5384 (N_5384,N_5159,N_5054);
and U5385 (N_5385,N_5095,N_5085);
nand U5386 (N_5386,N_5002,N_5134);
and U5387 (N_5387,N_5111,N_5062);
nand U5388 (N_5388,N_5155,N_5182);
and U5389 (N_5389,N_5048,N_5147);
and U5390 (N_5390,N_5147,N_5186);
nand U5391 (N_5391,N_5138,N_5121);
and U5392 (N_5392,N_5081,N_5045);
nor U5393 (N_5393,N_5008,N_5156);
nand U5394 (N_5394,N_5102,N_5133);
nor U5395 (N_5395,N_5185,N_5143);
xor U5396 (N_5396,N_5009,N_5118);
nand U5397 (N_5397,N_5007,N_5138);
xnor U5398 (N_5398,N_5119,N_5128);
nor U5399 (N_5399,N_5026,N_5028);
nand U5400 (N_5400,N_5234,N_5201);
xor U5401 (N_5401,N_5393,N_5240);
and U5402 (N_5402,N_5395,N_5295);
nor U5403 (N_5403,N_5398,N_5223);
nand U5404 (N_5404,N_5308,N_5213);
xnor U5405 (N_5405,N_5274,N_5389);
and U5406 (N_5406,N_5363,N_5376);
nor U5407 (N_5407,N_5337,N_5267);
xnor U5408 (N_5408,N_5345,N_5277);
or U5409 (N_5409,N_5280,N_5303);
xnor U5410 (N_5410,N_5388,N_5276);
and U5411 (N_5411,N_5379,N_5352);
and U5412 (N_5412,N_5243,N_5265);
xor U5413 (N_5413,N_5377,N_5219);
xor U5414 (N_5414,N_5296,N_5231);
xor U5415 (N_5415,N_5206,N_5214);
or U5416 (N_5416,N_5285,N_5220);
or U5417 (N_5417,N_5210,N_5362);
nand U5418 (N_5418,N_5329,N_5305);
and U5419 (N_5419,N_5390,N_5326);
nand U5420 (N_5420,N_5289,N_5358);
and U5421 (N_5421,N_5324,N_5271);
and U5422 (N_5422,N_5347,N_5331);
or U5423 (N_5423,N_5317,N_5222);
nor U5424 (N_5424,N_5349,N_5361);
xnor U5425 (N_5425,N_5301,N_5269);
or U5426 (N_5426,N_5380,N_5279);
xor U5427 (N_5427,N_5391,N_5228);
and U5428 (N_5428,N_5300,N_5351);
and U5429 (N_5429,N_5216,N_5330);
xnor U5430 (N_5430,N_5310,N_5292);
nand U5431 (N_5431,N_5397,N_5212);
and U5432 (N_5432,N_5350,N_5282);
nand U5433 (N_5433,N_5266,N_5281);
or U5434 (N_5434,N_5375,N_5316);
nor U5435 (N_5435,N_5236,N_5215);
or U5436 (N_5436,N_5381,N_5251);
nor U5437 (N_5437,N_5286,N_5354);
xnor U5438 (N_5438,N_5370,N_5338);
nor U5439 (N_5439,N_5378,N_5200);
or U5440 (N_5440,N_5257,N_5204);
and U5441 (N_5441,N_5217,N_5203);
and U5442 (N_5442,N_5304,N_5253);
xnor U5443 (N_5443,N_5270,N_5360);
or U5444 (N_5444,N_5320,N_5208);
and U5445 (N_5445,N_5278,N_5318);
or U5446 (N_5446,N_5374,N_5205);
xnor U5447 (N_5447,N_5249,N_5259);
nor U5448 (N_5448,N_5335,N_5365);
nor U5449 (N_5449,N_5252,N_5235);
and U5450 (N_5450,N_5342,N_5294);
nand U5451 (N_5451,N_5384,N_5232);
or U5452 (N_5452,N_5260,N_5230);
or U5453 (N_5453,N_5315,N_5328);
xor U5454 (N_5454,N_5334,N_5207);
and U5455 (N_5455,N_5211,N_5356);
xnor U5456 (N_5456,N_5246,N_5233);
and U5457 (N_5457,N_5238,N_5254);
nand U5458 (N_5458,N_5226,N_5367);
or U5459 (N_5459,N_5255,N_5312);
xnor U5460 (N_5460,N_5344,N_5307);
nor U5461 (N_5461,N_5290,N_5359);
xnor U5462 (N_5462,N_5373,N_5272);
or U5463 (N_5463,N_5386,N_5298);
or U5464 (N_5464,N_5250,N_5218);
nor U5465 (N_5465,N_5268,N_5368);
nand U5466 (N_5466,N_5369,N_5262);
nor U5467 (N_5467,N_5242,N_5340);
nor U5468 (N_5468,N_5396,N_5288);
or U5469 (N_5469,N_5364,N_5371);
nand U5470 (N_5470,N_5264,N_5322);
nand U5471 (N_5471,N_5333,N_5311);
nor U5472 (N_5472,N_5383,N_5357);
xnor U5473 (N_5473,N_5392,N_5323);
nand U5474 (N_5474,N_5343,N_5327);
and U5475 (N_5475,N_5224,N_5385);
xor U5476 (N_5476,N_5245,N_5399);
and U5477 (N_5477,N_5309,N_5202);
or U5478 (N_5478,N_5348,N_5325);
nor U5479 (N_5479,N_5244,N_5248);
and U5480 (N_5480,N_5256,N_5332);
and U5481 (N_5481,N_5275,N_5341);
xor U5482 (N_5482,N_5355,N_5319);
or U5483 (N_5483,N_5306,N_5263);
nor U5484 (N_5484,N_5394,N_5258);
and U5485 (N_5485,N_5239,N_5241);
nor U5486 (N_5486,N_5293,N_5209);
xnor U5487 (N_5487,N_5321,N_5299);
nand U5488 (N_5488,N_5261,N_5302);
nand U5489 (N_5489,N_5346,N_5382);
or U5490 (N_5490,N_5353,N_5336);
or U5491 (N_5491,N_5284,N_5229);
and U5492 (N_5492,N_5227,N_5221);
nor U5493 (N_5493,N_5291,N_5387);
nor U5494 (N_5494,N_5247,N_5237);
xnor U5495 (N_5495,N_5287,N_5273);
xor U5496 (N_5496,N_5283,N_5366);
and U5497 (N_5497,N_5313,N_5314);
nand U5498 (N_5498,N_5225,N_5372);
nor U5499 (N_5499,N_5297,N_5339);
nand U5500 (N_5500,N_5396,N_5256);
and U5501 (N_5501,N_5396,N_5287);
nand U5502 (N_5502,N_5298,N_5365);
and U5503 (N_5503,N_5287,N_5288);
and U5504 (N_5504,N_5324,N_5351);
nand U5505 (N_5505,N_5297,N_5361);
and U5506 (N_5506,N_5299,N_5351);
xor U5507 (N_5507,N_5277,N_5335);
nor U5508 (N_5508,N_5236,N_5342);
or U5509 (N_5509,N_5315,N_5398);
nor U5510 (N_5510,N_5377,N_5207);
and U5511 (N_5511,N_5329,N_5295);
xnor U5512 (N_5512,N_5369,N_5286);
nand U5513 (N_5513,N_5296,N_5271);
nand U5514 (N_5514,N_5324,N_5347);
or U5515 (N_5515,N_5359,N_5292);
and U5516 (N_5516,N_5226,N_5223);
or U5517 (N_5517,N_5379,N_5201);
nor U5518 (N_5518,N_5397,N_5346);
and U5519 (N_5519,N_5373,N_5225);
and U5520 (N_5520,N_5215,N_5287);
xnor U5521 (N_5521,N_5289,N_5297);
nand U5522 (N_5522,N_5389,N_5325);
or U5523 (N_5523,N_5244,N_5339);
and U5524 (N_5524,N_5342,N_5293);
or U5525 (N_5525,N_5257,N_5374);
nand U5526 (N_5526,N_5253,N_5333);
or U5527 (N_5527,N_5230,N_5239);
nor U5528 (N_5528,N_5268,N_5302);
or U5529 (N_5529,N_5227,N_5386);
and U5530 (N_5530,N_5290,N_5258);
or U5531 (N_5531,N_5291,N_5219);
and U5532 (N_5532,N_5320,N_5383);
and U5533 (N_5533,N_5328,N_5336);
or U5534 (N_5534,N_5260,N_5343);
nor U5535 (N_5535,N_5331,N_5375);
nor U5536 (N_5536,N_5309,N_5386);
xnor U5537 (N_5537,N_5217,N_5312);
xnor U5538 (N_5538,N_5317,N_5273);
nor U5539 (N_5539,N_5320,N_5248);
nor U5540 (N_5540,N_5301,N_5342);
nor U5541 (N_5541,N_5231,N_5214);
or U5542 (N_5542,N_5317,N_5358);
xnor U5543 (N_5543,N_5306,N_5359);
and U5544 (N_5544,N_5272,N_5326);
xnor U5545 (N_5545,N_5365,N_5218);
nand U5546 (N_5546,N_5240,N_5315);
and U5547 (N_5547,N_5274,N_5211);
nand U5548 (N_5548,N_5395,N_5360);
or U5549 (N_5549,N_5208,N_5339);
nor U5550 (N_5550,N_5381,N_5289);
nand U5551 (N_5551,N_5312,N_5261);
xnor U5552 (N_5552,N_5285,N_5320);
or U5553 (N_5553,N_5254,N_5295);
or U5554 (N_5554,N_5240,N_5288);
nor U5555 (N_5555,N_5366,N_5319);
or U5556 (N_5556,N_5232,N_5288);
xor U5557 (N_5557,N_5263,N_5374);
nor U5558 (N_5558,N_5220,N_5399);
and U5559 (N_5559,N_5399,N_5360);
nor U5560 (N_5560,N_5232,N_5386);
nor U5561 (N_5561,N_5210,N_5351);
nand U5562 (N_5562,N_5354,N_5201);
or U5563 (N_5563,N_5204,N_5201);
xor U5564 (N_5564,N_5218,N_5340);
xor U5565 (N_5565,N_5340,N_5215);
nor U5566 (N_5566,N_5289,N_5276);
or U5567 (N_5567,N_5396,N_5389);
or U5568 (N_5568,N_5342,N_5230);
nor U5569 (N_5569,N_5297,N_5245);
and U5570 (N_5570,N_5259,N_5278);
nor U5571 (N_5571,N_5305,N_5310);
nand U5572 (N_5572,N_5239,N_5201);
and U5573 (N_5573,N_5310,N_5317);
xor U5574 (N_5574,N_5284,N_5378);
and U5575 (N_5575,N_5239,N_5328);
and U5576 (N_5576,N_5389,N_5287);
or U5577 (N_5577,N_5394,N_5298);
and U5578 (N_5578,N_5380,N_5325);
nand U5579 (N_5579,N_5355,N_5203);
nor U5580 (N_5580,N_5388,N_5222);
and U5581 (N_5581,N_5376,N_5346);
nor U5582 (N_5582,N_5301,N_5345);
and U5583 (N_5583,N_5222,N_5319);
or U5584 (N_5584,N_5315,N_5384);
xnor U5585 (N_5585,N_5391,N_5383);
or U5586 (N_5586,N_5215,N_5208);
xnor U5587 (N_5587,N_5253,N_5222);
nand U5588 (N_5588,N_5257,N_5227);
nand U5589 (N_5589,N_5296,N_5358);
or U5590 (N_5590,N_5300,N_5244);
or U5591 (N_5591,N_5210,N_5296);
xor U5592 (N_5592,N_5281,N_5249);
or U5593 (N_5593,N_5271,N_5365);
or U5594 (N_5594,N_5392,N_5397);
nor U5595 (N_5595,N_5206,N_5339);
nor U5596 (N_5596,N_5259,N_5206);
nand U5597 (N_5597,N_5327,N_5206);
or U5598 (N_5598,N_5358,N_5347);
xnor U5599 (N_5599,N_5254,N_5235);
nand U5600 (N_5600,N_5585,N_5400);
and U5601 (N_5601,N_5412,N_5474);
and U5602 (N_5602,N_5464,N_5479);
and U5603 (N_5603,N_5458,N_5492);
nor U5604 (N_5604,N_5404,N_5524);
or U5605 (N_5605,N_5519,N_5537);
nor U5606 (N_5606,N_5454,N_5558);
xor U5607 (N_5607,N_5543,N_5551);
nand U5608 (N_5608,N_5583,N_5575);
or U5609 (N_5609,N_5573,N_5430);
nor U5610 (N_5610,N_5417,N_5507);
nand U5611 (N_5611,N_5520,N_5529);
xor U5612 (N_5612,N_5548,N_5594);
or U5613 (N_5613,N_5442,N_5418);
or U5614 (N_5614,N_5440,N_5406);
or U5615 (N_5615,N_5439,N_5505);
xnor U5616 (N_5616,N_5403,N_5441);
or U5617 (N_5617,N_5416,N_5574);
and U5618 (N_5618,N_5487,N_5553);
nand U5619 (N_5619,N_5556,N_5437);
xnor U5620 (N_5620,N_5523,N_5456);
nand U5621 (N_5621,N_5592,N_5436);
nand U5622 (N_5622,N_5434,N_5426);
xor U5623 (N_5623,N_5460,N_5545);
nor U5624 (N_5624,N_5517,N_5531);
nand U5625 (N_5625,N_5470,N_5569);
and U5626 (N_5626,N_5564,N_5457);
or U5627 (N_5627,N_5544,N_5424);
or U5628 (N_5628,N_5435,N_5473);
xor U5629 (N_5629,N_5444,N_5518);
and U5630 (N_5630,N_5550,N_5496);
xor U5631 (N_5631,N_5503,N_5485);
or U5632 (N_5632,N_5451,N_5552);
and U5633 (N_5633,N_5405,N_5576);
or U5634 (N_5634,N_5532,N_5565);
nand U5635 (N_5635,N_5528,N_5534);
nand U5636 (N_5636,N_5539,N_5504);
or U5637 (N_5637,N_5494,N_5411);
or U5638 (N_5638,N_5459,N_5579);
and U5639 (N_5639,N_5402,N_5509);
xor U5640 (N_5640,N_5567,N_5493);
and U5641 (N_5641,N_5431,N_5483);
or U5642 (N_5642,N_5535,N_5536);
xnor U5643 (N_5643,N_5508,N_5513);
xnor U5644 (N_5644,N_5433,N_5484);
xnor U5645 (N_5645,N_5486,N_5467);
nand U5646 (N_5646,N_5572,N_5480);
nor U5647 (N_5647,N_5407,N_5582);
and U5648 (N_5648,N_5596,N_5413);
nor U5649 (N_5649,N_5421,N_5559);
or U5650 (N_5650,N_5488,N_5581);
nor U5651 (N_5651,N_5547,N_5453);
and U5652 (N_5652,N_5477,N_5490);
nor U5653 (N_5653,N_5452,N_5530);
or U5654 (N_5654,N_5566,N_5538);
and U5655 (N_5655,N_5408,N_5465);
nand U5656 (N_5656,N_5481,N_5590);
nand U5657 (N_5657,N_5475,N_5587);
or U5658 (N_5658,N_5429,N_5591);
nor U5659 (N_5659,N_5571,N_5560);
and U5660 (N_5660,N_5506,N_5455);
nand U5661 (N_5661,N_5511,N_5462);
nor U5662 (N_5662,N_5562,N_5468);
or U5663 (N_5663,N_5414,N_5546);
and U5664 (N_5664,N_5522,N_5586);
nand U5665 (N_5665,N_5554,N_5515);
or U5666 (N_5666,N_5489,N_5449);
or U5667 (N_5667,N_5428,N_5447);
nand U5668 (N_5668,N_5526,N_5423);
and U5669 (N_5669,N_5472,N_5540);
nand U5670 (N_5670,N_5438,N_5570);
and U5671 (N_5671,N_5445,N_5478);
nand U5672 (N_5672,N_5598,N_5499);
and U5673 (N_5673,N_5555,N_5471);
xnor U5674 (N_5674,N_5425,N_5527);
or U5675 (N_5675,N_5415,N_5525);
or U5676 (N_5676,N_5512,N_5549);
nand U5677 (N_5677,N_5502,N_5580);
nor U5678 (N_5678,N_5577,N_5498);
and U5679 (N_5679,N_5561,N_5589);
and U5680 (N_5680,N_5469,N_5595);
and U5681 (N_5681,N_5495,N_5466);
and U5682 (N_5682,N_5491,N_5427);
or U5683 (N_5683,N_5584,N_5593);
or U5684 (N_5684,N_5500,N_5443);
nand U5685 (N_5685,N_5497,N_5410);
or U5686 (N_5686,N_5557,N_5599);
and U5687 (N_5687,N_5541,N_5542);
nand U5688 (N_5688,N_5432,N_5521);
nor U5689 (N_5689,N_5563,N_5461);
and U5690 (N_5690,N_5419,N_5501);
nand U5691 (N_5691,N_5482,N_5588);
nor U5692 (N_5692,N_5533,N_5514);
or U5693 (N_5693,N_5446,N_5516);
xor U5694 (N_5694,N_5450,N_5476);
and U5695 (N_5695,N_5578,N_5401);
or U5696 (N_5696,N_5597,N_5422);
nor U5697 (N_5697,N_5568,N_5448);
nand U5698 (N_5698,N_5463,N_5409);
or U5699 (N_5699,N_5510,N_5420);
or U5700 (N_5700,N_5441,N_5473);
or U5701 (N_5701,N_5536,N_5468);
nand U5702 (N_5702,N_5536,N_5547);
nand U5703 (N_5703,N_5513,N_5573);
nor U5704 (N_5704,N_5494,N_5519);
nor U5705 (N_5705,N_5465,N_5580);
xor U5706 (N_5706,N_5496,N_5546);
and U5707 (N_5707,N_5434,N_5495);
nor U5708 (N_5708,N_5560,N_5479);
xnor U5709 (N_5709,N_5554,N_5588);
nand U5710 (N_5710,N_5447,N_5425);
xnor U5711 (N_5711,N_5484,N_5548);
nand U5712 (N_5712,N_5408,N_5589);
and U5713 (N_5713,N_5410,N_5529);
nor U5714 (N_5714,N_5514,N_5564);
nand U5715 (N_5715,N_5470,N_5444);
and U5716 (N_5716,N_5521,N_5485);
or U5717 (N_5717,N_5598,N_5479);
xor U5718 (N_5718,N_5528,N_5432);
nand U5719 (N_5719,N_5563,N_5530);
or U5720 (N_5720,N_5561,N_5547);
nand U5721 (N_5721,N_5575,N_5537);
xor U5722 (N_5722,N_5404,N_5523);
or U5723 (N_5723,N_5585,N_5409);
xnor U5724 (N_5724,N_5422,N_5491);
and U5725 (N_5725,N_5427,N_5418);
and U5726 (N_5726,N_5429,N_5540);
xor U5727 (N_5727,N_5431,N_5475);
nand U5728 (N_5728,N_5451,N_5467);
or U5729 (N_5729,N_5524,N_5503);
nor U5730 (N_5730,N_5446,N_5557);
xnor U5731 (N_5731,N_5461,N_5591);
nand U5732 (N_5732,N_5439,N_5463);
and U5733 (N_5733,N_5449,N_5475);
and U5734 (N_5734,N_5517,N_5479);
and U5735 (N_5735,N_5561,N_5573);
xor U5736 (N_5736,N_5594,N_5543);
and U5737 (N_5737,N_5452,N_5568);
xor U5738 (N_5738,N_5464,N_5469);
and U5739 (N_5739,N_5431,N_5568);
nand U5740 (N_5740,N_5522,N_5527);
and U5741 (N_5741,N_5468,N_5439);
xor U5742 (N_5742,N_5400,N_5573);
or U5743 (N_5743,N_5488,N_5479);
nand U5744 (N_5744,N_5587,N_5552);
xnor U5745 (N_5745,N_5599,N_5429);
xor U5746 (N_5746,N_5403,N_5561);
nand U5747 (N_5747,N_5460,N_5483);
nor U5748 (N_5748,N_5489,N_5465);
nand U5749 (N_5749,N_5401,N_5545);
xor U5750 (N_5750,N_5592,N_5469);
xnor U5751 (N_5751,N_5434,N_5542);
nand U5752 (N_5752,N_5562,N_5490);
nand U5753 (N_5753,N_5523,N_5466);
or U5754 (N_5754,N_5528,N_5527);
or U5755 (N_5755,N_5444,N_5482);
nor U5756 (N_5756,N_5479,N_5515);
nand U5757 (N_5757,N_5551,N_5485);
or U5758 (N_5758,N_5570,N_5408);
or U5759 (N_5759,N_5452,N_5406);
nand U5760 (N_5760,N_5425,N_5512);
nand U5761 (N_5761,N_5474,N_5401);
or U5762 (N_5762,N_5416,N_5419);
xor U5763 (N_5763,N_5418,N_5561);
or U5764 (N_5764,N_5471,N_5503);
nor U5765 (N_5765,N_5478,N_5483);
xor U5766 (N_5766,N_5543,N_5407);
xnor U5767 (N_5767,N_5543,N_5433);
nor U5768 (N_5768,N_5591,N_5549);
nand U5769 (N_5769,N_5452,N_5544);
nand U5770 (N_5770,N_5438,N_5414);
or U5771 (N_5771,N_5432,N_5539);
nor U5772 (N_5772,N_5505,N_5454);
nand U5773 (N_5773,N_5475,N_5493);
nand U5774 (N_5774,N_5529,N_5444);
and U5775 (N_5775,N_5525,N_5537);
nand U5776 (N_5776,N_5563,N_5460);
or U5777 (N_5777,N_5579,N_5589);
and U5778 (N_5778,N_5485,N_5531);
xor U5779 (N_5779,N_5442,N_5498);
nor U5780 (N_5780,N_5589,N_5425);
nor U5781 (N_5781,N_5443,N_5520);
xnor U5782 (N_5782,N_5568,N_5547);
nor U5783 (N_5783,N_5428,N_5528);
or U5784 (N_5784,N_5430,N_5408);
nor U5785 (N_5785,N_5575,N_5493);
nor U5786 (N_5786,N_5552,N_5445);
xor U5787 (N_5787,N_5468,N_5453);
or U5788 (N_5788,N_5457,N_5532);
or U5789 (N_5789,N_5454,N_5494);
nor U5790 (N_5790,N_5413,N_5444);
nand U5791 (N_5791,N_5508,N_5558);
or U5792 (N_5792,N_5489,N_5452);
nand U5793 (N_5793,N_5462,N_5486);
or U5794 (N_5794,N_5403,N_5433);
and U5795 (N_5795,N_5403,N_5570);
nand U5796 (N_5796,N_5435,N_5463);
or U5797 (N_5797,N_5409,N_5482);
or U5798 (N_5798,N_5494,N_5444);
nand U5799 (N_5799,N_5501,N_5434);
xor U5800 (N_5800,N_5638,N_5775);
and U5801 (N_5801,N_5672,N_5746);
nand U5802 (N_5802,N_5695,N_5764);
nand U5803 (N_5803,N_5624,N_5777);
nor U5804 (N_5804,N_5651,N_5759);
nand U5805 (N_5805,N_5784,N_5761);
xnor U5806 (N_5806,N_5617,N_5608);
and U5807 (N_5807,N_5781,N_5694);
nand U5808 (N_5808,N_5686,N_5636);
xor U5809 (N_5809,N_5709,N_5690);
xor U5810 (N_5810,N_5696,N_5737);
nand U5811 (N_5811,N_5730,N_5606);
and U5812 (N_5812,N_5734,N_5741);
and U5813 (N_5813,N_5689,N_5665);
xor U5814 (N_5814,N_5646,N_5715);
and U5815 (N_5815,N_5799,N_5660);
or U5816 (N_5816,N_5693,N_5621);
xnor U5817 (N_5817,N_5722,N_5755);
and U5818 (N_5818,N_5684,N_5779);
nand U5819 (N_5819,N_5794,N_5749);
xnor U5820 (N_5820,N_5674,N_5787);
nor U5821 (N_5821,N_5616,N_5644);
and U5822 (N_5822,N_5654,N_5735);
xnor U5823 (N_5823,N_5685,N_5655);
and U5824 (N_5824,N_5704,N_5656);
nor U5825 (N_5825,N_5600,N_5700);
nand U5826 (N_5826,N_5783,N_5642);
nand U5827 (N_5827,N_5743,N_5745);
nor U5828 (N_5828,N_5632,N_5698);
nand U5829 (N_5829,N_5767,N_5723);
nand U5830 (N_5830,N_5776,N_5687);
or U5831 (N_5831,N_5659,N_5673);
nor U5832 (N_5832,N_5724,N_5748);
or U5833 (N_5833,N_5758,N_5782);
xnor U5834 (N_5834,N_5752,N_5631);
nand U5835 (N_5835,N_5765,N_5726);
and U5836 (N_5836,N_5653,N_5760);
xnor U5837 (N_5837,N_5742,N_5792);
nand U5838 (N_5838,N_5670,N_5729);
xor U5839 (N_5839,N_5603,N_5699);
and U5840 (N_5840,N_5721,N_5790);
nor U5841 (N_5841,N_5705,N_5680);
nand U5842 (N_5842,N_5733,N_5681);
and U5843 (N_5843,N_5763,N_5703);
and U5844 (N_5844,N_5645,N_5716);
and U5845 (N_5845,N_5697,N_5648);
xnor U5846 (N_5846,N_5641,N_5675);
nor U5847 (N_5847,N_5676,N_5797);
and U5848 (N_5848,N_5679,N_5702);
xor U5849 (N_5849,N_5612,N_5717);
and U5850 (N_5850,N_5618,N_5662);
xnor U5851 (N_5851,N_5605,N_5780);
nor U5852 (N_5852,N_5634,N_5643);
nand U5853 (N_5853,N_5762,N_5640);
and U5854 (N_5854,N_5772,N_5768);
or U5855 (N_5855,N_5701,N_5753);
nor U5856 (N_5856,N_5615,N_5630);
and U5857 (N_5857,N_5633,N_5778);
and U5858 (N_5858,N_5736,N_5789);
nor U5859 (N_5859,N_5607,N_5732);
and U5860 (N_5860,N_5744,N_5620);
nor U5861 (N_5861,N_5650,N_5718);
xor U5862 (N_5862,N_5738,N_5663);
and U5863 (N_5863,N_5739,N_5714);
and U5864 (N_5864,N_5667,N_5750);
nor U5865 (N_5865,N_5788,N_5731);
or U5866 (N_5866,N_5728,N_5658);
or U5867 (N_5867,N_5602,N_5691);
or U5868 (N_5868,N_5747,N_5706);
and U5869 (N_5869,N_5683,N_5629);
or U5870 (N_5870,N_5666,N_5601);
nand U5871 (N_5871,N_5637,N_5627);
xnor U5872 (N_5872,N_5708,N_5711);
nand U5873 (N_5873,N_5785,N_5719);
nand U5874 (N_5874,N_5725,N_5635);
nand U5875 (N_5875,N_5647,N_5771);
nor U5876 (N_5876,N_5611,N_5727);
xnor U5877 (N_5877,N_5626,N_5649);
and U5878 (N_5878,N_5639,N_5604);
xor U5879 (N_5879,N_5798,N_5710);
xor U5880 (N_5880,N_5609,N_5713);
nor U5881 (N_5881,N_5657,N_5628);
and U5882 (N_5882,N_5614,N_5664);
nor U5883 (N_5883,N_5692,N_5661);
xnor U5884 (N_5884,N_5712,N_5786);
and U5885 (N_5885,N_5774,N_5754);
and U5886 (N_5886,N_5791,N_5707);
and U5887 (N_5887,N_5668,N_5619);
and U5888 (N_5888,N_5677,N_5610);
xnor U5889 (N_5889,N_5751,N_5652);
and U5890 (N_5890,N_5769,N_5773);
nand U5891 (N_5891,N_5720,N_5757);
and U5892 (N_5892,N_5793,N_5766);
or U5893 (N_5893,N_5613,N_5740);
xnor U5894 (N_5894,N_5622,N_5756);
nand U5895 (N_5895,N_5625,N_5770);
nand U5896 (N_5896,N_5671,N_5678);
and U5897 (N_5897,N_5623,N_5669);
xor U5898 (N_5898,N_5688,N_5682);
and U5899 (N_5899,N_5796,N_5795);
nor U5900 (N_5900,N_5609,N_5757);
and U5901 (N_5901,N_5679,N_5674);
nor U5902 (N_5902,N_5621,N_5785);
or U5903 (N_5903,N_5746,N_5604);
nor U5904 (N_5904,N_5608,N_5690);
and U5905 (N_5905,N_5738,N_5668);
or U5906 (N_5906,N_5766,N_5790);
nand U5907 (N_5907,N_5726,N_5616);
nor U5908 (N_5908,N_5725,N_5638);
nand U5909 (N_5909,N_5639,N_5680);
nor U5910 (N_5910,N_5755,N_5621);
nand U5911 (N_5911,N_5750,N_5670);
and U5912 (N_5912,N_5678,N_5664);
xor U5913 (N_5913,N_5625,N_5710);
nand U5914 (N_5914,N_5732,N_5675);
nand U5915 (N_5915,N_5656,N_5680);
xor U5916 (N_5916,N_5623,N_5666);
nand U5917 (N_5917,N_5661,N_5662);
nor U5918 (N_5918,N_5732,N_5636);
or U5919 (N_5919,N_5740,N_5634);
nand U5920 (N_5920,N_5786,N_5682);
xor U5921 (N_5921,N_5688,N_5749);
xor U5922 (N_5922,N_5672,N_5700);
or U5923 (N_5923,N_5788,N_5638);
xnor U5924 (N_5924,N_5752,N_5722);
and U5925 (N_5925,N_5645,N_5734);
or U5926 (N_5926,N_5667,N_5674);
nor U5927 (N_5927,N_5747,N_5601);
nand U5928 (N_5928,N_5683,N_5752);
or U5929 (N_5929,N_5712,N_5743);
nand U5930 (N_5930,N_5679,N_5797);
and U5931 (N_5931,N_5747,N_5795);
or U5932 (N_5932,N_5675,N_5661);
nand U5933 (N_5933,N_5637,N_5796);
nand U5934 (N_5934,N_5631,N_5776);
xnor U5935 (N_5935,N_5636,N_5702);
xnor U5936 (N_5936,N_5707,N_5644);
nor U5937 (N_5937,N_5712,N_5640);
and U5938 (N_5938,N_5748,N_5727);
and U5939 (N_5939,N_5688,N_5715);
nand U5940 (N_5940,N_5776,N_5637);
xor U5941 (N_5941,N_5660,N_5795);
nand U5942 (N_5942,N_5737,N_5609);
and U5943 (N_5943,N_5662,N_5778);
nand U5944 (N_5944,N_5668,N_5690);
or U5945 (N_5945,N_5672,N_5701);
or U5946 (N_5946,N_5722,N_5778);
and U5947 (N_5947,N_5778,N_5779);
or U5948 (N_5948,N_5635,N_5766);
or U5949 (N_5949,N_5772,N_5675);
or U5950 (N_5950,N_5780,N_5757);
or U5951 (N_5951,N_5683,N_5627);
and U5952 (N_5952,N_5718,N_5608);
nand U5953 (N_5953,N_5666,N_5738);
nor U5954 (N_5954,N_5660,N_5748);
nand U5955 (N_5955,N_5690,N_5721);
nor U5956 (N_5956,N_5791,N_5705);
nand U5957 (N_5957,N_5778,N_5644);
or U5958 (N_5958,N_5734,N_5743);
xnor U5959 (N_5959,N_5623,N_5740);
nor U5960 (N_5960,N_5775,N_5635);
nand U5961 (N_5961,N_5623,N_5686);
nand U5962 (N_5962,N_5637,N_5739);
or U5963 (N_5963,N_5721,N_5662);
nor U5964 (N_5964,N_5719,N_5684);
or U5965 (N_5965,N_5621,N_5783);
nand U5966 (N_5966,N_5735,N_5646);
xnor U5967 (N_5967,N_5610,N_5653);
xor U5968 (N_5968,N_5765,N_5648);
and U5969 (N_5969,N_5699,N_5716);
xor U5970 (N_5970,N_5760,N_5788);
xnor U5971 (N_5971,N_5740,N_5797);
xnor U5972 (N_5972,N_5723,N_5781);
nand U5973 (N_5973,N_5740,N_5646);
or U5974 (N_5974,N_5661,N_5712);
xnor U5975 (N_5975,N_5711,N_5691);
nand U5976 (N_5976,N_5765,N_5712);
and U5977 (N_5977,N_5627,N_5619);
nand U5978 (N_5978,N_5639,N_5778);
xnor U5979 (N_5979,N_5693,N_5764);
nand U5980 (N_5980,N_5690,N_5629);
nor U5981 (N_5981,N_5681,N_5629);
or U5982 (N_5982,N_5611,N_5795);
or U5983 (N_5983,N_5753,N_5745);
or U5984 (N_5984,N_5641,N_5795);
nor U5985 (N_5985,N_5745,N_5621);
and U5986 (N_5986,N_5780,N_5787);
nand U5987 (N_5987,N_5736,N_5711);
and U5988 (N_5988,N_5687,N_5658);
and U5989 (N_5989,N_5745,N_5720);
or U5990 (N_5990,N_5730,N_5752);
xnor U5991 (N_5991,N_5698,N_5604);
nand U5992 (N_5992,N_5780,N_5637);
or U5993 (N_5993,N_5682,N_5670);
xnor U5994 (N_5994,N_5686,N_5743);
and U5995 (N_5995,N_5625,N_5649);
and U5996 (N_5996,N_5625,N_5707);
or U5997 (N_5997,N_5792,N_5631);
nor U5998 (N_5998,N_5745,N_5611);
nor U5999 (N_5999,N_5779,N_5769);
and U6000 (N_6000,N_5911,N_5807);
and U6001 (N_6001,N_5966,N_5940);
and U6002 (N_6002,N_5891,N_5865);
xor U6003 (N_6003,N_5840,N_5882);
nand U6004 (N_6004,N_5871,N_5879);
nand U6005 (N_6005,N_5820,N_5895);
nand U6006 (N_6006,N_5979,N_5814);
nor U6007 (N_6007,N_5866,N_5901);
xor U6008 (N_6008,N_5876,N_5809);
xnor U6009 (N_6009,N_5837,N_5877);
xnor U6010 (N_6010,N_5830,N_5961);
and U6011 (N_6011,N_5846,N_5917);
xnor U6012 (N_6012,N_5999,N_5887);
or U6013 (N_6013,N_5878,N_5982);
nor U6014 (N_6014,N_5897,N_5974);
nor U6015 (N_6015,N_5800,N_5947);
or U6016 (N_6016,N_5910,N_5896);
or U6017 (N_6017,N_5909,N_5852);
nor U6018 (N_6018,N_5936,N_5839);
nor U6019 (N_6019,N_5973,N_5953);
xnor U6020 (N_6020,N_5822,N_5843);
or U6021 (N_6021,N_5854,N_5811);
nor U6022 (N_6022,N_5905,N_5823);
or U6023 (N_6023,N_5874,N_5951);
nor U6024 (N_6024,N_5875,N_5934);
xor U6025 (N_6025,N_5838,N_5926);
nor U6026 (N_6026,N_5991,N_5819);
nor U6027 (N_6027,N_5826,N_5806);
or U6028 (N_6028,N_5930,N_5888);
nor U6029 (N_6029,N_5912,N_5922);
nand U6030 (N_6030,N_5935,N_5921);
and U6031 (N_6031,N_5928,N_5899);
or U6032 (N_6032,N_5802,N_5927);
or U6033 (N_6033,N_5968,N_5817);
xnor U6034 (N_6034,N_5872,N_5941);
xnor U6035 (N_6035,N_5808,N_5849);
nor U6036 (N_6036,N_5946,N_5913);
and U6037 (N_6037,N_5975,N_5932);
and U6038 (N_6038,N_5836,N_5864);
or U6039 (N_6039,N_5976,N_5933);
xnor U6040 (N_6040,N_5937,N_5825);
xor U6041 (N_6041,N_5850,N_5869);
and U6042 (N_6042,N_5831,N_5805);
xor U6043 (N_6043,N_5965,N_5944);
nor U6044 (N_6044,N_5907,N_5916);
nor U6045 (N_6045,N_5998,N_5980);
and U6046 (N_6046,N_5954,N_5952);
nor U6047 (N_6047,N_5983,N_5956);
and U6048 (N_6048,N_5860,N_5903);
and U6049 (N_6049,N_5915,N_5883);
or U6050 (N_6050,N_5851,N_5813);
xor U6051 (N_6051,N_5945,N_5943);
and U6052 (N_6052,N_5859,N_5950);
xor U6053 (N_6053,N_5925,N_5827);
nand U6054 (N_6054,N_5845,N_5893);
nand U6055 (N_6055,N_5918,N_5873);
nand U6056 (N_6056,N_5962,N_5994);
nand U6057 (N_6057,N_5995,N_5889);
or U6058 (N_6058,N_5942,N_5890);
nand U6059 (N_6059,N_5986,N_5862);
and U6060 (N_6060,N_5978,N_5870);
xor U6061 (N_6061,N_5969,N_5861);
and U6062 (N_6062,N_5902,N_5816);
and U6063 (N_6063,N_5858,N_5993);
nor U6064 (N_6064,N_5988,N_5923);
or U6065 (N_6065,N_5929,N_5931);
nand U6066 (N_6066,N_5863,N_5970);
xnor U6067 (N_6067,N_5920,N_5804);
nor U6068 (N_6068,N_5892,N_5924);
or U6069 (N_6069,N_5841,N_5960);
xnor U6070 (N_6070,N_5967,N_5985);
and U6071 (N_6071,N_5972,N_5853);
nor U6072 (N_6072,N_5880,N_5963);
xnor U6073 (N_6073,N_5914,N_5955);
xnor U6074 (N_6074,N_5803,N_5948);
nand U6075 (N_6075,N_5957,N_5958);
xor U6076 (N_6076,N_5977,N_5886);
and U6077 (N_6077,N_5992,N_5996);
xor U6078 (N_6078,N_5938,N_5919);
nor U6079 (N_6079,N_5959,N_5828);
nor U6080 (N_6080,N_5844,N_5939);
xnor U6081 (N_6081,N_5833,N_5867);
and U6082 (N_6082,N_5815,N_5981);
nand U6083 (N_6083,N_5964,N_5990);
and U6084 (N_6084,N_5997,N_5855);
xor U6085 (N_6085,N_5987,N_5885);
and U6086 (N_6086,N_5801,N_5842);
xnor U6087 (N_6087,N_5824,N_5904);
nor U6088 (N_6088,N_5848,N_5884);
and U6089 (N_6089,N_5810,N_5900);
nand U6090 (N_6090,N_5908,N_5984);
or U6091 (N_6091,N_5989,N_5821);
nand U6092 (N_6092,N_5818,N_5949);
xnor U6093 (N_6093,N_5971,N_5868);
xnor U6094 (N_6094,N_5834,N_5835);
or U6095 (N_6095,N_5812,N_5906);
or U6096 (N_6096,N_5829,N_5894);
nor U6097 (N_6097,N_5832,N_5857);
nand U6098 (N_6098,N_5898,N_5881);
nand U6099 (N_6099,N_5856,N_5847);
nor U6100 (N_6100,N_5874,N_5856);
nand U6101 (N_6101,N_5803,N_5958);
nor U6102 (N_6102,N_5861,N_5830);
or U6103 (N_6103,N_5863,N_5963);
or U6104 (N_6104,N_5997,N_5951);
nand U6105 (N_6105,N_5878,N_5815);
and U6106 (N_6106,N_5876,N_5977);
or U6107 (N_6107,N_5826,N_5836);
nand U6108 (N_6108,N_5982,N_5999);
xnor U6109 (N_6109,N_5807,N_5842);
and U6110 (N_6110,N_5896,N_5921);
nand U6111 (N_6111,N_5998,N_5898);
xnor U6112 (N_6112,N_5829,N_5846);
and U6113 (N_6113,N_5917,N_5819);
xor U6114 (N_6114,N_5998,N_5820);
and U6115 (N_6115,N_5822,N_5886);
nand U6116 (N_6116,N_5907,N_5885);
nor U6117 (N_6117,N_5877,N_5803);
or U6118 (N_6118,N_5924,N_5921);
nor U6119 (N_6119,N_5900,N_5982);
nor U6120 (N_6120,N_5956,N_5898);
or U6121 (N_6121,N_5875,N_5863);
xnor U6122 (N_6122,N_5805,N_5895);
nor U6123 (N_6123,N_5805,N_5834);
or U6124 (N_6124,N_5804,N_5932);
nand U6125 (N_6125,N_5860,N_5989);
or U6126 (N_6126,N_5877,N_5893);
nor U6127 (N_6127,N_5962,N_5893);
nand U6128 (N_6128,N_5850,N_5964);
or U6129 (N_6129,N_5955,N_5901);
xnor U6130 (N_6130,N_5956,N_5987);
and U6131 (N_6131,N_5818,N_5960);
xnor U6132 (N_6132,N_5840,N_5816);
and U6133 (N_6133,N_5870,N_5986);
xnor U6134 (N_6134,N_5952,N_5859);
nand U6135 (N_6135,N_5893,N_5816);
and U6136 (N_6136,N_5919,N_5811);
xnor U6137 (N_6137,N_5910,N_5834);
nand U6138 (N_6138,N_5878,N_5885);
xnor U6139 (N_6139,N_5998,N_5812);
or U6140 (N_6140,N_5971,N_5988);
or U6141 (N_6141,N_5831,N_5884);
nor U6142 (N_6142,N_5830,N_5857);
and U6143 (N_6143,N_5940,N_5978);
and U6144 (N_6144,N_5921,N_5836);
and U6145 (N_6145,N_5808,N_5958);
and U6146 (N_6146,N_5808,N_5873);
or U6147 (N_6147,N_5991,N_5919);
nand U6148 (N_6148,N_5832,N_5997);
xnor U6149 (N_6149,N_5823,N_5904);
and U6150 (N_6150,N_5985,N_5880);
and U6151 (N_6151,N_5955,N_5816);
or U6152 (N_6152,N_5963,N_5885);
nand U6153 (N_6153,N_5887,N_5954);
and U6154 (N_6154,N_5945,N_5938);
nand U6155 (N_6155,N_5894,N_5915);
nand U6156 (N_6156,N_5906,N_5860);
and U6157 (N_6157,N_5945,N_5999);
nand U6158 (N_6158,N_5813,N_5959);
nor U6159 (N_6159,N_5858,N_5886);
and U6160 (N_6160,N_5823,N_5874);
xnor U6161 (N_6161,N_5845,N_5933);
nor U6162 (N_6162,N_5904,N_5874);
or U6163 (N_6163,N_5972,N_5907);
and U6164 (N_6164,N_5952,N_5918);
nand U6165 (N_6165,N_5853,N_5958);
nor U6166 (N_6166,N_5889,N_5813);
and U6167 (N_6167,N_5989,N_5822);
and U6168 (N_6168,N_5813,N_5929);
or U6169 (N_6169,N_5932,N_5967);
nor U6170 (N_6170,N_5960,N_5898);
nor U6171 (N_6171,N_5984,N_5894);
and U6172 (N_6172,N_5956,N_5940);
and U6173 (N_6173,N_5986,N_5918);
and U6174 (N_6174,N_5919,N_5821);
nand U6175 (N_6175,N_5962,N_5858);
nor U6176 (N_6176,N_5916,N_5843);
xor U6177 (N_6177,N_5909,N_5806);
or U6178 (N_6178,N_5871,N_5809);
nand U6179 (N_6179,N_5985,N_5860);
xnor U6180 (N_6180,N_5984,N_5861);
and U6181 (N_6181,N_5820,N_5992);
xor U6182 (N_6182,N_5869,N_5923);
nand U6183 (N_6183,N_5985,N_5974);
nor U6184 (N_6184,N_5807,N_5946);
nor U6185 (N_6185,N_5925,N_5888);
or U6186 (N_6186,N_5986,N_5984);
and U6187 (N_6187,N_5913,N_5879);
and U6188 (N_6188,N_5803,N_5941);
and U6189 (N_6189,N_5932,N_5826);
nand U6190 (N_6190,N_5840,N_5827);
or U6191 (N_6191,N_5977,N_5802);
or U6192 (N_6192,N_5898,N_5824);
and U6193 (N_6193,N_5924,N_5917);
nor U6194 (N_6194,N_5894,N_5888);
or U6195 (N_6195,N_5906,N_5842);
and U6196 (N_6196,N_5910,N_5948);
or U6197 (N_6197,N_5971,N_5921);
and U6198 (N_6198,N_5971,N_5982);
xnor U6199 (N_6199,N_5985,N_5895);
xor U6200 (N_6200,N_6111,N_6156);
nor U6201 (N_6201,N_6060,N_6177);
and U6202 (N_6202,N_6121,N_6018);
nand U6203 (N_6203,N_6071,N_6074);
xor U6204 (N_6204,N_6098,N_6168);
and U6205 (N_6205,N_6178,N_6195);
nand U6206 (N_6206,N_6193,N_6009);
and U6207 (N_6207,N_6122,N_6145);
xnor U6208 (N_6208,N_6170,N_6065);
nor U6209 (N_6209,N_6093,N_6078);
and U6210 (N_6210,N_6107,N_6116);
or U6211 (N_6211,N_6128,N_6134);
xor U6212 (N_6212,N_6056,N_6023);
or U6213 (N_6213,N_6010,N_6186);
or U6214 (N_6214,N_6125,N_6095);
and U6215 (N_6215,N_6058,N_6040);
xnor U6216 (N_6216,N_6028,N_6029);
or U6217 (N_6217,N_6011,N_6072);
nand U6218 (N_6218,N_6114,N_6135);
nand U6219 (N_6219,N_6117,N_6006);
nand U6220 (N_6220,N_6039,N_6064);
and U6221 (N_6221,N_6090,N_6196);
nand U6222 (N_6222,N_6187,N_6008);
nand U6223 (N_6223,N_6052,N_6126);
or U6224 (N_6224,N_6034,N_6139);
xor U6225 (N_6225,N_6094,N_6015);
nor U6226 (N_6226,N_6081,N_6017);
and U6227 (N_6227,N_6147,N_6155);
xor U6228 (N_6228,N_6012,N_6199);
nand U6229 (N_6229,N_6099,N_6119);
or U6230 (N_6230,N_6025,N_6057);
nor U6231 (N_6231,N_6113,N_6016);
nand U6232 (N_6232,N_6005,N_6007);
or U6233 (N_6233,N_6059,N_6164);
and U6234 (N_6234,N_6150,N_6054);
or U6235 (N_6235,N_6141,N_6104);
nand U6236 (N_6236,N_6082,N_6001);
and U6237 (N_6237,N_6152,N_6146);
xor U6238 (N_6238,N_6143,N_6045);
xor U6239 (N_6239,N_6102,N_6192);
xnor U6240 (N_6240,N_6038,N_6036);
nand U6241 (N_6241,N_6030,N_6138);
nor U6242 (N_6242,N_6154,N_6130);
nor U6243 (N_6243,N_6167,N_6096);
nand U6244 (N_6244,N_6142,N_6066);
and U6245 (N_6245,N_6194,N_6123);
xnor U6246 (N_6246,N_6000,N_6031);
xor U6247 (N_6247,N_6159,N_6077);
nor U6248 (N_6248,N_6151,N_6061);
and U6249 (N_6249,N_6105,N_6115);
nand U6250 (N_6250,N_6086,N_6014);
and U6251 (N_6251,N_6033,N_6190);
nand U6252 (N_6252,N_6019,N_6024);
nor U6253 (N_6253,N_6003,N_6026);
and U6254 (N_6254,N_6174,N_6048);
and U6255 (N_6255,N_6118,N_6136);
xnor U6256 (N_6256,N_6120,N_6160);
and U6257 (N_6257,N_6181,N_6087);
or U6258 (N_6258,N_6137,N_6032);
nor U6259 (N_6259,N_6124,N_6129);
xnor U6260 (N_6260,N_6049,N_6173);
or U6261 (N_6261,N_6042,N_6103);
or U6262 (N_6262,N_6037,N_6108);
nor U6263 (N_6263,N_6166,N_6084);
and U6264 (N_6264,N_6161,N_6191);
xnor U6265 (N_6265,N_6070,N_6185);
nand U6266 (N_6266,N_6182,N_6163);
or U6267 (N_6267,N_6109,N_6097);
and U6268 (N_6268,N_6169,N_6165);
and U6269 (N_6269,N_6046,N_6189);
nand U6270 (N_6270,N_6002,N_6184);
and U6271 (N_6271,N_6100,N_6110);
nand U6272 (N_6272,N_6183,N_6132);
or U6273 (N_6273,N_6148,N_6080);
or U6274 (N_6274,N_6076,N_6176);
or U6275 (N_6275,N_6092,N_6179);
xnor U6276 (N_6276,N_6089,N_6069);
and U6277 (N_6277,N_6013,N_6022);
and U6278 (N_6278,N_6149,N_6133);
or U6279 (N_6279,N_6053,N_6062);
and U6280 (N_6280,N_6068,N_6088);
and U6281 (N_6281,N_6041,N_6075);
xor U6282 (N_6282,N_6063,N_6020);
nand U6283 (N_6283,N_6144,N_6044);
xnor U6284 (N_6284,N_6079,N_6047);
xor U6285 (N_6285,N_6027,N_6112);
xnor U6286 (N_6286,N_6198,N_6085);
nand U6287 (N_6287,N_6162,N_6067);
nand U6288 (N_6288,N_6171,N_6083);
or U6289 (N_6289,N_6157,N_6101);
nor U6290 (N_6290,N_6140,N_6197);
or U6291 (N_6291,N_6131,N_6175);
nand U6292 (N_6292,N_6021,N_6180);
xnor U6293 (N_6293,N_6073,N_6004);
nor U6294 (N_6294,N_6172,N_6158);
nor U6295 (N_6295,N_6091,N_6050);
xnor U6296 (N_6296,N_6188,N_6055);
nor U6297 (N_6297,N_6051,N_6106);
or U6298 (N_6298,N_6153,N_6035);
or U6299 (N_6299,N_6127,N_6043);
nand U6300 (N_6300,N_6181,N_6176);
xnor U6301 (N_6301,N_6061,N_6199);
xnor U6302 (N_6302,N_6072,N_6121);
nand U6303 (N_6303,N_6038,N_6027);
nand U6304 (N_6304,N_6028,N_6065);
nor U6305 (N_6305,N_6097,N_6022);
xor U6306 (N_6306,N_6058,N_6009);
xor U6307 (N_6307,N_6135,N_6063);
or U6308 (N_6308,N_6071,N_6141);
nor U6309 (N_6309,N_6018,N_6050);
or U6310 (N_6310,N_6131,N_6071);
and U6311 (N_6311,N_6197,N_6163);
nand U6312 (N_6312,N_6012,N_6165);
and U6313 (N_6313,N_6185,N_6129);
xor U6314 (N_6314,N_6048,N_6109);
nor U6315 (N_6315,N_6044,N_6003);
and U6316 (N_6316,N_6181,N_6067);
nand U6317 (N_6317,N_6000,N_6092);
or U6318 (N_6318,N_6157,N_6121);
xnor U6319 (N_6319,N_6034,N_6083);
nor U6320 (N_6320,N_6076,N_6185);
and U6321 (N_6321,N_6059,N_6162);
and U6322 (N_6322,N_6036,N_6129);
xor U6323 (N_6323,N_6042,N_6080);
or U6324 (N_6324,N_6066,N_6110);
nand U6325 (N_6325,N_6120,N_6042);
and U6326 (N_6326,N_6041,N_6033);
nor U6327 (N_6327,N_6076,N_6050);
and U6328 (N_6328,N_6184,N_6020);
and U6329 (N_6329,N_6194,N_6103);
and U6330 (N_6330,N_6049,N_6044);
nor U6331 (N_6331,N_6053,N_6103);
nor U6332 (N_6332,N_6150,N_6166);
nor U6333 (N_6333,N_6163,N_6053);
nand U6334 (N_6334,N_6172,N_6021);
or U6335 (N_6335,N_6167,N_6114);
nor U6336 (N_6336,N_6129,N_6163);
and U6337 (N_6337,N_6036,N_6197);
nor U6338 (N_6338,N_6080,N_6020);
or U6339 (N_6339,N_6070,N_6085);
xnor U6340 (N_6340,N_6143,N_6088);
xnor U6341 (N_6341,N_6074,N_6091);
xor U6342 (N_6342,N_6140,N_6037);
nor U6343 (N_6343,N_6125,N_6196);
nand U6344 (N_6344,N_6066,N_6059);
nand U6345 (N_6345,N_6033,N_6046);
nor U6346 (N_6346,N_6032,N_6178);
xor U6347 (N_6347,N_6076,N_6175);
and U6348 (N_6348,N_6113,N_6097);
nand U6349 (N_6349,N_6020,N_6000);
nor U6350 (N_6350,N_6111,N_6164);
nor U6351 (N_6351,N_6029,N_6054);
xor U6352 (N_6352,N_6128,N_6022);
and U6353 (N_6353,N_6047,N_6055);
xor U6354 (N_6354,N_6138,N_6107);
or U6355 (N_6355,N_6119,N_6137);
nor U6356 (N_6356,N_6122,N_6011);
nor U6357 (N_6357,N_6186,N_6023);
nand U6358 (N_6358,N_6083,N_6164);
xor U6359 (N_6359,N_6041,N_6190);
nor U6360 (N_6360,N_6059,N_6029);
xnor U6361 (N_6361,N_6065,N_6131);
nor U6362 (N_6362,N_6128,N_6162);
xor U6363 (N_6363,N_6107,N_6114);
nor U6364 (N_6364,N_6088,N_6063);
nor U6365 (N_6365,N_6097,N_6139);
nand U6366 (N_6366,N_6177,N_6180);
xor U6367 (N_6367,N_6117,N_6182);
nor U6368 (N_6368,N_6080,N_6171);
or U6369 (N_6369,N_6079,N_6045);
or U6370 (N_6370,N_6191,N_6045);
nor U6371 (N_6371,N_6190,N_6080);
and U6372 (N_6372,N_6137,N_6197);
nand U6373 (N_6373,N_6184,N_6111);
nor U6374 (N_6374,N_6073,N_6095);
and U6375 (N_6375,N_6020,N_6135);
and U6376 (N_6376,N_6057,N_6175);
or U6377 (N_6377,N_6142,N_6059);
and U6378 (N_6378,N_6095,N_6198);
or U6379 (N_6379,N_6104,N_6013);
and U6380 (N_6380,N_6011,N_6146);
nor U6381 (N_6381,N_6118,N_6000);
or U6382 (N_6382,N_6036,N_6064);
xor U6383 (N_6383,N_6185,N_6079);
nand U6384 (N_6384,N_6173,N_6016);
nor U6385 (N_6385,N_6010,N_6106);
and U6386 (N_6386,N_6118,N_6048);
nand U6387 (N_6387,N_6114,N_6006);
nor U6388 (N_6388,N_6095,N_6057);
xnor U6389 (N_6389,N_6141,N_6088);
nor U6390 (N_6390,N_6179,N_6029);
xor U6391 (N_6391,N_6089,N_6062);
and U6392 (N_6392,N_6134,N_6093);
nor U6393 (N_6393,N_6067,N_6080);
nor U6394 (N_6394,N_6170,N_6074);
nand U6395 (N_6395,N_6162,N_6058);
nor U6396 (N_6396,N_6196,N_6154);
nand U6397 (N_6397,N_6171,N_6059);
xor U6398 (N_6398,N_6148,N_6094);
nand U6399 (N_6399,N_6058,N_6098);
or U6400 (N_6400,N_6287,N_6291);
and U6401 (N_6401,N_6350,N_6337);
or U6402 (N_6402,N_6207,N_6324);
or U6403 (N_6403,N_6262,N_6354);
and U6404 (N_6404,N_6302,N_6227);
or U6405 (N_6405,N_6244,N_6214);
nand U6406 (N_6406,N_6383,N_6379);
nand U6407 (N_6407,N_6323,N_6378);
or U6408 (N_6408,N_6239,N_6327);
nor U6409 (N_6409,N_6377,N_6376);
nand U6410 (N_6410,N_6202,N_6226);
and U6411 (N_6411,N_6333,N_6209);
or U6412 (N_6412,N_6204,N_6271);
or U6413 (N_6413,N_6251,N_6300);
xor U6414 (N_6414,N_6265,N_6257);
nand U6415 (N_6415,N_6320,N_6396);
and U6416 (N_6416,N_6370,N_6297);
or U6417 (N_6417,N_6298,N_6341);
or U6418 (N_6418,N_6367,N_6335);
nor U6419 (N_6419,N_6311,N_6253);
or U6420 (N_6420,N_6384,N_6213);
nor U6421 (N_6421,N_6283,N_6373);
xnor U6422 (N_6422,N_6375,N_6263);
and U6423 (N_6423,N_6254,N_6313);
xnor U6424 (N_6424,N_6279,N_6280);
xor U6425 (N_6425,N_6229,N_6348);
and U6426 (N_6426,N_6306,N_6390);
nor U6427 (N_6427,N_6345,N_6234);
nand U6428 (N_6428,N_6289,N_6366);
or U6429 (N_6429,N_6203,N_6266);
nand U6430 (N_6430,N_6387,N_6381);
nor U6431 (N_6431,N_6332,N_6281);
xor U6432 (N_6432,N_6355,N_6394);
xor U6433 (N_6433,N_6309,N_6270);
nand U6434 (N_6434,N_6351,N_6317);
xnor U6435 (N_6435,N_6236,N_6395);
and U6436 (N_6436,N_6388,N_6307);
or U6437 (N_6437,N_6356,N_6328);
or U6438 (N_6438,N_6358,N_6397);
and U6439 (N_6439,N_6346,N_6264);
nor U6440 (N_6440,N_6347,N_6278);
nand U6441 (N_6441,N_6261,N_6331);
xor U6442 (N_6442,N_6343,N_6369);
xnor U6443 (N_6443,N_6259,N_6292);
xnor U6444 (N_6444,N_6267,N_6235);
or U6445 (N_6445,N_6205,N_6241);
nand U6446 (N_6446,N_6296,N_6200);
nand U6447 (N_6447,N_6305,N_6308);
xnor U6448 (N_6448,N_6326,N_6315);
nand U6449 (N_6449,N_6372,N_6238);
or U6450 (N_6450,N_6360,N_6359);
or U6451 (N_6451,N_6250,N_6294);
and U6452 (N_6452,N_6225,N_6230);
and U6453 (N_6453,N_6334,N_6392);
xor U6454 (N_6454,N_6243,N_6299);
nor U6455 (N_6455,N_6339,N_6398);
and U6456 (N_6456,N_6374,N_6389);
or U6457 (N_6457,N_6223,N_6304);
and U6458 (N_6458,N_6393,N_6368);
nand U6459 (N_6459,N_6314,N_6336);
xor U6460 (N_6460,N_6240,N_6217);
and U6461 (N_6461,N_6242,N_6237);
and U6462 (N_6462,N_6275,N_6208);
or U6463 (N_6463,N_6246,N_6211);
and U6464 (N_6464,N_6316,N_6386);
and U6465 (N_6465,N_6301,N_6293);
xnor U6466 (N_6466,N_6340,N_6277);
or U6467 (N_6467,N_6321,N_6318);
and U6468 (N_6468,N_6295,N_6269);
xnor U6469 (N_6469,N_6221,N_6288);
nor U6470 (N_6470,N_6276,N_6219);
nor U6471 (N_6471,N_6247,N_6371);
or U6472 (N_6472,N_6312,N_6206);
nor U6473 (N_6473,N_6285,N_6218);
nor U6474 (N_6474,N_6216,N_6361);
nand U6475 (N_6475,N_6310,N_6201);
nand U6476 (N_6476,N_6260,N_6258);
nand U6477 (N_6477,N_6357,N_6232);
xnor U6478 (N_6478,N_6215,N_6228);
nor U6479 (N_6479,N_6284,N_6268);
nor U6480 (N_6480,N_6224,N_6248);
or U6481 (N_6481,N_6290,N_6325);
nand U6482 (N_6482,N_6249,N_6303);
or U6483 (N_6483,N_6330,N_6319);
or U6484 (N_6484,N_6282,N_6364);
nand U6485 (N_6485,N_6353,N_6385);
and U6486 (N_6486,N_6272,N_6255);
and U6487 (N_6487,N_6210,N_6212);
and U6488 (N_6488,N_6222,N_6322);
xor U6489 (N_6489,N_6399,N_6273);
nand U6490 (N_6490,N_6274,N_6252);
and U6491 (N_6491,N_6362,N_6365);
nor U6492 (N_6492,N_6352,N_6329);
and U6493 (N_6493,N_6344,N_6245);
nor U6494 (N_6494,N_6286,N_6380);
nand U6495 (N_6495,N_6256,N_6231);
nand U6496 (N_6496,N_6349,N_6382);
xnor U6497 (N_6497,N_6338,N_6363);
or U6498 (N_6498,N_6391,N_6220);
xnor U6499 (N_6499,N_6342,N_6233);
or U6500 (N_6500,N_6323,N_6244);
or U6501 (N_6501,N_6369,N_6213);
and U6502 (N_6502,N_6217,N_6321);
nand U6503 (N_6503,N_6343,N_6279);
nor U6504 (N_6504,N_6269,N_6380);
xnor U6505 (N_6505,N_6344,N_6298);
xnor U6506 (N_6506,N_6349,N_6238);
xnor U6507 (N_6507,N_6343,N_6386);
and U6508 (N_6508,N_6301,N_6297);
nand U6509 (N_6509,N_6252,N_6316);
and U6510 (N_6510,N_6370,N_6342);
nand U6511 (N_6511,N_6233,N_6315);
xor U6512 (N_6512,N_6222,N_6287);
and U6513 (N_6513,N_6243,N_6251);
nor U6514 (N_6514,N_6317,N_6209);
or U6515 (N_6515,N_6318,N_6289);
or U6516 (N_6516,N_6268,N_6341);
or U6517 (N_6517,N_6271,N_6372);
nor U6518 (N_6518,N_6289,N_6352);
nor U6519 (N_6519,N_6266,N_6272);
nand U6520 (N_6520,N_6334,N_6214);
or U6521 (N_6521,N_6211,N_6383);
and U6522 (N_6522,N_6345,N_6302);
or U6523 (N_6523,N_6338,N_6381);
or U6524 (N_6524,N_6340,N_6286);
nand U6525 (N_6525,N_6396,N_6374);
xor U6526 (N_6526,N_6340,N_6292);
xnor U6527 (N_6527,N_6388,N_6315);
or U6528 (N_6528,N_6216,N_6380);
xor U6529 (N_6529,N_6358,N_6361);
or U6530 (N_6530,N_6213,N_6396);
or U6531 (N_6531,N_6254,N_6353);
nor U6532 (N_6532,N_6356,N_6348);
nand U6533 (N_6533,N_6268,N_6336);
or U6534 (N_6534,N_6344,N_6221);
nor U6535 (N_6535,N_6340,N_6351);
nand U6536 (N_6536,N_6276,N_6354);
or U6537 (N_6537,N_6333,N_6391);
and U6538 (N_6538,N_6259,N_6208);
and U6539 (N_6539,N_6310,N_6209);
xnor U6540 (N_6540,N_6390,N_6319);
nor U6541 (N_6541,N_6358,N_6357);
xnor U6542 (N_6542,N_6222,N_6323);
xnor U6543 (N_6543,N_6395,N_6335);
and U6544 (N_6544,N_6209,N_6297);
nor U6545 (N_6545,N_6300,N_6326);
nand U6546 (N_6546,N_6312,N_6297);
or U6547 (N_6547,N_6302,N_6256);
nand U6548 (N_6548,N_6255,N_6221);
xor U6549 (N_6549,N_6369,N_6385);
and U6550 (N_6550,N_6284,N_6221);
or U6551 (N_6551,N_6348,N_6299);
xnor U6552 (N_6552,N_6235,N_6367);
nand U6553 (N_6553,N_6397,N_6373);
nor U6554 (N_6554,N_6358,N_6317);
nand U6555 (N_6555,N_6224,N_6287);
or U6556 (N_6556,N_6234,N_6220);
or U6557 (N_6557,N_6372,N_6228);
and U6558 (N_6558,N_6218,N_6289);
or U6559 (N_6559,N_6335,N_6253);
or U6560 (N_6560,N_6376,N_6355);
or U6561 (N_6561,N_6271,N_6224);
nand U6562 (N_6562,N_6264,N_6243);
nor U6563 (N_6563,N_6249,N_6238);
nor U6564 (N_6564,N_6289,N_6225);
and U6565 (N_6565,N_6313,N_6206);
and U6566 (N_6566,N_6216,N_6292);
nand U6567 (N_6567,N_6242,N_6308);
and U6568 (N_6568,N_6352,N_6353);
xnor U6569 (N_6569,N_6380,N_6296);
xnor U6570 (N_6570,N_6282,N_6313);
or U6571 (N_6571,N_6328,N_6288);
xnor U6572 (N_6572,N_6265,N_6343);
nor U6573 (N_6573,N_6296,N_6259);
or U6574 (N_6574,N_6315,N_6377);
or U6575 (N_6575,N_6232,N_6223);
nor U6576 (N_6576,N_6232,N_6322);
and U6577 (N_6577,N_6365,N_6358);
nor U6578 (N_6578,N_6210,N_6387);
xor U6579 (N_6579,N_6292,N_6357);
nand U6580 (N_6580,N_6234,N_6344);
and U6581 (N_6581,N_6226,N_6384);
nand U6582 (N_6582,N_6362,N_6317);
nor U6583 (N_6583,N_6210,N_6222);
and U6584 (N_6584,N_6225,N_6375);
nand U6585 (N_6585,N_6257,N_6225);
nor U6586 (N_6586,N_6278,N_6227);
nand U6587 (N_6587,N_6343,N_6264);
nor U6588 (N_6588,N_6271,N_6294);
xor U6589 (N_6589,N_6206,N_6200);
xor U6590 (N_6590,N_6355,N_6369);
nand U6591 (N_6591,N_6237,N_6388);
or U6592 (N_6592,N_6310,N_6338);
or U6593 (N_6593,N_6215,N_6235);
nor U6594 (N_6594,N_6396,N_6245);
nor U6595 (N_6595,N_6248,N_6230);
xnor U6596 (N_6596,N_6319,N_6380);
nor U6597 (N_6597,N_6338,N_6345);
or U6598 (N_6598,N_6372,N_6267);
and U6599 (N_6599,N_6330,N_6365);
and U6600 (N_6600,N_6467,N_6450);
or U6601 (N_6601,N_6518,N_6521);
nand U6602 (N_6602,N_6446,N_6526);
and U6603 (N_6603,N_6488,N_6429);
xor U6604 (N_6604,N_6577,N_6505);
or U6605 (N_6605,N_6563,N_6411);
nor U6606 (N_6606,N_6543,N_6567);
xnor U6607 (N_6607,N_6586,N_6455);
nand U6608 (N_6608,N_6581,N_6404);
nand U6609 (N_6609,N_6512,N_6513);
nand U6610 (N_6610,N_6540,N_6576);
or U6611 (N_6611,N_6527,N_6470);
nand U6612 (N_6612,N_6444,N_6568);
nor U6613 (N_6613,N_6412,N_6421);
nor U6614 (N_6614,N_6517,N_6515);
or U6615 (N_6615,N_6508,N_6566);
or U6616 (N_6616,N_6445,N_6495);
nor U6617 (N_6617,N_6432,N_6402);
and U6618 (N_6618,N_6558,N_6442);
nor U6619 (N_6619,N_6551,N_6514);
and U6620 (N_6620,N_6548,N_6587);
and U6621 (N_6621,N_6502,N_6538);
or U6622 (N_6622,N_6554,N_6487);
nand U6623 (N_6623,N_6418,N_6591);
and U6624 (N_6624,N_6426,N_6557);
nor U6625 (N_6625,N_6535,N_6499);
or U6626 (N_6626,N_6539,N_6441);
or U6627 (N_6627,N_6560,N_6520);
or U6628 (N_6628,N_6546,N_6572);
and U6629 (N_6629,N_6471,N_6585);
xnor U6630 (N_6630,N_6473,N_6435);
nor U6631 (N_6631,N_6489,N_6443);
or U6632 (N_6632,N_6523,N_6462);
nor U6633 (N_6633,N_6598,N_6498);
nor U6634 (N_6634,N_6465,N_6536);
nor U6635 (N_6635,N_6436,N_6510);
nor U6636 (N_6636,N_6413,N_6545);
nor U6637 (N_6637,N_6427,N_6434);
nor U6638 (N_6638,N_6478,N_6476);
xor U6639 (N_6639,N_6532,N_6420);
and U6640 (N_6640,N_6570,N_6579);
xor U6641 (N_6641,N_6564,N_6501);
or U6642 (N_6642,N_6593,N_6485);
xnor U6643 (N_6643,N_6425,N_6533);
or U6644 (N_6644,N_6561,N_6562);
nand U6645 (N_6645,N_6463,N_6438);
nor U6646 (N_6646,N_6490,N_6409);
nor U6647 (N_6647,N_6453,N_6522);
nor U6648 (N_6648,N_6492,N_6537);
xor U6649 (N_6649,N_6559,N_6422);
nand U6650 (N_6650,N_6497,N_6457);
or U6651 (N_6651,N_6507,N_6483);
nor U6652 (N_6652,N_6542,N_6575);
xor U6653 (N_6653,N_6550,N_6574);
nor U6654 (N_6654,N_6408,N_6400);
xor U6655 (N_6655,N_6415,N_6494);
nor U6656 (N_6656,N_6479,N_6549);
nand U6657 (N_6657,N_6484,N_6590);
or U6658 (N_6658,N_6430,N_6416);
nor U6659 (N_6659,N_6401,N_6503);
and U6660 (N_6660,N_6582,N_6461);
nor U6661 (N_6661,N_6524,N_6424);
nand U6662 (N_6662,N_6486,N_6583);
and U6663 (N_6663,N_6403,N_6530);
xnor U6664 (N_6664,N_6448,N_6477);
nand U6665 (N_6665,N_6595,N_6459);
and U6666 (N_6666,N_6410,N_6468);
and U6667 (N_6667,N_6589,N_6454);
nor U6668 (N_6668,N_6553,N_6584);
and U6669 (N_6669,N_6592,N_6580);
nor U6670 (N_6670,N_6547,N_6417);
nor U6671 (N_6671,N_6599,N_6588);
nand U6672 (N_6672,N_6491,N_6519);
and U6673 (N_6673,N_6474,N_6475);
xnor U6674 (N_6674,N_6528,N_6596);
nand U6675 (N_6675,N_6481,N_6597);
nor U6676 (N_6676,N_6516,N_6423);
nor U6677 (N_6677,N_6573,N_6496);
and U6678 (N_6678,N_6556,N_6525);
and U6679 (N_6679,N_6544,N_6439);
xnor U6680 (N_6680,N_6452,N_6458);
nand U6681 (N_6681,N_6406,N_6594);
or U6682 (N_6682,N_6482,N_6509);
or U6683 (N_6683,N_6469,N_6433);
nor U6684 (N_6684,N_6437,N_6464);
nor U6685 (N_6685,N_6447,N_6531);
nand U6686 (N_6686,N_6571,N_6456);
nand U6687 (N_6687,N_6440,N_6500);
nor U6688 (N_6688,N_6472,N_6555);
nor U6689 (N_6689,N_6449,N_6405);
nor U6690 (N_6690,N_6466,N_6414);
nand U6691 (N_6691,N_6506,N_6407);
nor U6692 (N_6692,N_6569,N_6460);
and U6693 (N_6693,N_6565,N_6534);
and U6694 (N_6694,N_6578,N_6431);
nand U6695 (N_6695,N_6419,N_6480);
nor U6696 (N_6696,N_6493,N_6552);
or U6697 (N_6697,N_6541,N_6529);
nor U6698 (N_6698,N_6504,N_6511);
nand U6699 (N_6699,N_6428,N_6451);
and U6700 (N_6700,N_6565,N_6559);
and U6701 (N_6701,N_6479,N_6415);
xor U6702 (N_6702,N_6443,N_6404);
and U6703 (N_6703,N_6585,N_6506);
and U6704 (N_6704,N_6403,N_6566);
or U6705 (N_6705,N_6469,N_6497);
and U6706 (N_6706,N_6511,N_6561);
nand U6707 (N_6707,N_6497,N_6437);
nand U6708 (N_6708,N_6483,N_6557);
xor U6709 (N_6709,N_6430,N_6588);
nand U6710 (N_6710,N_6407,N_6431);
or U6711 (N_6711,N_6485,N_6403);
or U6712 (N_6712,N_6480,N_6416);
xor U6713 (N_6713,N_6510,N_6475);
xnor U6714 (N_6714,N_6553,N_6508);
and U6715 (N_6715,N_6587,N_6478);
or U6716 (N_6716,N_6583,N_6549);
and U6717 (N_6717,N_6542,N_6552);
nor U6718 (N_6718,N_6441,N_6579);
nor U6719 (N_6719,N_6587,N_6474);
xor U6720 (N_6720,N_6574,N_6489);
xnor U6721 (N_6721,N_6474,N_6411);
nand U6722 (N_6722,N_6538,N_6580);
or U6723 (N_6723,N_6527,N_6469);
xnor U6724 (N_6724,N_6575,N_6493);
and U6725 (N_6725,N_6481,N_6595);
xor U6726 (N_6726,N_6536,N_6554);
and U6727 (N_6727,N_6490,N_6476);
xor U6728 (N_6728,N_6432,N_6547);
xnor U6729 (N_6729,N_6474,N_6537);
or U6730 (N_6730,N_6484,N_6465);
nand U6731 (N_6731,N_6567,N_6589);
nor U6732 (N_6732,N_6539,N_6583);
nand U6733 (N_6733,N_6568,N_6541);
nor U6734 (N_6734,N_6564,N_6578);
nand U6735 (N_6735,N_6572,N_6465);
xnor U6736 (N_6736,N_6518,N_6443);
nor U6737 (N_6737,N_6431,N_6446);
nand U6738 (N_6738,N_6505,N_6485);
nand U6739 (N_6739,N_6438,N_6503);
nor U6740 (N_6740,N_6451,N_6494);
and U6741 (N_6741,N_6447,N_6416);
xor U6742 (N_6742,N_6565,N_6401);
nand U6743 (N_6743,N_6409,N_6586);
nand U6744 (N_6744,N_6496,N_6581);
and U6745 (N_6745,N_6564,N_6488);
nor U6746 (N_6746,N_6418,N_6544);
or U6747 (N_6747,N_6411,N_6446);
nand U6748 (N_6748,N_6412,N_6516);
and U6749 (N_6749,N_6559,N_6403);
or U6750 (N_6750,N_6554,N_6438);
nor U6751 (N_6751,N_6414,N_6500);
nor U6752 (N_6752,N_6452,N_6447);
nand U6753 (N_6753,N_6547,N_6503);
nor U6754 (N_6754,N_6587,N_6533);
nor U6755 (N_6755,N_6488,N_6515);
xor U6756 (N_6756,N_6569,N_6400);
nor U6757 (N_6757,N_6409,N_6540);
or U6758 (N_6758,N_6491,N_6474);
nand U6759 (N_6759,N_6569,N_6451);
and U6760 (N_6760,N_6555,N_6557);
or U6761 (N_6761,N_6517,N_6537);
nor U6762 (N_6762,N_6463,N_6576);
or U6763 (N_6763,N_6433,N_6588);
xor U6764 (N_6764,N_6593,N_6586);
or U6765 (N_6765,N_6588,N_6522);
and U6766 (N_6766,N_6512,N_6545);
nor U6767 (N_6767,N_6527,N_6518);
xnor U6768 (N_6768,N_6451,N_6427);
nor U6769 (N_6769,N_6516,N_6538);
xnor U6770 (N_6770,N_6428,N_6537);
nor U6771 (N_6771,N_6479,N_6487);
or U6772 (N_6772,N_6480,N_6576);
and U6773 (N_6773,N_6510,N_6593);
or U6774 (N_6774,N_6440,N_6405);
nand U6775 (N_6775,N_6408,N_6540);
and U6776 (N_6776,N_6575,N_6503);
or U6777 (N_6777,N_6467,N_6590);
and U6778 (N_6778,N_6458,N_6597);
nor U6779 (N_6779,N_6509,N_6493);
xnor U6780 (N_6780,N_6586,N_6471);
nand U6781 (N_6781,N_6495,N_6430);
nand U6782 (N_6782,N_6437,N_6447);
nor U6783 (N_6783,N_6591,N_6567);
or U6784 (N_6784,N_6418,N_6593);
nor U6785 (N_6785,N_6528,N_6408);
nand U6786 (N_6786,N_6599,N_6403);
nor U6787 (N_6787,N_6486,N_6483);
and U6788 (N_6788,N_6521,N_6496);
nor U6789 (N_6789,N_6583,N_6526);
nand U6790 (N_6790,N_6437,N_6569);
or U6791 (N_6791,N_6532,N_6453);
nand U6792 (N_6792,N_6595,N_6439);
or U6793 (N_6793,N_6555,N_6519);
or U6794 (N_6794,N_6433,N_6506);
nor U6795 (N_6795,N_6504,N_6408);
and U6796 (N_6796,N_6505,N_6563);
xnor U6797 (N_6797,N_6587,N_6420);
or U6798 (N_6798,N_6433,N_6557);
and U6799 (N_6799,N_6510,N_6425);
nand U6800 (N_6800,N_6687,N_6634);
xnor U6801 (N_6801,N_6690,N_6702);
and U6802 (N_6802,N_6652,N_6654);
nor U6803 (N_6803,N_6734,N_6655);
or U6804 (N_6804,N_6642,N_6676);
nand U6805 (N_6805,N_6738,N_6675);
nor U6806 (N_6806,N_6605,N_6680);
or U6807 (N_6807,N_6693,N_6722);
xor U6808 (N_6808,N_6658,N_6685);
xor U6809 (N_6809,N_6647,N_6691);
nand U6810 (N_6810,N_6653,N_6705);
nor U6811 (N_6811,N_6783,N_6606);
nand U6812 (N_6812,N_6657,N_6700);
nand U6813 (N_6813,N_6768,N_6712);
nor U6814 (N_6814,N_6604,N_6711);
xnor U6815 (N_6815,N_6651,N_6744);
xor U6816 (N_6816,N_6731,N_6785);
or U6817 (N_6817,N_6784,N_6786);
nand U6818 (N_6818,N_6706,N_6639);
or U6819 (N_6819,N_6646,N_6670);
nand U6820 (N_6820,N_6696,N_6627);
nand U6821 (N_6821,N_6767,N_6750);
or U6822 (N_6822,N_6704,N_6796);
xnor U6823 (N_6823,N_6667,N_6751);
xor U6824 (N_6824,N_6659,N_6716);
xnor U6825 (N_6825,N_6773,N_6798);
or U6826 (N_6826,N_6656,N_6795);
nand U6827 (N_6827,N_6683,N_6678);
and U6828 (N_6828,N_6707,N_6650);
nor U6829 (N_6829,N_6752,N_6625);
or U6830 (N_6830,N_6692,N_6746);
nor U6831 (N_6831,N_6660,N_6788);
or U6832 (N_6832,N_6761,N_6643);
nor U6833 (N_6833,N_6753,N_6677);
and U6834 (N_6834,N_6635,N_6648);
or U6835 (N_6835,N_6719,N_6756);
and U6836 (N_6836,N_6760,N_6739);
nor U6837 (N_6837,N_6787,N_6717);
xor U6838 (N_6838,N_6776,N_6799);
and U6839 (N_6839,N_6727,N_6743);
and U6840 (N_6840,N_6794,N_6689);
and U6841 (N_6841,N_6622,N_6765);
xor U6842 (N_6842,N_6669,N_6758);
nor U6843 (N_6843,N_6694,N_6674);
xnor U6844 (N_6844,N_6615,N_6736);
or U6845 (N_6845,N_6699,N_6620);
nand U6846 (N_6846,N_6695,N_6777);
or U6847 (N_6847,N_6762,N_6609);
nand U6848 (N_6848,N_6772,N_6632);
nand U6849 (N_6849,N_6698,N_6733);
nand U6850 (N_6850,N_6684,N_6770);
xor U6851 (N_6851,N_6797,N_6621);
xnor U6852 (N_6852,N_6771,N_6721);
xor U6853 (N_6853,N_6637,N_6790);
nor U6854 (N_6854,N_6741,N_6671);
xnor U6855 (N_6855,N_6723,N_6710);
xnor U6856 (N_6856,N_6740,N_6729);
or U6857 (N_6857,N_6601,N_6616);
xnor U6858 (N_6858,N_6630,N_6737);
or U6859 (N_6859,N_6602,N_6775);
and U6860 (N_6860,N_6633,N_6612);
nand U6861 (N_6861,N_6666,N_6754);
nor U6862 (N_6862,N_6610,N_6611);
and U6863 (N_6863,N_6766,N_6640);
nand U6864 (N_6864,N_6782,N_6781);
xor U6865 (N_6865,N_6703,N_6681);
nor U6866 (N_6866,N_6638,N_6780);
nor U6867 (N_6867,N_6774,N_6701);
xor U6868 (N_6868,N_6728,N_6645);
nand U6869 (N_6869,N_6789,N_6600);
xor U6870 (N_6870,N_6608,N_6749);
nand U6871 (N_6871,N_6715,N_6618);
nor U6872 (N_6872,N_6730,N_6614);
and U6873 (N_6873,N_6668,N_6623);
and U6874 (N_6874,N_6726,N_6742);
xnor U6875 (N_6875,N_6673,N_6763);
nor U6876 (N_6876,N_6755,N_6603);
nor U6877 (N_6877,N_6631,N_6713);
and U6878 (N_6878,N_6748,N_6661);
nand U6879 (N_6879,N_6613,N_6665);
or U6880 (N_6880,N_6663,N_6629);
and U6881 (N_6881,N_6714,N_6791);
nand U6882 (N_6882,N_6641,N_6686);
or U6883 (N_6883,N_6724,N_6697);
xor U6884 (N_6884,N_6607,N_6626);
or U6885 (N_6885,N_6778,N_6732);
and U6886 (N_6886,N_6725,N_6682);
nor U6887 (N_6887,N_6757,N_6708);
nand U6888 (N_6888,N_6720,N_6764);
and U6889 (N_6889,N_6644,N_6747);
and U6890 (N_6890,N_6649,N_6636);
nand U6891 (N_6891,N_6662,N_6745);
nor U6892 (N_6892,N_6735,N_6688);
or U6893 (N_6893,N_6672,N_6792);
nand U6894 (N_6894,N_6628,N_6617);
or U6895 (N_6895,N_6779,N_6619);
nand U6896 (N_6896,N_6709,N_6679);
nor U6897 (N_6897,N_6793,N_6769);
or U6898 (N_6898,N_6624,N_6718);
nand U6899 (N_6899,N_6759,N_6664);
and U6900 (N_6900,N_6693,N_6642);
nor U6901 (N_6901,N_6692,N_6666);
or U6902 (N_6902,N_6764,N_6747);
and U6903 (N_6903,N_6690,N_6782);
xnor U6904 (N_6904,N_6617,N_6727);
and U6905 (N_6905,N_6637,N_6635);
and U6906 (N_6906,N_6771,N_6617);
and U6907 (N_6907,N_6785,N_6708);
nand U6908 (N_6908,N_6683,N_6693);
or U6909 (N_6909,N_6759,N_6685);
nand U6910 (N_6910,N_6690,N_6614);
or U6911 (N_6911,N_6784,N_6641);
and U6912 (N_6912,N_6763,N_6685);
or U6913 (N_6913,N_6691,N_6792);
or U6914 (N_6914,N_6773,N_6693);
nor U6915 (N_6915,N_6651,N_6721);
xor U6916 (N_6916,N_6713,N_6718);
nand U6917 (N_6917,N_6633,N_6673);
nor U6918 (N_6918,N_6631,N_6797);
and U6919 (N_6919,N_6615,N_6690);
nor U6920 (N_6920,N_6797,N_6666);
xnor U6921 (N_6921,N_6603,N_6781);
and U6922 (N_6922,N_6619,N_6707);
or U6923 (N_6923,N_6706,N_6646);
xor U6924 (N_6924,N_6600,N_6684);
or U6925 (N_6925,N_6764,N_6609);
xor U6926 (N_6926,N_6736,N_6794);
xor U6927 (N_6927,N_6625,N_6740);
xnor U6928 (N_6928,N_6623,N_6680);
xnor U6929 (N_6929,N_6781,N_6633);
xnor U6930 (N_6930,N_6778,N_6635);
nand U6931 (N_6931,N_6792,N_6640);
xor U6932 (N_6932,N_6697,N_6695);
nand U6933 (N_6933,N_6729,N_6731);
nor U6934 (N_6934,N_6602,N_6797);
or U6935 (N_6935,N_6632,N_6614);
or U6936 (N_6936,N_6661,N_6782);
xor U6937 (N_6937,N_6627,N_6779);
nand U6938 (N_6938,N_6636,N_6697);
xor U6939 (N_6939,N_6695,N_6763);
or U6940 (N_6940,N_6656,N_6681);
xor U6941 (N_6941,N_6766,N_6637);
or U6942 (N_6942,N_6663,N_6665);
nor U6943 (N_6943,N_6644,N_6619);
and U6944 (N_6944,N_6640,N_6681);
or U6945 (N_6945,N_6651,N_6766);
xnor U6946 (N_6946,N_6728,N_6661);
xnor U6947 (N_6947,N_6604,N_6728);
and U6948 (N_6948,N_6610,N_6680);
nand U6949 (N_6949,N_6703,N_6763);
and U6950 (N_6950,N_6771,N_6601);
xor U6951 (N_6951,N_6724,N_6645);
nand U6952 (N_6952,N_6718,N_6665);
and U6953 (N_6953,N_6675,N_6623);
nand U6954 (N_6954,N_6718,N_6705);
nor U6955 (N_6955,N_6723,N_6769);
xor U6956 (N_6956,N_6749,N_6694);
nand U6957 (N_6957,N_6756,N_6600);
nor U6958 (N_6958,N_6698,N_6762);
xnor U6959 (N_6959,N_6789,N_6788);
nor U6960 (N_6960,N_6604,N_6701);
nor U6961 (N_6961,N_6649,N_6629);
and U6962 (N_6962,N_6615,N_6633);
nand U6963 (N_6963,N_6720,N_6633);
xor U6964 (N_6964,N_6744,N_6762);
nor U6965 (N_6965,N_6707,N_6794);
nand U6966 (N_6966,N_6641,N_6623);
nand U6967 (N_6967,N_6691,N_6796);
or U6968 (N_6968,N_6624,N_6746);
nor U6969 (N_6969,N_6694,N_6621);
or U6970 (N_6970,N_6682,N_6633);
xor U6971 (N_6971,N_6706,N_6746);
or U6972 (N_6972,N_6691,N_6634);
or U6973 (N_6973,N_6711,N_6702);
and U6974 (N_6974,N_6725,N_6758);
nor U6975 (N_6975,N_6689,N_6734);
nor U6976 (N_6976,N_6796,N_6617);
and U6977 (N_6977,N_6783,N_6671);
xor U6978 (N_6978,N_6642,N_6783);
xnor U6979 (N_6979,N_6782,N_6676);
xnor U6980 (N_6980,N_6788,N_6625);
or U6981 (N_6981,N_6613,N_6788);
nand U6982 (N_6982,N_6635,N_6679);
and U6983 (N_6983,N_6792,N_6687);
nor U6984 (N_6984,N_6607,N_6668);
or U6985 (N_6985,N_6628,N_6727);
nor U6986 (N_6986,N_6655,N_6700);
xor U6987 (N_6987,N_6799,N_6613);
xnor U6988 (N_6988,N_6631,N_6767);
or U6989 (N_6989,N_6767,N_6788);
nand U6990 (N_6990,N_6729,N_6719);
nand U6991 (N_6991,N_6676,N_6680);
nor U6992 (N_6992,N_6647,N_6632);
nand U6993 (N_6993,N_6607,N_6726);
xor U6994 (N_6994,N_6727,N_6771);
xor U6995 (N_6995,N_6690,N_6713);
xnor U6996 (N_6996,N_6672,N_6666);
nand U6997 (N_6997,N_6600,N_6740);
nand U6998 (N_6998,N_6764,N_6625);
and U6999 (N_6999,N_6720,N_6760);
nor U7000 (N_7000,N_6850,N_6970);
nand U7001 (N_7001,N_6994,N_6864);
and U7002 (N_7002,N_6833,N_6805);
nand U7003 (N_7003,N_6937,N_6809);
xor U7004 (N_7004,N_6844,N_6847);
or U7005 (N_7005,N_6973,N_6999);
or U7006 (N_7006,N_6991,N_6961);
xor U7007 (N_7007,N_6915,N_6884);
xor U7008 (N_7008,N_6846,N_6802);
and U7009 (N_7009,N_6814,N_6877);
xnor U7010 (N_7010,N_6906,N_6856);
and U7011 (N_7011,N_6863,N_6965);
xnor U7012 (N_7012,N_6917,N_6879);
nand U7013 (N_7013,N_6963,N_6807);
nor U7014 (N_7014,N_6813,N_6874);
or U7015 (N_7015,N_6876,N_6916);
and U7016 (N_7016,N_6895,N_6981);
or U7017 (N_7017,N_6966,N_6839);
nand U7018 (N_7018,N_6815,N_6806);
and U7019 (N_7019,N_6854,N_6891);
nor U7020 (N_7020,N_6931,N_6822);
xnor U7021 (N_7021,N_6871,N_6812);
xnor U7022 (N_7022,N_6945,N_6949);
or U7023 (N_7023,N_6942,N_6845);
or U7024 (N_7024,N_6926,N_6925);
nor U7025 (N_7025,N_6861,N_6941);
xor U7026 (N_7026,N_6971,N_6817);
or U7027 (N_7027,N_6972,N_6921);
nor U7028 (N_7028,N_6886,N_6855);
xnor U7029 (N_7029,N_6857,N_6920);
nor U7030 (N_7030,N_6842,N_6964);
nand U7031 (N_7031,N_6952,N_6902);
nor U7032 (N_7032,N_6859,N_6858);
xor U7033 (N_7033,N_6848,N_6948);
nand U7034 (N_7034,N_6967,N_6865);
or U7035 (N_7035,N_6830,N_6800);
nand U7036 (N_7036,N_6862,N_6831);
and U7037 (N_7037,N_6824,N_6987);
and U7038 (N_7038,N_6960,N_6943);
nor U7039 (N_7039,N_6982,N_6976);
and U7040 (N_7040,N_6889,N_6903);
xnor U7041 (N_7041,N_6868,N_6985);
nor U7042 (N_7042,N_6881,N_6899);
nand U7043 (N_7043,N_6922,N_6810);
and U7044 (N_7044,N_6969,N_6837);
nor U7045 (N_7045,N_6892,N_6979);
xnor U7046 (N_7046,N_6808,N_6897);
and U7047 (N_7047,N_6940,N_6811);
nor U7048 (N_7048,N_6851,N_6829);
or U7049 (N_7049,N_6935,N_6957);
xnor U7050 (N_7050,N_6992,N_6927);
xor U7051 (N_7051,N_6988,N_6959);
nor U7052 (N_7052,N_6888,N_6853);
and U7053 (N_7053,N_6849,N_6984);
and U7054 (N_7054,N_6803,N_6880);
nand U7055 (N_7055,N_6989,N_6983);
and U7056 (N_7056,N_6947,N_6887);
and U7057 (N_7057,N_6905,N_6914);
and U7058 (N_7058,N_6896,N_6997);
nor U7059 (N_7059,N_6913,N_6951);
xor U7060 (N_7060,N_6993,N_6866);
nand U7061 (N_7061,N_6954,N_6990);
and U7062 (N_7062,N_6933,N_6873);
and U7063 (N_7063,N_6827,N_6835);
xor U7064 (N_7064,N_6978,N_6924);
xnor U7065 (N_7065,N_6804,N_6834);
xor U7066 (N_7066,N_6878,N_6962);
or U7067 (N_7067,N_6826,N_6828);
nand U7068 (N_7068,N_6801,N_6843);
or U7069 (N_7069,N_6820,N_6898);
nand U7070 (N_7070,N_6919,N_6908);
or U7071 (N_7071,N_6821,N_6840);
and U7072 (N_7072,N_6841,N_6818);
or U7073 (N_7073,N_6883,N_6977);
nor U7074 (N_7074,N_6869,N_6956);
or U7075 (N_7075,N_6907,N_6932);
and U7076 (N_7076,N_6836,N_6901);
and U7077 (N_7077,N_6838,N_6852);
nor U7078 (N_7078,N_6998,N_6909);
or U7079 (N_7079,N_6934,N_6819);
xnor U7080 (N_7080,N_6928,N_6867);
nor U7081 (N_7081,N_6953,N_6939);
and U7082 (N_7082,N_6946,N_6816);
or U7083 (N_7083,N_6870,N_6955);
and U7084 (N_7084,N_6923,N_6825);
xnor U7085 (N_7085,N_6995,N_6950);
xor U7086 (N_7086,N_6894,N_6938);
or U7087 (N_7087,N_6912,N_6930);
nor U7088 (N_7088,N_6918,N_6996);
nand U7089 (N_7089,N_6986,N_6890);
xor U7090 (N_7090,N_6974,N_6911);
xor U7091 (N_7091,N_6980,N_6944);
or U7092 (N_7092,N_6904,N_6872);
nand U7093 (N_7093,N_6823,N_6875);
nand U7094 (N_7094,N_6929,N_6958);
or U7095 (N_7095,N_6975,N_6832);
nand U7096 (N_7096,N_6910,N_6893);
nand U7097 (N_7097,N_6936,N_6885);
or U7098 (N_7098,N_6900,N_6860);
xnor U7099 (N_7099,N_6968,N_6882);
or U7100 (N_7100,N_6920,N_6808);
nor U7101 (N_7101,N_6852,N_6844);
nor U7102 (N_7102,N_6901,N_6944);
xor U7103 (N_7103,N_6819,N_6915);
xnor U7104 (N_7104,N_6827,N_6836);
nor U7105 (N_7105,N_6897,N_6835);
nand U7106 (N_7106,N_6875,N_6864);
nor U7107 (N_7107,N_6818,N_6930);
xor U7108 (N_7108,N_6879,N_6874);
and U7109 (N_7109,N_6971,N_6888);
nor U7110 (N_7110,N_6976,N_6939);
nor U7111 (N_7111,N_6854,N_6864);
nor U7112 (N_7112,N_6881,N_6925);
nor U7113 (N_7113,N_6861,N_6919);
nor U7114 (N_7114,N_6867,N_6903);
or U7115 (N_7115,N_6892,N_6807);
xnor U7116 (N_7116,N_6962,N_6966);
nor U7117 (N_7117,N_6902,N_6960);
and U7118 (N_7118,N_6959,N_6935);
nand U7119 (N_7119,N_6864,N_6957);
and U7120 (N_7120,N_6883,N_6944);
or U7121 (N_7121,N_6871,N_6994);
nand U7122 (N_7122,N_6852,N_6865);
nor U7123 (N_7123,N_6803,N_6902);
nor U7124 (N_7124,N_6928,N_6917);
or U7125 (N_7125,N_6932,N_6809);
nand U7126 (N_7126,N_6966,N_6941);
and U7127 (N_7127,N_6899,N_6851);
xor U7128 (N_7128,N_6867,N_6817);
nor U7129 (N_7129,N_6812,N_6984);
and U7130 (N_7130,N_6829,N_6904);
nor U7131 (N_7131,N_6976,N_6928);
and U7132 (N_7132,N_6940,N_6997);
or U7133 (N_7133,N_6870,N_6863);
xnor U7134 (N_7134,N_6957,N_6868);
and U7135 (N_7135,N_6909,N_6958);
xor U7136 (N_7136,N_6982,N_6967);
nor U7137 (N_7137,N_6864,N_6800);
or U7138 (N_7138,N_6940,N_6847);
xnor U7139 (N_7139,N_6864,N_6956);
nand U7140 (N_7140,N_6839,N_6915);
nand U7141 (N_7141,N_6980,N_6836);
and U7142 (N_7142,N_6950,N_6997);
nand U7143 (N_7143,N_6973,N_6807);
nand U7144 (N_7144,N_6853,N_6902);
nand U7145 (N_7145,N_6828,N_6893);
or U7146 (N_7146,N_6815,N_6865);
and U7147 (N_7147,N_6988,N_6804);
nand U7148 (N_7148,N_6936,N_6925);
xor U7149 (N_7149,N_6869,N_6901);
xnor U7150 (N_7150,N_6859,N_6949);
xor U7151 (N_7151,N_6885,N_6812);
nand U7152 (N_7152,N_6840,N_6823);
xor U7153 (N_7153,N_6950,N_6817);
or U7154 (N_7154,N_6999,N_6840);
xnor U7155 (N_7155,N_6854,N_6899);
or U7156 (N_7156,N_6934,N_6935);
or U7157 (N_7157,N_6977,N_6891);
or U7158 (N_7158,N_6862,N_6996);
or U7159 (N_7159,N_6872,N_6964);
and U7160 (N_7160,N_6986,N_6984);
or U7161 (N_7161,N_6810,N_6888);
xnor U7162 (N_7162,N_6847,N_6843);
or U7163 (N_7163,N_6953,N_6880);
xor U7164 (N_7164,N_6918,N_6898);
nor U7165 (N_7165,N_6845,N_6992);
nand U7166 (N_7166,N_6901,N_6852);
or U7167 (N_7167,N_6926,N_6811);
nor U7168 (N_7168,N_6883,N_6987);
nor U7169 (N_7169,N_6935,N_6931);
or U7170 (N_7170,N_6990,N_6830);
and U7171 (N_7171,N_6947,N_6900);
nand U7172 (N_7172,N_6944,N_6808);
or U7173 (N_7173,N_6915,N_6828);
nand U7174 (N_7174,N_6944,N_6963);
or U7175 (N_7175,N_6813,N_6839);
xnor U7176 (N_7176,N_6845,N_6931);
and U7177 (N_7177,N_6878,N_6933);
xor U7178 (N_7178,N_6988,N_6971);
xnor U7179 (N_7179,N_6914,N_6989);
or U7180 (N_7180,N_6829,N_6818);
and U7181 (N_7181,N_6831,N_6854);
xor U7182 (N_7182,N_6870,N_6885);
nor U7183 (N_7183,N_6922,N_6967);
and U7184 (N_7184,N_6921,N_6906);
or U7185 (N_7185,N_6900,N_6964);
xnor U7186 (N_7186,N_6879,N_6979);
and U7187 (N_7187,N_6901,N_6980);
or U7188 (N_7188,N_6988,N_6897);
xnor U7189 (N_7189,N_6833,N_6994);
nor U7190 (N_7190,N_6966,N_6903);
nor U7191 (N_7191,N_6865,N_6825);
nor U7192 (N_7192,N_6851,N_6917);
nand U7193 (N_7193,N_6858,N_6830);
and U7194 (N_7194,N_6834,N_6863);
and U7195 (N_7195,N_6801,N_6987);
and U7196 (N_7196,N_6946,N_6818);
nand U7197 (N_7197,N_6976,N_6869);
nor U7198 (N_7198,N_6841,N_6968);
and U7199 (N_7199,N_6885,N_6862);
and U7200 (N_7200,N_7146,N_7083);
xnor U7201 (N_7201,N_7174,N_7089);
xor U7202 (N_7202,N_7004,N_7065);
or U7203 (N_7203,N_7030,N_7123);
xnor U7204 (N_7204,N_7061,N_7182);
nand U7205 (N_7205,N_7148,N_7104);
and U7206 (N_7206,N_7059,N_7100);
nor U7207 (N_7207,N_7190,N_7181);
nor U7208 (N_7208,N_7093,N_7041);
xor U7209 (N_7209,N_7109,N_7192);
xor U7210 (N_7210,N_7145,N_7157);
or U7211 (N_7211,N_7124,N_7026);
or U7212 (N_7212,N_7127,N_7150);
nor U7213 (N_7213,N_7153,N_7135);
xnor U7214 (N_7214,N_7014,N_7022);
and U7215 (N_7215,N_7169,N_7168);
and U7216 (N_7216,N_7062,N_7121);
nor U7217 (N_7217,N_7177,N_7042);
nand U7218 (N_7218,N_7043,N_7185);
and U7219 (N_7219,N_7032,N_7141);
xor U7220 (N_7220,N_7165,N_7092);
xnor U7221 (N_7221,N_7134,N_7113);
and U7222 (N_7222,N_7112,N_7198);
or U7223 (N_7223,N_7197,N_7051);
and U7224 (N_7224,N_7082,N_7088);
or U7225 (N_7225,N_7094,N_7117);
and U7226 (N_7226,N_7147,N_7012);
nand U7227 (N_7227,N_7005,N_7195);
or U7228 (N_7228,N_7008,N_7036);
xor U7229 (N_7229,N_7095,N_7047);
and U7230 (N_7230,N_7018,N_7154);
or U7231 (N_7231,N_7015,N_7156);
or U7232 (N_7232,N_7184,N_7140);
nand U7233 (N_7233,N_7081,N_7007);
and U7234 (N_7234,N_7163,N_7143);
nor U7235 (N_7235,N_7180,N_7063);
or U7236 (N_7236,N_7001,N_7045);
nand U7237 (N_7237,N_7017,N_7070);
xnor U7238 (N_7238,N_7085,N_7137);
or U7239 (N_7239,N_7126,N_7175);
and U7240 (N_7240,N_7166,N_7087);
and U7241 (N_7241,N_7131,N_7039);
or U7242 (N_7242,N_7074,N_7171);
nor U7243 (N_7243,N_7139,N_7172);
nor U7244 (N_7244,N_7019,N_7097);
nand U7245 (N_7245,N_7099,N_7013);
or U7246 (N_7246,N_7176,N_7102);
or U7247 (N_7247,N_7064,N_7114);
and U7248 (N_7248,N_7052,N_7132);
nand U7249 (N_7249,N_7167,N_7024);
and U7250 (N_7250,N_7084,N_7162);
or U7251 (N_7251,N_7038,N_7077);
nand U7252 (N_7252,N_7155,N_7069);
nand U7253 (N_7253,N_7129,N_7189);
and U7254 (N_7254,N_7199,N_7073);
or U7255 (N_7255,N_7053,N_7055);
or U7256 (N_7256,N_7149,N_7193);
and U7257 (N_7257,N_7009,N_7011);
xor U7258 (N_7258,N_7118,N_7152);
nand U7259 (N_7259,N_7159,N_7002);
xor U7260 (N_7260,N_7098,N_7142);
nor U7261 (N_7261,N_7136,N_7016);
xor U7262 (N_7262,N_7196,N_7031);
nor U7263 (N_7263,N_7071,N_7133);
and U7264 (N_7264,N_7068,N_7173);
or U7265 (N_7265,N_7080,N_7090);
and U7266 (N_7266,N_7108,N_7058);
xor U7267 (N_7267,N_7086,N_7122);
and U7268 (N_7268,N_7183,N_7194);
and U7269 (N_7269,N_7158,N_7048);
xnor U7270 (N_7270,N_7120,N_7054);
xor U7271 (N_7271,N_7107,N_7105);
nor U7272 (N_7272,N_7056,N_7191);
xor U7273 (N_7273,N_7021,N_7091);
or U7274 (N_7274,N_7067,N_7101);
and U7275 (N_7275,N_7078,N_7046);
xor U7276 (N_7276,N_7006,N_7186);
or U7277 (N_7277,N_7057,N_7040);
nor U7278 (N_7278,N_7044,N_7034);
or U7279 (N_7279,N_7144,N_7125);
nor U7280 (N_7280,N_7111,N_7066);
nand U7281 (N_7281,N_7119,N_7025);
or U7282 (N_7282,N_7110,N_7033);
nand U7283 (N_7283,N_7106,N_7187);
or U7284 (N_7284,N_7096,N_7023);
and U7285 (N_7285,N_7079,N_7050);
xnor U7286 (N_7286,N_7160,N_7115);
or U7287 (N_7287,N_7020,N_7049);
xnor U7288 (N_7288,N_7178,N_7161);
xnor U7289 (N_7289,N_7010,N_7072);
nor U7290 (N_7290,N_7000,N_7138);
xor U7291 (N_7291,N_7164,N_7103);
and U7292 (N_7292,N_7060,N_7027);
nor U7293 (N_7293,N_7028,N_7179);
or U7294 (N_7294,N_7128,N_7188);
xor U7295 (N_7295,N_7037,N_7003);
nor U7296 (N_7296,N_7029,N_7075);
and U7297 (N_7297,N_7076,N_7151);
nor U7298 (N_7298,N_7116,N_7035);
nor U7299 (N_7299,N_7130,N_7170);
nor U7300 (N_7300,N_7139,N_7123);
or U7301 (N_7301,N_7191,N_7028);
xor U7302 (N_7302,N_7034,N_7115);
xnor U7303 (N_7303,N_7112,N_7073);
and U7304 (N_7304,N_7011,N_7172);
and U7305 (N_7305,N_7029,N_7042);
and U7306 (N_7306,N_7063,N_7076);
nor U7307 (N_7307,N_7127,N_7183);
and U7308 (N_7308,N_7121,N_7059);
and U7309 (N_7309,N_7132,N_7033);
or U7310 (N_7310,N_7009,N_7160);
or U7311 (N_7311,N_7123,N_7067);
and U7312 (N_7312,N_7140,N_7078);
nor U7313 (N_7313,N_7045,N_7131);
or U7314 (N_7314,N_7151,N_7106);
or U7315 (N_7315,N_7071,N_7039);
xnor U7316 (N_7316,N_7025,N_7177);
nand U7317 (N_7317,N_7093,N_7028);
or U7318 (N_7318,N_7072,N_7030);
and U7319 (N_7319,N_7059,N_7094);
and U7320 (N_7320,N_7155,N_7071);
and U7321 (N_7321,N_7197,N_7036);
xnor U7322 (N_7322,N_7100,N_7058);
nand U7323 (N_7323,N_7177,N_7007);
or U7324 (N_7324,N_7092,N_7002);
xnor U7325 (N_7325,N_7004,N_7163);
and U7326 (N_7326,N_7080,N_7198);
and U7327 (N_7327,N_7124,N_7051);
nand U7328 (N_7328,N_7176,N_7060);
nor U7329 (N_7329,N_7088,N_7152);
or U7330 (N_7330,N_7119,N_7174);
and U7331 (N_7331,N_7060,N_7022);
xnor U7332 (N_7332,N_7159,N_7029);
nor U7333 (N_7333,N_7095,N_7063);
and U7334 (N_7334,N_7165,N_7046);
and U7335 (N_7335,N_7034,N_7099);
or U7336 (N_7336,N_7029,N_7027);
and U7337 (N_7337,N_7051,N_7049);
and U7338 (N_7338,N_7107,N_7073);
nand U7339 (N_7339,N_7092,N_7164);
nand U7340 (N_7340,N_7091,N_7001);
xnor U7341 (N_7341,N_7180,N_7108);
and U7342 (N_7342,N_7028,N_7196);
xnor U7343 (N_7343,N_7114,N_7009);
xnor U7344 (N_7344,N_7133,N_7171);
nand U7345 (N_7345,N_7048,N_7116);
or U7346 (N_7346,N_7185,N_7121);
nor U7347 (N_7347,N_7051,N_7133);
nor U7348 (N_7348,N_7113,N_7132);
nand U7349 (N_7349,N_7030,N_7055);
or U7350 (N_7350,N_7019,N_7096);
nor U7351 (N_7351,N_7117,N_7138);
or U7352 (N_7352,N_7001,N_7004);
nor U7353 (N_7353,N_7150,N_7105);
xor U7354 (N_7354,N_7199,N_7102);
and U7355 (N_7355,N_7008,N_7046);
xnor U7356 (N_7356,N_7094,N_7156);
nand U7357 (N_7357,N_7170,N_7057);
and U7358 (N_7358,N_7045,N_7130);
nor U7359 (N_7359,N_7151,N_7154);
nand U7360 (N_7360,N_7115,N_7179);
nor U7361 (N_7361,N_7134,N_7170);
nor U7362 (N_7362,N_7142,N_7139);
or U7363 (N_7363,N_7105,N_7026);
nor U7364 (N_7364,N_7128,N_7180);
xor U7365 (N_7365,N_7176,N_7042);
nand U7366 (N_7366,N_7153,N_7191);
or U7367 (N_7367,N_7108,N_7119);
and U7368 (N_7368,N_7044,N_7124);
nand U7369 (N_7369,N_7141,N_7121);
or U7370 (N_7370,N_7186,N_7188);
and U7371 (N_7371,N_7046,N_7118);
nor U7372 (N_7372,N_7167,N_7022);
nor U7373 (N_7373,N_7015,N_7104);
nand U7374 (N_7374,N_7178,N_7045);
nor U7375 (N_7375,N_7146,N_7044);
or U7376 (N_7376,N_7187,N_7140);
xnor U7377 (N_7377,N_7159,N_7174);
or U7378 (N_7378,N_7060,N_7061);
or U7379 (N_7379,N_7049,N_7113);
and U7380 (N_7380,N_7119,N_7125);
or U7381 (N_7381,N_7131,N_7109);
nor U7382 (N_7382,N_7071,N_7108);
and U7383 (N_7383,N_7151,N_7191);
nand U7384 (N_7384,N_7095,N_7154);
nor U7385 (N_7385,N_7124,N_7014);
nand U7386 (N_7386,N_7135,N_7182);
nand U7387 (N_7387,N_7192,N_7101);
or U7388 (N_7388,N_7122,N_7145);
or U7389 (N_7389,N_7158,N_7070);
and U7390 (N_7390,N_7045,N_7039);
and U7391 (N_7391,N_7074,N_7060);
xnor U7392 (N_7392,N_7061,N_7154);
nor U7393 (N_7393,N_7027,N_7023);
or U7394 (N_7394,N_7151,N_7034);
xnor U7395 (N_7395,N_7099,N_7087);
xnor U7396 (N_7396,N_7073,N_7058);
nor U7397 (N_7397,N_7097,N_7074);
nor U7398 (N_7398,N_7096,N_7025);
or U7399 (N_7399,N_7016,N_7178);
and U7400 (N_7400,N_7346,N_7320);
nor U7401 (N_7401,N_7214,N_7205);
or U7402 (N_7402,N_7302,N_7212);
nand U7403 (N_7403,N_7246,N_7343);
nand U7404 (N_7404,N_7216,N_7224);
nor U7405 (N_7405,N_7209,N_7325);
xnor U7406 (N_7406,N_7338,N_7377);
xnor U7407 (N_7407,N_7335,N_7387);
nand U7408 (N_7408,N_7311,N_7220);
nand U7409 (N_7409,N_7319,N_7266);
nor U7410 (N_7410,N_7213,N_7250);
nor U7411 (N_7411,N_7221,N_7210);
nand U7412 (N_7412,N_7299,N_7301);
and U7413 (N_7413,N_7310,N_7340);
or U7414 (N_7414,N_7264,N_7217);
xnor U7415 (N_7415,N_7358,N_7206);
nand U7416 (N_7416,N_7288,N_7287);
and U7417 (N_7417,N_7295,N_7394);
nand U7418 (N_7418,N_7279,N_7380);
nand U7419 (N_7419,N_7373,N_7366);
xor U7420 (N_7420,N_7370,N_7379);
xor U7421 (N_7421,N_7258,N_7284);
or U7422 (N_7422,N_7262,N_7291);
nor U7423 (N_7423,N_7215,N_7203);
or U7424 (N_7424,N_7344,N_7354);
nor U7425 (N_7425,N_7393,N_7378);
xor U7426 (N_7426,N_7290,N_7316);
nand U7427 (N_7427,N_7238,N_7371);
xnor U7428 (N_7428,N_7225,N_7355);
or U7429 (N_7429,N_7236,N_7244);
nand U7430 (N_7430,N_7322,N_7294);
nand U7431 (N_7431,N_7336,N_7383);
xor U7432 (N_7432,N_7324,N_7384);
and U7433 (N_7433,N_7234,N_7326);
nand U7434 (N_7434,N_7265,N_7286);
nor U7435 (N_7435,N_7235,N_7261);
xor U7436 (N_7436,N_7327,N_7204);
nand U7437 (N_7437,N_7259,N_7201);
nor U7438 (N_7438,N_7334,N_7277);
xnor U7439 (N_7439,N_7362,N_7218);
nand U7440 (N_7440,N_7247,N_7226);
nor U7441 (N_7441,N_7278,N_7321);
nor U7442 (N_7442,N_7388,N_7252);
xor U7443 (N_7443,N_7271,N_7254);
nor U7444 (N_7444,N_7331,N_7398);
nor U7445 (N_7445,N_7328,N_7323);
nand U7446 (N_7446,N_7267,N_7351);
xor U7447 (N_7447,N_7219,N_7240);
and U7448 (N_7448,N_7245,N_7239);
or U7449 (N_7449,N_7348,N_7395);
nand U7450 (N_7450,N_7298,N_7272);
or U7451 (N_7451,N_7303,N_7332);
nor U7452 (N_7452,N_7280,N_7337);
and U7453 (N_7453,N_7318,N_7367);
xor U7454 (N_7454,N_7296,N_7274);
nand U7455 (N_7455,N_7309,N_7306);
nand U7456 (N_7456,N_7372,N_7202);
nand U7457 (N_7457,N_7200,N_7356);
xor U7458 (N_7458,N_7232,N_7313);
and U7459 (N_7459,N_7256,N_7281);
nor U7460 (N_7460,N_7375,N_7263);
and U7461 (N_7461,N_7268,N_7282);
and U7462 (N_7462,N_7231,N_7386);
or U7463 (N_7463,N_7315,N_7364);
nor U7464 (N_7464,N_7369,N_7374);
xor U7465 (N_7465,N_7365,N_7211);
or U7466 (N_7466,N_7307,N_7243);
nand U7467 (N_7467,N_7260,N_7249);
nand U7468 (N_7468,N_7251,N_7352);
xor U7469 (N_7469,N_7359,N_7391);
nor U7470 (N_7470,N_7222,N_7349);
and U7471 (N_7471,N_7233,N_7330);
and U7472 (N_7472,N_7360,N_7257);
or U7473 (N_7473,N_7382,N_7289);
and U7474 (N_7474,N_7230,N_7385);
or U7475 (N_7475,N_7253,N_7275);
or U7476 (N_7476,N_7361,N_7329);
nor U7477 (N_7477,N_7223,N_7357);
nand U7478 (N_7478,N_7341,N_7363);
and U7479 (N_7479,N_7345,N_7397);
or U7480 (N_7480,N_7300,N_7207);
or U7481 (N_7481,N_7270,N_7376);
nor U7482 (N_7482,N_7227,N_7392);
and U7483 (N_7483,N_7276,N_7339);
and U7484 (N_7484,N_7350,N_7208);
xor U7485 (N_7485,N_7292,N_7242);
nand U7486 (N_7486,N_7368,N_7228);
xor U7487 (N_7487,N_7399,N_7283);
and U7488 (N_7488,N_7333,N_7269);
nand U7489 (N_7489,N_7237,N_7342);
and U7490 (N_7490,N_7293,N_7347);
xnor U7491 (N_7491,N_7241,N_7317);
xnor U7492 (N_7492,N_7229,N_7248);
nor U7493 (N_7493,N_7305,N_7390);
nand U7494 (N_7494,N_7273,N_7304);
nand U7495 (N_7495,N_7389,N_7312);
nor U7496 (N_7496,N_7285,N_7396);
xor U7497 (N_7497,N_7297,N_7308);
or U7498 (N_7498,N_7381,N_7353);
or U7499 (N_7499,N_7314,N_7255);
nor U7500 (N_7500,N_7261,N_7221);
nand U7501 (N_7501,N_7369,N_7390);
xor U7502 (N_7502,N_7343,N_7258);
and U7503 (N_7503,N_7311,N_7258);
or U7504 (N_7504,N_7270,N_7311);
xnor U7505 (N_7505,N_7223,N_7387);
and U7506 (N_7506,N_7276,N_7285);
or U7507 (N_7507,N_7350,N_7318);
nand U7508 (N_7508,N_7357,N_7299);
xor U7509 (N_7509,N_7270,N_7231);
nor U7510 (N_7510,N_7344,N_7333);
nor U7511 (N_7511,N_7214,N_7385);
xor U7512 (N_7512,N_7234,N_7266);
or U7513 (N_7513,N_7341,N_7234);
nand U7514 (N_7514,N_7250,N_7273);
or U7515 (N_7515,N_7318,N_7366);
or U7516 (N_7516,N_7389,N_7392);
and U7517 (N_7517,N_7282,N_7379);
xor U7518 (N_7518,N_7385,N_7334);
nor U7519 (N_7519,N_7295,N_7210);
nor U7520 (N_7520,N_7236,N_7271);
nand U7521 (N_7521,N_7210,N_7288);
and U7522 (N_7522,N_7264,N_7238);
and U7523 (N_7523,N_7219,N_7264);
nor U7524 (N_7524,N_7234,N_7287);
and U7525 (N_7525,N_7277,N_7222);
or U7526 (N_7526,N_7225,N_7238);
and U7527 (N_7527,N_7392,N_7230);
nor U7528 (N_7528,N_7394,N_7242);
xor U7529 (N_7529,N_7203,N_7320);
xor U7530 (N_7530,N_7284,N_7392);
and U7531 (N_7531,N_7205,N_7340);
and U7532 (N_7532,N_7263,N_7275);
or U7533 (N_7533,N_7263,N_7217);
xor U7534 (N_7534,N_7290,N_7390);
nor U7535 (N_7535,N_7286,N_7279);
or U7536 (N_7536,N_7229,N_7272);
xor U7537 (N_7537,N_7307,N_7248);
and U7538 (N_7538,N_7270,N_7303);
nand U7539 (N_7539,N_7340,N_7386);
and U7540 (N_7540,N_7389,N_7299);
or U7541 (N_7541,N_7296,N_7278);
xor U7542 (N_7542,N_7345,N_7344);
nor U7543 (N_7543,N_7387,N_7326);
nand U7544 (N_7544,N_7311,N_7249);
nor U7545 (N_7545,N_7233,N_7260);
xor U7546 (N_7546,N_7208,N_7229);
nand U7547 (N_7547,N_7279,N_7343);
xor U7548 (N_7548,N_7337,N_7293);
nor U7549 (N_7549,N_7244,N_7301);
or U7550 (N_7550,N_7211,N_7262);
or U7551 (N_7551,N_7312,N_7318);
nand U7552 (N_7552,N_7385,N_7285);
and U7553 (N_7553,N_7339,N_7372);
nand U7554 (N_7554,N_7372,N_7329);
nand U7555 (N_7555,N_7249,N_7381);
or U7556 (N_7556,N_7328,N_7382);
and U7557 (N_7557,N_7262,N_7296);
and U7558 (N_7558,N_7296,N_7268);
nor U7559 (N_7559,N_7315,N_7388);
and U7560 (N_7560,N_7306,N_7345);
xor U7561 (N_7561,N_7375,N_7348);
xnor U7562 (N_7562,N_7301,N_7395);
nor U7563 (N_7563,N_7200,N_7275);
nand U7564 (N_7564,N_7385,N_7329);
nand U7565 (N_7565,N_7224,N_7205);
xor U7566 (N_7566,N_7280,N_7395);
nor U7567 (N_7567,N_7342,N_7314);
nand U7568 (N_7568,N_7313,N_7246);
xnor U7569 (N_7569,N_7230,N_7352);
or U7570 (N_7570,N_7287,N_7259);
nand U7571 (N_7571,N_7245,N_7307);
xor U7572 (N_7572,N_7255,N_7335);
xnor U7573 (N_7573,N_7377,N_7378);
and U7574 (N_7574,N_7289,N_7335);
nor U7575 (N_7575,N_7324,N_7280);
nand U7576 (N_7576,N_7297,N_7371);
xor U7577 (N_7577,N_7235,N_7217);
and U7578 (N_7578,N_7361,N_7237);
nor U7579 (N_7579,N_7231,N_7263);
nor U7580 (N_7580,N_7312,N_7379);
nand U7581 (N_7581,N_7292,N_7240);
or U7582 (N_7582,N_7268,N_7287);
and U7583 (N_7583,N_7283,N_7389);
and U7584 (N_7584,N_7239,N_7220);
nor U7585 (N_7585,N_7208,N_7334);
and U7586 (N_7586,N_7244,N_7228);
nand U7587 (N_7587,N_7284,N_7249);
nor U7588 (N_7588,N_7291,N_7387);
and U7589 (N_7589,N_7250,N_7211);
nand U7590 (N_7590,N_7208,N_7372);
nand U7591 (N_7591,N_7285,N_7241);
nand U7592 (N_7592,N_7376,N_7230);
xnor U7593 (N_7593,N_7235,N_7325);
xnor U7594 (N_7594,N_7235,N_7336);
and U7595 (N_7595,N_7205,N_7231);
and U7596 (N_7596,N_7281,N_7371);
or U7597 (N_7597,N_7392,N_7220);
nor U7598 (N_7598,N_7345,N_7205);
and U7599 (N_7599,N_7378,N_7293);
xor U7600 (N_7600,N_7404,N_7550);
and U7601 (N_7601,N_7400,N_7434);
nor U7602 (N_7602,N_7411,N_7437);
nand U7603 (N_7603,N_7467,N_7545);
and U7604 (N_7604,N_7509,N_7512);
and U7605 (N_7605,N_7523,N_7458);
nand U7606 (N_7606,N_7419,N_7535);
and U7607 (N_7607,N_7551,N_7573);
nand U7608 (N_7608,N_7567,N_7455);
or U7609 (N_7609,N_7457,N_7585);
nor U7610 (N_7610,N_7529,N_7541);
xnor U7611 (N_7611,N_7469,N_7557);
or U7612 (N_7612,N_7408,N_7471);
nand U7613 (N_7613,N_7402,N_7576);
xnor U7614 (N_7614,N_7525,N_7559);
xnor U7615 (N_7615,N_7561,N_7492);
xor U7616 (N_7616,N_7426,N_7596);
or U7617 (N_7617,N_7444,N_7599);
xor U7618 (N_7618,N_7439,N_7597);
and U7619 (N_7619,N_7405,N_7425);
nor U7620 (N_7620,N_7486,N_7579);
nand U7621 (N_7621,N_7555,N_7450);
and U7622 (N_7622,N_7554,N_7429);
nor U7623 (N_7623,N_7410,N_7563);
or U7624 (N_7624,N_7590,N_7462);
xnor U7625 (N_7625,N_7575,N_7537);
and U7626 (N_7626,N_7443,N_7564);
or U7627 (N_7627,N_7552,N_7514);
nand U7628 (N_7628,N_7591,N_7530);
xor U7629 (N_7629,N_7453,N_7413);
or U7630 (N_7630,N_7586,N_7490);
nand U7631 (N_7631,N_7570,N_7473);
and U7632 (N_7632,N_7440,N_7528);
or U7633 (N_7633,N_7562,N_7474);
xor U7634 (N_7634,N_7589,N_7422);
and U7635 (N_7635,N_7519,N_7436);
nand U7636 (N_7636,N_7583,N_7578);
and U7637 (N_7637,N_7531,N_7544);
or U7638 (N_7638,N_7438,N_7584);
nor U7639 (N_7639,N_7558,N_7403);
xnor U7640 (N_7640,N_7595,N_7442);
xnor U7641 (N_7641,N_7475,N_7420);
nand U7642 (N_7642,N_7417,N_7421);
nor U7643 (N_7643,N_7432,N_7495);
xnor U7644 (N_7644,N_7581,N_7577);
xor U7645 (N_7645,N_7553,N_7415);
nor U7646 (N_7646,N_7502,N_7556);
nor U7647 (N_7647,N_7424,N_7435);
nand U7648 (N_7648,N_7503,N_7480);
xor U7649 (N_7649,N_7482,N_7401);
nor U7650 (N_7650,N_7454,N_7533);
or U7651 (N_7651,N_7511,N_7430);
nand U7652 (N_7652,N_7580,N_7526);
nor U7653 (N_7653,N_7542,N_7449);
nor U7654 (N_7654,N_7518,N_7461);
nor U7655 (N_7655,N_7441,N_7446);
nand U7656 (N_7656,N_7572,N_7451);
and U7657 (N_7657,N_7431,N_7464);
nor U7658 (N_7658,N_7409,N_7406);
and U7659 (N_7659,N_7499,N_7536);
nand U7660 (N_7660,N_7520,N_7510);
xnor U7661 (N_7661,N_7460,N_7485);
and U7662 (N_7662,N_7543,N_7539);
nand U7663 (N_7663,N_7497,N_7515);
nand U7664 (N_7664,N_7513,N_7414);
and U7665 (N_7665,N_7587,N_7517);
nand U7666 (N_7666,N_7433,N_7465);
nor U7667 (N_7667,N_7546,N_7560);
xor U7668 (N_7668,N_7516,N_7494);
or U7669 (N_7669,N_7427,N_7484);
nor U7670 (N_7670,N_7538,N_7508);
xnor U7671 (N_7671,N_7524,N_7452);
nand U7672 (N_7672,N_7483,N_7598);
xnor U7673 (N_7673,N_7593,N_7588);
and U7674 (N_7674,N_7493,N_7506);
and U7675 (N_7675,N_7447,N_7428);
nor U7676 (N_7676,N_7501,N_7488);
or U7677 (N_7677,N_7489,N_7448);
nor U7678 (N_7678,N_7416,N_7534);
nor U7679 (N_7679,N_7477,N_7412);
xor U7680 (N_7680,N_7568,N_7500);
and U7681 (N_7681,N_7527,N_7547);
nor U7682 (N_7682,N_7481,N_7466);
and U7683 (N_7683,N_7594,N_7549);
nor U7684 (N_7684,N_7476,N_7574);
and U7685 (N_7685,N_7496,N_7522);
xor U7686 (N_7686,N_7540,N_7487);
and U7687 (N_7687,N_7423,N_7472);
xnor U7688 (N_7688,N_7569,N_7505);
or U7689 (N_7689,N_7504,N_7521);
or U7690 (N_7690,N_7592,N_7582);
nor U7691 (N_7691,N_7445,N_7459);
nand U7692 (N_7692,N_7566,N_7407);
xnor U7693 (N_7693,N_7478,N_7468);
nor U7694 (N_7694,N_7507,N_7463);
or U7695 (N_7695,N_7456,N_7470);
and U7696 (N_7696,N_7532,N_7571);
or U7697 (N_7697,N_7565,N_7418);
or U7698 (N_7698,N_7491,N_7498);
xor U7699 (N_7699,N_7548,N_7479);
nor U7700 (N_7700,N_7560,N_7402);
nand U7701 (N_7701,N_7579,N_7576);
nor U7702 (N_7702,N_7599,N_7471);
xnor U7703 (N_7703,N_7525,N_7566);
xor U7704 (N_7704,N_7425,N_7539);
nand U7705 (N_7705,N_7569,N_7585);
nor U7706 (N_7706,N_7559,N_7541);
xor U7707 (N_7707,N_7449,N_7409);
or U7708 (N_7708,N_7413,N_7548);
nand U7709 (N_7709,N_7527,N_7421);
and U7710 (N_7710,N_7508,N_7422);
xor U7711 (N_7711,N_7416,N_7554);
xor U7712 (N_7712,N_7447,N_7534);
xnor U7713 (N_7713,N_7419,N_7420);
nor U7714 (N_7714,N_7545,N_7537);
nand U7715 (N_7715,N_7556,N_7535);
nand U7716 (N_7716,N_7557,N_7494);
and U7717 (N_7717,N_7582,N_7572);
or U7718 (N_7718,N_7590,N_7436);
and U7719 (N_7719,N_7487,N_7584);
or U7720 (N_7720,N_7423,N_7476);
xor U7721 (N_7721,N_7454,N_7450);
nand U7722 (N_7722,N_7550,N_7571);
nand U7723 (N_7723,N_7512,N_7490);
or U7724 (N_7724,N_7510,N_7508);
xor U7725 (N_7725,N_7435,N_7511);
or U7726 (N_7726,N_7445,N_7442);
or U7727 (N_7727,N_7460,N_7459);
nor U7728 (N_7728,N_7566,N_7484);
nand U7729 (N_7729,N_7577,N_7487);
and U7730 (N_7730,N_7471,N_7521);
xor U7731 (N_7731,N_7447,N_7569);
and U7732 (N_7732,N_7563,N_7504);
nand U7733 (N_7733,N_7506,N_7557);
nor U7734 (N_7734,N_7413,N_7584);
or U7735 (N_7735,N_7446,N_7589);
nand U7736 (N_7736,N_7594,N_7401);
and U7737 (N_7737,N_7494,N_7520);
nand U7738 (N_7738,N_7469,N_7470);
xor U7739 (N_7739,N_7507,N_7410);
and U7740 (N_7740,N_7524,N_7576);
and U7741 (N_7741,N_7541,N_7494);
xnor U7742 (N_7742,N_7565,N_7402);
or U7743 (N_7743,N_7560,N_7527);
and U7744 (N_7744,N_7445,N_7465);
or U7745 (N_7745,N_7423,N_7561);
and U7746 (N_7746,N_7439,N_7594);
nor U7747 (N_7747,N_7525,N_7575);
xnor U7748 (N_7748,N_7460,N_7476);
xnor U7749 (N_7749,N_7471,N_7440);
or U7750 (N_7750,N_7578,N_7465);
nor U7751 (N_7751,N_7407,N_7466);
nor U7752 (N_7752,N_7563,N_7485);
or U7753 (N_7753,N_7478,N_7421);
xnor U7754 (N_7754,N_7461,N_7439);
nor U7755 (N_7755,N_7419,N_7537);
and U7756 (N_7756,N_7559,N_7512);
or U7757 (N_7757,N_7475,N_7405);
or U7758 (N_7758,N_7439,N_7414);
nand U7759 (N_7759,N_7484,N_7500);
and U7760 (N_7760,N_7444,N_7536);
or U7761 (N_7761,N_7472,N_7507);
xnor U7762 (N_7762,N_7454,N_7461);
or U7763 (N_7763,N_7499,N_7480);
and U7764 (N_7764,N_7487,N_7436);
nor U7765 (N_7765,N_7531,N_7459);
or U7766 (N_7766,N_7509,N_7412);
or U7767 (N_7767,N_7464,N_7548);
xor U7768 (N_7768,N_7583,N_7567);
or U7769 (N_7769,N_7569,N_7504);
xor U7770 (N_7770,N_7513,N_7534);
nand U7771 (N_7771,N_7422,N_7492);
nand U7772 (N_7772,N_7500,N_7517);
or U7773 (N_7773,N_7464,N_7561);
nand U7774 (N_7774,N_7532,N_7466);
nor U7775 (N_7775,N_7422,N_7496);
nor U7776 (N_7776,N_7466,N_7458);
nor U7777 (N_7777,N_7546,N_7500);
and U7778 (N_7778,N_7500,N_7525);
xor U7779 (N_7779,N_7570,N_7407);
xor U7780 (N_7780,N_7484,N_7429);
and U7781 (N_7781,N_7576,N_7514);
nor U7782 (N_7782,N_7566,N_7557);
nor U7783 (N_7783,N_7517,N_7430);
or U7784 (N_7784,N_7535,N_7433);
and U7785 (N_7785,N_7493,N_7498);
nor U7786 (N_7786,N_7577,N_7403);
nand U7787 (N_7787,N_7576,N_7551);
xnor U7788 (N_7788,N_7436,N_7503);
or U7789 (N_7789,N_7511,N_7432);
nand U7790 (N_7790,N_7491,N_7520);
and U7791 (N_7791,N_7500,N_7491);
nand U7792 (N_7792,N_7571,N_7507);
or U7793 (N_7793,N_7450,N_7413);
and U7794 (N_7794,N_7598,N_7478);
and U7795 (N_7795,N_7483,N_7577);
nor U7796 (N_7796,N_7463,N_7488);
or U7797 (N_7797,N_7430,N_7539);
nor U7798 (N_7798,N_7514,N_7471);
xnor U7799 (N_7799,N_7551,N_7554);
nor U7800 (N_7800,N_7703,N_7698);
and U7801 (N_7801,N_7784,N_7690);
nand U7802 (N_7802,N_7630,N_7717);
nand U7803 (N_7803,N_7712,N_7661);
nand U7804 (N_7804,N_7707,N_7695);
nor U7805 (N_7805,N_7607,N_7723);
nor U7806 (N_7806,N_7665,N_7747);
or U7807 (N_7807,N_7671,N_7693);
xor U7808 (N_7808,N_7645,N_7746);
xor U7809 (N_7809,N_7676,N_7666);
nand U7810 (N_7810,N_7683,N_7663);
and U7811 (N_7811,N_7726,N_7793);
nand U7812 (N_7812,N_7625,N_7692);
nand U7813 (N_7813,N_7706,N_7759);
xor U7814 (N_7814,N_7684,N_7766);
nand U7815 (N_7815,N_7659,N_7700);
and U7816 (N_7816,N_7787,N_7752);
nor U7817 (N_7817,N_7791,N_7798);
or U7818 (N_7818,N_7624,N_7732);
xnor U7819 (N_7819,N_7674,N_7620);
and U7820 (N_7820,N_7739,N_7643);
nand U7821 (N_7821,N_7760,N_7646);
xnor U7822 (N_7822,N_7652,N_7672);
nand U7823 (N_7823,N_7713,N_7682);
and U7824 (N_7824,N_7776,N_7770);
nand U7825 (N_7825,N_7675,N_7755);
nand U7826 (N_7826,N_7678,N_7715);
nor U7827 (N_7827,N_7761,N_7753);
and U7828 (N_7828,N_7641,N_7681);
or U7829 (N_7829,N_7777,N_7694);
nand U7830 (N_7830,N_7704,N_7763);
xnor U7831 (N_7831,N_7685,N_7741);
xnor U7832 (N_7832,N_7740,N_7656);
nand U7833 (N_7833,N_7702,N_7628);
or U7834 (N_7834,N_7658,N_7719);
or U7835 (N_7835,N_7795,N_7792);
and U7836 (N_7836,N_7609,N_7637);
or U7837 (N_7837,N_7765,N_7764);
xor U7838 (N_7838,N_7610,N_7638);
or U7839 (N_7839,N_7626,N_7697);
nor U7840 (N_7840,N_7714,N_7633);
and U7841 (N_7841,N_7779,N_7686);
nor U7842 (N_7842,N_7757,N_7789);
and U7843 (N_7843,N_7794,N_7745);
nor U7844 (N_7844,N_7754,N_7606);
or U7845 (N_7845,N_7735,N_7632);
nor U7846 (N_7846,N_7605,N_7631);
xnor U7847 (N_7847,N_7736,N_7680);
nand U7848 (N_7848,N_7668,N_7748);
xnor U7849 (N_7849,N_7785,N_7710);
xnor U7850 (N_7850,N_7774,N_7679);
and U7851 (N_7851,N_7691,N_7662);
nor U7852 (N_7852,N_7602,N_7769);
and U7853 (N_7853,N_7660,N_7771);
or U7854 (N_7854,N_7640,N_7603);
nand U7855 (N_7855,N_7720,N_7782);
xor U7856 (N_7856,N_7687,N_7749);
nor U7857 (N_7857,N_7751,N_7613);
and U7858 (N_7858,N_7727,N_7621);
nor U7859 (N_7859,N_7619,N_7618);
and U7860 (N_7860,N_7716,N_7701);
and U7861 (N_7861,N_7742,N_7756);
nand U7862 (N_7862,N_7731,N_7758);
nor U7863 (N_7863,N_7750,N_7614);
nand U7864 (N_7864,N_7655,N_7711);
xor U7865 (N_7865,N_7616,N_7601);
nor U7866 (N_7866,N_7600,N_7725);
or U7867 (N_7867,N_7636,N_7728);
xnor U7868 (N_7868,N_7688,N_7737);
xnor U7869 (N_7869,N_7705,N_7762);
nand U7870 (N_7870,N_7604,N_7615);
and U7871 (N_7871,N_7608,N_7790);
and U7872 (N_7872,N_7670,N_7778);
nor U7873 (N_7873,N_7664,N_7730);
nor U7874 (N_7874,N_7654,N_7611);
nand U7875 (N_7875,N_7623,N_7648);
nand U7876 (N_7876,N_7721,N_7651);
and U7877 (N_7877,N_7667,N_7797);
or U7878 (N_7878,N_7709,N_7634);
xor U7879 (N_7879,N_7699,N_7649);
xnor U7880 (N_7880,N_7781,N_7647);
or U7881 (N_7881,N_7629,N_7627);
xnor U7882 (N_7882,N_7733,N_7642);
and U7883 (N_7883,N_7743,N_7796);
and U7884 (N_7884,N_7775,N_7689);
and U7885 (N_7885,N_7768,N_7780);
xnor U7886 (N_7886,N_7799,N_7729);
or U7887 (N_7887,N_7788,N_7696);
xnor U7888 (N_7888,N_7744,N_7650);
or U7889 (N_7889,N_7644,N_7639);
and U7890 (N_7890,N_7786,N_7722);
nor U7891 (N_7891,N_7738,N_7708);
and U7892 (N_7892,N_7677,N_7772);
or U7893 (N_7893,N_7724,N_7617);
xnor U7894 (N_7894,N_7734,N_7669);
nor U7895 (N_7895,N_7783,N_7657);
or U7896 (N_7896,N_7767,N_7635);
xor U7897 (N_7897,N_7773,N_7718);
or U7898 (N_7898,N_7622,N_7612);
xnor U7899 (N_7899,N_7653,N_7673);
or U7900 (N_7900,N_7785,N_7751);
and U7901 (N_7901,N_7761,N_7771);
xnor U7902 (N_7902,N_7630,N_7785);
xnor U7903 (N_7903,N_7617,N_7610);
nor U7904 (N_7904,N_7608,N_7700);
or U7905 (N_7905,N_7638,N_7645);
and U7906 (N_7906,N_7678,N_7641);
nand U7907 (N_7907,N_7751,N_7624);
or U7908 (N_7908,N_7631,N_7639);
xor U7909 (N_7909,N_7662,N_7652);
nor U7910 (N_7910,N_7622,N_7648);
or U7911 (N_7911,N_7780,N_7632);
nand U7912 (N_7912,N_7765,N_7649);
nor U7913 (N_7913,N_7662,N_7664);
nand U7914 (N_7914,N_7734,N_7606);
nor U7915 (N_7915,N_7607,N_7647);
or U7916 (N_7916,N_7680,N_7741);
nand U7917 (N_7917,N_7658,N_7664);
nand U7918 (N_7918,N_7749,N_7781);
and U7919 (N_7919,N_7600,N_7742);
or U7920 (N_7920,N_7657,N_7654);
and U7921 (N_7921,N_7658,N_7785);
and U7922 (N_7922,N_7764,N_7781);
xor U7923 (N_7923,N_7798,N_7754);
xor U7924 (N_7924,N_7671,N_7667);
and U7925 (N_7925,N_7622,N_7650);
xor U7926 (N_7926,N_7684,N_7739);
nor U7927 (N_7927,N_7721,N_7711);
nand U7928 (N_7928,N_7715,N_7636);
or U7929 (N_7929,N_7785,N_7794);
nor U7930 (N_7930,N_7652,N_7799);
or U7931 (N_7931,N_7716,N_7636);
or U7932 (N_7932,N_7707,N_7688);
and U7933 (N_7933,N_7699,N_7691);
and U7934 (N_7934,N_7796,N_7679);
or U7935 (N_7935,N_7757,N_7763);
or U7936 (N_7936,N_7677,N_7607);
nand U7937 (N_7937,N_7600,N_7781);
or U7938 (N_7938,N_7760,N_7697);
and U7939 (N_7939,N_7716,N_7642);
nand U7940 (N_7940,N_7722,N_7604);
or U7941 (N_7941,N_7788,N_7782);
and U7942 (N_7942,N_7714,N_7739);
nand U7943 (N_7943,N_7703,N_7606);
nand U7944 (N_7944,N_7672,N_7696);
or U7945 (N_7945,N_7702,N_7745);
nor U7946 (N_7946,N_7700,N_7713);
xor U7947 (N_7947,N_7742,N_7750);
xor U7948 (N_7948,N_7655,N_7699);
xnor U7949 (N_7949,N_7784,N_7712);
or U7950 (N_7950,N_7623,N_7713);
and U7951 (N_7951,N_7716,N_7688);
or U7952 (N_7952,N_7755,N_7749);
nor U7953 (N_7953,N_7711,N_7743);
and U7954 (N_7954,N_7673,N_7709);
xnor U7955 (N_7955,N_7623,N_7662);
and U7956 (N_7956,N_7604,N_7608);
and U7957 (N_7957,N_7614,N_7654);
nor U7958 (N_7958,N_7716,N_7682);
nand U7959 (N_7959,N_7772,N_7637);
and U7960 (N_7960,N_7780,N_7721);
or U7961 (N_7961,N_7636,N_7788);
or U7962 (N_7962,N_7670,N_7796);
xnor U7963 (N_7963,N_7659,N_7723);
xnor U7964 (N_7964,N_7647,N_7759);
or U7965 (N_7965,N_7754,N_7659);
and U7966 (N_7966,N_7602,N_7643);
or U7967 (N_7967,N_7636,N_7676);
and U7968 (N_7968,N_7718,N_7792);
nor U7969 (N_7969,N_7797,N_7639);
xor U7970 (N_7970,N_7766,N_7714);
nor U7971 (N_7971,N_7641,N_7698);
nor U7972 (N_7972,N_7636,N_7791);
and U7973 (N_7973,N_7747,N_7670);
and U7974 (N_7974,N_7711,N_7730);
or U7975 (N_7975,N_7798,N_7725);
and U7976 (N_7976,N_7776,N_7720);
xor U7977 (N_7977,N_7759,N_7652);
xnor U7978 (N_7978,N_7643,N_7693);
or U7979 (N_7979,N_7656,N_7752);
and U7980 (N_7980,N_7789,N_7657);
nand U7981 (N_7981,N_7657,N_7610);
nor U7982 (N_7982,N_7625,N_7777);
or U7983 (N_7983,N_7799,N_7764);
nor U7984 (N_7984,N_7685,N_7607);
nor U7985 (N_7985,N_7693,N_7656);
xnor U7986 (N_7986,N_7724,N_7737);
or U7987 (N_7987,N_7664,N_7614);
and U7988 (N_7988,N_7751,N_7611);
xnor U7989 (N_7989,N_7607,N_7697);
xnor U7990 (N_7990,N_7783,N_7729);
nand U7991 (N_7991,N_7737,N_7762);
xor U7992 (N_7992,N_7773,N_7602);
and U7993 (N_7993,N_7750,N_7735);
and U7994 (N_7994,N_7715,N_7781);
xor U7995 (N_7995,N_7796,N_7697);
nor U7996 (N_7996,N_7672,N_7779);
nor U7997 (N_7997,N_7756,N_7711);
nand U7998 (N_7998,N_7633,N_7732);
nor U7999 (N_7999,N_7626,N_7746);
nand U8000 (N_8000,N_7809,N_7870);
nand U8001 (N_8001,N_7894,N_7859);
or U8002 (N_8002,N_7899,N_7818);
xnor U8003 (N_8003,N_7992,N_7967);
xor U8004 (N_8004,N_7991,N_7934);
nor U8005 (N_8005,N_7984,N_7922);
nor U8006 (N_8006,N_7988,N_7808);
or U8007 (N_8007,N_7840,N_7960);
and U8008 (N_8008,N_7883,N_7918);
nor U8009 (N_8009,N_7920,N_7850);
xor U8010 (N_8010,N_7896,N_7907);
nor U8011 (N_8011,N_7949,N_7805);
and U8012 (N_8012,N_7893,N_7832);
xnor U8013 (N_8013,N_7955,N_7904);
nor U8014 (N_8014,N_7905,N_7956);
and U8015 (N_8015,N_7916,N_7810);
or U8016 (N_8016,N_7946,N_7813);
xnor U8017 (N_8017,N_7930,N_7932);
nand U8018 (N_8018,N_7990,N_7892);
nand U8019 (N_8019,N_7948,N_7997);
nand U8020 (N_8020,N_7915,N_7943);
or U8021 (N_8021,N_7817,N_7823);
xor U8022 (N_8022,N_7857,N_7868);
nor U8023 (N_8023,N_7906,N_7901);
nor U8024 (N_8024,N_7933,N_7875);
xnor U8025 (N_8025,N_7909,N_7942);
and U8026 (N_8026,N_7924,N_7878);
xnor U8027 (N_8027,N_7923,N_7839);
and U8028 (N_8028,N_7841,N_7958);
xor U8029 (N_8029,N_7854,N_7830);
nand U8030 (N_8030,N_7864,N_7911);
or U8031 (N_8031,N_7848,N_7996);
xor U8032 (N_8032,N_7941,N_7944);
nor U8033 (N_8033,N_7884,N_7998);
and U8034 (N_8034,N_7816,N_7889);
or U8035 (N_8035,N_7994,N_7903);
nor U8036 (N_8036,N_7925,N_7858);
xor U8037 (N_8037,N_7837,N_7975);
and U8038 (N_8038,N_7908,N_7953);
and U8039 (N_8039,N_7962,N_7807);
and U8040 (N_8040,N_7999,N_7844);
nand U8041 (N_8041,N_7867,N_7940);
nor U8042 (N_8042,N_7983,N_7959);
xnor U8043 (N_8043,N_7872,N_7866);
and U8044 (N_8044,N_7945,N_7853);
or U8045 (N_8045,N_7928,N_7833);
nand U8046 (N_8046,N_7973,N_7989);
xnor U8047 (N_8047,N_7880,N_7855);
nand U8048 (N_8048,N_7842,N_7828);
or U8049 (N_8049,N_7952,N_7968);
nor U8050 (N_8050,N_7897,N_7815);
xnor U8051 (N_8051,N_7985,N_7965);
xor U8052 (N_8052,N_7982,N_7898);
and U8053 (N_8053,N_7882,N_7829);
nand U8054 (N_8054,N_7860,N_7863);
nor U8055 (N_8055,N_7902,N_7927);
and U8056 (N_8056,N_7803,N_7871);
and U8057 (N_8057,N_7865,N_7887);
xor U8058 (N_8058,N_7938,N_7972);
xor U8059 (N_8059,N_7970,N_7976);
or U8060 (N_8060,N_7811,N_7879);
and U8061 (N_8061,N_7847,N_7914);
and U8062 (N_8062,N_7849,N_7993);
xnor U8063 (N_8063,N_7912,N_7822);
and U8064 (N_8064,N_7804,N_7939);
or U8065 (N_8065,N_7888,N_7935);
nand U8066 (N_8066,N_7886,N_7969);
and U8067 (N_8067,N_7845,N_7824);
xnor U8068 (N_8068,N_7913,N_7877);
or U8069 (N_8069,N_7986,N_7974);
nand U8070 (N_8070,N_7814,N_7802);
or U8071 (N_8071,N_7826,N_7820);
xnor U8072 (N_8072,N_7961,N_7836);
xnor U8073 (N_8073,N_7801,N_7862);
or U8074 (N_8074,N_7825,N_7869);
or U8075 (N_8075,N_7917,N_7978);
nand U8076 (N_8076,N_7885,N_7926);
nor U8077 (N_8077,N_7929,N_7947);
xnor U8078 (N_8078,N_7966,N_7838);
nor U8079 (N_8079,N_7891,N_7919);
nor U8080 (N_8080,N_7931,N_7979);
and U8081 (N_8081,N_7800,N_7987);
xor U8082 (N_8082,N_7950,N_7900);
nand U8083 (N_8083,N_7954,N_7895);
nor U8084 (N_8084,N_7921,N_7874);
nor U8085 (N_8085,N_7977,N_7821);
xor U8086 (N_8086,N_7861,N_7806);
and U8087 (N_8087,N_7852,N_7851);
and U8088 (N_8088,N_7981,N_7937);
and U8089 (N_8089,N_7834,N_7843);
nand U8090 (N_8090,N_7881,N_7835);
or U8091 (N_8091,N_7819,N_7980);
and U8092 (N_8092,N_7890,N_7873);
or U8093 (N_8093,N_7963,N_7971);
and U8094 (N_8094,N_7812,N_7910);
xnor U8095 (N_8095,N_7957,N_7995);
xor U8096 (N_8096,N_7951,N_7856);
nand U8097 (N_8097,N_7876,N_7827);
or U8098 (N_8098,N_7831,N_7846);
nand U8099 (N_8099,N_7936,N_7964);
xor U8100 (N_8100,N_7953,N_7812);
nor U8101 (N_8101,N_7883,N_7897);
nor U8102 (N_8102,N_7890,N_7959);
or U8103 (N_8103,N_7927,N_7886);
or U8104 (N_8104,N_7823,N_7839);
or U8105 (N_8105,N_7801,N_7929);
and U8106 (N_8106,N_7870,N_7961);
nand U8107 (N_8107,N_7833,N_7870);
nor U8108 (N_8108,N_7924,N_7949);
nor U8109 (N_8109,N_7941,N_7960);
xnor U8110 (N_8110,N_7935,N_7955);
or U8111 (N_8111,N_7933,N_7910);
xor U8112 (N_8112,N_7963,N_7992);
xor U8113 (N_8113,N_7919,N_7934);
or U8114 (N_8114,N_7850,N_7980);
or U8115 (N_8115,N_7834,N_7833);
and U8116 (N_8116,N_7984,N_7953);
nor U8117 (N_8117,N_7878,N_7867);
or U8118 (N_8118,N_7952,N_7908);
and U8119 (N_8119,N_7849,N_7956);
and U8120 (N_8120,N_7823,N_7853);
and U8121 (N_8121,N_7998,N_7850);
or U8122 (N_8122,N_7925,N_7918);
or U8123 (N_8123,N_7853,N_7880);
nand U8124 (N_8124,N_7885,N_7968);
and U8125 (N_8125,N_7901,N_7831);
nand U8126 (N_8126,N_7900,N_7889);
nor U8127 (N_8127,N_7888,N_7975);
nand U8128 (N_8128,N_7900,N_7957);
or U8129 (N_8129,N_7911,N_7917);
or U8130 (N_8130,N_7980,N_7909);
and U8131 (N_8131,N_7862,N_7891);
and U8132 (N_8132,N_7819,N_7858);
or U8133 (N_8133,N_7865,N_7944);
nand U8134 (N_8134,N_7881,N_7947);
nor U8135 (N_8135,N_7964,N_7999);
or U8136 (N_8136,N_7980,N_7840);
nor U8137 (N_8137,N_7932,N_7829);
and U8138 (N_8138,N_7906,N_7894);
nor U8139 (N_8139,N_7881,N_7885);
nor U8140 (N_8140,N_7856,N_7869);
or U8141 (N_8141,N_7902,N_7892);
and U8142 (N_8142,N_7847,N_7979);
xor U8143 (N_8143,N_7942,N_7874);
or U8144 (N_8144,N_7861,N_7989);
xnor U8145 (N_8145,N_7815,N_7844);
or U8146 (N_8146,N_7999,N_7828);
and U8147 (N_8147,N_7873,N_7888);
or U8148 (N_8148,N_7808,N_7834);
or U8149 (N_8149,N_7851,N_7829);
xnor U8150 (N_8150,N_7857,N_7941);
xnor U8151 (N_8151,N_7980,N_7803);
or U8152 (N_8152,N_7978,N_7909);
nor U8153 (N_8153,N_7975,N_7947);
nand U8154 (N_8154,N_7804,N_7997);
nand U8155 (N_8155,N_7979,N_7882);
nand U8156 (N_8156,N_7953,N_7829);
and U8157 (N_8157,N_7980,N_7861);
nand U8158 (N_8158,N_7973,N_7890);
or U8159 (N_8159,N_7996,N_7891);
xnor U8160 (N_8160,N_7964,N_7900);
or U8161 (N_8161,N_7932,N_7906);
xnor U8162 (N_8162,N_7818,N_7865);
nor U8163 (N_8163,N_7984,N_7949);
xnor U8164 (N_8164,N_7931,N_7821);
nand U8165 (N_8165,N_7815,N_7921);
nor U8166 (N_8166,N_7952,N_7812);
nand U8167 (N_8167,N_7811,N_7878);
nor U8168 (N_8168,N_7902,N_7907);
nand U8169 (N_8169,N_7971,N_7805);
and U8170 (N_8170,N_7898,N_7890);
or U8171 (N_8171,N_7804,N_7982);
nor U8172 (N_8172,N_7919,N_7852);
xnor U8173 (N_8173,N_7905,N_7930);
nand U8174 (N_8174,N_7957,N_7914);
or U8175 (N_8175,N_7885,N_7833);
and U8176 (N_8176,N_7833,N_7904);
nor U8177 (N_8177,N_7925,N_7901);
nor U8178 (N_8178,N_7985,N_7961);
and U8179 (N_8179,N_7941,N_7939);
nand U8180 (N_8180,N_7880,N_7912);
nand U8181 (N_8181,N_7944,N_7979);
xnor U8182 (N_8182,N_7885,N_7855);
or U8183 (N_8183,N_7893,N_7854);
nand U8184 (N_8184,N_7806,N_7871);
nor U8185 (N_8185,N_7900,N_7878);
or U8186 (N_8186,N_7822,N_7863);
xnor U8187 (N_8187,N_7822,N_7862);
and U8188 (N_8188,N_7991,N_7866);
nand U8189 (N_8189,N_7932,N_7806);
and U8190 (N_8190,N_7926,N_7873);
xor U8191 (N_8191,N_7824,N_7922);
nand U8192 (N_8192,N_7978,N_7971);
nor U8193 (N_8193,N_7981,N_7821);
xnor U8194 (N_8194,N_7830,N_7933);
or U8195 (N_8195,N_7863,N_7973);
nor U8196 (N_8196,N_7931,N_7918);
and U8197 (N_8197,N_7855,N_7815);
or U8198 (N_8198,N_7981,N_7851);
nor U8199 (N_8199,N_7929,N_7808);
nand U8200 (N_8200,N_8155,N_8178);
nor U8201 (N_8201,N_8168,N_8045);
nand U8202 (N_8202,N_8030,N_8127);
nand U8203 (N_8203,N_8106,N_8046);
or U8204 (N_8204,N_8174,N_8007);
xnor U8205 (N_8205,N_8105,N_8147);
or U8206 (N_8206,N_8038,N_8133);
xnor U8207 (N_8207,N_8083,N_8080);
and U8208 (N_8208,N_8092,N_8167);
or U8209 (N_8209,N_8116,N_8135);
xnor U8210 (N_8210,N_8042,N_8071);
xnor U8211 (N_8211,N_8000,N_8193);
nor U8212 (N_8212,N_8180,N_8094);
and U8213 (N_8213,N_8126,N_8025);
and U8214 (N_8214,N_8197,N_8048);
and U8215 (N_8215,N_8113,N_8063);
nor U8216 (N_8216,N_8043,N_8142);
xnor U8217 (N_8217,N_8010,N_8132);
and U8218 (N_8218,N_8187,N_8122);
xor U8219 (N_8219,N_8076,N_8152);
xnor U8220 (N_8220,N_8091,N_8172);
nor U8221 (N_8221,N_8103,N_8017);
or U8222 (N_8222,N_8096,N_8179);
nor U8223 (N_8223,N_8067,N_8065);
and U8224 (N_8224,N_8002,N_8018);
and U8225 (N_8225,N_8108,N_8049);
or U8226 (N_8226,N_8196,N_8124);
nand U8227 (N_8227,N_8123,N_8084);
nand U8228 (N_8228,N_8198,N_8166);
and U8229 (N_8229,N_8078,N_8064);
xnor U8230 (N_8230,N_8139,N_8060);
or U8231 (N_8231,N_8044,N_8016);
or U8232 (N_8232,N_8057,N_8115);
or U8233 (N_8233,N_8006,N_8011);
and U8234 (N_8234,N_8136,N_8144);
nor U8235 (N_8235,N_8099,N_8023);
nor U8236 (N_8236,N_8058,N_8192);
nor U8237 (N_8237,N_8062,N_8009);
nand U8238 (N_8238,N_8028,N_8075);
xor U8239 (N_8239,N_8027,N_8114);
xor U8240 (N_8240,N_8151,N_8101);
nor U8241 (N_8241,N_8169,N_8015);
nor U8242 (N_8242,N_8053,N_8183);
nor U8243 (N_8243,N_8047,N_8087);
and U8244 (N_8244,N_8081,N_8153);
nor U8245 (N_8245,N_8146,N_8110);
nor U8246 (N_8246,N_8148,N_8039);
or U8247 (N_8247,N_8014,N_8150);
or U8248 (N_8248,N_8111,N_8095);
nand U8249 (N_8249,N_8066,N_8164);
nand U8250 (N_8250,N_8182,N_8041);
and U8251 (N_8251,N_8161,N_8194);
nand U8252 (N_8252,N_8077,N_8074);
and U8253 (N_8253,N_8033,N_8154);
and U8254 (N_8254,N_8118,N_8158);
nand U8255 (N_8255,N_8032,N_8119);
or U8256 (N_8256,N_8162,N_8188);
xnor U8257 (N_8257,N_8001,N_8021);
and U8258 (N_8258,N_8037,N_8059);
xnor U8259 (N_8259,N_8013,N_8121);
or U8260 (N_8260,N_8003,N_8022);
xor U8261 (N_8261,N_8165,N_8035);
and U8262 (N_8262,N_8031,N_8051);
and U8263 (N_8263,N_8020,N_8145);
nand U8264 (N_8264,N_8120,N_8156);
nor U8265 (N_8265,N_8159,N_8189);
nand U8266 (N_8266,N_8079,N_8068);
nand U8267 (N_8267,N_8034,N_8185);
nor U8268 (N_8268,N_8131,N_8029);
or U8269 (N_8269,N_8190,N_8052);
nor U8270 (N_8270,N_8026,N_8024);
and U8271 (N_8271,N_8112,N_8008);
and U8272 (N_8272,N_8130,N_8171);
xor U8273 (N_8273,N_8098,N_8186);
xor U8274 (N_8274,N_8125,N_8019);
nor U8275 (N_8275,N_8070,N_8129);
and U8276 (N_8276,N_8086,N_8177);
or U8277 (N_8277,N_8104,N_8137);
and U8278 (N_8278,N_8072,N_8093);
or U8279 (N_8279,N_8004,N_8140);
nand U8280 (N_8280,N_8055,N_8175);
and U8281 (N_8281,N_8173,N_8088);
nand U8282 (N_8282,N_8097,N_8138);
or U8283 (N_8283,N_8181,N_8056);
nand U8284 (N_8284,N_8050,N_8100);
xnor U8285 (N_8285,N_8170,N_8134);
xor U8286 (N_8286,N_8061,N_8117);
and U8287 (N_8287,N_8085,N_8143);
or U8288 (N_8288,N_8082,N_8107);
nor U8289 (N_8289,N_8191,N_8005);
nand U8290 (N_8290,N_8195,N_8160);
and U8291 (N_8291,N_8141,N_8102);
nand U8292 (N_8292,N_8073,N_8149);
or U8293 (N_8293,N_8157,N_8012);
nor U8294 (N_8294,N_8199,N_8036);
xor U8295 (N_8295,N_8128,N_8040);
nor U8296 (N_8296,N_8054,N_8069);
or U8297 (N_8297,N_8109,N_8163);
nand U8298 (N_8298,N_8090,N_8089);
or U8299 (N_8299,N_8184,N_8176);
nand U8300 (N_8300,N_8197,N_8070);
nor U8301 (N_8301,N_8099,N_8056);
xnor U8302 (N_8302,N_8006,N_8199);
or U8303 (N_8303,N_8020,N_8182);
nand U8304 (N_8304,N_8113,N_8038);
and U8305 (N_8305,N_8150,N_8103);
nand U8306 (N_8306,N_8133,N_8175);
xnor U8307 (N_8307,N_8103,N_8128);
or U8308 (N_8308,N_8071,N_8151);
or U8309 (N_8309,N_8023,N_8186);
or U8310 (N_8310,N_8110,N_8068);
nand U8311 (N_8311,N_8114,N_8142);
nor U8312 (N_8312,N_8034,N_8188);
xnor U8313 (N_8313,N_8140,N_8181);
nand U8314 (N_8314,N_8117,N_8151);
xor U8315 (N_8315,N_8014,N_8082);
xor U8316 (N_8316,N_8106,N_8148);
or U8317 (N_8317,N_8096,N_8156);
nor U8318 (N_8318,N_8035,N_8025);
nor U8319 (N_8319,N_8136,N_8156);
xor U8320 (N_8320,N_8009,N_8087);
and U8321 (N_8321,N_8153,N_8063);
nor U8322 (N_8322,N_8106,N_8071);
nand U8323 (N_8323,N_8128,N_8011);
nand U8324 (N_8324,N_8161,N_8170);
nor U8325 (N_8325,N_8024,N_8143);
or U8326 (N_8326,N_8006,N_8182);
nor U8327 (N_8327,N_8136,N_8078);
or U8328 (N_8328,N_8066,N_8005);
nor U8329 (N_8329,N_8101,N_8131);
nor U8330 (N_8330,N_8015,N_8180);
nand U8331 (N_8331,N_8109,N_8098);
and U8332 (N_8332,N_8110,N_8162);
nor U8333 (N_8333,N_8085,N_8081);
and U8334 (N_8334,N_8186,N_8188);
and U8335 (N_8335,N_8148,N_8085);
nand U8336 (N_8336,N_8149,N_8057);
nor U8337 (N_8337,N_8151,N_8177);
nand U8338 (N_8338,N_8181,N_8139);
nand U8339 (N_8339,N_8048,N_8062);
xor U8340 (N_8340,N_8093,N_8149);
nand U8341 (N_8341,N_8157,N_8079);
nor U8342 (N_8342,N_8181,N_8183);
or U8343 (N_8343,N_8102,N_8043);
xor U8344 (N_8344,N_8181,N_8076);
nor U8345 (N_8345,N_8175,N_8110);
nor U8346 (N_8346,N_8198,N_8133);
xor U8347 (N_8347,N_8101,N_8146);
and U8348 (N_8348,N_8010,N_8149);
nand U8349 (N_8349,N_8015,N_8189);
or U8350 (N_8350,N_8080,N_8062);
nand U8351 (N_8351,N_8001,N_8119);
and U8352 (N_8352,N_8081,N_8064);
nand U8353 (N_8353,N_8049,N_8059);
and U8354 (N_8354,N_8036,N_8119);
xor U8355 (N_8355,N_8166,N_8169);
nor U8356 (N_8356,N_8196,N_8025);
nand U8357 (N_8357,N_8082,N_8144);
nand U8358 (N_8358,N_8198,N_8091);
xnor U8359 (N_8359,N_8100,N_8067);
and U8360 (N_8360,N_8096,N_8141);
or U8361 (N_8361,N_8143,N_8075);
or U8362 (N_8362,N_8185,N_8070);
nor U8363 (N_8363,N_8020,N_8076);
and U8364 (N_8364,N_8031,N_8185);
xor U8365 (N_8365,N_8123,N_8100);
or U8366 (N_8366,N_8059,N_8110);
and U8367 (N_8367,N_8185,N_8180);
xor U8368 (N_8368,N_8005,N_8121);
and U8369 (N_8369,N_8057,N_8163);
and U8370 (N_8370,N_8082,N_8137);
or U8371 (N_8371,N_8070,N_8058);
nor U8372 (N_8372,N_8191,N_8092);
xnor U8373 (N_8373,N_8163,N_8133);
nand U8374 (N_8374,N_8030,N_8181);
and U8375 (N_8375,N_8158,N_8126);
xnor U8376 (N_8376,N_8117,N_8149);
or U8377 (N_8377,N_8061,N_8185);
or U8378 (N_8378,N_8059,N_8022);
xor U8379 (N_8379,N_8058,N_8117);
xor U8380 (N_8380,N_8118,N_8018);
xor U8381 (N_8381,N_8165,N_8191);
and U8382 (N_8382,N_8104,N_8023);
nor U8383 (N_8383,N_8170,N_8073);
nand U8384 (N_8384,N_8071,N_8018);
or U8385 (N_8385,N_8182,N_8016);
nand U8386 (N_8386,N_8137,N_8018);
or U8387 (N_8387,N_8147,N_8120);
nor U8388 (N_8388,N_8159,N_8101);
nand U8389 (N_8389,N_8010,N_8140);
or U8390 (N_8390,N_8124,N_8182);
nor U8391 (N_8391,N_8025,N_8071);
xor U8392 (N_8392,N_8152,N_8065);
or U8393 (N_8393,N_8170,N_8097);
xnor U8394 (N_8394,N_8105,N_8057);
or U8395 (N_8395,N_8037,N_8139);
xor U8396 (N_8396,N_8184,N_8052);
nor U8397 (N_8397,N_8171,N_8107);
nor U8398 (N_8398,N_8084,N_8034);
nand U8399 (N_8399,N_8151,N_8083);
nand U8400 (N_8400,N_8360,N_8333);
xnor U8401 (N_8401,N_8350,N_8292);
and U8402 (N_8402,N_8338,N_8309);
nor U8403 (N_8403,N_8246,N_8210);
and U8404 (N_8404,N_8348,N_8240);
nor U8405 (N_8405,N_8353,N_8253);
nand U8406 (N_8406,N_8375,N_8344);
and U8407 (N_8407,N_8256,N_8318);
xnor U8408 (N_8408,N_8346,N_8284);
nand U8409 (N_8409,N_8233,N_8285);
and U8410 (N_8410,N_8308,N_8366);
xor U8411 (N_8411,N_8362,N_8295);
or U8412 (N_8412,N_8257,N_8393);
nand U8413 (N_8413,N_8316,N_8201);
or U8414 (N_8414,N_8207,N_8358);
and U8415 (N_8415,N_8381,N_8231);
or U8416 (N_8416,N_8315,N_8245);
and U8417 (N_8417,N_8216,N_8235);
and U8418 (N_8418,N_8218,N_8352);
and U8419 (N_8419,N_8277,N_8282);
and U8420 (N_8420,N_8329,N_8349);
nor U8421 (N_8421,N_8335,N_8331);
nand U8422 (N_8422,N_8242,N_8205);
xor U8423 (N_8423,N_8301,N_8307);
xnor U8424 (N_8424,N_8286,N_8363);
and U8425 (N_8425,N_8357,N_8265);
nand U8426 (N_8426,N_8370,N_8220);
or U8427 (N_8427,N_8356,N_8280);
and U8428 (N_8428,N_8336,N_8248);
or U8429 (N_8429,N_8342,N_8320);
and U8430 (N_8430,N_8274,N_8391);
xnor U8431 (N_8431,N_8281,N_8247);
nand U8432 (N_8432,N_8399,N_8398);
and U8433 (N_8433,N_8310,N_8317);
nand U8434 (N_8434,N_8289,N_8283);
or U8435 (N_8435,N_8387,N_8323);
and U8436 (N_8436,N_8373,N_8211);
and U8437 (N_8437,N_8337,N_8326);
nor U8438 (N_8438,N_8380,N_8293);
xor U8439 (N_8439,N_8252,N_8374);
nand U8440 (N_8440,N_8340,N_8367);
nand U8441 (N_8441,N_8251,N_8325);
xor U8442 (N_8442,N_8260,N_8266);
nand U8443 (N_8443,N_8296,N_8297);
and U8444 (N_8444,N_8278,N_8330);
or U8445 (N_8445,N_8345,N_8239);
nor U8446 (N_8446,N_8385,N_8376);
and U8447 (N_8447,N_8262,N_8324);
and U8448 (N_8448,N_8384,N_8206);
nand U8449 (N_8449,N_8254,N_8208);
nor U8450 (N_8450,N_8304,N_8229);
or U8451 (N_8451,N_8300,N_8202);
and U8452 (N_8452,N_8227,N_8294);
nand U8453 (N_8453,N_8312,N_8270);
or U8454 (N_8454,N_8321,N_8314);
xor U8455 (N_8455,N_8249,N_8311);
or U8456 (N_8456,N_8224,N_8361);
nand U8457 (N_8457,N_8302,N_8390);
nand U8458 (N_8458,N_8226,N_8327);
or U8459 (N_8459,N_8332,N_8223);
or U8460 (N_8460,N_8339,N_8264);
or U8461 (N_8461,N_8386,N_8371);
and U8462 (N_8462,N_8359,N_8268);
xor U8463 (N_8463,N_8319,N_8213);
nand U8464 (N_8464,N_8236,N_8379);
nor U8465 (N_8465,N_8214,N_8272);
xor U8466 (N_8466,N_8306,N_8238);
and U8467 (N_8467,N_8396,N_8389);
nor U8468 (N_8468,N_8343,N_8347);
or U8469 (N_8469,N_8368,N_8313);
or U8470 (N_8470,N_8275,N_8328);
nand U8471 (N_8471,N_8341,N_8276);
nand U8472 (N_8472,N_8291,N_8212);
nor U8473 (N_8473,N_8382,N_8222);
nand U8474 (N_8474,N_8243,N_8237);
nand U8475 (N_8475,N_8261,N_8241);
nand U8476 (N_8476,N_8299,N_8217);
and U8477 (N_8477,N_8225,N_8397);
nor U8478 (N_8478,N_8234,N_8395);
and U8479 (N_8479,N_8372,N_8228);
nand U8480 (N_8480,N_8271,N_8200);
xnor U8481 (N_8481,N_8322,N_8269);
or U8482 (N_8482,N_8219,N_8221);
nand U8483 (N_8483,N_8365,N_8394);
nand U8484 (N_8484,N_8369,N_8378);
or U8485 (N_8485,N_8303,N_8377);
nor U8486 (N_8486,N_8273,N_8258);
xor U8487 (N_8487,N_8244,N_8334);
or U8488 (N_8488,N_8351,N_8298);
xnor U8489 (N_8489,N_8232,N_8263);
xor U8490 (N_8490,N_8383,N_8290);
and U8491 (N_8491,N_8255,N_8230);
xnor U8492 (N_8492,N_8364,N_8215);
and U8493 (N_8493,N_8388,N_8259);
and U8494 (N_8494,N_8204,N_8288);
nor U8495 (N_8495,N_8203,N_8279);
nor U8496 (N_8496,N_8250,N_8392);
xor U8497 (N_8497,N_8354,N_8267);
and U8498 (N_8498,N_8209,N_8287);
nand U8499 (N_8499,N_8355,N_8305);
nand U8500 (N_8500,N_8377,N_8230);
nor U8501 (N_8501,N_8391,N_8338);
nor U8502 (N_8502,N_8399,N_8381);
or U8503 (N_8503,N_8377,N_8372);
or U8504 (N_8504,N_8299,N_8358);
and U8505 (N_8505,N_8252,N_8229);
xnor U8506 (N_8506,N_8326,N_8389);
xor U8507 (N_8507,N_8305,N_8396);
nand U8508 (N_8508,N_8300,N_8236);
nor U8509 (N_8509,N_8375,N_8386);
nand U8510 (N_8510,N_8368,N_8389);
xor U8511 (N_8511,N_8206,N_8340);
or U8512 (N_8512,N_8216,N_8280);
or U8513 (N_8513,N_8281,N_8232);
nand U8514 (N_8514,N_8361,N_8327);
xnor U8515 (N_8515,N_8234,N_8262);
or U8516 (N_8516,N_8223,N_8203);
xor U8517 (N_8517,N_8206,N_8288);
nand U8518 (N_8518,N_8206,N_8211);
or U8519 (N_8519,N_8390,N_8232);
or U8520 (N_8520,N_8386,N_8356);
or U8521 (N_8521,N_8290,N_8223);
nor U8522 (N_8522,N_8304,N_8266);
nor U8523 (N_8523,N_8282,N_8281);
or U8524 (N_8524,N_8316,N_8223);
xor U8525 (N_8525,N_8334,N_8344);
nor U8526 (N_8526,N_8318,N_8306);
nor U8527 (N_8527,N_8382,N_8320);
xor U8528 (N_8528,N_8203,N_8244);
nand U8529 (N_8529,N_8324,N_8387);
nand U8530 (N_8530,N_8377,N_8261);
nor U8531 (N_8531,N_8399,N_8230);
nand U8532 (N_8532,N_8386,N_8366);
xor U8533 (N_8533,N_8393,N_8371);
nand U8534 (N_8534,N_8267,N_8226);
and U8535 (N_8535,N_8230,N_8312);
nand U8536 (N_8536,N_8290,N_8309);
and U8537 (N_8537,N_8268,N_8239);
xor U8538 (N_8538,N_8297,N_8229);
or U8539 (N_8539,N_8318,N_8237);
and U8540 (N_8540,N_8390,N_8298);
and U8541 (N_8541,N_8268,N_8225);
nand U8542 (N_8542,N_8358,N_8397);
xor U8543 (N_8543,N_8377,N_8234);
xnor U8544 (N_8544,N_8317,N_8384);
xor U8545 (N_8545,N_8338,N_8396);
or U8546 (N_8546,N_8333,N_8322);
or U8547 (N_8547,N_8396,N_8372);
and U8548 (N_8548,N_8300,N_8337);
nor U8549 (N_8549,N_8286,N_8230);
nand U8550 (N_8550,N_8399,N_8303);
nand U8551 (N_8551,N_8264,N_8249);
nor U8552 (N_8552,N_8327,N_8350);
xor U8553 (N_8553,N_8301,N_8358);
nand U8554 (N_8554,N_8234,N_8346);
nand U8555 (N_8555,N_8225,N_8286);
or U8556 (N_8556,N_8303,N_8382);
nand U8557 (N_8557,N_8307,N_8338);
or U8558 (N_8558,N_8316,N_8228);
nand U8559 (N_8559,N_8238,N_8330);
or U8560 (N_8560,N_8375,N_8255);
and U8561 (N_8561,N_8386,N_8228);
xor U8562 (N_8562,N_8366,N_8343);
xnor U8563 (N_8563,N_8218,N_8284);
xnor U8564 (N_8564,N_8295,N_8290);
and U8565 (N_8565,N_8313,N_8220);
xnor U8566 (N_8566,N_8286,N_8354);
or U8567 (N_8567,N_8224,N_8339);
nand U8568 (N_8568,N_8292,N_8217);
nor U8569 (N_8569,N_8320,N_8310);
and U8570 (N_8570,N_8259,N_8227);
and U8571 (N_8571,N_8288,N_8228);
nor U8572 (N_8572,N_8354,N_8294);
or U8573 (N_8573,N_8299,N_8265);
or U8574 (N_8574,N_8363,N_8293);
xor U8575 (N_8575,N_8386,N_8344);
nand U8576 (N_8576,N_8344,N_8332);
nor U8577 (N_8577,N_8336,N_8252);
and U8578 (N_8578,N_8399,N_8227);
nand U8579 (N_8579,N_8224,N_8257);
nor U8580 (N_8580,N_8271,N_8248);
nor U8581 (N_8581,N_8381,N_8238);
nand U8582 (N_8582,N_8349,N_8345);
or U8583 (N_8583,N_8252,N_8382);
or U8584 (N_8584,N_8375,N_8265);
nand U8585 (N_8585,N_8337,N_8348);
and U8586 (N_8586,N_8221,N_8343);
nor U8587 (N_8587,N_8273,N_8395);
or U8588 (N_8588,N_8344,N_8351);
nor U8589 (N_8589,N_8287,N_8254);
xor U8590 (N_8590,N_8368,N_8360);
and U8591 (N_8591,N_8301,N_8399);
nor U8592 (N_8592,N_8270,N_8286);
nor U8593 (N_8593,N_8349,N_8213);
or U8594 (N_8594,N_8331,N_8340);
and U8595 (N_8595,N_8332,N_8378);
and U8596 (N_8596,N_8232,N_8301);
and U8597 (N_8597,N_8312,N_8263);
or U8598 (N_8598,N_8381,N_8207);
or U8599 (N_8599,N_8290,N_8224);
or U8600 (N_8600,N_8588,N_8536);
and U8601 (N_8601,N_8532,N_8413);
xor U8602 (N_8602,N_8489,N_8511);
xnor U8603 (N_8603,N_8432,N_8418);
nor U8604 (N_8604,N_8504,N_8550);
nor U8605 (N_8605,N_8499,N_8509);
nand U8606 (N_8606,N_8572,N_8575);
and U8607 (N_8607,N_8424,N_8444);
and U8608 (N_8608,N_8492,N_8515);
nor U8609 (N_8609,N_8480,N_8520);
nand U8610 (N_8610,N_8547,N_8516);
xnor U8611 (N_8611,N_8531,N_8401);
nand U8612 (N_8612,N_8574,N_8580);
or U8613 (N_8613,N_8420,N_8561);
nand U8614 (N_8614,N_8474,N_8417);
xnor U8615 (N_8615,N_8577,N_8522);
xnor U8616 (N_8616,N_8421,N_8579);
and U8617 (N_8617,N_8403,N_8568);
xnor U8618 (N_8618,N_8414,N_8528);
nand U8619 (N_8619,N_8517,N_8469);
nand U8620 (N_8620,N_8490,N_8422);
or U8621 (N_8621,N_8493,N_8497);
nand U8622 (N_8622,N_8491,N_8456);
nor U8623 (N_8623,N_8534,N_8518);
and U8624 (N_8624,N_8500,N_8448);
nor U8625 (N_8625,N_8440,N_8545);
nor U8626 (N_8626,N_8573,N_8569);
or U8627 (N_8627,N_8513,N_8533);
and U8628 (N_8628,N_8412,N_8478);
nor U8629 (N_8629,N_8481,N_8431);
nor U8630 (N_8630,N_8553,N_8584);
nand U8631 (N_8631,N_8484,N_8537);
or U8632 (N_8632,N_8597,N_8427);
nor U8633 (N_8633,N_8404,N_8514);
xor U8634 (N_8634,N_8461,N_8400);
or U8635 (N_8635,N_8529,N_8586);
nand U8636 (N_8636,N_8457,N_8555);
and U8637 (N_8637,N_8519,N_8433);
nor U8638 (N_8638,N_8472,N_8571);
nand U8639 (N_8639,N_8589,N_8566);
and U8640 (N_8640,N_8554,N_8479);
and U8641 (N_8641,N_8498,N_8523);
xnor U8642 (N_8642,N_8567,N_8423);
and U8643 (N_8643,N_8449,N_8544);
nor U8644 (N_8644,N_8596,N_8551);
or U8645 (N_8645,N_8512,N_8494);
or U8646 (N_8646,N_8446,N_8419);
nand U8647 (N_8647,N_8542,N_8443);
or U8648 (N_8648,N_8428,N_8510);
and U8649 (N_8649,N_8563,N_8447);
and U8650 (N_8650,N_8426,N_8408);
nand U8651 (N_8651,N_8546,N_8471);
or U8652 (N_8652,N_8496,N_8441);
nor U8653 (N_8653,N_8540,N_8436);
or U8654 (N_8654,N_8466,N_8486);
nor U8655 (N_8655,N_8530,N_8458);
nand U8656 (N_8656,N_8548,N_8525);
or U8657 (N_8657,N_8582,N_8488);
xnor U8658 (N_8658,N_8410,N_8508);
and U8659 (N_8659,N_8541,N_8442);
nor U8660 (N_8660,N_8592,N_8434);
and U8661 (N_8661,N_8465,N_8477);
xnor U8662 (N_8662,N_8587,N_8557);
nand U8663 (N_8663,N_8467,N_8459);
or U8664 (N_8664,N_8598,N_8460);
xor U8665 (N_8665,N_8565,N_8576);
and U8666 (N_8666,N_8556,N_8470);
and U8667 (N_8667,N_8570,N_8552);
nand U8668 (N_8668,N_8485,N_8411);
and U8669 (N_8669,N_8585,N_8503);
and U8670 (N_8670,N_8475,N_8591);
nand U8671 (N_8671,N_8437,N_8430);
nand U8672 (N_8672,N_8506,N_8558);
or U8673 (N_8673,N_8590,N_8524);
xnor U8674 (N_8674,N_8416,N_8463);
nand U8675 (N_8675,N_8483,N_8462);
xor U8676 (N_8676,N_8562,N_8539);
or U8677 (N_8677,N_8473,N_8450);
nor U8678 (N_8678,N_8445,N_8452);
nand U8679 (N_8679,N_8527,N_8564);
nand U8680 (N_8680,N_8405,N_8495);
xor U8681 (N_8681,N_8464,N_8581);
nor U8682 (N_8682,N_8502,N_8583);
xnor U8683 (N_8683,N_8468,N_8409);
or U8684 (N_8684,N_8559,N_8595);
nor U8685 (N_8685,N_8507,N_8487);
or U8686 (N_8686,N_8425,N_8593);
nor U8687 (N_8687,N_8439,N_8526);
nand U8688 (N_8688,N_8453,N_8476);
xor U8689 (N_8689,N_8560,N_8451);
xor U8690 (N_8690,N_8578,N_8599);
or U8691 (N_8691,N_8429,N_8501);
or U8692 (N_8692,N_8406,N_8415);
nand U8693 (N_8693,N_8455,N_8594);
nor U8694 (N_8694,N_8549,N_8535);
or U8695 (N_8695,N_8543,N_8454);
nor U8696 (N_8696,N_8521,N_8538);
or U8697 (N_8697,N_8435,N_8407);
nand U8698 (N_8698,N_8438,N_8482);
nand U8699 (N_8699,N_8402,N_8505);
xnor U8700 (N_8700,N_8586,N_8534);
nand U8701 (N_8701,N_8517,N_8555);
nand U8702 (N_8702,N_8453,N_8428);
or U8703 (N_8703,N_8487,N_8541);
nor U8704 (N_8704,N_8578,N_8505);
xor U8705 (N_8705,N_8489,N_8507);
xor U8706 (N_8706,N_8488,N_8595);
xnor U8707 (N_8707,N_8541,N_8581);
or U8708 (N_8708,N_8468,N_8528);
xnor U8709 (N_8709,N_8428,N_8557);
and U8710 (N_8710,N_8517,N_8592);
nor U8711 (N_8711,N_8581,N_8514);
and U8712 (N_8712,N_8469,N_8588);
and U8713 (N_8713,N_8581,N_8450);
or U8714 (N_8714,N_8531,N_8510);
nand U8715 (N_8715,N_8553,N_8483);
nor U8716 (N_8716,N_8546,N_8548);
xnor U8717 (N_8717,N_8466,N_8433);
or U8718 (N_8718,N_8575,N_8484);
nor U8719 (N_8719,N_8478,N_8499);
nor U8720 (N_8720,N_8443,N_8460);
or U8721 (N_8721,N_8462,N_8455);
xnor U8722 (N_8722,N_8507,N_8430);
nand U8723 (N_8723,N_8441,N_8587);
or U8724 (N_8724,N_8566,N_8514);
nand U8725 (N_8725,N_8494,N_8489);
xor U8726 (N_8726,N_8515,N_8569);
nor U8727 (N_8727,N_8479,N_8414);
nor U8728 (N_8728,N_8467,N_8587);
nand U8729 (N_8729,N_8514,N_8562);
or U8730 (N_8730,N_8596,N_8471);
nor U8731 (N_8731,N_8525,N_8572);
and U8732 (N_8732,N_8450,N_8582);
nand U8733 (N_8733,N_8484,N_8443);
nand U8734 (N_8734,N_8499,N_8588);
xnor U8735 (N_8735,N_8436,N_8521);
nand U8736 (N_8736,N_8464,N_8519);
nor U8737 (N_8737,N_8582,N_8550);
nor U8738 (N_8738,N_8438,N_8591);
nand U8739 (N_8739,N_8557,N_8546);
nor U8740 (N_8740,N_8583,N_8594);
nand U8741 (N_8741,N_8505,N_8467);
xor U8742 (N_8742,N_8426,N_8401);
nor U8743 (N_8743,N_8504,N_8409);
and U8744 (N_8744,N_8586,N_8563);
nand U8745 (N_8745,N_8484,N_8513);
nand U8746 (N_8746,N_8511,N_8499);
nand U8747 (N_8747,N_8569,N_8422);
nand U8748 (N_8748,N_8596,N_8591);
and U8749 (N_8749,N_8426,N_8566);
xnor U8750 (N_8750,N_8453,N_8545);
nor U8751 (N_8751,N_8565,N_8468);
xor U8752 (N_8752,N_8413,N_8558);
nand U8753 (N_8753,N_8438,N_8585);
nand U8754 (N_8754,N_8484,N_8439);
or U8755 (N_8755,N_8494,N_8561);
xor U8756 (N_8756,N_8432,N_8483);
or U8757 (N_8757,N_8511,N_8471);
nand U8758 (N_8758,N_8565,N_8597);
nand U8759 (N_8759,N_8434,N_8498);
or U8760 (N_8760,N_8534,N_8540);
nand U8761 (N_8761,N_8593,N_8490);
xnor U8762 (N_8762,N_8405,N_8401);
and U8763 (N_8763,N_8437,N_8543);
and U8764 (N_8764,N_8460,N_8456);
or U8765 (N_8765,N_8528,N_8456);
nand U8766 (N_8766,N_8486,N_8534);
or U8767 (N_8767,N_8412,N_8421);
nand U8768 (N_8768,N_8557,N_8461);
and U8769 (N_8769,N_8509,N_8422);
nand U8770 (N_8770,N_8529,N_8472);
or U8771 (N_8771,N_8421,N_8576);
xor U8772 (N_8772,N_8494,N_8496);
or U8773 (N_8773,N_8408,N_8503);
nor U8774 (N_8774,N_8567,N_8465);
or U8775 (N_8775,N_8506,N_8519);
nand U8776 (N_8776,N_8545,N_8500);
or U8777 (N_8777,N_8590,N_8485);
nor U8778 (N_8778,N_8559,N_8460);
nand U8779 (N_8779,N_8542,N_8586);
nor U8780 (N_8780,N_8581,N_8403);
nor U8781 (N_8781,N_8404,N_8490);
xor U8782 (N_8782,N_8405,N_8533);
nand U8783 (N_8783,N_8565,N_8554);
xor U8784 (N_8784,N_8513,N_8482);
nand U8785 (N_8785,N_8428,N_8478);
or U8786 (N_8786,N_8497,N_8433);
or U8787 (N_8787,N_8514,N_8567);
nor U8788 (N_8788,N_8466,N_8476);
and U8789 (N_8789,N_8410,N_8527);
and U8790 (N_8790,N_8514,N_8463);
nand U8791 (N_8791,N_8422,N_8477);
and U8792 (N_8792,N_8417,N_8585);
and U8793 (N_8793,N_8455,N_8422);
nand U8794 (N_8794,N_8499,N_8506);
xor U8795 (N_8795,N_8567,N_8490);
or U8796 (N_8796,N_8525,N_8500);
nand U8797 (N_8797,N_8582,N_8482);
and U8798 (N_8798,N_8508,N_8505);
xor U8799 (N_8799,N_8458,N_8525);
xor U8800 (N_8800,N_8681,N_8779);
nand U8801 (N_8801,N_8795,N_8704);
xnor U8802 (N_8802,N_8773,N_8609);
nor U8803 (N_8803,N_8613,N_8735);
nand U8804 (N_8804,N_8719,N_8635);
nand U8805 (N_8805,N_8710,N_8682);
and U8806 (N_8806,N_8686,N_8770);
nor U8807 (N_8807,N_8684,N_8783);
nand U8808 (N_8808,N_8623,N_8722);
or U8809 (N_8809,N_8756,N_8734);
xnor U8810 (N_8810,N_8705,N_8780);
nor U8811 (N_8811,N_8668,N_8644);
xor U8812 (N_8812,N_8607,N_8754);
nand U8813 (N_8813,N_8799,N_8778);
nor U8814 (N_8814,N_8655,N_8712);
nor U8815 (N_8815,N_8670,N_8709);
and U8816 (N_8816,N_8737,N_8765);
nand U8817 (N_8817,N_8660,N_8747);
and U8818 (N_8818,N_8726,N_8763);
nor U8819 (N_8819,N_8720,N_8600);
nor U8820 (N_8820,N_8624,N_8714);
nand U8821 (N_8821,N_8619,N_8713);
or U8822 (N_8822,N_8627,N_8757);
nand U8823 (N_8823,N_8614,N_8601);
nand U8824 (N_8824,N_8733,N_8741);
xor U8825 (N_8825,N_8758,N_8736);
or U8826 (N_8826,N_8611,N_8731);
and U8827 (N_8827,N_8698,N_8787);
xnor U8828 (N_8828,N_8716,N_8762);
or U8829 (N_8829,N_8798,N_8746);
xor U8830 (N_8830,N_8774,N_8729);
or U8831 (N_8831,N_8634,N_8771);
or U8832 (N_8832,N_8724,N_8694);
or U8833 (N_8833,N_8632,N_8687);
nand U8834 (N_8834,N_8761,N_8692);
or U8835 (N_8835,N_8671,N_8752);
and U8836 (N_8836,N_8631,N_8702);
xnor U8837 (N_8837,N_8633,N_8677);
nor U8838 (N_8838,N_8637,N_8739);
or U8839 (N_8839,N_8793,N_8683);
nor U8840 (N_8840,N_8777,N_8674);
xor U8841 (N_8841,N_8646,N_8603);
xnor U8842 (N_8842,N_8663,N_8753);
and U8843 (N_8843,N_8744,N_8703);
nor U8844 (N_8844,N_8768,N_8728);
xor U8845 (N_8845,N_8658,N_8662);
and U8846 (N_8846,N_8749,N_8653);
or U8847 (N_8847,N_8650,N_8708);
nand U8848 (N_8848,N_8678,N_8630);
and U8849 (N_8849,N_8654,N_8665);
xnor U8850 (N_8850,N_8732,N_8742);
and U8851 (N_8851,N_8680,N_8738);
nand U8852 (N_8852,N_8789,N_8782);
nor U8853 (N_8853,N_8786,N_8626);
nand U8854 (N_8854,N_8775,N_8664);
or U8855 (N_8855,N_8723,N_8750);
nor U8856 (N_8856,N_8755,N_8781);
nand U8857 (N_8857,N_8760,N_8673);
or U8858 (N_8858,N_8718,N_8791);
and U8859 (N_8859,N_8675,N_8639);
or U8860 (N_8860,N_8693,N_8797);
nand U8861 (N_8861,N_8676,N_8641);
nor U8862 (N_8862,N_8730,N_8743);
and U8863 (N_8863,N_8659,N_8657);
or U8864 (N_8864,N_8605,N_8651);
and U8865 (N_8865,N_8706,N_8608);
xnor U8866 (N_8866,N_8669,N_8690);
or U8867 (N_8867,N_8745,N_8604);
xnor U8868 (N_8868,N_8790,N_8636);
nand U8869 (N_8869,N_8602,N_8794);
xor U8870 (N_8870,N_8785,N_8764);
and U8871 (N_8871,N_8772,N_8751);
or U8872 (N_8872,N_8740,N_8645);
nand U8873 (N_8873,N_8784,N_8699);
nor U8874 (N_8874,N_8616,N_8796);
nor U8875 (N_8875,N_8647,N_8685);
nand U8876 (N_8876,N_8622,N_8721);
xnor U8877 (N_8877,N_8649,N_8615);
and U8878 (N_8878,N_8792,N_8767);
or U8879 (N_8879,N_8612,N_8725);
and U8880 (N_8880,N_8707,N_8620);
or U8881 (N_8881,N_8696,N_8691);
nand U8882 (N_8882,N_8640,N_8688);
nor U8883 (N_8883,N_8638,N_8629);
or U8884 (N_8884,N_8610,N_8695);
and U8885 (N_8885,N_8661,N_8625);
nor U8886 (N_8886,N_8618,N_8689);
xnor U8887 (N_8887,N_8656,N_8727);
xor U8888 (N_8888,N_8666,N_8606);
xor U8889 (N_8889,N_8759,N_8700);
xnor U8890 (N_8890,N_8697,N_8748);
xnor U8891 (N_8891,N_8766,N_8717);
nand U8892 (N_8892,N_8701,N_8617);
nor U8893 (N_8893,N_8776,N_8672);
nor U8894 (N_8894,N_8667,N_8652);
and U8895 (N_8895,N_8788,N_8715);
xnor U8896 (N_8896,N_8621,N_8769);
or U8897 (N_8897,N_8648,N_8628);
xnor U8898 (N_8898,N_8643,N_8642);
and U8899 (N_8899,N_8679,N_8711);
nor U8900 (N_8900,N_8789,N_8707);
nand U8901 (N_8901,N_8782,N_8710);
xor U8902 (N_8902,N_8660,N_8665);
and U8903 (N_8903,N_8793,N_8728);
or U8904 (N_8904,N_8770,N_8680);
or U8905 (N_8905,N_8697,N_8735);
nand U8906 (N_8906,N_8777,N_8788);
and U8907 (N_8907,N_8600,N_8633);
nand U8908 (N_8908,N_8628,N_8796);
nor U8909 (N_8909,N_8754,N_8640);
nand U8910 (N_8910,N_8663,N_8725);
nand U8911 (N_8911,N_8606,N_8734);
and U8912 (N_8912,N_8647,N_8764);
nand U8913 (N_8913,N_8799,N_8708);
xnor U8914 (N_8914,N_8622,N_8621);
and U8915 (N_8915,N_8719,N_8616);
nand U8916 (N_8916,N_8733,N_8725);
nor U8917 (N_8917,N_8610,N_8738);
and U8918 (N_8918,N_8649,N_8653);
xor U8919 (N_8919,N_8770,N_8742);
and U8920 (N_8920,N_8615,N_8769);
or U8921 (N_8921,N_8725,N_8666);
nand U8922 (N_8922,N_8652,N_8672);
and U8923 (N_8923,N_8731,N_8720);
or U8924 (N_8924,N_8616,N_8716);
and U8925 (N_8925,N_8720,N_8707);
or U8926 (N_8926,N_8732,N_8659);
nand U8927 (N_8927,N_8738,N_8685);
and U8928 (N_8928,N_8704,N_8734);
nor U8929 (N_8929,N_8608,N_8749);
and U8930 (N_8930,N_8710,N_8603);
nor U8931 (N_8931,N_8739,N_8796);
xor U8932 (N_8932,N_8667,N_8685);
nor U8933 (N_8933,N_8653,N_8786);
nand U8934 (N_8934,N_8658,N_8704);
nand U8935 (N_8935,N_8629,N_8616);
or U8936 (N_8936,N_8693,N_8672);
or U8937 (N_8937,N_8631,N_8637);
nand U8938 (N_8938,N_8744,N_8705);
nor U8939 (N_8939,N_8727,N_8618);
xnor U8940 (N_8940,N_8696,N_8682);
nor U8941 (N_8941,N_8688,N_8684);
and U8942 (N_8942,N_8681,N_8612);
and U8943 (N_8943,N_8737,N_8680);
and U8944 (N_8944,N_8600,N_8658);
xor U8945 (N_8945,N_8766,N_8740);
and U8946 (N_8946,N_8680,N_8684);
nand U8947 (N_8947,N_8715,N_8615);
or U8948 (N_8948,N_8748,N_8691);
xnor U8949 (N_8949,N_8689,N_8635);
or U8950 (N_8950,N_8760,N_8798);
nor U8951 (N_8951,N_8646,N_8752);
and U8952 (N_8952,N_8739,N_8774);
xnor U8953 (N_8953,N_8642,N_8646);
nand U8954 (N_8954,N_8756,N_8715);
nand U8955 (N_8955,N_8799,N_8601);
nand U8956 (N_8956,N_8681,N_8700);
xnor U8957 (N_8957,N_8765,N_8616);
xnor U8958 (N_8958,N_8751,N_8721);
nor U8959 (N_8959,N_8679,N_8645);
or U8960 (N_8960,N_8603,N_8618);
xor U8961 (N_8961,N_8673,N_8725);
nor U8962 (N_8962,N_8750,N_8680);
xor U8963 (N_8963,N_8725,N_8750);
xor U8964 (N_8964,N_8673,N_8762);
and U8965 (N_8965,N_8641,N_8748);
and U8966 (N_8966,N_8733,N_8652);
or U8967 (N_8967,N_8610,N_8728);
nor U8968 (N_8968,N_8608,N_8639);
and U8969 (N_8969,N_8783,N_8645);
nor U8970 (N_8970,N_8754,N_8636);
or U8971 (N_8971,N_8710,N_8613);
xnor U8972 (N_8972,N_8637,N_8777);
nand U8973 (N_8973,N_8604,N_8735);
or U8974 (N_8974,N_8772,N_8786);
and U8975 (N_8975,N_8618,N_8685);
xnor U8976 (N_8976,N_8719,N_8660);
nor U8977 (N_8977,N_8716,N_8612);
and U8978 (N_8978,N_8793,N_8686);
and U8979 (N_8979,N_8796,N_8775);
nor U8980 (N_8980,N_8603,N_8634);
and U8981 (N_8981,N_8621,N_8754);
or U8982 (N_8982,N_8655,N_8707);
nor U8983 (N_8983,N_8627,N_8606);
or U8984 (N_8984,N_8729,N_8601);
xor U8985 (N_8985,N_8780,N_8742);
nand U8986 (N_8986,N_8762,N_8638);
and U8987 (N_8987,N_8612,N_8785);
nor U8988 (N_8988,N_8764,N_8729);
nand U8989 (N_8989,N_8668,N_8754);
or U8990 (N_8990,N_8729,N_8609);
nor U8991 (N_8991,N_8760,N_8629);
xnor U8992 (N_8992,N_8748,N_8602);
nand U8993 (N_8993,N_8697,N_8722);
or U8994 (N_8994,N_8760,N_8656);
or U8995 (N_8995,N_8782,N_8722);
and U8996 (N_8996,N_8702,N_8710);
nand U8997 (N_8997,N_8711,N_8608);
nand U8998 (N_8998,N_8729,N_8634);
nand U8999 (N_8999,N_8694,N_8732);
or U9000 (N_9000,N_8869,N_8955);
and U9001 (N_9001,N_8854,N_8927);
nor U9002 (N_9002,N_8842,N_8861);
or U9003 (N_9003,N_8878,N_8896);
or U9004 (N_9004,N_8894,N_8828);
xnor U9005 (N_9005,N_8888,N_8941);
and U9006 (N_9006,N_8960,N_8841);
xnor U9007 (N_9007,N_8890,N_8997);
nor U9008 (N_9008,N_8931,N_8942);
or U9009 (N_9009,N_8994,N_8915);
or U9010 (N_9010,N_8911,N_8956);
nor U9011 (N_9011,N_8983,N_8933);
nor U9012 (N_9012,N_8918,N_8971);
nor U9013 (N_9013,N_8961,N_8907);
and U9014 (N_9014,N_8923,N_8990);
nor U9015 (N_9015,N_8967,N_8852);
nor U9016 (N_9016,N_8993,N_8995);
xor U9017 (N_9017,N_8953,N_8949);
or U9018 (N_9018,N_8935,N_8800);
nor U9019 (N_9019,N_8881,N_8908);
and U9020 (N_9020,N_8999,N_8932);
or U9021 (N_9021,N_8906,N_8959);
or U9022 (N_9022,N_8975,N_8872);
nand U9023 (N_9023,N_8801,N_8972);
xnor U9024 (N_9024,N_8851,N_8985);
or U9025 (N_9025,N_8807,N_8864);
nand U9026 (N_9026,N_8823,N_8880);
or U9027 (N_9027,N_8865,N_8847);
and U9028 (N_9028,N_8899,N_8969);
xnor U9029 (N_9029,N_8898,N_8853);
nand U9030 (N_9030,N_8947,N_8944);
xor U9031 (N_9031,N_8929,N_8860);
and U9032 (N_9032,N_8885,N_8982);
and U9033 (N_9033,N_8919,N_8824);
xor U9034 (N_9034,N_8876,N_8977);
or U9035 (N_9035,N_8958,N_8889);
nor U9036 (N_9036,N_8968,N_8815);
and U9037 (N_9037,N_8901,N_8886);
and U9038 (N_9038,N_8962,N_8980);
and U9039 (N_9039,N_8820,N_8914);
nand U9040 (N_9040,N_8809,N_8863);
nor U9041 (N_9041,N_8897,N_8875);
and U9042 (N_9042,N_8829,N_8979);
and U9043 (N_9043,N_8883,N_8964);
nor U9044 (N_9044,N_8974,N_8806);
xor U9045 (N_9045,N_8945,N_8804);
nand U9046 (N_9046,N_8939,N_8818);
and U9047 (N_9047,N_8849,N_8873);
xor U9048 (N_9048,N_8904,N_8805);
and U9049 (N_9049,N_8887,N_8871);
nor U9050 (N_9050,N_8819,N_8884);
xor U9051 (N_9051,N_8905,N_8821);
or U9052 (N_9052,N_8912,N_8848);
or U9053 (N_9053,N_8991,N_8830);
nand U9054 (N_9054,N_8943,N_8930);
xnor U9055 (N_9055,N_8840,N_8917);
nor U9056 (N_9056,N_8893,N_8817);
nor U9057 (N_9057,N_8855,N_8845);
or U9058 (N_9058,N_8965,N_8910);
nand U9059 (N_9059,N_8903,N_8836);
nand U9060 (N_9060,N_8822,N_8812);
xor U9061 (N_9061,N_8938,N_8992);
and U9062 (N_9062,N_8986,N_8867);
xnor U9063 (N_9063,N_8973,N_8835);
and U9064 (N_9064,N_8877,N_8837);
xor U9065 (N_9065,N_8989,N_8802);
or U9066 (N_9066,N_8952,N_8882);
xor U9067 (N_9067,N_8978,N_8866);
nand U9068 (N_9068,N_8843,N_8987);
nor U9069 (N_9069,N_8838,N_8936);
or U9070 (N_9070,N_8970,N_8921);
xor U9071 (N_9071,N_8862,N_8909);
and U9072 (N_9072,N_8874,N_8834);
nor U9073 (N_9073,N_8957,N_8966);
nor U9074 (N_9074,N_8856,N_8858);
or U9075 (N_9075,N_8839,N_8900);
and U9076 (N_9076,N_8844,N_8832);
or U9077 (N_9077,N_8826,N_8924);
nor U9078 (N_9078,N_8827,N_8963);
xor U9079 (N_9079,N_8868,N_8940);
and U9080 (N_9080,N_8846,N_8988);
nand U9081 (N_9081,N_8998,N_8996);
xnor U9082 (N_9082,N_8926,N_8925);
nor U9083 (N_9083,N_8976,N_8811);
xor U9084 (N_9084,N_8937,N_8870);
or U9085 (N_9085,N_8833,N_8803);
or U9086 (N_9086,N_8948,N_8814);
xnor U9087 (N_9087,N_8895,N_8954);
xor U9088 (N_9088,N_8891,N_8816);
and U9089 (N_9089,N_8920,N_8813);
nor U9090 (N_9090,N_8928,N_8808);
xor U9091 (N_9091,N_8951,N_8922);
nand U9092 (N_9092,N_8984,N_8892);
and U9093 (N_9093,N_8946,N_8825);
nand U9094 (N_9094,N_8913,N_8857);
and U9095 (N_9095,N_8950,N_8850);
nand U9096 (N_9096,N_8934,N_8879);
nor U9097 (N_9097,N_8859,N_8831);
and U9098 (N_9098,N_8810,N_8902);
xnor U9099 (N_9099,N_8916,N_8981);
and U9100 (N_9100,N_8821,N_8837);
nor U9101 (N_9101,N_8881,N_8842);
nand U9102 (N_9102,N_8823,N_8914);
xor U9103 (N_9103,N_8846,N_8995);
nor U9104 (N_9104,N_8872,N_8831);
or U9105 (N_9105,N_8845,N_8993);
and U9106 (N_9106,N_8884,N_8847);
nand U9107 (N_9107,N_8850,N_8804);
and U9108 (N_9108,N_8998,N_8896);
nor U9109 (N_9109,N_8970,N_8852);
and U9110 (N_9110,N_8981,N_8833);
or U9111 (N_9111,N_8917,N_8951);
and U9112 (N_9112,N_8973,N_8994);
and U9113 (N_9113,N_8903,N_8951);
nand U9114 (N_9114,N_8826,N_8837);
and U9115 (N_9115,N_8836,N_8816);
nand U9116 (N_9116,N_8956,N_8831);
or U9117 (N_9117,N_8906,N_8944);
or U9118 (N_9118,N_8960,N_8878);
nand U9119 (N_9119,N_8939,N_8950);
xor U9120 (N_9120,N_8840,N_8913);
or U9121 (N_9121,N_8865,N_8883);
or U9122 (N_9122,N_8955,N_8854);
nand U9123 (N_9123,N_8973,N_8903);
and U9124 (N_9124,N_8805,N_8802);
nor U9125 (N_9125,N_8817,N_8995);
nand U9126 (N_9126,N_8876,N_8829);
xor U9127 (N_9127,N_8874,N_8902);
or U9128 (N_9128,N_8903,N_8888);
and U9129 (N_9129,N_8877,N_8841);
nor U9130 (N_9130,N_8899,N_8998);
nor U9131 (N_9131,N_8917,N_8833);
xor U9132 (N_9132,N_8902,N_8961);
or U9133 (N_9133,N_8951,N_8807);
nand U9134 (N_9134,N_8813,N_8912);
xor U9135 (N_9135,N_8900,N_8855);
or U9136 (N_9136,N_8850,N_8986);
xor U9137 (N_9137,N_8934,N_8874);
nor U9138 (N_9138,N_8805,N_8979);
or U9139 (N_9139,N_8817,N_8948);
or U9140 (N_9140,N_8960,N_8981);
or U9141 (N_9141,N_8934,N_8951);
xor U9142 (N_9142,N_8815,N_8940);
and U9143 (N_9143,N_8983,N_8906);
xor U9144 (N_9144,N_8951,N_8945);
and U9145 (N_9145,N_8822,N_8862);
and U9146 (N_9146,N_8845,N_8801);
xnor U9147 (N_9147,N_8842,N_8963);
or U9148 (N_9148,N_8929,N_8988);
xor U9149 (N_9149,N_8895,N_8813);
nor U9150 (N_9150,N_8940,N_8812);
nor U9151 (N_9151,N_8826,N_8966);
and U9152 (N_9152,N_8910,N_8826);
and U9153 (N_9153,N_8974,N_8865);
xnor U9154 (N_9154,N_8818,N_8995);
nor U9155 (N_9155,N_8805,N_8989);
xnor U9156 (N_9156,N_8830,N_8864);
and U9157 (N_9157,N_8959,N_8971);
nor U9158 (N_9158,N_8907,N_8841);
nand U9159 (N_9159,N_8973,N_8953);
nor U9160 (N_9160,N_8983,N_8874);
xor U9161 (N_9161,N_8897,N_8830);
and U9162 (N_9162,N_8829,N_8955);
nor U9163 (N_9163,N_8834,N_8923);
nand U9164 (N_9164,N_8994,N_8933);
or U9165 (N_9165,N_8936,N_8893);
xnor U9166 (N_9166,N_8864,N_8884);
or U9167 (N_9167,N_8813,N_8937);
xor U9168 (N_9168,N_8990,N_8968);
or U9169 (N_9169,N_8962,N_8828);
or U9170 (N_9170,N_8952,N_8860);
xor U9171 (N_9171,N_8852,N_8839);
nor U9172 (N_9172,N_8904,N_8887);
nand U9173 (N_9173,N_8842,N_8800);
nand U9174 (N_9174,N_8990,N_8935);
xnor U9175 (N_9175,N_8838,N_8800);
or U9176 (N_9176,N_8837,N_8866);
nand U9177 (N_9177,N_8928,N_8931);
nor U9178 (N_9178,N_8889,N_8837);
nand U9179 (N_9179,N_8926,N_8902);
xnor U9180 (N_9180,N_8995,N_8899);
or U9181 (N_9181,N_8838,N_8997);
and U9182 (N_9182,N_8874,N_8954);
and U9183 (N_9183,N_8858,N_8986);
xor U9184 (N_9184,N_8819,N_8879);
nor U9185 (N_9185,N_8891,N_8855);
nor U9186 (N_9186,N_8885,N_8996);
nand U9187 (N_9187,N_8894,N_8866);
or U9188 (N_9188,N_8901,N_8995);
nand U9189 (N_9189,N_8899,N_8975);
nor U9190 (N_9190,N_8863,N_8848);
nor U9191 (N_9191,N_8865,N_8969);
xor U9192 (N_9192,N_8979,N_8817);
nand U9193 (N_9193,N_8930,N_8979);
and U9194 (N_9194,N_8918,N_8926);
nand U9195 (N_9195,N_8939,N_8848);
nand U9196 (N_9196,N_8930,N_8823);
nand U9197 (N_9197,N_8878,N_8996);
xor U9198 (N_9198,N_8891,N_8954);
nor U9199 (N_9199,N_8905,N_8899);
and U9200 (N_9200,N_9184,N_9095);
nand U9201 (N_9201,N_9139,N_9084);
nand U9202 (N_9202,N_9129,N_9058);
and U9203 (N_9203,N_9008,N_9038);
nor U9204 (N_9204,N_9002,N_9180);
xor U9205 (N_9205,N_9043,N_9020);
or U9206 (N_9206,N_9185,N_9155);
nand U9207 (N_9207,N_9081,N_9111);
nand U9208 (N_9208,N_9191,N_9103);
or U9209 (N_9209,N_9036,N_9074);
nor U9210 (N_9210,N_9161,N_9116);
nor U9211 (N_9211,N_9092,N_9153);
and U9212 (N_9212,N_9018,N_9170);
and U9213 (N_9213,N_9086,N_9156);
xor U9214 (N_9214,N_9113,N_9188);
xnor U9215 (N_9215,N_9104,N_9179);
or U9216 (N_9216,N_9112,N_9011);
or U9217 (N_9217,N_9187,N_9087);
nor U9218 (N_9218,N_9046,N_9101);
nor U9219 (N_9219,N_9026,N_9154);
or U9220 (N_9220,N_9067,N_9133);
xor U9221 (N_9221,N_9048,N_9182);
or U9222 (N_9222,N_9031,N_9000);
and U9223 (N_9223,N_9121,N_9013);
nor U9224 (N_9224,N_9198,N_9158);
nor U9225 (N_9225,N_9049,N_9091);
or U9226 (N_9226,N_9077,N_9119);
nand U9227 (N_9227,N_9063,N_9047);
nand U9228 (N_9228,N_9131,N_9093);
or U9229 (N_9229,N_9145,N_9085);
or U9230 (N_9230,N_9127,N_9022);
nand U9231 (N_9231,N_9078,N_9171);
or U9232 (N_9232,N_9199,N_9007);
or U9233 (N_9233,N_9105,N_9053);
or U9234 (N_9234,N_9073,N_9109);
nand U9235 (N_9235,N_9146,N_9189);
nand U9236 (N_9236,N_9122,N_9186);
nand U9237 (N_9237,N_9001,N_9066);
and U9238 (N_9238,N_9089,N_9037);
nor U9239 (N_9239,N_9166,N_9003);
xnor U9240 (N_9240,N_9094,N_9017);
nor U9241 (N_9241,N_9107,N_9079);
or U9242 (N_9242,N_9080,N_9172);
nand U9243 (N_9243,N_9052,N_9065);
or U9244 (N_9244,N_9135,N_9138);
and U9245 (N_9245,N_9019,N_9099);
nand U9246 (N_9246,N_9082,N_9176);
nor U9247 (N_9247,N_9056,N_9150);
xnor U9248 (N_9248,N_9123,N_9090);
or U9249 (N_9249,N_9132,N_9012);
nand U9250 (N_9250,N_9190,N_9054);
or U9251 (N_9251,N_9195,N_9169);
nor U9252 (N_9252,N_9004,N_9196);
or U9253 (N_9253,N_9192,N_9115);
nand U9254 (N_9254,N_9157,N_9027);
or U9255 (N_9255,N_9005,N_9042);
or U9256 (N_9256,N_9030,N_9024);
or U9257 (N_9257,N_9174,N_9194);
or U9258 (N_9258,N_9039,N_9168);
nor U9259 (N_9259,N_9028,N_9143);
nor U9260 (N_9260,N_9057,N_9147);
nand U9261 (N_9261,N_9126,N_9140);
or U9262 (N_9262,N_9137,N_9050);
xor U9263 (N_9263,N_9021,N_9088);
xor U9264 (N_9264,N_9118,N_9108);
xnor U9265 (N_9265,N_9059,N_9175);
or U9266 (N_9266,N_9102,N_9162);
and U9267 (N_9267,N_9100,N_9136);
and U9268 (N_9268,N_9183,N_9096);
and U9269 (N_9269,N_9193,N_9044);
nor U9270 (N_9270,N_9072,N_9159);
or U9271 (N_9271,N_9097,N_9144);
xor U9272 (N_9272,N_9141,N_9151);
or U9273 (N_9273,N_9040,N_9148);
nand U9274 (N_9274,N_9060,N_9164);
nor U9275 (N_9275,N_9098,N_9023);
nand U9276 (N_9276,N_9106,N_9177);
and U9277 (N_9277,N_9006,N_9173);
nor U9278 (N_9278,N_9142,N_9014);
nor U9279 (N_9279,N_9062,N_9016);
nand U9280 (N_9280,N_9120,N_9076);
nor U9281 (N_9281,N_9015,N_9070);
or U9282 (N_9282,N_9114,N_9110);
and U9283 (N_9283,N_9051,N_9083);
nand U9284 (N_9284,N_9068,N_9041);
xor U9285 (N_9285,N_9009,N_9178);
nor U9286 (N_9286,N_9045,N_9055);
and U9287 (N_9287,N_9069,N_9117);
and U9288 (N_9288,N_9181,N_9160);
or U9289 (N_9289,N_9149,N_9033);
xnor U9290 (N_9290,N_9125,N_9075);
nor U9291 (N_9291,N_9034,N_9064);
or U9292 (N_9292,N_9071,N_9128);
or U9293 (N_9293,N_9010,N_9025);
and U9294 (N_9294,N_9035,N_9167);
nor U9295 (N_9295,N_9197,N_9032);
nand U9296 (N_9296,N_9165,N_9163);
or U9297 (N_9297,N_9124,N_9152);
and U9298 (N_9298,N_9130,N_9134);
nand U9299 (N_9299,N_9061,N_9029);
nand U9300 (N_9300,N_9099,N_9067);
xor U9301 (N_9301,N_9064,N_9005);
nor U9302 (N_9302,N_9096,N_9071);
or U9303 (N_9303,N_9129,N_9075);
and U9304 (N_9304,N_9136,N_9156);
and U9305 (N_9305,N_9021,N_9150);
or U9306 (N_9306,N_9161,N_9085);
nand U9307 (N_9307,N_9192,N_9110);
nor U9308 (N_9308,N_9041,N_9151);
or U9309 (N_9309,N_9181,N_9062);
or U9310 (N_9310,N_9093,N_9120);
nor U9311 (N_9311,N_9127,N_9152);
or U9312 (N_9312,N_9137,N_9127);
xnor U9313 (N_9313,N_9090,N_9051);
nand U9314 (N_9314,N_9159,N_9054);
nor U9315 (N_9315,N_9047,N_9045);
nor U9316 (N_9316,N_9000,N_9054);
and U9317 (N_9317,N_9008,N_9119);
nor U9318 (N_9318,N_9176,N_9017);
nand U9319 (N_9319,N_9078,N_9060);
nand U9320 (N_9320,N_9017,N_9153);
nand U9321 (N_9321,N_9165,N_9091);
nor U9322 (N_9322,N_9064,N_9053);
and U9323 (N_9323,N_9100,N_9121);
or U9324 (N_9324,N_9127,N_9083);
nor U9325 (N_9325,N_9072,N_9068);
xor U9326 (N_9326,N_9000,N_9049);
xnor U9327 (N_9327,N_9134,N_9027);
nor U9328 (N_9328,N_9085,N_9092);
nand U9329 (N_9329,N_9004,N_9014);
and U9330 (N_9330,N_9100,N_9159);
nor U9331 (N_9331,N_9088,N_9110);
and U9332 (N_9332,N_9185,N_9070);
nor U9333 (N_9333,N_9088,N_9116);
or U9334 (N_9334,N_9197,N_9199);
nand U9335 (N_9335,N_9074,N_9094);
xor U9336 (N_9336,N_9007,N_9013);
or U9337 (N_9337,N_9066,N_9053);
xor U9338 (N_9338,N_9180,N_9102);
nor U9339 (N_9339,N_9140,N_9163);
nor U9340 (N_9340,N_9085,N_9055);
and U9341 (N_9341,N_9059,N_9163);
and U9342 (N_9342,N_9018,N_9017);
or U9343 (N_9343,N_9012,N_9136);
nor U9344 (N_9344,N_9026,N_9140);
nand U9345 (N_9345,N_9051,N_9132);
nand U9346 (N_9346,N_9063,N_9115);
or U9347 (N_9347,N_9064,N_9111);
xor U9348 (N_9348,N_9021,N_9004);
and U9349 (N_9349,N_9025,N_9084);
and U9350 (N_9350,N_9024,N_9158);
and U9351 (N_9351,N_9078,N_9046);
and U9352 (N_9352,N_9057,N_9024);
nor U9353 (N_9353,N_9033,N_9041);
nand U9354 (N_9354,N_9179,N_9054);
nor U9355 (N_9355,N_9173,N_9072);
nor U9356 (N_9356,N_9181,N_9057);
or U9357 (N_9357,N_9131,N_9116);
or U9358 (N_9358,N_9008,N_9022);
nor U9359 (N_9359,N_9138,N_9044);
nand U9360 (N_9360,N_9101,N_9125);
nor U9361 (N_9361,N_9145,N_9065);
nor U9362 (N_9362,N_9080,N_9155);
and U9363 (N_9363,N_9073,N_9013);
and U9364 (N_9364,N_9117,N_9153);
or U9365 (N_9365,N_9092,N_9120);
or U9366 (N_9366,N_9103,N_9132);
and U9367 (N_9367,N_9136,N_9154);
and U9368 (N_9368,N_9044,N_9128);
nand U9369 (N_9369,N_9112,N_9124);
nand U9370 (N_9370,N_9004,N_9162);
and U9371 (N_9371,N_9118,N_9055);
and U9372 (N_9372,N_9122,N_9117);
nand U9373 (N_9373,N_9057,N_9176);
or U9374 (N_9374,N_9076,N_9074);
nand U9375 (N_9375,N_9191,N_9175);
and U9376 (N_9376,N_9153,N_9094);
nor U9377 (N_9377,N_9103,N_9021);
or U9378 (N_9378,N_9042,N_9150);
xnor U9379 (N_9379,N_9083,N_9110);
nand U9380 (N_9380,N_9181,N_9030);
and U9381 (N_9381,N_9032,N_9036);
xnor U9382 (N_9382,N_9127,N_9091);
or U9383 (N_9383,N_9012,N_9174);
nor U9384 (N_9384,N_9149,N_9123);
nand U9385 (N_9385,N_9028,N_9106);
nor U9386 (N_9386,N_9154,N_9059);
nor U9387 (N_9387,N_9014,N_9173);
and U9388 (N_9388,N_9000,N_9066);
or U9389 (N_9389,N_9024,N_9034);
nor U9390 (N_9390,N_9049,N_9043);
xnor U9391 (N_9391,N_9075,N_9014);
xnor U9392 (N_9392,N_9159,N_9077);
nand U9393 (N_9393,N_9020,N_9053);
nor U9394 (N_9394,N_9166,N_9131);
or U9395 (N_9395,N_9126,N_9059);
nand U9396 (N_9396,N_9168,N_9170);
nor U9397 (N_9397,N_9109,N_9172);
xnor U9398 (N_9398,N_9076,N_9124);
nand U9399 (N_9399,N_9120,N_9036);
xor U9400 (N_9400,N_9274,N_9331);
xor U9401 (N_9401,N_9302,N_9234);
and U9402 (N_9402,N_9367,N_9242);
or U9403 (N_9403,N_9324,N_9254);
xnor U9404 (N_9404,N_9230,N_9250);
and U9405 (N_9405,N_9259,N_9294);
and U9406 (N_9406,N_9384,N_9399);
nor U9407 (N_9407,N_9265,N_9396);
nor U9408 (N_9408,N_9239,N_9201);
xnor U9409 (N_9409,N_9363,N_9394);
or U9410 (N_9410,N_9269,N_9385);
xor U9411 (N_9411,N_9272,N_9372);
and U9412 (N_9412,N_9225,N_9317);
nand U9413 (N_9413,N_9296,N_9270);
and U9414 (N_9414,N_9267,N_9348);
and U9415 (N_9415,N_9316,N_9304);
xor U9416 (N_9416,N_9379,N_9223);
nor U9417 (N_9417,N_9214,N_9358);
xnor U9418 (N_9418,N_9361,N_9397);
xor U9419 (N_9419,N_9247,N_9387);
nand U9420 (N_9420,N_9307,N_9373);
nand U9421 (N_9421,N_9381,N_9325);
xnor U9422 (N_9422,N_9318,N_9392);
and U9423 (N_9423,N_9278,N_9374);
nand U9424 (N_9424,N_9208,N_9284);
nor U9425 (N_9425,N_9355,N_9389);
or U9426 (N_9426,N_9257,N_9268);
or U9427 (N_9427,N_9335,N_9398);
nor U9428 (N_9428,N_9292,N_9228);
nor U9429 (N_9429,N_9386,N_9341);
nor U9430 (N_9430,N_9283,N_9288);
nand U9431 (N_9431,N_9306,N_9333);
and U9432 (N_9432,N_9285,N_9376);
or U9433 (N_9433,N_9210,N_9320);
nor U9434 (N_9434,N_9298,N_9312);
nor U9435 (N_9435,N_9339,N_9258);
nand U9436 (N_9436,N_9291,N_9264);
or U9437 (N_9437,N_9319,N_9248);
xnor U9438 (N_9438,N_9351,N_9233);
or U9439 (N_9439,N_9226,N_9238);
xnor U9440 (N_9440,N_9327,N_9217);
and U9441 (N_9441,N_9219,N_9383);
nor U9442 (N_9442,N_9364,N_9299);
nand U9443 (N_9443,N_9357,N_9345);
or U9444 (N_9444,N_9368,N_9289);
or U9445 (N_9445,N_9220,N_9252);
and U9446 (N_9446,N_9260,N_9315);
and U9447 (N_9447,N_9300,N_9343);
nor U9448 (N_9448,N_9359,N_9277);
or U9449 (N_9449,N_9213,N_9303);
or U9450 (N_9450,N_9310,N_9309);
xor U9451 (N_9451,N_9236,N_9246);
xnor U9452 (N_9452,N_9311,N_9275);
nand U9453 (N_9453,N_9337,N_9243);
or U9454 (N_9454,N_9377,N_9271);
nor U9455 (N_9455,N_9273,N_9293);
or U9456 (N_9456,N_9360,N_9224);
and U9457 (N_9457,N_9338,N_9356);
or U9458 (N_9458,N_9349,N_9218);
nand U9459 (N_9459,N_9314,N_9366);
or U9460 (N_9460,N_9216,N_9221);
nand U9461 (N_9461,N_9342,N_9211);
xnor U9462 (N_9462,N_9207,N_9380);
or U9463 (N_9463,N_9346,N_9329);
nand U9464 (N_9464,N_9388,N_9227);
nor U9465 (N_9465,N_9229,N_9393);
nand U9466 (N_9466,N_9204,N_9261);
nor U9467 (N_9467,N_9305,N_9202);
nand U9468 (N_9468,N_9215,N_9352);
xnor U9469 (N_9469,N_9231,N_9321);
nand U9470 (N_9470,N_9256,N_9281);
nand U9471 (N_9471,N_9326,N_9232);
nand U9472 (N_9472,N_9370,N_9263);
nand U9473 (N_9473,N_9390,N_9301);
or U9474 (N_9474,N_9212,N_9336);
or U9475 (N_9475,N_9295,N_9245);
nor U9476 (N_9476,N_9313,N_9276);
or U9477 (N_9477,N_9235,N_9240);
nor U9478 (N_9478,N_9395,N_9369);
and U9479 (N_9479,N_9266,N_9244);
xor U9480 (N_9480,N_9222,N_9353);
nand U9481 (N_9481,N_9382,N_9262);
nor U9482 (N_9482,N_9290,N_9297);
or U9483 (N_9483,N_9209,N_9251);
nor U9484 (N_9484,N_9200,N_9347);
or U9485 (N_9485,N_9280,N_9241);
or U9486 (N_9486,N_9322,N_9332);
nor U9487 (N_9487,N_9350,N_9323);
and U9488 (N_9488,N_9279,N_9328);
nor U9489 (N_9489,N_9206,N_9308);
or U9490 (N_9490,N_9334,N_9282);
xnor U9491 (N_9491,N_9391,N_9330);
nand U9492 (N_9492,N_9340,N_9354);
nor U9493 (N_9493,N_9378,N_9365);
xnor U9494 (N_9494,N_9344,N_9287);
or U9495 (N_9495,N_9249,N_9286);
or U9496 (N_9496,N_9255,N_9253);
nand U9497 (N_9497,N_9362,N_9203);
xor U9498 (N_9498,N_9371,N_9237);
nor U9499 (N_9499,N_9205,N_9375);
and U9500 (N_9500,N_9237,N_9291);
and U9501 (N_9501,N_9376,N_9273);
or U9502 (N_9502,N_9366,N_9336);
and U9503 (N_9503,N_9236,N_9390);
nor U9504 (N_9504,N_9347,N_9310);
nor U9505 (N_9505,N_9325,N_9374);
nor U9506 (N_9506,N_9391,N_9398);
and U9507 (N_9507,N_9291,N_9261);
or U9508 (N_9508,N_9327,N_9310);
or U9509 (N_9509,N_9220,N_9333);
nand U9510 (N_9510,N_9262,N_9212);
and U9511 (N_9511,N_9335,N_9316);
nor U9512 (N_9512,N_9300,N_9295);
nor U9513 (N_9513,N_9311,N_9362);
or U9514 (N_9514,N_9270,N_9245);
or U9515 (N_9515,N_9307,N_9337);
nor U9516 (N_9516,N_9272,N_9341);
nor U9517 (N_9517,N_9285,N_9216);
or U9518 (N_9518,N_9311,N_9394);
and U9519 (N_9519,N_9253,N_9272);
or U9520 (N_9520,N_9239,N_9360);
nor U9521 (N_9521,N_9350,N_9211);
xor U9522 (N_9522,N_9321,N_9289);
xor U9523 (N_9523,N_9234,N_9379);
nand U9524 (N_9524,N_9245,N_9200);
or U9525 (N_9525,N_9356,N_9263);
or U9526 (N_9526,N_9385,N_9225);
nor U9527 (N_9527,N_9208,N_9392);
or U9528 (N_9528,N_9345,N_9361);
or U9529 (N_9529,N_9220,N_9315);
or U9530 (N_9530,N_9246,N_9324);
xnor U9531 (N_9531,N_9386,N_9336);
or U9532 (N_9532,N_9386,N_9211);
nor U9533 (N_9533,N_9324,N_9216);
nor U9534 (N_9534,N_9323,N_9340);
nor U9535 (N_9535,N_9345,N_9395);
and U9536 (N_9536,N_9246,N_9240);
nor U9537 (N_9537,N_9282,N_9386);
xnor U9538 (N_9538,N_9229,N_9295);
or U9539 (N_9539,N_9203,N_9279);
or U9540 (N_9540,N_9379,N_9215);
and U9541 (N_9541,N_9328,N_9315);
nor U9542 (N_9542,N_9254,N_9371);
and U9543 (N_9543,N_9245,N_9383);
nor U9544 (N_9544,N_9313,N_9241);
nand U9545 (N_9545,N_9213,N_9262);
nor U9546 (N_9546,N_9277,N_9236);
nand U9547 (N_9547,N_9317,N_9356);
and U9548 (N_9548,N_9373,N_9381);
nand U9549 (N_9549,N_9223,N_9397);
xor U9550 (N_9550,N_9367,N_9268);
xor U9551 (N_9551,N_9211,N_9205);
and U9552 (N_9552,N_9265,N_9235);
or U9553 (N_9553,N_9393,N_9352);
xnor U9554 (N_9554,N_9241,N_9333);
xnor U9555 (N_9555,N_9293,N_9263);
nand U9556 (N_9556,N_9394,N_9238);
xnor U9557 (N_9557,N_9228,N_9207);
nand U9558 (N_9558,N_9243,N_9371);
nor U9559 (N_9559,N_9347,N_9357);
nand U9560 (N_9560,N_9297,N_9398);
nand U9561 (N_9561,N_9298,N_9279);
or U9562 (N_9562,N_9240,N_9223);
xor U9563 (N_9563,N_9217,N_9281);
or U9564 (N_9564,N_9399,N_9233);
and U9565 (N_9565,N_9302,N_9372);
nand U9566 (N_9566,N_9249,N_9243);
nor U9567 (N_9567,N_9342,N_9271);
nor U9568 (N_9568,N_9211,N_9225);
nor U9569 (N_9569,N_9270,N_9343);
or U9570 (N_9570,N_9238,N_9254);
or U9571 (N_9571,N_9314,N_9273);
nand U9572 (N_9572,N_9218,N_9261);
xor U9573 (N_9573,N_9220,N_9399);
or U9574 (N_9574,N_9242,N_9380);
nand U9575 (N_9575,N_9294,N_9265);
xor U9576 (N_9576,N_9321,N_9369);
or U9577 (N_9577,N_9310,N_9257);
nor U9578 (N_9578,N_9319,N_9370);
xor U9579 (N_9579,N_9233,N_9264);
nor U9580 (N_9580,N_9371,N_9353);
xor U9581 (N_9581,N_9262,N_9366);
nand U9582 (N_9582,N_9328,N_9332);
and U9583 (N_9583,N_9283,N_9209);
nand U9584 (N_9584,N_9357,N_9231);
nor U9585 (N_9585,N_9332,N_9275);
nor U9586 (N_9586,N_9281,N_9201);
or U9587 (N_9587,N_9282,N_9244);
and U9588 (N_9588,N_9211,N_9308);
nor U9589 (N_9589,N_9342,N_9322);
xnor U9590 (N_9590,N_9241,N_9210);
nand U9591 (N_9591,N_9278,N_9259);
nand U9592 (N_9592,N_9237,N_9350);
and U9593 (N_9593,N_9326,N_9322);
and U9594 (N_9594,N_9385,N_9214);
and U9595 (N_9595,N_9201,N_9358);
or U9596 (N_9596,N_9357,N_9211);
nand U9597 (N_9597,N_9317,N_9224);
or U9598 (N_9598,N_9378,N_9360);
and U9599 (N_9599,N_9222,N_9339);
nor U9600 (N_9600,N_9446,N_9421);
nor U9601 (N_9601,N_9416,N_9538);
nand U9602 (N_9602,N_9408,N_9597);
xnor U9603 (N_9603,N_9546,N_9482);
xor U9604 (N_9604,N_9519,N_9447);
and U9605 (N_9605,N_9543,N_9526);
xnor U9606 (N_9606,N_9427,N_9590);
or U9607 (N_9607,N_9593,N_9485);
xor U9608 (N_9608,N_9440,N_9414);
and U9609 (N_9609,N_9400,N_9545);
and U9610 (N_9610,N_9551,N_9566);
nor U9611 (N_9611,N_9452,N_9514);
nand U9612 (N_9612,N_9422,N_9418);
nor U9613 (N_9613,N_9415,N_9419);
and U9614 (N_9614,N_9495,N_9588);
nand U9615 (N_9615,N_9560,N_9402);
xnor U9616 (N_9616,N_9576,N_9473);
and U9617 (N_9617,N_9476,N_9556);
nor U9618 (N_9618,N_9437,N_9504);
nor U9619 (N_9619,N_9596,N_9497);
xnor U9620 (N_9620,N_9413,N_9466);
and U9621 (N_9621,N_9570,N_9405);
nand U9622 (N_9622,N_9487,N_9434);
or U9623 (N_9623,N_9537,N_9587);
or U9624 (N_9624,N_9586,N_9534);
nor U9625 (N_9625,N_9459,N_9591);
nand U9626 (N_9626,N_9594,N_9449);
xor U9627 (N_9627,N_9502,N_9505);
or U9628 (N_9628,N_9598,N_9554);
xor U9629 (N_9629,N_9469,N_9571);
and U9630 (N_9630,N_9508,N_9544);
and U9631 (N_9631,N_9595,N_9532);
nand U9632 (N_9632,N_9577,N_9444);
nand U9633 (N_9633,N_9456,N_9409);
nor U9634 (N_9634,N_9585,N_9484);
xnor U9635 (N_9635,N_9455,N_9489);
nor U9636 (N_9636,N_9483,N_9461);
or U9637 (N_9637,N_9531,N_9478);
nor U9638 (N_9638,N_9525,N_9507);
nor U9639 (N_9639,N_9499,N_9488);
and U9640 (N_9640,N_9559,N_9511);
xor U9641 (N_9641,N_9486,N_9548);
xor U9642 (N_9642,N_9438,N_9510);
nand U9643 (N_9643,N_9472,N_9540);
or U9644 (N_9644,N_9549,N_9501);
nand U9645 (N_9645,N_9578,N_9480);
xor U9646 (N_9646,N_9442,N_9599);
nand U9647 (N_9647,N_9411,N_9584);
or U9648 (N_9648,N_9443,N_9536);
xnor U9649 (N_9649,N_9517,N_9404);
xnor U9650 (N_9650,N_9568,N_9521);
and U9651 (N_9651,N_9417,N_9403);
and U9652 (N_9652,N_9454,N_9462);
xnor U9653 (N_9653,N_9445,N_9474);
nor U9654 (N_9654,N_9569,N_9516);
or U9655 (N_9655,N_9428,N_9439);
and U9656 (N_9656,N_9471,N_9581);
xor U9657 (N_9657,N_9492,N_9406);
and U9658 (N_9658,N_9432,N_9458);
nor U9659 (N_9659,N_9436,N_9592);
nor U9660 (N_9660,N_9574,N_9564);
nor U9661 (N_9661,N_9448,N_9523);
nand U9662 (N_9662,N_9522,N_9460);
xor U9663 (N_9663,N_9496,N_9457);
nand U9664 (N_9664,N_9425,N_9431);
and U9665 (N_9665,N_9450,N_9401);
or U9666 (N_9666,N_9407,N_9557);
xnor U9667 (N_9667,N_9552,N_9430);
nand U9668 (N_9668,N_9493,N_9481);
and U9669 (N_9669,N_9589,N_9524);
and U9670 (N_9670,N_9435,N_9561);
and U9671 (N_9671,N_9558,N_9498);
and U9672 (N_9672,N_9451,N_9542);
nor U9673 (N_9673,N_9470,N_9467);
or U9674 (N_9674,N_9465,N_9506);
and U9675 (N_9675,N_9494,N_9580);
xor U9676 (N_9676,N_9475,N_9520);
nand U9677 (N_9677,N_9572,N_9553);
nor U9678 (N_9678,N_9528,N_9565);
or U9679 (N_9679,N_9575,N_9412);
nor U9680 (N_9680,N_9420,N_9562);
and U9681 (N_9681,N_9463,N_9563);
or U9682 (N_9682,N_9530,N_9433);
xor U9683 (N_9683,N_9426,N_9555);
or U9684 (N_9684,N_9464,N_9509);
or U9685 (N_9685,N_9477,N_9500);
nand U9686 (N_9686,N_9518,N_9513);
and U9687 (N_9687,N_9567,N_9490);
xor U9688 (N_9688,N_9429,N_9503);
nand U9689 (N_9689,N_9535,N_9491);
xor U9690 (N_9690,N_9515,N_9547);
xor U9691 (N_9691,N_9468,N_9512);
xor U9692 (N_9692,N_9410,N_9550);
xnor U9693 (N_9693,N_9527,N_9424);
nand U9694 (N_9694,N_9539,N_9479);
and U9695 (N_9695,N_9423,N_9533);
nor U9696 (N_9696,N_9579,N_9453);
xnor U9697 (N_9697,N_9583,N_9573);
nor U9698 (N_9698,N_9541,N_9441);
xor U9699 (N_9699,N_9582,N_9529);
or U9700 (N_9700,N_9453,N_9473);
xnor U9701 (N_9701,N_9529,N_9574);
nand U9702 (N_9702,N_9426,N_9560);
xor U9703 (N_9703,N_9523,N_9556);
or U9704 (N_9704,N_9401,N_9530);
nor U9705 (N_9705,N_9554,N_9501);
or U9706 (N_9706,N_9462,N_9439);
and U9707 (N_9707,N_9454,N_9505);
or U9708 (N_9708,N_9414,N_9450);
nor U9709 (N_9709,N_9499,N_9456);
or U9710 (N_9710,N_9488,N_9538);
and U9711 (N_9711,N_9563,N_9565);
nor U9712 (N_9712,N_9508,N_9459);
and U9713 (N_9713,N_9460,N_9583);
and U9714 (N_9714,N_9507,N_9429);
or U9715 (N_9715,N_9587,N_9434);
nand U9716 (N_9716,N_9556,N_9535);
and U9717 (N_9717,N_9450,N_9531);
or U9718 (N_9718,N_9496,N_9487);
nand U9719 (N_9719,N_9492,N_9481);
xnor U9720 (N_9720,N_9403,N_9455);
or U9721 (N_9721,N_9496,N_9505);
xor U9722 (N_9722,N_9525,N_9414);
and U9723 (N_9723,N_9430,N_9428);
nand U9724 (N_9724,N_9423,N_9583);
nor U9725 (N_9725,N_9517,N_9565);
or U9726 (N_9726,N_9581,N_9504);
xnor U9727 (N_9727,N_9535,N_9504);
nor U9728 (N_9728,N_9536,N_9555);
and U9729 (N_9729,N_9482,N_9443);
and U9730 (N_9730,N_9578,N_9452);
nand U9731 (N_9731,N_9484,N_9532);
nand U9732 (N_9732,N_9451,N_9587);
xnor U9733 (N_9733,N_9488,N_9551);
nand U9734 (N_9734,N_9527,N_9500);
nand U9735 (N_9735,N_9445,N_9488);
nor U9736 (N_9736,N_9476,N_9483);
and U9737 (N_9737,N_9555,N_9497);
xor U9738 (N_9738,N_9519,N_9524);
or U9739 (N_9739,N_9566,N_9422);
or U9740 (N_9740,N_9576,N_9423);
nor U9741 (N_9741,N_9536,N_9541);
nand U9742 (N_9742,N_9415,N_9527);
xor U9743 (N_9743,N_9529,N_9539);
or U9744 (N_9744,N_9442,N_9592);
nor U9745 (N_9745,N_9567,N_9478);
nand U9746 (N_9746,N_9443,N_9450);
nor U9747 (N_9747,N_9553,N_9411);
nand U9748 (N_9748,N_9432,N_9461);
and U9749 (N_9749,N_9580,N_9482);
or U9750 (N_9750,N_9594,N_9559);
and U9751 (N_9751,N_9412,N_9567);
and U9752 (N_9752,N_9406,N_9434);
xor U9753 (N_9753,N_9419,N_9406);
nand U9754 (N_9754,N_9431,N_9474);
nand U9755 (N_9755,N_9429,N_9471);
or U9756 (N_9756,N_9451,N_9447);
xor U9757 (N_9757,N_9514,N_9588);
nor U9758 (N_9758,N_9474,N_9450);
nand U9759 (N_9759,N_9594,N_9499);
and U9760 (N_9760,N_9412,N_9440);
and U9761 (N_9761,N_9520,N_9511);
xor U9762 (N_9762,N_9546,N_9424);
nand U9763 (N_9763,N_9444,N_9459);
or U9764 (N_9764,N_9430,N_9544);
xnor U9765 (N_9765,N_9446,N_9408);
and U9766 (N_9766,N_9583,N_9448);
nor U9767 (N_9767,N_9596,N_9403);
nor U9768 (N_9768,N_9509,N_9588);
xor U9769 (N_9769,N_9497,N_9583);
nand U9770 (N_9770,N_9466,N_9592);
nand U9771 (N_9771,N_9502,N_9442);
and U9772 (N_9772,N_9505,N_9463);
or U9773 (N_9773,N_9537,N_9516);
nand U9774 (N_9774,N_9594,N_9526);
xor U9775 (N_9775,N_9501,N_9564);
nor U9776 (N_9776,N_9441,N_9533);
xor U9777 (N_9777,N_9596,N_9511);
nand U9778 (N_9778,N_9595,N_9410);
xor U9779 (N_9779,N_9526,N_9430);
and U9780 (N_9780,N_9423,N_9549);
xor U9781 (N_9781,N_9500,N_9441);
nor U9782 (N_9782,N_9578,N_9515);
and U9783 (N_9783,N_9559,N_9437);
nand U9784 (N_9784,N_9413,N_9550);
nor U9785 (N_9785,N_9574,N_9442);
nand U9786 (N_9786,N_9410,N_9594);
nand U9787 (N_9787,N_9472,N_9421);
or U9788 (N_9788,N_9406,N_9545);
or U9789 (N_9789,N_9425,N_9454);
xnor U9790 (N_9790,N_9400,N_9527);
and U9791 (N_9791,N_9473,N_9401);
xor U9792 (N_9792,N_9475,N_9563);
and U9793 (N_9793,N_9439,N_9515);
xor U9794 (N_9794,N_9404,N_9470);
nor U9795 (N_9795,N_9424,N_9418);
and U9796 (N_9796,N_9450,N_9405);
nor U9797 (N_9797,N_9446,N_9471);
nor U9798 (N_9798,N_9429,N_9418);
and U9799 (N_9799,N_9498,N_9497);
and U9800 (N_9800,N_9688,N_9670);
nand U9801 (N_9801,N_9634,N_9636);
xnor U9802 (N_9802,N_9727,N_9739);
xor U9803 (N_9803,N_9775,N_9686);
and U9804 (N_9804,N_9612,N_9735);
nor U9805 (N_9805,N_9678,N_9745);
xor U9806 (N_9806,N_9650,N_9667);
xor U9807 (N_9807,N_9681,N_9607);
nor U9808 (N_9808,N_9608,N_9647);
xnor U9809 (N_9809,N_9764,N_9654);
and U9810 (N_9810,N_9716,N_9763);
xnor U9811 (N_9811,N_9628,N_9731);
xor U9812 (N_9812,N_9640,N_9722);
nor U9813 (N_9813,N_9777,N_9749);
nand U9814 (N_9814,N_9637,N_9776);
and U9815 (N_9815,N_9684,N_9736);
or U9816 (N_9816,N_9699,N_9672);
nor U9817 (N_9817,N_9798,N_9754);
nor U9818 (N_9818,N_9632,N_9700);
xnor U9819 (N_9819,N_9767,N_9796);
nor U9820 (N_9820,N_9741,N_9685);
or U9821 (N_9821,N_9664,N_9631);
xnor U9822 (N_9822,N_9698,N_9615);
nor U9823 (N_9823,N_9617,N_9778);
nor U9824 (N_9824,N_9750,N_9605);
or U9825 (N_9825,N_9641,N_9768);
nand U9826 (N_9826,N_9740,N_9758);
nor U9827 (N_9827,N_9712,N_9620);
or U9828 (N_9828,N_9600,N_9680);
nor U9829 (N_9829,N_9705,N_9765);
nor U9830 (N_9830,N_9694,N_9610);
nor U9831 (N_9831,N_9662,N_9773);
xnor U9832 (N_9832,N_9625,N_9645);
nand U9833 (N_9833,N_9623,N_9665);
xor U9834 (N_9834,N_9709,N_9788);
and U9835 (N_9835,N_9744,N_9791);
nand U9836 (N_9836,N_9674,N_9639);
or U9837 (N_9837,N_9710,N_9762);
or U9838 (N_9838,N_9683,N_9718);
nand U9839 (N_9839,N_9633,N_9785);
nor U9840 (N_9840,N_9792,N_9748);
or U9841 (N_9841,N_9757,N_9751);
and U9842 (N_9842,N_9738,N_9687);
xnor U9843 (N_9843,N_9653,N_9626);
xnor U9844 (N_9844,N_9658,N_9769);
and U9845 (N_9845,N_9734,N_9659);
xnor U9846 (N_9846,N_9782,N_9780);
or U9847 (N_9847,N_9614,N_9787);
nand U9848 (N_9848,N_9714,N_9789);
nand U9849 (N_9849,N_9675,N_9717);
and U9850 (N_9850,N_9635,N_9725);
xor U9851 (N_9851,N_9690,N_9649);
xnor U9852 (N_9852,N_9799,N_9661);
xnor U9853 (N_9853,N_9630,N_9794);
or U9854 (N_9854,N_9697,N_9756);
nor U9855 (N_9855,N_9779,N_9793);
nor U9856 (N_9856,N_9715,N_9668);
or U9857 (N_9857,N_9618,N_9703);
nor U9858 (N_9858,N_9604,N_9646);
xnor U9859 (N_9859,N_9644,N_9719);
nor U9860 (N_9860,N_9629,N_9676);
xor U9861 (N_9861,N_9651,N_9797);
and U9862 (N_9862,N_9622,N_9656);
xor U9863 (N_9863,N_9708,N_9729);
nor U9864 (N_9864,N_9746,N_9781);
and U9865 (N_9865,N_9648,N_9737);
or U9866 (N_9866,N_9755,N_9742);
or U9867 (N_9867,N_9603,N_9673);
xor U9868 (N_9868,N_9652,N_9624);
xor U9869 (N_9869,N_9795,N_9692);
nand U9870 (N_9870,N_9702,N_9772);
xor U9871 (N_9871,N_9677,N_9753);
or U9872 (N_9872,N_9611,N_9691);
or U9873 (N_9873,N_9761,N_9730);
nand U9874 (N_9874,N_9627,N_9657);
nand U9875 (N_9875,N_9752,N_9783);
nor U9876 (N_9876,N_9726,N_9696);
xnor U9877 (N_9877,N_9771,N_9679);
and U9878 (N_9878,N_9760,N_9619);
and U9879 (N_9879,N_9682,N_9669);
and U9880 (N_9880,N_9671,N_9606);
and U9881 (N_9881,N_9663,N_9786);
nand U9882 (N_9882,N_9720,N_9643);
or U9883 (N_9883,N_9609,N_9602);
and U9884 (N_9884,N_9747,N_9723);
or U9885 (N_9885,N_9732,N_9613);
xnor U9886 (N_9886,N_9733,N_9784);
xnor U9887 (N_9887,N_9689,N_9695);
and U9888 (N_9888,N_9655,N_9770);
or U9889 (N_9889,N_9766,N_9701);
nor U9890 (N_9890,N_9711,N_9660);
nand U9891 (N_9891,N_9790,N_9616);
xnor U9892 (N_9892,N_9706,N_9774);
or U9893 (N_9893,N_9713,N_9642);
or U9894 (N_9894,N_9743,N_9728);
nand U9895 (N_9895,N_9704,N_9693);
xnor U9896 (N_9896,N_9724,N_9666);
nand U9897 (N_9897,N_9707,N_9759);
xor U9898 (N_9898,N_9601,N_9621);
nand U9899 (N_9899,N_9638,N_9721);
nor U9900 (N_9900,N_9766,N_9780);
xnor U9901 (N_9901,N_9678,N_9795);
nor U9902 (N_9902,N_9627,N_9702);
nor U9903 (N_9903,N_9785,N_9721);
xor U9904 (N_9904,N_9673,N_9662);
nor U9905 (N_9905,N_9704,N_9797);
nand U9906 (N_9906,N_9662,N_9653);
and U9907 (N_9907,N_9765,N_9759);
and U9908 (N_9908,N_9737,N_9707);
or U9909 (N_9909,N_9760,N_9798);
and U9910 (N_9910,N_9603,N_9667);
nand U9911 (N_9911,N_9613,N_9713);
or U9912 (N_9912,N_9644,N_9656);
and U9913 (N_9913,N_9742,N_9623);
nand U9914 (N_9914,N_9707,N_9718);
nor U9915 (N_9915,N_9709,N_9785);
or U9916 (N_9916,N_9677,N_9638);
xnor U9917 (N_9917,N_9684,N_9738);
nand U9918 (N_9918,N_9757,N_9708);
and U9919 (N_9919,N_9722,N_9653);
xnor U9920 (N_9920,N_9795,N_9710);
nand U9921 (N_9921,N_9690,N_9656);
nor U9922 (N_9922,N_9685,N_9659);
or U9923 (N_9923,N_9708,N_9675);
xor U9924 (N_9924,N_9696,N_9743);
or U9925 (N_9925,N_9696,N_9722);
and U9926 (N_9926,N_9743,N_9753);
nand U9927 (N_9927,N_9698,N_9601);
and U9928 (N_9928,N_9729,N_9650);
nor U9929 (N_9929,N_9716,N_9700);
xnor U9930 (N_9930,N_9654,N_9708);
nand U9931 (N_9931,N_9648,N_9641);
nand U9932 (N_9932,N_9773,N_9768);
xor U9933 (N_9933,N_9760,N_9736);
and U9934 (N_9934,N_9682,N_9708);
nand U9935 (N_9935,N_9690,N_9630);
xor U9936 (N_9936,N_9756,N_9630);
or U9937 (N_9937,N_9750,N_9742);
xnor U9938 (N_9938,N_9778,N_9688);
and U9939 (N_9939,N_9636,N_9790);
or U9940 (N_9940,N_9657,N_9684);
nor U9941 (N_9941,N_9767,N_9712);
or U9942 (N_9942,N_9691,N_9629);
xor U9943 (N_9943,N_9681,N_9639);
xnor U9944 (N_9944,N_9705,N_9618);
nand U9945 (N_9945,N_9772,N_9725);
xnor U9946 (N_9946,N_9787,N_9678);
nand U9947 (N_9947,N_9612,N_9770);
nor U9948 (N_9948,N_9771,N_9668);
or U9949 (N_9949,N_9656,N_9724);
and U9950 (N_9950,N_9637,N_9614);
nor U9951 (N_9951,N_9682,N_9703);
xnor U9952 (N_9952,N_9611,N_9747);
and U9953 (N_9953,N_9757,N_9707);
and U9954 (N_9954,N_9733,N_9731);
or U9955 (N_9955,N_9681,N_9694);
nor U9956 (N_9956,N_9615,N_9749);
and U9957 (N_9957,N_9719,N_9720);
and U9958 (N_9958,N_9779,N_9667);
and U9959 (N_9959,N_9690,N_9741);
nor U9960 (N_9960,N_9647,N_9654);
nor U9961 (N_9961,N_9755,N_9665);
and U9962 (N_9962,N_9778,N_9783);
or U9963 (N_9963,N_9676,N_9734);
or U9964 (N_9964,N_9666,N_9639);
xor U9965 (N_9965,N_9616,N_9655);
or U9966 (N_9966,N_9685,N_9629);
nand U9967 (N_9967,N_9786,N_9648);
nand U9968 (N_9968,N_9756,N_9775);
nand U9969 (N_9969,N_9729,N_9763);
nand U9970 (N_9970,N_9799,N_9664);
and U9971 (N_9971,N_9727,N_9635);
or U9972 (N_9972,N_9659,N_9704);
nand U9973 (N_9973,N_9785,N_9692);
or U9974 (N_9974,N_9791,N_9611);
and U9975 (N_9975,N_9690,N_9786);
nand U9976 (N_9976,N_9718,N_9744);
nor U9977 (N_9977,N_9757,N_9684);
or U9978 (N_9978,N_9649,N_9729);
or U9979 (N_9979,N_9678,N_9749);
and U9980 (N_9980,N_9734,N_9632);
nand U9981 (N_9981,N_9759,N_9703);
nand U9982 (N_9982,N_9678,N_9798);
nor U9983 (N_9983,N_9796,N_9682);
nor U9984 (N_9984,N_9687,N_9795);
nor U9985 (N_9985,N_9756,N_9668);
nor U9986 (N_9986,N_9689,N_9741);
or U9987 (N_9987,N_9715,N_9684);
and U9988 (N_9988,N_9608,N_9719);
and U9989 (N_9989,N_9744,N_9724);
and U9990 (N_9990,N_9681,N_9612);
or U9991 (N_9991,N_9711,N_9747);
or U9992 (N_9992,N_9675,N_9728);
nor U9993 (N_9993,N_9611,N_9740);
and U9994 (N_9994,N_9620,N_9680);
nor U9995 (N_9995,N_9724,N_9732);
xor U9996 (N_9996,N_9626,N_9688);
nand U9997 (N_9997,N_9738,N_9637);
or U9998 (N_9998,N_9747,N_9674);
nor U9999 (N_9999,N_9626,N_9780);
nand U10000 (N_10000,N_9833,N_9985);
or U10001 (N_10001,N_9821,N_9955);
or U10002 (N_10002,N_9855,N_9818);
nor U10003 (N_10003,N_9824,N_9811);
or U10004 (N_10004,N_9988,N_9822);
and U10005 (N_10005,N_9928,N_9970);
and U10006 (N_10006,N_9838,N_9954);
xnor U10007 (N_10007,N_9974,N_9914);
nor U10008 (N_10008,N_9925,N_9885);
and U10009 (N_10009,N_9829,N_9981);
nor U10010 (N_10010,N_9860,N_9912);
nand U10011 (N_10011,N_9964,N_9979);
and U10012 (N_10012,N_9962,N_9938);
nor U10013 (N_10013,N_9966,N_9908);
nand U10014 (N_10014,N_9987,N_9997);
or U10015 (N_10015,N_9924,N_9884);
and U10016 (N_10016,N_9982,N_9871);
xnor U10017 (N_10017,N_9853,N_9913);
nand U10018 (N_10018,N_9986,N_9959);
nor U10019 (N_10019,N_9946,N_9990);
and U10020 (N_10020,N_9900,N_9907);
and U10021 (N_10021,N_9933,N_9803);
nand U10022 (N_10022,N_9842,N_9800);
nor U10023 (N_10023,N_9841,N_9866);
nand U10024 (N_10024,N_9864,N_9875);
nand U10025 (N_10025,N_9832,N_9975);
nand U10026 (N_10026,N_9854,N_9816);
or U10027 (N_10027,N_9950,N_9968);
xor U10028 (N_10028,N_9919,N_9857);
nand U10029 (N_10029,N_9993,N_9805);
or U10030 (N_10030,N_9813,N_9906);
xor U10031 (N_10031,N_9936,N_9939);
or U10032 (N_10032,N_9980,N_9889);
nor U10033 (N_10033,N_9953,N_9899);
nor U10034 (N_10034,N_9896,N_9848);
or U10035 (N_10035,N_9940,N_9886);
nor U10036 (N_10036,N_9807,N_9969);
xor U10037 (N_10037,N_9991,N_9870);
xor U10038 (N_10038,N_9934,N_9910);
and U10039 (N_10039,N_9835,N_9941);
xnor U10040 (N_10040,N_9909,N_9817);
nor U10041 (N_10041,N_9911,N_9892);
and U10042 (N_10042,N_9883,N_9869);
nor U10043 (N_10043,N_9947,N_9808);
xor U10044 (N_10044,N_9978,N_9830);
nor U10045 (N_10045,N_9876,N_9996);
nand U10046 (N_10046,N_9961,N_9897);
nand U10047 (N_10047,N_9998,N_9823);
nor U10048 (N_10048,N_9944,N_9918);
nor U10049 (N_10049,N_9927,N_9880);
or U10050 (N_10050,N_9867,N_9862);
and U10051 (N_10051,N_9949,N_9951);
nor U10052 (N_10052,N_9917,N_9973);
and U10053 (N_10053,N_9844,N_9921);
nand U10054 (N_10054,N_9971,N_9868);
nand U10055 (N_10055,N_9815,N_9904);
nand U10056 (N_10056,N_9846,N_9967);
nor U10057 (N_10057,N_9812,N_9804);
or U10058 (N_10058,N_9992,N_9887);
xnor U10059 (N_10059,N_9849,N_9852);
nand U10060 (N_10060,N_9827,N_9888);
nand U10061 (N_10061,N_9895,N_9810);
xnor U10062 (N_10062,N_9859,N_9916);
and U10063 (N_10063,N_9882,N_9814);
nor U10064 (N_10064,N_9977,N_9929);
or U10065 (N_10065,N_9836,N_9865);
nand U10066 (N_10066,N_9999,N_9843);
nor U10067 (N_10067,N_9972,N_9920);
xor U10068 (N_10068,N_9948,N_9893);
and U10069 (N_10069,N_9994,N_9930);
and U10070 (N_10070,N_9922,N_9989);
and U10071 (N_10071,N_9881,N_9845);
nor U10072 (N_10072,N_9861,N_9801);
xnor U10073 (N_10073,N_9809,N_9945);
nand U10074 (N_10074,N_9856,N_9965);
and U10075 (N_10075,N_9976,N_9963);
nand U10076 (N_10076,N_9958,N_9937);
nor U10077 (N_10077,N_9890,N_9995);
or U10078 (N_10078,N_9831,N_9863);
and U10079 (N_10079,N_9879,N_9834);
nand U10080 (N_10080,N_9903,N_9905);
nor U10081 (N_10081,N_9931,N_9942);
xnor U10082 (N_10082,N_9837,N_9874);
and U10083 (N_10083,N_9901,N_9872);
and U10084 (N_10084,N_9935,N_9902);
nand U10085 (N_10085,N_9873,N_9957);
or U10086 (N_10086,N_9983,N_9851);
xnor U10087 (N_10087,N_9894,N_9926);
nor U10088 (N_10088,N_9819,N_9932);
and U10089 (N_10089,N_9915,N_9877);
or U10090 (N_10090,N_9923,N_9984);
and U10091 (N_10091,N_9802,N_9898);
or U10092 (N_10092,N_9943,N_9956);
nand U10093 (N_10093,N_9826,N_9847);
and U10094 (N_10094,N_9878,N_9806);
nor U10095 (N_10095,N_9840,N_9825);
and U10096 (N_10096,N_9839,N_9820);
nand U10097 (N_10097,N_9850,N_9960);
nor U10098 (N_10098,N_9828,N_9858);
nor U10099 (N_10099,N_9952,N_9891);
nor U10100 (N_10100,N_9978,N_9836);
nand U10101 (N_10101,N_9992,N_9849);
xnor U10102 (N_10102,N_9905,N_9837);
xor U10103 (N_10103,N_9883,N_9921);
nand U10104 (N_10104,N_9961,N_9902);
and U10105 (N_10105,N_9961,N_9899);
nand U10106 (N_10106,N_9806,N_9866);
xor U10107 (N_10107,N_9985,N_9959);
and U10108 (N_10108,N_9972,N_9851);
or U10109 (N_10109,N_9844,N_9857);
nand U10110 (N_10110,N_9876,N_9806);
nand U10111 (N_10111,N_9868,N_9922);
and U10112 (N_10112,N_9918,N_9900);
or U10113 (N_10113,N_9855,N_9877);
nor U10114 (N_10114,N_9996,N_9968);
nor U10115 (N_10115,N_9879,N_9997);
and U10116 (N_10116,N_9905,N_9860);
nand U10117 (N_10117,N_9904,N_9901);
xor U10118 (N_10118,N_9991,N_9886);
and U10119 (N_10119,N_9924,N_9849);
nand U10120 (N_10120,N_9900,N_9849);
nand U10121 (N_10121,N_9976,N_9827);
or U10122 (N_10122,N_9812,N_9970);
xor U10123 (N_10123,N_9914,N_9800);
nand U10124 (N_10124,N_9986,N_9873);
or U10125 (N_10125,N_9843,N_9844);
and U10126 (N_10126,N_9828,N_9814);
xor U10127 (N_10127,N_9893,N_9927);
xor U10128 (N_10128,N_9837,N_9818);
xor U10129 (N_10129,N_9867,N_9877);
or U10130 (N_10130,N_9982,N_9934);
nand U10131 (N_10131,N_9967,N_9912);
or U10132 (N_10132,N_9909,N_9982);
nor U10133 (N_10133,N_9890,N_9804);
nor U10134 (N_10134,N_9834,N_9886);
xor U10135 (N_10135,N_9947,N_9806);
xnor U10136 (N_10136,N_9989,N_9841);
and U10137 (N_10137,N_9833,N_9883);
or U10138 (N_10138,N_9964,N_9839);
and U10139 (N_10139,N_9836,N_9820);
nor U10140 (N_10140,N_9816,N_9814);
xor U10141 (N_10141,N_9858,N_9919);
nand U10142 (N_10142,N_9831,N_9994);
xnor U10143 (N_10143,N_9852,N_9954);
nand U10144 (N_10144,N_9880,N_9980);
nor U10145 (N_10145,N_9957,N_9931);
and U10146 (N_10146,N_9804,N_9990);
nand U10147 (N_10147,N_9939,N_9980);
nor U10148 (N_10148,N_9988,N_9969);
nor U10149 (N_10149,N_9948,N_9821);
and U10150 (N_10150,N_9879,N_9981);
and U10151 (N_10151,N_9827,N_9823);
and U10152 (N_10152,N_9907,N_9940);
nand U10153 (N_10153,N_9920,N_9852);
nand U10154 (N_10154,N_9908,N_9871);
nor U10155 (N_10155,N_9901,N_9819);
or U10156 (N_10156,N_9865,N_9980);
xnor U10157 (N_10157,N_9805,N_9907);
xnor U10158 (N_10158,N_9985,N_9963);
xnor U10159 (N_10159,N_9962,N_9932);
nand U10160 (N_10160,N_9948,N_9808);
xnor U10161 (N_10161,N_9954,N_9951);
xor U10162 (N_10162,N_9965,N_9828);
nor U10163 (N_10163,N_9924,N_9843);
xor U10164 (N_10164,N_9887,N_9828);
and U10165 (N_10165,N_9883,N_9931);
nand U10166 (N_10166,N_9919,N_9881);
nand U10167 (N_10167,N_9920,N_9943);
and U10168 (N_10168,N_9961,N_9819);
nor U10169 (N_10169,N_9879,N_9957);
nand U10170 (N_10170,N_9835,N_9976);
or U10171 (N_10171,N_9858,N_9988);
nor U10172 (N_10172,N_9967,N_9830);
or U10173 (N_10173,N_9922,N_9885);
xor U10174 (N_10174,N_9942,N_9824);
xnor U10175 (N_10175,N_9967,N_9954);
xnor U10176 (N_10176,N_9802,N_9953);
and U10177 (N_10177,N_9923,N_9960);
or U10178 (N_10178,N_9817,N_9834);
or U10179 (N_10179,N_9968,N_9862);
and U10180 (N_10180,N_9950,N_9826);
xor U10181 (N_10181,N_9865,N_9921);
xor U10182 (N_10182,N_9846,N_9976);
or U10183 (N_10183,N_9858,N_9935);
nor U10184 (N_10184,N_9889,N_9916);
and U10185 (N_10185,N_9971,N_9837);
or U10186 (N_10186,N_9911,N_9917);
and U10187 (N_10187,N_9978,N_9957);
xnor U10188 (N_10188,N_9965,N_9986);
nor U10189 (N_10189,N_9942,N_9974);
xor U10190 (N_10190,N_9857,N_9870);
or U10191 (N_10191,N_9878,N_9812);
xor U10192 (N_10192,N_9882,N_9830);
nand U10193 (N_10193,N_9801,N_9832);
or U10194 (N_10194,N_9897,N_9954);
xor U10195 (N_10195,N_9903,N_9954);
nand U10196 (N_10196,N_9898,N_9924);
or U10197 (N_10197,N_9874,N_9813);
or U10198 (N_10198,N_9961,N_9841);
nor U10199 (N_10199,N_9861,N_9899);
nand U10200 (N_10200,N_10055,N_10023);
or U10201 (N_10201,N_10065,N_10025);
nand U10202 (N_10202,N_10045,N_10111);
and U10203 (N_10203,N_10004,N_10140);
and U10204 (N_10204,N_10096,N_10020);
nor U10205 (N_10205,N_10048,N_10156);
xnor U10206 (N_10206,N_10099,N_10176);
xnor U10207 (N_10207,N_10181,N_10087);
xnor U10208 (N_10208,N_10119,N_10137);
nand U10209 (N_10209,N_10159,N_10038);
or U10210 (N_10210,N_10194,N_10064);
nor U10211 (N_10211,N_10125,N_10115);
nor U10212 (N_10212,N_10017,N_10146);
and U10213 (N_10213,N_10067,N_10081);
and U10214 (N_10214,N_10129,N_10030);
xnor U10215 (N_10215,N_10161,N_10006);
xnor U10216 (N_10216,N_10121,N_10116);
xnor U10217 (N_10217,N_10080,N_10155);
nand U10218 (N_10218,N_10012,N_10027);
or U10219 (N_10219,N_10084,N_10154);
and U10220 (N_10220,N_10082,N_10110);
or U10221 (N_10221,N_10092,N_10132);
nor U10222 (N_10222,N_10097,N_10160);
nor U10223 (N_10223,N_10001,N_10056);
nor U10224 (N_10224,N_10089,N_10197);
nor U10225 (N_10225,N_10144,N_10033);
nand U10226 (N_10226,N_10177,N_10173);
or U10227 (N_10227,N_10126,N_10141);
nand U10228 (N_10228,N_10073,N_10085);
and U10229 (N_10229,N_10094,N_10013);
or U10230 (N_10230,N_10036,N_10124);
or U10231 (N_10231,N_10196,N_10042);
nor U10232 (N_10232,N_10068,N_10058);
nand U10233 (N_10233,N_10118,N_10083);
or U10234 (N_10234,N_10152,N_10180);
and U10235 (N_10235,N_10077,N_10106);
or U10236 (N_10236,N_10172,N_10108);
or U10237 (N_10237,N_10088,N_10185);
nand U10238 (N_10238,N_10102,N_10044);
or U10239 (N_10239,N_10003,N_10158);
nand U10240 (N_10240,N_10117,N_10043);
nand U10241 (N_10241,N_10014,N_10000);
or U10242 (N_10242,N_10188,N_10070);
xnor U10243 (N_10243,N_10112,N_10162);
nor U10244 (N_10244,N_10079,N_10198);
and U10245 (N_10245,N_10100,N_10105);
nand U10246 (N_10246,N_10130,N_10074);
and U10247 (N_10247,N_10095,N_10147);
nand U10248 (N_10248,N_10035,N_10031);
nand U10249 (N_10249,N_10078,N_10028);
or U10250 (N_10250,N_10007,N_10011);
nor U10251 (N_10251,N_10053,N_10069);
xnor U10252 (N_10252,N_10150,N_10157);
or U10253 (N_10253,N_10024,N_10131);
nor U10254 (N_10254,N_10167,N_10050);
and U10255 (N_10255,N_10143,N_10063);
nor U10256 (N_10256,N_10049,N_10184);
and U10257 (N_10257,N_10002,N_10114);
and U10258 (N_10258,N_10142,N_10145);
and U10259 (N_10259,N_10166,N_10047);
or U10260 (N_10260,N_10059,N_10135);
or U10261 (N_10261,N_10021,N_10107);
and U10262 (N_10262,N_10005,N_10093);
or U10263 (N_10263,N_10109,N_10098);
and U10264 (N_10264,N_10062,N_10171);
and U10265 (N_10265,N_10149,N_10182);
xor U10266 (N_10266,N_10133,N_10008);
nand U10267 (N_10267,N_10057,N_10039);
and U10268 (N_10268,N_10113,N_10015);
nand U10269 (N_10269,N_10122,N_10040);
nand U10270 (N_10270,N_10060,N_10029);
xor U10271 (N_10271,N_10032,N_10075);
xnor U10272 (N_10272,N_10189,N_10187);
and U10273 (N_10273,N_10153,N_10127);
nor U10274 (N_10274,N_10136,N_10018);
xnor U10275 (N_10275,N_10168,N_10183);
nand U10276 (N_10276,N_10178,N_10016);
nor U10277 (N_10277,N_10164,N_10123);
xnor U10278 (N_10278,N_10151,N_10175);
xor U10279 (N_10279,N_10054,N_10170);
xnor U10280 (N_10280,N_10010,N_10134);
nor U10281 (N_10281,N_10051,N_10046);
nor U10282 (N_10282,N_10179,N_10199);
xor U10283 (N_10283,N_10086,N_10138);
or U10284 (N_10284,N_10034,N_10165);
or U10285 (N_10285,N_10019,N_10128);
and U10286 (N_10286,N_10193,N_10076);
nand U10287 (N_10287,N_10104,N_10066);
and U10288 (N_10288,N_10120,N_10190);
xor U10289 (N_10289,N_10090,N_10052);
xor U10290 (N_10290,N_10169,N_10191);
and U10291 (N_10291,N_10091,N_10009);
nor U10292 (N_10292,N_10186,N_10071);
and U10293 (N_10293,N_10174,N_10022);
nor U10294 (N_10294,N_10041,N_10139);
nor U10295 (N_10295,N_10163,N_10072);
nand U10296 (N_10296,N_10103,N_10061);
xnor U10297 (N_10297,N_10195,N_10148);
nand U10298 (N_10298,N_10101,N_10192);
or U10299 (N_10299,N_10037,N_10026);
and U10300 (N_10300,N_10106,N_10169);
and U10301 (N_10301,N_10136,N_10040);
xnor U10302 (N_10302,N_10116,N_10192);
or U10303 (N_10303,N_10057,N_10028);
nand U10304 (N_10304,N_10075,N_10089);
or U10305 (N_10305,N_10193,N_10127);
nor U10306 (N_10306,N_10061,N_10022);
nor U10307 (N_10307,N_10001,N_10042);
xnor U10308 (N_10308,N_10152,N_10134);
nand U10309 (N_10309,N_10074,N_10058);
and U10310 (N_10310,N_10083,N_10145);
nor U10311 (N_10311,N_10120,N_10106);
nand U10312 (N_10312,N_10131,N_10077);
nand U10313 (N_10313,N_10152,N_10064);
nand U10314 (N_10314,N_10070,N_10088);
or U10315 (N_10315,N_10075,N_10193);
and U10316 (N_10316,N_10192,N_10196);
nor U10317 (N_10317,N_10154,N_10106);
nand U10318 (N_10318,N_10070,N_10122);
and U10319 (N_10319,N_10141,N_10082);
xnor U10320 (N_10320,N_10189,N_10180);
xnor U10321 (N_10321,N_10088,N_10194);
and U10322 (N_10322,N_10018,N_10053);
nor U10323 (N_10323,N_10153,N_10182);
nor U10324 (N_10324,N_10059,N_10000);
nand U10325 (N_10325,N_10021,N_10028);
and U10326 (N_10326,N_10188,N_10040);
or U10327 (N_10327,N_10156,N_10080);
nor U10328 (N_10328,N_10032,N_10169);
nor U10329 (N_10329,N_10092,N_10112);
xnor U10330 (N_10330,N_10017,N_10030);
nand U10331 (N_10331,N_10176,N_10097);
xnor U10332 (N_10332,N_10060,N_10197);
nor U10333 (N_10333,N_10126,N_10188);
or U10334 (N_10334,N_10087,N_10032);
nand U10335 (N_10335,N_10005,N_10063);
xor U10336 (N_10336,N_10151,N_10196);
nor U10337 (N_10337,N_10125,N_10179);
or U10338 (N_10338,N_10073,N_10170);
nand U10339 (N_10339,N_10068,N_10010);
xor U10340 (N_10340,N_10092,N_10047);
and U10341 (N_10341,N_10043,N_10014);
xnor U10342 (N_10342,N_10173,N_10140);
xnor U10343 (N_10343,N_10169,N_10023);
and U10344 (N_10344,N_10180,N_10029);
nor U10345 (N_10345,N_10151,N_10116);
or U10346 (N_10346,N_10190,N_10122);
or U10347 (N_10347,N_10093,N_10148);
nand U10348 (N_10348,N_10051,N_10171);
and U10349 (N_10349,N_10180,N_10177);
nand U10350 (N_10350,N_10025,N_10066);
nand U10351 (N_10351,N_10134,N_10139);
nand U10352 (N_10352,N_10127,N_10164);
or U10353 (N_10353,N_10033,N_10131);
xor U10354 (N_10354,N_10003,N_10160);
and U10355 (N_10355,N_10073,N_10118);
nor U10356 (N_10356,N_10043,N_10167);
and U10357 (N_10357,N_10007,N_10165);
nand U10358 (N_10358,N_10019,N_10097);
or U10359 (N_10359,N_10133,N_10117);
or U10360 (N_10360,N_10076,N_10030);
nand U10361 (N_10361,N_10117,N_10091);
nand U10362 (N_10362,N_10182,N_10010);
xor U10363 (N_10363,N_10026,N_10029);
or U10364 (N_10364,N_10009,N_10081);
nand U10365 (N_10365,N_10095,N_10025);
nor U10366 (N_10366,N_10112,N_10005);
xnor U10367 (N_10367,N_10019,N_10176);
and U10368 (N_10368,N_10153,N_10165);
xor U10369 (N_10369,N_10146,N_10082);
and U10370 (N_10370,N_10094,N_10176);
nand U10371 (N_10371,N_10012,N_10098);
and U10372 (N_10372,N_10042,N_10033);
and U10373 (N_10373,N_10129,N_10148);
or U10374 (N_10374,N_10044,N_10170);
or U10375 (N_10375,N_10034,N_10097);
and U10376 (N_10376,N_10143,N_10021);
and U10377 (N_10377,N_10172,N_10072);
xor U10378 (N_10378,N_10108,N_10000);
nand U10379 (N_10379,N_10049,N_10106);
or U10380 (N_10380,N_10016,N_10084);
or U10381 (N_10381,N_10175,N_10113);
xor U10382 (N_10382,N_10158,N_10115);
or U10383 (N_10383,N_10135,N_10188);
and U10384 (N_10384,N_10129,N_10095);
xor U10385 (N_10385,N_10001,N_10124);
nor U10386 (N_10386,N_10024,N_10184);
nor U10387 (N_10387,N_10185,N_10022);
and U10388 (N_10388,N_10171,N_10192);
nor U10389 (N_10389,N_10099,N_10158);
and U10390 (N_10390,N_10105,N_10079);
xnor U10391 (N_10391,N_10174,N_10026);
or U10392 (N_10392,N_10001,N_10040);
or U10393 (N_10393,N_10082,N_10181);
or U10394 (N_10394,N_10195,N_10039);
nand U10395 (N_10395,N_10100,N_10031);
and U10396 (N_10396,N_10130,N_10075);
xnor U10397 (N_10397,N_10058,N_10081);
nor U10398 (N_10398,N_10196,N_10107);
xnor U10399 (N_10399,N_10080,N_10184);
and U10400 (N_10400,N_10373,N_10209);
and U10401 (N_10401,N_10271,N_10272);
xnor U10402 (N_10402,N_10320,N_10364);
nand U10403 (N_10403,N_10232,N_10252);
and U10404 (N_10404,N_10306,N_10262);
nand U10405 (N_10405,N_10315,N_10326);
or U10406 (N_10406,N_10205,N_10259);
xor U10407 (N_10407,N_10291,N_10263);
nor U10408 (N_10408,N_10212,N_10229);
or U10409 (N_10409,N_10250,N_10357);
and U10410 (N_10410,N_10362,N_10280);
xor U10411 (N_10411,N_10254,N_10388);
and U10412 (N_10412,N_10313,N_10219);
nand U10413 (N_10413,N_10312,N_10398);
or U10414 (N_10414,N_10243,N_10375);
and U10415 (N_10415,N_10275,N_10374);
nor U10416 (N_10416,N_10257,N_10247);
or U10417 (N_10417,N_10296,N_10227);
nor U10418 (N_10418,N_10359,N_10222);
or U10419 (N_10419,N_10385,N_10300);
nand U10420 (N_10420,N_10349,N_10307);
xor U10421 (N_10421,N_10293,N_10303);
nand U10422 (N_10422,N_10305,N_10365);
nand U10423 (N_10423,N_10282,N_10234);
and U10424 (N_10424,N_10288,N_10347);
xnor U10425 (N_10425,N_10322,N_10346);
nand U10426 (N_10426,N_10204,N_10342);
nand U10427 (N_10427,N_10336,N_10202);
xnor U10428 (N_10428,N_10258,N_10399);
nor U10429 (N_10429,N_10338,N_10390);
nand U10430 (N_10430,N_10201,N_10290);
nand U10431 (N_10431,N_10239,N_10397);
nand U10432 (N_10432,N_10333,N_10294);
or U10433 (N_10433,N_10215,N_10200);
nand U10434 (N_10434,N_10265,N_10238);
or U10435 (N_10435,N_10292,N_10248);
xor U10436 (N_10436,N_10356,N_10353);
nand U10437 (N_10437,N_10345,N_10330);
xnor U10438 (N_10438,N_10331,N_10233);
nor U10439 (N_10439,N_10376,N_10270);
and U10440 (N_10440,N_10381,N_10279);
xor U10441 (N_10441,N_10264,N_10278);
or U10442 (N_10442,N_10335,N_10207);
or U10443 (N_10443,N_10389,N_10277);
nor U10444 (N_10444,N_10253,N_10379);
or U10445 (N_10445,N_10273,N_10268);
and U10446 (N_10446,N_10318,N_10255);
nand U10447 (N_10447,N_10220,N_10392);
or U10448 (N_10448,N_10334,N_10350);
and U10449 (N_10449,N_10236,N_10358);
nor U10450 (N_10450,N_10340,N_10395);
or U10451 (N_10451,N_10383,N_10304);
and U10452 (N_10452,N_10355,N_10321);
nand U10453 (N_10453,N_10394,N_10206);
or U10454 (N_10454,N_10391,N_10244);
nand U10455 (N_10455,N_10285,N_10241);
xnor U10456 (N_10456,N_10323,N_10302);
xnor U10457 (N_10457,N_10245,N_10319);
xnor U10458 (N_10458,N_10351,N_10308);
nor U10459 (N_10459,N_10328,N_10289);
nor U10460 (N_10460,N_10377,N_10286);
nand U10461 (N_10461,N_10203,N_10295);
or U10462 (N_10462,N_10208,N_10283);
nand U10463 (N_10463,N_10281,N_10210);
or U10464 (N_10464,N_10343,N_10325);
nand U10465 (N_10465,N_10231,N_10276);
xnor U10466 (N_10466,N_10235,N_10225);
nor U10467 (N_10467,N_10299,N_10297);
or U10468 (N_10468,N_10329,N_10216);
nor U10469 (N_10469,N_10382,N_10266);
xor U10470 (N_10470,N_10256,N_10274);
or U10471 (N_10471,N_10301,N_10217);
xnor U10472 (N_10472,N_10367,N_10332);
nand U10473 (N_10473,N_10309,N_10371);
and U10474 (N_10474,N_10230,N_10361);
xnor U10475 (N_10475,N_10354,N_10363);
nor U10476 (N_10476,N_10251,N_10372);
xnor U10477 (N_10477,N_10387,N_10267);
nand U10478 (N_10478,N_10226,N_10224);
or U10479 (N_10479,N_10284,N_10228);
nand U10480 (N_10480,N_10240,N_10368);
and U10481 (N_10481,N_10242,N_10298);
or U10482 (N_10482,N_10369,N_10211);
nor U10483 (N_10483,N_10213,N_10339);
xnor U10484 (N_10484,N_10380,N_10370);
or U10485 (N_10485,N_10393,N_10360);
and U10486 (N_10486,N_10344,N_10348);
nor U10487 (N_10487,N_10218,N_10341);
nand U10488 (N_10488,N_10337,N_10384);
nor U10489 (N_10489,N_10237,N_10260);
xnor U10490 (N_10490,N_10324,N_10396);
nand U10491 (N_10491,N_10246,N_10316);
nor U10492 (N_10492,N_10311,N_10249);
xnor U10493 (N_10493,N_10269,N_10310);
nand U10494 (N_10494,N_10287,N_10386);
nor U10495 (N_10495,N_10221,N_10317);
and U10496 (N_10496,N_10378,N_10327);
or U10497 (N_10497,N_10214,N_10314);
xnor U10498 (N_10498,N_10261,N_10352);
and U10499 (N_10499,N_10366,N_10223);
or U10500 (N_10500,N_10334,N_10381);
xor U10501 (N_10501,N_10315,N_10220);
nand U10502 (N_10502,N_10316,N_10323);
and U10503 (N_10503,N_10379,N_10316);
xor U10504 (N_10504,N_10304,N_10204);
xor U10505 (N_10505,N_10301,N_10266);
xnor U10506 (N_10506,N_10368,N_10258);
and U10507 (N_10507,N_10375,N_10235);
or U10508 (N_10508,N_10398,N_10336);
xor U10509 (N_10509,N_10243,N_10215);
xnor U10510 (N_10510,N_10369,N_10288);
and U10511 (N_10511,N_10299,N_10310);
xnor U10512 (N_10512,N_10307,N_10362);
or U10513 (N_10513,N_10357,N_10364);
nand U10514 (N_10514,N_10280,N_10310);
nor U10515 (N_10515,N_10299,N_10320);
nand U10516 (N_10516,N_10208,N_10391);
nand U10517 (N_10517,N_10376,N_10222);
or U10518 (N_10518,N_10326,N_10202);
and U10519 (N_10519,N_10329,N_10332);
nor U10520 (N_10520,N_10245,N_10371);
and U10521 (N_10521,N_10270,N_10310);
and U10522 (N_10522,N_10201,N_10210);
xor U10523 (N_10523,N_10397,N_10242);
nor U10524 (N_10524,N_10227,N_10235);
nor U10525 (N_10525,N_10316,N_10380);
nor U10526 (N_10526,N_10296,N_10254);
nand U10527 (N_10527,N_10228,N_10283);
nor U10528 (N_10528,N_10256,N_10288);
xnor U10529 (N_10529,N_10281,N_10303);
nand U10530 (N_10530,N_10365,N_10348);
nor U10531 (N_10531,N_10201,N_10303);
nor U10532 (N_10532,N_10363,N_10236);
nand U10533 (N_10533,N_10371,N_10292);
and U10534 (N_10534,N_10268,N_10286);
or U10535 (N_10535,N_10217,N_10276);
or U10536 (N_10536,N_10309,N_10313);
and U10537 (N_10537,N_10397,N_10282);
and U10538 (N_10538,N_10308,N_10210);
xnor U10539 (N_10539,N_10339,N_10205);
nand U10540 (N_10540,N_10325,N_10237);
xor U10541 (N_10541,N_10200,N_10203);
or U10542 (N_10542,N_10385,N_10290);
or U10543 (N_10543,N_10394,N_10301);
or U10544 (N_10544,N_10275,N_10306);
and U10545 (N_10545,N_10300,N_10365);
xor U10546 (N_10546,N_10342,N_10279);
nand U10547 (N_10547,N_10383,N_10261);
or U10548 (N_10548,N_10214,N_10230);
or U10549 (N_10549,N_10241,N_10373);
and U10550 (N_10550,N_10373,N_10376);
xor U10551 (N_10551,N_10300,N_10353);
nand U10552 (N_10552,N_10329,N_10204);
or U10553 (N_10553,N_10386,N_10231);
xnor U10554 (N_10554,N_10297,N_10293);
nor U10555 (N_10555,N_10335,N_10233);
and U10556 (N_10556,N_10393,N_10361);
xnor U10557 (N_10557,N_10360,N_10269);
nand U10558 (N_10558,N_10255,N_10219);
and U10559 (N_10559,N_10308,N_10226);
nand U10560 (N_10560,N_10354,N_10334);
nor U10561 (N_10561,N_10248,N_10309);
nor U10562 (N_10562,N_10363,N_10320);
and U10563 (N_10563,N_10287,N_10327);
nand U10564 (N_10564,N_10363,N_10331);
or U10565 (N_10565,N_10225,N_10312);
nand U10566 (N_10566,N_10205,N_10388);
or U10567 (N_10567,N_10375,N_10390);
or U10568 (N_10568,N_10314,N_10343);
xnor U10569 (N_10569,N_10202,N_10249);
and U10570 (N_10570,N_10334,N_10260);
and U10571 (N_10571,N_10284,N_10377);
nand U10572 (N_10572,N_10206,N_10399);
nor U10573 (N_10573,N_10345,N_10248);
and U10574 (N_10574,N_10271,N_10277);
xor U10575 (N_10575,N_10219,N_10363);
xor U10576 (N_10576,N_10265,N_10385);
and U10577 (N_10577,N_10289,N_10258);
or U10578 (N_10578,N_10236,N_10223);
nor U10579 (N_10579,N_10388,N_10374);
and U10580 (N_10580,N_10266,N_10216);
nand U10581 (N_10581,N_10222,N_10233);
nor U10582 (N_10582,N_10344,N_10249);
nor U10583 (N_10583,N_10255,N_10204);
nor U10584 (N_10584,N_10317,N_10279);
nand U10585 (N_10585,N_10357,N_10279);
nand U10586 (N_10586,N_10371,N_10258);
and U10587 (N_10587,N_10302,N_10218);
nor U10588 (N_10588,N_10296,N_10329);
or U10589 (N_10589,N_10396,N_10376);
nand U10590 (N_10590,N_10304,N_10265);
nor U10591 (N_10591,N_10285,N_10333);
or U10592 (N_10592,N_10389,N_10347);
and U10593 (N_10593,N_10343,N_10382);
or U10594 (N_10594,N_10374,N_10235);
and U10595 (N_10595,N_10209,N_10393);
or U10596 (N_10596,N_10360,N_10334);
and U10597 (N_10597,N_10360,N_10283);
or U10598 (N_10598,N_10351,N_10240);
nor U10599 (N_10599,N_10390,N_10302);
and U10600 (N_10600,N_10423,N_10513);
or U10601 (N_10601,N_10452,N_10419);
or U10602 (N_10602,N_10562,N_10592);
xnor U10603 (N_10603,N_10576,N_10572);
nor U10604 (N_10604,N_10460,N_10433);
xor U10605 (N_10605,N_10570,N_10546);
and U10606 (N_10606,N_10468,N_10422);
nor U10607 (N_10607,N_10580,N_10434);
and U10608 (N_10608,N_10547,N_10517);
nand U10609 (N_10609,N_10537,N_10494);
nand U10610 (N_10610,N_10578,N_10443);
nor U10611 (N_10611,N_10441,N_10463);
xor U10612 (N_10612,N_10448,N_10490);
nor U10613 (N_10613,N_10535,N_10473);
and U10614 (N_10614,N_10530,N_10588);
nand U10615 (N_10615,N_10451,N_10557);
or U10616 (N_10616,N_10539,N_10488);
nor U10617 (N_10617,N_10543,N_10558);
xnor U10618 (N_10618,N_10408,N_10507);
or U10619 (N_10619,N_10511,N_10401);
xor U10620 (N_10620,N_10476,N_10516);
xnor U10621 (N_10621,N_10538,N_10548);
xor U10622 (N_10622,N_10523,N_10484);
and U10623 (N_10623,N_10594,N_10501);
xnor U10624 (N_10624,N_10591,N_10565);
and U10625 (N_10625,N_10426,N_10575);
nor U10626 (N_10626,N_10446,N_10462);
nand U10627 (N_10627,N_10403,N_10552);
nand U10628 (N_10628,N_10550,N_10458);
or U10629 (N_10629,N_10514,N_10568);
nor U10630 (N_10630,N_10406,N_10472);
xor U10631 (N_10631,N_10508,N_10470);
or U10632 (N_10632,N_10553,N_10402);
and U10633 (N_10633,N_10429,N_10521);
xnor U10634 (N_10634,N_10481,N_10482);
and U10635 (N_10635,N_10589,N_10499);
nand U10636 (N_10636,N_10556,N_10442);
nor U10637 (N_10637,N_10559,N_10461);
or U10638 (N_10638,N_10524,N_10542);
nand U10639 (N_10639,N_10497,N_10456);
nand U10640 (N_10640,N_10420,N_10487);
or U10641 (N_10641,N_10489,N_10454);
nand U10642 (N_10642,N_10438,N_10596);
or U10643 (N_10643,N_10503,N_10549);
or U10644 (N_10644,N_10571,N_10525);
or U10645 (N_10645,N_10417,N_10449);
nand U10646 (N_10646,N_10566,N_10409);
nand U10647 (N_10647,N_10432,N_10486);
xnor U10648 (N_10648,N_10540,N_10581);
or U10649 (N_10649,N_10455,N_10551);
and U10650 (N_10650,N_10431,N_10522);
xnor U10651 (N_10651,N_10416,N_10512);
and U10652 (N_10652,N_10541,N_10453);
nand U10653 (N_10653,N_10424,N_10509);
and U10654 (N_10654,N_10555,N_10593);
xnor U10655 (N_10655,N_10532,N_10407);
nor U10656 (N_10656,N_10413,N_10465);
nor U10657 (N_10657,N_10436,N_10595);
or U10658 (N_10658,N_10506,N_10518);
xnor U10659 (N_10659,N_10444,N_10527);
nand U10660 (N_10660,N_10475,N_10469);
or U10661 (N_10661,N_10439,N_10437);
xnor U10662 (N_10662,N_10585,N_10582);
nor U10663 (N_10663,N_10466,N_10586);
nor U10664 (N_10664,N_10561,N_10405);
nor U10665 (N_10665,N_10598,N_10400);
or U10666 (N_10666,N_10564,N_10440);
or U10667 (N_10667,N_10428,N_10471);
and U10668 (N_10668,N_10464,N_10412);
nand U10669 (N_10669,N_10536,N_10404);
nor U10670 (N_10670,N_10599,N_10545);
and U10671 (N_10671,N_10474,N_10563);
nor U10672 (N_10672,N_10567,N_10410);
or U10673 (N_10673,N_10435,N_10583);
nand U10674 (N_10674,N_10579,N_10483);
or U10675 (N_10675,N_10520,N_10477);
and U10676 (N_10676,N_10418,N_10574);
or U10677 (N_10677,N_10529,N_10496);
nor U10678 (N_10678,N_10528,N_10573);
xnor U10679 (N_10679,N_10415,N_10533);
or U10680 (N_10680,N_10531,N_10479);
nor U10681 (N_10681,N_10554,N_10498);
and U10682 (N_10682,N_10457,N_10500);
or U10683 (N_10683,N_10414,N_10450);
and U10684 (N_10684,N_10430,N_10491);
or U10685 (N_10685,N_10534,N_10478);
and U10686 (N_10686,N_10495,N_10519);
and U10687 (N_10687,N_10515,N_10492);
xnor U10688 (N_10688,N_10485,N_10421);
nor U10689 (N_10689,N_10587,N_10577);
nor U10690 (N_10690,N_10544,N_10502);
nand U10691 (N_10691,N_10447,N_10493);
xor U10692 (N_10692,N_10597,N_10560);
or U10693 (N_10693,N_10505,N_10425);
or U10694 (N_10694,N_10510,N_10526);
xnor U10695 (N_10695,N_10467,N_10411);
nand U10696 (N_10696,N_10504,N_10569);
nand U10697 (N_10697,N_10480,N_10584);
xnor U10698 (N_10698,N_10459,N_10590);
and U10699 (N_10699,N_10427,N_10445);
nor U10700 (N_10700,N_10411,N_10545);
and U10701 (N_10701,N_10514,N_10541);
or U10702 (N_10702,N_10554,N_10439);
nand U10703 (N_10703,N_10461,N_10458);
and U10704 (N_10704,N_10461,N_10573);
or U10705 (N_10705,N_10404,N_10466);
and U10706 (N_10706,N_10512,N_10586);
nand U10707 (N_10707,N_10455,N_10496);
and U10708 (N_10708,N_10517,N_10531);
xnor U10709 (N_10709,N_10432,N_10442);
and U10710 (N_10710,N_10551,N_10458);
nor U10711 (N_10711,N_10440,N_10497);
xnor U10712 (N_10712,N_10513,N_10475);
xnor U10713 (N_10713,N_10514,N_10565);
nor U10714 (N_10714,N_10424,N_10551);
or U10715 (N_10715,N_10557,N_10441);
or U10716 (N_10716,N_10569,N_10452);
nand U10717 (N_10717,N_10424,N_10536);
xnor U10718 (N_10718,N_10465,N_10420);
nand U10719 (N_10719,N_10529,N_10530);
xor U10720 (N_10720,N_10479,N_10591);
or U10721 (N_10721,N_10587,N_10502);
nor U10722 (N_10722,N_10536,N_10416);
or U10723 (N_10723,N_10563,N_10418);
or U10724 (N_10724,N_10566,N_10545);
nor U10725 (N_10725,N_10479,N_10400);
and U10726 (N_10726,N_10451,N_10538);
nor U10727 (N_10727,N_10446,N_10416);
xor U10728 (N_10728,N_10430,N_10499);
or U10729 (N_10729,N_10435,N_10488);
xnor U10730 (N_10730,N_10497,N_10523);
or U10731 (N_10731,N_10488,N_10404);
nor U10732 (N_10732,N_10447,N_10401);
or U10733 (N_10733,N_10548,N_10409);
and U10734 (N_10734,N_10546,N_10410);
or U10735 (N_10735,N_10539,N_10540);
and U10736 (N_10736,N_10428,N_10432);
nor U10737 (N_10737,N_10554,N_10558);
xnor U10738 (N_10738,N_10422,N_10444);
and U10739 (N_10739,N_10424,N_10569);
nor U10740 (N_10740,N_10527,N_10491);
nand U10741 (N_10741,N_10487,N_10493);
or U10742 (N_10742,N_10469,N_10471);
xor U10743 (N_10743,N_10438,N_10486);
and U10744 (N_10744,N_10576,N_10477);
xor U10745 (N_10745,N_10507,N_10450);
nor U10746 (N_10746,N_10434,N_10502);
or U10747 (N_10747,N_10570,N_10583);
and U10748 (N_10748,N_10443,N_10448);
or U10749 (N_10749,N_10468,N_10461);
and U10750 (N_10750,N_10586,N_10434);
nor U10751 (N_10751,N_10527,N_10583);
nand U10752 (N_10752,N_10556,N_10444);
or U10753 (N_10753,N_10580,N_10561);
or U10754 (N_10754,N_10492,N_10570);
nand U10755 (N_10755,N_10556,N_10485);
or U10756 (N_10756,N_10424,N_10402);
nand U10757 (N_10757,N_10590,N_10426);
nand U10758 (N_10758,N_10412,N_10575);
and U10759 (N_10759,N_10465,N_10587);
or U10760 (N_10760,N_10446,N_10562);
nor U10761 (N_10761,N_10447,N_10436);
and U10762 (N_10762,N_10514,N_10521);
nor U10763 (N_10763,N_10544,N_10400);
and U10764 (N_10764,N_10423,N_10555);
and U10765 (N_10765,N_10444,N_10592);
nor U10766 (N_10766,N_10439,N_10546);
xnor U10767 (N_10767,N_10428,N_10583);
or U10768 (N_10768,N_10465,N_10519);
xor U10769 (N_10769,N_10533,N_10599);
xor U10770 (N_10770,N_10425,N_10592);
or U10771 (N_10771,N_10575,N_10511);
nand U10772 (N_10772,N_10520,N_10537);
xor U10773 (N_10773,N_10549,N_10582);
nor U10774 (N_10774,N_10531,N_10587);
and U10775 (N_10775,N_10525,N_10457);
nor U10776 (N_10776,N_10429,N_10569);
and U10777 (N_10777,N_10443,N_10474);
nand U10778 (N_10778,N_10537,N_10401);
or U10779 (N_10779,N_10563,N_10531);
or U10780 (N_10780,N_10556,N_10472);
xor U10781 (N_10781,N_10453,N_10438);
or U10782 (N_10782,N_10455,N_10510);
nor U10783 (N_10783,N_10541,N_10424);
xor U10784 (N_10784,N_10498,N_10474);
nand U10785 (N_10785,N_10481,N_10414);
nand U10786 (N_10786,N_10457,N_10466);
xor U10787 (N_10787,N_10403,N_10448);
xor U10788 (N_10788,N_10407,N_10499);
and U10789 (N_10789,N_10426,N_10442);
xor U10790 (N_10790,N_10510,N_10446);
or U10791 (N_10791,N_10591,N_10451);
nor U10792 (N_10792,N_10521,N_10411);
xor U10793 (N_10793,N_10529,N_10548);
nand U10794 (N_10794,N_10434,N_10404);
and U10795 (N_10795,N_10568,N_10501);
nor U10796 (N_10796,N_10503,N_10480);
and U10797 (N_10797,N_10466,N_10563);
or U10798 (N_10798,N_10447,N_10405);
and U10799 (N_10799,N_10583,N_10521);
or U10800 (N_10800,N_10790,N_10689);
nor U10801 (N_10801,N_10629,N_10756);
or U10802 (N_10802,N_10789,N_10691);
or U10803 (N_10803,N_10670,N_10616);
or U10804 (N_10804,N_10640,N_10698);
and U10805 (N_10805,N_10633,N_10755);
nand U10806 (N_10806,N_10617,N_10664);
and U10807 (N_10807,N_10721,N_10605);
nand U10808 (N_10808,N_10602,N_10742);
nand U10809 (N_10809,N_10711,N_10621);
nor U10810 (N_10810,N_10739,N_10730);
xor U10811 (N_10811,N_10705,N_10646);
nand U10812 (N_10812,N_10626,N_10672);
and U10813 (N_10813,N_10759,N_10679);
or U10814 (N_10814,N_10684,N_10775);
and U10815 (N_10815,N_10671,N_10728);
and U10816 (N_10816,N_10787,N_10763);
nor U10817 (N_10817,N_10611,N_10638);
or U10818 (N_10818,N_10645,N_10761);
nand U10819 (N_10819,N_10639,N_10627);
nor U10820 (N_10820,N_10753,N_10666);
or U10821 (N_10821,N_10771,N_10600);
nor U10822 (N_10822,N_10752,N_10700);
xor U10823 (N_10823,N_10612,N_10681);
xnor U10824 (N_10824,N_10734,N_10604);
and U10825 (N_10825,N_10783,N_10647);
and U10826 (N_10826,N_10714,N_10786);
xnor U10827 (N_10827,N_10675,N_10662);
nand U10828 (N_10828,N_10634,N_10660);
nand U10829 (N_10829,N_10701,N_10674);
nor U10830 (N_10830,N_10614,N_10729);
and U10831 (N_10831,N_10668,N_10732);
nand U10832 (N_10832,N_10650,N_10607);
xor U10833 (N_10833,N_10685,N_10657);
nand U10834 (N_10834,N_10619,N_10628);
and U10835 (N_10835,N_10798,N_10618);
xor U10836 (N_10836,N_10613,N_10696);
or U10837 (N_10837,N_10750,N_10770);
xor U10838 (N_10838,N_10661,N_10731);
nor U10839 (N_10839,N_10688,N_10765);
xor U10840 (N_10840,N_10768,N_10720);
and U10841 (N_10841,N_10623,N_10766);
nand U10842 (N_10842,N_10717,N_10776);
nand U10843 (N_10843,N_10649,N_10682);
and U10844 (N_10844,N_10788,N_10779);
nand U10845 (N_10845,N_10757,N_10725);
and U10846 (N_10846,N_10778,N_10769);
and U10847 (N_10847,N_10620,N_10697);
nand U10848 (N_10848,N_10652,N_10694);
nor U10849 (N_10849,N_10601,N_10784);
nand U10850 (N_10850,N_10665,N_10635);
nand U10851 (N_10851,N_10631,N_10738);
xor U10852 (N_10852,N_10773,N_10749);
xor U10853 (N_10853,N_10777,N_10658);
nand U10854 (N_10854,N_10699,N_10710);
nand U10855 (N_10855,N_10683,N_10726);
xnor U10856 (N_10856,N_10767,N_10736);
nor U10857 (N_10857,N_10719,N_10608);
or U10858 (N_10858,N_10764,N_10642);
xnor U10859 (N_10859,N_10792,N_10606);
xnor U10860 (N_10860,N_10722,N_10706);
xnor U10861 (N_10861,N_10795,N_10758);
nor U10862 (N_10862,N_10751,N_10702);
and U10863 (N_10863,N_10667,N_10630);
or U10864 (N_10864,N_10740,N_10609);
and U10865 (N_10865,N_10796,N_10793);
nor U10866 (N_10866,N_10708,N_10727);
xnor U10867 (N_10867,N_10718,N_10754);
and U10868 (N_10868,N_10680,N_10676);
nand U10869 (N_10869,N_10655,N_10760);
or U10870 (N_10870,N_10715,N_10644);
xnor U10871 (N_10871,N_10632,N_10677);
and U10872 (N_10872,N_10772,N_10704);
nor U10873 (N_10873,N_10774,N_10690);
xor U10874 (N_10874,N_10762,N_10678);
nor U10875 (N_10875,N_10724,N_10799);
or U10876 (N_10876,N_10692,N_10748);
and U10877 (N_10877,N_10673,N_10741);
xor U10878 (N_10878,N_10735,N_10636);
nor U10879 (N_10879,N_10797,N_10785);
and U10880 (N_10880,N_10791,N_10780);
nor U10881 (N_10881,N_10693,N_10695);
and U10882 (N_10882,N_10643,N_10733);
nand U10883 (N_10883,N_10713,N_10745);
or U10884 (N_10884,N_10737,N_10641);
nor U10885 (N_10885,N_10637,N_10651);
xor U10886 (N_10886,N_10782,N_10653);
nor U10887 (N_10887,N_10747,N_10794);
and U10888 (N_10888,N_10624,N_10686);
or U10889 (N_10889,N_10712,N_10603);
xor U10890 (N_10890,N_10659,N_10716);
nor U10891 (N_10891,N_10622,N_10663);
or U10892 (N_10892,N_10744,N_10654);
and U10893 (N_10893,N_10707,N_10743);
and U10894 (N_10894,N_10656,N_10610);
nor U10895 (N_10895,N_10625,N_10648);
nor U10896 (N_10896,N_10723,N_10781);
xnor U10897 (N_10897,N_10746,N_10687);
nand U10898 (N_10898,N_10669,N_10709);
or U10899 (N_10899,N_10615,N_10703);
nand U10900 (N_10900,N_10683,N_10658);
nand U10901 (N_10901,N_10687,N_10693);
xnor U10902 (N_10902,N_10766,N_10722);
nor U10903 (N_10903,N_10695,N_10651);
nand U10904 (N_10904,N_10774,N_10738);
and U10905 (N_10905,N_10626,N_10616);
nor U10906 (N_10906,N_10763,N_10653);
nor U10907 (N_10907,N_10681,N_10772);
nand U10908 (N_10908,N_10776,N_10701);
xnor U10909 (N_10909,N_10633,N_10605);
or U10910 (N_10910,N_10773,N_10737);
or U10911 (N_10911,N_10770,N_10613);
or U10912 (N_10912,N_10785,N_10726);
nor U10913 (N_10913,N_10740,N_10679);
nand U10914 (N_10914,N_10610,N_10789);
and U10915 (N_10915,N_10714,N_10725);
or U10916 (N_10916,N_10715,N_10786);
nor U10917 (N_10917,N_10699,N_10644);
nor U10918 (N_10918,N_10639,N_10749);
nand U10919 (N_10919,N_10616,N_10774);
nand U10920 (N_10920,N_10715,N_10705);
or U10921 (N_10921,N_10656,N_10680);
or U10922 (N_10922,N_10688,N_10660);
or U10923 (N_10923,N_10766,N_10640);
and U10924 (N_10924,N_10723,N_10738);
nand U10925 (N_10925,N_10715,N_10615);
or U10926 (N_10926,N_10739,N_10793);
nor U10927 (N_10927,N_10782,N_10798);
nand U10928 (N_10928,N_10639,N_10651);
xnor U10929 (N_10929,N_10609,N_10757);
and U10930 (N_10930,N_10781,N_10755);
nor U10931 (N_10931,N_10648,N_10709);
and U10932 (N_10932,N_10603,N_10791);
nand U10933 (N_10933,N_10686,N_10740);
and U10934 (N_10934,N_10726,N_10724);
or U10935 (N_10935,N_10783,N_10734);
xor U10936 (N_10936,N_10622,N_10786);
or U10937 (N_10937,N_10703,N_10762);
and U10938 (N_10938,N_10724,N_10795);
or U10939 (N_10939,N_10648,N_10731);
and U10940 (N_10940,N_10661,N_10788);
and U10941 (N_10941,N_10720,N_10607);
nor U10942 (N_10942,N_10673,N_10712);
nand U10943 (N_10943,N_10795,N_10768);
or U10944 (N_10944,N_10679,N_10723);
nor U10945 (N_10945,N_10665,N_10708);
and U10946 (N_10946,N_10604,N_10770);
or U10947 (N_10947,N_10645,N_10621);
nor U10948 (N_10948,N_10640,N_10722);
xnor U10949 (N_10949,N_10695,N_10738);
nor U10950 (N_10950,N_10685,N_10607);
xnor U10951 (N_10951,N_10782,N_10793);
xor U10952 (N_10952,N_10740,N_10724);
nand U10953 (N_10953,N_10641,N_10787);
and U10954 (N_10954,N_10611,N_10704);
xnor U10955 (N_10955,N_10633,N_10798);
nand U10956 (N_10956,N_10669,N_10642);
and U10957 (N_10957,N_10668,N_10611);
nor U10958 (N_10958,N_10704,N_10634);
nor U10959 (N_10959,N_10688,N_10622);
and U10960 (N_10960,N_10672,N_10719);
nand U10961 (N_10961,N_10635,N_10727);
xor U10962 (N_10962,N_10776,N_10685);
xor U10963 (N_10963,N_10732,N_10700);
xnor U10964 (N_10964,N_10700,N_10672);
and U10965 (N_10965,N_10754,N_10674);
xnor U10966 (N_10966,N_10779,N_10667);
nor U10967 (N_10967,N_10627,N_10678);
xor U10968 (N_10968,N_10768,N_10674);
or U10969 (N_10969,N_10639,N_10666);
or U10970 (N_10970,N_10647,N_10667);
nor U10971 (N_10971,N_10729,N_10714);
nor U10972 (N_10972,N_10689,N_10631);
or U10973 (N_10973,N_10739,N_10662);
xnor U10974 (N_10974,N_10640,N_10663);
nand U10975 (N_10975,N_10647,N_10709);
and U10976 (N_10976,N_10640,N_10732);
or U10977 (N_10977,N_10720,N_10764);
nand U10978 (N_10978,N_10784,N_10685);
xor U10979 (N_10979,N_10716,N_10780);
nand U10980 (N_10980,N_10771,N_10604);
and U10981 (N_10981,N_10794,N_10613);
nand U10982 (N_10982,N_10776,N_10732);
and U10983 (N_10983,N_10618,N_10665);
or U10984 (N_10984,N_10789,N_10755);
or U10985 (N_10985,N_10707,N_10745);
nand U10986 (N_10986,N_10757,N_10722);
nand U10987 (N_10987,N_10789,N_10796);
and U10988 (N_10988,N_10629,N_10742);
or U10989 (N_10989,N_10740,N_10745);
nor U10990 (N_10990,N_10653,N_10704);
nor U10991 (N_10991,N_10691,N_10710);
and U10992 (N_10992,N_10741,N_10668);
nor U10993 (N_10993,N_10665,N_10641);
nor U10994 (N_10994,N_10783,N_10661);
nand U10995 (N_10995,N_10695,N_10677);
and U10996 (N_10996,N_10744,N_10755);
and U10997 (N_10997,N_10616,N_10791);
or U10998 (N_10998,N_10787,N_10748);
nand U10999 (N_10999,N_10701,N_10602);
and U11000 (N_11000,N_10980,N_10911);
nor U11001 (N_11001,N_10825,N_10815);
nand U11002 (N_11002,N_10881,N_10889);
xnor U11003 (N_11003,N_10966,N_10840);
and U11004 (N_11004,N_10894,N_10874);
xor U11005 (N_11005,N_10865,N_10992);
or U11006 (N_11006,N_10996,N_10871);
nand U11007 (N_11007,N_10899,N_10985);
nand U11008 (N_11008,N_10901,N_10941);
or U11009 (N_11009,N_10998,N_10895);
or U11010 (N_11010,N_10858,N_10991);
xor U11011 (N_11011,N_10801,N_10999);
and U11012 (N_11012,N_10893,N_10818);
nand U11013 (N_11013,N_10988,N_10957);
or U11014 (N_11014,N_10967,N_10882);
and U11015 (N_11015,N_10890,N_10832);
xnor U11016 (N_11016,N_10886,N_10974);
nor U11017 (N_11017,N_10860,N_10955);
nor U11018 (N_11018,N_10912,N_10908);
and U11019 (N_11019,N_10961,N_10896);
xor U11020 (N_11020,N_10969,N_10829);
or U11021 (N_11021,N_10934,N_10936);
and U11022 (N_11022,N_10855,N_10960);
xor U11023 (N_11023,N_10875,N_10852);
nor U11024 (N_11024,N_10831,N_10953);
or U11025 (N_11025,N_10971,N_10869);
and U11026 (N_11026,N_10888,N_10931);
nor U11027 (N_11027,N_10986,N_10826);
and U11028 (N_11028,N_10977,N_10823);
or U11029 (N_11029,N_10820,N_10859);
and U11030 (N_11030,N_10834,N_10905);
or U11031 (N_11031,N_10868,N_10959);
and U11032 (N_11032,N_10997,N_10973);
nand U11033 (N_11033,N_10812,N_10811);
and U11034 (N_11034,N_10947,N_10981);
nand U11035 (N_11035,N_10849,N_10824);
and U11036 (N_11036,N_10809,N_10958);
nand U11037 (N_11037,N_10923,N_10925);
xor U11038 (N_11038,N_10841,N_10983);
or U11039 (N_11039,N_10845,N_10951);
xor U11040 (N_11040,N_10975,N_10900);
and U11041 (N_11041,N_10844,N_10990);
nor U11042 (N_11042,N_10827,N_10927);
xor U11043 (N_11043,N_10919,N_10880);
xnor U11044 (N_11044,N_10968,N_10857);
nand U11045 (N_11045,N_10839,N_10984);
nor U11046 (N_11046,N_10906,N_10939);
or U11047 (N_11047,N_10805,N_10982);
and U11048 (N_11048,N_10879,N_10822);
or U11049 (N_11049,N_10819,N_10989);
xnor U11050 (N_11050,N_10856,N_10924);
or U11051 (N_11051,N_10804,N_10816);
and U11052 (N_11052,N_10943,N_10942);
nor U11053 (N_11053,N_10861,N_10814);
xor U11054 (N_11054,N_10902,N_10870);
xnor U11055 (N_11055,N_10883,N_10876);
or U11056 (N_11056,N_10897,N_10828);
nand U11057 (N_11057,N_10863,N_10945);
xor U11058 (N_11058,N_10938,N_10910);
xor U11059 (N_11059,N_10836,N_10949);
nor U11060 (N_11060,N_10930,N_10956);
xor U11061 (N_11061,N_10914,N_10850);
nand U11062 (N_11062,N_10847,N_10921);
xor U11063 (N_11063,N_10922,N_10918);
xnor U11064 (N_11064,N_10948,N_10995);
and U11065 (N_11065,N_10846,N_10937);
xor U11066 (N_11066,N_10813,N_10810);
xnor U11067 (N_11067,N_10913,N_10821);
or U11068 (N_11068,N_10873,N_10970);
nor U11069 (N_11069,N_10892,N_10932);
nor U11070 (N_11070,N_10802,N_10867);
nor U11071 (N_11071,N_10891,N_10920);
or U11072 (N_11072,N_10926,N_10866);
xor U11073 (N_11073,N_10915,N_10806);
and U11074 (N_11074,N_10994,N_10917);
nor U11075 (N_11075,N_10993,N_10887);
and U11076 (N_11076,N_10837,N_10979);
or U11077 (N_11077,N_10935,N_10987);
nand U11078 (N_11078,N_10972,N_10853);
nand U11079 (N_11079,N_10872,N_10835);
nor U11080 (N_11080,N_10877,N_10940);
or U11081 (N_11081,N_10929,N_10944);
and U11082 (N_11082,N_10952,N_10898);
xor U11083 (N_11083,N_10817,N_10904);
xor U11084 (N_11084,N_10854,N_10884);
nor U11085 (N_11085,N_10848,N_10976);
nand U11086 (N_11086,N_10808,N_10800);
nand U11087 (N_11087,N_10843,N_10907);
xnor U11088 (N_11088,N_10803,N_10807);
nor U11089 (N_11089,N_10833,N_10964);
and U11090 (N_11090,N_10928,N_10954);
or U11091 (N_11091,N_10978,N_10862);
and U11092 (N_11092,N_10933,N_10909);
and U11093 (N_11093,N_10962,N_10851);
xnor U11094 (N_11094,N_10946,N_10885);
xnor U11095 (N_11095,N_10878,N_10838);
xor U11096 (N_11096,N_10965,N_10830);
nor U11097 (N_11097,N_10842,N_10963);
or U11098 (N_11098,N_10864,N_10903);
nand U11099 (N_11099,N_10950,N_10916);
and U11100 (N_11100,N_10886,N_10968);
xnor U11101 (N_11101,N_10956,N_10959);
nor U11102 (N_11102,N_10807,N_10884);
nor U11103 (N_11103,N_10917,N_10974);
nand U11104 (N_11104,N_10917,N_10869);
or U11105 (N_11105,N_10967,N_10954);
xor U11106 (N_11106,N_10970,N_10871);
or U11107 (N_11107,N_10846,N_10885);
xnor U11108 (N_11108,N_10994,N_10860);
xnor U11109 (N_11109,N_10822,N_10942);
nand U11110 (N_11110,N_10926,N_10863);
nand U11111 (N_11111,N_10919,N_10864);
and U11112 (N_11112,N_10980,N_10940);
nor U11113 (N_11113,N_10960,N_10937);
or U11114 (N_11114,N_10815,N_10980);
and U11115 (N_11115,N_10964,N_10829);
and U11116 (N_11116,N_10951,N_10817);
and U11117 (N_11117,N_10994,N_10996);
nand U11118 (N_11118,N_10967,N_10955);
nor U11119 (N_11119,N_10991,N_10804);
nand U11120 (N_11120,N_10817,N_10912);
and U11121 (N_11121,N_10924,N_10897);
nor U11122 (N_11122,N_10958,N_10896);
and U11123 (N_11123,N_10977,N_10841);
and U11124 (N_11124,N_10923,N_10910);
nor U11125 (N_11125,N_10828,N_10860);
nor U11126 (N_11126,N_10967,N_10813);
and U11127 (N_11127,N_10950,N_10901);
nor U11128 (N_11128,N_10809,N_10845);
xor U11129 (N_11129,N_10968,N_10889);
or U11130 (N_11130,N_10924,N_10958);
or U11131 (N_11131,N_10995,N_10828);
nor U11132 (N_11132,N_10879,N_10903);
or U11133 (N_11133,N_10997,N_10908);
or U11134 (N_11134,N_10955,N_10985);
and U11135 (N_11135,N_10866,N_10861);
nand U11136 (N_11136,N_10811,N_10958);
or U11137 (N_11137,N_10936,N_10884);
xor U11138 (N_11138,N_10975,N_10833);
xor U11139 (N_11139,N_10964,N_10938);
xnor U11140 (N_11140,N_10925,N_10958);
or U11141 (N_11141,N_10903,N_10899);
nand U11142 (N_11142,N_10928,N_10933);
nand U11143 (N_11143,N_10995,N_10896);
and U11144 (N_11144,N_10824,N_10901);
or U11145 (N_11145,N_10801,N_10962);
or U11146 (N_11146,N_10993,N_10882);
or U11147 (N_11147,N_10881,N_10821);
nor U11148 (N_11148,N_10993,N_10862);
xnor U11149 (N_11149,N_10957,N_10856);
and U11150 (N_11150,N_10983,N_10925);
and U11151 (N_11151,N_10886,N_10920);
or U11152 (N_11152,N_10841,N_10835);
xnor U11153 (N_11153,N_10842,N_10993);
nor U11154 (N_11154,N_10833,N_10994);
nor U11155 (N_11155,N_10957,N_10854);
and U11156 (N_11156,N_10844,N_10840);
nor U11157 (N_11157,N_10857,N_10850);
nor U11158 (N_11158,N_10920,N_10814);
nor U11159 (N_11159,N_10959,N_10958);
or U11160 (N_11160,N_10802,N_10847);
nand U11161 (N_11161,N_10986,N_10825);
nor U11162 (N_11162,N_10927,N_10876);
and U11163 (N_11163,N_10831,N_10925);
or U11164 (N_11164,N_10956,N_10990);
nor U11165 (N_11165,N_10807,N_10808);
or U11166 (N_11166,N_10887,N_10858);
nand U11167 (N_11167,N_10886,N_10947);
nor U11168 (N_11168,N_10926,N_10859);
or U11169 (N_11169,N_10943,N_10986);
and U11170 (N_11170,N_10866,N_10893);
nand U11171 (N_11171,N_10919,N_10883);
or U11172 (N_11172,N_10898,N_10808);
nor U11173 (N_11173,N_10863,N_10886);
nand U11174 (N_11174,N_10979,N_10818);
nand U11175 (N_11175,N_10998,N_10876);
nor U11176 (N_11176,N_10953,N_10922);
xor U11177 (N_11177,N_10922,N_10936);
nand U11178 (N_11178,N_10923,N_10850);
nor U11179 (N_11179,N_10897,N_10886);
and U11180 (N_11180,N_10961,N_10839);
or U11181 (N_11181,N_10826,N_10983);
and U11182 (N_11182,N_10930,N_10894);
and U11183 (N_11183,N_10879,N_10821);
nor U11184 (N_11184,N_10828,N_10856);
xor U11185 (N_11185,N_10836,N_10961);
and U11186 (N_11186,N_10949,N_10950);
nor U11187 (N_11187,N_10923,N_10854);
or U11188 (N_11188,N_10907,N_10970);
xnor U11189 (N_11189,N_10955,N_10961);
xnor U11190 (N_11190,N_10869,N_10972);
xnor U11191 (N_11191,N_10986,N_10944);
or U11192 (N_11192,N_10833,N_10872);
nor U11193 (N_11193,N_10836,N_10857);
nand U11194 (N_11194,N_10840,N_10951);
and U11195 (N_11195,N_10983,N_10894);
xnor U11196 (N_11196,N_10842,N_10903);
nor U11197 (N_11197,N_10995,N_10998);
or U11198 (N_11198,N_10911,N_10844);
or U11199 (N_11199,N_10831,N_10899);
nor U11200 (N_11200,N_11077,N_11065);
or U11201 (N_11201,N_11022,N_11036);
or U11202 (N_11202,N_11106,N_11051);
or U11203 (N_11203,N_11026,N_11030);
nor U11204 (N_11204,N_11061,N_11156);
nor U11205 (N_11205,N_11098,N_11023);
and U11206 (N_11206,N_11064,N_11018);
and U11207 (N_11207,N_11148,N_11172);
nor U11208 (N_11208,N_11048,N_11021);
xor U11209 (N_11209,N_11181,N_11152);
nor U11210 (N_11210,N_11096,N_11121);
nor U11211 (N_11211,N_11076,N_11131);
nand U11212 (N_11212,N_11185,N_11058);
and U11213 (N_11213,N_11147,N_11078);
and U11214 (N_11214,N_11039,N_11145);
nor U11215 (N_11215,N_11006,N_11081);
and U11216 (N_11216,N_11128,N_11107);
or U11217 (N_11217,N_11103,N_11166);
nand U11218 (N_11218,N_11117,N_11001);
xor U11219 (N_11219,N_11045,N_11084);
nand U11220 (N_11220,N_11020,N_11151);
nor U11221 (N_11221,N_11071,N_11097);
nor U11222 (N_11222,N_11052,N_11146);
or U11223 (N_11223,N_11080,N_11126);
nand U11224 (N_11224,N_11004,N_11028);
or U11225 (N_11225,N_11090,N_11016);
or U11226 (N_11226,N_11118,N_11101);
nor U11227 (N_11227,N_11127,N_11113);
or U11228 (N_11228,N_11089,N_11184);
xor U11229 (N_11229,N_11025,N_11199);
nand U11230 (N_11230,N_11034,N_11136);
nor U11231 (N_11231,N_11179,N_11187);
xor U11232 (N_11232,N_11158,N_11150);
xor U11233 (N_11233,N_11019,N_11180);
or U11234 (N_11234,N_11057,N_11086);
and U11235 (N_11235,N_11153,N_11091);
and U11236 (N_11236,N_11056,N_11190);
nand U11237 (N_11237,N_11119,N_11130);
nand U11238 (N_11238,N_11196,N_11168);
and U11239 (N_11239,N_11124,N_11014);
and U11240 (N_11240,N_11099,N_11120);
xnor U11241 (N_11241,N_11161,N_11007);
and U11242 (N_11242,N_11157,N_11198);
and U11243 (N_11243,N_11109,N_11194);
nor U11244 (N_11244,N_11085,N_11108);
or U11245 (N_11245,N_11027,N_11040);
and U11246 (N_11246,N_11009,N_11188);
or U11247 (N_11247,N_11134,N_11002);
xnor U11248 (N_11248,N_11024,N_11060);
nor U11249 (N_11249,N_11195,N_11169);
or U11250 (N_11250,N_11160,N_11053);
nor U11251 (N_11251,N_11037,N_11178);
nor U11252 (N_11252,N_11093,N_11139);
and U11253 (N_11253,N_11186,N_11079);
and U11254 (N_11254,N_11137,N_11046);
nor U11255 (N_11255,N_11141,N_11059);
nor U11256 (N_11256,N_11092,N_11115);
xnor U11257 (N_11257,N_11133,N_11110);
nand U11258 (N_11258,N_11135,N_11069);
xnor U11259 (N_11259,N_11197,N_11149);
nor U11260 (N_11260,N_11100,N_11038);
or U11261 (N_11261,N_11042,N_11005);
or U11262 (N_11262,N_11155,N_11044);
or U11263 (N_11263,N_11050,N_11105);
nand U11264 (N_11264,N_11162,N_11174);
xnor U11265 (N_11265,N_11088,N_11144);
xor U11266 (N_11266,N_11003,N_11031);
and U11267 (N_11267,N_11191,N_11017);
and U11268 (N_11268,N_11011,N_11111);
and U11269 (N_11269,N_11125,N_11013);
and U11270 (N_11270,N_11192,N_11083);
nor U11271 (N_11271,N_11104,N_11123);
xor U11272 (N_11272,N_11182,N_11138);
nor U11273 (N_11273,N_11183,N_11033);
nand U11274 (N_11274,N_11072,N_11129);
nand U11275 (N_11275,N_11140,N_11068);
or U11276 (N_11276,N_11176,N_11012);
or U11277 (N_11277,N_11116,N_11102);
xnor U11278 (N_11278,N_11015,N_11122);
xnor U11279 (N_11279,N_11047,N_11189);
nor U11280 (N_11280,N_11043,N_11029);
nand U11281 (N_11281,N_11175,N_11055);
nor U11282 (N_11282,N_11067,N_11041);
xnor U11283 (N_11283,N_11054,N_11154);
nor U11284 (N_11284,N_11032,N_11143);
or U11285 (N_11285,N_11010,N_11193);
xnor U11286 (N_11286,N_11035,N_11177);
nor U11287 (N_11287,N_11171,N_11163);
and U11288 (N_11288,N_11087,N_11164);
and U11289 (N_11289,N_11062,N_11049);
nor U11290 (N_11290,N_11073,N_11112);
or U11291 (N_11291,N_11159,N_11114);
xnor U11292 (N_11292,N_11165,N_11094);
and U11293 (N_11293,N_11075,N_11142);
and U11294 (N_11294,N_11095,N_11167);
nor U11295 (N_11295,N_11063,N_11000);
xnor U11296 (N_11296,N_11170,N_11132);
xor U11297 (N_11297,N_11066,N_11008);
or U11298 (N_11298,N_11082,N_11074);
or U11299 (N_11299,N_11070,N_11173);
or U11300 (N_11300,N_11186,N_11194);
or U11301 (N_11301,N_11027,N_11051);
and U11302 (N_11302,N_11171,N_11013);
and U11303 (N_11303,N_11178,N_11005);
xnor U11304 (N_11304,N_11181,N_11025);
and U11305 (N_11305,N_11000,N_11120);
nor U11306 (N_11306,N_11013,N_11020);
nand U11307 (N_11307,N_11038,N_11171);
nor U11308 (N_11308,N_11105,N_11095);
nor U11309 (N_11309,N_11051,N_11020);
and U11310 (N_11310,N_11055,N_11015);
nor U11311 (N_11311,N_11084,N_11124);
nand U11312 (N_11312,N_11141,N_11183);
xnor U11313 (N_11313,N_11089,N_11136);
nand U11314 (N_11314,N_11197,N_11040);
nand U11315 (N_11315,N_11021,N_11162);
or U11316 (N_11316,N_11042,N_11017);
xnor U11317 (N_11317,N_11036,N_11066);
nand U11318 (N_11318,N_11073,N_11132);
nor U11319 (N_11319,N_11027,N_11165);
nand U11320 (N_11320,N_11181,N_11086);
and U11321 (N_11321,N_11136,N_11031);
and U11322 (N_11322,N_11043,N_11126);
nand U11323 (N_11323,N_11041,N_11161);
nor U11324 (N_11324,N_11063,N_11009);
and U11325 (N_11325,N_11009,N_11178);
or U11326 (N_11326,N_11040,N_11152);
nor U11327 (N_11327,N_11129,N_11163);
xor U11328 (N_11328,N_11072,N_11135);
xor U11329 (N_11329,N_11074,N_11025);
nor U11330 (N_11330,N_11188,N_11161);
nand U11331 (N_11331,N_11191,N_11147);
or U11332 (N_11332,N_11054,N_11151);
nand U11333 (N_11333,N_11087,N_11055);
or U11334 (N_11334,N_11069,N_11180);
and U11335 (N_11335,N_11005,N_11055);
xnor U11336 (N_11336,N_11123,N_11053);
nand U11337 (N_11337,N_11068,N_11035);
and U11338 (N_11338,N_11149,N_11073);
xnor U11339 (N_11339,N_11025,N_11147);
nor U11340 (N_11340,N_11003,N_11110);
xnor U11341 (N_11341,N_11012,N_11090);
xor U11342 (N_11342,N_11070,N_11130);
xor U11343 (N_11343,N_11054,N_11183);
nand U11344 (N_11344,N_11052,N_11171);
nor U11345 (N_11345,N_11041,N_11199);
and U11346 (N_11346,N_11058,N_11164);
or U11347 (N_11347,N_11126,N_11087);
or U11348 (N_11348,N_11008,N_11077);
nor U11349 (N_11349,N_11155,N_11025);
xor U11350 (N_11350,N_11035,N_11136);
or U11351 (N_11351,N_11193,N_11154);
nor U11352 (N_11352,N_11025,N_11095);
or U11353 (N_11353,N_11073,N_11038);
nor U11354 (N_11354,N_11101,N_11023);
nand U11355 (N_11355,N_11023,N_11163);
or U11356 (N_11356,N_11077,N_11086);
or U11357 (N_11357,N_11087,N_11149);
and U11358 (N_11358,N_11021,N_11146);
nand U11359 (N_11359,N_11188,N_11026);
nor U11360 (N_11360,N_11046,N_11009);
and U11361 (N_11361,N_11183,N_11199);
nor U11362 (N_11362,N_11127,N_11034);
xor U11363 (N_11363,N_11182,N_11145);
or U11364 (N_11364,N_11072,N_11145);
and U11365 (N_11365,N_11096,N_11024);
nor U11366 (N_11366,N_11032,N_11129);
nand U11367 (N_11367,N_11140,N_11046);
nand U11368 (N_11368,N_11023,N_11121);
or U11369 (N_11369,N_11155,N_11034);
nor U11370 (N_11370,N_11032,N_11106);
and U11371 (N_11371,N_11116,N_11064);
and U11372 (N_11372,N_11181,N_11083);
and U11373 (N_11373,N_11003,N_11152);
nor U11374 (N_11374,N_11080,N_11059);
or U11375 (N_11375,N_11073,N_11179);
xor U11376 (N_11376,N_11191,N_11068);
or U11377 (N_11377,N_11064,N_11143);
or U11378 (N_11378,N_11172,N_11083);
and U11379 (N_11379,N_11030,N_11172);
or U11380 (N_11380,N_11169,N_11052);
nor U11381 (N_11381,N_11046,N_11176);
nand U11382 (N_11382,N_11052,N_11090);
xor U11383 (N_11383,N_11075,N_11091);
xor U11384 (N_11384,N_11092,N_11061);
xnor U11385 (N_11385,N_11164,N_11024);
xnor U11386 (N_11386,N_11043,N_11196);
and U11387 (N_11387,N_11074,N_11024);
nor U11388 (N_11388,N_11068,N_11041);
nor U11389 (N_11389,N_11010,N_11186);
nor U11390 (N_11390,N_11054,N_11166);
or U11391 (N_11391,N_11125,N_11024);
or U11392 (N_11392,N_11092,N_11147);
nor U11393 (N_11393,N_11044,N_11160);
and U11394 (N_11394,N_11134,N_11108);
and U11395 (N_11395,N_11026,N_11160);
nor U11396 (N_11396,N_11071,N_11129);
xor U11397 (N_11397,N_11199,N_11071);
nor U11398 (N_11398,N_11147,N_11010);
or U11399 (N_11399,N_11020,N_11148);
xnor U11400 (N_11400,N_11347,N_11280);
nor U11401 (N_11401,N_11307,N_11265);
and U11402 (N_11402,N_11366,N_11261);
xor U11403 (N_11403,N_11335,N_11250);
xor U11404 (N_11404,N_11223,N_11201);
nand U11405 (N_11405,N_11383,N_11233);
or U11406 (N_11406,N_11288,N_11329);
or U11407 (N_11407,N_11282,N_11334);
and U11408 (N_11408,N_11306,N_11377);
nor U11409 (N_11409,N_11246,N_11369);
or U11410 (N_11410,N_11279,N_11331);
and U11411 (N_11411,N_11228,N_11296);
nand U11412 (N_11412,N_11337,N_11254);
nor U11413 (N_11413,N_11385,N_11338);
and U11414 (N_11414,N_11322,N_11248);
and U11415 (N_11415,N_11237,N_11242);
or U11416 (N_11416,N_11356,N_11325);
and U11417 (N_11417,N_11318,N_11283);
nor U11418 (N_11418,N_11263,N_11285);
xnor U11419 (N_11419,N_11372,N_11214);
xor U11420 (N_11420,N_11238,N_11308);
xor U11421 (N_11421,N_11274,N_11290);
nand U11422 (N_11422,N_11231,N_11204);
nand U11423 (N_11423,N_11346,N_11378);
xnor U11424 (N_11424,N_11361,N_11273);
and U11425 (N_11425,N_11235,N_11374);
xor U11426 (N_11426,N_11386,N_11368);
nor U11427 (N_11427,N_11312,N_11332);
nand U11428 (N_11428,N_11256,N_11216);
and U11429 (N_11429,N_11300,N_11303);
nand U11430 (N_11430,N_11375,N_11211);
nand U11431 (N_11431,N_11230,N_11328);
nand U11432 (N_11432,N_11222,N_11387);
and U11433 (N_11433,N_11269,N_11350);
nand U11434 (N_11434,N_11244,N_11252);
or U11435 (N_11435,N_11299,N_11394);
nor U11436 (N_11436,N_11349,N_11388);
nand U11437 (N_11437,N_11258,N_11260);
xor U11438 (N_11438,N_11357,N_11355);
nand U11439 (N_11439,N_11381,N_11240);
and U11440 (N_11440,N_11320,N_11391);
nand U11441 (N_11441,N_11339,N_11389);
or U11442 (N_11442,N_11321,N_11379);
nand U11443 (N_11443,N_11371,N_11207);
xor U11444 (N_11444,N_11373,N_11324);
or U11445 (N_11445,N_11259,N_11284);
or U11446 (N_11446,N_11390,N_11219);
nand U11447 (N_11447,N_11249,N_11293);
nand U11448 (N_11448,N_11313,N_11251);
or U11449 (N_11449,N_11370,N_11270);
or U11450 (N_11450,N_11205,N_11236);
or U11451 (N_11451,N_11212,N_11351);
nor U11452 (N_11452,N_11395,N_11227);
and U11453 (N_11453,N_11229,N_11363);
nor U11454 (N_11454,N_11327,N_11297);
nor U11455 (N_11455,N_11217,N_11317);
xnor U11456 (N_11456,N_11276,N_11315);
and U11457 (N_11457,N_11319,N_11243);
and U11458 (N_11458,N_11220,N_11336);
xor U11459 (N_11459,N_11267,N_11399);
or U11460 (N_11460,N_11342,N_11302);
or U11461 (N_11461,N_11365,N_11364);
nand U11462 (N_11462,N_11213,N_11310);
nand U11463 (N_11463,N_11330,N_11358);
and U11464 (N_11464,N_11239,N_11367);
or U11465 (N_11465,N_11396,N_11380);
or U11466 (N_11466,N_11354,N_11255);
or U11467 (N_11467,N_11289,N_11352);
or U11468 (N_11468,N_11295,N_11376);
or U11469 (N_11469,N_11304,N_11359);
and U11470 (N_11470,N_11215,N_11247);
xor U11471 (N_11471,N_11298,N_11275);
nand U11472 (N_11472,N_11266,N_11286);
nand U11473 (N_11473,N_11203,N_11262);
nor U11474 (N_11474,N_11221,N_11333);
and U11475 (N_11475,N_11323,N_11206);
nand U11476 (N_11476,N_11314,N_11292);
xor U11477 (N_11477,N_11344,N_11341);
or U11478 (N_11478,N_11208,N_11340);
nand U11479 (N_11479,N_11316,N_11362);
xnor U11480 (N_11480,N_11360,N_11278);
nor U11481 (N_11481,N_11305,N_11268);
or U11482 (N_11482,N_11253,N_11202);
nor U11483 (N_11483,N_11245,N_11345);
xor U11484 (N_11484,N_11209,N_11210);
or U11485 (N_11485,N_11200,N_11398);
nor U11486 (N_11486,N_11226,N_11225);
and U11487 (N_11487,N_11281,N_11392);
xnor U11488 (N_11488,N_11272,N_11287);
nand U11489 (N_11489,N_11382,N_11232);
or U11490 (N_11490,N_11353,N_11277);
and U11491 (N_11491,N_11271,N_11326);
or U11492 (N_11492,N_11311,N_11309);
nand U11493 (N_11493,N_11343,N_11301);
and U11494 (N_11494,N_11234,N_11241);
nor U11495 (N_11495,N_11224,N_11218);
nand U11496 (N_11496,N_11257,N_11291);
nand U11497 (N_11497,N_11294,N_11348);
nor U11498 (N_11498,N_11393,N_11397);
xnor U11499 (N_11499,N_11264,N_11384);
nor U11500 (N_11500,N_11320,N_11209);
nand U11501 (N_11501,N_11209,N_11280);
nand U11502 (N_11502,N_11394,N_11338);
and U11503 (N_11503,N_11299,N_11215);
nor U11504 (N_11504,N_11384,N_11346);
and U11505 (N_11505,N_11201,N_11393);
nand U11506 (N_11506,N_11382,N_11200);
or U11507 (N_11507,N_11203,N_11339);
xor U11508 (N_11508,N_11352,N_11375);
nand U11509 (N_11509,N_11242,N_11238);
or U11510 (N_11510,N_11384,N_11379);
xor U11511 (N_11511,N_11244,N_11259);
and U11512 (N_11512,N_11350,N_11349);
and U11513 (N_11513,N_11228,N_11274);
or U11514 (N_11514,N_11205,N_11370);
or U11515 (N_11515,N_11365,N_11293);
or U11516 (N_11516,N_11340,N_11310);
xor U11517 (N_11517,N_11357,N_11338);
xnor U11518 (N_11518,N_11339,N_11259);
nand U11519 (N_11519,N_11223,N_11248);
and U11520 (N_11520,N_11369,N_11200);
nand U11521 (N_11521,N_11340,N_11391);
and U11522 (N_11522,N_11228,N_11384);
or U11523 (N_11523,N_11370,N_11302);
xor U11524 (N_11524,N_11390,N_11381);
nor U11525 (N_11525,N_11383,N_11362);
or U11526 (N_11526,N_11370,N_11251);
nand U11527 (N_11527,N_11380,N_11214);
and U11528 (N_11528,N_11241,N_11316);
nor U11529 (N_11529,N_11339,N_11379);
or U11530 (N_11530,N_11383,N_11215);
nand U11531 (N_11531,N_11379,N_11375);
nor U11532 (N_11532,N_11289,N_11220);
xnor U11533 (N_11533,N_11204,N_11385);
and U11534 (N_11534,N_11294,N_11307);
and U11535 (N_11535,N_11201,N_11213);
and U11536 (N_11536,N_11218,N_11324);
xor U11537 (N_11537,N_11350,N_11265);
nor U11538 (N_11538,N_11269,N_11347);
nand U11539 (N_11539,N_11229,N_11218);
xnor U11540 (N_11540,N_11259,N_11367);
xor U11541 (N_11541,N_11270,N_11265);
nand U11542 (N_11542,N_11306,N_11320);
and U11543 (N_11543,N_11274,N_11310);
xor U11544 (N_11544,N_11213,N_11237);
or U11545 (N_11545,N_11238,N_11261);
and U11546 (N_11546,N_11254,N_11397);
or U11547 (N_11547,N_11319,N_11326);
nor U11548 (N_11548,N_11343,N_11250);
nand U11549 (N_11549,N_11290,N_11313);
and U11550 (N_11550,N_11397,N_11244);
nand U11551 (N_11551,N_11202,N_11307);
xor U11552 (N_11552,N_11350,N_11251);
or U11553 (N_11553,N_11268,N_11279);
nand U11554 (N_11554,N_11252,N_11220);
nand U11555 (N_11555,N_11374,N_11385);
nand U11556 (N_11556,N_11299,N_11283);
xnor U11557 (N_11557,N_11372,N_11361);
nor U11558 (N_11558,N_11262,N_11217);
xor U11559 (N_11559,N_11398,N_11341);
xnor U11560 (N_11560,N_11300,N_11365);
nand U11561 (N_11561,N_11244,N_11391);
nor U11562 (N_11562,N_11257,N_11246);
or U11563 (N_11563,N_11340,N_11362);
xnor U11564 (N_11564,N_11246,N_11309);
xor U11565 (N_11565,N_11320,N_11258);
or U11566 (N_11566,N_11223,N_11216);
and U11567 (N_11567,N_11317,N_11233);
nand U11568 (N_11568,N_11215,N_11228);
or U11569 (N_11569,N_11316,N_11389);
xnor U11570 (N_11570,N_11377,N_11200);
nand U11571 (N_11571,N_11245,N_11295);
xnor U11572 (N_11572,N_11379,N_11264);
xor U11573 (N_11573,N_11240,N_11242);
xnor U11574 (N_11574,N_11233,N_11273);
xnor U11575 (N_11575,N_11335,N_11219);
and U11576 (N_11576,N_11294,N_11389);
nor U11577 (N_11577,N_11227,N_11289);
nand U11578 (N_11578,N_11339,N_11320);
nand U11579 (N_11579,N_11295,N_11303);
nand U11580 (N_11580,N_11237,N_11218);
xnor U11581 (N_11581,N_11232,N_11356);
xnor U11582 (N_11582,N_11366,N_11285);
and U11583 (N_11583,N_11254,N_11317);
or U11584 (N_11584,N_11203,N_11382);
xnor U11585 (N_11585,N_11317,N_11271);
nor U11586 (N_11586,N_11344,N_11370);
nand U11587 (N_11587,N_11360,N_11307);
and U11588 (N_11588,N_11392,N_11275);
xnor U11589 (N_11589,N_11230,N_11218);
nand U11590 (N_11590,N_11333,N_11204);
nand U11591 (N_11591,N_11252,N_11371);
xnor U11592 (N_11592,N_11311,N_11374);
xnor U11593 (N_11593,N_11373,N_11229);
nand U11594 (N_11594,N_11308,N_11376);
nor U11595 (N_11595,N_11383,N_11367);
or U11596 (N_11596,N_11375,N_11393);
xor U11597 (N_11597,N_11310,N_11353);
nor U11598 (N_11598,N_11344,N_11202);
xor U11599 (N_11599,N_11379,N_11341);
nand U11600 (N_11600,N_11499,N_11494);
nand U11601 (N_11601,N_11532,N_11403);
nand U11602 (N_11602,N_11477,N_11470);
and U11603 (N_11603,N_11414,N_11581);
xor U11604 (N_11604,N_11540,N_11524);
nand U11605 (N_11605,N_11554,N_11510);
xnor U11606 (N_11606,N_11424,N_11575);
xor U11607 (N_11607,N_11522,N_11549);
nand U11608 (N_11608,N_11405,N_11415);
nand U11609 (N_11609,N_11421,N_11533);
nor U11610 (N_11610,N_11400,N_11488);
xor U11611 (N_11611,N_11482,N_11550);
xor U11612 (N_11612,N_11473,N_11465);
or U11613 (N_11613,N_11478,N_11570);
and U11614 (N_11614,N_11588,N_11489);
or U11615 (N_11615,N_11515,N_11481);
nor U11616 (N_11616,N_11485,N_11506);
nand U11617 (N_11617,N_11419,N_11483);
or U11618 (N_11618,N_11525,N_11541);
xnor U11619 (N_11619,N_11449,N_11546);
nor U11620 (N_11620,N_11571,N_11574);
or U11621 (N_11621,N_11437,N_11530);
and U11622 (N_11622,N_11544,N_11486);
or U11623 (N_11623,N_11531,N_11561);
and U11624 (N_11624,N_11517,N_11459);
xnor U11625 (N_11625,N_11504,N_11402);
nand U11626 (N_11626,N_11534,N_11568);
nand U11627 (N_11627,N_11591,N_11444);
xor U11628 (N_11628,N_11466,N_11420);
or U11629 (N_11629,N_11505,N_11468);
nor U11630 (N_11630,N_11422,N_11401);
and U11631 (N_11631,N_11440,N_11539);
xnor U11632 (N_11632,N_11586,N_11573);
nor U11633 (N_11633,N_11582,N_11427);
nand U11634 (N_11634,N_11527,N_11442);
or U11635 (N_11635,N_11460,N_11500);
nand U11636 (N_11636,N_11594,N_11455);
nor U11637 (N_11637,N_11454,N_11431);
xnor U11638 (N_11638,N_11491,N_11547);
and U11639 (N_11639,N_11543,N_11426);
or U11640 (N_11640,N_11425,N_11433);
or U11641 (N_11641,N_11452,N_11597);
nand U11642 (N_11642,N_11471,N_11556);
nand U11643 (N_11643,N_11560,N_11578);
or U11644 (N_11644,N_11520,N_11559);
xnor U11645 (N_11645,N_11404,N_11490);
and U11646 (N_11646,N_11448,N_11598);
nor U11647 (N_11647,N_11416,N_11567);
or U11648 (N_11648,N_11487,N_11406);
xnor U11649 (N_11649,N_11476,N_11495);
or U11650 (N_11650,N_11585,N_11479);
nor U11651 (N_11651,N_11469,N_11577);
xor U11652 (N_11652,N_11592,N_11595);
nand U11653 (N_11653,N_11423,N_11501);
xor U11654 (N_11654,N_11496,N_11445);
or U11655 (N_11655,N_11498,N_11456);
xnor U11656 (N_11656,N_11536,N_11587);
nor U11657 (N_11657,N_11518,N_11572);
and U11658 (N_11658,N_11590,N_11516);
and U11659 (N_11659,N_11474,N_11493);
nor U11660 (N_11660,N_11583,N_11432);
xnor U11661 (N_11661,N_11563,N_11472);
nand U11662 (N_11662,N_11410,N_11458);
or U11663 (N_11663,N_11438,N_11508);
nor U11664 (N_11664,N_11555,N_11565);
nand U11665 (N_11665,N_11509,N_11542);
xor U11666 (N_11666,N_11413,N_11464);
nor U11667 (N_11667,N_11519,N_11407);
and U11668 (N_11668,N_11521,N_11579);
and U11669 (N_11669,N_11580,N_11450);
and U11670 (N_11670,N_11523,N_11463);
or U11671 (N_11671,N_11439,N_11457);
or U11672 (N_11672,N_11441,N_11562);
and U11673 (N_11673,N_11511,N_11428);
nor U11674 (N_11674,N_11513,N_11553);
xnor U11675 (N_11675,N_11566,N_11453);
xor U11676 (N_11676,N_11412,N_11529);
xor U11677 (N_11677,N_11545,N_11502);
xnor U11678 (N_11678,N_11430,N_11484);
or U11679 (N_11679,N_11480,N_11557);
nand U11680 (N_11680,N_11507,N_11446);
nand U11681 (N_11681,N_11447,N_11564);
nand U11682 (N_11682,N_11552,N_11408);
nand U11683 (N_11683,N_11569,N_11451);
and U11684 (N_11684,N_11526,N_11548);
or U11685 (N_11685,N_11462,N_11435);
nor U11686 (N_11686,N_11558,N_11475);
xnor U11687 (N_11687,N_11512,N_11584);
or U11688 (N_11688,N_11497,N_11418);
nand U11689 (N_11689,N_11576,N_11411);
nor U11690 (N_11690,N_11537,N_11535);
nor U11691 (N_11691,N_11461,N_11599);
nor U11692 (N_11692,N_11596,N_11429);
nand U11693 (N_11693,N_11538,N_11492);
xnor U11694 (N_11694,N_11467,N_11514);
xor U11695 (N_11695,N_11589,N_11593);
and U11696 (N_11696,N_11551,N_11503);
xnor U11697 (N_11697,N_11417,N_11436);
xor U11698 (N_11698,N_11528,N_11434);
nor U11699 (N_11699,N_11443,N_11409);
or U11700 (N_11700,N_11496,N_11407);
nor U11701 (N_11701,N_11551,N_11457);
xnor U11702 (N_11702,N_11455,N_11528);
and U11703 (N_11703,N_11512,N_11402);
nor U11704 (N_11704,N_11413,N_11589);
nand U11705 (N_11705,N_11457,N_11441);
nand U11706 (N_11706,N_11535,N_11407);
nor U11707 (N_11707,N_11458,N_11594);
nand U11708 (N_11708,N_11490,N_11505);
nand U11709 (N_11709,N_11435,N_11524);
xor U11710 (N_11710,N_11595,N_11516);
or U11711 (N_11711,N_11492,N_11477);
nand U11712 (N_11712,N_11443,N_11583);
nor U11713 (N_11713,N_11484,N_11564);
or U11714 (N_11714,N_11584,N_11523);
xor U11715 (N_11715,N_11598,N_11465);
nor U11716 (N_11716,N_11512,N_11405);
and U11717 (N_11717,N_11598,N_11528);
or U11718 (N_11718,N_11566,N_11458);
and U11719 (N_11719,N_11419,N_11451);
nor U11720 (N_11720,N_11438,N_11466);
nand U11721 (N_11721,N_11583,N_11469);
nand U11722 (N_11722,N_11596,N_11403);
nor U11723 (N_11723,N_11495,N_11568);
xnor U11724 (N_11724,N_11573,N_11451);
or U11725 (N_11725,N_11552,N_11566);
nor U11726 (N_11726,N_11410,N_11446);
or U11727 (N_11727,N_11593,N_11425);
or U11728 (N_11728,N_11459,N_11511);
xor U11729 (N_11729,N_11528,N_11479);
or U11730 (N_11730,N_11533,N_11497);
nand U11731 (N_11731,N_11553,N_11469);
xor U11732 (N_11732,N_11443,N_11524);
and U11733 (N_11733,N_11577,N_11412);
nand U11734 (N_11734,N_11419,N_11431);
nand U11735 (N_11735,N_11516,N_11519);
or U11736 (N_11736,N_11552,N_11548);
or U11737 (N_11737,N_11463,N_11483);
nand U11738 (N_11738,N_11439,N_11508);
or U11739 (N_11739,N_11484,N_11533);
nor U11740 (N_11740,N_11478,N_11476);
or U11741 (N_11741,N_11564,N_11438);
nor U11742 (N_11742,N_11539,N_11430);
or U11743 (N_11743,N_11570,N_11466);
and U11744 (N_11744,N_11533,N_11510);
nand U11745 (N_11745,N_11405,N_11416);
nor U11746 (N_11746,N_11488,N_11535);
xnor U11747 (N_11747,N_11501,N_11594);
xnor U11748 (N_11748,N_11541,N_11476);
or U11749 (N_11749,N_11497,N_11542);
nor U11750 (N_11750,N_11449,N_11575);
and U11751 (N_11751,N_11426,N_11457);
nor U11752 (N_11752,N_11481,N_11595);
nor U11753 (N_11753,N_11476,N_11461);
and U11754 (N_11754,N_11537,N_11456);
xnor U11755 (N_11755,N_11413,N_11417);
xnor U11756 (N_11756,N_11477,N_11532);
or U11757 (N_11757,N_11527,N_11518);
nand U11758 (N_11758,N_11510,N_11468);
nand U11759 (N_11759,N_11583,N_11473);
nor U11760 (N_11760,N_11522,N_11493);
nor U11761 (N_11761,N_11448,N_11473);
nand U11762 (N_11762,N_11565,N_11571);
or U11763 (N_11763,N_11506,N_11574);
nand U11764 (N_11764,N_11428,N_11540);
and U11765 (N_11765,N_11504,N_11570);
xor U11766 (N_11766,N_11499,N_11501);
or U11767 (N_11767,N_11550,N_11539);
xor U11768 (N_11768,N_11587,N_11483);
xor U11769 (N_11769,N_11431,N_11571);
nand U11770 (N_11770,N_11553,N_11538);
xnor U11771 (N_11771,N_11562,N_11427);
nor U11772 (N_11772,N_11517,N_11536);
and U11773 (N_11773,N_11423,N_11559);
nor U11774 (N_11774,N_11509,N_11451);
or U11775 (N_11775,N_11407,N_11478);
xor U11776 (N_11776,N_11456,N_11552);
and U11777 (N_11777,N_11446,N_11574);
nand U11778 (N_11778,N_11450,N_11481);
and U11779 (N_11779,N_11576,N_11413);
nand U11780 (N_11780,N_11549,N_11561);
and U11781 (N_11781,N_11487,N_11556);
and U11782 (N_11782,N_11558,N_11515);
and U11783 (N_11783,N_11433,N_11415);
nand U11784 (N_11784,N_11559,N_11477);
xnor U11785 (N_11785,N_11508,N_11424);
or U11786 (N_11786,N_11591,N_11468);
nand U11787 (N_11787,N_11502,N_11596);
nor U11788 (N_11788,N_11531,N_11476);
xnor U11789 (N_11789,N_11439,N_11567);
and U11790 (N_11790,N_11584,N_11520);
xor U11791 (N_11791,N_11508,N_11422);
xor U11792 (N_11792,N_11597,N_11533);
nor U11793 (N_11793,N_11533,N_11424);
xor U11794 (N_11794,N_11553,N_11413);
nand U11795 (N_11795,N_11595,N_11494);
nor U11796 (N_11796,N_11416,N_11596);
nor U11797 (N_11797,N_11552,N_11430);
and U11798 (N_11798,N_11594,N_11461);
nor U11799 (N_11799,N_11582,N_11468);
and U11800 (N_11800,N_11749,N_11701);
nor U11801 (N_11801,N_11615,N_11774);
xor U11802 (N_11802,N_11628,N_11721);
and U11803 (N_11803,N_11799,N_11620);
nand U11804 (N_11804,N_11785,N_11736);
xnor U11805 (N_11805,N_11798,N_11662);
and U11806 (N_11806,N_11696,N_11626);
nor U11807 (N_11807,N_11748,N_11653);
nor U11808 (N_11808,N_11625,N_11663);
nand U11809 (N_11809,N_11641,N_11611);
nor U11810 (N_11810,N_11601,N_11673);
xnor U11811 (N_11811,N_11718,N_11649);
and U11812 (N_11812,N_11618,N_11691);
xor U11813 (N_11813,N_11672,N_11670);
nor U11814 (N_11814,N_11656,N_11660);
xnor U11815 (N_11815,N_11684,N_11766);
nor U11816 (N_11816,N_11737,N_11770);
nand U11817 (N_11817,N_11730,N_11768);
or U11818 (N_11818,N_11624,N_11747);
and U11819 (N_11819,N_11795,N_11610);
and U11820 (N_11820,N_11733,N_11723);
nand U11821 (N_11821,N_11681,N_11644);
or U11822 (N_11822,N_11778,N_11651);
nor U11823 (N_11823,N_11665,N_11658);
nand U11824 (N_11824,N_11762,N_11603);
nand U11825 (N_11825,N_11694,N_11609);
xnor U11826 (N_11826,N_11635,N_11607);
nor U11827 (N_11827,N_11765,N_11784);
or U11828 (N_11828,N_11771,N_11600);
nor U11829 (N_11829,N_11605,N_11753);
or U11830 (N_11830,N_11712,N_11621);
or U11831 (N_11831,N_11654,N_11752);
nand U11832 (N_11832,N_11783,N_11622);
or U11833 (N_11833,N_11743,N_11714);
nand U11834 (N_11834,N_11623,N_11698);
nor U11835 (N_11835,N_11773,N_11686);
and U11836 (N_11836,N_11751,N_11619);
nand U11837 (N_11837,N_11715,N_11614);
or U11838 (N_11838,N_11638,N_11728);
xor U11839 (N_11839,N_11627,N_11682);
nor U11840 (N_11840,N_11740,N_11708);
or U11841 (N_11841,N_11634,N_11772);
nor U11842 (N_11842,N_11727,N_11717);
or U11843 (N_11843,N_11674,N_11687);
nand U11844 (N_11844,N_11731,N_11685);
nand U11845 (N_11845,N_11713,N_11657);
and U11846 (N_11846,N_11790,N_11739);
and U11847 (N_11847,N_11667,N_11652);
or U11848 (N_11848,N_11629,N_11647);
nor U11849 (N_11849,N_11704,N_11763);
nand U11850 (N_11850,N_11631,N_11645);
and U11851 (N_11851,N_11756,N_11726);
nand U11852 (N_11852,N_11732,N_11659);
nor U11853 (N_11853,N_11767,N_11754);
or U11854 (N_11854,N_11705,N_11683);
or U11855 (N_11855,N_11604,N_11668);
and U11856 (N_11856,N_11745,N_11710);
nor U11857 (N_11857,N_11782,N_11760);
or U11858 (N_11858,N_11655,N_11786);
or U11859 (N_11859,N_11779,N_11664);
nor U11860 (N_11860,N_11676,N_11720);
nor U11861 (N_11861,N_11797,N_11702);
nand U11862 (N_11862,N_11688,N_11769);
and U11863 (N_11863,N_11725,N_11764);
nor U11864 (N_11864,N_11675,N_11792);
xnor U11865 (N_11865,N_11787,N_11690);
nor U11866 (N_11866,N_11613,N_11643);
nand U11867 (N_11867,N_11709,N_11716);
nand U11868 (N_11868,N_11793,N_11695);
or U11869 (N_11869,N_11679,N_11750);
xnor U11870 (N_11870,N_11780,N_11776);
nand U11871 (N_11871,N_11707,N_11666);
or U11872 (N_11872,N_11755,N_11757);
nand U11873 (N_11873,N_11616,N_11632);
and U11874 (N_11874,N_11630,N_11661);
and U11875 (N_11875,N_11692,N_11791);
and U11876 (N_11876,N_11648,N_11636);
or U11877 (N_11877,N_11608,N_11680);
nand U11878 (N_11878,N_11699,N_11724);
nor U11879 (N_11879,N_11788,N_11612);
nor U11880 (N_11880,N_11650,N_11642);
nand U11881 (N_11881,N_11678,N_11741);
nand U11882 (N_11882,N_11700,N_11775);
and U11883 (N_11883,N_11759,N_11734);
and U11884 (N_11884,N_11617,N_11639);
and U11885 (N_11885,N_11758,N_11719);
and U11886 (N_11886,N_11689,N_11633);
nor U11887 (N_11887,N_11746,N_11777);
or U11888 (N_11888,N_11693,N_11706);
or U11889 (N_11889,N_11671,N_11602);
or U11890 (N_11890,N_11637,N_11781);
or U11891 (N_11891,N_11703,N_11729);
nand U11892 (N_11892,N_11677,N_11796);
xor U11893 (N_11893,N_11742,N_11697);
nor U11894 (N_11894,N_11794,N_11606);
nand U11895 (N_11895,N_11669,N_11738);
nand U11896 (N_11896,N_11722,N_11744);
and U11897 (N_11897,N_11711,N_11789);
nand U11898 (N_11898,N_11735,N_11761);
xnor U11899 (N_11899,N_11646,N_11640);
xnor U11900 (N_11900,N_11654,N_11743);
nand U11901 (N_11901,N_11643,N_11690);
nor U11902 (N_11902,N_11655,N_11742);
nor U11903 (N_11903,N_11635,N_11638);
or U11904 (N_11904,N_11606,N_11662);
xnor U11905 (N_11905,N_11690,N_11634);
xnor U11906 (N_11906,N_11670,N_11637);
nand U11907 (N_11907,N_11615,N_11677);
and U11908 (N_11908,N_11795,N_11792);
nor U11909 (N_11909,N_11798,N_11778);
or U11910 (N_11910,N_11666,N_11646);
nor U11911 (N_11911,N_11610,N_11648);
xor U11912 (N_11912,N_11757,N_11751);
nor U11913 (N_11913,N_11631,N_11625);
and U11914 (N_11914,N_11617,N_11640);
nand U11915 (N_11915,N_11785,N_11739);
xor U11916 (N_11916,N_11753,N_11721);
and U11917 (N_11917,N_11752,N_11715);
nor U11918 (N_11918,N_11735,N_11673);
nand U11919 (N_11919,N_11750,N_11664);
or U11920 (N_11920,N_11714,N_11746);
and U11921 (N_11921,N_11706,N_11761);
or U11922 (N_11922,N_11779,N_11648);
and U11923 (N_11923,N_11675,N_11788);
nor U11924 (N_11924,N_11728,N_11712);
nor U11925 (N_11925,N_11669,N_11686);
nor U11926 (N_11926,N_11774,N_11633);
nand U11927 (N_11927,N_11704,N_11683);
and U11928 (N_11928,N_11656,N_11602);
nor U11929 (N_11929,N_11651,N_11698);
xnor U11930 (N_11930,N_11765,N_11797);
nand U11931 (N_11931,N_11766,N_11773);
or U11932 (N_11932,N_11748,N_11727);
xor U11933 (N_11933,N_11686,N_11713);
nor U11934 (N_11934,N_11779,N_11767);
or U11935 (N_11935,N_11773,N_11681);
and U11936 (N_11936,N_11722,N_11726);
and U11937 (N_11937,N_11747,N_11707);
and U11938 (N_11938,N_11788,N_11621);
and U11939 (N_11939,N_11753,N_11676);
or U11940 (N_11940,N_11701,N_11665);
and U11941 (N_11941,N_11724,N_11694);
nand U11942 (N_11942,N_11618,N_11740);
nor U11943 (N_11943,N_11613,N_11744);
nand U11944 (N_11944,N_11648,N_11658);
nand U11945 (N_11945,N_11679,N_11778);
xnor U11946 (N_11946,N_11713,N_11784);
or U11947 (N_11947,N_11629,N_11609);
nor U11948 (N_11948,N_11763,N_11780);
nor U11949 (N_11949,N_11647,N_11742);
nand U11950 (N_11950,N_11720,N_11642);
and U11951 (N_11951,N_11735,N_11639);
xnor U11952 (N_11952,N_11667,N_11794);
and U11953 (N_11953,N_11760,N_11626);
and U11954 (N_11954,N_11665,N_11789);
xor U11955 (N_11955,N_11622,N_11795);
xnor U11956 (N_11956,N_11769,N_11658);
nand U11957 (N_11957,N_11680,N_11715);
nor U11958 (N_11958,N_11743,N_11696);
xnor U11959 (N_11959,N_11707,N_11654);
nor U11960 (N_11960,N_11784,N_11741);
and U11961 (N_11961,N_11789,N_11784);
xnor U11962 (N_11962,N_11683,N_11719);
and U11963 (N_11963,N_11774,N_11693);
xor U11964 (N_11964,N_11636,N_11632);
nand U11965 (N_11965,N_11677,N_11726);
and U11966 (N_11966,N_11709,N_11724);
xor U11967 (N_11967,N_11723,N_11608);
and U11968 (N_11968,N_11607,N_11661);
and U11969 (N_11969,N_11630,N_11770);
or U11970 (N_11970,N_11795,N_11733);
or U11971 (N_11971,N_11675,N_11733);
nor U11972 (N_11972,N_11778,N_11661);
and U11973 (N_11973,N_11780,N_11636);
or U11974 (N_11974,N_11600,N_11680);
nor U11975 (N_11975,N_11614,N_11794);
nand U11976 (N_11976,N_11720,N_11643);
or U11977 (N_11977,N_11719,N_11665);
and U11978 (N_11978,N_11651,N_11603);
nor U11979 (N_11979,N_11740,N_11739);
nor U11980 (N_11980,N_11777,N_11726);
nand U11981 (N_11981,N_11660,N_11706);
or U11982 (N_11982,N_11770,N_11738);
nand U11983 (N_11983,N_11728,N_11737);
or U11984 (N_11984,N_11779,N_11606);
or U11985 (N_11985,N_11753,N_11671);
xnor U11986 (N_11986,N_11670,N_11786);
nor U11987 (N_11987,N_11749,N_11706);
nand U11988 (N_11988,N_11776,N_11772);
xor U11989 (N_11989,N_11677,N_11674);
xnor U11990 (N_11990,N_11778,N_11635);
xor U11991 (N_11991,N_11660,N_11662);
nor U11992 (N_11992,N_11702,N_11709);
or U11993 (N_11993,N_11681,N_11677);
xnor U11994 (N_11994,N_11611,N_11798);
and U11995 (N_11995,N_11758,N_11740);
or U11996 (N_11996,N_11656,N_11647);
nand U11997 (N_11997,N_11624,N_11686);
or U11998 (N_11998,N_11724,N_11784);
nand U11999 (N_11999,N_11612,N_11628);
nor U12000 (N_12000,N_11864,N_11886);
xor U12001 (N_12001,N_11917,N_11806);
nand U12002 (N_12002,N_11874,N_11908);
nor U12003 (N_12003,N_11941,N_11840);
and U12004 (N_12004,N_11932,N_11897);
and U12005 (N_12005,N_11924,N_11817);
or U12006 (N_12006,N_11851,N_11849);
xnor U12007 (N_12007,N_11947,N_11820);
xnor U12008 (N_12008,N_11831,N_11813);
nor U12009 (N_12009,N_11926,N_11828);
xor U12010 (N_12010,N_11920,N_11929);
nor U12011 (N_12011,N_11988,N_11890);
xor U12012 (N_12012,N_11974,N_11899);
xnor U12013 (N_12013,N_11962,N_11844);
and U12014 (N_12014,N_11855,N_11867);
and U12015 (N_12015,N_11933,N_11980);
xor U12016 (N_12016,N_11945,N_11959);
or U12017 (N_12017,N_11903,N_11937);
nor U12018 (N_12018,N_11948,N_11839);
nor U12019 (N_12019,N_11905,N_11868);
nor U12020 (N_12020,N_11989,N_11836);
xor U12021 (N_12021,N_11845,N_11990);
and U12022 (N_12022,N_11964,N_11860);
nand U12023 (N_12023,N_11846,N_11858);
and U12024 (N_12024,N_11803,N_11826);
nor U12025 (N_12025,N_11950,N_11808);
and U12026 (N_12026,N_11877,N_11812);
xor U12027 (N_12027,N_11983,N_11818);
nand U12028 (N_12028,N_11965,N_11979);
nor U12029 (N_12029,N_11879,N_11912);
and U12030 (N_12030,N_11958,N_11889);
nand U12031 (N_12031,N_11807,N_11862);
nor U12032 (N_12032,N_11935,N_11998);
or U12033 (N_12033,N_11943,N_11910);
or U12034 (N_12034,N_11859,N_11837);
nand U12035 (N_12035,N_11938,N_11916);
xor U12036 (N_12036,N_11982,N_11940);
xnor U12037 (N_12037,N_11829,N_11825);
xnor U12038 (N_12038,N_11966,N_11819);
and U12039 (N_12039,N_11995,N_11892);
nor U12040 (N_12040,N_11913,N_11880);
nor U12041 (N_12041,N_11805,N_11976);
and U12042 (N_12042,N_11883,N_11885);
or U12043 (N_12043,N_11878,N_11971);
xnor U12044 (N_12044,N_11814,N_11918);
nor U12045 (N_12045,N_11848,N_11978);
and U12046 (N_12046,N_11866,N_11810);
nor U12047 (N_12047,N_11884,N_11875);
nor U12048 (N_12048,N_11843,N_11835);
or U12049 (N_12049,N_11833,N_11972);
nor U12050 (N_12050,N_11949,N_11800);
and U12051 (N_12051,N_11994,N_11816);
nor U12052 (N_12052,N_11987,N_11975);
nor U12053 (N_12053,N_11985,N_11928);
xnor U12054 (N_12054,N_11871,N_11991);
or U12055 (N_12055,N_11847,N_11857);
nor U12056 (N_12056,N_11952,N_11852);
or U12057 (N_12057,N_11997,N_11901);
and U12058 (N_12058,N_11919,N_11863);
xor U12059 (N_12059,N_11931,N_11973);
and U12060 (N_12060,N_11834,N_11838);
and U12061 (N_12061,N_11832,N_11930);
xnor U12062 (N_12062,N_11873,N_11856);
or U12063 (N_12063,N_11957,N_11977);
and U12064 (N_12064,N_11893,N_11921);
xor U12065 (N_12065,N_11969,N_11954);
xnor U12066 (N_12066,N_11984,N_11904);
nand U12067 (N_12067,N_11895,N_11865);
or U12068 (N_12068,N_11992,N_11922);
xnor U12069 (N_12069,N_11881,N_11955);
nor U12070 (N_12070,N_11996,N_11967);
and U12071 (N_12071,N_11861,N_11809);
nor U12072 (N_12072,N_11815,N_11927);
nor U12073 (N_12073,N_11827,N_11824);
nand U12074 (N_12074,N_11934,N_11801);
nor U12075 (N_12075,N_11963,N_11970);
xor U12076 (N_12076,N_11870,N_11909);
or U12077 (N_12077,N_11999,N_11906);
nor U12078 (N_12078,N_11986,N_11936);
and U12079 (N_12079,N_11894,N_11821);
nand U12080 (N_12080,N_11902,N_11915);
nand U12081 (N_12081,N_11946,N_11842);
nand U12082 (N_12082,N_11898,N_11968);
xnor U12083 (N_12083,N_11888,N_11939);
or U12084 (N_12084,N_11853,N_11914);
and U12085 (N_12085,N_11956,N_11896);
xor U12086 (N_12086,N_11811,N_11802);
and U12087 (N_12087,N_11961,N_11882);
nor U12088 (N_12088,N_11854,N_11953);
nand U12089 (N_12089,N_11900,N_11925);
or U12090 (N_12090,N_11960,N_11923);
nand U12091 (N_12091,N_11876,N_11823);
and U12092 (N_12092,N_11981,N_11822);
or U12093 (N_12093,N_11804,N_11944);
or U12094 (N_12094,N_11907,N_11993);
xnor U12095 (N_12095,N_11891,N_11872);
xnor U12096 (N_12096,N_11911,N_11869);
nor U12097 (N_12097,N_11841,N_11850);
nor U12098 (N_12098,N_11887,N_11830);
xnor U12099 (N_12099,N_11942,N_11951);
or U12100 (N_12100,N_11974,N_11956);
nor U12101 (N_12101,N_11907,N_11991);
or U12102 (N_12102,N_11802,N_11963);
nand U12103 (N_12103,N_11832,N_11855);
and U12104 (N_12104,N_11928,N_11810);
or U12105 (N_12105,N_11996,N_11813);
and U12106 (N_12106,N_11978,N_11823);
nand U12107 (N_12107,N_11828,N_11996);
and U12108 (N_12108,N_11983,N_11948);
nand U12109 (N_12109,N_11943,N_11963);
nor U12110 (N_12110,N_11882,N_11993);
and U12111 (N_12111,N_11973,N_11831);
and U12112 (N_12112,N_11848,N_11833);
and U12113 (N_12113,N_11919,N_11839);
and U12114 (N_12114,N_11849,N_11861);
or U12115 (N_12115,N_11854,N_11832);
nor U12116 (N_12116,N_11914,N_11888);
and U12117 (N_12117,N_11952,N_11853);
or U12118 (N_12118,N_11996,N_11809);
xnor U12119 (N_12119,N_11802,N_11858);
xor U12120 (N_12120,N_11989,N_11930);
nand U12121 (N_12121,N_11825,N_11862);
or U12122 (N_12122,N_11813,N_11927);
nor U12123 (N_12123,N_11950,N_11937);
or U12124 (N_12124,N_11941,N_11928);
or U12125 (N_12125,N_11992,N_11902);
xnor U12126 (N_12126,N_11996,N_11979);
or U12127 (N_12127,N_11882,N_11922);
and U12128 (N_12128,N_11944,N_11818);
nor U12129 (N_12129,N_11941,N_11938);
xnor U12130 (N_12130,N_11853,N_11962);
nor U12131 (N_12131,N_11926,N_11813);
or U12132 (N_12132,N_11804,N_11852);
and U12133 (N_12133,N_11928,N_11822);
or U12134 (N_12134,N_11947,N_11883);
and U12135 (N_12135,N_11932,N_11849);
nor U12136 (N_12136,N_11867,N_11896);
xor U12137 (N_12137,N_11934,N_11933);
xor U12138 (N_12138,N_11922,N_11997);
nor U12139 (N_12139,N_11861,N_11911);
nand U12140 (N_12140,N_11825,N_11952);
and U12141 (N_12141,N_11876,N_11956);
nor U12142 (N_12142,N_11960,N_11823);
xnor U12143 (N_12143,N_11978,N_11961);
or U12144 (N_12144,N_11952,N_11996);
or U12145 (N_12145,N_11874,N_11881);
nor U12146 (N_12146,N_11912,N_11826);
or U12147 (N_12147,N_11970,N_11894);
or U12148 (N_12148,N_11898,N_11919);
nor U12149 (N_12149,N_11856,N_11928);
xor U12150 (N_12150,N_11974,N_11811);
xor U12151 (N_12151,N_11896,N_11962);
nand U12152 (N_12152,N_11968,N_11828);
or U12153 (N_12153,N_11946,N_11921);
nand U12154 (N_12154,N_11882,N_11865);
and U12155 (N_12155,N_11951,N_11929);
nand U12156 (N_12156,N_11900,N_11837);
and U12157 (N_12157,N_11959,N_11871);
and U12158 (N_12158,N_11878,N_11943);
nand U12159 (N_12159,N_11989,N_11962);
xor U12160 (N_12160,N_11822,N_11983);
nand U12161 (N_12161,N_11811,N_11971);
or U12162 (N_12162,N_11886,N_11815);
nor U12163 (N_12163,N_11844,N_11863);
nor U12164 (N_12164,N_11808,N_11812);
nand U12165 (N_12165,N_11960,N_11940);
or U12166 (N_12166,N_11964,N_11869);
xnor U12167 (N_12167,N_11968,N_11925);
nand U12168 (N_12168,N_11838,N_11821);
or U12169 (N_12169,N_11980,N_11849);
or U12170 (N_12170,N_11833,N_11805);
or U12171 (N_12171,N_11899,N_11819);
nor U12172 (N_12172,N_11822,N_11952);
and U12173 (N_12173,N_11838,N_11968);
xor U12174 (N_12174,N_11907,N_11910);
or U12175 (N_12175,N_11949,N_11950);
or U12176 (N_12176,N_11826,N_11973);
nor U12177 (N_12177,N_11851,N_11942);
and U12178 (N_12178,N_11819,N_11852);
nand U12179 (N_12179,N_11918,N_11838);
nor U12180 (N_12180,N_11864,N_11942);
and U12181 (N_12181,N_11932,N_11804);
nand U12182 (N_12182,N_11810,N_11830);
nand U12183 (N_12183,N_11998,N_11804);
or U12184 (N_12184,N_11935,N_11864);
xor U12185 (N_12185,N_11804,N_11848);
nor U12186 (N_12186,N_11946,N_11848);
or U12187 (N_12187,N_11974,N_11880);
nand U12188 (N_12188,N_11846,N_11986);
xnor U12189 (N_12189,N_11990,N_11957);
or U12190 (N_12190,N_11835,N_11825);
nand U12191 (N_12191,N_11966,N_11892);
nand U12192 (N_12192,N_11872,N_11934);
xnor U12193 (N_12193,N_11846,N_11955);
or U12194 (N_12194,N_11887,N_11915);
and U12195 (N_12195,N_11844,N_11819);
or U12196 (N_12196,N_11900,N_11885);
and U12197 (N_12197,N_11892,N_11853);
or U12198 (N_12198,N_11998,N_11809);
and U12199 (N_12199,N_11976,N_11973);
xnor U12200 (N_12200,N_12192,N_12182);
and U12201 (N_12201,N_12093,N_12042);
nand U12202 (N_12202,N_12024,N_12161);
nor U12203 (N_12203,N_12012,N_12013);
or U12204 (N_12204,N_12140,N_12098);
nand U12205 (N_12205,N_12178,N_12084);
xor U12206 (N_12206,N_12145,N_12076);
and U12207 (N_12207,N_12194,N_12100);
or U12208 (N_12208,N_12168,N_12048);
and U12209 (N_12209,N_12169,N_12191);
or U12210 (N_12210,N_12156,N_12111);
or U12211 (N_12211,N_12125,N_12190);
nor U12212 (N_12212,N_12027,N_12081);
nand U12213 (N_12213,N_12059,N_12108);
or U12214 (N_12214,N_12018,N_12011);
and U12215 (N_12215,N_12044,N_12116);
nand U12216 (N_12216,N_12133,N_12109);
nor U12217 (N_12217,N_12001,N_12032);
and U12218 (N_12218,N_12034,N_12175);
and U12219 (N_12219,N_12056,N_12157);
or U12220 (N_12220,N_12086,N_12113);
nor U12221 (N_12221,N_12138,N_12083);
and U12222 (N_12222,N_12047,N_12104);
xor U12223 (N_12223,N_12030,N_12170);
and U12224 (N_12224,N_12160,N_12126);
nor U12225 (N_12225,N_12000,N_12110);
and U12226 (N_12226,N_12091,N_12071);
and U12227 (N_12227,N_12015,N_12054);
nand U12228 (N_12228,N_12118,N_12065);
nand U12229 (N_12229,N_12005,N_12082);
and U12230 (N_12230,N_12007,N_12112);
nor U12231 (N_12231,N_12151,N_12099);
xor U12232 (N_12232,N_12102,N_12080);
nand U12233 (N_12233,N_12185,N_12119);
and U12234 (N_12234,N_12193,N_12021);
or U12235 (N_12235,N_12003,N_12010);
nand U12236 (N_12236,N_12107,N_12051);
or U12237 (N_12237,N_12096,N_12198);
and U12238 (N_12238,N_12045,N_12006);
nor U12239 (N_12239,N_12094,N_12130);
nor U12240 (N_12240,N_12022,N_12167);
or U12241 (N_12241,N_12124,N_12199);
nand U12242 (N_12242,N_12123,N_12017);
nor U12243 (N_12243,N_12163,N_12055);
nand U12244 (N_12244,N_12074,N_12152);
xor U12245 (N_12245,N_12149,N_12014);
and U12246 (N_12246,N_12155,N_12035);
nor U12247 (N_12247,N_12064,N_12128);
and U12248 (N_12248,N_12101,N_12088);
nand U12249 (N_12249,N_12079,N_12127);
and U12250 (N_12250,N_12066,N_12136);
or U12251 (N_12251,N_12115,N_12186);
and U12252 (N_12252,N_12176,N_12172);
or U12253 (N_12253,N_12154,N_12179);
nand U12254 (N_12254,N_12144,N_12039);
xor U12255 (N_12255,N_12016,N_12050);
nor U12256 (N_12256,N_12180,N_12078);
or U12257 (N_12257,N_12070,N_12135);
nand U12258 (N_12258,N_12106,N_12117);
xnor U12259 (N_12259,N_12103,N_12146);
nor U12260 (N_12260,N_12060,N_12142);
xnor U12261 (N_12261,N_12114,N_12129);
xnor U12262 (N_12262,N_12026,N_12025);
or U12263 (N_12263,N_12147,N_12038);
nor U12264 (N_12264,N_12037,N_12073);
or U12265 (N_12265,N_12077,N_12004);
nand U12266 (N_12266,N_12177,N_12046);
nor U12267 (N_12267,N_12150,N_12183);
xnor U12268 (N_12268,N_12195,N_12033);
or U12269 (N_12269,N_12139,N_12087);
or U12270 (N_12270,N_12181,N_12019);
and U12271 (N_12271,N_12062,N_12174);
xnor U12272 (N_12272,N_12008,N_12159);
xor U12273 (N_12273,N_12072,N_12075);
xnor U12274 (N_12274,N_12092,N_12188);
xor U12275 (N_12275,N_12061,N_12189);
or U12276 (N_12276,N_12120,N_12097);
nand U12277 (N_12277,N_12153,N_12041);
or U12278 (N_12278,N_12009,N_12067);
and U12279 (N_12279,N_12095,N_12052);
nand U12280 (N_12280,N_12069,N_12029);
xnor U12281 (N_12281,N_12141,N_12057);
nand U12282 (N_12282,N_12187,N_12162);
nand U12283 (N_12283,N_12132,N_12121);
or U12284 (N_12284,N_12173,N_12184);
nand U12285 (N_12285,N_12040,N_12143);
and U12286 (N_12286,N_12197,N_12166);
or U12287 (N_12287,N_12063,N_12028);
xnor U12288 (N_12288,N_12137,N_12089);
xnor U12289 (N_12289,N_12122,N_12134);
and U12290 (N_12290,N_12068,N_12164);
nor U12291 (N_12291,N_12058,N_12085);
or U12292 (N_12292,N_12196,N_12036);
nand U12293 (N_12293,N_12090,N_12165);
nor U12294 (N_12294,N_12023,N_12148);
or U12295 (N_12295,N_12049,N_12020);
nand U12296 (N_12296,N_12105,N_12043);
xnor U12297 (N_12297,N_12031,N_12131);
nor U12298 (N_12298,N_12158,N_12053);
or U12299 (N_12299,N_12171,N_12002);
nor U12300 (N_12300,N_12097,N_12125);
and U12301 (N_12301,N_12004,N_12089);
or U12302 (N_12302,N_12097,N_12021);
xnor U12303 (N_12303,N_12077,N_12013);
nor U12304 (N_12304,N_12017,N_12193);
or U12305 (N_12305,N_12115,N_12036);
nand U12306 (N_12306,N_12153,N_12098);
xor U12307 (N_12307,N_12066,N_12006);
or U12308 (N_12308,N_12142,N_12084);
or U12309 (N_12309,N_12159,N_12152);
and U12310 (N_12310,N_12031,N_12066);
nor U12311 (N_12311,N_12150,N_12040);
and U12312 (N_12312,N_12196,N_12017);
xor U12313 (N_12313,N_12036,N_12027);
nand U12314 (N_12314,N_12014,N_12039);
and U12315 (N_12315,N_12032,N_12107);
and U12316 (N_12316,N_12145,N_12040);
nor U12317 (N_12317,N_12009,N_12134);
nand U12318 (N_12318,N_12085,N_12038);
or U12319 (N_12319,N_12074,N_12016);
or U12320 (N_12320,N_12173,N_12099);
nor U12321 (N_12321,N_12164,N_12044);
nand U12322 (N_12322,N_12163,N_12192);
xor U12323 (N_12323,N_12090,N_12068);
and U12324 (N_12324,N_12131,N_12156);
xnor U12325 (N_12325,N_12125,N_12130);
or U12326 (N_12326,N_12068,N_12190);
nand U12327 (N_12327,N_12099,N_12181);
or U12328 (N_12328,N_12152,N_12008);
and U12329 (N_12329,N_12070,N_12090);
or U12330 (N_12330,N_12016,N_12022);
or U12331 (N_12331,N_12017,N_12045);
or U12332 (N_12332,N_12159,N_12029);
nor U12333 (N_12333,N_12007,N_12122);
and U12334 (N_12334,N_12115,N_12183);
nor U12335 (N_12335,N_12168,N_12020);
xnor U12336 (N_12336,N_12055,N_12082);
nor U12337 (N_12337,N_12136,N_12032);
or U12338 (N_12338,N_12129,N_12107);
nand U12339 (N_12339,N_12164,N_12119);
nor U12340 (N_12340,N_12115,N_12177);
or U12341 (N_12341,N_12096,N_12032);
nand U12342 (N_12342,N_12103,N_12139);
nand U12343 (N_12343,N_12055,N_12136);
or U12344 (N_12344,N_12035,N_12128);
or U12345 (N_12345,N_12006,N_12069);
or U12346 (N_12346,N_12105,N_12009);
nand U12347 (N_12347,N_12079,N_12014);
xnor U12348 (N_12348,N_12069,N_12158);
and U12349 (N_12349,N_12187,N_12148);
nand U12350 (N_12350,N_12151,N_12049);
nor U12351 (N_12351,N_12197,N_12091);
and U12352 (N_12352,N_12056,N_12072);
or U12353 (N_12353,N_12089,N_12027);
nand U12354 (N_12354,N_12125,N_12128);
and U12355 (N_12355,N_12038,N_12032);
xnor U12356 (N_12356,N_12095,N_12067);
xor U12357 (N_12357,N_12177,N_12194);
nand U12358 (N_12358,N_12116,N_12163);
nor U12359 (N_12359,N_12154,N_12137);
or U12360 (N_12360,N_12150,N_12076);
or U12361 (N_12361,N_12148,N_12176);
and U12362 (N_12362,N_12168,N_12166);
or U12363 (N_12363,N_12175,N_12170);
or U12364 (N_12364,N_12050,N_12147);
nand U12365 (N_12365,N_12085,N_12159);
nor U12366 (N_12366,N_12058,N_12046);
nor U12367 (N_12367,N_12076,N_12102);
xor U12368 (N_12368,N_12016,N_12189);
nor U12369 (N_12369,N_12128,N_12111);
xor U12370 (N_12370,N_12077,N_12164);
xnor U12371 (N_12371,N_12199,N_12185);
xor U12372 (N_12372,N_12015,N_12055);
and U12373 (N_12373,N_12082,N_12196);
nor U12374 (N_12374,N_12158,N_12102);
xnor U12375 (N_12375,N_12011,N_12159);
and U12376 (N_12376,N_12100,N_12064);
nand U12377 (N_12377,N_12191,N_12022);
nand U12378 (N_12378,N_12171,N_12144);
nand U12379 (N_12379,N_12010,N_12173);
or U12380 (N_12380,N_12093,N_12065);
and U12381 (N_12381,N_12146,N_12099);
xnor U12382 (N_12382,N_12135,N_12195);
xor U12383 (N_12383,N_12037,N_12194);
or U12384 (N_12384,N_12035,N_12070);
nor U12385 (N_12385,N_12152,N_12168);
or U12386 (N_12386,N_12146,N_12046);
nand U12387 (N_12387,N_12176,N_12013);
nand U12388 (N_12388,N_12051,N_12019);
xor U12389 (N_12389,N_12006,N_12084);
and U12390 (N_12390,N_12007,N_12188);
nor U12391 (N_12391,N_12045,N_12186);
xor U12392 (N_12392,N_12177,N_12118);
xnor U12393 (N_12393,N_12029,N_12030);
nor U12394 (N_12394,N_12097,N_12157);
nand U12395 (N_12395,N_12050,N_12068);
or U12396 (N_12396,N_12181,N_12198);
xor U12397 (N_12397,N_12130,N_12085);
and U12398 (N_12398,N_12135,N_12069);
xor U12399 (N_12399,N_12053,N_12104);
nor U12400 (N_12400,N_12358,N_12287);
and U12401 (N_12401,N_12316,N_12261);
or U12402 (N_12402,N_12298,N_12228);
or U12403 (N_12403,N_12279,N_12259);
nand U12404 (N_12404,N_12224,N_12368);
nor U12405 (N_12405,N_12321,N_12348);
nand U12406 (N_12406,N_12255,N_12380);
xor U12407 (N_12407,N_12375,N_12285);
xor U12408 (N_12408,N_12342,N_12339);
or U12409 (N_12409,N_12341,N_12208);
and U12410 (N_12410,N_12349,N_12294);
and U12411 (N_12411,N_12314,N_12374);
nand U12412 (N_12412,N_12300,N_12328);
nor U12413 (N_12413,N_12258,N_12383);
or U12414 (N_12414,N_12264,N_12276);
nand U12415 (N_12415,N_12325,N_12360);
and U12416 (N_12416,N_12397,N_12211);
or U12417 (N_12417,N_12290,N_12332);
nand U12418 (N_12418,N_12233,N_12366);
xnor U12419 (N_12419,N_12256,N_12353);
and U12420 (N_12420,N_12393,N_12371);
nand U12421 (N_12421,N_12370,N_12334);
nand U12422 (N_12422,N_12241,N_12356);
or U12423 (N_12423,N_12372,N_12230);
and U12424 (N_12424,N_12311,N_12379);
or U12425 (N_12425,N_12203,N_12364);
and U12426 (N_12426,N_12308,N_12257);
xnor U12427 (N_12427,N_12326,N_12369);
nand U12428 (N_12428,N_12317,N_12340);
nand U12429 (N_12429,N_12347,N_12283);
or U12430 (N_12430,N_12204,N_12363);
xor U12431 (N_12431,N_12329,N_12267);
nand U12432 (N_12432,N_12221,N_12333);
and U12433 (N_12433,N_12337,N_12307);
nand U12434 (N_12434,N_12253,N_12205);
nor U12435 (N_12435,N_12206,N_12274);
nor U12436 (N_12436,N_12207,N_12319);
nor U12437 (N_12437,N_12273,N_12249);
nor U12438 (N_12438,N_12373,N_12216);
nor U12439 (N_12439,N_12245,N_12306);
and U12440 (N_12440,N_12376,N_12244);
and U12441 (N_12441,N_12362,N_12323);
and U12442 (N_12442,N_12243,N_12234);
or U12443 (N_12443,N_12262,N_12248);
nor U12444 (N_12444,N_12335,N_12266);
nand U12445 (N_12445,N_12247,N_12275);
nand U12446 (N_12446,N_12202,N_12301);
nand U12447 (N_12447,N_12215,N_12304);
or U12448 (N_12448,N_12312,N_12214);
xnor U12449 (N_12449,N_12390,N_12354);
or U12450 (N_12450,N_12310,N_12392);
and U12451 (N_12451,N_12291,N_12303);
nor U12452 (N_12452,N_12269,N_12394);
nand U12453 (N_12453,N_12263,N_12239);
nand U12454 (N_12454,N_12280,N_12391);
nand U12455 (N_12455,N_12336,N_12254);
nand U12456 (N_12456,N_12265,N_12399);
nand U12457 (N_12457,N_12386,N_12223);
nand U12458 (N_12458,N_12252,N_12227);
nand U12459 (N_12459,N_12331,N_12351);
nor U12460 (N_12460,N_12213,N_12309);
nor U12461 (N_12461,N_12367,N_12271);
and U12462 (N_12462,N_12286,N_12246);
nand U12463 (N_12463,N_12382,N_12289);
nor U12464 (N_12464,N_12250,N_12299);
and U12465 (N_12465,N_12365,N_12388);
or U12466 (N_12466,N_12218,N_12377);
and U12467 (N_12467,N_12352,N_12219);
nand U12468 (N_12468,N_12229,N_12357);
and U12469 (N_12469,N_12209,N_12385);
and U12470 (N_12470,N_12315,N_12355);
xor U12471 (N_12471,N_12200,N_12361);
or U12472 (N_12472,N_12201,N_12330);
and U12473 (N_12473,N_12359,N_12378);
or U12474 (N_12474,N_12389,N_12231);
xnor U12475 (N_12475,N_12384,N_12345);
xnor U12476 (N_12476,N_12350,N_12292);
or U12477 (N_12477,N_12346,N_12270);
xnor U12478 (N_12478,N_12284,N_12235);
or U12479 (N_12479,N_12281,N_12322);
and U12480 (N_12480,N_12305,N_12288);
or U12481 (N_12481,N_12225,N_12242);
and U12482 (N_12482,N_12327,N_12295);
nand U12483 (N_12483,N_12268,N_12220);
and U12484 (N_12484,N_12237,N_12297);
nand U12485 (N_12485,N_12344,N_12296);
nor U12486 (N_12486,N_12396,N_12251);
nor U12487 (N_12487,N_12210,N_12232);
nor U12488 (N_12488,N_12212,N_12238);
and U12489 (N_12489,N_12338,N_12236);
or U12490 (N_12490,N_12320,N_12381);
nand U12491 (N_12491,N_12217,N_12226);
nor U12492 (N_12492,N_12222,N_12272);
and U12493 (N_12493,N_12277,N_12278);
nand U12494 (N_12494,N_12324,N_12282);
or U12495 (N_12495,N_12240,N_12343);
and U12496 (N_12496,N_12395,N_12318);
nor U12497 (N_12497,N_12302,N_12260);
or U12498 (N_12498,N_12398,N_12387);
or U12499 (N_12499,N_12313,N_12293);
and U12500 (N_12500,N_12336,N_12253);
nor U12501 (N_12501,N_12209,N_12301);
or U12502 (N_12502,N_12371,N_12215);
nand U12503 (N_12503,N_12338,N_12330);
xnor U12504 (N_12504,N_12301,N_12314);
or U12505 (N_12505,N_12386,N_12299);
nor U12506 (N_12506,N_12301,N_12357);
xnor U12507 (N_12507,N_12369,N_12230);
and U12508 (N_12508,N_12286,N_12369);
or U12509 (N_12509,N_12304,N_12240);
nor U12510 (N_12510,N_12333,N_12283);
and U12511 (N_12511,N_12301,N_12210);
nor U12512 (N_12512,N_12241,N_12251);
and U12513 (N_12513,N_12355,N_12275);
and U12514 (N_12514,N_12297,N_12338);
and U12515 (N_12515,N_12205,N_12393);
nand U12516 (N_12516,N_12339,N_12373);
and U12517 (N_12517,N_12274,N_12332);
or U12518 (N_12518,N_12271,N_12377);
nand U12519 (N_12519,N_12270,N_12227);
nor U12520 (N_12520,N_12390,N_12301);
or U12521 (N_12521,N_12223,N_12311);
and U12522 (N_12522,N_12328,N_12343);
xnor U12523 (N_12523,N_12399,N_12380);
and U12524 (N_12524,N_12377,N_12351);
or U12525 (N_12525,N_12233,N_12336);
xnor U12526 (N_12526,N_12249,N_12229);
and U12527 (N_12527,N_12317,N_12293);
nor U12528 (N_12528,N_12240,N_12312);
and U12529 (N_12529,N_12233,N_12231);
nand U12530 (N_12530,N_12379,N_12216);
nand U12531 (N_12531,N_12267,N_12322);
xnor U12532 (N_12532,N_12295,N_12234);
nor U12533 (N_12533,N_12379,N_12279);
and U12534 (N_12534,N_12364,N_12224);
nand U12535 (N_12535,N_12363,N_12370);
nor U12536 (N_12536,N_12379,N_12364);
nand U12537 (N_12537,N_12201,N_12216);
xor U12538 (N_12538,N_12274,N_12289);
nor U12539 (N_12539,N_12359,N_12395);
nand U12540 (N_12540,N_12329,N_12336);
or U12541 (N_12541,N_12326,N_12365);
xnor U12542 (N_12542,N_12345,N_12214);
xnor U12543 (N_12543,N_12229,N_12295);
and U12544 (N_12544,N_12283,N_12315);
nand U12545 (N_12545,N_12318,N_12227);
and U12546 (N_12546,N_12309,N_12278);
or U12547 (N_12547,N_12289,N_12203);
nand U12548 (N_12548,N_12297,N_12224);
nor U12549 (N_12549,N_12325,N_12337);
or U12550 (N_12550,N_12235,N_12269);
xor U12551 (N_12551,N_12320,N_12288);
nand U12552 (N_12552,N_12243,N_12235);
and U12553 (N_12553,N_12369,N_12204);
and U12554 (N_12554,N_12359,N_12233);
and U12555 (N_12555,N_12227,N_12246);
and U12556 (N_12556,N_12232,N_12361);
and U12557 (N_12557,N_12252,N_12361);
nand U12558 (N_12558,N_12215,N_12302);
or U12559 (N_12559,N_12295,N_12286);
nand U12560 (N_12560,N_12296,N_12385);
and U12561 (N_12561,N_12285,N_12298);
nor U12562 (N_12562,N_12349,N_12357);
nor U12563 (N_12563,N_12333,N_12206);
or U12564 (N_12564,N_12301,N_12374);
nor U12565 (N_12565,N_12309,N_12368);
and U12566 (N_12566,N_12201,N_12204);
xnor U12567 (N_12567,N_12225,N_12335);
nand U12568 (N_12568,N_12312,N_12389);
nand U12569 (N_12569,N_12330,N_12264);
nor U12570 (N_12570,N_12228,N_12313);
nor U12571 (N_12571,N_12379,N_12307);
and U12572 (N_12572,N_12362,N_12380);
nand U12573 (N_12573,N_12262,N_12338);
or U12574 (N_12574,N_12394,N_12309);
nand U12575 (N_12575,N_12203,N_12327);
xnor U12576 (N_12576,N_12326,N_12384);
nor U12577 (N_12577,N_12205,N_12283);
and U12578 (N_12578,N_12308,N_12269);
nand U12579 (N_12579,N_12315,N_12266);
or U12580 (N_12580,N_12237,N_12286);
and U12581 (N_12581,N_12308,N_12362);
nor U12582 (N_12582,N_12343,N_12391);
nor U12583 (N_12583,N_12382,N_12277);
or U12584 (N_12584,N_12268,N_12234);
or U12585 (N_12585,N_12325,N_12306);
xor U12586 (N_12586,N_12358,N_12215);
xor U12587 (N_12587,N_12276,N_12321);
or U12588 (N_12588,N_12261,N_12288);
or U12589 (N_12589,N_12320,N_12342);
and U12590 (N_12590,N_12302,N_12228);
and U12591 (N_12591,N_12303,N_12261);
nand U12592 (N_12592,N_12313,N_12387);
nand U12593 (N_12593,N_12257,N_12261);
nor U12594 (N_12594,N_12346,N_12257);
xor U12595 (N_12595,N_12396,N_12316);
nand U12596 (N_12596,N_12329,N_12292);
and U12597 (N_12597,N_12302,N_12331);
nand U12598 (N_12598,N_12344,N_12346);
and U12599 (N_12599,N_12237,N_12260);
nand U12600 (N_12600,N_12411,N_12509);
nand U12601 (N_12601,N_12578,N_12461);
xor U12602 (N_12602,N_12455,N_12424);
or U12603 (N_12603,N_12561,N_12527);
xnor U12604 (N_12604,N_12420,N_12504);
or U12605 (N_12605,N_12524,N_12535);
nor U12606 (N_12606,N_12454,N_12562);
or U12607 (N_12607,N_12494,N_12404);
nand U12608 (N_12608,N_12441,N_12466);
and U12609 (N_12609,N_12556,N_12512);
or U12610 (N_12610,N_12481,N_12479);
xor U12611 (N_12611,N_12532,N_12475);
and U12612 (N_12612,N_12521,N_12470);
nor U12613 (N_12613,N_12518,N_12443);
nand U12614 (N_12614,N_12526,N_12588);
xor U12615 (N_12615,N_12472,N_12408);
nand U12616 (N_12616,N_12585,N_12410);
nand U12617 (N_12617,N_12540,N_12457);
nor U12618 (N_12618,N_12570,N_12467);
xnor U12619 (N_12619,N_12477,N_12566);
nand U12620 (N_12620,N_12440,N_12548);
nor U12621 (N_12621,N_12418,N_12568);
nor U12622 (N_12622,N_12513,N_12510);
nor U12623 (N_12623,N_12516,N_12537);
and U12624 (N_12624,N_12499,N_12407);
nor U12625 (N_12625,N_12565,N_12575);
xnor U12626 (N_12626,N_12544,N_12473);
and U12627 (N_12627,N_12431,N_12413);
xor U12628 (N_12628,N_12584,N_12591);
nor U12629 (N_12629,N_12459,N_12458);
or U12630 (N_12630,N_12547,N_12492);
nor U12631 (N_12631,N_12495,N_12563);
nand U12632 (N_12632,N_12442,N_12416);
nor U12633 (N_12633,N_12496,N_12511);
nor U12634 (N_12634,N_12403,N_12469);
xnor U12635 (N_12635,N_12488,N_12425);
or U12636 (N_12636,N_12464,N_12572);
xnor U12637 (N_12637,N_12531,N_12595);
nand U12638 (N_12638,N_12439,N_12414);
xnor U12639 (N_12639,N_12599,N_12446);
or U12640 (N_12640,N_12430,N_12541);
nor U12641 (N_12641,N_12447,N_12533);
xor U12642 (N_12642,N_12596,N_12589);
xor U12643 (N_12643,N_12522,N_12560);
nand U12644 (N_12644,N_12412,N_12536);
nor U12645 (N_12645,N_12497,N_12471);
or U12646 (N_12646,N_12480,N_12582);
or U12647 (N_12647,N_12580,N_12483);
xnor U12648 (N_12648,N_12487,N_12543);
nand U12649 (N_12649,N_12465,N_12505);
and U12650 (N_12650,N_12590,N_12448);
nand U12651 (N_12651,N_12426,N_12415);
nor U12652 (N_12652,N_12550,N_12493);
or U12653 (N_12653,N_12546,N_12555);
nand U12654 (N_12654,N_12569,N_12592);
nand U12655 (N_12655,N_12525,N_12553);
nor U12656 (N_12656,N_12490,N_12476);
nand U12657 (N_12657,N_12500,N_12437);
and U12658 (N_12658,N_12463,N_12539);
and U12659 (N_12659,N_12549,N_12597);
nor U12660 (N_12660,N_12583,N_12552);
nand U12661 (N_12661,N_12406,N_12434);
xor U12662 (N_12662,N_12567,N_12489);
and U12663 (N_12663,N_12402,N_12460);
xor U12664 (N_12664,N_12484,N_12528);
nand U12665 (N_12665,N_12514,N_12571);
nor U12666 (N_12666,N_12506,N_12538);
xnor U12667 (N_12667,N_12558,N_12557);
or U12668 (N_12668,N_12577,N_12587);
or U12669 (N_12669,N_12502,N_12445);
and U12670 (N_12670,N_12574,N_12468);
nand U12671 (N_12671,N_12529,N_12433);
nor U12672 (N_12672,N_12405,N_12559);
nand U12673 (N_12673,N_12486,N_12427);
or U12674 (N_12674,N_12444,N_12429);
nor U12675 (N_12675,N_12594,N_12573);
or U12676 (N_12676,N_12520,N_12564);
or U12677 (N_12677,N_12491,N_12432);
or U12678 (N_12678,N_12422,N_12436);
nor U12679 (N_12679,N_12474,N_12507);
or U12680 (N_12680,N_12598,N_12417);
or U12681 (N_12681,N_12428,N_12435);
or U12682 (N_12682,N_12508,N_12438);
nor U12683 (N_12683,N_12554,N_12530);
nor U12684 (N_12684,N_12453,N_12503);
or U12685 (N_12685,N_12519,N_12581);
nand U12686 (N_12686,N_12485,N_12593);
and U12687 (N_12687,N_12456,N_12409);
or U12688 (N_12688,N_12586,N_12579);
or U12689 (N_12689,N_12449,N_12423);
or U12690 (N_12690,N_12400,N_12545);
xor U12691 (N_12691,N_12515,N_12498);
nor U12692 (N_12692,N_12478,N_12401);
or U12693 (N_12693,N_12451,N_12462);
and U12694 (N_12694,N_12419,N_12542);
or U12695 (N_12695,N_12421,N_12551);
xnor U12696 (N_12696,N_12523,N_12452);
nor U12697 (N_12697,N_12450,N_12576);
or U12698 (N_12698,N_12517,N_12534);
nor U12699 (N_12699,N_12482,N_12501);
or U12700 (N_12700,N_12415,N_12521);
or U12701 (N_12701,N_12547,N_12456);
nand U12702 (N_12702,N_12453,N_12573);
nor U12703 (N_12703,N_12463,N_12530);
and U12704 (N_12704,N_12498,N_12474);
nor U12705 (N_12705,N_12598,N_12461);
nand U12706 (N_12706,N_12556,N_12498);
or U12707 (N_12707,N_12494,N_12492);
and U12708 (N_12708,N_12444,N_12506);
nand U12709 (N_12709,N_12471,N_12504);
xor U12710 (N_12710,N_12493,N_12522);
nand U12711 (N_12711,N_12594,N_12423);
xnor U12712 (N_12712,N_12508,N_12412);
xor U12713 (N_12713,N_12427,N_12571);
nand U12714 (N_12714,N_12582,N_12558);
nand U12715 (N_12715,N_12461,N_12437);
nand U12716 (N_12716,N_12577,N_12586);
xor U12717 (N_12717,N_12481,N_12528);
xor U12718 (N_12718,N_12540,N_12589);
nor U12719 (N_12719,N_12482,N_12440);
and U12720 (N_12720,N_12587,N_12584);
nand U12721 (N_12721,N_12589,N_12541);
and U12722 (N_12722,N_12511,N_12469);
xor U12723 (N_12723,N_12558,N_12559);
and U12724 (N_12724,N_12481,N_12502);
and U12725 (N_12725,N_12427,N_12424);
or U12726 (N_12726,N_12416,N_12593);
and U12727 (N_12727,N_12570,N_12583);
and U12728 (N_12728,N_12566,N_12598);
and U12729 (N_12729,N_12437,N_12433);
and U12730 (N_12730,N_12402,N_12514);
or U12731 (N_12731,N_12542,N_12416);
or U12732 (N_12732,N_12429,N_12488);
xnor U12733 (N_12733,N_12478,N_12529);
or U12734 (N_12734,N_12569,N_12461);
or U12735 (N_12735,N_12425,N_12568);
xnor U12736 (N_12736,N_12446,N_12475);
xor U12737 (N_12737,N_12414,N_12517);
xnor U12738 (N_12738,N_12494,N_12451);
xor U12739 (N_12739,N_12404,N_12484);
or U12740 (N_12740,N_12429,N_12453);
nand U12741 (N_12741,N_12472,N_12556);
or U12742 (N_12742,N_12485,N_12547);
nand U12743 (N_12743,N_12450,N_12440);
xor U12744 (N_12744,N_12450,N_12585);
xnor U12745 (N_12745,N_12457,N_12482);
and U12746 (N_12746,N_12477,N_12498);
or U12747 (N_12747,N_12520,N_12471);
nand U12748 (N_12748,N_12595,N_12408);
or U12749 (N_12749,N_12412,N_12598);
nand U12750 (N_12750,N_12468,N_12428);
nor U12751 (N_12751,N_12423,N_12516);
nand U12752 (N_12752,N_12482,N_12568);
or U12753 (N_12753,N_12436,N_12421);
nor U12754 (N_12754,N_12499,N_12561);
xnor U12755 (N_12755,N_12532,N_12513);
nor U12756 (N_12756,N_12545,N_12559);
nor U12757 (N_12757,N_12514,N_12475);
and U12758 (N_12758,N_12485,N_12521);
and U12759 (N_12759,N_12474,N_12592);
nor U12760 (N_12760,N_12547,N_12520);
xnor U12761 (N_12761,N_12529,N_12560);
nand U12762 (N_12762,N_12470,N_12440);
nor U12763 (N_12763,N_12514,N_12517);
or U12764 (N_12764,N_12593,N_12480);
nor U12765 (N_12765,N_12479,N_12552);
xor U12766 (N_12766,N_12556,N_12586);
and U12767 (N_12767,N_12476,N_12544);
xor U12768 (N_12768,N_12522,N_12458);
and U12769 (N_12769,N_12558,N_12419);
xor U12770 (N_12770,N_12446,N_12526);
and U12771 (N_12771,N_12525,N_12524);
and U12772 (N_12772,N_12443,N_12550);
nand U12773 (N_12773,N_12529,N_12462);
and U12774 (N_12774,N_12442,N_12535);
xnor U12775 (N_12775,N_12415,N_12514);
or U12776 (N_12776,N_12468,N_12501);
nor U12777 (N_12777,N_12552,N_12427);
nand U12778 (N_12778,N_12412,N_12466);
nand U12779 (N_12779,N_12488,N_12435);
nand U12780 (N_12780,N_12467,N_12583);
nand U12781 (N_12781,N_12516,N_12585);
or U12782 (N_12782,N_12520,N_12422);
and U12783 (N_12783,N_12449,N_12537);
or U12784 (N_12784,N_12516,N_12476);
and U12785 (N_12785,N_12571,N_12466);
xnor U12786 (N_12786,N_12462,N_12471);
nand U12787 (N_12787,N_12502,N_12444);
and U12788 (N_12788,N_12472,N_12456);
or U12789 (N_12789,N_12473,N_12445);
xor U12790 (N_12790,N_12448,N_12406);
nor U12791 (N_12791,N_12420,N_12523);
or U12792 (N_12792,N_12590,N_12581);
or U12793 (N_12793,N_12506,N_12508);
nand U12794 (N_12794,N_12591,N_12423);
and U12795 (N_12795,N_12565,N_12555);
xor U12796 (N_12796,N_12455,N_12567);
or U12797 (N_12797,N_12509,N_12582);
nand U12798 (N_12798,N_12433,N_12591);
nor U12799 (N_12799,N_12462,N_12416);
nand U12800 (N_12800,N_12759,N_12656);
nor U12801 (N_12801,N_12643,N_12629);
or U12802 (N_12802,N_12620,N_12625);
and U12803 (N_12803,N_12623,N_12631);
nor U12804 (N_12804,N_12709,N_12779);
nor U12805 (N_12805,N_12677,N_12712);
nand U12806 (N_12806,N_12770,N_12644);
nor U12807 (N_12807,N_12756,N_12765);
or U12808 (N_12808,N_12793,N_12668);
xnor U12809 (N_12809,N_12601,N_12727);
nand U12810 (N_12810,N_12664,N_12760);
nand U12811 (N_12811,N_12790,N_12688);
nor U12812 (N_12812,N_12730,N_12784);
nand U12813 (N_12813,N_12660,N_12799);
or U12814 (N_12814,N_12610,N_12692);
or U12815 (N_12815,N_12788,N_12714);
nor U12816 (N_12816,N_12605,N_12674);
xnor U12817 (N_12817,N_12641,N_12676);
nand U12818 (N_12818,N_12675,N_12780);
nor U12819 (N_12819,N_12711,N_12723);
or U12820 (N_12820,N_12689,N_12744);
or U12821 (N_12821,N_12651,N_12606);
xnor U12822 (N_12822,N_12632,N_12761);
xnor U12823 (N_12823,N_12786,N_12671);
and U12824 (N_12824,N_12769,N_12719);
or U12825 (N_12825,N_12763,N_12791);
nor U12826 (N_12826,N_12745,N_12696);
or U12827 (N_12827,N_12737,N_12762);
and U12828 (N_12828,N_12713,N_12720);
nor U12829 (N_12829,N_12774,N_12750);
nand U12830 (N_12830,N_12646,N_12691);
nor U12831 (N_12831,N_12652,N_12742);
nor U12832 (N_12832,N_12650,N_12670);
xor U12833 (N_12833,N_12721,N_12628);
or U12834 (N_12834,N_12642,N_12658);
and U12835 (N_12835,N_12722,N_12697);
and U12836 (N_12836,N_12752,N_12653);
or U12837 (N_12837,N_12639,N_12715);
nor U12838 (N_12838,N_12754,N_12731);
nand U12839 (N_12839,N_12699,N_12751);
nand U12840 (N_12840,N_12796,N_12798);
nor U12841 (N_12841,N_12782,N_12704);
xnor U12842 (N_12842,N_12789,N_12797);
nor U12843 (N_12843,N_12661,N_12776);
xnor U12844 (N_12844,N_12706,N_12647);
nor U12845 (N_12845,N_12729,N_12705);
nor U12846 (N_12846,N_12621,N_12702);
nor U12847 (N_12847,N_12627,N_12667);
nor U12848 (N_12848,N_12794,N_12739);
nand U12849 (N_12849,N_12710,N_12766);
nand U12850 (N_12850,N_12600,N_12672);
and U12851 (N_12851,N_12666,N_12686);
or U12852 (N_12852,N_12637,N_12662);
xor U12853 (N_12853,N_12783,N_12778);
xnor U12854 (N_12854,N_12734,N_12613);
nor U12855 (N_12855,N_12685,N_12680);
and U12856 (N_12856,N_12619,N_12787);
and U12857 (N_12857,N_12693,N_12669);
nor U12858 (N_12858,N_12648,N_12771);
nor U12859 (N_12859,N_12792,N_12645);
and U12860 (N_12860,N_12682,N_12728);
and U12861 (N_12861,N_12681,N_12636);
nor U12862 (N_12862,N_12700,N_12725);
nor U12863 (N_12863,N_12733,N_12736);
and U12864 (N_12864,N_12795,N_12755);
nand U12865 (N_12865,N_12701,N_12768);
or U12866 (N_12866,N_12757,N_12602);
nor U12867 (N_12867,N_12740,N_12694);
xnor U12868 (N_12868,N_12718,N_12659);
nand U12869 (N_12869,N_12683,N_12614);
xor U12870 (N_12870,N_12684,N_12748);
or U12871 (N_12871,N_12758,N_12615);
and U12872 (N_12872,N_12777,N_12603);
xnor U12873 (N_12873,N_12735,N_12633);
xnor U12874 (N_12874,N_12630,N_12611);
and U12875 (N_12875,N_12673,N_12663);
and U12876 (N_12876,N_12608,N_12624);
nand U12877 (N_12877,N_12687,N_12716);
nand U12878 (N_12878,N_12781,N_12635);
and U12879 (N_12879,N_12665,N_12678);
and U12880 (N_12880,N_12738,N_12764);
xnor U12881 (N_12881,N_12612,N_12657);
and U12882 (N_12882,N_12707,N_12640);
xor U12883 (N_12883,N_12717,N_12604);
nand U12884 (N_12884,N_12626,N_12732);
and U12885 (N_12885,N_12654,N_12617);
xnor U12886 (N_12886,N_12679,N_12618);
nor U12887 (N_12887,N_12607,N_12622);
and U12888 (N_12888,N_12698,N_12616);
nor U12889 (N_12889,N_12749,N_12726);
xnor U12890 (N_12890,N_12773,N_12767);
xnor U12891 (N_12891,N_12634,N_12746);
nand U12892 (N_12892,N_12703,N_12785);
nand U12893 (N_12893,N_12609,N_12741);
xnor U12894 (N_12894,N_12695,N_12775);
nand U12895 (N_12895,N_12753,N_12747);
and U12896 (N_12896,N_12690,N_12649);
xor U12897 (N_12897,N_12724,N_12772);
nor U12898 (N_12898,N_12708,N_12638);
nand U12899 (N_12899,N_12655,N_12743);
or U12900 (N_12900,N_12637,N_12712);
nand U12901 (N_12901,N_12650,N_12713);
nand U12902 (N_12902,N_12785,N_12603);
xnor U12903 (N_12903,N_12770,N_12727);
nand U12904 (N_12904,N_12703,N_12654);
or U12905 (N_12905,N_12728,N_12774);
nand U12906 (N_12906,N_12730,N_12679);
nor U12907 (N_12907,N_12698,N_12615);
nand U12908 (N_12908,N_12748,N_12645);
nor U12909 (N_12909,N_12622,N_12654);
xor U12910 (N_12910,N_12705,N_12604);
xnor U12911 (N_12911,N_12674,N_12607);
or U12912 (N_12912,N_12672,N_12733);
nor U12913 (N_12913,N_12705,N_12654);
xnor U12914 (N_12914,N_12619,N_12790);
or U12915 (N_12915,N_12631,N_12789);
or U12916 (N_12916,N_12787,N_12644);
or U12917 (N_12917,N_12704,N_12662);
nor U12918 (N_12918,N_12799,N_12756);
nor U12919 (N_12919,N_12750,N_12722);
and U12920 (N_12920,N_12753,N_12752);
or U12921 (N_12921,N_12753,N_12708);
nor U12922 (N_12922,N_12750,N_12690);
xor U12923 (N_12923,N_12611,N_12691);
or U12924 (N_12924,N_12678,N_12605);
nor U12925 (N_12925,N_12775,N_12705);
and U12926 (N_12926,N_12740,N_12664);
and U12927 (N_12927,N_12778,N_12744);
or U12928 (N_12928,N_12726,N_12795);
xor U12929 (N_12929,N_12648,N_12620);
nor U12930 (N_12930,N_12605,N_12718);
nor U12931 (N_12931,N_12609,N_12712);
nor U12932 (N_12932,N_12767,N_12692);
and U12933 (N_12933,N_12642,N_12704);
or U12934 (N_12934,N_12691,N_12795);
nand U12935 (N_12935,N_12775,N_12625);
xnor U12936 (N_12936,N_12655,N_12682);
nand U12937 (N_12937,N_12770,N_12613);
or U12938 (N_12938,N_12657,N_12729);
or U12939 (N_12939,N_12667,N_12739);
and U12940 (N_12940,N_12641,N_12669);
nand U12941 (N_12941,N_12646,N_12780);
xor U12942 (N_12942,N_12715,N_12745);
nor U12943 (N_12943,N_12630,N_12696);
or U12944 (N_12944,N_12722,N_12776);
or U12945 (N_12945,N_12643,N_12616);
and U12946 (N_12946,N_12613,N_12716);
nand U12947 (N_12947,N_12738,N_12664);
or U12948 (N_12948,N_12742,N_12663);
nor U12949 (N_12949,N_12789,N_12610);
nor U12950 (N_12950,N_12658,N_12666);
xnor U12951 (N_12951,N_12729,N_12630);
xnor U12952 (N_12952,N_12686,N_12721);
and U12953 (N_12953,N_12604,N_12745);
or U12954 (N_12954,N_12765,N_12741);
xnor U12955 (N_12955,N_12601,N_12770);
or U12956 (N_12956,N_12733,N_12739);
or U12957 (N_12957,N_12694,N_12629);
xor U12958 (N_12958,N_12636,N_12721);
nand U12959 (N_12959,N_12697,N_12749);
xnor U12960 (N_12960,N_12696,N_12739);
and U12961 (N_12961,N_12707,N_12627);
nand U12962 (N_12962,N_12784,N_12721);
nor U12963 (N_12963,N_12724,N_12745);
nand U12964 (N_12964,N_12630,N_12752);
nand U12965 (N_12965,N_12684,N_12612);
nor U12966 (N_12966,N_12769,N_12717);
nor U12967 (N_12967,N_12648,N_12758);
or U12968 (N_12968,N_12725,N_12761);
and U12969 (N_12969,N_12794,N_12720);
or U12970 (N_12970,N_12602,N_12689);
nand U12971 (N_12971,N_12784,N_12742);
nor U12972 (N_12972,N_12750,N_12604);
nor U12973 (N_12973,N_12670,N_12764);
nor U12974 (N_12974,N_12796,N_12688);
nor U12975 (N_12975,N_12741,N_12753);
xor U12976 (N_12976,N_12716,N_12727);
or U12977 (N_12977,N_12644,N_12778);
nand U12978 (N_12978,N_12727,N_12717);
and U12979 (N_12979,N_12787,N_12654);
nor U12980 (N_12980,N_12734,N_12695);
nor U12981 (N_12981,N_12685,N_12682);
xor U12982 (N_12982,N_12636,N_12690);
xnor U12983 (N_12983,N_12612,N_12689);
nor U12984 (N_12984,N_12786,N_12620);
nand U12985 (N_12985,N_12711,N_12693);
nand U12986 (N_12986,N_12682,N_12665);
and U12987 (N_12987,N_12731,N_12635);
or U12988 (N_12988,N_12725,N_12646);
or U12989 (N_12989,N_12722,N_12771);
nand U12990 (N_12990,N_12650,N_12666);
xor U12991 (N_12991,N_12788,N_12710);
and U12992 (N_12992,N_12638,N_12785);
and U12993 (N_12993,N_12759,N_12760);
and U12994 (N_12994,N_12791,N_12765);
xnor U12995 (N_12995,N_12704,N_12627);
xor U12996 (N_12996,N_12738,N_12676);
nor U12997 (N_12997,N_12705,N_12785);
xor U12998 (N_12998,N_12646,N_12756);
nand U12999 (N_12999,N_12751,N_12723);
or U13000 (N_13000,N_12832,N_12879);
nand U13001 (N_13001,N_12961,N_12871);
nor U13002 (N_13002,N_12849,N_12842);
nor U13003 (N_13003,N_12900,N_12895);
or U13004 (N_13004,N_12894,N_12998);
nand U13005 (N_13005,N_12927,N_12860);
or U13006 (N_13006,N_12887,N_12815);
nor U13007 (N_13007,N_12876,N_12833);
nand U13008 (N_13008,N_12996,N_12977);
nand U13009 (N_13009,N_12918,N_12899);
nor U13010 (N_13010,N_12829,N_12821);
and U13011 (N_13011,N_12892,N_12969);
xor U13012 (N_13012,N_12956,N_12932);
or U13013 (N_13013,N_12960,N_12855);
nor U13014 (N_13014,N_12859,N_12917);
nor U13015 (N_13015,N_12968,N_12913);
or U13016 (N_13016,N_12869,N_12803);
or U13017 (N_13017,N_12920,N_12931);
or U13018 (N_13018,N_12810,N_12962);
and U13019 (N_13019,N_12885,N_12883);
and U13020 (N_13020,N_12906,N_12959);
nor U13021 (N_13021,N_12828,N_12915);
or U13022 (N_13022,N_12835,N_12807);
xor U13023 (N_13023,N_12991,N_12862);
nor U13024 (N_13024,N_12904,N_12800);
nor U13025 (N_13025,N_12980,N_12973);
nor U13026 (N_13026,N_12929,N_12878);
or U13027 (N_13027,N_12943,N_12908);
and U13028 (N_13028,N_12861,N_12978);
or U13029 (N_13029,N_12901,N_12847);
nand U13030 (N_13030,N_12804,N_12999);
nor U13031 (N_13031,N_12986,N_12825);
xnor U13032 (N_13032,N_12930,N_12814);
or U13033 (N_13033,N_12924,N_12845);
nand U13034 (N_13034,N_12976,N_12928);
xnor U13035 (N_13035,N_12897,N_12873);
nor U13036 (N_13036,N_12801,N_12942);
nor U13037 (N_13037,N_12818,N_12851);
xnor U13038 (N_13038,N_12870,N_12830);
or U13039 (N_13039,N_12819,N_12853);
xor U13040 (N_13040,N_12993,N_12837);
and U13041 (N_13041,N_12914,N_12974);
xor U13042 (N_13042,N_12933,N_12891);
nor U13043 (N_13043,N_12858,N_12946);
nand U13044 (N_13044,N_12990,N_12912);
and U13045 (N_13045,N_12981,N_12963);
nor U13046 (N_13046,N_12872,N_12827);
or U13047 (N_13047,N_12941,N_12983);
nor U13048 (N_13048,N_12957,N_12936);
nand U13049 (N_13049,N_12857,N_12984);
nand U13050 (N_13050,N_12854,N_12903);
or U13051 (N_13051,N_12948,N_12867);
or U13052 (N_13052,N_12822,N_12839);
xor U13053 (N_13053,N_12886,N_12806);
nor U13054 (N_13054,N_12898,N_12964);
or U13055 (N_13055,N_12923,N_12919);
or U13056 (N_13056,N_12884,N_12826);
and U13057 (N_13057,N_12850,N_12965);
or U13058 (N_13058,N_12840,N_12893);
xor U13059 (N_13059,N_12848,N_12813);
xor U13060 (N_13060,N_12890,N_12947);
xor U13061 (N_13061,N_12951,N_12809);
nor U13062 (N_13062,N_12910,N_12967);
nand U13063 (N_13063,N_12875,N_12966);
or U13064 (N_13064,N_12882,N_12868);
nor U13065 (N_13065,N_12805,N_12856);
nand U13066 (N_13066,N_12972,N_12877);
nand U13067 (N_13067,N_12922,N_12911);
or U13068 (N_13068,N_12926,N_12866);
nor U13069 (N_13069,N_12985,N_12896);
nor U13070 (N_13070,N_12907,N_12952);
xor U13071 (N_13071,N_12823,N_12958);
nor U13072 (N_13072,N_12874,N_12989);
nor U13073 (N_13073,N_12987,N_12979);
nor U13074 (N_13074,N_12953,N_12816);
nand U13075 (N_13075,N_12955,N_12844);
xnor U13076 (N_13076,N_12880,N_12905);
xor U13077 (N_13077,N_12925,N_12949);
and U13078 (N_13078,N_12846,N_12888);
nor U13079 (N_13079,N_12889,N_12802);
nand U13080 (N_13080,N_12834,N_12881);
nand U13081 (N_13081,N_12935,N_12864);
nor U13082 (N_13082,N_12863,N_12944);
nand U13083 (N_13083,N_12820,N_12940);
xnor U13084 (N_13084,N_12950,N_12817);
nand U13085 (N_13085,N_12938,N_12988);
nor U13086 (N_13086,N_12902,N_12945);
xor U13087 (N_13087,N_12970,N_12831);
and U13088 (N_13088,N_12934,N_12909);
and U13089 (N_13089,N_12971,N_12997);
nand U13090 (N_13090,N_12954,N_12808);
nor U13091 (N_13091,N_12995,N_12937);
or U13092 (N_13092,N_12994,N_12975);
or U13093 (N_13093,N_12812,N_12939);
or U13094 (N_13094,N_12841,N_12916);
nand U13095 (N_13095,N_12865,N_12921);
nor U13096 (N_13096,N_12992,N_12811);
nand U13097 (N_13097,N_12852,N_12824);
or U13098 (N_13098,N_12982,N_12838);
or U13099 (N_13099,N_12836,N_12843);
nand U13100 (N_13100,N_12900,N_12961);
nand U13101 (N_13101,N_12997,N_12878);
nor U13102 (N_13102,N_12838,N_12984);
and U13103 (N_13103,N_12874,N_12923);
nor U13104 (N_13104,N_12834,N_12953);
nand U13105 (N_13105,N_12884,N_12976);
xnor U13106 (N_13106,N_12964,N_12930);
nand U13107 (N_13107,N_12872,N_12928);
nor U13108 (N_13108,N_12861,N_12940);
nand U13109 (N_13109,N_12889,N_12922);
nand U13110 (N_13110,N_12956,N_12900);
or U13111 (N_13111,N_12806,N_12871);
nand U13112 (N_13112,N_12973,N_12872);
and U13113 (N_13113,N_12929,N_12937);
nand U13114 (N_13114,N_12971,N_12998);
and U13115 (N_13115,N_12943,N_12946);
nand U13116 (N_13116,N_12890,N_12925);
and U13117 (N_13117,N_12861,N_12922);
nor U13118 (N_13118,N_12826,N_12861);
or U13119 (N_13119,N_12906,N_12886);
or U13120 (N_13120,N_12815,N_12866);
xnor U13121 (N_13121,N_12973,N_12956);
or U13122 (N_13122,N_12802,N_12821);
or U13123 (N_13123,N_12855,N_12801);
or U13124 (N_13124,N_12947,N_12928);
nor U13125 (N_13125,N_12978,N_12945);
nor U13126 (N_13126,N_12814,N_12823);
nand U13127 (N_13127,N_12853,N_12837);
xor U13128 (N_13128,N_12910,N_12801);
and U13129 (N_13129,N_12946,N_12806);
or U13130 (N_13130,N_12962,N_12954);
or U13131 (N_13131,N_12978,N_12822);
and U13132 (N_13132,N_12939,N_12898);
xnor U13133 (N_13133,N_12893,N_12890);
or U13134 (N_13134,N_12953,N_12913);
and U13135 (N_13135,N_12985,N_12821);
nand U13136 (N_13136,N_12876,N_12927);
and U13137 (N_13137,N_12873,N_12933);
nor U13138 (N_13138,N_12832,N_12818);
and U13139 (N_13139,N_12816,N_12893);
or U13140 (N_13140,N_12822,N_12819);
and U13141 (N_13141,N_12864,N_12829);
and U13142 (N_13142,N_12845,N_12964);
and U13143 (N_13143,N_12987,N_12830);
nand U13144 (N_13144,N_12860,N_12828);
or U13145 (N_13145,N_12956,N_12967);
and U13146 (N_13146,N_12898,N_12847);
and U13147 (N_13147,N_12829,N_12919);
nor U13148 (N_13148,N_12877,N_12983);
nand U13149 (N_13149,N_12881,N_12961);
and U13150 (N_13150,N_12820,N_12978);
xnor U13151 (N_13151,N_12916,N_12860);
nor U13152 (N_13152,N_12913,N_12982);
and U13153 (N_13153,N_12962,N_12948);
or U13154 (N_13154,N_12879,N_12942);
and U13155 (N_13155,N_12874,N_12848);
xnor U13156 (N_13156,N_12819,N_12831);
nor U13157 (N_13157,N_12886,N_12960);
xor U13158 (N_13158,N_12935,N_12973);
or U13159 (N_13159,N_12920,N_12836);
xnor U13160 (N_13160,N_12884,N_12932);
nand U13161 (N_13161,N_12945,N_12920);
xor U13162 (N_13162,N_12994,N_12887);
and U13163 (N_13163,N_12803,N_12838);
or U13164 (N_13164,N_12979,N_12959);
nand U13165 (N_13165,N_12827,N_12922);
or U13166 (N_13166,N_12870,N_12965);
xnor U13167 (N_13167,N_12841,N_12853);
and U13168 (N_13168,N_12876,N_12811);
and U13169 (N_13169,N_12959,N_12965);
nor U13170 (N_13170,N_12851,N_12847);
nor U13171 (N_13171,N_12852,N_12940);
or U13172 (N_13172,N_12919,N_12979);
and U13173 (N_13173,N_12941,N_12907);
nor U13174 (N_13174,N_12842,N_12946);
or U13175 (N_13175,N_12944,N_12974);
nor U13176 (N_13176,N_12880,N_12953);
xnor U13177 (N_13177,N_12994,N_12939);
xnor U13178 (N_13178,N_12925,N_12980);
nand U13179 (N_13179,N_12824,N_12948);
or U13180 (N_13180,N_12928,N_12933);
and U13181 (N_13181,N_12910,N_12855);
or U13182 (N_13182,N_12848,N_12919);
nor U13183 (N_13183,N_12915,N_12929);
xnor U13184 (N_13184,N_12949,N_12920);
and U13185 (N_13185,N_12944,N_12913);
and U13186 (N_13186,N_12956,N_12879);
nand U13187 (N_13187,N_12866,N_12876);
nand U13188 (N_13188,N_12931,N_12894);
nor U13189 (N_13189,N_12905,N_12859);
nand U13190 (N_13190,N_12871,N_12891);
nand U13191 (N_13191,N_12827,N_12807);
nor U13192 (N_13192,N_12859,N_12989);
and U13193 (N_13193,N_12890,N_12884);
nand U13194 (N_13194,N_12838,N_12998);
and U13195 (N_13195,N_12861,N_12952);
or U13196 (N_13196,N_12921,N_12993);
or U13197 (N_13197,N_12802,N_12936);
nand U13198 (N_13198,N_12986,N_12861);
or U13199 (N_13199,N_12987,N_12996);
nor U13200 (N_13200,N_13012,N_13181);
nor U13201 (N_13201,N_13150,N_13189);
or U13202 (N_13202,N_13165,N_13031);
nor U13203 (N_13203,N_13171,N_13042);
nand U13204 (N_13204,N_13036,N_13019);
or U13205 (N_13205,N_13123,N_13086);
xnor U13206 (N_13206,N_13060,N_13184);
or U13207 (N_13207,N_13063,N_13175);
xor U13208 (N_13208,N_13152,N_13136);
nand U13209 (N_13209,N_13172,N_13061);
nor U13210 (N_13210,N_13056,N_13114);
nor U13211 (N_13211,N_13021,N_13053);
nor U13212 (N_13212,N_13049,N_13182);
or U13213 (N_13213,N_13134,N_13174);
nand U13214 (N_13214,N_13074,N_13149);
or U13215 (N_13215,N_13026,N_13162);
or U13216 (N_13216,N_13046,N_13105);
xor U13217 (N_13217,N_13194,N_13138);
nand U13218 (N_13218,N_13109,N_13160);
nor U13219 (N_13219,N_13128,N_13115);
nand U13220 (N_13220,N_13020,N_13108);
nand U13221 (N_13221,N_13062,N_13052);
and U13222 (N_13222,N_13185,N_13028);
nand U13223 (N_13223,N_13085,N_13142);
nor U13224 (N_13224,N_13163,N_13016);
or U13225 (N_13225,N_13018,N_13039);
nor U13226 (N_13226,N_13041,N_13089);
nand U13227 (N_13227,N_13083,N_13111);
nand U13228 (N_13228,N_13169,N_13179);
and U13229 (N_13229,N_13176,N_13195);
xnor U13230 (N_13230,N_13067,N_13094);
nor U13231 (N_13231,N_13084,N_13047);
or U13232 (N_13232,N_13054,N_13102);
xor U13233 (N_13233,N_13193,N_13075);
nor U13234 (N_13234,N_13071,N_13013);
xor U13235 (N_13235,N_13113,N_13091);
or U13236 (N_13236,N_13166,N_13095);
nor U13237 (N_13237,N_13130,N_13096);
xor U13238 (N_13238,N_13186,N_13139);
xnor U13239 (N_13239,N_13058,N_13079);
xnor U13240 (N_13240,N_13196,N_13069);
xor U13241 (N_13241,N_13100,N_13192);
or U13242 (N_13242,N_13043,N_13072);
or U13243 (N_13243,N_13155,N_13168);
nor U13244 (N_13244,N_13001,N_13147);
and U13245 (N_13245,N_13158,N_13064);
and U13246 (N_13246,N_13187,N_13038);
or U13247 (N_13247,N_13077,N_13017);
nand U13248 (N_13248,N_13118,N_13051);
and U13249 (N_13249,N_13104,N_13198);
xor U13250 (N_13250,N_13112,N_13164);
and U13251 (N_13251,N_13010,N_13059);
and U13252 (N_13252,N_13098,N_13143);
nand U13253 (N_13253,N_13180,N_13173);
nor U13254 (N_13254,N_13022,N_13119);
nand U13255 (N_13255,N_13027,N_13090);
and U13256 (N_13256,N_13005,N_13023);
nor U13257 (N_13257,N_13127,N_13199);
xnor U13258 (N_13258,N_13066,N_13146);
nor U13259 (N_13259,N_13070,N_13153);
or U13260 (N_13260,N_13110,N_13093);
xnor U13261 (N_13261,N_13004,N_13092);
nor U13262 (N_13262,N_13024,N_13002);
nor U13263 (N_13263,N_13121,N_13088);
nand U13264 (N_13264,N_13131,N_13057);
nand U13265 (N_13265,N_13190,N_13133);
and U13266 (N_13266,N_13145,N_13122);
xnor U13267 (N_13267,N_13040,N_13030);
or U13268 (N_13268,N_13135,N_13120);
or U13269 (N_13269,N_13144,N_13197);
or U13270 (N_13270,N_13178,N_13101);
nor U13271 (N_13271,N_13034,N_13125);
nand U13272 (N_13272,N_13183,N_13029);
xnor U13273 (N_13273,N_13124,N_13156);
and U13274 (N_13274,N_13032,N_13106);
nor U13275 (N_13275,N_13033,N_13014);
xor U13276 (N_13276,N_13003,N_13161);
xnor U13277 (N_13277,N_13132,N_13117);
or U13278 (N_13278,N_13068,N_13103);
xnor U13279 (N_13279,N_13006,N_13048);
nor U13280 (N_13280,N_13129,N_13116);
xor U13281 (N_13281,N_13087,N_13154);
nor U13282 (N_13282,N_13141,N_13009);
and U13283 (N_13283,N_13082,N_13177);
xor U13284 (N_13284,N_13076,N_13159);
nand U13285 (N_13285,N_13073,N_13137);
or U13286 (N_13286,N_13099,N_13148);
and U13287 (N_13287,N_13188,N_13081);
nand U13288 (N_13288,N_13080,N_13170);
xnor U13289 (N_13289,N_13167,N_13015);
nand U13290 (N_13290,N_13191,N_13157);
or U13291 (N_13291,N_13037,N_13107);
or U13292 (N_13292,N_13097,N_13025);
xnor U13293 (N_13293,N_13126,N_13000);
and U13294 (N_13294,N_13078,N_13050);
xor U13295 (N_13295,N_13151,N_13055);
nand U13296 (N_13296,N_13045,N_13008);
or U13297 (N_13297,N_13044,N_13140);
xor U13298 (N_13298,N_13035,N_13007);
xor U13299 (N_13299,N_13011,N_13065);
xor U13300 (N_13300,N_13088,N_13069);
or U13301 (N_13301,N_13101,N_13007);
or U13302 (N_13302,N_13116,N_13198);
nand U13303 (N_13303,N_13038,N_13178);
nor U13304 (N_13304,N_13005,N_13152);
nor U13305 (N_13305,N_13069,N_13195);
nand U13306 (N_13306,N_13159,N_13173);
and U13307 (N_13307,N_13136,N_13045);
nor U13308 (N_13308,N_13162,N_13176);
nor U13309 (N_13309,N_13159,N_13051);
or U13310 (N_13310,N_13032,N_13158);
nand U13311 (N_13311,N_13084,N_13175);
nor U13312 (N_13312,N_13099,N_13052);
and U13313 (N_13313,N_13032,N_13183);
nand U13314 (N_13314,N_13120,N_13142);
and U13315 (N_13315,N_13121,N_13197);
nor U13316 (N_13316,N_13123,N_13174);
xor U13317 (N_13317,N_13119,N_13175);
xnor U13318 (N_13318,N_13091,N_13045);
or U13319 (N_13319,N_13077,N_13141);
xor U13320 (N_13320,N_13045,N_13117);
and U13321 (N_13321,N_13090,N_13055);
nand U13322 (N_13322,N_13098,N_13090);
or U13323 (N_13323,N_13046,N_13123);
or U13324 (N_13324,N_13018,N_13041);
nor U13325 (N_13325,N_13094,N_13190);
or U13326 (N_13326,N_13050,N_13033);
nand U13327 (N_13327,N_13090,N_13149);
xnor U13328 (N_13328,N_13165,N_13016);
xnor U13329 (N_13329,N_13130,N_13018);
or U13330 (N_13330,N_13045,N_13152);
nor U13331 (N_13331,N_13112,N_13159);
nand U13332 (N_13332,N_13074,N_13053);
nand U13333 (N_13333,N_13181,N_13118);
and U13334 (N_13334,N_13097,N_13118);
or U13335 (N_13335,N_13176,N_13136);
xnor U13336 (N_13336,N_13128,N_13006);
nand U13337 (N_13337,N_13199,N_13196);
nand U13338 (N_13338,N_13170,N_13043);
or U13339 (N_13339,N_13056,N_13078);
or U13340 (N_13340,N_13165,N_13012);
nor U13341 (N_13341,N_13124,N_13180);
nand U13342 (N_13342,N_13106,N_13068);
or U13343 (N_13343,N_13154,N_13127);
or U13344 (N_13344,N_13023,N_13050);
nand U13345 (N_13345,N_13132,N_13024);
or U13346 (N_13346,N_13036,N_13060);
xor U13347 (N_13347,N_13062,N_13028);
and U13348 (N_13348,N_13098,N_13169);
nand U13349 (N_13349,N_13034,N_13095);
nand U13350 (N_13350,N_13021,N_13064);
xnor U13351 (N_13351,N_13042,N_13113);
nor U13352 (N_13352,N_13183,N_13033);
or U13353 (N_13353,N_13139,N_13151);
and U13354 (N_13354,N_13133,N_13012);
or U13355 (N_13355,N_13070,N_13097);
and U13356 (N_13356,N_13054,N_13122);
xor U13357 (N_13357,N_13194,N_13167);
or U13358 (N_13358,N_13071,N_13145);
xnor U13359 (N_13359,N_13134,N_13180);
xnor U13360 (N_13360,N_13051,N_13043);
or U13361 (N_13361,N_13071,N_13109);
and U13362 (N_13362,N_13045,N_13167);
or U13363 (N_13363,N_13100,N_13087);
nand U13364 (N_13364,N_13159,N_13043);
nor U13365 (N_13365,N_13117,N_13134);
nor U13366 (N_13366,N_13184,N_13172);
xnor U13367 (N_13367,N_13018,N_13138);
xor U13368 (N_13368,N_13058,N_13096);
or U13369 (N_13369,N_13185,N_13003);
xor U13370 (N_13370,N_13114,N_13042);
or U13371 (N_13371,N_13139,N_13046);
and U13372 (N_13372,N_13171,N_13007);
nor U13373 (N_13373,N_13150,N_13130);
or U13374 (N_13374,N_13068,N_13132);
xor U13375 (N_13375,N_13032,N_13013);
and U13376 (N_13376,N_13150,N_13014);
and U13377 (N_13377,N_13016,N_13105);
and U13378 (N_13378,N_13178,N_13043);
xnor U13379 (N_13379,N_13005,N_13164);
or U13380 (N_13380,N_13044,N_13156);
nand U13381 (N_13381,N_13124,N_13157);
and U13382 (N_13382,N_13032,N_13079);
xor U13383 (N_13383,N_13067,N_13058);
nor U13384 (N_13384,N_13100,N_13171);
and U13385 (N_13385,N_13037,N_13044);
and U13386 (N_13386,N_13168,N_13083);
xor U13387 (N_13387,N_13058,N_13031);
and U13388 (N_13388,N_13139,N_13039);
xnor U13389 (N_13389,N_13009,N_13024);
or U13390 (N_13390,N_13091,N_13187);
nand U13391 (N_13391,N_13019,N_13052);
xor U13392 (N_13392,N_13012,N_13033);
nand U13393 (N_13393,N_13030,N_13004);
nor U13394 (N_13394,N_13074,N_13060);
xor U13395 (N_13395,N_13086,N_13193);
nor U13396 (N_13396,N_13188,N_13115);
nand U13397 (N_13397,N_13147,N_13071);
nor U13398 (N_13398,N_13192,N_13012);
xor U13399 (N_13399,N_13093,N_13124);
nor U13400 (N_13400,N_13283,N_13361);
or U13401 (N_13401,N_13261,N_13342);
nand U13402 (N_13402,N_13387,N_13217);
nor U13403 (N_13403,N_13391,N_13231);
nor U13404 (N_13404,N_13330,N_13305);
and U13405 (N_13405,N_13357,N_13273);
nand U13406 (N_13406,N_13275,N_13352);
xnor U13407 (N_13407,N_13284,N_13326);
xor U13408 (N_13408,N_13346,N_13208);
or U13409 (N_13409,N_13263,N_13392);
nand U13410 (N_13410,N_13218,N_13382);
nand U13411 (N_13411,N_13223,N_13246);
or U13412 (N_13412,N_13227,N_13201);
and U13413 (N_13413,N_13235,N_13203);
and U13414 (N_13414,N_13258,N_13270);
and U13415 (N_13415,N_13397,N_13359);
nor U13416 (N_13416,N_13210,N_13206);
and U13417 (N_13417,N_13215,N_13287);
nor U13418 (N_13418,N_13225,N_13276);
or U13419 (N_13419,N_13345,N_13328);
nor U13420 (N_13420,N_13380,N_13351);
or U13421 (N_13421,N_13333,N_13377);
or U13422 (N_13422,N_13375,N_13306);
xor U13423 (N_13423,N_13323,N_13362);
xnor U13424 (N_13424,N_13388,N_13230);
xor U13425 (N_13425,N_13335,N_13253);
nor U13426 (N_13426,N_13316,N_13302);
or U13427 (N_13427,N_13300,N_13288);
nand U13428 (N_13428,N_13282,N_13200);
nor U13429 (N_13429,N_13264,N_13356);
nand U13430 (N_13430,N_13394,N_13340);
or U13431 (N_13431,N_13204,N_13292);
nand U13432 (N_13432,N_13386,N_13374);
nor U13433 (N_13433,N_13219,N_13398);
nand U13434 (N_13434,N_13224,N_13220);
nand U13435 (N_13435,N_13370,N_13266);
xor U13436 (N_13436,N_13293,N_13265);
nand U13437 (N_13437,N_13389,N_13228);
and U13438 (N_13438,N_13232,N_13298);
nand U13439 (N_13439,N_13331,N_13247);
or U13440 (N_13440,N_13205,N_13343);
or U13441 (N_13441,N_13222,N_13327);
nor U13442 (N_13442,N_13202,N_13390);
xnor U13443 (N_13443,N_13260,N_13319);
or U13444 (N_13444,N_13256,N_13339);
nand U13445 (N_13445,N_13286,N_13216);
nand U13446 (N_13446,N_13274,N_13369);
nand U13447 (N_13447,N_13229,N_13254);
nor U13448 (N_13448,N_13249,N_13322);
or U13449 (N_13449,N_13372,N_13350);
xor U13450 (N_13450,N_13347,N_13295);
nor U13451 (N_13451,N_13294,N_13334);
nor U13452 (N_13452,N_13364,N_13373);
and U13453 (N_13453,N_13271,N_13239);
or U13454 (N_13454,N_13209,N_13259);
xnor U13455 (N_13455,N_13257,N_13312);
or U13456 (N_13456,N_13252,N_13221);
or U13457 (N_13457,N_13353,N_13344);
or U13458 (N_13458,N_13381,N_13255);
nand U13459 (N_13459,N_13337,N_13280);
nand U13460 (N_13460,N_13384,N_13336);
and U13461 (N_13461,N_13355,N_13285);
nand U13462 (N_13462,N_13234,N_13368);
nand U13463 (N_13463,N_13395,N_13301);
xor U13464 (N_13464,N_13308,N_13279);
or U13465 (N_13465,N_13315,N_13396);
nand U13466 (N_13466,N_13236,N_13248);
and U13467 (N_13467,N_13251,N_13211);
nand U13468 (N_13468,N_13367,N_13358);
xor U13469 (N_13469,N_13329,N_13289);
and U13470 (N_13470,N_13318,N_13349);
or U13471 (N_13471,N_13297,N_13291);
xor U13472 (N_13472,N_13233,N_13341);
nand U13473 (N_13473,N_13314,N_13354);
or U13474 (N_13474,N_13237,N_13304);
nand U13475 (N_13475,N_13376,N_13393);
xnor U13476 (N_13476,N_13240,N_13250);
nor U13477 (N_13477,N_13348,N_13338);
nand U13478 (N_13478,N_13360,N_13321);
xor U13479 (N_13479,N_13207,N_13272);
or U13480 (N_13480,N_13307,N_13243);
xor U13481 (N_13481,N_13214,N_13244);
or U13482 (N_13482,N_13399,N_13281);
xnor U13483 (N_13483,N_13371,N_13303);
nand U13484 (N_13484,N_13226,N_13277);
nand U13485 (N_13485,N_13379,N_13290);
xnor U13486 (N_13486,N_13242,N_13299);
or U13487 (N_13487,N_13332,N_13325);
or U13488 (N_13488,N_13313,N_13212);
xnor U13489 (N_13489,N_13363,N_13311);
xor U13490 (N_13490,N_13238,N_13245);
xor U13491 (N_13491,N_13262,N_13320);
nand U13492 (N_13492,N_13296,N_13267);
and U13493 (N_13493,N_13309,N_13269);
and U13494 (N_13494,N_13241,N_13378);
and U13495 (N_13495,N_13213,N_13310);
and U13496 (N_13496,N_13385,N_13268);
and U13497 (N_13497,N_13383,N_13366);
nor U13498 (N_13498,N_13317,N_13365);
and U13499 (N_13499,N_13278,N_13324);
nand U13500 (N_13500,N_13237,N_13294);
xor U13501 (N_13501,N_13337,N_13398);
or U13502 (N_13502,N_13245,N_13304);
and U13503 (N_13503,N_13270,N_13301);
nand U13504 (N_13504,N_13275,N_13344);
or U13505 (N_13505,N_13347,N_13387);
xnor U13506 (N_13506,N_13382,N_13248);
nand U13507 (N_13507,N_13234,N_13274);
or U13508 (N_13508,N_13242,N_13313);
xnor U13509 (N_13509,N_13201,N_13322);
nor U13510 (N_13510,N_13264,N_13232);
nand U13511 (N_13511,N_13280,N_13380);
or U13512 (N_13512,N_13355,N_13348);
or U13513 (N_13513,N_13342,N_13232);
xor U13514 (N_13514,N_13361,N_13383);
and U13515 (N_13515,N_13272,N_13269);
and U13516 (N_13516,N_13296,N_13361);
nor U13517 (N_13517,N_13379,N_13316);
xnor U13518 (N_13518,N_13391,N_13371);
nand U13519 (N_13519,N_13335,N_13215);
or U13520 (N_13520,N_13379,N_13388);
nand U13521 (N_13521,N_13397,N_13376);
nor U13522 (N_13522,N_13274,N_13381);
nand U13523 (N_13523,N_13387,N_13343);
or U13524 (N_13524,N_13313,N_13374);
nand U13525 (N_13525,N_13291,N_13325);
nand U13526 (N_13526,N_13270,N_13387);
nor U13527 (N_13527,N_13224,N_13345);
nor U13528 (N_13528,N_13259,N_13331);
nand U13529 (N_13529,N_13357,N_13286);
nand U13530 (N_13530,N_13345,N_13219);
or U13531 (N_13531,N_13303,N_13209);
nor U13532 (N_13532,N_13304,N_13321);
nor U13533 (N_13533,N_13204,N_13262);
or U13534 (N_13534,N_13343,N_13253);
xnor U13535 (N_13535,N_13271,N_13365);
nor U13536 (N_13536,N_13242,N_13315);
nor U13537 (N_13537,N_13216,N_13232);
nor U13538 (N_13538,N_13234,N_13272);
nor U13539 (N_13539,N_13238,N_13352);
nor U13540 (N_13540,N_13380,N_13315);
or U13541 (N_13541,N_13381,N_13219);
or U13542 (N_13542,N_13303,N_13391);
and U13543 (N_13543,N_13321,N_13278);
or U13544 (N_13544,N_13248,N_13283);
or U13545 (N_13545,N_13387,N_13221);
or U13546 (N_13546,N_13318,N_13389);
xor U13547 (N_13547,N_13391,N_13264);
and U13548 (N_13548,N_13346,N_13398);
or U13549 (N_13549,N_13331,N_13385);
and U13550 (N_13550,N_13201,N_13386);
and U13551 (N_13551,N_13203,N_13299);
xnor U13552 (N_13552,N_13237,N_13218);
or U13553 (N_13553,N_13225,N_13209);
and U13554 (N_13554,N_13206,N_13363);
and U13555 (N_13555,N_13311,N_13373);
xor U13556 (N_13556,N_13317,N_13343);
nand U13557 (N_13557,N_13229,N_13393);
or U13558 (N_13558,N_13256,N_13235);
or U13559 (N_13559,N_13308,N_13392);
xnor U13560 (N_13560,N_13282,N_13251);
or U13561 (N_13561,N_13247,N_13235);
nor U13562 (N_13562,N_13352,N_13315);
xor U13563 (N_13563,N_13201,N_13262);
or U13564 (N_13564,N_13368,N_13243);
or U13565 (N_13565,N_13339,N_13323);
xnor U13566 (N_13566,N_13213,N_13246);
and U13567 (N_13567,N_13243,N_13373);
xor U13568 (N_13568,N_13292,N_13373);
nand U13569 (N_13569,N_13375,N_13253);
and U13570 (N_13570,N_13362,N_13266);
nor U13571 (N_13571,N_13360,N_13201);
or U13572 (N_13572,N_13223,N_13332);
or U13573 (N_13573,N_13311,N_13318);
nor U13574 (N_13574,N_13344,N_13349);
or U13575 (N_13575,N_13386,N_13223);
nor U13576 (N_13576,N_13357,N_13389);
nor U13577 (N_13577,N_13321,N_13333);
nand U13578 (N_13578,N_13227,N_13267);
nor U13579 (N_13579,N_13341,N_13394);
and U13580 (N_13580,N_13297,N_13369);
and U13581 (N_13581,N_13275,N_13205);
or U13582 (N_13582,N_13319,N_13287);
nor U13583 (N_13583,N_13395,N_13389);
and U13584 (N_13584,N_13241,N_13337);
nor U13585 (N_13585,N_13256,N_13376);
xor U13586 (N_13586,N_13389,N_13398);
and U13587 (N_13587,N_13361,N_13322);
nand U13588 (N_13588,N_13361,N_13390);
and U13589 (N_13589,N_13368,N_13257);
xnor U13590 (N_13590,N_13285,N_13368);
and U13591 (N_13591,N_13221,N_13392);
or U13592 (N_13592,N_13360,N_13311);
and U13593 (N_13593,N_13271,N_13371);
and U13594 (N_13594,N_13362,N_13360);
nor U13595 (N_13595,N_13278,N_13380);
xor U13596 (N_13596,N_13386,N_13227);
nand U13597 (N_13597,N_13295,N_13398);
xor U13598 (N_13598,N_13314,N_13255);
nor U13599 (N_13599,N_13266,N_13398);
or U13600 (N_13600,N_13472,N_13479);
xor U13601 (N_13601,N_13489,N_13585);
and U13602 (N_13602,N_13471,N_13475);
xnor U13603 (N_13603,N_13454,N_13430);
nand U13604 (N_13604,N_13488,N_13580);
nor U13605 (N_13605,N_13405,N_13566);
or U13606 (N_13606,N_13438,N_13451);
and U13607 (N_13607,N_13443,N_13495);
or U13608 (N_13608,N_13450,N_13587);
xor U13609 (N_13609,N_13555,N_13568);
nand U13610 (N_13610,N_13499,N_13422);
xnor U13611 (N_13611,N_13485,N_13403);
xor U13612 (N_13612,N_13433,N_13515);
and U13613 (N_13613,N_13426,N_13462);
and U13614 (N_13614,N_13506,N_13458);
and U13615 (N_13615,N_13514,N_13494);
nor U13616 (N_13616,N_13464,N_13554);
or U13617 (N_13617,N_13551,N_13559);
xnor U13618 (N_13618,N_13572,N_13571);
nor U13619 (N_13619,N_13511,N_13440);
nand U13620 (N_13620,N_13500,N_13432);
nor U13621 (N_13621,N_13498,N_13492);
nand U13622 (N_13622,N_13546,N_13519);
nor U13623 (N_13623,N_13524,N_13549);
nand U13624 (N_13624,N_13463,N_13491);
and U13625 (N_13625,N_13595,N_13408);
or U13626 (N_13626,N_13547,N_13483);
nor U13627 (N_13627,N_13477,N_13532);
and U13628 (N_13628,N_13482,N_13556);
nand U13629 (N_13629,N_13558,N_13428);
nor U13630 (N_13630,N_13545,N_13493);
nand U13631 (N_13631,N_13529,N_13550);
and U13632 (N_13632,N_13552,N_13570);
xor U13633 (N_13633,N_13419,N_13478);
xnor U13634 (N_13634,N_13468,N_13518);
and U13635 (N_13635,N_13502,N_13473);
nor U13636 (N_13636,N_13431,N_13577);
and U13637 (N_13637,N_13588,N_13581);
xor U13638 (N_13638,N_13429,N_13578);
or U13639 (N_13639,N_13423,N_13439);
nor U13640 (N_13640,N_13575,N_13560);
nor U13641 (N_13641,N_13427,N_13593);
xnor U13642 (N_13642,N_13448,N_13536);
xor U13643 (N_13643,N_13574,N_13548);
nand U13644 (N_13644,N_13533,N_13516);
and U13645 (N_13645,N_13517,N_13467);
xnor U13646 (N_13646,N_13481,N_13437);
and U13647 (N_13647,N_13424,N_13401);
or U13648 (N_13648,N_13522,N_13459);
and U13649 (N_13649,N_13525,N_13508);
and U13650 (N_13650,N_13456,N_13460);
nor U13651 (N_13651,N_13597,N_13410);
or U13652 (N_13652,N_13445,N_13404);
or U13653 (N_13653,N_13444,N_13461);
or U13654 (N_13654,N_13531,N_13591);
and U13655 (N_13655,N_13469,N_13453);
or U13656 (N_13656,N_13496,N_13474);
nand U13657 (N_13657,N_13513,N_13447);
xor U13658 (N_13658,N_13407,N_13527);
or U13659 (N_13659,N_13490,N_13598);
or U13660 (N_13660,N_13567,N_13402);
nand U13661 (N_13661,N_13586,N_13435);
nor U13662 (N_13662,N_13563,N_13539);
or U13663 (N_13663,N_13530,N_13557);
xnor U13664 (N_13664,N_13409,N_13512);
or U13665 (N_13665,N_13504,N_13418);
xnor U13666 (N_13666,N_13579,N_13582);
nand U13667 (N_13667,N_13564,N_13420);
nor U13668 (N_13668,N_13434,N_13484);
and U13669 (N_13669,N_13411,N_13592);
nand U13670 (N_13670,N_13505,N_13520);
xor U13671 (N_13671,N_13449,N_13521);
nor U13672 (N_13672,N_13415,N_13470);
nor U13673 (N_13673,N_13501,N_13466);
nor U13674 (N_13674,N_13446,N_13486);
or U13675 (N_13675,N_13457,N_13526);
and U13676 (N_13676,N_13476,N_13565);
xor U13677 (N_13677,N_13503,N_13590);
xor U13678 (N_13678,N_13510,N_13507);
nor U13679 (N_13679,N_13561,N_13425);
nor U13680 (N_13680,N_13417,N_13562);
xor U13681 (N_13681,N_13487,N_13441);
nor U13682 (N_13682,N_13596,N_13535);
and U13683 (N_13683,N_13414,N_13465);
or U13684 (N_13684,N_13480,N_13589);
xnor U13685 (N_13685,N_13436,N_13537);
nor U13686 (N_13686,N_13455,N_13583);
and U13687 (N_13687,N_13413,N_13442);
xnor U13688 (N_13688,N_13576,N_13544);
nor U13689 (N_13689,N_13540,N_13412);
or U13690 (N_13690,N_13523,N_13599);
and U13691 (N_13691,N_13421,N_13569);
nor U13692 (N_13692,N_13584,N_13406);
nor U13693 (N_13693,N_13452,N_13528);
nor U13694 (N_13694,N_13594,N_13553);
nand U13695 (N_13695,N_13573,N_13542);
xnor U13696 (N_13696,N_13400,N_13509);
nor U13697 (N_13697,N_13534,N_13497);
and U13698 (N_13698,N_13543,N_13538);
nor U13699 (N_13699,N_13541,N_13416);
and U13700 (N_13700,N_13442,N_13481);
nor U13701 (N_13701,N_13451,N_13548);
or U13702 (N_13702,N_13508,N_13461);
nor U13703 (N_13703,N_13448,N_13566);
and U13704 (N_13704,N_13554,N_13530);
or U13705 (N_13705,N_13473,N_13416);
or U13706 (N_13706,N_13431,N_13495);
or U13707 (N_13707,N_13459,N_13536);
or U13708 (N_13708,N_13401,N_13433);
and U13709 (N_13709,N_13488,N_13558);
xnor U13710 (N_13710,N_13433,N_13426);
or U13711 (N_13711,N_13524,N_13400);
nand U13712 (N_13712,N_13406,N_13472);
and U13713 (N_13713,N_13485,N_13447);
nand U13714 (N_13714,N_13510,N_13413);
nand U13715 (N_13715,N_13583,N_13458);
and U13716 (N_13716,N_13501,N_13419);
nor U13717 (N_13717,N_13553,N_13482);
and U13718 (N_13718,N_13522,N_13473);
xor U13719 (N_13719,N_13558,N_13490);
xor U13720 (N_13720,N_13427,N_13464);
or U13721 (N_13721,N_13450,N_13421);
xor U13722 (N_13722,N_13477,N_13507);
and U13723 (N_13723,N_13496,N_13561);
and U13724 (N_13724,N_13573,N_13554);
and U13725 (N_13725,N_13485,N_13475);
and U13726 (N_13726,N_13412,N_13534);
nand U13727 (N_13727,N_13518,N_13528);
nor U13728 (N_13728,N_13513,N_13473);
and U13729 (N_13729,N_13560,N_13500);
or U13730 (N_13730,N_13432,N_13497);
and U13731 (N_13731,N_13564,N_13585);
and U13732 (N_13732,N_13593,N_13536);
nand U13733 (N_13733,N_13576,N_13469);
and U13734 (N_13734,N_13534,N_13463);
nand U13735 (N_13735,N_13496,N_13597);
xnor U13736 (N_13736,N_13408,N_13507);
nor U13737 (N_13737,N_13518,N_13562);
xor U13738 (N_13738,N_13452,N_13548);
nor U13739 (N_13739,N_13514,N_13572);
nor U13740 (N_13740,N_13532,N_13402);
and U13741 (N_13741,N_13400,N_13438);
and U13742 (N_13742,N_13547,N_13567);
xnor U13743 (N_13743,N_13567,N_13459);
and U13744 (N_13744,N_13482,N_13513);
xnor U13745 (N_13745,N_13487,N_13575);
or U13746 (N_13746,N_13599,N_13557);
xor U13747 (N_13747,N_13567,N_13523);
and U13748 (N_13748,N_13405,N_13538);
and U13749 (N_13749,N_13592,N_13468);
nand U13750 (N_13750,N_13562,N_13580);
or U13751 (N_13751,N_13433,N_13418);
xnor U13752 (N_13752,N_13496,N_13542);
and U13753 (N_13753,N_13432,N_13469);
nand U13754 (N_13754,N_13559,N_13490);
nor U13755 (N_13755,N_13504,N_13524);
or U13756 (N_13756,N_13411,N_13539);
nor U13757 (N_13757,N_13499,N_13527);
nand U13758 (N_13758,N_13480,N_13501);
xnor U13759 (N_13759,N_13497,N_13496);
nand U13760 (N_13760,N_13503,N_13448);
nor U13761 (N_13761,N_13407,N_13439);
xnor U13762 (N_13762,N_13591,N_13540);
and U13763 (N_13763,N_13482,N_13425);
nand U13764 (N_13764,N_13506,N_13424);
xor U13765 (N_13765,N_13545,N_13490);
or U13766 (N_13766,N_13565,N_13448);
xor U13767 (N_13767,N_13475,N_13415);
and U13768 (N_13768,N_13539,N_13594);
xor U13769 (N_13769,N_13590,N_13514);
nand U13770 (N_13770,N_13402,N_13494);
or U13771 (N_13771,N_13500,N_13598);
and U13772 (N_13772,N_13449,N_13519);
xor U13773 (N_13773,N_13459,N_13423);
and U13774 (N_13774,N_13463,N_13413);
and U13775 (N_13775,N_13514,N_13554);
or U13776 (N_13776,N_13447,N_13499);
nor U13777 (N_13777,N_13469,N_13470);
nand U13778 (N_13778,N_13526,N_13484);
or U13779 (N_13779,N_13521,N_13469);
xor U13780 (N_13780,N_13579,N_13588);
nor U13781 (N_13781,N_13416,N_13579);
nor U13782 (N_13782,N_13539,N_13534);
nor U13783 (N_13783,N_13432,N_13450);
nor U13784 (N_13784,N_13463,N_13432);
nor U13785 (N_13785,N_13551,N_13415);
nor U13786 (N_13786,N_13588,N_13584);
xnor U13787 (N_13787,N_13496,N_13490);
nand U13788 (N_13788,N_13498,N_13543);
xor U13789 (N_13789,N_13523,N_13571);
nand U13790 (N_13790,N_13493,N_13566);
nor U13791 (N_13791,N_13596,N_13560);
nand U13792 (N_13792,N_13555,N_13412);
nand U13793 (N_13793,N_13406,N_13533);
nand U13794 (N_13794,N_13570,N_13544);
nand U13795 (N_13795,N_13425,N_13464);
nor U13796 (N_13796,N_13462,N_13571);
nand U13797 (N_13797,N_13475,N_13431);
nor U13798 (N_13798,N_13420,N_13525);
xor U13799 (N_13799,N_13506,N_13532);
or U13800 (N_13800,N_13666,N_13623);
or U13801 (N_13801,N_13751,N_13627);
nor U13802 (N_13802,N_13658,N_13639);
or U13803 (N_13803,N_13670,N_13711);
xnor U13804 (N_13804,N_13777,N_13667);
xor U13805 (N_13805,N_13741,N_13608);
and U13806 (N_13806,N_13668,N_13761);
and U13807 (N_13807,N_13774,N_13795);
and U13808 (N_13808,N_13674,N_13604);
xnor U13809 (N_13809,N_13675,N_13643);
nand U13810 (N_13810,N_13695,N_13747);
and U13811 (N_13811,N_13794,N_13651);
or U13812 (N_13812,N_13646,N_13681);
or U13813 (N_13813,N_13775,N_13657);
nand U13814 (N_13814,N_13776,N_13699);
or U13815 (N_13815,N_13697,N_13745);
or U13816 (N_13816,N_13626,N_13602);
nand U13817 (N_13817,N_13738,N_13728);
nor U13818 (N_13818,N_13678,N_13734);
and U13819 (N_13819,N_13625,N_13731);
nand U13820 (N_13820,N_13705,N_13750);
and U13821 (N_13821,N_13641,N_13630);
nor U13822 (N_13822,N_13661,N_13649);
or U13823 (N_13823,N_13732,N_13727);
or U13824 (N_13824,N_13790,N_13619);
xnor U13825 (N_13825,N_13621,N_13698);
nand U13826 (N_13826,N_13696,N_13700);
or U13827 (N_13827,N_13612,N_13720);
xor U13828 (N_13828,N_13671,N_13740);
or U13829 (N_13829,N_13605,N_13633);
and U13830 (N_13830,N_13615,N_13798);
nor U13831 (N_13831,N_13701,N_13781);
and U13832 (N_13832,N_13660,N_13760);
nand U13833 (N_13833,N_13616,N_13758);
nor U13834 (N_13834,N_13749,N_13632);
and U13835 (N_13835,N_13610,N_13736);
nor U13836 (N_13836,N_13769,N_13709);
and U13837 (N_13837,N_13694,N_13611);
nor U13838 (N_13838,N_13676,N_13680);
nand U13839 (N_13839,N_13702,N_13664);
nand U13840 (N_13840,N_13785,N_13692);
nand U13841 (N_13841,N_13725,N_13669);
or U13842 (N_13842,N_13723,N_13620);
nor U13843 (N_13843,N_13786,N_13659);
xnor U13844 (N_13844,N_13706,N_13782);
or U13845 (N_13845,N_13622,N_13679);
xnor U13846 (N_13846,N_13724,N_13772);
or U13847 (N_13847,N_13743,N_13744);
nor U13848 (N_13848,N_13756,N_13609);
or U13849 (N_13849,N_13644,N_13793);
xor U13850 (N_13850,N_13606,N_13716);
or U13851 (N_13851,N_13759,N_13682);
nand U13852 (N_13852,N_13719,N_13693);
or U13853 (N_13853,N_13607,N_13613);
or U13854 (N_13854,N_13665,N_13770);
or U13855 (N_13855,N_13757,N_13754);
nand U13856 (N_13856,N_13636,N_13746);
xnor U13857 (N_13857,N_13784,N_13642);
or U13858 (N_13858,N_13687,N_13788);
nor U13859 (N_13859,N_13708,N_13799);
nand U13860 (N_13860,N_13763,N_13653);
and U13861 (N_13861,N_13603,N_13647);
nor U13862 (N_13862,N_13710,N_13787);
nor U13863 (N_13863,N_13648,N_13766);
nor U13864 (N_13864,N_13650,N_13634);
nand U13865 (N_13865,N_13718,N_13635);
and U13866 (N_13866,N_13640,N_13614);
nor U13867 (N_13867,N_13739,N_13624);
or U13868 (N_13868,N_13655,N_13663);
xor U13869 (N_13869,N_13629,N_13689);
nand U13870 (N_13870,N_13673,N_13762);
xnor U13871 (N_13871,N_13737,N_13628);
nor U13872 (N_13872,N_13765,N_13733);
nor U13873 (N_13873,N_13780,N_13672);
and U13874 (N_13874,N_13637,N_13771);
or U13875 (N_13875,N_13729,N_13645);
nand U13876 (N_13876,N_13783,N_13755);
nand U13877 (N_13877,N_13791,N_13638);
xnor U13878 (N_13878,N_13730,N_13721);
nor U13879 (N_13879,N_13704,N_13789);
or U13880 (N_13880,N_13684,N_13714);
or U13881 (N_13881,N_13742,N_13601);
nor U13882 (N_13882,N_13764,N_13717);
xor U13883 (N_13883,N_13715,N_13712);
and U13884 (N_13884,N_13726,N_13600);
nand U13885 (N_13885,N_13691,N_13722);
or U13886 (N_13886,N_13748,N_13685);
and U13887 (N_13887,N_13618,N_13796);
nor U13888 (N_13888,N_13713,N_13768);
and U13889 (N_13889,N_13767,N_13688);
nor U13890 (N_13890,N_13683,N_13773);
nor U13891 (N_13891,N_13690,N_13753);
or U13892 (N_13892,N_13662,N_13654);
nand U13893 (N_13893,N_13735,N_13617);
or U13894 (N_13894,N_13797,N_13686);
nor U13895 (N_13895,N_13656,N_13703);
nand U13896 (N_13896,N_13707,N_13778);
nor U13897 (N_13897,N_13792,N_13752);
nor U13898 (N_13898,N_13779,N_13677);
and U13899 (N_13899,N_13631,N_13652);
or U13900 (N_13900,N_13644,N_13693);
and U13901 (N_13901,N_13614,N_13766);
or U13902 (N_13902,N_13758,N_13697);
nor U13903 (N_13903,N_13761,N_13701);
nor U13904 (N_13904,N_13600,N_13683);
nand U13905 (N_13905,N_13688,N_13630);
nand U13906 (N_13906,N_13740,N_13718);
nor U13907 (N_13907,N_13736,N_13659);
xor U13908 (N_13908,N_13625,N_13642);
nand U13909 (N_13909,N_13769,N_13641);
xor U13910 (N_13910,N_13766,N_13617);
or U13911 (N_13911,N_13711,N_13688);
or U13912 (N_13912,N_13677,N_13703);
nand U13913 (N_13913,N_13669,N_13774);
nor U13914 (N_13914,N_13678,N_13604);
or U13915 (N_13915,N_13773,N_13676);
or U13916 (N_13916,N_13698,N_13663);
or U13917 (N_13917,N_13668,N_13654);
nor U13918 (N_13918,N_13707,N_13726);
xor U13919 (N_13919,N_13698,N_13636);
nand U13920 (N_13920,N_13733,N_13647);
nor U13921 (N_13921,N_13615,N_13655);
nand U13922 (N_13922,N_13749,N_13786);
nor U13923 (N_13923,N_13668,N_13614);
nand U13924 (N_13924,N_13602,N_13769);
nor U13925 (N_13925,N_13724,N_13756);
or U13926 (N_13926,N_13748,N_13628);
or U13927 (N_13927,N_13661,N_13733);
and U13928 (N_13928,N_13600,N_13649);
nand U13929 (N_13929,N_13695,N_13772);
and U13930 (N_13930,N_13601,N_13776);
or U13931 (N_13931,N_13713,N_13709);
nand U13932 (N_13932,N_13684,N_13661);
xnor U13933 (N_13933,N_13612,N_13699);
nand U13934 (N_13934,N_13698,N_13692);
nor U13935 (N_13935,N_13775,N_13669);
nor U13936 (N_13936,N_13606,N_13729);
xnor U13937 (N_13937,N_13617,N_13762);
nand U13938 (N_13938,N_13739,N_13774);
or U13939 (N_13939,N_13743,N_13701);
nor U13940 (N_13940,N_13680,N_13704);
nand U13941 (N_13941,N_13773,N_13630);
nor U13942 (N_13942,N_13776,N_13608);
and U13943 (N_13943,N_13674,N_13794);
xnor U13944 (N_13944,N_13618,N_13600);
nand U13945 (N_13945,N_13671,N_13722);
or U13946 (N_13946,N_13728,N_13648);
nand U13947 (N_13947,N_13666,N_13701);
and U13948 (N_13948,N_13667,N_13721);
nand U13949 (N_13949,N_13656,N_13671);
nand U13950 (N_13950,N_13729,N_13735);
xor U13951 (N_13951,N_13728,N_13680);
xor U13952 (N_13952,N_13612,N_13731);
nor U13953 (N_13953,N_13752,N_13795);
xor U13954 (N_13954,N_13750,N_13741);
and U13955 (N_13955,N_13621,N_13756);
or U13956 (N_13956,N_13793,N_13647);
or U13957 (N_13957,N_13712,N_13783);
xnor U13958 (N_13958,N_13687,N_13756);
or U13959 (N_13959,N_13752,N_13788);
nor U13960 (N_13960,N_13797,N_13654);
nor U13961 (N_13961,N_13668,N_13656);
xor U13962 (N_13962,N_13706,N_13630);
and U13963 (N_13963,N_13649,N_13754);
nor U13964 (N_13964,N_13776,N_13694);
and U13965 (N_13965,N_13730,N_13714);
and U13966 (N_13966,N_13673,N_13661);
nor U13967 (N_13967,N_13726,N_13670);
xor U13968 (N_13968,N_13685,N_13683);
nand U13969 (N_13969,N_13698,N_13750);
xor U13970 (N_13970,N_13708,N_13633);
nand U13971 (N_13971,N_13738,N_13623);
nand U13972 (N_13972,N_13701,N_13703);
or U13973 (N_13973,N_13704,N_13644);
and U13974 (N_13974,N_13613,N_13642);
and U13975 (N_13975,N_13785,N_13632);
nand U13976 (N_13976,N_13632,N_13686);
xor U13977 (N_13977,N_13620,N_13693);
nor U13978 (N_13978,N_13620,N_13702);
nand U13979 (N_13979,N_13755,N_13728);
nor U13980 (N_13980,N_13649,N_13747);
nand U13981 (N_13981,N_13635,N_13727);
nand U13982 (N_13982,N_13726,N_13720);
xor U13983 (N_13983,N_13723,N_13643);
and U13984 (N_13984,N_13670,N_13777);
nand U13985 (N_13985,N_13626,N_13787);
nor U13986 (N_13986,N_13679,N_13746);
nand U13987 (N_13987,N_13677,N_13777);
nor U13988 (N_13988,N_13713,N_13725);
nand U13989 (N_13989,N_13608,N_13616);
nor U13990 (N_13990,N_13792,N_13656);
or U13991 (N_13991,N_13688,N_13677);
or U13992 (N_13992,N_13752,N_13607);
nor U13993 (N_13993,N_13742,N_13772);
nand U13994 (N_13994,N_13643,N_13630);
and U13995 (N_13995,N_13741,N_13740);
or U13996 (N_13996,N_13778,N_13704);
nor U13997 (N_13997,N_13784,N_13617);
xnor U13998 (N_13998,N_13689,N_13710);
xnor U13999 (N_13999,N_13652,N_13624);
nand U14000 (N_14000,N_13893,N_13935);
and U14001 (N_14001,N_13986,N_13804);
nand U14002 (N_14002,N_13852,N_13884);
or U14003 (N_14003,N_13947,N_13888);
and U14004 (N_14004,N_13818,N_13970);
xnor U14005 (N_14005,N_13922,N_13892);
nor U14006 (N_14006,N_13900,N_13927);
nor U14007 (N_14007,N_13955,N_13940);
or U14008 (N_14008,N_13913,N_13853);
xor U14009 (N_14009,N_13875,N_13857);
xor U14010 (N_14010,N_13824,N_13999);
nor U14011 (N_14011,N_13915,N_13863);
or U14012 (N_14012,N_13899,N_13815);
and U14013 (N_14013,N_13801,N_13904);
xor U14014 (N_14014,N_13805,N_13968);
or U14015 (N_14015,N_13943,N_13909);
and U14016 (N_14016,N_13994,N_13916);
xnor U14017 (N_14017,N_13860,N_13845);
nand U14018 (N_14018,N_13856,N_13836);
or U14019 (N_14019,N_13880,N_13809);
and U14020 (N_14020,N_13847,N_13978);
and U14021 (N_14021,N_13816,N_13918);
nand U14022 (N_14022,N_13972,N_13907);
nor U14023 (N_14023,N_13969,N_13963);
nand U14024 (N_14024,N_13912,N_13841);
nand U14025 (N_14025,N_13976,N_13806);
or U14026 (N_14026,N_13830,N_13924);
nand U14027 (N_14027,N_13903,N_13842);
or U14028 (N_14028,N_13967,N_13944);
xnor U14029 (N_14029,N_13862,N_13866);
nor U14030 (N_14030,N_13835,N_13973);
nor U14031 (N_14031,N_13960,N_13920);
or U14032 (N_14032,N_13895,N_13854);
nand U14033 (N_14033,N_13810,N_13929);
nand U14034 (N_14034,N_13873,N_13989);
and U14035 (N_14035,N_13933,N_13825);
nand U14036 (N_14036,N_13984,N_13951);
nor U14037 (N_14037,N_13829,N_13874);
and U14038 (N_14038,N_13908,N_13870);
or U14039 (N_14039,N_13838,N_13872);
and U14040 (N_14040,N_13931,N_13998);
and U14041 (N_14041,N_13941,N_13821);
nor U14042 (N_14042,N_13983,N_13966);
or U14043 (N_14043,N_13831,N_13822);
or U14044 (N_14044,N_13932,N_13921);
nor U14045 (N_14045,N_13877,N_13811);
xor U14046 (N_14046,N_13869,N_13991);
nor U14047 (N_14047,N_13982,N_13819);
nand U14048 (N_14048,N_13923,N_13887);
or U14049 (N_14049,N_13981,N_13987);
and U14050 (N_14050,N_13925,N_13910);
or U14051 (N_14051,N_13988,N_13843);
or U14052 (N_14052,N_13800,N_13889);
or U14053 (N_14053,N_13846,N_13848);
xor U14054 (N_14054,N_13997,N_13855);
nand U14055 (N_14055,N_13990,N_13861);
nand U14056 (N_14056,N_13864,N_13917);
or U14057 (N_14057,N_13992,N_13979);
xor U14058 (N_14058,N_13890,N_13993);
or U14059 (N_14059,N_13839,N_13911);
or U14060 (N_14060,N_13956,N_13803);
and U14061 (N_14061,N_13939,N_13868);
and U14062 (N_14062,N_13958,N_13820);
nor U14063 (N_14063,N_13977,N_13882);
xor U14064 (N_14064,N_13948,N_13928);
xnor U14065 (N_14065,N_13826,N_13971);
and U14066 (N_14066,N_13914,N_13949);
or U14067 (N_14067,N_13885,N_13942);
nand U14068 (N_14068,N_13946,N_13813);
or U14069 (N_14069,N_13891,N_13926);
and U14070 (N_14070,N_13980,N_13867);
nor U14071 (N_14071,N_13954,N_13901);
or U14072 (N_14072,N_13844,N_13812);
nor U14073 (N_14073,N_13837,N_13965);
nand U14074 (N_14074,N_13883,N_13957);
xnor U14075 (N_14075,N_13902,N_13961);
nor U14076 (N_14076,N_13950,N_13814);
xnor U14077 (N_14077,N_13871,N_13985);
or U14078 (N_14078,N_13930,N_13938);
nand U14079 (N_14079,N_13851,N_13876);
nand U14080 (N_14080,N_13996,N_13840);
or U14081 (N_14081,N_13832,N_13897);
nand U14082 (N_14082,N_13934,N_13896);
xor U14083 (N_14083,N_13886,N_13859);
and U14084 (N_14084,N_13833,N_13905);
xnor U14085 (N_14085,N_13879,N_13849);
nand U14086 (N_14086,N_13802,N_13962);
and U14087 (N_14087,N_13817,N_13823);
and U14088 (N_14088,N_13881,N_13850);
nor U14089 (N_14089,N_13834,N_13858);
or U14090 (N_14090,N_13975,N_13959);
and U14091 (N_14091,N_13828,N_13964);
nand U14092 (N_14092,N_13827,N_13995);
nor U14093 (N_14093,N_13945,N_13878);
nand U14094 (N_14094,N_13898,N_13894);
and U14095 (N_14095,N_13865,N_13906);
nand U14096 (N_14096,N_13937,N_13974);
nor U14097 (N_14097,N_13952,N_13919);
or U14098 (N_14098,N_13936,N_13807);
or U14099 (N_14099,N_13953,N_13808);
xnor U14100 (N_14100,N_13995,N_13833);
nor U14101 (N_14101,N_13945,N_13968);
nand U14102 (N_14102,N_13978,N_13841);
nor U14103 (N_14103,N_13806,N_13948);
nor U14104 (N_14104,N_13812,N_13843);
and U14105 (N_14105,N_13882,N_13975);
nand U14106 (N_14106,N_13895,N_13971);
xor U14107 (N_14107,N_13993,N_13970);
nand U14108 (N_14108,N_13832,N_13931);
xnor U14109 (N_14109,N_13993,N_13880);
or U14110 (N_14110,N_13914,N_13966);
nand U14111 (N_14111,N_13847,N_13855);
or U14112 (N_14112,N_13984,N_13822);
nand U14113 (N_14113,N_13916,N_13966);
nor U14114 (N_14114,N_13982,N_13936);
nand U14115 (N_14115,N_13828,N_13938);
and U14116 (N_14116,N_13965,N_13988);
nor U14117 (N_14117,N_13943,N_13833);
and U14118 (N_14118,N_13863,N_13974);
and U14119 (N_14119,N_13907,N_13895);
and U14120 (N_14120,N_13982,N_13879);
and U14121 (N_14121,N_13987,N_13911);
or U14122 (N_14122,N_13984,N_13863);
or U14123 (N_14123,N_13989,N_13835);
nor U14124 (N_14124,N_13818,N_13878);
nand U14125 (N_14125,N_13854,N_13980);
xnor U14126 (N_14126,N_13882,N_13859);
nor U14127 (N_14127,N_13835,N_13932);
nor U14128 (N_14128,N_13896,N_13989);
nor U14129 (N_14129,N_13977,N_13812);
nand U14130 (N_14130,N_13945,N_13857);
nand U14131 (N_14131,N_13992,N_13823);
nor U14132 (N_14132,N_13948,N_13879);
nor U14133 (N_14133,N_13975,N_13877);
xnor U14134 (N_14134,N_13863,N_13819);
xor U14135 (N_14135,N_13957,N_13804);
and U14136 (N_14136,N_13996,N_13807);
nand U14137 (N_14137,N_13989,N_13984);
nor U14138 (N_14138,N_13841,N_13995);
or U14139 (N_14139,N_13907,N_13836);
and U14140 (N_14140,N_13899,N_13914);
xnor U14141 (N_14141,N_13966,N_13929);
and U14142 (N_14142,N_13971,N_13972);
or U14143 (N_14143,N_13920,N_13866);
nor U14144 (N_14144,N_13948,N_13891);
or U14145 (N_14145,N_13801,N_13810);
or U14146 (N_14146,N_13945,N_13880);
nor U14147 (N_14147,N_13978,N_13901);
nor U14148 (N_14148,N_13916,N_13987);
or U14149 (N_14149,N_13988,N_13882);
and U14150 (N_14150,N_13962,N_13855);
nand U14151 (N_14151,N_13970,N_13932);
or U14152 (N_14152,N_13948,N_13973);
xnor U14153 (N_14153,N_13895,N_13959);
and U14154 (N_14154,N_13949,N_13994);
or U14155 (N_14155,N_13928,N_13880);
nor U14156 (N_14156,N_13902,N_13854);
nor U14157 (N_14157,N_13982,N_13994);
or U14158 (N_14158,N_13878,N_13897);
nor U14159 (N_14159,N_13988,N_13907);
nor U14160 (N_14160,N_13945,N_13822);
nor U14161 (N_14161,N_13968,N_13885);
nand U14162 (N_14162,N_13903,N_13949);
xnor U14163 (N_14163,N_13930,N_13902);
or U14164 (N_14164,N_13852,N_13914);
nand U14165 (N_14165,N_13897,N_13824);
or U14166 (N_14166,N_13909,N_13806);
nor U14167 (N_14167,N_13828,N_13918);
nor U14168 (N_14168,N_13981,N_13892);
xor U14169 (N_14169,N_13943,N_13824);
or U14170 (N_14170,N_13866,N_13909);
or U14171 (N_14171,N_13800,N_13851);
nor U14172 (N_14172,N_13857,N_13961);
nand U14173 (N_14173,N_13853,N_13994);
and U14174 (N_14174,N_13930,N_13803);
nor U14175 (N_14175,N_13900,N_13951);
xnor U14176 (N_14176,N_13839,N_13933);
nor U14177 (N_14177,N_13976,N_13851);
nor U14178 (N_14178,N_13863,N_13922);
nor U14179 (N_14179,N_13971,N_13954);
nand U14180 (N_14180,N_13958,N_13856);
or U14181 (N_14181,N_13865,N_13879);
nor U14182 (N_14182,N_13831,N_13914);
or U14183 (N_14183,N_13819,N_13854);
and U14184 (N_14184,N_13984,N_13844);
xnor U14185 (N_14185,N_13989,N_13800);
nand U14186 (N_14186,N_13936,N_13803);
nand U14187 (N_14187,N_13872,N_13933);
or U14188 (N_14188,N_13909,N_13844);
nor U14189 (N_14189,N_13908,N_13802);
xnor U14190 (N_14190,N_13941,N_13833);
nor U14191 (N_14191,N_13959,N_13912);
or U14192 (N_14192,N_13830,N_13872);
and U14193 (N_14193,N_13993,N_13867);
nand U14194 (N_14194,N_13864,N_13953);
and U14195 (N_14195,N_13893,N_13930);
nor U14196 (N_14196,N_13814,N_13991);
nor U14197 (N_14197,N_13920,N_13832);
xnor U14198 (N_14198,N_13979,N_13903);
and U14199 (N_14199,N_13908,N_13881);
nand U14200 (N_14200,N_14021,N_14107);
and U14201 (N_14201,N_14024,N_14053);
and U14202 (N_14202,N_14143,N_14169);
nand U14203 (N_14203,N_14076,N_14132);
xor U14204 (N_14204,N_14036,N_14046);
and U14205 (N_14205,N_14101,N_14002);
nor U14206 (N_14206,N_14114,N_14080);
xnor U14207 (N_14207,N_14019,N_14195);
or U14208 (N_14208,N_14042,N_14164);
or U14209 (N_14209,N_14057,N_14189);
and U14210 (N_14210,N_14193,N_14004);
and U14211 (N_14211,N_14069,N_14026);
or U14212 (N_14212,N_14064,N_14000);
xnor U14213 (N_14213,N_14075,N_14198);
nand U14214 (N_14214,N_14171,N_14194);
xnor U14215 (N_14215,N_14027,N_14056);
xnor U14216 (N_14216,N_14175,N_14172);
nor U14217 (N_14217,N_14054,N_14108);
xnor U14218 (N_14218,N_14095,N_14071);
nor U14219 (N_14219,N_14059,N_14181);
nor U14220 (N_14220,N_14050,N_14159);
nand U14221 (N_14221,N_14158,N_14082);
and U14222 (N_14222,N_14037,N_14131);
xor U14223 (N_14223,N_14190,N_14063);
and U14224 (N_14224,N_14188,N_14051);
xor U14225 (N_14225,N_14070,N_14003);
nor U14226 (N_14226,N_14178,N_14096);
nor U14227 (N_14227,N_14091,N_14090);
nor U14228 (N_14228,N_14162,N_14110);
nor U14229 (N_14229,N_14014,N_14136);
and U14230 (N_14230,N_14078,N_14166);
or U14231 (N_14231,N_14105,N_14129);
nor U14232 (N_14232,N_14119,N_14155);
xnor U14233 (N_14233,N_14160,N_14147);
xnor U14234 (N_14234,N_14066,N_14135);
nor U14235 (N_14235,N_14020,N_14140);
and U14236 (N_14236,N_14098,N_14030);
and U14237 (N_14237,N_14044,N_14170);
xnor U14238 (N_14238,N_14065,N_14009);
xnor U14239 (N_14239,N_14029,N_14097);
nand U14240 (N_14240,N_14123,N_14055);
xnor U14241 (N_14241,N_14137,N_14047);
and U14242 (N_14242,N_14127,N_14043);
xor U14243 (N_14243,N_14045,N_14111);
or U14244 (N_14244,N_14017,N_14049);
or U14245 (N_14245,N_14052,N_14102);
or U14246 (N_14246,N_14139,N_14034);
or U14247 (N_14247,N_14041,N_14118);
nor U14248 (N_14248,N_14035,N_14145);
and U14249 (N_14249,N_14073,N_14089);
nand U14250 (N_14250,N_14199,N_14077);
or U14251 (N_14251,N_14025,N_14163);
xor U14252 (N_14252,N_14109,N_14174);
or U14253 (N_14253,N_14022,N_14013);
and U14254 (N_14254,N_14005,N_14016);
nand U14255 (N_14255,N_14149,N_14150);
or U14256 (N_14256,N_14018,N_14072);
and U14257 (N_14257,N_14176,N_14134);
nand U14258 (N_14258,N_14039,N_14100);
xor U14259 (N_14259,N_14001,N_14006);
xnor U14260 (N_14260,N_14186,N_14165);
xnor U14261 (N_14261,N_14184,N_14128);
or U14262 (N_14262,N_14148,N_14130);
xnor U14263 (N_14263,N_14168,N_14141);
nand U14264 (N_14264,N_14125,N_14048);
or U14265 (N_14265,N_14106,N_14083);
nor U14266 (N_14266,N_14117,N_14023);
nand U14267 (N_14267,N_14104,N_14152);
xnor U14268 (N_14268,N_14144,N_14113);
nand U14269 (N_14269,N_14183,N_14093);
nor U14270 (N_14270,N_14116,N_14010);
xnor U14271 (N_14271,N_14173,N_14028);
and U14272 (N_14272,N_14038,N_14099);
nor U14273 (N_14273,N_14180,N_14032);
or U14274 (N_14274,N_14015,N_14031);
xnor U14275 (N_14275,N_14121,N_14007);
nor U14276 (N_14276,N_14068,N_14033);
and U14277 (N_14277,N_14085,N_14084);
xor U14278 (N_14278,N_14086,N_14191);
xor U14279 (N_14279,N_14196,N_14154);
or U14280 (N_14280,N_14185,N_14187);
nand U14281 (N_14281,N_14179,N_14088);
and U14282 (N_14282,N_14012,N_14120);
and U14283 (N_14283,N_14011,N_14167);
nand U14284 (N_14284,N_14060,N_14103);
and U14285 (N_14285,N_14087,N_14079);
xor U14286 (N_14286,N_14074,N_14142);
and U14287 (N_14287,N_14197,N_14067);
xor U14288 (N_14288,N_14156,N_14115);
nor U14289 (N_14289,N_14008,N_14081);
xnor U14290 (N_14290,N_14161,N_14112);
xnor U14291 (N_14291,N_14122,N_14061);
xor U14292 (N_14292,N_14138,N_14192);
nand U14293 (N_14293,N_14133,N_14040);
or U14294 (N_14294,N_14126,N_14182);
xnor U14295 (N_14295,N_14124,N_14151);
nor U14296 (N_14296,N_14153,N_14146);
nor U14297 (N_14297,N_14058,N_14094);
and U14298 (N_14298,N_14062,N_14092);
and U14299 (N_14299,N_14177,N_14157);
and U14300 (N_14300,N_14017,N_14028);
xnor U14301 (N_14301,N_14109,N_14081);
nor U14302 (N_14302,N_14111,N_14130);
nor U14303 (N_14303,N_14048,N_14007);
nor U14304 (N_14304,N_14062,N_14186);
and U14305 (N_14305,N_14189,N_14168);
and U14306 (N_14306,N_14058,N_14138);
nor U14307 (N_14307,N_14139,N_14118);
nor U14308 (N_14308,N_14089,N_14054);
or U14309 (N_14309,N_14070,N_14167);
nor U14310 (N_14310,N_14112,N_14148);
nor U14311 (N_14311,N_14005,N_14148);
or U14312 (N_14312,N_14120,N_14075);
and U14313 (N_14313,N_14052,N_14007);
xor U14314 (N_14314,N_14009,N_14191);
and U14315 (N_14315,N_14087,N_14104);
or U14316 (N_14316,N_14125,N_14083);
and U14317 (N_14317,N_14164,N_14185);
nor U14318 (N_14318,N_14006,N_14038);
nor U14319 (N_14319,N_14061,N_14194);
and U14320 (N_14320,N_14078,N_14197);
xnor U14321 (N_14321,N_14196,N_14021);
or U14322 (N_14322,N_14179,N_14125);
nand U14323 (N_14323,N_14101,N_14019);
and U14324 (N_14324,N_14110,N_14197);
or U14325 (N_14325,N_14199,N_14115);
nand U14326 (N_14326,N_14047,N_14005);
nand U14327 (N_14327,N_14100,N_14129);
xor U14328 (N_14328,N_14004,N_14009);
nand U14329 (N_14329,N_14074,N_14000);
or U14330 (N_14330,N_14141,N_14115);
and U14331 (N_14331,N_14085,N_14145);
nand U14332 (N_14332,N_14045,N_14060);
and U14333 (N_14333,N_14090,N_14096);
or U14334 (N_14334,N_14142,N_14055);
xor U14335 (N_14335,N_14183,N_14078);
and U14336 (N_14336,N_14110,N_14106);
or U14337 (N_14337,N_14044,N_14090);
xor U14338 (N_14338,N_14169,N_14054);
and U14339 (N_14339,N_14083,N_14095);
xor U14340 (N_14340,N_14189,N_14047);
nor U14341 (N_14341,N_14167,N_14042);
xnor U14342 (N_14342,N_14013,N_14075);
nand U14343 (N_14343,N_14164,N_14130);
nor U14344 (N_14344,N_14169,N_14027);
xor U14345 (N_14345,N_14133,N_14185);
nand U14346 (N_14346,N_14120,N_14156);
or U14347 (N_14347,N_14163,N_14185);
nand U14348 (N_14348,N_14062,N_14113);
and U14349 (N_14349,N_14098,N_14108);
and U14350 (N_14350,N_14076,N_14135);
xor U14351 (N_14351,N_14190,N_14001);
nand U14352 (N_14352,N_14166,N_14137);
nor U14353 (N_14353,N_14061,N_14015);
and U14354 (N_14354,N_14031,N_14187);
nor U14355 (N_14355,N_14048,N_14121);
or U14356 (N_14356,N_14195,N_14099);
or U14357 (N_14357,N_14020,N_14178);
and U14358 (N_14358,N_14182,N_14145);
xnor U14359 (N_14359,N_14080,N_14181);
and U14360 (N_14360,N_14020,N_14074);
nand U14361 (N_14361,N_14029,N_14121);
nor U14362 (N_14362,N_14047,N_14067);
xor U14363 (N_14363,N_14132,N_14041);
xnor U14364 (N_14364,N_14046,N_14146);
or U14365 (N_14365,N_14026,N_14030);
or U14366 (N_14366,N_14014,N_14079);
or U14367 (N_14367,N_14144,N_14049);
or U14368 (N_14368,N_14116,N_14126);
nor U14369 (N_14369,N_14133,N_14178);
nor U14370 (N_14370,N_14143,N_14167);
or U14371 (N_14371,N_14034,N_14118);
or U14372 (N_14372,N_14166,N_14163);
or U14373 (N_14373,N_14046,N_14013);
or U14374 (N_14374,N_14116,N_14111);
nor U14375 (N_14375,N_14017,N_14145);
and U14376 (N_14376,N_14066,N_14030);
and U14377 (N_14377,N_14029,N_14106);
nor U14378 (N_14378,N_14090,N_14081);
and U14379 (N_14379,N_14158,N_14052);
or U14380 (N_14380,N_14093,N_14080);
nand U14381 (N_14381,N_14165,N_14148);
and U14382 (N_14382,N_14085,N_14111);
and U14383 (N_14383,N_14016,N_14115);
xor U14384 (N_14384,N_14016,N_14101);
nand U14385 (N_14385,N_14083,N_14182);
nor U14386 (N_14386,N_14122,N_14130);
nor U14387 (N_14387,N_14143,N_14078);
and U14388 (N_14388,N_14159,N_14040);
or U14389 (N_14389,N_14107,N_14003);
xor U14390 (N_14390,N_14021,N_14063);
nand U14391 (N_14391,N_14087,N_14125);
and U14392 (N_14392,N_14103,N_14143);
and U14393 (N_14393,N_14133,N_14076);
nor U14394 (N_14394,N_14077,N_14025);
xnor U14395 (N_14395,N_14065,N_14139);
and U14396 (N_14396,N_14014,N_14115);
nor U14397 (N_14397,N_14130,N_14065);
xnor U14398 (N_14398,N_14038,N_14094);
xor U14399 (N_14399,N_14082,N_14094);
nand U14400 (N_14400,N_14336,N_14382);
nor U14401 (N_14401,N_14377,N_14335);
xor U14402 (N_14402,N_14272,N_14303);
or U14403 (N_14403,N_14386,N_14290);
or U14404 (N_14404,N_14304,N_14298);
and U14405 (N_14405,N_14380,N_14326);
or U14406 (N_14406,N_14322,N_14393);
xnor U14407 (N_14407,N_14242,N_14338);
xor U14408 (N_14408,N_14390,N_14247);
nand U14409 (N_14409,N_14324,N_14256);
or U14410 (N_14410,N_14277,N_14248);
xor U14411 (N_14411,N_14399,N_14270);
xnor U14412 (N_14412,N_14346,N_14226);
nor U14413 (N_14413,N_14325,N_14213);
and U14414 (N_14414,N_14251,N_14265);
and U14415 (N_14415,N_14269,N_14327);
and U14416 (N_14416,N_14207,N_14315);
nand U14417 (N_14417,N_14283,N_14358);
or U14418 (N_14418,N_14359,N_14373);
and U14419 (N_14419,N_14218,N_14212);
xnor U14420 (N_14420,N_14253,N_14299);
or U14421 (N_14421,N_14246,N_14287);
nor U14422 (N_14422,N_14214,N_14211);
or U14423 (N_14423,N_14289,N_14334);
and U14424 (N_14424,N_14329,N_14293);
and U14425 (N_14425,N_14232,N_14309);
xnor U14426 (N_14426,N_14233,N_14361);
and U14427 (N_14427,N_14305,N_14268);
xnor U14428 (N_14428,N_14220,N_14343);
or U14429 (N_14429,N_14202,N_14347);
nor U14430 (N_14430,N_14206,N_14267);
and U14431 (N_14431,N_14344,N_14281);
xnor U14432 (N_14432,N_14271,N_14200);
or U14433 (N_14433,N_14376,N_14208);
and U14434 (N_14434,N_14288,N_14294);
and U14435 (N_14435,N_14307,N_14262);
and U14436 (N_14436,N_14222,N_14254);
xnor U14437 (N_14437,N_14229,N_14260);
or U14438 (N_14438,N_14363,N_14286);
or U14439 (N_14439,N_14278,N_14204);
or U14440 (N_14440,N_14354,N_14261);
or U14441 (N_14441,N_14319,N_14342);
and U14442 (N_14442,N_14350,N_14371);
xnor U14443 (N_14443,N_14209,N_14235);
xnor U14444 (N_14444,N_14317,N_14306);
xor U14445 (N_14445,N_14215,N_14383);
and U14446 (N_14446,N_14321,N_14362);
xnor U14447 (N_14447,N_14355,N_14366);
xnor U14448 (N_14448,N_14263,N_14273);
nand U14449 (N_14449,N_14302,N_14227);
nor U14450 (N_14450,N_14332,N_14291);
and U14451 (N_14451,N_14391,N_14374);
nor U14452 (N_14452,N_14387,N_14388);
nor U14453 (N_14453,N_14384,N_14238);
nor U14454 (N_14454,N_14244,N_14368);
xnor U14455 (N_14455,N_14234,N_14308);
or U14456 (N_14456,N_14210,N_14280);
nor U14457 (N_14457,N_14348,N_14240);
and U14458 (N_14458,N_14241,N_14351);
or U14459 (N_14459,N_14323,N_14300);
or U14460 (N_14460,N_14396,N_14340);
nor U14461 (N_14461,N_14360,N_14284);
or U14462 (N_14462,N_14345,N_14236);
and U14463 (N_14463,N_14341,N_14356);
nor U14464 (N_14464,N_14311,N_14274);
xnor U14465 (N_14465,N_14297,N_14301);
or U14466 (N_14466,N_14276,N_14398);
and U14467 (N_14467,N_14320,N_14367);
or U14468 (N_14468,N_14378,N_14352);
nor U14469 (N_14469,N_14252,N_14372);
nand U14470 (N_14470,N_14219,N_14225);
nand U14471 (N_14471,N_14279,N_14205);
xor U14472 (N_14472,N_14318,N_14385);
xnor U14473 (N_14473,N_14237,N_14369);
nand U14474 (N_14474,N_14394,N_14259);
and U14475 (N_14475,N_14264,N_14313);
and U14476 (N_14476,N_14243,N_14395);
nor U14477 (N_14477,N_14365,N_14257);
xnor U14478 (N_14478,N_14389,N_14310);
xnor U14479 (N_14479,N_14249,N_14203);
nor U14480 (N_14480,N_14231,N_14250);
xor U14481 (N_14481,N_14266,N_14333);
xnor U14482 (N_14482,N_14216,N_14217);
nand U14483 (N_14483,N_14282,N_14328);
and U14484 (N_14484,N_14296,N_14292);
xnor U14485 (N_14485,N_14223,N_14364);
and U14486 (N_14486,N_14397,N_14339);
and U14487 (N_14487,N_14239,N_14379);
xnor U14488 (N_14488,N_14224,N_14353);
nor U14489 (N_14489,N_14312,N_14392);
or U14490 (N_14490,N_14349,N_14221);
and U14491 (N_14491,N_14375,N_14228);
nor U14492 (N_14492,N_14331,N_14230);
xor U14493 (N_14493,N_14370,N_14201);
nor U14494 (N_14494,N_14255,N_14295);
nor U14495 (N_14495,N_14275,N_14357);
nor U14496 (N_14496,N_14314,N_14330);
nor U14497 (N_14497,N_14258,N_14245);
nand U14498 (N_14498,N_14337,N_14316);
nand U14499 (N_14499,N_14285,N_14381);
nand U14500 (N_14500,N_14379,N_14247);
xor U14501 (N_14501,N_14249,N_14286);
nor U14502 (N_14502,N_14385,N_14272);
nor U14503 (N_14503,N_14200,N_14267);
nand U14504 (N_14504,N_14342,N_14302);
nand U14505 (N_14505,N_14335,N_14261);
or U14506 (N_14506,N_14276,N_14310);
or U14507 (N_14507,N_14288,N_14395);
xnor U14508 (N_14508,N_14210,N_14232);
nand U14509 (N_14509,N_14374,N_14307);
and U14510 (N_14510,N_14286,N_14372);
nor U14511 (N_14511,N_14200,N_14218);
nand U14512 (N_14512,N_14268,N_14209);
and U14513 (N_14513,N_14309,N_14350);
or U14514 (N_14514,N_14371,N_14216);
nand U14515 (N_14515,N_14377,N_14315);
and U14516 (N_14516,N_14322,N_14239);
or U14517 (N_14517,N_14204,N_14395);
nand U14518 (N_14518,N_14208,N_14341);
and U14519 (N_14519,N_14393,N_14270);
xor U14520 (N_14520,N_14269,N_14220);
and U14521 (N_14521,N_14324,N_14382);
nand U14522 (N_14522,N_14386,N_14281);
nor U14523 (N_14523,N_14316,N_14292);
and U14524 (N_14524,N_14371,N_14221);
or U14525 (N_14525,N_14387,N_14299);
or U14526 (N_14526,N_14356,N_14359);
xnor U14527 (N_14527,N_14210,N_14383);
nand U14528 (N_14528,N_14352,N_14379);
nor U14529 (N_14529,N_14346,N_14237);
nand U14530 (N_14530,N_14228,N_14342);
nand U14531 (N_14531,N_14341,N_14223);
nand U14532 (N_14532,N_14293,N_14238);
xor U14533 (N_14533,N_14208,N_14232);
nand U14534 (N_14534,N_14225,N_14391);
nor U14535 (N_14535,N_14227,N_14313);
nand U14536 (N_14536,N_14267,N_14293);
xnor U14537 (N_14537,N_14311,N_14303);
xor U14538 (N_14538,N_14323,N_14308);
nand U14539 (N_14539,N_14324,N_14251);
nand U14540 (N_14540,N_14348,N_14278);
xnor U14541 (N_14541,N_14203,N_14294);
nor U14542 (N_14542,N_14265,N_14247);
or U14543 (N_14543,N_14276,N_14301);
nor U14544 (N_14544,N_14258,N_14267);
nor U14545 (N_14545,N_14218,N_14372);
xnor U14546 (N_14546,N_14249,N_14325);
or U14547 (N_14547,N_14316,N_14223);
nor U14548 (N_14548,N_14326,N_14384);
nor U14549 (N_14549,N_14299,N_14338);
and U14550 (N_14550,N_14298,N_14219);
xnor U14551 (N_14551,N_14252,N_14266);
xnor U14552 (N_14552,N_14387,N_14369);
nand U14553 (N_14553,N_14310,N_14378);
nor U14554 (N_14554,N_14213,N_14361);
or U14555 (N_14555,N_14323,N_14261);
nor U14556 (N_14556,N_14251,N_14360);
xnor U14557 (N_14557,N_14233,N_14239);
and U14558 (N_14558,N_14340,N_14279);
xor U14559 (N_14559,N_14395,N_14213);
xnor U14560 (N_14560,N_14277,N_14256);
and U14561 (N_14561,N_14282,N_14369);
nor U14562 (N_14562,N_14327,N_14328);
or U14563 (N_14563,N_14213,N_14353);
xnor U14564 (N_14564,N_14340,N_14315);
nor U14565 (N_14565,N_14223,N_14398);
and U14566 (N_14566,N_14339,N_14398);
xnor U14567 (N_14567,N_14351,N_14296);
or U14568 (N_14568,N_14251,N_14366);
or U14569 (N_14569,N_14257,N_14232);
or U14570 (N_14570,N_14270,N_14316);
and U14571 (N_14571,N_14306,N_14396);
or U14572 (N_14572,N_14234,N_14353);
and U14573 (N_14573,N_14203,N_14208);
and U14574 (N_14574,N_14348,N_14357);
or U14575 (N_14575,N_14228,N_14320);
and U14576 (N_14576,N_14277,N_14211);
or U14577 (N_14577,N_14379,N_14360);
nand U14578 (N_14578,N_14249,N_14279);
xnor U14579 (N_14579,N_14231,N_14267);
nor U14580 (N_14580,N_14315,N_14367);
and U14581 (N_14581,N_14390,N_14374);
xnor U14582 (N_14582,N_14352,N_14389);
or U14583 (N_14583,N_14396,N_14256);
or U14584 (N_14584,N_14373,N_14289);
or U14585 (N_14585,N_14291,N_14278);
or U14586 (N_14586,N_14249,N_14244);
nand U14587 (N_14587,N_14336,N_14292);
nand U14588 (N_14588,N_14232,N_14393);
xnor U14589 (N_14589,N_14383,N_14208);
nand U14590 (N_14590,N_14226,N_14397);
xor U14591 (N_14591,N_14290,N_14343);
nand U14592 (N_14592,N_14278,N_14372);
or U14593 (N_14593,N_14324,N_14205);
or U14594 (N_14594,N_14261,N_14276);
or U14595 (N_14595,N_14364,N_14275);
nand U14596 (N_14596,N_14387,N_14207);
and U14597 (N_14597,N_14385,N_14289);
or U14598 (N_14598,N_14323,N_14202);
and U14599 (N_14599,N_14272,N_14237);
xnor U14600 (N_14600,N_14426,N_14511);
xor U14601 (N_14601,N_14585,N_14575);
and U14602 (N_14602,N_14478,N_14464);
or U14603 (N_14603,N_14481,N_14566);
nor U14604 (N_14604,N_14451,N_14550);
nor U14605 (N_14605,N_14554,N_14433);
nor U14606 (N_14606,N_14423,N_14516);
nor U14607 (N_14607,N_14514,N_14567);
nand U14608 (N_14608,N_14509,N_14557);
and U14609 (N_14609,N_14402,N_14515);
xor U14610 (N_14610,N_14545,N_14519);
and U14611 (N_14611,N_14489,N_14421);
nor U14612 (N_14612,N_14496,N_14458);
nor U14613 (N_14613,N_14574,N_14487);
and U14614 (N_14614,N_14408,N_14562);
xor U14615 (N_14615,N_14595,N_14417);
nand U14616 (N_14616,N_14599,N_14494);
xor U14617 (N_14617,N_14459,N_14460);
or U14618 (N_14618,N_14527,N_14578);
xnor U14619 (N_14619,N_14500,N_14555);
and U14620 (N_14620,N_14541,N_14439);
xnor U14621 (N_14621,N_14449,N_14467);
nand U14622 (N_14622,N_14420,N_14530);
xnor U14623 (N_14623,N_14484,N_14534);
or U14624 (N_14624,N_14446,N_14539);
or U14625 (N_14625,N_14404,N_14597);
and U14626 (N_14626,N_14422,N_14559);
nor U14627 (N_14627,N_14431,N_14512);
or U14628 (N_14628,N_14589,N_14440);
and U14629 (N_14629,N_14490,N_14468);
or U14630 (N_14630,N_14533,N_14419);
nor U14631 (N_14631,N_14453,N_14418);
and U14632 (N_14632,N_14588,N_14565);
nand U14633 (N_14633,N_14401,N_14476);
and U14634 (N_14634,N_14450,N_14549);
nor U14635 (N_14635,N_14444,N_14522);
or U14636 (N_14636,N_14482,N_14445);
nor U14637 (N_14637,N_14488,N_14492);
and U14638 (N_14638,N_14593,N_14413);
and U14639 (N_14639,N_14412,N_14443);
or U14640 (N_14640,N_14579,N_14448);
and U14641 (N_14641,N_14465,N_14592);
xnor U14642 (N_14642,N_14480,N_14462);
and U14643 (N_14643,N_14581,N_14596);
and U14644 (N_14644,N_14583,N_14580);
xor U14645 (N_14645,N_14466,N_14531);
and U14646 (N_14646,N_14457,N_14523);
and U14647 (N_14647,N_14403,N_14456);
or U14648 (N_14648,N_14504,N_14517);
or U14649 (N_14649,N_14409,N_14493);
nor U14650 (N_14650,N_14598,N_14437);
and U14651 (N_14651,N_14473,N_14524);
nand U14652 (N_14652,N_14415,N_14501);
nor U14653 (N_14653,N_14560,N_14432);
or U14654 (N_14654,N_14442,N_14411);
xor U14655 (N_14655,N_14532,N_14498);
and U14656 (N_14656,N_14435,N_14590);
nand U14657 (N_14657,N_14556,N_14438);
nor U14658 (N_14658,N_14572,N_14552);
or U14659 (N_14659,N_14513,N_14571);
nor U14660 (N_14660,N_14591,N_14508);
xnor U14661 (N_14661,N_14528,N_14400);
xor U14662 (N_14662,N_14461,N_14452);
nor U14663 (N_14663,N_14497,N_14470);
xnor U14664 (N_14664,N_14469,N_14410);
xnor U14665 (N_14665,N_14455,N_14507);
and U14666 (N_14666,N_14548,N_14542);
or U14667 (N_14667,N_14485,N_14483);
or U14668 (N_14668,N_14474,N_14434);
xor U14669 (N_14669,N_14405,N_14547);
nand U14670 (N_14670,N_14594,N_14520);
nor U14671 (N_14671,N_14526,N_14553);
and U14672 (N_14672,N_14568,N_14586);
xnor U14673 (N_14673,N_14551,N_14577);
xor U14674 (N_14674,N_14538,N_14563);
nand U14675 (N_14675,N_14475,N_14576);
nor U14676 (N_14676,N_14441,N_14569);
and U14677 (N_14677,N_14428,N_14477);
nor U14678 (N_14678,N_14529,N_14510);
and U14679 (N_14679,N_14587,N_14570);
and U14680 (N_14680,N_14499,N_14424);
or U14681 (N_14681,N_14425,N_14430);
nand U14682 (N_14682,N_14502,N_14471);
xor U14683 (N_14683,N_14479,N_14561);
nor U14684 (N_14684,N_14414,N_14564);
and U14685 (N_14685,N_14427,N_14518);
or U14686 (N_14686,N_14536,N_14506);
nor U14687 (N_14687,N_14544,N_14486);
or U14688 (N_14688,N_14573,N_14429);
or U14689 (N_14689,N_14463,N_14540);
nand U14690 (N_14690,N_14454,N_14407);
and U14691 (N_14691,N_14525,N_14584);
nand U14692 (N_14692,N_14406,N_14495);
xor U14693 (N_14693,N_14472,N_14546);
nand U14694 (N_14694,N_14543,N_14503);
or U14695 (N_14695,N_14521,N_14582);
nand U14696 (N_14696,N_14535,N_14537);
xnor U14697 (N_14697,N_14436,N_14491);
and U14698 (N_14698,N_14558,N_14447);
xnor U14699 (N_14699,N_14505,N_14416);
xor U14700 (N_14700,N_14492,N_14473);
nor U14701 (N_14701,N_14505,N_14563);
and U14702 (N_14702,N_14545,N_14443);
and U14703 (N_14703,N_14508,N_14587);
or U14704 (N_14704,N_14509,N_14482);
nor U14705 (N_14705,N_14466,N_14439);
nor U14706 (N_14706,N_14494,N_14522);
and U14707 (N_14707,N_14503,N_14518);
and U14708 (N_14708,N_14409,N_14502);
xnor U14709 (N_14709,N_14517,N_14456);
nor U14710 (N_14710,N_14503,N_14429);
nor U14711 (N_14711,N_14551,N_14424);
or U14712 (N_14712,N_14461,N_14493);
or U14713 (N_14713,N_14452,N_14490);
nand U14714 (N_14714,N_14426,N_14580);
and U14715 (N_14715,N_14442,N_14434);
nor U14716 (N_14716,N_14515,N_14501);
nand U14717 (N_14717,N_14492,N_14480);
nand U14718 (N_14718,N_14503,N_14434);
xnor U14719 (N_14719,N_14561,N_14500);
or U14720 (N_14720,N_14484,N_14598);
nor U14721 (N_14721,N_14428,N_14526);
and U14722 (N_14722,N_14439,N_14409);
nor U14723 (N_14723,N_14505,N_14421);
xor U14724 (N_14724,N_14411,N_14477);
or U14725 (N_14725,N_14582,N_14434);
nor U14726 (N_14726,N_14492,N_14594);
xor U14727 (N_14727,N_14496,N_14554);
or U14728 (N_14728,N_14568,N_14442);
nor U14729 (N_14729,N_14470,N_14423);
and U14730 (N_14730,N_14448,N_14582);
nor U14731 (N_14731,N_14581,N_14448);
or U14732 (N_14732,N_14431,N_14591);
and U14733 (N_14733,N_14468,N_14478);
or U14734 (N_14734,N_14489,N_14415);
xnor U14735 (N_14735,N_14587,N_14543);
nor U14736 (N_14736,N_14554,N_14508);
nand U14737 (N_14737,N_14540,N_14588);
nor U14738 (N_14738,N_14571,N_14556);
xnor U14739 (N_14739,N_14535,N_14464);
and U14740 (N_14740,N_14502,N_14496);
or U14741 (N_14741,N_14458,N_14586);
and U14742 (N_14742,N_14444,N_14459);
nor U14743 (N_14743,N_14400,N_14571);
nor U14744 (N_14744,N_14493,N_14537);
or U14745 (N_14745,N_14462,N_14588);
or U14746 (N_14746,N_14516,N_14481);
nand U14747 (N_14747,N_14427,N_14481);
nor U14748 (N_14748,N_14473,N_14571);
xor U14749 (N_14749,N_14465,N_14572);
nor U14750 (N_14750,N_14552,N_14489);
and U14751 (N_14751,N_14467,N_14470);
and U14752 (N_14752,N_14580,N_14431);
nor U14753 (N_14753,N_14535,N_14586);
or U14754 (N_14754,N_14473,N_14547);
and U14755 (N_14755,N_14459,N_14474);
and U14756 (N_14756,N_14404,N_14491);
or U14757 (N_14757,N_14570,N_14496);
nand U14758 (N_14758,N_14537,N_14459);
or U14759 (N_14759,N_14583,N_14555);
nand U14760 (N_14760,N_14575,N_14445);
nor U14761 (N_14761,N_14401,N_14473);
nand U14762 (N_14762,N_14565,N_14507);
nand U14763 (N_14763,N_14443,N_14442);
or U14764 (N_14764,N_14493,N_14438);
and U14765 (N_14765,N_14427,N_14449);
and U14766 (N_14766,N_14527,N_14403);
xor U14767 (N_14767,N_14585,N_14449);
and U14768 (N_14768,N_14416,N_14421);
nand U14769 (N_14769,N_14427,N_14436);
xnor U14770 (N_14770,N_14503,N_14561);
or U14771 (N_14771,N_14459,N_14442);
or U14772 (N_14772,N_14445,N_14549);
or U14773 (N_14773,N_14407,N_14423);
nor U14774 (N_14774,N_14462,N_14553);
or U14775 (N_14775,N_14510,N_14492);
xnor U14776 (N_14776,N_14426,N_14460);
and U14777 (N_14777,N_14401,N_14582);
xnor U14778 (N_14778,N_14528,N_14437);
nor U14779 (N_14779,N_14553,N_14541);
or U14780 (N_14780,N_14557,N_14570);
nor U14781 (N_14781,N_14470,N_14474);
and U14782 (N_14782,N_14524,N_14582);
nand U14783 (N_14783,N_14422,N_14504);
nand U14784 (N_14784,N_14454,N_14518);
nand U14785 (N_14785,N_14430,N_14429);
and U14786 (N_14786,N_14404,N_14497);
or U14787 (N_14787,N_14415,N_14448);
xor U14788 (N_14788,N_14461,N_14581);
or U14789 (N_14789,N_14411,N_14456);
or U14790 (N_14790,N_14446,N_14409);
xnor U14791 (N_14791,N_14514,N_14444);
or U14792 (N_14792,N_14458,N_14539);
nand U14793 (N_14793,N_14577,N_14582);
xor U14794 (N_14794,N_14465,N_14599);
nor U14795 (N_14795,N_14448,N_14447);
and U14796 (N_14796,N_14416,N_14588);
xnor U14797 (N_14797,N_14573,N_14539);
and U14798 (N_14798,N_14463,N_14423);
or U14799 (N_14799,N_14539,N_14449);
or U14800 (N_14800,N_14635,N_14723);
and U14801 (N_14801,N_14659,N_14686);
and U14802 (N_14802,N_14794,N_14614);
and U14803 (N_14803,N_14766,N_14606);
xor U14804 (N_14804,N_14715,N_14797);
nor U14805 (N_14805,N_14758,N_14754);
nor U14806 (N_14806,N_14701,N_14664);
and U14807 (N_14807,N_14739,N_14662);
or U14808 (N_14808,N_14734,N_14781);
and U14809 (N_14809,N_14740,N_14655);
nand U14810 (N_14810,N_14728,N_14700);
and U14811 (N_14811,N_14705,N_14730);
or U14812 (N_14812,N_14769,N_14764);
and U14813 (N_14813,N_14663,N_14691);
nand U14814 (N_14814,N_14759,N_14735);
and U14815 (N_14815,N_14760,N_14631);
xor U14816 (N_14816,N_14775,N_14677);
nor U14817 (N_14817,N_14768,N_14637);
and U14818 (N_14818,N_14651,N_14668);
xnor U14819 (N_14819,N_14741,N_14776);
nor U14820 (N_14820,N_14656,N_14630);
nor U14821 (N_14821,N_14788,N_14678);
and U14822 (N_14822,N_14688,N_14761);
or U14823 (N_14823,N_14698,N_14608);
nand U14824 (N_14824,N_14763,N_14667);
or U14825 (N_14825,N_14699,N_14619);
and U14826 (N_14826,N_14719,N_14640);
nor U14827 (N_14827,N_14680,N_14658);
and U14828 (N_14828,N_14789,N_14687);
and U14829 (N_14829,N_14799,N_14648);
and U14830 (N_14830,N_14620,N_14634);
nand U14831 (N_14831,N_14646,N_14777);
or U14832 (N_14832,N_14750,N_14603);
xor U14833 (N_14833,N_14600,N_14676);
nand U14834 (N_14834,N_14612,N_14706);
nor U14835 (N_14835,N_14737,N_14792);
nor U14836 (N_14836,N_14743,N_14649);
nand U14837 (N_14837,N_14738,N_14736);
and U14838 (N_14838,N_14773,N_14616);
and U14839 (N_14839,N_14770,N_14650);
and U14840 (N_14840,N_14641,N_14704);
nand U14841 (N_14841,N_14628,N_14692);
and U14842 (N_14842,N_14765,N_14783);
nor U14843 (N_14843,N_14729,N_14710);
nor U14844 (N_14844,N_14786,N_14601);
nor U14845 (N_14845,N_14756,N_14689);
or U14846 (N_14846,N_14711,N_14731);
or U14847 (N_14847,N_14751,N_14696);
and U14848 (N_14848,N_14671,N_14717);
nor U14849 (N_14849,N_14609,N_14618);
xor U14850 (N_14850,N_14748,N_14657);
nand U14851 (N_14851,N_14654,N_14798);
xor U14852 (N_14852,N_14610,N_14685);
and U14853 (N_14853,N_14702,N_14774);
nor U14854 (N_14854,N_14666,N_14714);
or U14855 (N_14855,N_14690,N_14644);
nand U14856 (N_14856,N_14726,N_14716);
nor U14857 (N_14857,N_14779,N_14670);
nand U14858 (N_14858,N_14742,N_14626);
or U14859 (N_14859,N_14604,N_14707);
and U14860 (N_14860,N_14684,N_14643);
xnor U14861 (N_14861,N_14673,N_14694);
xnor U14862 (N_14862,N_14732,N_14745);
or U14863 (N_14863,N_14636,N_14629);
xor U14864 (N_14864,N_14669,N_14771);
or U14865 (N_14865,N_14725,N_14672);
nand U14866 (N_14866,N_14713,N_14793);
or U14867 (N_14867,N_14722,N_14703);
or U14868 (N_14868,N_14755,N_14660);
nand U14869 (N_14869,N_14780,N_14796);
nand U14870 (N_14870,N_14605,N_14682);
and U14871 (N_14871,N_14749,N_14791);
nand U14872 (N_14872,N_14645,N_14784);
or U14873 (N_14873,N_14639,N_14622);
or U14874 (N_14874,N_14661,N_14683);
nor U14875 (N_14875,N_14762,N_14615);
nand U14876 (N_14876,N_14625,N_14721);
nor U14877 (N_14877,N_14693,N_14744);
and U14878 (N_14878,N_14785,N_14733);
or U14879 (N_14879,N_14647,N_14632);
xor U14880 (N_14880,N_14697,N_14679);
xor U14881 (N_14881,N_14633,N_14790);
and U14882 (N_14882,N_14767,N_14757);
nor U14883 (N_14883,N_14627,N_14624);
or U14884 (N_14884,N_14665,N_14746);
or U14885 (N_14885,N_14652,N_14753);
or U14886 (N_14886,N_14752,N_14607);
xnor U14887 (N_14887,N_14675,N_14720);
and U14888 (N_14888,N_14617,N_14724);
or U14889 (N_14889,N_14642,N_14795);
xor U14890 (N_14890,N_14602,N_14653);
nor U14891 (N_14891,N_14611,N_14695);
and U14892 (N_14892,N_14709,N_14621);
and U14893 (N_14893,N_14623,N_14772);
and U14894 (N_14894,N_14747,N_14782);
nor U14895 (N_14895,N_14778,N_14712);
xor U14896 (N_14896,N_14638,N_14708);
nand U14897 (N_14897,N_14674,N_14613);
and U14898 (N_14898,N_14727,N_14681);
or U14899 (N_14899,N_14718,N_14787);
or U14900 (N_14900,N_14751,N_14727);
nand U14901 (N_14901,N_14702,N_14786);
nor U14902 (N_14902,N_14671,N_14672);
xnor U14903 (N_14903,N_14634,N_14746);
and U14904 (N_14904,N_14765,N_14623);
nor U14905 (N_14905,N_14758,N_14780);
nor U14906 (N_14906,N_14774,N_14734);
xnor U14907 (N_14907,N_14709,N_14689);
nor U14908 (N_14908,N_14743,N_14715);
nand U14909 (N_14909,N_14670,N_14646);
or U14910 (N_14910,N_14739,N_14710);
nand U14911 (N_14911,N_14685,N_14696);
xnor U14912 (N_14912,N_14762,N_14782);
nand U14913 (N_14913,N_14602,N_14771);
and U14914 (N_14914,N_14723,N_14738);
or U14915 (N_14915,N_14616,N_14769);
nand U14916 (N_14916,N_14723,N_14733);
nand U14917 (N_14917,N_14787,N_14700);
xnor U14918 (N_14918,N_14647,N_14710);
or U14919 (N_14919,N_14622,N_14646);
nor U14920 (N_14920,N_14627,N_14745);
or U14921 (N_14921,N_14670,N_14626);
xor U14922 (N_14922,N_14755,N_14647);
nand U14923 (N_14923,N_14601,N_14673);
nand U14924 (N_14924,N_14731,N_14719);
and U14925 (N_14925,N_14651,N_14709);
and U14926 (N_14926,N_14721,N_14614);
nor U14927 (N_14927,N_14609,N_14737);
nor U14928 (N_14928,N_14646,N_14613);
or U14929 (N_14929,N_14734,N_14605);
xor U14930 (N_14930,N_14743,N_14767);
xnor U14931 (N_14931,N_14706,N_14641);
nand U14932 (N_14932,N_14789,N_14622);
nor U14933 (N_14933,N_14729,N_14725);
xor U14934 (N_14934,N_14628,N_14640);
and U14935 (N_14935,N_14659,N_14799);
xor U14936 (N_14936,N_14698,N_14799);
xnor U14937 (N_14937,N_14719,N_14603);
nor U14938 (N_14938,N_14635,N_14609);
and U14939 (N_14939,N_14720,N_14648);
xnor U14940 (N_14940,N_14708,N_14691);
and U14941 (N_14941,N_14649,N_14727);
nand U14942 (N_14942,N_14759,N_14683);
and U14943 (N_14943,N_14663,N_14701);
or U14944 (N_14944,N_14777,N_14735);
nand U14945 (N_14945,N_14667,N_14781);
nand U14946 (N_14946,N_14718,N_14703);
nor U14947 (N_14947,N_14616,N_14727);
or U14948 (N_14948,N_14674,N_14669);
xnor U14949 (N_14949,N_14657,N_14751);
nand U14950 (N_14950,N_14711,N_14766);
or U14951 (N_14951,N_14685,N_14664);
and U14952 (N_14952,N_14799,N_14623);
xor U14953 (N_14953,N_14715,N_14649);
xor U14954 (N_14954,N_14674,N_14786);
nand U14955 (N_14955,N_14701,N_14798);
nand U14956 (N_14956,N_14621,N_14730);
xor U14957 (N_14957,N_14675,N_14702);
xnor U14958 (N_14958,N_14781,N_14755);
xnor U14959 (N_14959,N_14729,N_14683);
and U14960 (N_14960,N_14615,N_14683);
and U14961 (N_14961,N_14606,N_14698);
or U14962 (N_14962,N_14699,N_14693);
nand U14963 (N_14963,N_14757,N_14789);
nor U14964 (N_14964,N_14787,N_14606);
nor U14965 (N_14965,N_14724,N_14666);
xnor U14966 (N_14966,N_14709,N_14631);
xor U14967 (N_14967,N_14677,N_14671);
nand U14968 (N_14968,N_14743,N_14728);
nand U14969 (N_14969,N_14786,N_14730);
nand U14970 (N_14970,N_14756,N_14732);
nand U14971 (N_14971,N_14604,N_14716);
or U14972 (N_14972,N_14764,N_14786);
nor U14973 (N_14973,N_14704,N_14723);
or U14974 (N_14974,N_14775,N_14687);
xor U14975 (N_14975,N_14683,N_14655);
xnor U14976 (N_14976,N_14656,N_14633);
xor U14977 (N_14977,N_14702,N_14744);
or U14978 (N_14978,N_14609,N_14745);
xor U14979 (N_14979,N_14731,N_14734);
nor U14980 (N_14980,N_14676,N_14765);
nor U14981 (N_14981,N_14719,N_14725);
and U14982 (N_14982,N_14719,N_14680);
or U14983 (N_14983,N_14767,N_14626);
nand U14984 (N_14984,N_14626,N_14719);
xnor U14985 (N_14985,N_14706,N_14635);
xnor U14986 (N_14986,N_14781,N_14646);
or U14987 (N_14987,N_14794,N_14685);
and U14988 (N_14988,N_14761,N_14729);
nor U14989 (N_14989,N_14626,N_14672);
nand U14990 (N_14990,N_14668,N_14680);
nand U14991 (N_14991,N_14644,N_14630);
and U14992 (N_14992,N_14667,N_14725);
xor U14993 (N_14993,N_14620,N_14676);
xor U14994 (N_14994,N_14765,N_14678);
xnor U14995 (N_14995,N_14659,N_14625);
xor U14996 (N_14996,N_14700,N_14679);
or U14997 (N_14997,N_14665,N_14797);
nand U14998 (N_14998,N_14654,N_14731);
or U14999 (N_14999,N_14668,N_14770);
and UO_0 (O_0,N_14862,N_14922);
or UO_1 (O_1,N_14964,N_14874);
nand UO_2 (O_2,N_14974,N_14944);
and UO_3 (O_3,N_14811,N_14971);
and UO_4 (O_4,N_14838,N_14917);
xor UO_5 (O_5,N_14826,N_14854);
nand UO_6 (O_6,N_14904,N_14932);
nand UO_7 (O_7,N_14924,N_14941);
nand UO_8 (O_8,N_14880,N_14873);
nor UO_9 (O_9,N_14882,N_14956);
nor UO_10 (O_10,N_14966,N_14951);
nand UO_11 (O_11,N_14913,N_14995);
nand UO_12 (O_12,N_14909,N_14803);
and UO_13 (O_13,N_14939,N_14822);
nand UO_14 (O_14,N_14918,N_14884);
xnor UO_15 (O_15,N_14858,N_14827);
and UO_16 (O_16,N_14887,N_14997);
nand UO_17 (O_17,N_14875,N_14921);
xor UO_18 (O_18,N_14849,N_14891);
nor UO_19 (O_19,N_14804,N_14871);
nor UO_20 (O_20,N_14840,N_14863);
or UO_21 (O_21,N_14890,N_14970);
xor UO_22 (O_22,N_14923,N_14812);
or UO_23 (O_23,N_14865,N_14846);
or UO_24 (O_24,N_14876,N_14906);
or UO_25 (O_25,N_14843,N_14911);
xor UO_26 (O_26,N_14817,N_14965);
and UO_27 (O_27,N_14929,N_14809);
nor UO_28 (O_28,N_14950,N_14893);
nor UO_29 (O_29,N_14936,N_14926);
or UO_30 (O_30,N_14975,N_14988);
or UO_31 (O_31,N_14859,N_14930);
nand UO_32 (O_32,N_14973,N_14832);
or UO_33 (O_33,N_14872,N_14903);
and UO_34 (O_34,N_14928,N_14842);
and UO_35 (O_35,N_14902,N_14994);
nand UO_36 (O_36,N_14894,N_14801);
xnor UO_37 (O_37,N_14955,N_14855);
xor UO_38 (O_38,N_14828,N_14853);
nor UO_39 (O_39,N_14807,N_14948);
nor UO_40 (O_40,N_14881,N_14883);
or UO_41 (O_41,N_14987,N_14866);
or UO_42 (O_42,N_14857,N_14996);
nand UO_43 (O_43,N_14877,N_14969);
nor UO_44 (O_44,N_14813,N_14805);
nand UO_45 (O_45,N_14919,N_14823);
or UO_46 (O_46,N_14868,N_14999);
nor UO_47 (O_47,N_14914,N_14824);
nand UO_48 (O_48,N_14934,N_14885);
or UO_49 (O_49,N_14931,N_14816);
xor UO_50 (O_50,N_14980,N_14852);
or UO_51 (O_51,N_14830,N_14986);
or UO_52 (O_52,N_14952,N_14864);
xnor UO_53 (O_53,N_14897,N_14837);
nand UO_54 (O_54,N_14833,N_14836);
xor UO_55 (O_55,N_14869,N_14947);
nor UO_56 (O_56,N_14898,N_14963);
xnor UO_57 (O_57,N_14960,N_14810);
and UO_58 (O_58,N_14856,N_14938);
or UO_59 (O_59,N_14845,N_14886);
nor UO_60 (O_60,N_14896,N_14900);
nor UO_61 (O_61,N_14982,N_14920);
nor UO_62 (O_62,N_14962,N_14984);
xnor UO_63 (O_63,N_14895,N_14957);
nor UO_64 (O_64,N_14925,N_14989);
or UO_65 (O_65,N_14814,N_14972);
or UO_66 (O_66,N_14977,N_14953);
and UO_67 (O_67,N_14933,N_14800);
nand UO_68 (O_68,N_14968,N_14927);
and UO_69 (O_69,N_14889,N_14907);
and UO_70 (O_70,N_14818,N_14831);
nand UO_71 (O_71,N_14878,N_14888);
nor UO_72 (O_72,N_14958,N_14981);
nand UO_73 (O_73,N_14835,N_14867);
and UO_74 (O_74,N_14820,N_14979);
and UO_75 (O_75,N_14916,N_14829);
nand UO_76 (O_76,N_14954,N_14841);
nand UO_77 (O_77,N_14976,N_14912);
nor UO_78 (O_78,N_14990,N_14991);
or UO_79 (O_79,N_14808,N_14992);
nand UO_80 (O_80,N_14839,N_14993);
or UO_81 (O_81,N_14985,N_14848);
xnor UO_82 (O_82,N_14943,N_14870);
xor UO_83 (O_83,N_14940,N_14847);
or UO_84 (O_84,N_14915,N_14942);
or UO_85 (O_85,N_14959,N_14910);
and UO_86 (O_86,N_14851,N_14945);
and UO_87 (O_87,N_14905,N_14983);
and UO_88 (O_88,N_14844,N_14899);
xnor UO_89 (O_89,N_14850,N_14815);
xor UO_90 (O_90,N_14825,N_14937);
or UO_91 (O_91,N_14819,N_14834);
xnor UO_92 (O_92,N_14935,N_14892);
or UO_93 (O_93,N_14998,N_14901);
nor UO_94 (O_94,N_14879,N_14961);
and UO_95 (O_95,N_14860,N_14978);
nor UO_96 (O_96,N_14802,N_14908);
and UO_97 (O_97,N_14946,N_14861);
xor UO_98 (O_98,N_14806,N_14967);
nor UO_99 (O_99,N_14949,N_14821);
or UO_100 (O_100,N_14927,N_14918);
nand UO_101 (O_101,N_14952,N_14852);
nor UO_102 (O_102,N_14947,N_14835);
nor UO_103 (O_103,N_14986,N_14835);
nor UO_104 (O_104,N_14919,N_14963);
nor UO_105 (O_105,N_14993,N_14849);
nor UO_106 (O_106,N_14842,N_14940);
and UO_107 (O_107,N_14922,N_14880);
and UO_108 (O_108,N_14892,N_14992);
xnor UO_109 (O_109,N_14986,N_14870);
or UO_110 (O_110,N_14855,N_14995);
nand UO_111 (O_111,N_14970,N_14877);
xnor UO_112 (O_112,N_14980,N_14837);
xnor UO_113 (O_113,N_14845,N_14839);
xnor UO_114 (O_114,N_14933,N_14816);
xnor UO_115 (O_115,N_14813,N_14851);
and UO_116 (O_116,N_14860,N_14940);
or UO_117 (O_117,N_14977,N_14878);
and UO_118 (O_118,N_14835,N_14937);
or UO_119 (O_119,N_14955,N_14981);
and UO_120 (O_120,N_14965,N_14960);
and UO_121 (O_121,N_14965,N_14959);
xor UO_122 (O_122,N_14975,N_14937);
nand UO_123 (O_123,N_14926,N_14903);
or UO_124 (O_124,N_14888,N_14866);
or UO_125 (O_125,N_14856,N_14829);
nand UO_126 (O_126,N_14939,N_14885);
and UO_127 (O_127,N_14845,N_14928);
and UO_128 (O_128,N_14993,N_14866);
and UO_129 (O_129,N_14902,N_14990);
xor UO_130 (O_130,N_14969,N_14875);
nor UO_131 (O_131,N_14964,N_14872);
xor UO_132 (O_132,N_14943,N_14906);
nor UO_133 (O_133,N_14891,N_14842);
xnor UO_134 (O_134,N_14805,N_14946);
nor UO_135 (O_135,N_14857,N_14960);
and UO_136 (O_136,N_14873,N_14932);
nand UO_137 (O_137,N_14928,N_14926);
nand UO_138 (O_138,N_14925,N_14854);
and UO_139 (O_139,N_14842,N_14800);
nor UO_140 (O_140,N_14951,N_14932);
or UO_141 (O_141,N_14956,N_14877);
nor UO_142 (O_142,N_14891,N_14988);
xnor UO_143 (O_143,N_14899,N_14873);
or UO_144 (O_144,N_14991,N_14856);
and UO_145 (O_145,N_14883,N_14911);
nand UO_146 (O_146,N_14827,N_14958);
nor UO_147 (O_147,N_14874,N_14834);
xnor UO_148 (O_148,N_14912,N_14966);
or UO_149 (O_149,N_14809,N_14873);
nor UO_150 (O_150,N_14967,N_14846);
nand UO_151 (O_151,N_14929,N_14965);
or UO_152 (O_152,N_14832,N_14916);
nand UO_153 (O_153,N_14926,N_14834);
nand UO_154 (O_154,N_14834,N_14984);
and UO_155 (O_155,N_14840,N_14930);
or UO_156 (O_156,N_14909,N_14889);
xnor UO_157 (O_157,N_14909,N_14899);
or UO_158 (O_158,N_14996,N_14885);
xor UO_159 (O_159,N_14881,N_14813);
and UO_160 (O_160,N_14843,N_14866);
xnor UO_161 (O_161,N_14826,N_14989);
xor UO_162 (O_162,N_14823,N_14942);
nor UO_163 (O_163,N_14847,N_14918);
nand UO_164 (O_164,N_14905,N_14990);
nand UO_165 (O_165,N_14870,N_14834);
nor UO_166 (O_166,N_14956,N_14836);
or UO_167 (O_167,N_14994,N_14895);
xnor UO_168 (O_168,N_14967,N_14982);
and UO_169 (O_169,N_14973,N_14842);
or UO_170 (O_170,N_14906,N_14814);
nand UO_171 (O_171,N_14828,N_14903);
nor UO_172 (O_172,N_14936,N_14800);
and UO_173 (O_173,N_14936,N_14854);
nor UO_174 (O_174,N_14860,N_14851);
nor UO_175 (O_175,N_14811,N_14934);
nor UO_176 (O_176,N_14867,N_14956);
and UO_177 (O_177,N_14912,N_14884);
nand UO_178 (O_178,N_14829,N_14847);
nand UO_179 (O_179,N_14906,N_14850);
xor UO_180 (O_180,N_14844,N_14876);
nor UO_181 (O_181,N_14905,N_14919);
and UO_182 (O_182,N_14995,N_14836);
and UO_183 (O_183,N_14975,N_14990);
xor UO_184 (O_184,N_14804,N_14915);
xnor UO_185 (O_185,N_14843,N_14863);
xor UO_186 (O_186,N_14910,N_14898);
xnor UO_187 (O_187,N_14882,N_14800);
xor UO_188 (O_188,N_14865,N_14931);
nor UO_189 (O_189,N_14996,N_14901);
or UO_190 (O_190,N_14848,N_14952);
xnor UO_191 (O_191,N_14888,N_14967);
xnor UO_192 (O_192,N_14999,N_14852);
and UO_193 (O_193,N_14923,N_14818);
nand UO_194 (O_194,N_14946,N_14865);
or UO_195 (O_195,N_14902,N_14934);
and UO_196 (O_196,N_14943,N_14845);
or UO_197 (O_197,N_14858,N_14863);
and UO_198 (O_198,N_14900,N_14878);
nand UO_199 (O_199,N_14956,N_14805);
xor UO_200 (O_200,N_14803,N_14974);
nand UO_201 (O_201,N_14818,N_14904);
xor UO_202 (O_202,N_14804,N_14813);
nor UO_203 (O_203,N_14905,N_14883);
xnor UO_204 (O_204,N_14958,N_14934);
or UO_205 (O_205,N_14993,N_14970);
nand UO_206 (O_206,N_14878,N_14853);
and UO_207 (O_207,N_14870,N_14902);
and UO_208 (O_208,N_14859,N_14951);
or UO_209 (O_209,N_14885,N_14831);
xor UO_210 (O_210,N_14845,N_14851);
and UO_211 (O_211,N_14801,N_14870);
nand UO_212 (O_212,N_14879,N_14905);
or UO_213 (O_213,N_14817,N_14824);
xnor UO_214 (O_214,N_14888,N_14840);
and UO_215 (O_215,N_14915,N_14934);
nor UO_216 (O_216,N_14867,N_14862);
nand UO_217 (O_217,N_14932,N_14943);
or UO_218 (O_218,N_14987,N_14961);
xnor UO_219 (O_219,N_14850,N_14814);
nand UO_220 (O_220,N_14961,N_14868);
nor UO_221 (O_221,N_14880,N_14924);
and UO_222 (O_222,N_14925,N_14907);
nor UO_223 (O_223,N_14857,N_14904);
nand UO_224 (O_224,N_14918,N_14839);
nand UO_225 (O_225,N_14927,N_14920);
nand UO_226 (O_226,N_14824,N_14959);
and UO_227 (O_227,N_14946,N_14991);
xnor UO_228 (O_228,N_14990,N_14970);
xor UO_229 (O_229,N_14915,N_14925);
and UO_230 (O_230,N_14879,N_14820);
nor UO_231 (O_231,N_14829,N_14923);
nor UO_232 (O_232,N_14996,N_14916);
xor UO_233 (O_233,N_14962,N_14870);
or UO_234 (O_234,N_14845,N_14808);
or UO_235 (O_235,N_14826,N_14945);
nand UO_236 (O_236,N_14869,N_14973);
xnor UO_237 (O_237,N_14915,N_14974);
and UO_238 (O_238,N_14843,N_14939);
nor UO_239 (O_239,N_14978,N_14904);
xor UO_240 (O_240,N_14924,N_14931);
and UO_241 (O_241,N_14937,N_14883);
or UO_242 (O_242,N_14913,N_14986);
xnor UO_243 (O_243,N_14874,N_14990);
nor UO_244 (O_244,N_14954,N_14940);
and UO_245 (O_245,N_14898,N_14808);
nand UO_246 (O_246,N_14858,N_14950);
or UO_247 (O_247,N_14898,N_14863);
xnor UO_248 (O_248,N_14874,N_14974);
and UO_249 (O_249,N_14813,N_14848);
nor UO_250 (O_250,N_14904,N_14862);
and UO_251 (O_251,N_14915,N_14865);
or UO_252 (O_252,N_14816,N_14889);
and UO_253 (O_253,N_14850,N_14833);
nand UO_254 (O_254,N_14806,N_14807);
xnor UO_255 (O_255,N_14828,N_14819);
nand UO_256 (O_256,N_14987,N_14806);
xor UO_257 (O_257,N_14820,N_14891);
nor UO_258 (O_258,N_14823,N_14868);
or UO_259 (O_259,N_14972,N_14966);
nand UO_260 (O_260,N_14981,N_14970);
nor UO_261 (O_261,N_14987,N_14883);
or UO_262 (O_262,N_14903,N_14982);
or UO_263 (O_263,N_14879,N_14933);
nor UO_264 (O_264,N_14910,N_14951);
nor UO_265 (O_265,N_14823,N_14907);
nand UO_266 (O_266,N_14990,N_14886);
and UO_267 (O_267,N_14804,N_14818);
or UO_268 (O_268,N_14933,N_14825);
xnor UO_269 (O_269,N_14957,N_14821);
nand UO_270 (O_270,N_14963,N_14987);
nand UO_271 (O_271,N_14893,N_14866);
xor UO_272 (O_272,N_14994,N_14966);
xor UO_273 (O_273,N_14916,N_14991);
and UO_274 (O_274,N_14960,N_14992);
or UO_275 (O_275,N_14962,N_14930);
nor UO_276 (O_276,N_14852,N_14833);
nand UO_277 (O_277,N_14981,N_14865);
and UO_278 (O_278,N_14995,N_14877);
and UO_279 (O_279,N_14844,N_14963);
xnor UO_280 (O_280,N_14844,N_14912);
or UO_281 (O_281,N_14851,N_14999);
nand UO_282 (O_282,N_14846,N_14863);
nor UO_283 (O_283,N_14966,N_14883);
xnor UO_284 (O_284,N_14933,N_14928);
nor UO_285 (O_285,N_14878,N_14834);
or UO_286 (O_286,N_14974,N_14970);
and UO_287 (O_287,N_14989,N_14993);
and UO_288 (O_288,N_14807,N_14856);
nand UO_289 (O_289,N_14801,N_14948);
nor UO_290 (O_290,N_14998,N_14875);
xnor UO_291 (O_291,N_14987,N_14895);
nand UO_292 (O_292,N_14990,N_14920);
nand UO_293 (O_293,N_14847,N_14969);
xor UO_294 (O_294,N_14931,N_14948);
nand UO_295 (O_295,N_14810,N_14812);
xor UO_296 (O_296,N_14939,N_14944);
nand UO_297 (O_297,N_14903,N_14824);
or UO_298 (O_298,N_14930,N_14807);
nand UO_299 (O_299,N_14945,N_14871);
xnor UO_300 (O_300,N_14961,N_14948);
or UO_301 (O_301,N_14888,N_14863);
or UO_302 (O_302,N_14964,N_14891);
nand UO_303 (O_303,N_14941,N_14986);
nor UO_304 (O_304,N_14850,N_14855);
or UO_305 (O_305,N_14860,N_14837);
nor UO_306 (O_306,N_14872,N_14868);
xor UO_307 (O_307,N_14963,N_14918);
nand UO_308 (O_308,N_14907,N_14953);
or UO_309 (O_309,N_14945,N_14901);
xnor UO_310 (O_310,N_14856,N_14839);
nor UO_311 (O_311,N_14984,N_14996);
xor UO_312 (O_312,N_14848,N_14824);
nand UO_313 (O_313,N_14834,N_14817);
and UO_314 (O_314,N_14972,N_14815);
and UO_315 (O_315,N_14809,N_14968);
or UO_316 (O_316,N_14964,N_14867);
nand UO_317 (O_317,N_14891,N_14889);
nor UO_318 (O_318,N_14909,N_14865);
xnor UO_319 (O_319,N_14804,N_14957);
and UO_320 (O_320,N_14855,N_14992);
nand UO_321 (O_321,N_14950,N_14920);
xnor UO_322 (O_322,N_14828,N_14944);
nand UO_323 (O_323,N_14819,N_14919);
and UO_324 (O_324,N_14982,N_14892);
or UO_325 (O_325,N_14858,N_14961);
and UO_326 (O_326,N_14926,N_14959);
xor UO_327 (O_327,N_14876,N_14917);
or UO_328 (O_328,N_14952,N_14851);
nor UO_329 (O_329,N_14922,N_14800);
nand UO_330 (O_330,N_14883,N_14826);
or UO_331 (O_331,N_14926,N_14814);
nor UO_332 (O_332,N_14844,N_14823);
nor UO_333 (O_333,N_14902,N_14961);
nand UO_334 (O_334,N_14836,N_14823);
nand UO_335 (O_335,N_14958,N_14884);
nor UO_336 (O_336,N_14937,N_14946);
nand UO_337 (O_337,N_14951,N_14914);
nor UO_338 (O_338,N_14891,N_14934);
nand UO_339 (O_339,N_14946,N_14878);
nand UO_340 (O_340,N_14933,N_14896);
nor UO_341 (O_341,N_14848,N_14838);
nand UO_342 (O_342,N_14843,N_14822);
and UO_343 (O_343,N_14979,N_14987);
nor UO_344 (O_344,N_14906,N_14898);
and UO_345 (O_345,N_14991,N_14825);
and UO_346 (O_346,N_14999,N_14830);
or UO_347 (O_347,N_14889,N_14823);
nand UO_348 (O_348,N_14851,N_14850);
nand UO_349 (O_349,N_14916,N_14843);
or UO_350 (O_350,N_14887,N_14954);
nand UO_351 (O_351,N_14992,N_14984);
and UO_352 (O_352,N_14918,N_14897);
or UO_353 (O_353,N_14824,N_14909);
nand UO_354 (O_354,N_14908,N_14927);
nor UO_355 (O_355,N_14990,N_14844);
nand UO_356 (O_356,N_14989,N_14918);
xor UO_357 (O_357,N_14809,N_14944);
or UO_358 (O_358,N_14941,N_14847);
nand UO_359 (O_359,N_14929,N_14851);
nand UO_360 (O_360,N_14973,N_14935);
nor UO_361 (O_361,N_14854,N_14827);
nand UO_362 (O_362,N_14997,N_14842);
nand UO_363 (O_363,N_14989,N_14953);
or UO_364 (O_364,N_14883,N_14944);
nand UO_365 (O_365,N_14985,N_14895);
nor UO_366 (O_366,N_14829,N_14867);
and UO_367 (O_367,N_14841,N_14816);
nand UO_368 (O_368,N_14949,N_14935);
xnor UO_369 (O_369,N_14979,N_14800);
or UO_370 (O_370,N_14820,N_14807);
xor UO_371 (O_371,N_14911,N_14831);
xnor UO_372 (O_372,N_14943,N_14914);
xnor UO_373 (O_373,N_14932,N_14890);
or UO_374 (O_374,N_14938,N_14903);
nand UO_375 (O_375,N_14811,N_14821);
nand UO_376 (O_376,N_14839,N_14800);
and UO_377 (O_377,N_14941,N_14926);
and UO_378 (O_378,N_14809,N_14941);
xnor UO_379 (O_379,N_14869,N_14868);
and UO_380 (O_380,N_14916,N_14949);
nand UO_381 (O_381,N_14851,N_14859);
nand UO_382 (O_382,N_14913,N_14822);
or UO_383 (O_383,N_14814,N_14981);
or UO_384 (O_384,N_14994,N_14886);
nand UO_385 (O_385,N_14908,N_14895);
and UO_386 (O_386,N_14956,N_14860);
nand UO_387 (O_387,N_14884,N_14849);
xnor UO_388 (O_388,N_14800,N_14923);
or UO_389 (O_389,N_14959,N_14881);
nand UO_390 (O_390,N_14826,N_14872);
and UO_391 (O_391,N_14928,N_14932);
and UO_392 (O_392,N_14884,N_14882);
or UO_393 (O_393,N_14864,N_14927);
nand UO_394 (O_394,N_14849,N_14932);
nor UO_395 (O_395,N_14972,N_14818);
or UO_396 (O_396,N_14911,N_14866);
and UO_397 (O_397,N_14996,N_14838);
or UO_398 (O_398,N_14921,N_14978);
or UO_399 (O_399,N_14837,N_14859);
nor UO_400 (O_400,N_14863,N_14934);
nor UO_401 (O_401,N_14998,N_14832);
and UO_402 (O_402,N_14942,N_14844);
or UO_403 (O_403,N_14945,N_14859);
nor UO_404 (O_404,N_14872,N_14835);
xnor UO_405 (O_405,N_14831,N_14907);
nand UO_406 (O_406,N_14973,N_14910);
and UO_407 (O_407,N_14869,N_14833);
or UO_408 (O_408,N_14884,N_14890);
xor UO_409 (O_409,N_14948,N_14873);
nand UO_410 (O_410,N_14890,N_14871);
xnor UO_411 (O_411,N_14925,N_14922);
xor UO_412 (O_412,N_14812,N_14900);
nor UO_413 (O_413,N_14860,N_14941);
or UO_414 (O_414,N_14959,N_14999);
nand UO_415 (O_415,N_14844,N_14868);
nand UO_416 (O_416,N_14866,N_14991);
xnor UO_417 (O_417,N_14976,N_14823);
and UO_418 (O_418,N_14945,N_14908);
xor UO_419 (O_419,N_14829,N_14910);
nor UO_420 (O_420,N_14985,N_14839);
nand UO_421 (O_421,N_14864,N_14800);
nand UO_422 (O_422,N_14872,N_14960);
nor UO_423 (O_423,N_14922,N_14807);
or UO_424 (O_424,N_14976,N_14937);
xor UO_425 (O_425,N_14820,N_14856);
xnor UO_426 (O_426,N_14806,N_14949);
nor UO_427 (O_427,N_14939,N_14880);
or UO_428 (O_428,N_14852,N_14808);
and UO_429 (O_429,N_14973,N_14820);
nor UO_430 (O_430,N_14976,N_14894);
or UO_431 (O_431,N_14976,N_14842);
xnor UO_432 (O_432,N_14862,N_14947);
nand UO_433 (O_433,N_14984,N_14994);
nor UO_434 (O_434,N_14934,N_14824);
nand UO_435 (O_435,N_14890,N_14997);
xnor UO_436 (O_436,N_14810,N_14805);
and UO_437 (O_437,N_14950,N_14998);
nand UO_438 (O_438,N_14924,N_14953);
xor UO_439 (O_439,N_14868,N_14927);
and UO_440 (O_440,N_14824,N_14805);
xnor UO_441 (O_441,N_14964,N_14857);
or UO_442 (O_442,N_14846,N_14853);
nand UO_443 (O_443,N_14897,N_14861);
and UO_444 (O_444,N_14874,N_14879);
nand UO_445 (O_445,N_14944,N_14872);
nor UO_446 (O_446,N_14843,N_14997);
nand UO_447 (O_447,N_14865,N_14918);
and UO_448 (O_448,N_14819,N_14939);
or UO_449 (O_449,N_14996,N_14918);
nor UO_450 (O_450,N_14949,N_14957);
xor UO_451 (O_451,N_14889,N_14810);
and UO_452 (O_452,N_14971,N_14849);
xor UO_453 (O_453,N_14888,N_14852);
or UO_454 (O_454,N_14979,N_14830);
or UO_455 (O_455,N_14818,N_14925);
and UO_456 (O_456,N_14970,N_14953);
xor UO_457 (O_457,N_14978,N_14891);
or UO_458 (O_458,N_14875,N_14851);
nor UO_459 (O_459,N_14903,N_14998);
nor UO_460 (O_460,N_14976,N_14857);
and UO_461 (O_461,N_14885,N_14946);
nor UO_462 (O_462,N_14966,N_14886);
and UO_463 (O_463,N_14922,N_14883);
or UO_464 (O_464,N_14967,N_14957);
nor UO_465 (O_465,N_14809,N_14811);
nor UO_466 (O_466,N_14967,N_14917);
or UO_467 (O_467,N_14933,N_14876);
nor UO_468 (O_468,N_14982,N_14895);
nand UO_469 (O_469,N_14833,N_14870);
and UO_470 (O_470,N_14975,N_14978);
and UO_471 (O_471,N_14860,N_14821);
xor UO_472 (O_472,N_14838,N_14958);
nand UO_473 (O_473,N_14855,N_14802);
or UO_474 (O_474,N_14889,N_14842);
and UO_475 (O_475,N_14899,N_14883);
nor UO_476 (O_476,N_14958,N_14945);
or UO_477 (O_477,N_14819,N_14835);
nand UO_478 (O_478,N_14970,N_14954);
nor UO_479 (O_479,N_14904,N_14916);
xnor UO_480 (O_480,N_14964,N_14979);
xor UO_481 (O_481,N_14931,N_14845);
nand UO_482 (O_482,N_14886,N_14913);
or UO_483 (O_483,N_14974,N_14854);
or UO_484 (O_484,N_14985,N_14811);
nand UO_485 (O_485,N_14972,N_14849);
xnor UO_486 (O_486,N_14878,N_14845);
or UO_487 (O_487,N_14872,N_14811);
nor UO_488 (O_488,N_14894,N_14887);
and UO_489 (O_489,N_14978,N_14977);
xor UO_490 (O_490,N_14868,N_14871);
nand UO_491 (O_491,N_14996,N_14886);
nor UO_492 (O_492,N_14808,N_14871);
xnor UO_493 (O_493,N_14861,N_14848);
and UO_494 (O_494,N_14842,N_14902);
nor UO_495 (O_495,N_14813,N_14866);
or UO_496 (O_496,N_14933,N_14969);
or UO_497 (O_497,N_14869,N_14801);
or UO_498 (O_498,N_14829,N_14933);
nand UO_499 (O_499,N_14987,N_14965);
nand UO_500 (O_500,N_14827,N_14955);
xnor UO_501 (O_501,N_14907,N_14863);
nor UO_502 (O_502,N_14956,N_14871);
nand UO_503 (O_503,N_14888,N_14907);
nand UO_504 (O_504,N_14891,N_14864);
or UO_505 (O_505,N_14813,N_14849);
or UO_506 (O_506,N_14829,N_14969);
or UO_507 (O_507,N_14984,N_14885);
and UO_508 (O_508,N_14814,N_14812);
or UO_509 (O_509,N_14951,N_14890);
or UO_510 (O_510,N_14964,N_14920);
and UO_511 (O_511,N_14952,N_14986);
or UO_512 (O_512,N_14943,N_14915);
xor UO_513 (O_513,N_14816,N_14838);
nand UO_514 (O_514,N_14822,N_14842);
nor UO_515 (O_515,N_14974,N_14941);
xnor UO_516 (O_516,N_14977,N_14962);
nor UO_517 (O_517,N_14853,N_14824);
xnor UO_518 (O_518,N_14892,N_14942);
nor UO_519 (O_519,N_14824,N_14960);
and UO_520 (O_520,N_14895,N_14892);
nand UO_521 (O_521,N_14860,N_14969);
nand UO_522 (O_522,N_14839,N_14931);
or UO_523 (O_523,N_14807,N_14933);
or UO_524 (O_524,N_14881,N_14905);
xor UO_525 (O_525,N_14908,N_14843);
and UO_526 (O_526,N_14839,N_14808);
xnor UO_527 (O_527,N_14814,N_14815);
nand UO_528 (O_528,N_14858,N_14880);
or UO_529 (O_529,N_14808,N_14818);
and UO_530 (O_530,N_14866,N_14895);
and UO_531 (O_531,N_14835,N_14965);
and UO_532 (O_532,N_14937,N_14985);
nor UO_533 (O_533,N_14870,N_14889);
and UO_534 (O_534,N_14966,N_14989);
and UO_535 (O_535,N_14858,N_14965);
and UO_536 (O_536,N_14809,N_14957);
and UO_537 (O_537,N_14925,N_14879);
xor UO_538 (O_538,N_14988,N_14810);
or UO_539 (O_539,N_14802,N_14919);
and UO_540 (O_540,N_14941,N_14817);
xor UO_541 (O_541,N_14844,N_14955);
or UO_542 (O_542,N_14885,N_14926);
nand UO_543 (O_543,N_14863,N_14890);
nor UO_544 (O_544,N_14913,N_14918);
nand UO_545 (O_545,N_14815,N_14877);
nand UO_546 (O_546,N_14928,N_14900);
and UO_547 (O_547,N_14949,N_14853);
and UO_548 (O_548,N_14824,N_14889);
and UO_549 (O_549,N_14875,N_14920);
nor UO_550 (O_550,N_14852,N_14990);
xnor UO_551 (O_551,N_14979,N_14842);
or UO_552 (O_552,N_14944,N_14857);
nor UO_553 (O_553,N_14910,N_14926);
and UO_554 (O_554,N_14814,N_14837);
nor UO_555 (O_555,N_14863,N_14857);
xnor UO_556 (O_556,N_14844,N_14861);
and UO_557 (O_557,N_14977,N_14917);
or UO_558 (O_558,N_14918,N_14975);
nand UO_559 (O_559,N_14936,N_14967);
or UO_560 (O_560,N_14844,N_14970);
nor UO_561 (O_561,N_14971,N_14801);
or UO_562 (O_562,N_14872,N_14917);
or UO_563 (O_563,N_14837,N_14827);
or UO_564 (O_564,N_14801,N_14988);
and UO_565 (O_565,N_14801,N_14954);
nand UO_566 (O_566,N_14917,N_14981);
and UO_567 (O_567,N_14855,N_14810);
and UO_568 (O_568,N_14991,N_14961);
nor UO_569 (O_569,N_14949,N_14830);
and UO_570 (O_570,N_14869,N_14806);
nor UO_571 (O_571,N_14933,N_14860);
and UO_572 (O_572,N_14812,N_14857);
nor UO_573 (O_573,N_14895,N_14991);
nor UO_574 (O_574,N_14851,N_14971);
nand UO_575 (O_575,N_14932,N_14967);
nor UO_576 (O_576,N_14916,N_14926);
nor UO_577 (O_577,N_14955,N_14924);
xor UO_578 (O_578,N_14875,N_14999);
nand UO_579 (O_579,N_14917,N_14881);
nand UO_580 (O_580,N_14922,N_14893);
and UO_581 (O_581,N_14983,N_14867);
nand UO_582 (O_582,N_14821,N_14988);
xor UO_583 (O_583,N_14948,N_14930);
nor UO_584 (O_584,N_14952,N_14951);
xor UO_585 (O_585,N_14925,N_14858);
and UO_586 (O_586,N_14912,N_14876);
nor UO_587 (O_587,N_14810,N_14985);
nor UO_588 (O_588,N_14808,N_14973);
or UO_589 (O_589,N_14832,N_14872);
or UO_590 (O_590,N_14992,N_14943);
and UO_591 (O_591,N_14860,N_14944);
xor UO_592 (O_592,N_14855,N_14869);
nor UO_593 (O_593,N_14911,N_14988);
nand UO_594 (O_594,N_14964,N_14858);
nand UO_595 (O_595,N_14984,N_14804);
nor UO_596 (O_596,N_14807,N_14973);
nand UO_597 (O_597,N_14910,N_14849);
nand UO_598 (O_598,N_14949,N_14891);
or UO_599 (O_599,N_14907,N_14943);
and UO_600 (O_600,N_14888,N_14936);
xor UO_601 (O_601,N_14880,N_14877);
and UO_602 (O_602,N_14872,N_14890);
nor UO_603 (O_603,N_14867,N_14973);
or UO_604 (O_604,N_14824,N_14990);
or UO_605 (O_605,N_14958,N_14930);
nor UO_606 (O_606,N_14813,N_14971);
nor UO_607 (O_607,N_14829,N_14990);
xor UO_608 (O_608,N_14857,N_14845);
nand UO_609 (O_609,N_14906,N_14920);
and UO_610 (O_610,N_14819,N_14941);
or UO_611 (O_611,N_14950,N_14901);
nand UO_612 (O_612,N_14870,N_14925);
and UO_613 (O_613,N_14941,N_14982);
xnor UO_614 (O_614,N_14872,N_14918);
xnor UO_615 (O_615,N_14883,N_14980);
xnor UO_616 (O_616,N_14997,N_14892);
and UO_617 (O_617,N_14835,N_14856);
and UO_618 (O_618,N_14815,N_14947);
xnor UO_619 (O_619,N_14830,N_14881);
nor UO_620 (O_620,N_14953,N_14839);
xnor UO_621 (O_621,N_14885,N_14879);
nand UO_622 (O_622,N_14833,N_14878);
and UO_623 (O_623,N_14880,N_14932);
nor UO_624 (O_624,N_14936,N_14871);
nor UO_625 (O_625,N_14930,N_14980);
xnor UO_626 (O_626,N_14917,N_14932);
nor UO_627 (O_627,N_14969,N_14988);
or UO_628 (O_628,N_14815,N_14809);
nand UO_629 (O_629,N_14960,N_14864);
nand UO_630 (O_630,N_14997,N_14885);
xnor UO_631 (O_631,N_14918,N_14814);
nand UO_632 (O_632,N_14813,N_14977);
and UO_633 (O_633,N_14919,N_14892);
or UO_634 (O_634,N_14809,N_14923);
nand UO_635 (O_635,N_14984,N_14906);
nor UO_636 (O_636,N_14819,N_14984);
nor UO_637 (O_637,N_14959,N_14846);
or UO_638 (O_638,N_14943,N_14989);
xnor UO_639 (O_639,N_14927,N_14988);
nor UO_640 (O_640,N_14859,N_14936);
nor UO_641 (O_641,N_14950,N_14913);
nor UO_642 (O_642,N_14999,N_14859);
or UO_643 (O_643,N_14960,N_14818);
nand UO_644 (O_644,N_14900,N_14807);
or UO_645 (O_645,N_14854,N_14812);
xnor UO_646 (O_646,N_14873,N_14901);
xnor UO_647 (O_647,N_14888,N_14912);
nor UO_648 (O_648,N_14977,N_14901);
nand UO_649 (O_649,N_14888,N_14817);
xnor UO_650 (O_650,N_14849,N_14970);
xnor UO_651 (O_651,N_14995,N_14814);
nand UO_652 (O_652,N_14915,N_14894);
nand UO_653 (O_653,N_14909,N_14998);
xor UO_654 (O_654,N_14870,N_14850);
and UO_655 (O_655,N_14855,N_14934);
and UO_656 (O_656,N_14983,N_14852);
nand UO_657 (O_657,N_14919,N_14962);
or UO_658 (O_658,N_14999,N_14805);
or UO_659 (O_659,N_14890,N_14990);
nor UO_660 (O_660,N_14869,N_14966);
nor UO_661 (O_661,N_14800,N_14850);
nor UO_662 (O_662,N_14891,N_14908);
xor UO_663 (O_663,N_14812,N_14976);
xor UO_664 (O_664,N_14856,N_14908);
or UO_665 (O_665,N_14979,N_14943);
and UO_666 (O_666,N_14929,N_14985);
xor UO_667 (O_667,N_14872,N_14991);
xnor UO_668 (O_668,N_14826,N_14891);
or UO_669 (O_669,N_14872,N_14876);
and UO_670 (O_670,N_14935,N_14885);
or UO_671 (O_671,N_14809,N_14947);
nor UO_672 (O_672,N_14812,N_14893);
or UO_673 (O_673,N_14892,N_14943);
nand UO_674 (O_674,N_14901,N_14918);
or UO_675 (O_675,N_14997,N_14973);
xor UO_676 (O_676,N_14952,N_14899);
and UO_677 (O_677,N_14827,N_14927);
nor UO_678 (O_678,N_14916,N_14897);
nand UO_679 (O_679,N_14821,N_14825);
and UO_680 (O_680,N_14999,N_14908);
and UO_681 (O_681,N_14976,N_14900);
and UO_682 (O_682,N_14940,N_14865);
or UO_683 (O_683,N_14943,N_14913);
and UO_684 (O_684,N_14806,N_14839);
nand UO_685 (O_685,N_14842,N_14871);
and UO_686 (O_686,N_14974,N_14878);
nand UO_687 (O_687,N_14841,N_14907);
and UO_688 (O_688,N_14989,N_14895);
nor UO_689 (O_689,N_14899,N_14938);
nor UO_690 (O_690,N_14811,N_14932);
xnor UO_691 (O_691,N_14816,N_14818);
or UO_692 (O_692,N_14816,N_14888);
and UO_693 (O_693,N_14879,N_14977);
xnor UO_694 (O_694,N_14808,N_14959);
nor UO_695 (O_695,N_14997,N_14907);
xor UO_696 (O_696,N_14856,N_14905);
or UO_697 (O_697,N_14819,N_14826);
xor UO_698 (O_698,N_14900,N_14876);
xor UO_699 (O_699,N_14905,N_14826);
nor UO_700 (O_700,N_14972,N_14802);
nor UO_701 (O_701,N_14932,N_14962);
and UO_702 (O_702,N_14837,N_14854);
xor UO_703 (O_703,N_14914,N_14986);
xor UO_704 (O_704,N_14876,N_14915);
xnor UO_705 (O_705,N_14839,N_14952);
nand UO_706 (O_706,N_14812,N_14985);
xor UO_707 (O_707,N_14854,N_14934);
and UO_708 (O_708,N_14909,N_14958);
or UO_709 (O_709,N_14978,N_14866);
nand UO_710 (O_710,N_14919,N_14874);
nand UO_711 (O_711,N_14853,N_14881);
nor UO_712 (O_712,N_14804,N_14910);
nand UO_713 (O_713,N_14919,N_14880);
and UO_714 (O_714,N_14955,N_14873);
and UO_715 (O_715,N_14877,N_14827);
and UO_716 (O_716,N_14927,N_14835);
nand UO_717 (O_717,N_14826,N_14955);
nand UO_718 (O_718,N_14901,N_14903);
and UO_719 (O_719,N_14962,N_14862);
nand UO_720 (O_720,N_14940,N_14806);
nor UO_721 (O_721,N_14934,N_14952);
and UO_722 (O_722,N_14834,N_14853);
or UO_723 (O_723,N_14808,N_14835);
xor UO_724 (O_724,N_14980,N_14993);
nor UO_725 (O_725,N_14856,N_14898);
nor UO_726 (O_726,N_14848,N_14890);
nor UO_727 (O_727,N_14843,N_14938);
nor UO_728 (O_728,N_14883,N_14967);
xnor UO_729 (O_729,N_14944,N_14940);
or UO_730 (O_730,N_14833,N_14955);
nand UO_731 (O_731,N_14989,N_14974);
nand UO_732 (O_732,N_14930,N_14835);
xnor UO_733 (O_733,N_14876,N_14845);
and UO_734 (O_734,N_14806,N_14907);
and UO_735 (O_735,N_14841,N_14940);
nand UO_736 (O_736,N_14800,N_14867);
xnor UO_737 (O_737,N_14955,N_14961);
xnor UO_738 (O_738,N_14882,N_14836);
nand UO_739 (O_739,N_14986,N_14805);
xor UO_740 (O_740,N_14861,N_14833);
and UO_741 (O_741,N_14992,N_14805);
xor UO_742 (O_742,N_14863,N_14852);
nor UO_743 (O_743,N_14800,N_14949);
and UO_744 (O_744,N_14825,N_14849);
xnor UO_745 (O_745,N_14976,N_14892);
nand UO_746 (O_746,N_14990,N_14816);
and UO_747 (O_747,N_14860,N_14926);
xor UO_748 (O_748,N_14888,N_14910);
nor UO_749 (O_749,N_14915,N_14882);
or UO_750 (O_750,N_14842,N_14989);
nand UO_751 (O_751,N_14812,N_14890);
xnor UO_752 (O_752,N_14993,N_14968);
and UO_753 (O_753,N_14910,N_14824);
nor UO_754 (O_754,N_14964,N_14981);
nand UO_755 (O_755,N_14931,N_14861);
xor UO_756 (O_756,N_14811,N_14823);
nand UO_757 (O_757,N_14932,N_14907);
nor UO_758 (O_758,N_14989,N_14818);
nand UO_759 (O_759,N_14851,N_14959);
nand UO_760 (O_760,N_14814,N_14810);
and UO_761 (O_761,N_14837,N_14824);
nor UO_762 (O_762,N_14945,N_14890);
nor UO_763 (O_763,N_14858,N_14949);
and UO_764 (O_764,N_14947,N_14831);
nor UO_765 (O_765,N_14934,N_14832);
and UO_766 (O_766,N_14925,N_14902);
xor UO_767 (O_767,N_14855,N_14978);
and UO_768 (O_768,N_14888,N_14812);
nor UO_769 (O_769,N_14990,N_14870);
and UO_770 (O_770,N_14833,N_14801);
nand UO_771 (O_771,N_14880,N_14916);
nand UO_772 (O_772,N_14960,N_14997);
nor UO_773 (O_773,N_14955,N_14990);
or UO_774 (O_774,N_14894,N_14893);
nor UO_775 (O_775,N_14938,N_14915);
xnor UO_776 (O_776,N_14967,N_14991);
nand UO_777 (O_777,N_14996,N_14861);
and UO_778 (O_778,N_14887,N_14912);
or UO_779 (O_779,N_14946,N_14965);
xor UO_780 (O_780,N_14815,N_14847);
xnor UO_781 (O_781,N_14886,N_14951);
nor UO_782 (O_782,N_14987,N_14996);
nand UO_783 (O_783,N_14942,N_14928);
nor UO_784 (O_784,N_14931,N_14965);
nand UO_785 (O_785,N_14982,N_14907);
xnor UO_786 (O_786,N_14849,N_14871);
nor UO_787 (O_787,N_14963,N_14988);
xor UO_788 (O_788,N_14857,N_14875);
nand UO_789 (O_789,N_14945,N_14979);
and UO_790 (O_790,N_14950,N_14898);
xnor UO_791 (O_791,N_14804,N_14986);
xor UO_792 (O_792,N_14974,N_14875);
xnor UO_793 (O_793,N_14944,N_14834);
or UO_794 (O_794,N_14801,N_14994);
xnor UO_795 (O_795,N_14915,N_14855);
or UO_796 (O_796,N_14832,N_14833);
nand UO_797 (O_797,N_14917,N_14887);
nand UO_798 (O_798,N_14945,N_14981);
nor UO_799 (O_799,N_14889,N_14937);
xnor UO_800 (O_800,N_14881,N_14982);
or UO_801 (O_801,N_14957,N_14884);
nand UO_802 (O_802,N_14918,N_14955);
or UO_803 (O_803,N_14834,N_14841);
or UO_804 (O_804,N_14862,N_14966);
or UO_805 (O_805,N_14832,N_14921);
nor UO_806 (O_806,N_14802,N_14833);
or UO_807 (O_807,N_14888,N_14860);
or UO_808 (O_808,N_14884,N_14947);
and UO_809 (O_809,N_14825,N_14872);
nor UO_810 (O_810,N_14901,N_14820);
xnor UO_811 (O_811,N_14959,N_14954);
nand UO_812 (O_812,N_14899,N_14872);
or UO_813 (O_813,N_14999,N_14876);
nor UO_814 (O_814,N_14967,N_14954);
nor UO_815 (O_815,N_14812,N_14972);
or UO_816 (O_816,N_14961,N_14831);
xor UO_817 (O_817,N_14902,N_14864);
or UO_818 (O_818,N_14818,N_14998);
nor UO_819 (O_819,N_14930,N_14969);
or UO_820 (O_820,N_14900,N_14835);
and UO_821 (O_821,N_14963,N_14809);
and UO_822 (O_822,N_14936,N_14801);
or UO_823 (O_823,N_14815,N_14982);
nand UO_824 (O_824,N_14878,N_14828);
or UO_825 (O_825,N_14831,N_14834);
and UO_826 (O_826,N_14953,N_14899);
or UO_827 (O_827,N_14913,N_14830);
xnor UO_828 (O_828,N_14810,N_14948);
nand UO_829 (O_829,N_14857,N_14895);
nor UO_830 (O_830,N_14836,N_14953);
nand UO_831 (O_831,N_14977,N_14906);
nand UO_832 (O_832,N_14814,N_14872);
nor UO_833 (O_833,N_14800,N_14871);
nand UO_834 (O_834,N_14825,N_14943);
or UO_835 (O_835,N_14890,N_14859);
and UO_836 (O_836,N_14828,N_14833);
and UO_837 (O_837,N_14808,N_14934);
xor UO_838 (O_838,N_14847,N_14884);
xor UO_839 (O_839,N_14845,N_14975);
nor UO_840 (O_840,N_14917,N_14877);
xor UO_841 (O_841,N_14935,N_14874);
nand UO_842 (O_842,N_14916,N_14978);
nor UO_843 (O_843,N_14901,N_14967);
nand UO_844 (O_844,N_14854,N_14855);
xnor UO_845 (O_845,N_14995,N_14946);
xnor UO_846 (O_846,N_14857,N_14983);
or UO_847 (O_847,N_14872,N_14864);
xnor UO_848 (O_848,N_14940,N_14923);
or UO_849 (O_849,N_14818,N_14886);
nor UO_850 (O_850,N_14998,N_14810);
nand UO_851 (O_851,N_14809,N_14996);
nand UO_852 (O_852,N_14943,N_14948);
or UO_853 (O_853,N_14972,N_14911);
or UO_854 (O_854,N_14853,N_14898);
xor UO_855 (O_855,N_14875,N_14900);
and UO_856 (O_856,N_14855,N_14904);
nand UO_857 (O_857,N_14854,N_14902);
and UO_858 (O_858,N_14823,N_14805);
and UO_859 (O_859,N_14836,N_14942);
nand UO_860 (O_860,N_14912,N_14914);
nor UO_861 (O_861,N_14883,N_14891);
or UO_862 (O_862,N_14990,N_14894);
and UO_863 (O_863,N_14970,N_14846);
and UO_864 (O_864,N_14850,N_14927);
nand UO_865 (O_865,N_14869,N_14823);
and UO_866 (O_866,N_14919,N_14916);
and UO_867 (O_867,N_14989,N_14871);
and UO_868 (O_868,N_14922,N_14977);
nor UO_869 (O_869,N_14824,N_14991);
nor UO_870 (O_870,N_14852,N_14935);
nor UO_871 (O_871,N_14937,N_14847);
nor UO_872 (O_872,N_14886,N_14861);
and UO_873 (O_873,N_14971,N_14987);
and UO_874 (O_874,N_14924,N_14821);
xnor UO_875 (O_875,N_14956,N_14898);
nand UO_876 (O_876,N_14813,N_14963);
and UO_877 (O_877,N_14865,N_14906);
nor UO_878 (O_878,N_14863,N_14940);
nand UO_879 (O_879,N_14997,N_14918);
nand UO_880 (O_880,N_14836,N_14920);
or UO_881 (O_881,N_14880,N_14854);
xor UO_882 (O_882,N_14900,N_14989);
or UO_883 (O_883,N_14870,N_14950);
nor UO_884 (O_884,N_14815,N_14845);
xnor UO_885 (O_885,N_14847,N_14998);
or UO_886 (O_886,N_14931,N_14977);
nand UO_887 (O_887,N_14929,N_14874);
or UO_888 (O_888,N_14876,N_14987);
xor UO_889 (O_889,N_14903,N_14990);
nand UO_890 (O_890,N_14985,N_14942);
or UO_891 (O_891,N_14970,N_14823);
nor UO_892 (O_892,N_14972,N_14888);
nand UO_893 (O_893,N_14878,N_14849);
xor UO_894 (O_894,N_14831,N_14812);
xor UO_895 (O_895,N_14921,N_14882);
xnor UO_896 (O_896,N_14942,N_14890);
nor UO_897 (O_897,N_14920,N_14874);
nand UO_898 (O_898,N_14956,N_14847);
xor UO_899 (O_899,N_14903,N_14912);
nand UO_900 (O_900,N_14997,N_14855);
nand UO_901 (O_901,N_14945,N_14906);
and UO_902 (O_902,N_14909,N_14954);
nand UO_903 (O_903,N_14896,N_14865);
xnor UO_904 (O_904,N_14949,N_14870);
xnor UO_905 (O_905,N_14821,N_14857);
nand UO_906 (O_906,N_14886,N_14894);
and UO_907 (O_907,N_14827,N_14807);
and UO_908 (O_908,N_14847,N_14960);
or UO_909 (O_909,N_14804,N_14902);
xnor UO_910 (O_910,N_14978,N_14973);
or UO_911 (O_911,N_14847,N_14975);
xor UO_912 (O_912,N_14864,N_14985);
or UO_913 (O_913,N_14858,N_14804);
and UO_914 (O_914,N_14880,N_14953);
and UO_915 (O_915,N_14806,N_14942);
and UO_916 (O_916,N_14893,N_14966);
or UO_917 (O_917,N_14891,N_14933);
nor UO_918 (O_918,N_14899,N_14871);
nor UO_919 (O_919,N_14918,N_14946);
or UO_920 (O_920,N_14812,N_14887);
or UO_921 (O_921,N_14958,N_14886);
or UO_922 (O_922,N_14956,N_14991);
or UO_923 (O_923,N_14937,N_14848);
and UO_924 (O_924,N_14816,N_14886);
nand UO_925 (O_925,N_14857,N_14945);
or UO_926 (O_926,N_14987,N_14885);
xnor UO_927 (O_927,N_14867,N_14884);
and UO_928 (O_928,N_14891,N_14970);
or UO_929 (O_929,N_14824,N_14862);
and UO_930 (O_930,N_14935,N_14952);
or UO_931 (O_931,N_14808,N_14844);
and UO_932 (O_932,N_14817,N_14805);
nor UO_933 (O_933,N_14850,N_14966);
and UO_934 (O_934,N_14990,N_14826);
nor UO_935 (O_935,N_14936,N_14965);
nand UO_936 (O_936,N_14851,N_14955);
or UO_937 (O_937,N_14861,N_14824);
nor UO_938 (O_938,N_14976,N_14973);
nand UO_939 (O_939,N_14945,N_14891);
and UO_940 (O_940,N_14954,N_14816);
or UO_941 (O_941,N_14967,N_14818);
and UO_942 (O_942,N_14950,N_14854);
nor UO_943 (O_943,N_14888,N_14802);
and UO_944 (O_944,N_14862,N_14917);
or UO_945 (O_945,N_14832,N_14917);
and UO_946 (O_946,N_14891,N_14865);
or UO_947 (O_947,N_14964,N_14987);
nand UO_948 (O_948,N_14826,N_14837);
xor UO_949 (O_949,N_14998,N_14914);
and UO_950 (O_950,N_14889,N_14953);
xnor UO_951 (O_951,N_14958,N_14849);
nor UO_952 (O_952,N_14877,N_14826);
or UO_953 (O_953,N_14923,N_14846);
nor UO_954 (O_954,N_14965,N_14845);
and UO_955 (O_955,N_14903,N_14875);
nand UO_956 (O_956,N_14911,N_14800);
nor UO_957 (O_957,N_14889,N_14967);
and UO_958 (O_958,N_14953,N_14936);
and UO_959 (O_959,N_14809,N_14825);
and UO_960 (O_960,N_14830,N_14937);
nand UO_961 (O_961,N_14837,N_14907);
xnor UO_962 (O_962,N_14826,N_14907);
or UO_963 (O_963,N_14809,N_14932);
and UO_964 (O_964,N_14880,N_14982);
and UO_965 (O_965,N_14951,N_14955);
nand UO_966 (O_966,N_14838,N_14899);
nor UO_967 (O_967,N_14843,N_14809);
xnor UO_968 (O_968,N_14935,N_14903);
nand UO_969 (O_969,N_14875,N_14924);
nand UO_970 (O_970,N_14819,N_14885);
xnor UO_971 (O_971,N_14957,N_14846);
or UO_972 (O_972,N_14859,N_14953);
xnor UO_973 (O_973,N_14903,N_14818);
and UO_974 (O_974,N_14918,N_14819);
nor UO_975 (O_975,N_14891,N_14924);
nor UO_976 (O_976,N_14898,N_14962);
or UO_977 (O_977,N_14880,N_14888);
nor UO_978 (O_978,N_14953,N_14938);
or UO_979 (O_979,N_14857,N_14806);
nor UO_980 (O_980,N_14935,N_14989);
or UO_981 (O_981,N_14923,N_14917);
nand UO_982 (O_982,N_14866,N_14811);
xor UO_983 (O_983,N_14971,N_14959);
and UO_984 (O_984,N_14845,N_14858);
xnor UO_985 (O_985,N_14922,N_14863);
or UO_986 (O_986,N_14862,N_14909);
and UO_987 (O_987,N_14817,N_14884);
and UO_988 (O_988,N_14812,N_14951);
or UO_989 (O_989,N_14952,N_14835);
nor UO_990 (O_990,N_14954,N_14838);
nand UO_991 (O_991,N_14842,N_14860);
nor UO_992 (O_992,N_14911,N_14987);
xor UO_993 (O_993,N_14877,N_14805);
xor UO_994 (O_994,N_14989,N_14959);
and UO_995 (O_995,N_14892,N_14838);
xnor UO_996 (O_996,N_14907,N_14941);
or UO_997 (O_997,N_14803,N_14874);
nand UO_998 (O_998,N_14897,N_14933);
or UO_999 (O_999,N_14841,N_14992);
xnor UO_1000 (O_1000,N_14930,N_14935);
or UO_1001 (O_1001,N_14964,N_14988);
nand UO_1002 (O_1002,N_14816,N_14877);
and UO_1003 (O_1003,N_14940,N_14962);
and UO_1004 (O_1004,N_14970,N_14854);
xor UO_1005 (O_1005,N_14876,N_14875);
and UO_1006 (O_1006,N_14876,N_14907);
nor UO_1007 (O_1007,N_14932,N_14944);
and UO_1008 (O_1008,N_14834,N_14850);
and UO_1009 (O_1009,N_14881,N_14983);
or UO_1010 (O_1010,N_14978,N_14822);
or UO_1011 (O_1011,N_14932,N_14860);
and UO_1012 (O_1012,N_14908,N_14809);
or UO_1013 (O_1013,N_14942,N_14954);
nand UO_1014 (O_1014,N_14802,N_14925);
and UO_1015 (O_1015,N_14990,N_14976);
nand UO_1016 (O_1016,N_14903,N_14819);
xor UO_1017 (O_1017,N_14971,N_14932);
nor UO_1018 (O_1018,N_14988,N_14852);
and UO_1019 (O_1019,N_14966,N_14957);
and UO_1020 (O_1020,N_14991,N_14876);
xor UO_1021 (O_1021,N_14974,N_14939);
nor UO_1022 (O_1022,N_14972,N_14937);
or UO_1023 (O_1023,N_14908,N_14893);
nor UO_1024 (O_1024,N_14988,N_14984);
or UO_1025 (O_1025,N_14916,N_14840);
xor UO_1026 (O_1026,N_14847,N_14954);
or UO_1027 (O_1027,N_14920,N_14815);
nor UO_1028 (O_1028,N_14802,N_14885);
nor UO_1029 (O_1029,N_14817,N_14966);
nand UO_1030 (O_1030,N_14836,N_14843);
nand UO_1031 (O_1031,N_14946,N_14982);
nor UO_1032 (O_1032,N_14835,N_14997);
and UO_1033 (O_1033,N_14887,N_14862);
nor UO_1034 (O_1034,N_14906,N_14810);
and UO_1035 (O_1035,N_14872,N_14819);
and UO_1036 (O_1036,N_14911,N_14823);
and UO_1037 (O_1037,N_14886,N_14808);
or UO_1038 (O_1038,N_14881,N_14999);
xnor UO_1039 (O_1039,N_14884,N_14836);
xnor UO_1040 (O_1040,N_14808,N_14918);
or UO_1041 (O_1041,N_14976,N_14939);
or UO_1042 (O_1042,N_14896,N_14849);
nand UO_1043 (O_1043,N_14888,N_14832);
and UO_1044 (O_1044,N_14845,N_14944);
nand UO_1045 (O_1045,N_14905,N_14837);
xnor UO_1046 (O_1046,N_14866,N_14855);
or UO_1047 (O_1047,N_14984,N_14985);
xnor UO_1048 (O_1048,N_14855,N_14975);
and UO_1049 (O_1049,N_14996,N_14945);
and UO_1050 (O_1050,N_14945,N_14939);
nor UO_1051 (O_1051,N_14993,N_14871);
nor UO_1052 (O_1052,N_14824,N_14863);
nor UO_1053 (O_1053,N_14864,N_14932);
xor UO_1054 (O_1054,N_14832,N_14854);
xor UO_1055 (O_1055,N_14920,N_14900);
xor UO_1056 (O_1056,N_14948,N_14903);
and UO_1057 (O_1057,N_14835,N_14964);
nand UO_1058 (O_1058,N_14897,N_14950);
nand UO_1059 (O_1059,N_14924,N_14935);
xor UO_1060 (O_1060,N_14990,N_14972);
nand UO_1061 (O_1061,N_14875,N_14843);
nand UO_1062 (O_1062,N_14804,N_14838);
and UO_1063 (O_1063,N_14947,N_14861);
nor UO_1064 (O_1064,N_14902,N_14812);
and UO_1065 (O_1065,N_14975,N_14996);
or UO_1066 (O_1066,N_14840,N_14910);
nor UO_1067 (O_1067,N_14834,N_14906);
nor UO_1068 (O_1068,N_14895,N_14972);
nand UO_1069 (O_1069,N_14819,N_14995);
xor UO_1070 (O_1070,N_14913,N_14971);
and UO_1071 (O_1071,N_14917,N_14946);
nand UO_1072 (O_1072,N_14901,N_14965);
or UO_1073 (O_1073,N_14810,N_14832);
xnor UO_1074 (O_1074,N_14840,N_14914);
nor UO_1075 (O_1075,N_14833,N_14831);
xnor UO_1076 (O_1076,N_14903,N_14814);
and UO_1077 (O_1077,N_14844,N_14996);
nor UO_1078 (O_1078,N_14949,N_14847);
nand UO_1079 (O_1079,N_14967,N_14838);
or UO_1080 (O_1080,N_14818,N_14982);
or UO_1081 (O_1081,N_14877,N_14983);
nand UO_1082 (O_1082,N_14849,N_14895);
or UO_1083 (O_1083,N_14905,N_14997);
nor UO_1084 (O_1084,N_14840,N_14978);
and UO_1085 (O_1085,N_14827,N_14961);
and UO_1086 (O_1086,N_14987,N_14886);
nand UO_1087 (O_1087,N_14809,N_14805);
and UO_1088 (O_1088,N_14845,N_14882);
xor UO_1089 (O_1089,N_14912,N_14920);
and UO_1090 (O_1090,N_14888,N_14956);
nor UO_1091 (O_1091,N_14934,N_14833);
nand UO_1092 (O_1092,N_14994,N_14936);
nand UO_1093 (O_1093,N_14918,N_14864);
and UO_1094 (O_1094,N_14908,N_14939);
nand UO_1095 (O_1095,N_14896,N_14947);
xnor UO_1096 (O_1096,N_14909,N_14853);
xor UO_1097 (O_1097,N_14967,N_14925);
and UO_1098 (O_1098,N_14900,N_14911);
xnor UO_1099 (O_1099,N_14848,N_14989);
and UO_1100 (O_1100,N_14954,N_14844);
nor UO_1101 (O_1101,N_14801,N_14929);
nor UO_1102 (O_1102,N_14855,N_14951);
nand UO_1103 (O_1103,N_14971,N_14896);
nand UO_1104 (O_1104,N_14882,N_14840);
or UO_1105 (O_1105,N_14982,N_14877);
or UO_1106 (O_1106,N_14952,N_14827);
and UO_1107 (O_1107,N_14900,N_14926);
nand UO_1108 (O_1108,N_14840,N_14936);
nand UO_1109 (O_1109,N_14970,N_14973);
or UO_1110 (O_1110,N_14834,N_14820);
and UO_1111 (O_1111,N_14846,N_14885);
nand UO_1112 (O_1112,N_14976,N_14964);
or UO_1113 (O_1113,N_14943,N_14883);
nor UO_1114 (O_1114,N_14972,N_14967);
and UO_1115 (O_1115,N_14801,N_14912);
xnor UO_1116 (O_1116,N_14945,N_14810);
and UO_1117 (O_1117,N_14848,N_14836);
and UO_1118 (O_1118,N_14816,N_14960);
xnor UO_1119 (O_1119,N_14989,N_14978);
or UO_1120 (O_1120,N_14949,N_14931);
xor UO_1121 (O_1121,N_14980,N_14884);
nor UO_1122 (O_1122,N_14995,N_14823);
or UO_1123 (O_1123,N_14991,N_14852);
or UO_1124 (O_1124,N_14951,N_14872);
nor UO_1125 (O_1125,N_14839,N_14824);
and UO_1126 (O_1126,N_14862,N_14829);
nor UO_1127 (O_1127,N_14859,N_14899);
or UO_1128 (O_1128,N_14861,N_14877);
nand UO_1129 (O_1129,N_14877,N_14989);
or UO_1130 (O_1130,N_14969,N_14820);
and UO_1131 (O_1131,N_14926,N_14845);
or UO_1132 (O_1132,N_14803,N_14942);
nor UO_1133 (O_1133,N_14851,N_14895);
and UO_1134 (O_1134,N_14829,N_14848);
nor UO_1135 (O_1135,N_14940,N_14918);
and UO_1136 (O_1136,N_14891,N_14984);
nor UO_1137 (O_1137,N_14876,N_14810);
or UO_1138 (O_1138,N_14933,N_14836);
nand UO_1139 (O_1139,N_14930,N_14920);
nor UO_1140 (O_1140,N_14875,N_14835);
xnor UO_1141 (O_1141,N_14944,N_14967);
and UO_1142 (O_1142,N_14838,N_14975);
nor UO_1143 (O_1143,N_14960,N_14995);
or UO_1144 (O_1144,N_14862,N_14908);
or UO_1145 (O_1145,N_14855,N_14878);
xnor UO_1146 (O_1146,N_14988,N_14848);
nor UO_1147 (O_1147,N_14899,N_14823);
and UO_1148 (O_1148,N_14954,N_14962);
xor UO_1149 (O_1149,N_14891,N_14877);
or UO_1150 (O_1150,N_14996,N_14938);
nand UO_1151 (O_1151,N_14949,N_14869);
nor UO_1152 (O_1152,N_14912,N_14917);
or UO_1153 (O_1153,N_14996,N_14876);
or UO_1154 (O_1154,N_14866,N_14944);
or UO_1155 (O_1155,N_14926,N_14882);
nor UO_1156 (O_1156,N_14904,N_14974);
nand UO_1157 (O_1157,N_14803,N_14806);
and UO_1158 (O_1158,N_14972,N_14867);
nor UO_1159 (O_1159,N_14882,N_14838);
or UO_1160 (O_1160,N_14814,N_14859);
xnor UO_1161 (O_1161,N_14812,N_14944);
xor UO_1162 (O_1162,N_14800,N_14919);
and UO_1163 (O_1163,N_14871,N_14847);
nand UO_1164 (O_1164,N_14885,N_14904);
nor UO_1165 (O_1165,N_14903,N_14840);
or UO_1166 (O_1166,N_14829,N_14807);
or UO_1167 (O_1167,N_14848,N_14802);
nor UO_1168 (O_1168,N_14871,N_14998);
and UO_1169 (O_1169,N_14871,N_14987);
and UO_1170 (O_1170,N_14929,N_14880);
or UO_1171 (O_1171,N_14935,N_14945);
xnor UO_1172 (O_1172,N_14957,N_14862);
or UO_1173 (O_1173,N_14823,N_14950);
and UO_1174 (O_1174,N_14984,N_14821);
xnor UO_1175 (O_1175,N_14916,N_14835);
nand UO_1176 (O_1176,N_14828,N_14969);
xnor UO_1177 (O_1177,N_14981,N_14891);
xnor UO_1178 (O_1178,N_14882,N_14843);
or UO_1179 (O_1179,N_14936,N_14918);
xnor UO_1180 (O_1180,N_14831,N_14938);
nand UO_1181 (O_1181,N_14925,N_14853);
nor UO_1182 (O_1182,N_14805,N_14907);
nor UO_1183 (O_1183,N_14805,N_14991);
nand UO_1184 (O_1184,N_14935,N_14833);
xor UO_1185 (O_1185,N_14848,N_14977);
nor UO_1186 (O_1186,N_14871,N_14932);
nand UO_1187 (O_1187,N_14835,N_14896);
nor UO_1188 (O_1188,N_14896,N_14872);
nand UO_1189 (O_1189,N_14965,N_14919);
nor UO_1190 (O_1190,N_14969,N_14894);
or UO_1191 (O_1191,N_14858,N_14986);
or UO_1192 (O_1192,N_14974,N_14826);
or UO_1193 (O_1193,N_14859,N_14956);
nor UO_1194 (O_1194,N_14864,N_14978);
xnor UO_1195 (O_1195,N_14862,N_14893);
xor UO_1196 (O_1196,N_14885,N_14800);
nand UO_1197 (O_1197,N_14945,N_14870);
xnor UO_1198 (O_1198,N_14975,N_14946);
or UO_1199 (O_1199,N_14880,N_14987);
or UO_1200 (O_1200,N_14847,N_14955);
xor UO_1201 (O_1201,N_14982,N_14871);
or UO_1202 (O_1202,N_14888,N_14829);
nand UO_1203 (O_1203,N_14954,N_14896);
or UO_1204 (O_1204,N_14971,N_14917);
xnor UO_1205 (O_1205,N_14809,N_14942);
and UO_1206 (O_1206,N_14849,N_14851);
nand UO_1207 (O_1207,N_14801,N_14958);
xor UO_1208 (O_1208,N_14840,N_14977);
and UO_1209 (O_1209,N_14969,N_14842);
nor UO_1210 (O_1210,N_14941,N_14920);
nor UO_1211 (O_1211,N_14804,N_14932);
xor UO_1212 (O_1212,N_14977,N_14839);
and UO_1213 (O_1213,N_14884,N_14830);
nand UO_1214 (O_1214,N_14838,N_14998);
and UO_1215 (O_1215,N_14971,N_14962);
nand UO_1216 (O_1216,N_14832,N_14882);
nor UO_1217 (O_1217,N_14843,N_14990);
or UO_1218 (O_1218,N_14871,N_14841);
nor UO_1219 (O_1219,N_14936,N_14858);
nand UO_1220 (O_1220,N_14916,N_14944);
or UO_1221 (O_1221,N_14921,N_14847);
and UO_1222 (O_1222,N_14992,N_14950);
nor UO_1223 (O_1223,N_14875,N_14858);
and UO_1224 (O_1224,N_14830,N_14854);
xor UO_1225 (O_1225,N_14853,N_14899);
xor UO_1226 (O_1226,N_14927,N_14979);
or UO_1227 (O_1227,N_14995,N_14945);
xor UO_1228 (O_1228,N_14911,N_14934);
or UO_1229 (O_1229,N_14934,N_14880);
nand UO_1230 (O_1230,N_14845,N_14942);
or UO_1231 (O_1231,N_14983,N_14915);
nand UO_1232 (O_1232,N_14836,N_14854);
nor UO_1233 (O_1233,N_14972,N_14949);
and UO_1234 (O_1234,N_14801,N_14817);
and UO_1235 (O_1235,N_14837,N_14960);
nand UO_1236 (O_1236,N_14811,N_14842);
and UO_1237 (O_1237,N_14841,N_14809);
xor UO_1238 (O_1238,N_14974,N_14937);
xor UO_1239 (O_1239,N_14890,N_14877);
xnor UO_1240 (O_1240,N_14927,N_14980);
xnor UO_1241 (O_1241,N_14980,N_14996);
nor UO_1242 (O_1242,N_14971,N_14875);
nor UO_1243 (O_1243,N_14918,N_14920);
nand UO_1244 (O_1244,N_14865,N_14852);
nor UO_1245 (O_1245,N_14900,N_14806);
xnor UO_1246 (O_1246,N_14826,N_14890);
nand UO_1247 (O_1247,N_14806,N_14963);
or UO_1248 (O_1248,N_14965,N_14829);
and UO_1249 (O_1249,N_14953,N_14944);
nand UO_1250 (O_1250,N_14969,N_14954);
nand UO_1251 (O_1251,N_14928,N_14963);
nand UO_1252 (O_1252,N_14873,N_14804);
nand UO_1253 (O_1253,N_14895,N_14810);
nor UO_1254 (O_1254,N_14938,N_14829);
nand UO_1255 (O_1255,N_14917,N_14905);
or UO_1256 (O_1256,N_14831,N_14840);
nor UO_1257 (O_1257,N_14925,N_14960);
and UO_1258 (O_1258,N_14828,N_14968);
xor UO_1259 (O_1259,N_14802,N_14902);
nor UO_1260 (O_1260,N_14917,N_14803);
nor UO_1261 (O_1261,N_14833,N_14804);
or UO_1262 (O_1262,N_14959,N_14871);
or UO_1263 (O_1263,N_14849,N_14848);
nor UO_1264 (O_1264,N_14964,N_14882);
nand UO_1265 (O_1265,N_14990,N_14978);
xor UO_1266 (O_1266,N_14972,N_14947);
nor UO_1267 (O_1267,N_14948,N_14836);
nand UO_1268 (O_1268,N_14852,N_14903);
or UO_1269 (O_1269,N_14817,N_14848);
xnor UO_1270 (O_1270,N_14881,N_14973);
xor UO_1271 (O_1271,N_14920,N_14976);
nand UO_1272 (O_1272,N_14820,N_14885);
nand UO_1273 (O_1273,N_14812,N_14984);
nor UO_1274 (O_1274,N_14802,N_14963);
nand UO_1275 (O_1275,N_14887,N_14841);
or UO_1276 (O_1276,N_14857,N_14999);
nand UO_1277 (O_1277,N_14982,N_14985);
xor UO_1278 (O_1278,N_14968,N_14942);
nor UO_1279 (O_1279,N_14899,N_14955);
xnor UO_1280 (O_1280,N_14902,N_14801);
nand UO_1281 (O_1281,N_14949,N_14979);
xor UO_1282 (O_1282,N_14912,N_14951);
xnor UO_1283 (O_1283,N_14999,N_14998);
nor UO_1284 (O_1284,N_14932,N_14826);
and UO_1285 (O_1285,N_14869,N_14908);
nor UO_1286 (O_1286,N_14874,N_14862);
or UO_1287 (O_1287,N_14858,N_14824);
nor UO_1288 (O_1288,N_14916,N_14995);
xor UO_1289 (O_1289,N_14849,N_14999);
xor UO_1290 (O_1290,N_14950,N_14831);
xor UO_1291 (O_1291,N_14990,N_14822);
and UO_1292 (O_1292,N_14970,N_14922);
xnor UO_1293 (O_1293,N_14912,N_14853);
xor UO_1294 (O_1294,N_14861,N_14962);
and UO_1295 (O_1295,N_14955,N_14929);
or UO_1296 (O_1296,N_14873,N_14906);
nor UO_1297 (O_1297,N_14885,N_14912);
and UO_1298 (O_1298,N_14996,N_14880);
and UO_1299 (O_1299,N_14907,N_14990);
nand UO_1300 (O_1300,N_14805,N_14938);
nor UO_1301 (O_1301,N_14908,N_14824);
and UO_1302 (O_1302,N_14984,N_14987);
or UO_1303 (O_1303,N_14891,N_14853);
and UO_1304 (O_1304,N_14830,N_14899);
nand UO_1305 (O_1305,N_14994,N_14907);
nand UO_1306 (O_1306,N_14840,N_14853);
xnor UO_1307 (O_1307,N_14926,N_14867);
xor UO_1308 (O_1308,N_14900,N_14871);
or UO_1309 (O_1309,N_14906,N_14851);
and UO_1310 (O_1310,N_14840,N_14933);
nor UO_1311 (O_1311,N_14823,N_14827);
nor UO_1312 (O_1312,N_14838,N_14809);
and UO_1313 (O_1313,N_14852,N_14950);
and UO_1314 (O_1314,N_14971,N_14946);
nor UO_1315 (O_1315,N_14917,N_14939);
and UO_1316 (O_1316,N_14993,N_14920);
xnor UO_1317 (O_1317,N_14977,N_14950);
nand UO_1318 (O_1318,N_14903,N_14925);
or UO_1319 (O_1319,N_14991,N_14832);
nor UO_1320 (O_1320,N_14833,N_14952);
or UO_1321 (O_1321,N_14886,N_14908);
nor UO_1322 (O_1322,N_14996,N_14982);
xor UO_1323 (O_1323,N_14820,N_14947);
xnor UO_1324 (O_1324,N_14872,N_14816);
nor UO_1325 (O_1325,N_14865,N_14803);
and UO_1326 (O_1326,N_14944,N_14880);
or UO_1327 (O_1327,N_14956,N_14937);
or UO_1328 (O_1328,N_14920,N_14929);
nor UO_1329 (O_1329,N_14877,N_14961);
nand UO_1330 (O_1330,N_14900,N_14881);
nand UO_1331 (O_1331,N_14810,N_14965);
or UO_1332 (O_1332,N_14851,N_14985);
nor UO_1333 (O_1333,N_14989,N_14986);
xnor UO_1334 (O_1334,N_14854,N_14875);
xnor UO_1335 (O_1335,N_14893,N_14884);
nand UO_1336 (O_1336,N_14981,N_14864);
or UO_1337 (O_1337,N_14949,N_14857);
or UO_1338 (O_1338,N_14863,N_14887);
or UO_1339 (O_1339,N_14809,N_14877);
xor UO_1340 (O_1340,N_14925,N_14815);
or UO_1341 (O_1341,N_14974,N_14999);
xnor UO_1342 (O_1342,N_14888,N_14941);
and UO_1343 (O_1343,N_14956,N_14831);
nor UO_1344 (O_1344,N_14878,N_14979);
and UO_1345 (O_1345,N_14863,N_14913);
xnor UO_1346 (O_1346,N_14888,N_14943);
xor UO_1347 (O_1347,N_14865,N_14960);
nor UO_1348 (O_1348,N_14819,N_14934);
or UO_1349 (O_1349,N_14977,N_14959);
and UO_1350 (O_1350,N_14832,N_14994);
xnor UO_1351 (O_1351,N_14850,N_14810);
and UO_1352 (O_1352,N_14826,N_14836);
nor UO_1353 (O_1353,N_14990,N_14954);
or UO_1354 (O_1354,N_14958,N_14892);
or UO_1355 (O_1355,N_14868,N_14905);
xnor UO_1356 (O_1356,N_14879,N_14900);
nand UO_1357 (O_1357,N_14843,N_14927);
nand UO_1358 (O_1358,N_14870,N_14928);
and UO_1359 (O_1359,N_14818,N_14820);
nand UO_1360 (O_1360,N_14896,N_14884);
or UO_1361 (O_1361,N_14918,N_14985);
nor UO_1362 (O_1362,N_14833,N_14906);
xor UO_1363 (O_1363,N_14838,N_14821);
nor UO_1364 (O_1364,N_14920,N_14923);
or UO_1365 (O_1365,N_14859,N_14839);
nor UO_1366 (O_1366,N_14942,N_14832);
nor UO_1367 (O_1367,N_14984,N_14968);
nor UO_1368 (O_1368,N_14894,N_14941);
nand UO_1369 (O_1369,N_14842,N_14950);
and UO_1370 (O_1370,N_14826,N_14831);
xor UO_1371 (O_1371,N_14822,N_14994);
nor UO_1372 (O_1372,N_14837,N_14977);
and UO_1373 (O_1373,N_14989,N_14908);
nor UO_1374 (O_1374,N_14909,N_14920);
nor UO_1375 (O_1375,N_14925,N_14817);
nand UO_1376 (O_1376,N_14866,N_14834);
and UO_1377 (O_1377,N_14935,N_14846);
or UO_1378 (O_1378,N_14859,N_14984);
nand UO_1379 (O_1379,N_14957,N_14961);
nand UO_1380 (O_1380,N_14877,N_14818);
and UO_1381 (O_1381,N_14934,N_14840);
and UO_1382 (O_1382,N_14815,N_14980);
nand UO_1383 (O_1383,N_14884,N_14915);
or UO_1384 (O_1384,N_14947,N_14854);
and UO_1385 (O_1385,N_14977,N_14989);
or UO_1386 (O_1386,N_14874,N_14840);
and UO_1387 (O_1387,N_14800,N_14997);
xor UO_1388 (O_1388,N_14910,N_14981);
nor UO_1389 (O_1389,N_14973,N_14897);
or UO_1390 (O_1390,N_14865,N_14939);
and UO_1391 (O_1391,N_14984,N_14901);
nor UO_1392 (O_1392,N_14987,N_14836);
xnor UO_1393 (O_1393,N_14821,N_14895);
nand UO_1394 (O_1394,N_14940,N_14872);
or UO_1395 (O_1395,N_14917,N_14826);
nand UO_1396 (O_1396,N_14923,N_14856);
nor UO_1397 (O_1397,N_14934,N_14815);
nor UO_1398 (O_1398,N_14965,N_14851);
xnor UO_1399 (O_1399,N_14841,N_14933);
xor UO_1400 (O_1400,N_14843,N_14825);
and UO_1401 (O_1401,N_14834,N_14869);
nor UO_1402 (O_1402,N_14850,N_14817);
and UO_1403 (O_1403,N_14940,N_14867);
nor UO_1404 (O_1404,N_14941,N_14881);
nand UO_1405 (O_1405,N_14910,N_14833);
nand UO_1406 (O_1406,N_14908,N_14840);
nor UO_1407 (O_1407,N_14978,N_14844);
xnor UO_1408 (O_1408,N_14906,N_14816);
nor UO_1409 (O_1409,N_14845,N_14990);
nand UO_1410 (O_1410,N_14906,N_14970);
xnor UO_1411 (O_1411,N_14888,N_14903);
xnor UO_1412 (O_1412,N_14952,N_14884);
and UO_1413 (O_1413,N_14933,N_14894);
nand UO_1414 (O_1414,N_14993,N_14831);
and UO_1415 (O_1415,N_14913,N_14800);
nand UO_1416 (O_1416,N_14925,N_14928);
or UO_1417 (O_1417,N_14920,N_14980);
xor UO_1418 (O_1418,N_14848,N_14832);
nor UO_1419 (O_1419,N_14884,N_14837);
xor UO_1420 (O_1420,N_14999,N_14923);
nand UO_1421 (O_1421,N_14956,N_14965);
and UO_1422 (O_1422,N_14909,N_14916);
or UO_1423 (O_1423,N_14804,N_14975);
and UO_1424 (O_1424,N_14994,N_14970);
nand UO_1425 (O_1425,N_14839,N_14945);
nor UO_1426 (O_1426,N_14940,N_14820);
nor UO_1427 (O_1427,N_14872,N_14937);
nor UO_1428 (O_1428,N_14869,N_14993);
nor UO_1429 (O_1429,N_14934,N_14988);
xor UO_1430 (O_1430,N_14968,N_14949);
nor UO_1431 (O_1431,N_14993,N_14997);
and UO_1432 (O_1432,N_14821,N_14874);
and UO_1433 (O_1433,N_14874,N_14905);
xor UO_1434 (O_1434,N_14846,N_14905);
or UO_1435 (O_1435,N_14855,N_14965);
nand UO_1436 (O_1436,N_14907,N_14879);
or UO_1437 (O_1437,N_14843,N_14979);
nor UO_1438 (O_1438,N_14865,N_14811);
nor UO_1439 (O_1439,N_14850,N_14904);
nand UO_1440 (O_1440,N_14983,N_14953);
nand UO_1441 (O_1441,N_14854,N_14829);
nor UO_1442 (O_1442,N_14835,N_14922);
or UO_1443 (O_1443,N_14843,N_14925);
and UO_1444 (O_1444,N_14800,N_14992);
or UO_1445 (O_1445,N_14872,N_14863);
xor UO_1446 (O_1446,N_14944,N_14982);
and UO_1447 (O_1447,N_14884,N_14841);
xor UO_1448 (O_1448,N_14852,N_14877);
or UO_1449 (O_1449,N_14829,N_14993);
or UO_1450 (O_1450,N_14904,N_14836);
or UO_1451 (O_1451,N_14964,N_14821);
nand UO_1452 (O_1452,N_14935,N_14921);
or UO_1453 (O_1453,N_14891,N_14926);
xnor UO_1454 (O_1454,N_14953,N_14826);
nand UO_1455 (O_1455,N_14952,N_14808);
nand UO_1456 (O_1456,N_14883,N_14846);
nand UO_1457 (O_1457,N_14971,N_14933);
nor UO_1458 (O_1458,N_14939,N_14970);
and UO_1459 (O_1459,N_14898,N_14870);
nor UO_1460 (O_1460,N_14949,N_14844);
xnor UO_1461 (O_1461,N_14946,N_14880);
nand UO_1462 (O_1462,N_14872,N_14839);
nor UO_1463 (O_1463,N_14843,N_14973);
or UO_1464 (O_1464,N_14890,N_14907);
nor UO_1465 (O_1465,N_14930,N_14858);
nand UO_1466 (O_1466,N_14964,N_14972);
nor UO_1467 (O_1467,N_14871,N_14862);
nor UO_1468 (O_1468,N_14858,N_14903);
nand UO_1469 (O_1469,N_14939,N_14881);
xor UO_1470 (O_1470,N_14947,N_14910);
or UO_1471 (O_1471,N_14896,N_14937);
nand UO_1472 (O_1472,N_14937,N_14803);
xor UO_1473 (O_1473,N_14943,N_14971);
and UO_1474 (O_1474,N_14971,N_14852);
xor UO_1475 (O_1475,N_14929,N_14919);
xor UO_1476 (O_1476,N_14814,N_14802);
or UO_1477 (O_1477,N_14945,N_14848);
or UO_1478 (O_1478,N_14932,N_14940);
and UO_1479 (O_1479,N_14821,N_14963);
and UO_1480 (O_1480,N_14802,N_14842);
and UO_1481 (O_1481,N_14874,N_14916);
nand UO_1482 (O_1482,N_14834,N_14868);
or UO_1483 (O_1483,N_14993,N_14861);
xor UO_1484 (O_1484,N_14926,N_14895);
nor UO_1485 (O_1485,N_14915,N_14930);
xnor UO_1486 (O_1486,N_14958,N_14816);
and UO_1487 (O_1487,N_14978,N_14956);
nor UO_1488 (O_1488,N_14803,N_14948);
and UO_1489 (O_1489,N_14834,N_14832);
nand UO_1490 (O_1490,N_14902,N_14816);
xor UO_1491 (O_1491,N_14816,N_14923);
and UO_1492 (O_1492,N_14985,N_14818);
nand UO_1493 (O_1493,N_14834,N_14875);
nand UO_1494 (O_1494,N_14991,N_14984);
and UO_1495 (O_1495,N_14885,N_14944);
xnor UO_1496 (O_1496,N_14913,N_14990);
and UO_1497 (O_1497,N_14970,N_14967);
or UO_1498 (O_1498,N_14884,N_14965);
and UO_1499 (O_1499,N_14952,N_14868);
nor UO_1500 (O_1500,N_14955,N_14811);
nand UO_1501 (O_1501,N_14883,N_14914);
nand UO_1502 (O_1502,N_14911,N_14852);
nor UO_1503 (O_1503,N_14836,N_14860);
or UO_1504 (O_1504,N_14820,N_14902);
xor UO_1505 (O_1505,N_14973,N_14865);
xor UO_1506 (O_1506,N_14839,N_14923);
or UO_1507 (O_1507,N_14857,N_14965);
and UO_1508 (O_1508,N_14950,N_14905);
xor UO_1509 (O_1509,N_14907,N_14804);
or UO_1510 (O_1510,N_14838,N_14824);
nor UO_1511 (O_1511,N_14883,N_14816);
nand UO_1512 (O_1512,N_14908,N_14988);
nand UO_1513 (O_1513,N_14842,N_14887);
and UO_1514 (O_1514,N_14930,N_14918);
nor UO_1515 (O_1515,N_14820,N_14930);
or UO_1516 (O_1516,N_14833,N_14841);
and UO_1517 (O_1517,N_14858,N_14988);
xor UO_1518 (O_1518,N_14850,N_14897);
and UO_1519 (O_1519,N_14893,N_14918);
and UO_1520 (O_1520,N_14830,N_14891);
nand UO_1521 (O_1521,N_14967,N_14937);
nand UO_1522 (O_1522,N_14996,N_14841);
nor UO_1523 (O_1523,N_14938,N_14812);
xor UO_1524 (O_1524,N_14900,N_14839);
nand UO_1525 (O_1525,N_14882,N_14948);
nor UO_1526 (O_1526,N_14908,N_14924);
or UO_1527 (O_1527,N_14970,N_14856);
or UO_1528 (O_1528,N_14858,N_14947);
and UO_1529 (O_1529,N_14822,N_14804);
nand UO_1530 (O_1530,N_14913,N_14956);
and UO_1531 (O_1531,N_14927,N_14889);
nand UO_1532 (O_1532,N_14890,N_14830);
or UO_1533 (O_1533,N_14950,N_14872);
or UO_1534 (O_1534,N_14826,N_14902);
nand UO_1535 (O_1535,N_14937,N_14990);
nor UO_1536 (O_1536,N_14868,N_14929);
nor UO_1537 (O_1537,N_14977,N_14832);
nand UO_1538 (O_1538,N_14853,N_14945);
or UO_1539 (O_1539,N_14911,N_14979);
or UO_1540 (O_1540,N_14878,N_14889);
and UO_1541 (O_1541,N_14807,N_14907);
nor UO_1542 (O_1542,N_14861,N_14938);
or UO_1543 (O_1543,N_14999,N_14996);
or UO_1544 (O_1544,N_14978,N_14808);
or UO_1545 (O_1545,N_14965,N_14895);
xnor UO_1546 (O_1546,N_14851,N_14841);
nand UO_1547 (O_1547,N_14809,N_14880);
nand UO_1548 (O_1548,N_14807,N_14925);
and UO_1549 (O_1549,N_14852,N_14959);
nand UO_1550 (O_1550,N_14930,N_14838);
nand UO_1551 (O_1551,N_14921,N_14967);
nor UO_1552 (O_1552,N_14917,N_14913);
and UO_1553 (O_1553,N_14828,N_14894);
xnor UO_1554 (O_1554,N_14964,N_14936);
and UO_1555 (O_1555,N_14906,N_14953);
nor UO_1556 (O_1556,N_14911,N_14973);
or UO_1557 (O_1557,N_14909,N_14805);
nor UO_1558 (O_1558,N_14845,N_14905);
xor UO_1559 (O_1559,N_14816,N_14919);
and UO_1560 (O_1560,N_14803,N_14986);
nor UO_1561 (O_1561,N_14985,N_14935);
xor UO_1562 (O_1562,N_14921,N_14924);
nor UO_1563 (O_1563,N_14958,N_14975);
or UO_1564 (O_1564,N_14811,N_14927);
nor UO_1565 (O_1565,N_14919,N_14820);
nor UO_1566 (O_1566,N_14823,N_14910);
nand UO_1567 (O_1567,N_14977,N_14943);
nand UO_1568 (O_1568,N_14893,N_14979);
nor UO_1569 (O_1569,N_14911,N_14809);
and UO_1570 (O_1570,N_14870,N_14851);
nor UO_1571 (O_1571,N_14873,N_14954);
nand UO_1572 (O_1572,N_14901,N_14898);
or UO_1573 (O_1573,N_14816,N_14852);
nor UO_1574 (O_1574,N_14923,N_14836);
and UO_1575 (O_1575,N_14961,N_14962);
nor UO_1576 (O_1576,N_14902,N_14918);
nor UO_1577 (O_1577,N_14844,N_14839);
and UO_1578 (O_1578,N_14860,N_14826);
xor UO_1579 (O_1579,N_14982,N_14976);
xor UO_1580 (O_1580,N_14834,N_14903);
nor UO_1581 (O_1581,N_14818,N_14887);
and UO_1582 (O_1582,N_14914,N_14961);
or UO_1583 (O_1583,N_14899,N_14942);
nand UO_1584 (O_1584,N_14908,N_14990);
or UO_1585 (O_1585,N_14957,N_14828);
or UO_1586 (O_1586,N_14961,N_14800);
nand UO_1587 (O_1587,N_14905,N_14839);
xnor UO_1588 (O_1588,N_14928,N_14865);
nor UO_1589 (O_1589,N_14884,N_14813);
or UO_1590 (O_1590,N_14862,N_14825);
xor UO_1591 (O_1591,N_14977,N_14819);
and UO_1592 (O_1592,N_14901,N_14994);
and UO_1593 (O_1593,N_14854,N_14975);
or UO_1594 (O_1594,N_14858,N_14892);
nand UO_1595 (O_1595,N_14829,N_14801);
xor UO_1596 (O_1596,N_14936,N_14821);
nor UO_1597 (O_1597,N_14918,N_14938);
nor UO_1598 (O_1598,N_14879,N_14924);
and UO_1599 (O_1599,N_14920,N_14958);
nor UO_1600 (O_1600,N_14849,N_14915);
and UO_1601 (O_1601,N_14978,N_14880);
or UO_1602 (O_1602,N_14986,N_14833);
and UO_1603 (O_1603,N_14912,N_14915);
nor UO_1604 (O_1604,N_14825,N_14956);
nor UO_1605 (O_1605,N_14846,N_14918);
nor UO_1606 (O_1606,N_14980,N_14923);
xor UO_1607 (O_1607,N_14896,N_14862);
xnor UO_1608 (O_1608,N_14856,N_14810);
nand UO_1609 (O_1609,N_14919,N_14992);
xnor UO_1610 (O_1610,N_14912,N_14985);
or UO_1611 (O_1611,N_14866,N_14979);
xnor UO_1612 (O_1612,N_14811,N_14917);
nand UO_1613 (O_1613,N_14953,N_14802);
nand UO_1614 (O_1614,N_14886,N_14887);
or UO_1615 (O_1615,N_14836,N_14877);
nand UO_1616 (O_1616,N_14937,N_14828);
and UO_1617 (O_1617,N_14930,N_14818);
nand UO_1618 (O_1618,N_14853,N_14826);
and UO_1619 (O_1619,N_14884,N_14894);
xor UO_1620 (O_1620,N_14930,N_14942);
or UO_1621 (O_1621,N_14947,N_14906);
or UO_1622 (O_1622,N_14990,N_14945);
or UO_1623 (O_1623,N_14841,N_14987);
or UO_1624 (O_1624,N_14957,N_14857);
and UO_1625 (O_1625,N_14876,N_14897);
xnor UO_1626 (O_1626,N_14985,N_14845);
xnor UO_1627 (O_1627,N_14929,N_14988);
or UO_1628 (O_1628,N_14924,N_14896);
nand UO_1629 (O_1629,N_14955,N_14807);
nor UO_1630 (O_1630,N_14894,N_14814);
nand UO_1631 (O_1631,N_14917,N_14856);
nand UO_1632 (O_1632,N_14817,N_14979);
nor UO_1633 (O_1633,N_14808,N_14897);
nand UO_1634 (O_1634,N_14899,N_14805);
nor UO_1635 (O_1635,N_14992,N_14967);
nand UO_1636 (O_1636,N_14827,N_14800);
and UO_1637 (O_1637,N_14819,N_14959);
and UO_1638 (O_1638,N_14953,N_14843);
nand UO_1639 (O_1639,N_14986,N_14812);
and UO_1640 (O_1640,N_14991,N_14919);
nand UO_1641 (O_1641,N_14913,N_14931);
xnor UO_1642 (O_1642,N_14999,N_14942);
xnor UO_1643 (O_1643,N_14805,N_14801);
and UO_1644 (O_1644,N_14919,N_14899);
nor UO_1645 (O_1645,N_14860,N_14901);
or UO_1646 (O_1646,N_14877,N_14974);
or UO_1647 (O_1647,N_14956,N_14922);
or UO_1648 (O_1648,N_14964,N_14961);
xnor UO_1649 (O_1649,N_14881,N_14945);
nor UO_1650 (O_1650,N_14800,N_14841);
and UO_1651 (O_1651,N_14861,N_14903);
xnor UO_1652 (O_1652,N_14838,N_14812);
xnor UO_1653 (O_1653,N_14820,N_14970);
and UO_1654 (O_1654,N_14891,N_14997);
nor UO_1655 (O_1655,N_14917,N_14885);
and UO_1656 (O_1656,N_14978,N_14884);
nor UO_1657 (O_1657,N_14824,N_14869);
nor UO_1658 (O_1658,N_14876,N_14925);
or UO_1659 (O_1659,N_14949,N_14811);
nand UO_1660 (O_1660,N_14894,N_14819);
and UO_1661 (O_1661,N_14872,N_14941);
or UO_1662 (O_1662,N_14955,N_14888);
and UO_1663 (O_1663,N_14896,N_14991);
nor UO_1664 (O_1664,N_14936,N_14977);
xor UO_1665 (O_1665,N_14935,N_14959);
xnor UO_1666 (O_1666,N_14917,N_14965);
xor UO_1667 (O_1667,N_14874,N_14901);
nand UO_1668 (O_1668,N_14891,N_14833);
and UO_1669 (O_1669,N_14889,N_14956);
and UO_1670 (O_1670,N_14856,N_14854);
and UO_1671 (O_1671,N_14878,N_14917);
and UO_1672 (O_1672,N_14978,N_14945);
xor UO_1673 (O_1673,N_14817,N_14949);
nor UO_1674 (O_1674,N_14869,N_14800);
nor UO_1675 (O_1675,N_14983,N_14856);
nand UO_1676 (O_1676,N_14887,N_14926);
xnor UO_1677 (O_1677,N_14988,N_14913);
nor UO_1678 (O_1678,N_14823,N_14955);
nor UO_1679 (O_1679,N_14855,N_14897);
xnor UO_1680 (O_1680,N_14988,N_14922);
and UO_1681 (O_1681,N_14838,N_14854);
nand UO_1682 (O_1682,N_14824,N_14977);
xor UO_1683 (O_1683,N_14862,N_14895);
or UO_1684 (O_1684,N_14809,N_14975);
and UO_1685 (O_1685,N_14951,N_14928);
xnor UO_1686 (O_1686,N_14931,N_14903);
and UO_1687 (O_1687,N_14932,N_14885);
nand UO_1688 (O_1688,N_14916,N_14968);
nor UO_1689 (O_1689,N_14879,N_14996);
or UO_1690 (O_1690,N_14905,N_14930);
or UO_1691 (O_1691,N_14830,N_14869);
nor UO_1692 (O_1692,N_14985,N_14840);
or UO_1693 (O_1693,N_14891,N_14923);
xnor UO_1694 (O_1694,N_14950,N_14800);
xor UO_1695 (O_1695,N_14986,N_14815);
nand UO_1696 (O_1696,N_14928,N_14840);
xor UO_1697 (O_1697,N_14859,N_14898);
nor UO_1698 (O_1698,N_14984,N_14871);
nor UO_1699 (O_1699,N_14860,N_14925);
or UO_1700 (O_1700,N_14914,N_14870);
nor UO_1701 (O_1701,N_14989,N_14963);
nor UO_1702 (O_1702,N_14855,N_14814);
and UO_1703 (O_1703,N_14928,N_14983);
xor UO_1704 (O_1704,N_14952,N_14965);
or UO_1705 (O_1705,N_14954,N_14998);
and UO_1706 (O_1706,N_14816,N_14826);
nor UO_1707 (O_1707,N_14893,N_14920);
xnor UO_1708 (O_1708,N_14900,N_14820);
or UO_1709 (O_1709,N_14958,N_14834);
xor UO_1710 (O_1710,N_14811,N_14968);
nor UO_1711 (O_1711,N_14983,N_14869);
or UO_1712 (O_1712,N_14893,N_14906);
and UO_1713 (O_1713,N_14937,N_14804);
xnor UO_1714 (O_1714,N_14982,N_14963);
or UO_1715 (O_1715,N_14998,N_14941);
nor UO_1716 (O_1716,N_14811,N_14987);
or UO_1717 (O_1717,N_14899,N_14967);
nor UO_1718 (O_1718,N_14966,N_14802);
or UO_1719 (O_1719,N_14818,N_14995);
nand UO_1720 (O_1720,N_14989,N_14894);
and UO_1721 (O_1721,N_14824,N_14877);
xnor UO_1722 (O_1722,N_14943,N_14818);
and UO_1723 (O_1723,N_14867,N_14902);
xnor UO_1724 (O_1724,N_14885,N_14930);
and UO_1725 (O_1725,N_14811,N_14925);
and UO_1726 (O_1726,N_14892,N_14805);
xor UO_1727 (O_1727,N_14837,N_14989);
nor UO_1728 (O_1728,N_14829,N_14806);
xnor UO_1729 (O_1729,N_14961,N_14972);
nor UO_1730 (O_1730,N_14863,N_14937);
or UO_1731 (O_1731,N_14972,N_14890);
nand UO_1732 (O_1732,N_14823,N_14813);
nor UO_1733 (O_1733,N_14990,N_14953);
nor UO_1734 (O_1734,N_14979,N_14864);
nor UO_1735 (O_1735,N_14993,N_14870);
xnor UO_1736 (O_1736,N_14896,N_14829);
or UO_1737 (O_1737,N_14953,N_14882);
xnor UO_1738 (O_1738,N_14916,N_14929);
xor UO_1739 (O_1739,N_14956,N_14800);
xor UO_1740 (O_1740,N_14966,N_14924);
nand UO_1741 (O_1741,N_14933,N_14866);
nand UO_1742 (O_1742,N_14825,N_14986);
or UO_1743 (O_1743,N_14944,N_14800);
nor UO_1744 (O_1744,N_14879,N_14846);
nand UO_1745 (O_1745,N_14933,N_14828);
nand UO_1746 (O_1746,N_14896,N_14918);
or UO_1747 (O_1747,N_14877,N_14813);
xnor UO_1748 (O_1748,N_14830,N_14825);
or UO_1749 (O_1749,N_14863,N_14918);
xor UO_1750 (O_1750,N_14949,N_14900);
and UO_1751 (O_1751,N_14956,N_14855);
nand UO_1752 (O_1752,N_14819,N_14836);
nand UO_1753 (O_1753,N_14809,N_14998);
xnor UO_1754 (O_1754,N_14804,N_14904);
or UO_1755 (O_1755,N_14986,N_14976);
nor UO_1756 (O_1756,N_14957,N_14984);
nor UO_1757 (O_1757,N_14963,N_14839);
and UO_1758 (O_1758,N_14894,N_14934);
or UO_1759 (O_1759,N_14974,N_14943);
nand UO_1760 (O_1760,N_14844,N_14857);
xnor UO_1761 (O_1761,N_14937,N_14910);
and UO_1762 (O_1762,N_14915,N_14829);
xnor UO_1763 (O_1763,N_14898,N_14824);
nor UO_1764 (O_1764,N_14932,N_14853);
and UO_1765 (O_1765,N_14980,N_14808);
nor UO_1766 (O_1766,N_14942,N_14810);
nor UO_1767 (O_1767,N_14922,N_14923);
and UO_1768 (O_1768,N_14801,N_14953);
xnor UO_1769 (O_1769,N_14950,N_14841);
and UO_1770 (O_1770,N_14869,N_14939);
or UO_1771 (O_1771,N_14894,N_14820);
or UO_1772 (O_1772,N_14904,N_14907);
nand UO_1773 (O_1773,N_14898,N_14960);
nor UO_1774 (O_1774,N_14996,N_14883);
xnor UO_1775 (O_1775,N_14806,N_14931);
nand UO_1776 (O_1776,N_14883,N_14959);
nand UO_1777 (O_1777,N_14847,N_14801);
nand UO_1778 (O_1778,N_14813,N_14864);
or UO_1779 (O_1779,N_14896,N_14801);
nand UO_1780 (O_1780,N_14802,N_14844);
nor UO_1781 (O_1781,N_14981,N_14830);
or UO_1782 (O_1782,N_14864,N_14907);
nor UO_1783 (O_1783,N_14834,N_14916);
nand UO_1784 (O_1784,N_14946,N_14854);
nor UO_1785 (O_1785,N_14966,N_14929);
and UO_1786 (O_1786,N_14986,N_14899);
xnor UO_1787 (O_1787,N_14934,N_14878);
or UO_1788 (O_1788,N_14947,N_14874);
and UO_1789 (O_1789,N_14819,N_14890);
nand UO_1790 (O_1790,N_14978,N_14923);
nor UO_1791 (O_1791,N_14858,N_14921);
nand UO_1792 (O_1792,N_14864,N_14946);
xor UO_1793 (O_1793,N_14881,N_14974);
nor UO_1794 (O_1794,N_14961,N_14898);
nor UO_1795 (O_1795,N_14991,N_14887);
xor UO_1796 (O_1796,N_14822,N_14948);
and UO_1797 (O_1797,N_14876,N_14866);
or UO_1798 (O_1798,N_14932,N_14908);
nor UO_1799 (O_1799,N_14852,N_14824);
and UO_1800 (O_1800,N_14859,N_14981);
or UO_1801 (O_1801,N_14999,N_14949);
nand UO_1802 (O_1802,N_14993,N_14953);
nor UO_1803 (O_1803,N_14977,N_14993);
nor UO_1804 (O_1804,N_14922,N_14924);
nor UO_1805 (O_1805,N_14910,N_14827);
or UO_1806 (O_1806,N_14965,N_14804);
or UO_1807 (O_1807,N_14901,N_14849);
nand UO_1808 (O_1808,N_14918,N_14806);
nor UO_1809 (O_1809,N_14960,N_14884);
or UO_1810 (O_1810,N_14824,N_14832);
nand UO_1811 (O_1811,N_14854,N_14858);
nand UO_1812 (O_1812,N_14829,N_14912);
nand UO_1813 (O_1813,N_14805,N_14915);
or UO_1814 (O_1814,N_14988,N_14937);
nor UO_1815 (O_1815,N_14920,N_14838);
xor UO_1816 (O_1816,N_14820,N_14844);
and UO_1817 (O_1817,N_14809,N_14807);
nand UO_1818 (O_1818,N_14964,N_14935);
xnor UO_1819 (O_1819,N_14852,N_14944);
or UO_1820 (O_1820,N_14826,N_14815);
and UO_1821 (O_1821,N_14953,N_14947);
xnor UO_1822 (O_1822,N_14822,N_14856);
nor UO_1823 (O_1823,N_14940,N_14947);
nor UO_1824 (O_1824,N_14862,N_14912);
nor UO_1825 (O_1825,N_14845,N_14813);
nor UO_1826 (O_1826,N_14883,N_14809);
nand UO_1827 (O_1827,N_14995,N_14894);
and UO_1828 (O_1828,N_14916,N_14935);
nor UO_1829 (O_1829,N_14997,N_14946);
xnor UO_1830 (O_1830,N_14889,N_14955);
and UO_1831 (O_1831,N_14897,N_14806);
and UO_1832 (O_1832,N_14828,N_14993);
nand UO_1833 (O_1833,N_14903,N_14984);
or UO_1834 (O_1834,N_14805,N_14872);
nand UO_1835 (O_1835,N_14913,N_14856);
or UO_1836 (O_1836,N_14953,N_14879);
and UO_1837 (O_1837,N_14817,N_14827);
nor UO_1838 (O_1838,N_14860,N_14914);
and UO_1839 (O_1839,N_14986,N_14979);
nand UO_1840 (O_1840,N_14946,N_14988);
xnor UO_1841 (O_1841,N_14882,N_14937);
xnor UO_1842 (O_1842,N_14804,N_14850);
or UO_1843 (O_1843,N_14873,N_14980);
nand UO_1844 (O_1844,N_14975,N_14989);
nor UO_1845 (O_1845,N_14882,N_14972);
nand UO_1846 (O_1846,N_14848,N_14881);
nor UO_1847 (O_1847,N_14903,N_14987);
nand UO_1848 (O_1848,N_14923,N_14857);
nand UO_1849 (O_1849,N_14824,N_14974);
and UO_1850 (O_1850,N_14922,N_14936);
xor UO_1851 (O_1851,N_14918,N_14995);
nor UO_1852 (O_1852,N_14864,N_14904);
nand UO_1853 (O_1853,N_14806,N_14947);
or UO_1854 (O_1854,N_14851,N_14825);
nand UO_1855 (O_1855,N_14887,N_14918);
and UO_1856 (O_1856,N_14843,N_14845);
nor UO_1857 (O_1857,N_14852,N_14932);
and UO_1858 (O_1858,N_14982,N_14842);
nand UO_1859 (O_1859,N_14946,N_14844);
xnor UO_1860 (O_1860,N_14922,N_14861);
and UO_1861 (O_1861,N_14932,N_14998);
nor UO_1862 (O_1862,N_14982,N_14912);
nor UO_1863 (O_1863,N_14896,N_14871);
and UO_1864 (O_1864,N_14887,N_14932);
and UO_1865 (O_1865,N_14827,N_14912);
nand UO_1866 (O_1866,N_14848,N_14961);
nor UO_1867 (O_1867,N_14874,N_14897);
or UO_1868 (O_1868,N_14868,N_14824);
or UO_1869 (O_1869,N_14820,N_14881);
and UO_1870 (O_1870,N_14810,N_14914);
xnor UO_1871 (O_1871,N_14856,N_14932);
and UO_1872 (O_1872,N_14936,N_14868);
xor UO_1873 (O_1873,N_14957,N_14860);
nor UO_1874 (O_1874,N_14876,N_14903);
xor UO_1875 (O_1875,N_14806,N_14828);
xnor UO_1876 (O_1876,N_14916,N_14805);
nand UO_1877 (O_1877,N_14861,N_14987);
xor UO_1878 (O_1878,N_14993,N_14891);
nand UO_1879 (O_1879,N_14948,N_14998);
and UO_1880 (O_1880,N_14871,N_14944);
and UO_1881 (O_1881,N_14824,N_14900);
xor UO_1882 (O_1882,N_14968,N_14986);
nand UO_1883 (O_1883,N_14984,N_14851);
xor UO_1884 (O_1884,N_14933,N_14839);
nor UO_1885 (O_1885,N_14861,N_14894);
or UO_1886 (O_1886,N_14936,N_14828);
nand UO_1887 (O_1887,N_14820,N_14923);
and UO_1888 (O_1888,N_14834,N_14930);
nand UO_1889 (O_1889,N_14942,N_14982);
nand UO_1890 (O_1890,N_14995,N_14997);
nor UO_1891 (O_1891,N_14850,N_14845);
or UO_1892 (O_1892,N_14802,N_14961);
or UO_1893 (O_1893,N_14817,N_14893);
nand UO_1894 (O_1894,N_14972,N_14944);
nand UO_1895 (O_1895,N_14961,N_14804);
nor UO_1896 (O_1896,N_14914,N_14927);
xor UO_1897 (O_1897,N_14866,N_14912);
nand UO_1898 (O_1898,N_14909,N_14881);
or UO_1899 (O_1899,N_14876,N_14911);
or UO_1900 (O_1900,N_14802,N_14977);
nand UO_1901 (O_1901,N_14989,N_14924);
nand UO_1902 (O_1902,N_14803,N_14916);
nand UO_1903 (O_1903,N_14823,N_14804);
or UO_1904 (O_1904,N_14817,N_14872);
or UO_1905 (O_1905,N_14963,N_14835);
or UO_1906 (O_1906,N_14976,N_14801);
and UO_1907 (O_1907,N_14977,N_14955);
nand UO_1908 (O_1908,N_14853,N_14929);
and UO_1909 (O_1909,N_14966,N_14829);
nor UO_1910 (O_1910,N_14847,N_14910);
or UO_1911 (O_1911,N_14842,N_14914);
nand UO_1912 (O_1912,N_14963,N_14926);
xor UO_1913 (O_1913,N_14909,N_14985);
xor UO_1914 (O_1914,N_14848,N_14986);
or UO_1915 (O_1915,N_14886,N_14800);
xnor UO_1916 (O_1916,N_14956,N_14975);
nand UO_1917 (O_1917,N_14809,N_14879);
nand UO_1918 (O_1918,N_14950,N_14907);
xor UO_1919 (O_1919,N_14928,N_14861);
nand UO_1920 (O_1920,N_14988,N_14931);
xor UO_1921 (O_1921,N_14830,N_14885);
nor UO_1922 (O_1922,N_14899,N_14984);
and UO_1923 (O_1923,N_14879,N_14840);
and UO_1924 (O_1924,N_14868,N_14870);
or UO_1925 (O_1925,N_14910,N_14924);
nor UO_1926 (O_1926,N_14881,N_14953);
and UO_1927 (O_1927,N_14915,N_14809);
or UO_1928 (O_1928,N_14995,N_14807);
or UO_1929 (O_1929,N_14955,N_14982);
nor UO_1930 (O_1930,N_14912,N_14992);
and UO_1931 (O_1931,N_14802,N_14841);
nand UO_1932 (O_1932,N_14983,N_14981);
nor UO_1933 (O_1933,N_14975,N_14976);
or UO_1934 (O_1934,N_14984,N_14800);
or UO_1935 (O_1935,N_14916,N_14946);
or UO_1936 (O_1936,N_14857,N_14893);
and UO_1937 (O_1937,N_14876,N_14939);
or UO_1938 (O_1938,N_14805,N_14860);
nand UO_1939 (O_1939,N_14971,N_14843);
or UO_1940 (O_1940,N_14836,N_14950);
xnor UO_1941 (O_1941,N_14863,N_14828);
and UO_1942 (O_1942,N_14888,N_14806);
xnor UO_1943 (O_1943,N_14801,N_14883);
nor UO_1944 (O_1944,N_14967,N_14909);
xnor UO_1945 (O_1945,N_14864,N_14833);
xor UO_1946 (O_1946,N_14960,N_14862);
and UO_1947 (O_1947,N_14840,N_14924);
or UO_1948 (O_1948,N_14993,N_14808);
nor UO_1949 (O_1949,N_14813,N_14855);
xor UO_1950 (O_1950,N_14995,N_14938);
nand UO_1951 (O_1951,N_14855,N_14863);
or UO_1952 (O_1952,N_14840,N_14809);
nor UO_1953 (O_1953,N_14921,N_14913);
and UO_1954 (O_1954,N_14955,N_14870);
nand UO_1955 (O_1955,N_14933,N_14811);
xnor UO_1956 (O_1956,N_14954,N_14907);
and UO_1957 (O_1957,N_14850,N_14907);
nor UO_1958 (O_1958,N_14862,N_14807);
or UO_1959 (O_1959,N_14811,N_14918);
and UO_1960 (O_1960,N_14844,N_14956);
nor UO_1961 (O_1961,N_14816,N_14857);
nand UO_1962 (O_1962,N_14932,N_14991);
and UO_1963 (O_1963,N_14810,N_14843);
or UO_1964 (O_1964,N_14967,N_14906);
or UO_1965 (O_1965,N_14908,N_14850);
xor UO_1966 (O_1966,N_14871,N_14970);
xor UO_1967 (O_1967,N_14902,N_14915);
and UO_1968 (O_1968,N_14820,N_14886);
and UO_1969 (O_1969,N_14868,N_14913);
nand UO_1970 (O_1970,N_14905,N_14834);
nor UO_1971 (O_1971,N_14884,N_14901);
nand UO_1972 (O_1972,N_14997,N_14844);
nand UO_1973 (O_1973,N_14860,N_14829);
or UO_1974 (O_1974,N_14908,N_14815);
nand UO_1975 (O_1975,N_14807,N_14897);
nor UO_1976 (O_1976,N_14990,N_14891);
or UO_1977 (O_1977,N_14951,N_14875);
and UO_1978 (O_1978,N_14972,N_14832);
or UO_1979 (O_1979,N_14955,N_14876);
xor UO_1980 (O_1980,N_14961,N_14932);
nand UO_1981 (O_1981,N_14805,N_14933);
or UO_1982 (O_1982,N_14978,N_14915);
nand UO_1983 (O_1983,N_14845,N_14844);
or UO_1984 (O_1984,N_14825,N_14833);
nor UO_1985 (O_1985,N_14959,N_14874);
nand UO_1986 (O_1986,N_14933,N_14966);
nand UO_1987 (O_1987,N_14877,N_14883);
nand UO_1988 (O_1988,N_14909,N_14939);
and UO_1989 (O_1989,N_14855,N_14972);
or UO_1990 (O_1990,N_14930,N_14865);
nor UO_1991 (O_1991,N_14997,N_14812);
or UO_1992 (O_1992,N_14973,N_14902);
and UO_1993 (O_1993,N_14978,N_14863);
nor UO_1994 (O_1994,N_14991,N_14947);
and UO_1995 (O_1995,N_14910,N_14876);
or UO_1996 (O_1996,N_14887,N_14901);
or UO_1997 (O_1997,N_14802,N_14806);
or UO_1998 (O_1998,N_14902,N_14929);
xnor UO_1999 (O_1999,N_14803,N_14922);
endmodule