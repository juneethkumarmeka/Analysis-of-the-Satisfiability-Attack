module basic_500_3000_500_30_levels_1xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_123,In_280);
or U1 (N_1,In_93,In_329);
nand U2 (N_2,In_384,In_21);
and U3 (N_3,In_327,In_416);
nor U4 (N_4,In_496,In_288);
nor U5 (N_5,In_170,In_96);
nand U6 (N_6,In_336,In_372);
nor U7 (N_7,In_253,In_197);
and U8 (N_8,In_192,In_162);
nand U9 (N_9,In_465,In_23);
nor U10 (N_10,In_155,In_490);
nand U11 (N_11,In_29,In_491);
or U12 (N_12,In_326,In_273);
xor U13 (N_13,In_11,In_215);
nand U14 (N_14,In_432,In_417);
nor U15 (N_15,In_146,In_359);
and U16 (N_16,In_232,In_3);
or U17 (N_17,In_363,In_430);
and U18 (N_18,In_339,In_173);
nand U19 (N_19,In_221,In_51);
and U20 (N_20,In_191,In_44);
or U21 (N_21,In_394,In_337);
nor U22 (N_22,In_182,In_412);
nor U23 (N_23,In_46,In_18);
and U24 (N_24,In_494,In_189);
and U25 (N_25,In_467,In_345);
nand U26 (N_26,In_214,In_357);
nor U27 (N_27,In_449,In_356);
or U28 (N_28,In_233,In_208);
nand U29 (N_29,In_27,In_84);
or U30 (N_30,In_385,In_87);
or U31 (N_31,In_330,In_53);
and U32 (N_32,In_195,In_309);
or U33 (N_33,In_142,In_2);
or U34 (N_34,In_335,In_271);
xnor U35 (N_35,In_325,In_350);
or U36 (N_36,In_301,In_20);
nor U37 (N_37,In_113,In_145);
nor U38 (N_38,In_386,In_423);
nor U39 (N_39,In_133,In_441);
and U40 (N_40,In_461,In_67);
or U41 (N_41,In_442,In_239);
and U42 (N_42,In_495,In_242);
or U43 (N_43,In_184,In_311);
and U44 (N_44,In_475,In_230);
nand U45 (N_45,In_76,In_315);
nor U46 (N_46,In_167,In_78);
nand U47 (N_47,In_234,In_422);
or U48 (N_48,In_160,In_287);
or U49 (N_49,In_274,In_185);
and U50 (N_50,In_306,In_203);
or U51 (N_51,In_246,In_59);
and U52 (N_52,In_199,In_318);
and U53 (N_53,In_131,In_135);
nand U54 (N_54,In_60,In_171);
nor U55 (N_55,In_138,In_437);
nand U56 (N_56,In_209,In_291);
and U57 (N_57,In_499,In_341);
nand U58 (N_58,In_344,In_360);
and U59 (N_59,In_174,In_43);
nor U60 (N_60,In_56,In_383);
or U61 (N_61,In_440,In_117);
or U62 (N_62,In_408,In_397);
and U63 (N_63,In_438,In_85);
and U64 (N_64,In_127,In_295);
or U65 (N_65,In_57,In_211);
or U66 (N_66,In_16,In_451);
nor U67 (N_67,In_71,In_258);
nor U68 (N_68,In_260,In_433);
or U69 (N_69,In_130,In_453);
or U70 (N_70,In_388,In_139);
nor U71 (N_71,In_459,In_460);
nor U72 (N_72,In_498,In_338);
or U73 (N_73,In_47,In_143);
or U74 (N_74,In_126,In_163);
or U75 (N_75,In_452,In_282);
or U76 (N_76,In_390,In_122);
or U77 (N_77,In_104,In_366);
or U78 (N_78,In_1,In_275);
and U79 (N_79,In_148,In_41);
or U80 (N_80,In_375,In_92);
nor U81 (N_81,In_5,In_198);
nor U82 (N_82,In_448,In_89);
and U83 (N_83,In_88,In_103);
or U84 (N_84,In_264,In_395);
and U85 (N_85,In_314,In_472);
nor U86 (N_86,In_178,In_4);
xnor U87 (N_87,In_302,In_231);
and U88 (N_88,In_420,In_63);
nor U89 (N_89,In_458,In_70);
or U90 (N_90,In_293,In_358);
nand U91 (N_91,In_129,In_187);
nand U92 (N_92,In_79,In_400);
nand U93 (N_93,In_474,In_380);
nor U94 (N_94,In_477,In_201);
or U95 (N_95,In_106,In_473);
or U96 (N_96,In_66,In_493);
or U97 (N_97,In_176,In_166);
nand U98 (N_98,In_277,In_444);
or U99 (N_99,In_310,In_406);
or U100 (N_100,In_333,In_379);
nand U101 (N_101,In_118,In_31);
or U102 (N_102,N_52,N_32);
nand U103 (N_103,N_34,In_405);
and U104 (N_104,In_352,In_402);
nor U105 (N_105,N_33,In_265);
nor U106 (N_106,N_76,N_38);
nand U107 (N_107,In_398,N_59);
and U108 (N_108,In_48,In_393);
or U109 (N_109,N_99,In_238);
nor U110 (N_110,In_248,In_7);
nor U111 (N_111,In_81,In_382);
nor U112 (N_112,In_252,In_164);
and U113 (N_113,In_147,N_24);
or U114 (N_114,In_153,N_14);
nand U115 (N_115,N_41,In_488);
nor U116 (N_116,In_37,In_200);
and U117 (N_117,In_454,In_290);
or U118 (N_118,In_346,In_140);
or U119 (N_119,N_70,N_25);
and U120 (N_120,In_245,N_7);
nor U121 (N_121,In_367,In_342);
or U122 (N_122,N_37,In_466);
and U123 (N_123,In_55,N_86);
or U124 (N_124,In_308,N_43);
and U125 (N_125,In_125,In_447);
nand U126 (N_126,In_332,In_156);
or U127 (N_127,In_255,In_285);
or U128 (N_128,In_268,In_36);
and U129 (N_129,N_36,In_168);
nand U130 (N_130,In_387,N_21);
or U131 (N_131,In_183,In_431);
xnor U132 (N_132,In_128,N_80);
nand U133 (N_133,In_38,In_377);
or U134 (N_134,In_241,N_87);
nor U135 (N_135,In_223,N_61);
nor U136 (N_136,In_227,In_476);
and U137 (N_137,In_415,In_492);
or U138 (N_138,In_483,In_58);
or U139 (N_139,N_82,In_105);
nor U140 (N_140,N_1,In_124);
nor U141 (N_141,In_108,In_312);
xnor U142 (N_142,In_80,N_53);
and U143 (N_143,N_69,In_334);
nor U144 (N_144,In_13,In_361);
nor U145 (N_145,In_40,In_267);
nand U146 (N_146,N_97,N_74);
nor U147 (N_147,In_300,In_299);
nand U148 (N_148,In_369,N_62);
nor U149 (N_149,In_455,In_62);
and U150 (N_150,In_292,In_100);
and U151 (N_151,In_74,N_77);
nand U152 (N_152,In_481,In_355);
nor U153 (N_153,N_18,In_77);
and U154 (N_154,In_73,In_217);
and U155 (N_155,In_487,In_463);
nor U156 (N_156,In_82,In_364);
or U157 (N_157,In_10,In_95);
and U158 (N_158,In_320,In_194);
nand U159 (N_159,In_206,N_92);
nor U160 (N_160,In_303,N_8);
nor U161 (N_161,In_436,In_204);
or U162 (N_162,In_159,In_322);
nor U163 (N_163,In_428,N_98);
nand U164 (N_164,N_54,N_27);
and U165 (N_165,In_278,N_95);
nand U166 (N_166,In_179,In_317);
and U167 (N_167,N_63,In_497);
or U168 (N_168,In_484,In_224);
and U169 (N_169,In_137,N_45);
or U170 (N_170,In_33,N_19);
and U171 (N_171,N_22,N_35);
nand U172 (N_172,In_279,In_257);
nor U173 (N_173,N_81,In_216);
xnor U174 (N_174,In_281,In_32);
or U175 (N_175,N_93,In_354);
and U176 (N_176,In_482,In_353);
xnor U177 (N_177,In_426,In_45);
and U178 (N_178,In_266,In_376);
or U179 (N_179,In_110,In_237);
nand U180 (N_180,In_434,N_58);
and U181 (N_181,In_17,In_323);
and U182 (N_182,In_172,N_91);
or U183 (N_183,N_51,In_429);
and U184 (N_184,In_6,In_119);
or U185 (N_185,In_262,In_362);
or U186 (N_186,N_26,In_371);
and U187 (N_187,In_349,In_331);
nand U188 (N_188,In_283,N_73);
or U189 (N_189,In_413,In_435);
nand U190 (N_190,In_39,In_403);
nor U191 (N_191,In_114,In_480);
nor U192 (N_192,In_324,N_68);
nand U193 (N_193,In_165,In_389);
nor U194 (N_194,In_343,In_263);
or U195 (N_195,In_478,In_69);
or U196 (N_196,N_4,In_236);
or U197 (N_197,In_83,In_181);
or U198 (N_198,In_348,N_12);
nand U199 (N_199,In_180,In_276);
and U200 (N_200,In_425,N_42);
nor U201 (N_201,In_90,In_97);
nand U202 (N_202,In_418,N_55);
nand U203 (N_203,N_194,In_22);
and U204 (N_204,In_414,N_169);
nand U205 (N_205,In_469,In_154);
xor U206 (N_206,In_25,In_298);
nor U207 (N_207,In_404,In_294);
and U208 (N_208,N_168,N_153);
nand U209 (N_209,N_176,N_142);
or U210 (N_210,N_196,In_190);
and U211 (N_211,In_392,In_24);
nor U212 (N_212,N_132,In_101);
nand U213 (N_213,N_119,In_297);
nand U214 (N_214,In_340,In_107);
nand U215 (N_215,N_181,In_289);
nor U216 (N_216,In_411,In_243);
or U217 (N_217,N_50,In_235);
nor U218 (N_218,In_468,In_35);
or U219 (N_219,In_479,N_118);
nor U220 (N_220,In_109,N_171);
nand U221 (N_221,In_254,N_154);
nand U222 (N_222,In_112,N_151);
nor U223 (N_223,In_446,In_284);
and U224 (N_224,In_188,N_163);
nor U225 (N_225,N_23,N_170);
nor U226 (N_226,N_110,In_196);
and U227 (N_227,In_419,N_39);
nor U228 (N_228,N_109,In_319);
and U229 (N_229,N_100,N_120);
nand U230 (N_230,In_116,In_244);
nand U231 (N_231,N_10,N_195);
nor U232 (N_232,In_229,N_65);
nand U233 (N_233,In_65,In_439);
or U234 (N_234,N_79,In_205);
and U235 (N_235,N_64,N_0);
nand U236 (N_236,In_175,In_373);
or U237 (N_237,In_307,N_164);
and U238 (N_238,N_130,N_133);
and U239 (N_239,N_159,In_136);
or U240 (N_240,N_75,N_106);
and U241 (N_241,N_139,N_141);
nor U242 (N_242,N_67,N_11);
nor U243 (N_243,In_132,N_13);
or U244 (N_244,In_249,N_192);
or U245 (N_245,N_5,N_29);
nor U246 (N_246,In_157,In_251);
and U247 (N_247,N_197,In_49);
nand U248 (N_248,In_489,In_94);
nor U249 (N_249,N_15,N_47);
nor U250 (N_250,N_78,In_218);
or U251 (N_251,N_174,In_226);
or U252 (N_252,N_112,N_150);
nand U253 (N_253,N_162,In_378);
nor U254 (N_254,N_175,In_259);
nor U255 (N_255,N_193,N_85);
nor U256 (N_256,In_261,N_188);
nor U257 (N_257,N_137,In_250);
or U258 (N_258,N_147,In_391);
nand U259 (N_259,N_185,In_61);
or U260 (N_260,N_105,In_99);
nor U261 (N_261,In_91,N_126);
or U262 (N_262,N_161,In_381);
nor U263 (N_263,N_155,N_122);
nand U264 (N_264,N_9,N_104);
nand U265 (N_265,N_66,N_186);
nor U266 (N_266,N_89,N_44);
nor U267 (N_267,N_3,In_54);
nor U268 (N_268,In_68,In_328);
nor U269 (N_269,N_72,In_485);
or U270 (N_270,In_410,N_128);
nand U271 (N_271,In_401,In_50);
nor U272 (N_272,N_28,In_286);
or U273 (N_273,In_72,In_213);
and U274 (N_274,In_150,N_17);
and U275 (N_275,In_470,In_409);
nor U276 (N_276,N_125,In_151);
and U277 (N_277,N_40,In_269);
nor U278 (N_278,N_180,N_143);
and U279 (N_279,N_179,N_116);
nor U280 (N_280,In_0,N_16);
or U281 (N_281,In_296,N_145);
nor U282 (N_282,In_149,In_427);
nor U283 (N_283,N_184,N_30);
nand U284 (N_284,N_148,In_365);
or U285 (N_285,In_186,N_6);
or U286 (N_286,In_34,N_107);
and U287 (N_287,In_445,In_210);
nand U288 (N_288,In_8,In_202);
nor U289 (N_289,N_101,In_222);
or U290 (N_290,N_46,In_26);
and U291 (N_291,In_321,N_108);
and U292 (N_292,In_30,N_71);
and U293 (N_293,In_225,N_20);
nor U294 (N_294,N_102,N_88);
nand U295 (N_295,N_199,N_113);
or U296 (N_296,N_152,In_111);
and U297 (N_297,In_368,N_129);
nand U298 (N_298,N_187,In_86);
nand U299 (N_299,In_456,N_198);
and U300 (N_300,N_262,N_265);
or U301 (N_301,N_215,N_56);
nand U302 (N_302,N_298,N_253);
or U303 (N_303,In_12,In_14);
nor U304 (N_304,In_270,N_124);
and U305 (N_305,N_138,N_260);
nor U306 (N_306,N_299,N_227);
nor U307 (N_307,N_271,N_208);
nor U308 (N_308,In_313,N_203);
or U309 (N_309,N_252,N_231);
nand U310 (N_310,N_140,In_407);
and U311 (N_311,N_280,N_177);
and U312 (N_312,In_9,N_156);
nand U313 (N_313,N_48,In_161);
nand U314 (N_314,In_399,N_228);
or U315 (N_315,N_272,N_31);
nand U316 (N_316,N_189,In_134);
nor U317 (N_317,In_443,N_294);
nand U318 (N_318,In_421,N_229);
nand U319 (N_319,In_374,In_240);
nor U320 (N_320,In_457,In_220);
nand U321 (N_321,In_486,N_247);
nand U322 (N_322,N_284,N_269);
nand U323 (N_323,N_166,N_244);
and U324 (N_324,N_274,N_165);
nand U325 (N_325,N_144,N_259);
nor U326 (N_326,N_240,In_193);
nor U327 (N_327,N_266,N_264);
nor U328 (N_328,N_182,N_202);
nand U329 (N_329,N_209,N_158);
nand U330 (N_330,N_277,N_117);
nand U331 (N_331,N_246,In_64);
nor U332 (N_332,In_396,N_257);
nor U333 (N_333,N_273,N_217);
nor U334 (N_334,In_75,N_251);
and U335 (N_335,In_471,In_424);
and U336 (N_336,N_210,N_218);
nand U337 (N_337,N_254,In_158);
and U338 (N_338,N_127,N_183);
nand U339 (N_339,N_238,N_49);
or U340 (N_340,N_289,In_272);
xor U341 (N_341,In_228,In_169);
and U342 (N_342,N_256,In_28);
and U343 (N_343,In_207,N_224);
and U344 (N_344,N_296,N_222);
and U345 (N_345,N_114,N_236);
or U346 (N_346,N_221,N_57);
nor U347 (N_347,N_239,In_305);
or U348 (N_348,N_167,N_206);
nand U349 (N_349,N_103,N_258);
or U350 (N_350,N_241,N_207);
and U351 (N_351,N_232,N_245);
and U352 (N_352,In_351,N_263);
and U353 (N_353,In_15,N_235);
xor U354 (N_354,N_111,In_19);
or U355 (N_355,N_94,N_157);
nor U356 (N_356,N_205,N_276);
or U357 (N_357,In_115,N_226);
nand U358 (N_358,N_60,N_290);
nor U359 (N_359,N_297,N_115);
nor U360 (N_360,N_295,N_204);
or U361 (N_361,In_42,In_256);
nand U362 (N_362,In_247,N_243);
and U363 (N_363,N_237,N_131);
and U364 (N_364,N_286,N_83);
nor U365 (N_365,N_250,N_134);
nand U366 (N_366,N_214,In_464);
nand U367 (N_367,N_255,N_190);
or U368 (N_368,N_136,N_220);
and U369 (N_369,N_292,N_200);
and U370 (N_370,In_347,In_120);
nand U371 (N_371,N_212,N_275);
and U372 (N_372,N_283,In_212);
and U373 (N_373,In_152,N_248);
and U374 (N_374,N_293,N_149);
and U375 (N_375,N_211,N_287);
nand U376 (N_376,In_219,In_141);
nand U377 (N_377,N_201,N_291);
or U378 (N_378,In_462,N_121);
nor U379 (N_379,In_98,N_279);
nor U380 (N_380,N_230,In_304);
and U381 (N_381,In_121,In_177);
nand U382 (N_382,N_135,N_285);
nor U383 (N_383,N_223,N_191);
and U384 (N_384,N_261,N_216);
or U385 (N_385,N_282,N_173);
and U386 (N_386,N_219,N_2);
and U387 (N_387,In_52,N_96);
and U388 (N_388,N_84,N_213);
or U389 (N_389,In_144,N_267);
nor U390 (N_390,In_102,N_178);
or U391 (N_391,N_281,N_146);
nor U392 (N_392,N_268,N_288);
nand U393 (N_393,N_233,N_160);
and U394 (N_394,N_225,N_172);
or U395 (N_395,In_316,In_450);
or U396 (N_396,N_234,N_270);
nand U397 (N_397,N_90,N_123);
nor U398 (N_398,In_370,N_249);
or U399 (N_399,N_278,N_242);
nand U400 (N_400,N_367,N_324);
and U401 (N_401,N_346,N_343);
or U402 (N_402,N_308,N_335);
and U403 (N_403,N_326,N_301);
or U404 (N_404,N_336,N_358);
and U405 (N_405,N_386,N_322);
nor U406 (N_406,N_319,N_376);
nor U407 (N_407,N_398,N_368);
nor U408 (N_408,N_300,N_330);
or U409 (N_409,N_369,N_381);
and U410 (N_410,N_312,N_375);
nand U411 (N_411,N_366,N_378);
and U412 (N_412,N_341,N_362);
nor U413 (N_413,N_342,N_339);
or U414 (N_414,N_349,N_327);
and U415 (N_415,N_390,N_313);
nand U416 (N_416,N_302,N_389);
nor U417 (N_417,N_393,N_354);
or U418 (N_418,N_310,N_334);
nand U419 (N_419,N_303,N_328);
nand U420 (N_420,N_352,N_387);
nand U421 (N_421,N_304,N_379);
and U422 (N_422,N_384,N_355);
or U423 (N_423,N_314,N_382);
and U424 (N_424,N_338,N_329);
and U425 (N_425,N_332,N_394);
nor U426 (N_426,N_325,N_385);
or U427 (N_427,N_315,N_388);
and U428 (N_428,N_320,N_370);
and U429 (N_429,N_323,N_305);
nor U430 (N_430,N_331,N_356);
nand U431 (N_431,N_377,N_371);
nor U432 (N_432,N_374,N_306);
nand U433 (N_433,N_360,N_372);
and U434 (N_434,N_359,N_392);
or U435 (N_435,N_307,N_373);
and U436 (N_436,N_395,N_345);
nand U437 (N_437,N_316,N_357);
nand U438 (N_438,N_383,N_318);
nor U439 (N_439,N_311,N_361);
nand U440 (N_440,N_397,N_350);
nand U441 (N_441,N_364,N_340);
nor U442 (N_442,N_396,N_353);
or U443 (N_443,N_365,N_309);
nand U444 (N_444,N_348,N_347);
or U445 (N_445,N_399,N_380);
nand U446 (N_446,N_337,N_321);
nand U447 (N_447,N_363,N_317);
or U448 (N_448,N_391,N_344);
or U449 (N_449,N_351,N_333);
nand U450 (N_450,N_395,N_367);
xnor U451 (N_451,N_330,N_362);
nor U452 (N_452,N_322,N_393);
nor U453 (N_453,N_348,N_334);
and U454 (N_454,N_318,N_356);
nor U455 (N_455,N_345,N_393);
and U456 (N_456,N_362,N_333);
and U457 (N_457,N_310,N_337);
and U458 (N_458,N_365,N_302);
nor U459 (N_459,N_306,N_311);
and U460 (N_460,N_384,N_307);
or U461 (N_461,N_367,N_317);
nor U462 (N_462,N_370,N_348);
and U463 (N_463,N_305,N_315);
nand U464 (N_464,N_300,N_317);
or U465 (N_465,N_335,N_397);
and U466 (N_466,N_390,N_394);
nand U467 (N_467,N_335,N_358);
nand U468 (N_468,N_359,N_386);
or U469 (N_469,N_302,N_384);
nand U470 (N_470,N_378,N_306);
and U471 (N_471,N_347,N_374);
and U472 (N_472,N_391,N_305);
or U473 (N_473,N_363,N_324);
or U474 (N_474,N_314,N_319);
nand U475 (N_475,N_331,N_341);
nand U476 (N_476,N_342,N_393);
nor U477 (N_477,N_374,N_386);
or U478 (N_478,N_341,N_322);
nor U479 (N_479,N_382,N_373);
nor U480 (N_480,N_338,N_371);
or U481 (N_481,N_343,N_304);
nand U482 (N_482,N_366,N_396);
nand U483 (N_483,N_309,N_351);
xor U484 (N_484,N_345,N_338);
nand U485 (N_485,N_333,N_344);
and U486 (N_486,N_386,N_372);
nor U487 (N_487,N_343,N_313);
nand U488 (N_488,N_399,N_303);
or U489 (N_489,N_349,N_387);
nor U490 (N_490,N_314,N_379);
or U491 (N_491,N_364,N_300);
and U492 (N_492,N_364,N_376);
nor U493 (N_493,N_365,N_371);
nor U494 (N_494,N_344,N_325);
or U495 (N_495,N_386,N_363);
or U496 (N_496,N_350,N_347);
or U497 (N_497,N_316,N_390);
nand U498 (N_498,N_355,N_332);
or U499 (N_499,N_326,N_310);
nand U500 (N_500,N_422,N_487);
nand U501 (N_501,N_405,N_431);
or U502 (N_502,N_401,N_410);
or U503 (N_503,N_406,N_420);
or U504 (N_504,N_433,N_428);
or U505 (N_505,N_400,N_455);
nand U506 (N_506,N_463,N_438);
xor U507 (N_507,N_423,N_489);
nand U508 (N_508,N_496,N_478);
nand U509 (N_509,N_464,N_453);
nand U510 (N_510,N_414,N_408);
nor U511 (N_511,N_475,N_403);
nor U512 (N_512,N_418,N_454);
nand U513 (N_513,N_426,N_415);
nor U514 (N_514,N_411,N_476);
or U515 (N_515,N_457,N_473);
and U516 (N_516,N_448,N_485);
nor U517 (N_517,N_446,N_467);
nand U518 (N_518,N_439,N_481);
or U519 (N_519,N_429,N_409);
and U520 (N_520,N_440,N_459);
and U521 (N_521,N_425,N_483);
nor U522 (N_522,N_421,N_465);
or U523 (N_523,N_416,N_437);
nor U524 (N_524,N_436,N_460);
and U525 (N_525,N_486,N_469);
and U526 (N_526,N_461,N_468);
and U527 (N_527,N_484,N_443);
nor U528 (N_528,N_471,N_492);
or U529 (N_529,N_434,N_449);
and U530 (N_530,N_402,N_407);
nand U531 (N_531,N_477,N_490);
nand U532 (N_532,N_430,N_419);
or U533 (N_533,N_488,N_444);
nor U534 (N_534,N_470,N_452);
nor U535 (N_535,N_451,N_447);
nand U536 (N_536,N_479,N_491);
nand U537 (N_537,N_404,N_442);
or U538 (N_538,N_494,N_499);
nor U539 (N_539,N_435,N_466);
and U540 (N_540,N_480,N_482);
or U541 (N_541,N_497,N_472);
and U542 (N_542,N_427,N_495);
nand U543 (N_543,N_462,N_413);
nor U544 (N_544,N_456,N_412);
nor U545 (N_545,N_445,N_450);
nand U546 (N_546,N_417,N_432);
nor U547 (N_547,N_474,N_498);
nand U548 (N_548,N_424,N_458);
nor U549 (N_549,N_441,N_493);
or U550 (N_550,N_498,N_454);
nor U551 (N_551,N_474,N_452);
nor U552 (N_552,N_412,N_478);
and U553 (N_553,N_432,N_461);
and U554 (N_554,N_424,N_485);
nand U555 (N_555,N_425,N_466);
or U556 (N_556,N_487,N_418);
nand U557 (N_557,N_461,N_497);
or U558 (N_558,N_419,N_485);
or U559 (N_559,N_481,N_437);
xnor U560 (N_560,N_479,N_403);
and U561 (N_561,N_450,N_462);
and U562 (N_562,N_446,N_491);
nand U563 (N_563,N_492,N_443);
and U564 (N_564,N_457,N_407);
nand U565 (N_565,N_449,N_464);
nor U566 (N_566,N_430,N_422);
nor U567 (N_567,N_427,N_487);
or U568 (N_568,N_477,N_496);
nand U569 (N_569,N_441,N_474);
or U570 (N_570,N_484,N_452);
nand U571 (N_571,N_471,N_469);
or U572 (N_572,N_411,N_416);
and U573 (N_573,N_495,N_479);
nor U574 (N_574,N_435,N_457);
nand U575 (N_575,N_484,N_445);
and U576 (N_576,N_453,N_462);
and U577 (N_577,N_440,N_474);
nand U578 (N_578,N_436,N_448);
nor U579 (N_579,N_499,N_414);
or U580 (N_580,N_490,N_449);
nand U581 (N_581,N_478,N_427);
and U582 (N_582,N_493,N_431);
nor U583 (N_583,N_423,N_498);
nor U584 (N_584,N_474,N_445);
nor U585 (N_585,N_487,N_462);
and U586 (N_586,N_486,N_416);
and U587 (N_587,N_458,N_483);
nand U588 (N_588,N_499,N_438);
and U589 (N_589,N_463,N_477);
or U590 (N_590,N_418,N_406);
nor U591 (N_591,N_403,N_413);
nand U592 (N_592,N_448,N_408);
or U593 (N_593,N_442,N_402);
or U594 (N_594,N_497,N_469);
nand U595 (N_595,N_452,N_447);
nor U596 (N_596,N_400,N_489);
or U597 (N_597,N_417,N_486);
nor U598 (N_598,N_444,N_449);
or U599 (N_599,N_449,N_422);
and U600 (N_600,N_576,N_572);
and U601 (N_601,N_546,N_525);
and U602 (N_602,N_555,N_539);
or U603 (N_603,N_573,N_533);
nand U604 (N_604,N_591,N_550);
and U605 (N_605,N_592,N_540);
or U606 (N_606,N_562,N_547);
nand U607 (N_607,N_597,N_569);
nor U608 (N_608,N_508,N_524);
or U609 (N_609,N_589,N_537);
nand U610 (N_610,N_544,N_521);
or U611 (N_611,N_581,N_574);
and U612 (N_612,N_568,N_541);
or U613 (N_613,N_575,N_536);
or U614 (N_614,N_580,N_507);
nand U615 (N_615,N_560,N_523);
nand U616 (N_616,N_528,N_558);
nor U617 (N_617,N_512,N_509);
or U618 (N_618,N_584,N_516);
and U619 (N_619,N_513,N_566);
or U620 (N_620,N_594,N_511);
nand U621 (N_621,N_595,N_593);
nand U622 (N_622,N_563,N_518);
or U623 (N_623,N_510,N_543);
nor U624 (N_624,N_531,N_517);
and U625 (N_625,N_545,N_538);
nand U626 (N_626,N_514,N_557);
nor U627 (N_627,N_503,N_582);
nand U628 (N_628,N_583,N_542);
nand U629 (N_629,N_578,N_588);
nor U630 (N_630,N_552,N_548);
nor U631 (N_631,N_579,N_504);
nand U632 (N_632,N_519,N_553);
nand U633 (N_633,N_586,N_534);
or U634 (N_634,N_501,N_500);
and U635 (N_635,N_564,N_515);
and U636 (N_636,N_526,N_520);
nor U637 (N_637,N_598,N_530);
nor U638 (N_638,N_590,N_532);
nand U639 (N_639,N_551,N_559);
nand U640 (N_640,N_506,N_599);
nor U641 (N_641,N_549,N_561);
nor U642 (N_642,N_567,N_585);
and U643 (N_643,N_529,N_565);
and U644 (N_644,N_505,N_554);
or U645 (N_645,N_596,N_522);
and U646 (N_646,N_502,N_571);
or U647 (N_647,N_556,N_527);
nand U648 (N_648,N_535,N_577);
or U649 (N_649,N_570,N_587);
and U650 (N_650,N_501,N_518);
and U651 (N_651,N_554,N_510);
nand U652 (N_652,N_534,N_599);
and U653 (N_653,N_572,N_533);
or U654 (N_654,N_571,N_575);
or U655 (N_655,N_549,N_531);
and U656 (N_656,N_560,N_588);
nand U657 (N_657,N_511,N_508);
nand U658 (N_658,N_507,N_544);
nor U659 (N_659,N_594,N_591);
nand U660 (N_660,N_588,N_512);
or U661 (N_661,N_533,N_550);
nor U662 (N_662,N_575,N_538);
and U663 (N_663,N_599,N_573);
or U664 (N_664,N_581,N_564);
nor U665 (N_665,N_513,N_563);
or U666 (N_666,N_527,N_576);
and U667 (N_667,N_574,N_508);
or U668 (N_668,N_520,N_518);
and U669 (N_669,N_582,N_588);
or U670 (N_670,N_585,N_557);
and U671 (N_671,N_574,N_547);
or U672 (N_672,N_517,N_553);
or U673 (N_673,N_569,N_521);
nor U674 (N_674,N_502,N_501);
nor U675 (N_675,N_577,N_541);
and U676 (N_676,N_539,N_552);
and U677 (N_677,N_567,N_568);
nand U678 (N_678,N_573,N_530);
and U679 (N_679,N_556,N_503);
or U680 (N_680,N_502,N_504);
and U681 (N_681,N_535,N_512);
or U682 (N_682,N_502,N_587);
or U683 (N_683,N_537,N_541);
or U684 (N_684,N_589,N_521);
nand U685 (N_685,N_593,N_546);
nor U686 (N_686,N_555,N_554);
and U687 (N_687,N_560,N_568);
and U688 (N_688,N_595,N_581);
xor U689 (N_689,N_553,N_511);
nor U690 (N_690,N_514,N_526);
nor U691 (N_691,N_517,N_596);
nor U692 (N_692,N_562,N_567);
and U693 (N_693,N_570,N_565);
nor U694 (N_694,N_569,N_517);
and U695 (N_695,N_542,N_527);
or U696 (N_696,N_553,N_552);
nand U697 (N_697,N_532,N_566);
nor U698 (N_698,N_511,N_565);
nand U699 (N_699,N_573,N_539);
and U700 (N_700,N_677,N_647);
nand U701 (N_701,N_644,N_621);
or U702 (N_702,N_678,N_641);
nand U703 (N_703,N_608,N_606);
nand U704 (N_704,N_661,N_642);
or U705 (N_705,N_638,N_663);
nor U706 (N_706,N_626,N_658);
nand U707 (N_707,N_696,N_679);
or U708 (N_708,N_698,N_690);
nor U709 (N_709,N_654,N_657);
nor U710 (N_710,N_664,N_695);
nor U711 (N_711,N_692,N_610);
and U712 (N_712,N_650,N_612);
or U713 (N_713,N_633,N_659);
or U714 (N_714,N_613,N_660);
or U715 (N_715,N_699,N_646);
nand U716 (N_716,N_671,N_601);
and U717 (N_717,N_645,N_685);
and U718 (N_718,N_652,N_649);
nand U719 (N_719,N_609,N_617);
or U720 (N_720,N_635,N_682);
nor U721 (N_721,N_683,N_623);
and U722 (N_722,N_668,N_605);
and U723 (N_723,N_672,N_628);
and U724 (N_724,N_607,N_630);
or U725 (N_725,N_656,N_600);
nand U726 (N_726,N_670,N_653);
nor U727 (N_727,N_643,N_639);
or U728 (N_728,N_674,N_624);
and U729 (N_729,N_603,N_693);
nor U730 (N_730,N_634,N_619);
nand U731 (N_731,N_620,N_629);
nand U732 (N_732,N_680,N_627);
or U733 (N_733,N_684,N_681);
and U734 (N_734,N_662,N_694);
nand U735 (N_735,N_614,N_697);
nand U736 (N_736,N_636,N_675);
and U737 (N_737,N_689,N_632);
nand U738 (N_738,N_687,N_640);
nor U739 (N_739,N_618,N_666);
nand U740 (N_740,N_648,N_615);
and U741 (N_741,N_625,N_616);
or U742 (N_742,N_655,N_676);
or U743 (N_743,N_602,N_604);
nand U744 (N_744,N_631,N_637);
and U745 (N_745,N_667,N_611);
nand U746 (N_746,N_688,N_691);
nand U747 (N_747,N_622,N_673);
nand U748 (N_748,N_651,N_686);
and U749 (N_749,N_665,N_669);
nand U750 (N_750,N_639,N_666);
or U751 (N_751,N_646,N_622);
nand U752 (N_752,N_695,N_606);
or U753 (N_753,N_680,N_645);
or U754 (N_754,N_667,N_616);
and U755 (N_755,N_679,N_645);
nand U756 (N_756,N_605,N_695);
nand U757 (N_757,N_674,N_629);
or U758 (N_758,N_689,N_661);
nor U759 (N_759,N_613,N_642);
and U760 (N_760,N_670,N_629);
and U761 (N_761,N_673,N_635);
or U762 (N_762,N_683,N_696);
and U763 (N_763,N_640,N_671);
or U764 (N_764,N_676,N_603);
or U765 (N_765,N_628,N_601);
nor U766 (N_766,N_609,N_610);
and U767 (N_767,N_641,N_606);
nor U768 (N_768,N_685,N_663);
or U769 (N_769,N_635,N_698);
and U770 (N_770,N_686,N_613);
nor U771 (N_771,N_618,N_616);
and U772 (N_772,N_674,N_631);
nand U773 (N_773,N_658,N_622);
nor U774 (N_774,N_673,N_697);
nor U775 (N_775,N_626,N_624);
or U776 (N_776,N_687,N_659);
or U777 (N_777,N_656,N_640);
nor U778 (N_778,N_647,N_646);
nor U779 (N_779,N_656,N_677);
nand U780 (N_780,N_695,N_639);
nand U781 (N_781,N_653,N_613);
nand U782 (N_782,N_639,N_690);
and U783 (N_783,N_605,N_649);
nand U784 (N_784,N_607,N_690);
or U785 (N_785,N_671,N_674);
and U786 (N_786,N_649,N_687);
nand U787 (N_787,N_605,N_614);
nand U788 (N_788,N_610,N_615);
nor U789 (N_789,N_649,N_680);
nor U790 (N_790,N_684,N_665);
and U791 (N_791,N_629,N_628);
or U792 (N_792,N_663,N_606);
and U793 (N_793,N_645,N_697);
or U794 (N_794,N_607,N_615);
or U795 (N_795,N_654,N_665);
nor U796 (N_796,N_603,N_649);
or U797 (N_797,N_690,N_623);
and U798 (N_798,N_627,N_662);
nor U799 (N_799,N_674,N_681);
or U800 (N_800,N_770,N_795);
nor U801 (N_801,N_778,N_760);
and U802 (N_802,N_796,N_718);
nand U803 (N_803,N_713,N_752);
and U804 (N_804,N_777,N_774);
nand U805 (N_805,N_734,N_705);
and U806 (N_806,N_726,N_746);
or U807 (N_807,N_712,N_716);
and U808 (N_808,N_749,N_724);
nand U809 (N_809,N_769,N_761);
or U810 (N_810,N_754,N_727);
nor U811 (N_811,N_725,N_775);
and U812 (N_812,N_700,N_717);
nor U813 (N_813,N_737,N_745);
xnor U814 (N_814,N_767,N_787);
nor U815 (N_815,N_758,N_783);
nor U816 (N_816,N_711,N_728);
nand U817 (N_817,N_715,N_750);
nor U818 (N_818,N_784,N_731);
nor U819 (N_819,N_781,N_766);
or U820 (N_820,N_772,N_751);
or U821 (N_821,N_779,N_788);
nor U822 (N_822,N_723,N_768);
and U823 (N_823,N_736,N_753);
and U824 (N_824,N_797,N_748);
or U825 (N_825,N_730,N_729);
or U826 (N_826,N_756,N_791);
or U827 (N_827,N_743,N_710);
nand U828 (N_828,N_719,N_764);
xnor U829 (N_829,N_733,N_785);
nor U830 (N_830,N_701,N_776);
nor U831 (N_831,N_763,N_706);
xor U832 (N_832,N_782,N_738);
nor U833 (N_833,N_722,N_732);
nand U834 (N_834,N_799,N_735);
and U835 (N_835,N_740,N_786);
nor U836 (N_836,N_762,N_720);
or U837 (N_837,N_707,N_747);
nand U838 (N_838,N_798,N_789);
or U839 (N_839,N_757,N_780);
nand U840 (N_840,N_792,N_704);
and U841 (N_841,N_773,N_703);
nor U842 (N_842,N_721,N_741);
and U843 (N_843,N_742,N_744);
and U844 (N_844,N_759,N_708);
nor U845 (N_845,N_771,N_755);
and U846 (N_846,N_739,N_709);
or U847 (N_847,N_794,N_765);
or U848 (N_848,N_790,N_702);
xor U849 (N_849,N_714,N_793);
and U850 (N_850,N_749,N_753);
and U851 (N_851,N_733,N_778);
or U852 (N_852,N_736,N_733);
and U853 (N_853,N_772,N_707);
nand U854 (N_854,N_795,N_797);
nand U855 (N_855,N_777,N_713);
nor U856 (N_856,N_788,N_701);
and U857 (N_857,N_733,N_795);
and U858 (N_858,N_763,N_753);
nor U859 (N_859,N_736,N_705);
nand U860 (N_860,N_719,N_728);
nor U861 (N_861,N_774,N_778);
and U862 (N_862,N_773,N_729);
or U863 (N_863,N_707,N_718);
or U864 (N_864,N_714,N_788);
nor U865 (N_865,N_764,N_703);
nand U866 (N_866,N_789,N_716);
nor U867 (N_867,N_716,N_780);
or U868 (N_868,N_795,N_742);
nor U869 (N_869,N_739,N_795);
and U870 (N_870,N_783,N_780);
nand U871 (N_871,N_793,N_730);
nand U872 (N_872,N_796,N_777);
or U873 (N_873,N_706,N_757);
or U874 (N_874,N_776,N_735);
nand U875 (N_875,N_717,N_758);
and U876 (N_876,N_751,N_739);
nor U877 (N_877,N_749,N_719);
nand U878 (N_878,N_796,N_789);
and U879 (N_879,N_711,N_710);
nor U880 (N_880,N_716,N_709);
nor U881 (N_881,N_741,N_730);
nor U882 (N_882,N_721,N_789);
nand U883 (N_883,N_769,N_719);
or U884 (N_884,N_797,N_770);
and U885 (N_885,N_740,N_763);
nand U886 (N_886,N_715,N_703);
and U887 (N_887,N_765,N_725);
nor U888 (N_888,N_711,N_763);
or U889 (N_889,N_748,N_790);
and U890 (N_890,N_701,N_737);
and U891 (N_891,N_789,N_707);
or U892 (N_892,N_727,N_752);
nand U893 (N_893,N_761,N_717);
nor U894 (N_894,N_723,N_730);
nor U895 (N_895,N_798,N_778);
nor U896 (N_896,N_705,N_744);
or U897 (N_897,N_779,N_756);
or U898 (N_898,N_738,N_785);
nor U899 (N_899,N_701,N_708);
or U900 (N_900,N_840,N_850);
or U901 (N_901,N_889,N_883);
nor U902 (N_902,N_828,N_870);
or U903 (N_903,N_896,N_837);
nand U904 (N_904,N_801,N_859);
and U905 (N_905,N_876,N_842);
nor U906 (N_906,N_861,N_818);
or U907 (N_907,N_862,N_858);
nand U908 (N_908,N_874,N_817);
or U909 (N_909,N_891,N_833);
nand U910 (N_910,N_802,N_822);
nor U911 (N_911,N_823,N_807);
and U912 (N_912,N_879,N_846);
nor U913 (N_913,N_814,N_897);
nand U914 (N_914,N_866,N_831);
nand U915 (N_915,N_830,N_852);
or U916 (N_916,N_881,N_860);
or U917 (N_917,N_853,N_893);
nor U918 (N_918,N_899,N_834);
nand U919 (N_919,N_829,N_886);
nand U920 (N_920,N_884,N_895);
nor U921 (N_921,N_868,N_836);
nor U922 (N_922,N_841,N_890);
or U923 (N_923,N_839,N_878);
nand U924 (N_924,N_810,N_875);
and U925 (N_925,N_885,N_844);
or U926 (N_926,N_894,N_892);
and U927 (N_927,N_812,N_819);
nor U928 (N_928,N_804,N_863);
or U929 (N_929,N_813,N_882);
nor U930 (N_930,N_898,N_869);
and U931 (N_931,N_851,N_816);
or U932 (N_932,N_815,N_827);
nand U933 (N_933,N_872,N_887);
or U934 (N_934,N_888,N_877);
nand U935 (N_935,N_847,N_800);
and U936 (N_936,N_803,N_809);
or U937 (N_937,N_805,N_806);
nor U938 (N_938,N_826,N_871);
nor U939 (N_939,N_843,N_857);
nand U940 (N_940,N_820,N_854);
and U941 (N_941,N_880,N_838);
nand U942 (N_942,N_848,N_849);
or U943 (N_943,N_824,N_873);
and U944 (N_944,N_865,N_864);
and U945 (N_945,N_845,N_867);
nor U946 (N_946,N_821,N_856);
nand U947 (N_947,N_832,N_825);
nor U948 (N_948,N_835,N_808);
nor U949 (N_949,N_811,N_855);
and U950 (N_950,N_835,N_875);
or U951 (N_951,N_811,N_825);
or U952 (N_952,N_867,N_830);
nor U953 (N_953,N_853,N_819);
and U954 (N_954,N_877,N_859);
and U955 (N_955,N_841,N_855);
and U956 (N_956,N_866,N_822);
nand U957 (N_957,N_820,N_819);
and U958 (N_958,N_827,N_876);
nand U959 (N_959,N_896,N_847);
or U960 (N_960,N_897,N_898);
nand U961 (N_961,N_890,N_817);
nor U962 (N_962,N_827,N_889);
nor U963 (N_963,N_899,N_860);
nand U964 (N_964,N_885,N_812);
nor U965 (N_965,N_873,N_837);
and U966 (N_966,N_877,N_875);
or U967 (N_967,N_862,N_856);
and U968 (N_968,N_817,N_875);
or U969 (N_969,N_863,N_867);
or U970 (N_970,N_820,N_865);
nor U971 (N_971,N_857,N_807);
or U972 (N_972,N_847,N_848);
or U973 (N_973,N_845,N_869);
nand U974 (N_974,N_861,N_837);
nand U975 (N_975,N_835,N_853);
and U976 (N_976,N_807,N_885);
xor U977 (N_977,N_828,N_819);
or U978 (N_978,N_869,N_887);
and U979 (N_979,N_899,N_810);
nor U980 (N_980,N_868,N_857);
and U981 (N_981,N_809,N_831);
nor U982 (N_982,N_870,N_853);
nand U983 (N_983,N_853,N_848);
nand U984 (N_984,N_890,N_893);
or U985 (N_985,N_847,N_859);
and U986 (N_986,N_862,N_815);
nor U987 (N_987,N_821,N_818);
nor U988 (N_988,N_899,N_882);
or U989 (N_989,N_824,N_835);
or U990 (N_990,N_831,N_897);
nand U991 (N_991,N_810,N_874);
or U992 (N_992,N_876,N_863);
nor U993 (N_993,N_881,N_891);
or U994 (N_994,N_885,N_852);
nor U995 (N_995,N_831,N_800);
and U996 (N_996,N_842,N_895);
and U997 (N_997,N_883,N_873);
nand U998 (N_998,N_822,N_886);
and U999 (N_999,N_851,N_872);
nor U1000 (N_1000,N_954,N_974);
and U1001 (N_1001,N_935,N_916);
or U1002 (N_1002,N_943,N_977);
and U1003 (N_1003,N_988,N_957);
nor U1004 (N_1004,N_989,N_992);
or U1005 (N_1005,N_956,N_959);
nand U1006 (N_1006,N_993,N_901);
and U1007 (N_1007,N_990,N_928);
and U1008 (N_1008,N_965,N_925);
and U1009 (N_1009,N_921,N_994);
nand U1010 (N_1010,N_930,N_955);
and U1011 (N_1011,N_927,N_960);
nand U1012 (N_1012,N_922,N_953);
or U1013 (N_1013,N_917,N_906);
nand U1014 (N_1014,N_948,N_910);
or U1015 (N_1015,N_966,N_939);
nand U1016 (N_1016,N_982,N_940);
nand U1017 (N_1017,N_946,N_914);
or U1018 (N_1018,N_942,N_972);
nor U1019 (N_1019,N_996,N_950);
and U1020 (N_1020,N_947,N_980);
and U1021 (N_1021,N_924,N_912);
nand U1022 (N_1022,N_918,N_981);
and U1023 (N_1023,N_911,N_976);
and U1024 (N_1024,N_937,N_920);
and U1025 (N_1025,N_936,N_961);
nand U1026 (N_1026,N_978,N_951);
nand U1027 (N_1027,N_984,N_997);
and U1028 (N_1028,N_934,N_986);
and U1029 (N_1029,N_971,N_931);
nand U1030 (N_1030,N_949,N_983);
nor U1031 (N_1031,N_926,N_915);
and U1032 (N_1032,N_970,N_933);
nand U1033 (N_1033,N_913,N_932);
and U1034 (N_1034,N_905,N_938);
or U1035 (N_1035,N_969,N_929);
nand U1036 (N_1036,N_958,N_967);
and U1037 (N_1037,N_945,N_987);
nor U1038 (N_1038,N_903,N_995);
nor U1039 (N_1039,N_907,N_998);
or U1040 (N_1040,N_902,N_941);
and U1041 (N_1041,N_923,N_975);
or U1042 (N_1042,N_900,N_973);
and U1043 (N_1043,N_904,N_908);
or U1044 (N_1044,N_919,N_963);
or U1045 (N_1045,N_964,N_985);
nor U1046 (N_1046,N_991,N_944);
nand U1047 (N_1047,N_952,N_968);
and U1048 (N_1048,N_962,N_999);
and U1049 (N_1049,N_909,N_979);
and U1050 (N_1050,N_914,N_936);
nor U1051 (N_1051,N_941,N_908);
and U1052 (N_1052,N_948,N_928);
or U1053 (N_1053,N_909,N_993);
or U1054 (N_1054,N_996,N_982);
nor U1055 (N_1055,N_973,N_993);
nor U1056 (N_1056,N_910,N_919);
nor U1057 (N_1057,N_987,N_934);
and U1058 (N_1058,N_999,N_922);
and U1059 (N_1059,N_986,N_927);
nor U1060 (N_1060,N_938,N_970);
and U1061 (N_1061,N_907,N_978);
and U1062 (N_1062,N_939,N_904);
or U1063 (N_1063,N_961,N_988);
and U1064 (N_1064,N_943,N_934);
nor U1065 (N_1065,N_992,N_958);
nand U1066 (N_1066,N_977,N_910);
or U1067 (N_1067,N_983,N_920);
and U1068 (N_1068,N_919,N_924);
nor U1069 (N_1069,N_903,N_949);
nor U1070 (N_1070,N_978,N_926);
and U1071 (N_1071,N_962,N_959);
nand U1072 (N_1072,N_924,N_901);
or U1073 (N_1073,N_974,N_979);
or U1074 (N_1074,N_972,N_981);
nor U1075 (N_1075,N_954,N_934);
and U1076 (N_1076,N_968,N_993);
and U1077 (N_1077,N_955,N_979);
or U1078 (N_1078,N_951,N_934);
or U1079 (N_1079,N_901,N_974);
and U1080 (N_1080,N_912,N_963);
nor U1081 (N_1081,N_988,N_940);
nor U1082 (N_1082,N_957,N_943);
nand U1083 (N_1083,N_911,N_997);
or U1084 (N_1084,N_965,N_930);
nor U1085 (N_1085,N_906,N_963);
nor U1086 (N_1086,N_919,N_906);
nor U1087 (N_1087,N_936,N_988);
nand U1088 (N_1088,N_964,N_950);
and U1089 (N_1089,N_995,N_976);
and U1090 (N_1090,N_912,N_920);
or U1091 (N_1091,N_964,N_938);
or U1092 (N_1092,N_989,N_959);
nor U1093 (N_1093,N_990,N_944);
or U1094 (N_1094,N_996,N_997);
or U1095 (N_1095,N_993,N_904);
and U1096 (N_1096,N_970,N_931);
and U1097 (N_1097,N_952,N_935);
and U1098 (N_1098,N_994,N_956);
nand U1099 (N_1099,N_986,N_913);
and U1100 (N_1100,N_1032,N_1054);
nor U1101 (N_1101,N_1001,N_1025);
nor U1102 (N_1102,N_1019,N_1085);
nor U1103 (N_1103,N_1066,N_1013);
nand U1104 (N_1104,N_1090,N_1069);
nor U1105 (N_1105,N_1089,N_1075);
or U1106 (N_1106,N_1059,N_1092);
or U1107 (N_1107,N_1036,N_1060);
nor U1108 (N_1108,N_1015,N_1061);
nand U1109 (N_1109,N_1065,N_1020);
or U1110 (N_1110,N_1047,N_1000);
and U1111 (N_1111,N_1080,N_1033);
nand U1112 (N_1112,N_1028,N_1055);
nand U1113 (N_1113,N_1037,N_1039);
nand U1114 (N_1114,N_1008,N_1004);
nor U1115 (N_1115,N_1067,N_1035);
nor U1116 (N_1116,N_1043,N_1094);
or U1117 (N_1117,N_1082,N_1083);
nor U1118 (N_1118,N_1009,N_1062);
nand U1119 (N_1119,N_1003,N_1081);
nor U1120 (N_1120,N_1063,N_1005);
and U1121 (N_1121,N_1058,N_1002);
or U1122 (N_1122,N_1068,N_1014);
and U1123 (N_1123,N_1064,N_1031);
nand U1124 (N_1124,N_1057,N_1016);
or U1125 (N_1125,N_1098,N_1018);
nand U1126 (N_1126,N_1097,N_1029);
nand U1127 (N_1127,N_1088,N_1091);
and U1128 (N_1128,N_1022,N_1044);
and U1129 (N_1129,N_1076,N_1038);
or U1130 (N_1130,N_1079,N_1021);
nand U1131 (N_1131,N_1041,N_1049);
nand U1132 (N_1132,N_1023,N_1086);
nand U1133 (N_1133,N_1045,N_1072);
nor U1134 (N_1134,N_1074,N_1078);
and U1135 (N_1135,N_1042,N_1099);
or U1136 (N_1136,N_1027,N_1046);
nor U1137 (N_1137,N_1050,N_1095);
nor U1138 (N_1138,N_1077,N_1051);
nand U1139 (N_1139,N_1070,N_1096);
or U1140 (N_1140,N_1034,N_1006);
and U1141 (N_1141,N_1048,N_1017);
nand U1142 (N_1142,N_1040,N_1052);
and U1143 (N_1143,N_1026,N_1011);
or U1144 (N_1144,N_1087,N_1053);
and U1145 (N_1145,N_1024,N_1012);
and U1146 (N_1146,N_1073,N_1010);
nor U1147 (N_1147,N_1030,N_1093);
nor U1148 (N_1148,N_1056,N_1084);
nand U1149 (N_1149,N_1007,N_1071);
nor U1150 (N_1150,N_1018,N_1085);
or U1151 (N_1151,N_1003,N_1011);
or U1152 (N_1152,N_1021,N_1014);
nor U1153 (N_1153,N_1054,N_1014);
or U1154 (N_1154,N_1007,N_1008);
nand U1155 (N_1155,N_1052,N_1085);
nand U1156 (N_1156,N_1005,N_1072);
nor U1157 (N_1157,N_1009,N_1091);
nand U1158 (N_1158,N_1069,N_1005);
nor U1159 (N_1159,N_1012,N_1029);
or U1160 (N_1160,N_1097,N_1093);
or U1161 (N_1161,N_1066,N_1078);
and U1162 (N_1162,N_1047,N_1022);
nor U1163 (N_1163,N_1069,N_1097);
and U1164 (N_1164,N_1045,N_1090);
nor U1165 (N_1165,N_1061,N_1014);
and U1166 (N_1166,N_1065,N_1017);
nor U1167 (N_1167,N_1012,N_1055);
or U1168 (N_1168,N_1058,N_1080);
nand U1169 (N_1169,N_1096,N_1093);
nand U1170 (N_1170,N_1094,N_1037);
and U1171 (N_1171,N_1023,N_1096);
nor U1172 (N_1172,N_1068,N_1057);
nor U1173 (N_1173,N_1023,N_1016);
or U1174 (N_1174,N_1018,N_1089);
and U1175 (N_1175,N_1081,N_1043);
nand U1176 (N_1176,N_1007,N_1018);
and U1177 (N_1177,N_1015,N_1005);
or U1178 (N_1178,N_1090,N_1009);
nand U1179 (N_1179,N_1063,N_1045);
or U1180 (N_1180,N_1085,N_1088);
and U1181 (N_1181,N_1096,N_1069);
nand U1182 (N_1182,N_1053,N_1054);
nand U1183 (N_1183,N_1070,N_1018);
and U1184 (N_1184,N_1081,N_1084);
nand U1185 (N_1185,N_1060,N_1013);
nor U1186 (N_1186,N_1011,N_1001);
nand U1187 (N_1187,N_1012,N_1034);
xnor U1188 (N_1188,N_1082,N_1084);
nand U1189 (N_1189,N_1067,N_1093);
or U1190 (N_1190,N_1096,N_1047);
and U1191 (N_1191,N_1002,N_1004);
or U1192 (N_1192,N_1020,N_1027);
and U1193 (N_1193,N_1054,N_1036);
and U1194 (N_1194,N_1000,N_1092);
or U1195 (N_1195,N_1028,N_1075);
nand U1196 (N_1196,N_1028,N_1093);
nand U1197 (N_1197,N_1002,N_1046);
or U1198 (N_1198,N_1021,N_1057);
nand U1199 (N_1199,N_1028,N_1002);
nor U1200 (N_1200,N_1151,N_1119);
or U1201 (N_1201,N_1149,N_1158);
nor U1202 (N_1202,N_1178,N_1120);
and U1203 (N_1203,N_1131,N_1127);
nor U1204 (N_1204,N_1116,N_1150);
nand U1205 (N_1205,N_1161,N_1136);
and U1206 (N_1206,N_1137,N_1189);
nand U1207 (N_1207,N_1174,N_1142);
and U1208 (N_1208,N_1160,N_1141);
or U1209 (N_1209,N_1115,N_1176);
or U1210 (N_1210,N_1130,N_1187);
nor U1211 (N_1211,N_1125,N_1193);
xor U1212 (N_1212,N_1169,N_1152);
or U1213 (N_1213,N_1162,N_1113);
nand U1214 (N_1214,N_1110,N_1121);
or U1215 (N_1215,N_1170,N_1177);
nand U1216 (N_1216,N_1199,N_1139);
nand U1217 (N_1217,N_1167,N_1103);
nand U1218 (N_1218,N_1179,N_1146);
or U1219 (N_1219,N_1107,N_1126);
and U1220 (N_1220,N_1145,N_1155);
and U1221 (N_1221,N_1117,N_1147);
nor U1222 (N_1222,N_1123,N_1192);
or U1223 (N_1223,N_1191,N_1132);
nor U1224 (N_1224,N_1109,N_1184);
or U1225 (N_1225,N_1180,N_1194);
nor U1226 (N_1226,N_1181,N_1106);
and U1227 (N_1227,N_1190,N_1112);
nor U1228 (N_1228,N_1159,N_1171);
and U1229 (N_1229,N_1148,N_1166);
nand U1230 (N_1230,N_1122,N_1173);
nor U1231 (N_1231,N_1165,N_1111);
and U1232 (N_1232,N_1183,N_1108);
nor U1233 (N_1233,N_1196,N_1134);
nor U1234 (N_1234,N_1140,N_1154);
or U1235 (N_1235,N_1197,N_1156);
nand U1236 (N_1236,N_1198,N_1105);
xnor U1237 (N_1237,N_1143,N_1124);
or U1238 (N_1238,N_1114,N_1195);
nor U1239 (N_1239,N_1144,N_1153);
or U1240 (N_1240,N_1172,N_1101);
or U1241 (N_1241,N_1102,N_1175);
or U1242 (N_1242,N_1182,N_1163);
nor U1243 (N_1243,N_1157,N_1185);
and U1244 (N_1244,N_1186,N_1138);
nor U1245 (N_1245,N_1188,N_1168);
and U1246 (N_1246,N_1135,N_1104);
nor U1247 (N_1247,N_1129,N_1133);
nand U1248 (N_1248,N_1164,N_1128);
nand U1249 (N_1249,N_1100,N_1118);
and U1250 (N_1250,N_1191,N_1194);
nand U1251 (N_1251,N_1105,N_1154);
or U1252 (N_1252,N_1115,N_1186);
and U1253 (N_1253,N_1178,N_1164);
nor U1254 (N_1254,N_1174,N_1172);
and U1255 (N_1255,N_1194,N_1140);
or U1256 (N_1256,N_1181,N_1103);
xnor U1257 (N_1257,N_1145,N_1186);
nor U1258 (N_1258,N_1132,N_1134);
nor U1259 (N_1259,N_1187,N_1197);
nand U1260 (N_1260,N_1127,N_1162);
and U1261 (N_1261,N_1141,N_1184);
and U1262 (N_1262,N_1114,N_1141);
nand U1263 (N_1263,N_1115,N_1178);
nor U1264 (N_1264,N_1120,N_1102);
and U1265 (N_1265,N_1117,N_1112);
or U1266 (N_1266,N_1188,N_1194);
nand U1267 (N_1267,N_1195,N_1107);
and U1268 (N_1268,N_1118,N_1194);
nor U1269 (N_1269,N_1153,N_1181);
or U1270 (N_1270,N_1137,N_1174);
nor U1271 (N_1271,N_1153,N_1189);
nand U1272 (N_1272,N_1164,N_1182);
nand U1273 (N_1273,N_1172,N_1125);
nand U1274 (N_1274,N_1111,N_1119);
or U1275 (N_1275,N_1159,N_1184);
or U1276 (N_1276,N_1183,N_1188);
and U1277 (N_1277,N_1128,N_1176);
or U1278 (N_1278,N_1146,N_1147);
nor U1279 (N_1279,N_1124,N_1187);
nor U1280 (N_1280,N_1162,N_1153);
nand U1281 (N_1281,N_1183,N_1143);
nand U1282 (N_1282,N_1127,N_1152);
nor U1283 (N_1283,N_1120,N_1140);
or U1284 (N_1284,N_1198,N_1154);
nor U1285 (N_1285,N_1126,N_1185);
and U1286 (N_1286,N_1100,N_1146);
nand U1287 (N_1287,N_1123,N_1129);
and U1288 (N_1288,N_1149,N_1137);
nor U1289 (N_1289,N_1154,N_1115);
and U1290 (N_1290,N_1170,N_1112);
or U1291 (N_1291,N_1102,N_1104);
nor U1292 (N_1292,N_1116,N_1186);
and U1293 (N_1293,N_1196,N_1133);
or U1294 (N_1294,N_1149,N_1118);
nor U1295 (N_1295,N_1150,N_1195);
and U1296 (N_1296,N_1103,N_1185);
and U1297 (N_1297,N_1155,N_1177);
nor U1298 (N_1298,N_1117,N_1185);
or U1299 (N_1299,N_1133,N_1121);
nor U1300 (N_1300,N_1228,N_1206);
nand U1301 (N_1301,N_1292,N_1204);
nor U1302 (N_1302,N_1284,N_1257);
nor U1303 (N_1303,N_1288,N_1200);
or U1304 (N_1304,N_1263,N_1245);
and U1305 (N_1305,N_1217,N_1213);
nand U1306 (N_1306,N_1272,N_1259);
and U1307 (N_1307,N_1248,N_1238);
and U1308 (N_1308,N_1207,N_1255);
nor U1309 (N_1309,N_1244,N_1254);
nand U1310 (N_1310,N_1222,N_1246);
nor U1311 (N_1311,N_1201,N_1275);
nor U1312 (N_1312,N_1289,N_1237);
or U1313 (N_1313,N_1294,N_1266);
or U1314 (N_1314,N_1277,N_1282);
or U1315 (N_1315,N_1240,N_1247);
nand U1316 (N_1316,N_1216,N_1283);
and U1317 (N_1317,N_1256,N_1202);
or U1318 (N_1318,N_1230,N_1208);
nand U1319 (N_1319,N_1205,N_1270);
nand U1320 (N_1320,N_1295,N_1210);
or U1321 (N_1321,N_1251,N_1220);
or U1322 (N_1322,N_1279,N_1224);
xor U1323 (N_1323,N_1232,N_1274);
and U1324 (N_1324,N_1223,N_1226);
or U1325 (N_1325,N_1268,N_1241);
nand U1326 (N_1326,N_1293,N_1233);
and U1327 (N_1327,N_1265,N_1219);
nand U1328 (N_1328,N_1273,N_1296);
and U1329 (N_1329,N_1229,N_1299);
and U1330 (N_1330,N_1214,N_1227);
nand U1331 (N_1331,N_1235,N_1212);
nand U1332 (N_1332,N_1242,N_1203);
nor U1333 (N_1333,N_1271,N_1211);
xnor U1334 (N_1334,N_1258,N_1234);
or U1335 (N_1335,N_1286,N_1215);
or U1336 (N_1336,N_1218,N_1225);
and U1337 (N_1337,N_1278,N_1285);
nand U1338 (N_1338,N_1221,N_1269);
and U1339 (N_1339,N_1239,N_1281);
nand U1340 (N_1340,N_1260,N_1298);
nor U1341 (N_1341,N_1236,N_1209);
nor U1342 (N_1342,N_1267,N_1261);
nand U1343 (N_1343,N_1291,N_1252);
nor U1344 (N_1344,N_1253,N_1287);
nor U1345 (N_1345,N_1262,N_1231);
or U1346 (N_1346,N_1250,N_1280);
and U1347 (N_1347,N_1243,N_1276);
and U1348 (N_1348,N_1290,N_1249);
nand U1349 (N_1349,N_1297,N_1264);
nor U1350 (N_1350,N_1266,N_1259);
nor U1351 (N_1351,N_1230,N_1287);
and U1352 (N_1352,N_1228,N_1217);
or U1353 (N_1353,N_1214,N_1228);
nor U1354 (N_1354,N_1296,N_1219);
nor U1355 (N_1355,N_1260,N_1208);
or U1356 (N_1356,N_1228,N_1226);
nand U1357 (N_1357,N_1230,N_1265);
or U1358 (N_1358,N_1270,N_1259);
or U1359 (N_1359,N_1251,N_1275);
and U1360 (N_1360,N_1298,N_1286);
nand U1361 (N_1361,N_1289,N_1287);
or U1362 (N_1362,N_1244,N_1223);
or U1363 (N_1363,N_1239,N_1235);
nor U1364 (N_1364,N_1208,N_1261);
nor U1365 (N_1365,N_1287,N_1223);
nor U1366 (N_1366,N_1291,N_1246);
xor U1367 (N_1367,N_1281,N_1228);
nor U1368 (N_1368,N_1216,N_1296);
or U1369 (N_1369,N_1251,N_1268);
nand U1370 (N_1370,N_1276,N_1266);
or U1371 (N_1371,N_1218,N_1295);
and U1372 (N_1372,N_1201,N_1258);
or U1373 (N_1373,N_1239,N_1225);
or U1374 (N_1374,N_1255,N_1233);
xor U1375 (N_1375,N_1212,N_1229);
nor U1376 (N_1376,N_1286,N_1246);
or U1377 (N_1377,N_1263,N_1223);
nand U1378 (N_1378,N_1299,N_1266);
and U1379 (N_1379,N_1278,N_1261);
nand U1380 (N_1380,N_1280,N_1208);
nand U1381 (N_1381,N_1296,N_1222);
or U1382 (N_1382,N_1280,N_1206);
and U1383 (N_1383,N_1276,N_1236);
or U1384 (N_1384,N_1283,N_1249);
or U1385 (N_1385,N_1240,N_1252);
nand U1386 (N_1386,N_1289,N_1265);
and U1387 (N_1387,N_1264,N_1293);
nand U1388 (N_1388,N_1272,N_1207);
or U1389 (N_1389,N_1216,N_1243);
nand U1390 (N_1390,N_1256,N_1272);
nand U1391 (N_1391,N_1202,N_1253);
and U1392 (N_1392,N_1270,N_1225);
nor U1393 (N_1393,N_1261,N_1275);
nand U1394 (N_1394,N_1217,N_1206);
nand U1395 (N_1395,N_1283,N_1218);
nand U1396 (N_1396,N_1261,N_1236);
nand U1397 (N_1397,N_1244,N_1219);
nand U1398 (N_1398,N_1232,N_1280);
nor U1399 (N_1399,N_1248,N_1211);
and U1400 (N_1400,N_1342,N_1314);
nor U1401 (N_1401,N_1304,N_1329);
xnor U1402 (N_1402,N_1372,N_1376);
nor U1403 (N_1403,N_1374,N_1363);
nand U1404 (N_1404,N_1375,N_1357);
nor U1405 (N_1405,N_1350,N_1378);
nor U1406 (N_1406,N_1356,N_1339);
nand U1407 (N_1407,N_1340,N_1393);
nor U1408 (N_1408,N_1365,N_1353);
and U1409 (N_1409,N_1377,N_1300);
or U1410 (N_1410,N_1351,N_1327);
nor U1411 (N_1411,N_1328,N_1334);
nor U1412 (N_1412,N_1325,N_1320);
or U1413 (N_1413,N_1383,N_1366);
nor U1414 (N_1414,N_1367,N_1326);
nor U1415 (N_1415,N_1312,N_1370);
nor U1416 (N_1416,N_1362,N_1315);
and U1417 (N_1417,N_1310,N_1371);
nand U1418 (N_1418,N_1324,N_1360);
nor U1419 (N_1419,N_1332,N_1346);
nor U1420 (N_1420,N_1317,N_1380);
nor U1421 (N_1421,N_1311,N_1349);
or U1422 (N_1422,N_1358,N_1382);
or U1423 (N_1423,N_1348,N_1384);
and U1424 (N_1424,N_1345,N_1308);
or U1425 (N_1425,N_1323,N_1335);
nor U1426 (N_1426,N_1337,N_1387);
nor U1427 (N_1427,N_1313,N_1305);
nand U1428 (N_1428,N_1397,N_1399);
or U1429 (N_1429,N_1373,N_1390);
nor U1430 (N_1430,N_1319,N_1364);
or U1431 (N_1431,N_1386,N_1391);
nand U1432 (N_1432,N_1321,N_1306);
nand U1433 (N_1433,N_1318,N_1394);
nor U1434 (N_1434,N_1396,N_1368);
nand U1435 (N_1435,N_1354,N_1316);
or U1436 (N_1436,N_1389,N_1381);
nand U1437 (N_1437,N_1388,N_1338);
nand U1438 (N_1438,N_1361,N_1369);
or U1439 (N_1439,N_1330,N_1303);
and U1440 (N_1440,N_1302,N_1359);
nand U1441 (N_1441,N_1331,N_1352);
nand U1442 (N_1442,N_1336,N_1385);
and U1443 (N_1443,N_1333,N_1395);
nor U1444 (N_1444,N_1307,N_1398);
and U1445 (N_1445,N_1322,N_1341);
nor U1446 (N_1446,N_1355,N_1392);
nor U1447 (N_1447,N_1344,N_1379);
nand U1448 (N_1448,N_1347,N_1309);
nor U1449 (N_1449,N_1343,N_1301);
and U1450 (N_1450,N_1324,N_1304);
or U1451 (N_1451,N_1357,N_1309);
and U1452 (N_1452,N_1320,N_1378);
and U1453 (N_1453,N_1344,N_1317);
nor U1454 (N_1454,N_1327,N_1357);
nand U1455 (N_1455,N_1300,N_1394);
nor U1456 (N_1456,N_1377,N_1320);
and U1457 (N_1457,N_1316,N_1375);
nor U1458 (N_1458,N_1359,N_1310);
or U1459 (N_1459,N_1301,N_1303);
nand U1460 (N_1460,N_1394,N_1373);
nor U1461 (N_1461,N_1315,N_1396);
and U1462 (N_1462,N_1313,N_1334);
nand U1463 (N_1463,N_1352,N_1321);
nand U1464 (N_1464,N_1340,N_1310);
nand U1465 (N_1465,N_1309,N_1368);
or U1466 (N_1466,N_1352,N_1382);
nand U1467 (N_1467,N_1322,N_1308);
or U1468 (N_1468,N_1315,N_1393);
and U1469 (N_1469,N_1333,N_1301);
or U1470 (N_1470,N_1319,N_1321);
nor U1471 (N_1471,N_1390,N_1388);
or U1472 (N_1472,N_1366,N_1304);
nor U1473 (N_1473,N_1391,N_1375);
or U1474 (N_1474,N_1316,N_1313);
and U1475 (N_1475,N_1372,N_1375);
nand U1476 (N_1476,N_1337,N_1311);
xor U1477 (N_1477,N_1396,N_1330);
nor U1478 (N_1478,N_1346,N_1395);
nand U1479 (N_1479,N_1335,N_1307);
nor U1480 (N_1480,N_1318,N_1361);
and U1481 (N_1481,N_1303,N_1320);
nor U1482 (N_1482,N_1321,N_1399);
and U1483 (N_1483,N_1308,N_1310);
nand U1484 (N_1484,N_1399,N_1330);
nand U1485 (N_1485,N_1302,N_1351);
and U1486 (N_1486,N_1342,N_1376);
or U1487 (N_1487,N_1319,N_1396);
nor U1488 (N_1488,N_1388,N_1366);
nand U1489 (N_1489,N_1392,N_1332);
or U1490 (N_1490,N_1304,N_1368);
nand U1491 (N_1491,N_1300,N_1340);
nor U1492 (N_1492,N_1385,N_1395);
nor U1493 (N_1493,N_1376,N_1384);
nand U1494 (N_1494,N_1319,N_1383);
nand U1495 (N_1495,N_1331,N_1361);
and U1496 (N_1496,N_1334,N_1347);
and U1497 (N_1497,N_1385,N_1362);
or U1498 (N_1498,N_1314,N_1307);
nand U1499 (N_1499,N_1381,N_1355);
or U1500 (N_1500,N_1499,N_1484);
or U1501 (N_1501,N_1440,N_1458);
or U1502 (N_1502,N_1491,N_1456);
and U1503 (N_1503,N_1413,N_1414);
or U1504 (N_1504,N_1416,N_1481);
nor U1505 (N_1505,N_1452,N_1429);
and U1506 (N_1506,N_1477,N_1442);
nor U1507 (N_1507,N_1462,N_1451);
nor U1508 (N_1508,N_1447,N_1431);
nand U1509 (N_1509,N_1479,N_1423);
and U1510 (N_1510,N_1426,N_1478);
and U1511 (N_1511,N_1444,N_1428);
nand U1512 (N_1512,N_1417,N_1469);
and U1513 (N_1513,N_1492,N_1437);
nor U1514 (N_1514,N_1403,N_1438);
nor U1515 (N_1515,N_1471,N_1483);
nor U1516 (N_1516,N_1496,N_1455);
nor U1517 (N_1517,N_1405,N_1486);
and U1518 (N_1518,N_1432,N_1445);
and U1519 (N_1519,N_1480,N_1488);
nand U1520 (N_1520,N_1402,N_1436);
nand U1521 (N_1521,N_1422,N_1421);
nor U1522 (N_1522,N_1474,N_1485);
nand U1523 (N_1523,N_1461,N_1419);
nor U1524 (N_1524,N_1408,N_1441);
nor U1525 (N_1525,N_1410,N_1439);
or U1526 (N_1526,N_1404,N_1424);
and U1527 (N_1527,N_1450,N_1427);
nor U1528 (N_1528,N_1464,N_1446);
and U1529 (N_1529,N_1459,N_1487);
and U1530 (N_1530,N_1415,N_1490);
nand U1531 (N_1531,N_1406,N_1453);
and U1532 (N_1532,N_1435,N_1467);
xnor U1533 (N_1533,N_1489,N_1430);
and U1534 (N_1534,N_1412,N_1457);
nor U1535 (N_1535,N_1448,N_1466);
nor U1536 (N_1536,N_1468,N_1401);
nor U1537 (N_1537,N_1470,N_1409);
and U1538 (N_1538,N_1476,N_1420);
or U1539 (N_1539,N_1495,N_1400);
and U1540 (N_1540,N_1443,N_1454);
nor U1541 (N_1541,N_1465,N_1460);
nor U1542 (N_1542,N_1449,N_1482);
nand U1543 (N_1543,N_1411,N_1433);
nand U1544 (N_1544,N_1497,N_1493);
xor U1545 (N_1545,N_1407,N_1463);
nor U1546 (N_1546,N_1473,N_1425);
or U1547 (N_1547,N_1494,N_1498);
or U1548 (N_1548,N_1472,N_1475);
and U1549 (N_1549,N_1434,N_1418);
nor U1550 (N_1550,N_1438,N_1450);
and U1551 (N_1551,N_1448,N_1445);
nor U1552 (N_1552,N_1469,N_1438);
nand U1553 (N_1553,N_1439,N_1426);
and U1554 (N_1554,N_1409,N_1407);
nor U1555 (N_1555,N_1464,N_1405);
nand U1556 (N_1556,N_1421,N_1408);
or U1557 (N_1557,N_1433,N_1496);
or U1558 (N_1558,N_1483,N_1453);
or U1559 (N_1559,N_1433,N_1451);
or U1560 (N_1560,N_1491,N_1438);
nor U1561 (N_1561,N_1436,N_1412);
nor U1562 (N_1562,N_1408,N_1483);
nand U1563 (N_1563,N_1492,N_1465);
and U1564 (N_1564,N_1427,N_1423);
nand U1565 (N_1565,N_1444,N_1432);
and U1566 (N_1566,N_1420,N_1434);
nor U1567 (N_1567,N_1486,N_1442);
nand U1568 (N_1568,N_1427,N_1444);
and U1569 (N_1569,N_1480,N_1404);
and U1570 (N_1570,N_1448,N_1497);
xor U1571 (N_1571,N_1476,N_1435);
and U1572 (N_1572,N_1422,N_1428);
nand U1573 (N_1573,N_1409,N_1490);
nor U1574 (N_1574,N_1411,N_1458);
nor U1575 (N_1575,N_1409,N_1442);
or U1576 (N_1576,N_1459,N_1409);
or U1577 (N_1577,N_1414,N_1422);
or U1578 (N_1578,N_1498,N_1448);
or U1579 (N_1579,N_1437,N_1499);
nor U1580 (N_1580,N_1416,N_1434);
or U1581 (N_1581,N_1402,N_1416);
or U1582 (N_1582,N_1474,N_1406);
nand U1583 (N_1583,N_1466,N_1498);
or U1584 (N_1584,N_1405,N_1456);
nor U1585 (N_1585,N_1440,N_1400);
nor U1586 (N_1586,N_1488,N_1445);
nand U1587 (N_1587,N_1422,N_1458);
nand U1588 (N_1588,N_1479,N_1482);
or U1589 (N_1589,N_1405,N_1458);
or U1590 (N_1590,N_1415,N_1477);
or U1591 (N_1591,N_1435,N_1481);
or U1592 (N_1592,N_1460,N_1435);
and U1593 (N_1593,N_1455,N_1450);
nor U1594 (N_1594,N_1481,N_1476);
nand U1595 (N_1595,N_1415,N_1479);
nand U1596 (N_1596,N_1487,N_1471);
or U1597 (N_1597,N_1478,N_1416);
and U1598 (N_1598,N_1407,N_1486);
nand U1599 (N_1599,N_1449,N_1470);
or U1600 (N_1600,N_1533,N_1537);
nand U1601 (N_1601,N_1561,N_1586);
nor U1602 (N_1602,N_1535,N_1552);
nand U1603 (N_1603,N_1587,N_1572);
or U1604 (N_1604,N_1526,N_1544);
and U1605 (N_1605,N_1527,N_1545);
and U1606 (N_1606,N_1588,N_1574);
nand U1607 (N_1607,N_1540,N_1518);
nand U1608 (N_1608,N_1560,N_1542);
nand U1609 (N_1609,N_1551,N_1503);
and U1610 (N_1610,N_1510,N_1534);
nor U1611 (N_1611,N_1570,N_1531);
xor U1612 (N_1612,N_1591,N_1549);
nor U1613 (N_1613,N_1564,N_1559);
nand U1614 (N_1614,N_1541,N_1562);
or U1615 (N_1615,N_1543,N_1505);
nand U1616 (N_1616,N_1500,N_1528);
nor U1617 (N_1617,N_1585,N_1512);
nor U1618 (N_1618,N_1556,N_1536);
and U1619 (N_1619,N_1599,N_1568);
and U1620 (N_1620,N_1558,N_1565);
or U1621 (N_1621,N_1519,N_1594);
or U1622 (N_1622,N_1515,N_1567);
or U1623 (N_1623,N_1555,N_1569);
and U1624 (N_1624,N_1516,N_1554);
nor U1625 (N_1625,N_1580,N_1584);
nand U1626 (N_1626,N_1563,N_1547);
nand U1627 (N_1627,N_1538,N_1507);
xor U1628 (N_1628,N_1532,N_1597);
nand U1629 (N_1629,N_1546,N_1504);
and U1630 (N_1630,N_1509,N_1598);
nor U1631 (N_1631,N_1539,N_1596);
and U1632 (N_1632,N_1576,N_1511);
nor U1633 (N_1633,N_1514,N_1522);
or U1634 (N_1634,N_1583,N_1550);
nor U1635 (N_1635,N_1517,N_1578);
nor U1636 (N_1636,N_1593,N_1521);
and U1637 (N_1637,N_1595,N_1502);
nor U1638 (N_1638,N_1525,N_1566);
and U1639 (N_1639,N_1592,N_1506);
or U1640 (N_1640,N_1548,N_1557);
and U1641 (N_1641,N_1523,N_1573);
nor U1642 (N_1642,N_1581,N_1520);
or U1643 (N_1643,N_1513,N_1553);
nor U1644 (N_1644,N_1524,N_1579);
nand U1645 (N_1645,N_1501,N_1508);
nand U1646 (N_1646,N_1589,N_1582);
or U1647 (N_1647,N_1575,N_1577);
nand U1648 (N_1648,N_1590,N_1529);
or U1649 (N_1649,N_1530,N_1571);
nor U1650 (N_1650,N_1528,N_1549);
nor U1651 (N_1651,N_1585,N_1559);
and U1652 (N_1652,N_1542,N_1537);
nand U1653 (N_1653,N_1590,N_1518);
nand U1654 (N_1654,N_1554,N_1599);
nand U1655 (N_1655,N_1582,N_1520);
and U1656 (N_1656,N_1512,N_1552);
or U1657 (N_1657,N_1556,N_1563);
nor U1658 (N_1658,N_1589,N_1579);
nand U1659 (N_1659,N_1561,N_1575);
or U1660 (N_1660,N_1559,N_1597);
nor U1661 (N_1661,N_1584,N_1535);
and U1662 (N_1662,N_1594,N_1539);
nor U1663 (N_1663,N_1530,N_1508);
nand U1664 (N_1664,N_1574,N_1509);
nand U1665 (N_1665,N_1562,N_1543);
nand U1666 (N_1666,N_1553,N_1557);
or U1667 (N_1667,N_1597,N_1567);
nor U1668 (N_1668,N_1545,N_1534);
nand U1669 (N_1669,N_1576,N_1562);
or U1670 (N_1670,N_1506,N_1573);
nor U1671 (N_1671,N_1522,N_1543);
nor U1672 (N_1672,N_1511,N_1567);
nor U1673 (N_1673,N_1513,N_1598);
xnor U1674 (N_1674,N_1563,N_1523);
nand U1675 (N_1675,N_1535,N_1513);
or U1676 (N_1676,N_1556,N_1597);
or U1677 (N_1677,N_1531,N_1532);
and U1678 (N_1678,N_1593,N_1567);
nand U1679 (N_1679,N_1590,N_1547);
nand U1680 (N_1680,N_1506,N_1576);
nor U1681 (N_1681,N_1534,N_1515);
nand U1682 (N_1682,N_1579,N_1548);
nor U1683 (N_1683,N_1577,N_1507);
or U1684 (N_1684,N_1534,N_1501);
nand U1685 (N_1685,N_1568,N_1589);
nand U1686 (N_1686,N_1565,N_1560);
nor U1687 (N_1687,N_1561,N_1583);
and U1688 (N_1688,N_1582,N_1528);
and U1689 (N_1689,N_1536,N_1552);
and U1690 (N_1690,N_1559,N_1501);
nand U1691 (N_1691,N_1523,N_1594);
or U1692 (N_1692,N_1503,N_1500);
and U1693 (N_1693,N_1526,N_1511);
nand U1694 (N_1694,N_1592,N_1599);
nor U1695 (N_1695,N_1561,N_1507);
or U1696 (N_1696,N_1567,N_1568);
nand U1697 (N_1697,N_1537,N_1532);
nor U1698 (N_1698,N_1520,N_1532);
nor U1699 (N_1699,N_1559,N_1565);
or U1700 (N_1700,N_1601,N_1612);
and U1701 (N_1701,N_1658,N_1674);
or U1702 (N_1702,N_1651,N_1625);
nor U1703 (N_1703,N_1619,N_1662);
and U1704 (N_1704,N_1655,N_1668);
or U1705 (N_1705,N_1606,N_1664);
nand U1706 (N_1706,N_1663,N_1614);
nand U1707 (N_1707,N_1689,N_1621);
and U1708 (N_1708,N_1684,N_1649);
or U1709 (N_1709,N_1670,N_1616);
and U1710 (N_1710,N_1698,N_1696);
or U1711 (N_1711,N_1682,N_1644);
nor U1712 (N_1712,N_1659,N_1678);
nand U1713 (N_1713,N_1694,N_1675);
nor U1714 (N_1714,N_1665,N_1634);
and U1715 (N_1715,N_1691,N_1666);
and U1716 (N_1716,N_1636,N_1650);
and U1717 (N_1717,N_1603,N_1638);
or U1718 (N_1718,N_1692,N_1620);
or U1719 (N_1719,N_1680,N_1607);
nand U1720 (N_1720,N_1640,N_1673);
and U1721 (N_1721,N_1671,N_1669);
and U1722 (N_1722,N_1693,N_1645);
and U1723 (N_1723,N_1629,N_1667);
nand U1724 (N_1724,N_1617,N_1653);
nand U1725 (N_1725,N_1622,N_1641);
or U1726 (N_1726,N_1605,N_1643);
and U1727 (N_1727,N_1626,N_1635);
nand U1728 (N_1728,N_1646,N_1611);
and U1729 (N_1729,N_1627,N_1654);
nand U1730 (N_1730,N_1639,N_1647);
and U1731 (N_1731,N_1683,N_1624);
and U1732 (N_1732,N_1699,N_1628);
nor U1733 (N_1733,N_1676,N_1687);
or U1734 (N_1734,N_1633,N_1602);
or U1735 (N_1735,N_1686,N_1608);
nor U1736 (N_1736,N_1618,N_1632);
and U1737 (N_1737,N_1623,N_1609);
nor U1738 (N_1738,N_1672,N_1690);
nor U1739 (N_1739,N_1610,N_1615);
nand U1740 (N_1740,N_1642,N_1630);
nor U1741 (N_1741,N_1661,N_1660);
and U1742 (N_1742,N_1681,N_1652);
and U1743 (N_1743,N_1697,N_1648);
or U1744 (N_1744,N_1677,N_1657);
nand U1745 (N_1745,N_1637,N_1613);
or U1746 (N_1746,N_1688,N_1685);
or U1747 (N_1747,N_1600,N_1695);
or U1748 (N_1748,N_1656,N_1631);
and U1749 (N_1749,N_1679,N_1604);
nor U1750 (N_1750,N_1665,N_1652);
and U1751 (N_1751,N_1613,N_1617);
nand U1752 (N_1752,N_1617,N_1657);
and U1753 (N_1753,N_1657,N_1698);
nor U1754 (N_1754,N_1622,N_1684);
or U1755 (N_1755,N_1622,N_1600);
nand U1756 (N_1756,N_1669,N_1635);
nor U1757 (N_1757,N_1690,N_1662);
nand U1758 (N_1758,N_1639,N_1619);
nand U1759 (N_1759,N_1665,N_1654);
nor U1760 (N_1760,N_1619,N_1667);
nor U1761 (N_1761,N_1689,N_1686);
or U1762 (N_1762,N_1695,N_1683);
and U1763 (N_1763,N_1641,N_1627);
nand U1764 (N_1764,N_1635,N_1629);
nand U1765 (N_1765,N_1613,N_1614);
or U1766 (N_1766,N_1647,N_1603);
or U1767 (N_1767,N_1677,N_1664);
nor U1768 (N_1768,N_1612,N_1687);
or U1769 (N_1769,N_1627,N_1655);
or U1770 (N_1770,N_1609,N_1687);
or U1771 (N_1771,N_1610,N_1648);
nor U1772 (N_1772,N_1663,N_1690);
or U1773 (N_1773,N_1685,N_1609);
and U1774 (N_1774,N_1698,N_1617);
nand U1775 (N_1775,N_1664,N_1652);
nand U1776 (N_1776,N_1621,N_1675);
and U1777 (N_1777,N_1636,N_1655);
and U1778 (N_1778,N_1695,N_1637);
xor U1779 (N_1779,N_1686,N_1600);
xor U1780 (N_1780,N_1656,N_1614);
or U1781 (N_1781,N_1652,N_1653);
nor U1782 (N_1782,N_1662,N_1655);
or U1783 (N_1783,N_1609,N_1641);
nand U1784 (N_1784,N_1620,N_1610);
and U1785 (N_1785,N_1655,N_1624);
nor U1786 (N_1786,N_1652,N_1614);
and U1787 (N_1787,N_1679,N_1636);
or U1788 (N_1788,N_1628,N_1666);
or U1789 (N_1789,N_1684,N_1624);
and U1790 (N_1790,N_1615,N_1649);
or U1791 (N_1791,N_1618,N_1615);
nor U1792 (N_1792,N_1696,N_1660);
and U1793 (N_1793,N_1681,N_1661);
and U1794 (N_1794,N_1664,N_1691);
nor U1795 (N_1795,N_1669,N_1684);
nor U1796 (N_1796,N_1618,N_1656);
and U1797 (N_1797,N_1642,N_1622);
or U1798 (N_1798,N_1691,N_1677);
nor U1799 (N_1799,N_1680,N_1656);
or U1800 (N_1800,N_1703,N_1733);
and U1801 (N_1801,N_1717,N_1721);
or U1802 (N_1802,N_1759,N_1799);
or U1803 (N_1803,N_1724,N_1773);
nand U1804 (N_1804,N_1719,N_1727);
nor U1805 (N_1805,N_1765,N_1778);
and U1806 (N_1806,N_1742,N_1757);
and U1807 (N_1807,N_1711,N_1755);
or U1808 (N_1808,N_1787,N_1732);
and U1809 (N_1809,N_1739,N_1726);
and U1810 (N_1810,N_1731,N_1709);
nor U1811 (N_1811,N_1798,N_1793);
or U1812 (N_1812,N_1720,N_1725);
or U1813 (N_1813,N_1714,N_1792);
nand U1814 (N_1814,N_1741,N_1769);
or U1815 (N_1815,N_1772,N_1786);
nor U1816 (N_1816,N_1785,N_1788);
or U1817 (N_1817,N_1749,N_1752);
and U1818 (N_1818,N_1723,N_1780);
nand U1819 (N_1819,N_1735,N_1710);
nand U1820 (N_1820,N_1747,N_1761);
and U1821 (N_1821,N_1784,N_1702);
nand U1822 (N_1822,N_1750,N_1771);
or U1823 (N_1823,N_1791,N_1748);
nand U1824 (N_1824,N_1704,N_1753);
and U1825 (N_1825,N_1751,N_1715);
nor U1826 (N_1826,N_1775,N_1796);
nor U1827 (N_1827,N_1743,N_1766);
and U1828 (N_1828,N_1701,N_1740);
nand U1829 (N_1829,N_1707,N_1728);
or U1830 (N_1830,N_1794,N_1734);
nand U1831 (N_1831,N_1718,N_1737);
nand U1832 (N_1832,N_1713,N_1746);
or U1833 (N_1833,N_1779,N_1797);
or U1834 (N_1834,N_1768,N_1763);
and U1835 (N_1835,N_1760,N_1764);
or U1836 (N_1836,N_1782,N_1790);
nor U1837 (N_1837,N_1745,N_1770);
or U1838 (N_1838,N_1783,N_1744);
nor U1839 (N_1839,N_1729,N_1781);
and U1840 (N_1840,N_1706,N_1758);
nor U1841 (N_1841,N_1795,N_1722);
or U1842 (N_1842,N_1762,N_1754);
nor U1843 (N_1843,N_1712,N_1774);
and U1844 (N_1844,N_1767,N_1700);
nor U1845 (N_1845,N_1736,N_1777);
or U1846 (N_1846,N_1738,N_1730);
nand U1847 (N_1847,N_1789,N_1776);
nand U1848 (N_1848,N_1708,N_1716);
and U1849 (N_1849,N_1756,N_1705);
and U1850 (N_1850,N_1763,N_1712);
and U1851 (N_1851,N_1775,N_1734);
or U1852 (N_1852,N_1794,N_1768);
nand U1853 (N_1853,N_1719,N_1722);
nor U1854 (N_1854,N_1748,N_1790);
nand U1855 (N_1855,N_1720,N_1782);
nand U1856 (N_1856,N_1766,N_1750);
nand U1857 (N_1857,N_1718,N_1720);
and U1858 (N_1858,N_1705,N_1741);
nand U1859 (N_1859,N_1759,N_1755);
nor U1860 (N_1860,N_1715,N_1796);
nor U1861 (N_1861,N_1751,N_1708);
nor U1862 (N_1862,N_1702,N_1730);
nor U1863 (N_1863,N_1732,N_1701);
or U1864 (N_1864,N_1785,N_1789);
nor U1865 (N_1865,N_1782,N_1778);
and U1866 (N_1866,N_1767,N_1749);
or U1867 (N_1867,N_1789,N_1732);
or U1868 (N_1868,N_1759,N_1789);
or U1869 (N_1869,N_1713,N_1707);
nand U1870 (N_1870,N_1780,N_1755);
or U1871 (N_1871,N_1702,N_1709);
nand U1872 (N_1872,N_1765,N_1752);
or U1873 (N_1873,N_1757,N_1785);
nand U1874 (N_1874,N_1769,N_1718);
and U1875 (N_1875,N_1731,N_1720);
or U1876 (N_1876,N_1737,N_1723);
nor U1877 (N_1877,N_1746,N_1741);
and U1878 (N_1878,N_1771,N_1772);
and U1879 (N_1879,N_1718,N_1792);
nand U1880 (N_1880,N_1759,N_1728);
and U1881 (N_1881,N_1705,N_1766);
and U1882 (N_1882,N_1714,N_1795);
nand U1883 (N_1883,N_1790,N_1742);
or U1884 (N_1884,N_1720,N_1743);
and U1885 (N_1885,N_1732,N_1751);
or U1886 (N_1886,N_1785,N_1742);
or U1887 (N_1887,N_1763,N_1743);
or U1888 (N_1888,N_1750,N_1759);
or U1889 (N_1889,N_1782,N_1753);
or U1890 (N_1890,N_1750,N_1704);
nor U1891 (N_1891,N_1728,N_1793);
and U1892 (N_1892,N_1718,N_1705);
nor U1893 (N_1893,N_1715,N_1705);
and U1894 (N_1894,N_1703,N_1783);
or U1895 (N_1895,N_1726,N_1736);
nor U1896 (N_1896,N_1798,N_1733);
nand U1897 (N_1897,N_1728,N_1767);
and U1898 (N_1898,N_1763,N_1720);
nor U1899 (N_1899,N_1728,N_1773);
nor U1900 (N_1900,N_1862,N_1883);
nand U1901 (N_1901,N_1836,N_1875);
nand U1902 (N_1902,N_1843,N_1861);
nand U1903 (N_1903,N_1848,N_1867);
or U1904 (N_1904,N_1874,N_1827);
nand U1905 (N_1905,N_1855,N_1898);
and U1906 (N_1906,N_1873,N_1805);
nand U1907 (N_1907,N_1820,N_1870);
and U1908 (N_1908,N_1829,N_1824);
xnor U1909 (N_1909,N_1877,N_1886);
nor U1910 (N_1910,N_1859,N_1895);
and U1911 (N_1911,N_1888,N_1806);
nor U1912 (N_1912,N_1825,N_1852);
nor U1913 (N_1913,N_1822,N_1863);
or U1914 (N_1914,N_1865,N_1838);
nand U1915 (N_1915,N_1834,N_1882);
nor U1916 (N_1916,N_1821,N_1800);
nor U1917 (N_1917,N_1860,N_1845);
or U1918 (N_1918,N_1815,N_1811);
and U1919 (N_1919,N_1828,N_1835);
nand U1920 (N_1920,N_1830,N_1823);
nor U1921 (N_1921,N_1831,N_1819);
nand U1922 (N_1922,N_1872,N_1833);
or U1923 (N_1923,N_1816,N_1808);
nand U1924 (N_1924,N_1891,N_1841);
nor U1925 (N_1925,N_1818,N_1880);
nand U1926 (N_1926,N_1812,N_1817);
or U1927 (N_1927,N_1890,N_1826);
nor U1928 (N_1928,N_1846,N_1858);
nand U1929 (N_1929,N_1804,N_1851);
or U1930 (N_1930,N_1813,N_1840);
nand U1931 (N_1931,N_1837,N_1887);
and U1932 (N_1932,N_1839,N_1885);
and U1933 (N_1933,N_1893,N_1856);
nor U1934 (N_1934,N_1894,N_1802);
nor U1935 (N_1935,N_1853,N_1842);
nand U1936 (N_1936,N_1884,N_1897);
xor U1937 (N_1937,N_1869,N_1832);
or U1938 (N_1938,N_1809,N_1889);
nor U1939 (N_1939,N_1868,N_1864);
nor U1940 (N_1940,N_1899,N_1857);
and U1941 (N_1941,N_1871,N_1866);
or U1942 (N_1942,N_1854,N_1892);
and U1943 (N_1943,N_1878,N_1881);
and U1944 (N_1944,N_1849,N_1876);
and U1945 (N_1945,N_1844,N_1879);
nor U1946 (N_1946,N_1803,N_1801);
nor U1947 (N_1947,N_1814,N_1850);
and U1948 (N_1948,N_1847,N_1810);
and U1949 (N_1949,N_1807,N_1896);
and U1950 (N_1950,N_1883,N_1823);
xnor U1951 (N_1951,N_1890,N_1862);
and U1952 (N_1952,N_1893,N_1853);
nor U1953 (N_1953,N_1811,N_1848);
nand U1954 (N_1954,N_1855,N_1834);
nand U1955 (N_1955,N_1864,N_1845);
or U1956 (N_1956,N_1870,N_1839);
nor U1957 (N_1957,N_1893,N_1894);
and U1958 (N_1958,N_1815,N_1861);
and U1959 (N_1959,N_1862,N_1821);
and U1960 (N_1960,N_1843,N_1872);
nand U1961 (N_1961,N_1846,N_1873);
nand U1962 (N_1962,N_1839,N_1858);
nor U1963 (N_1963,N_1818,N_1826);
nor U1964 (N_1964,N_1806,N_1823);
or U1965 (N_1965,N_1843,N_1800);
and U1966 (N_1966,N_1859,N_1896);
or U1967 (N_1967,N_1821,N_1861);
nand U1968 (N_1968,N_1815,N_1853);
and U1969 (N_1969,N_1877,N_1831);
or U1970 (N_1970,N_1807,N_1858);
nor U1971 (N_1971,N_1802,N_1886);
nor U1972 (N_1972,N_1838,N_1843);
nor U1973 (N_1973,N_1897,N_1868);
and U1974 (N_1974,N_1886,N_1822);
nor U1975 (N_1975,N_1877,N_1891);
nand U1976 (N_1976,N_1810,N_1891);
nand U1977 (N_1977,N_1823,N_1864);
and U1978 (N_1978,N_1881,N_1817);
and U1979 (N_1979,N_1841,N_1874);
nand U1980 (N_1980,N_1881,N_1875);
and U1981 (N_1981,N_1800,N_1841);
and U1982 (N_1982,N_1821,N_1828);
or U1983 (N_1983,N_1813,N_1838);
or U1984 (N_1984,N_1830,N_1867);
or U1985 (N_1985,N_1865,N_1818);
or U1986 (N_1986,N_1897,N_1866);
nand U1987 (N_1987,N_1825,N_1822);
or U1988 (N_1988,N_1881,N_1845);
nand U1989 (N_1989,N_1875,N_1871);
and U1990 (N_1990,N_1823,N_1844);
nand U1991 (N_1991,N_1864,N_1861);
nand U1992 (N_1992,N_1876,N_1800);
nand U1993 (N_1993,N_1800,N_1835);
nand U1994 (N_1994,N_1877,N_1813);
nor U1995 (N_1995,N_1878,N_1867);
nor U1996 (N_1996,N_1842,N_1832);
or U1997 (N_1997,N_1808,N_1821);
nor U1998 (N_1998,N_1880,N_1899);
nor U1999 (N_1999,N_1851,N_1848);
nand U2000 (N_2000,N_1930,N_1922);
nand U2001 (N_2001,N_1912,N_1965);
or U2002 (N_2002,N_1935,N_1953);
nand U2003 (N_2003,N_1915,N_1990);
or U2004 (N_2004,N_1909,N_1906);
or U2005 (N_2005,N_1975,N_1947);
and U2006 (N_2006,N_1997,N_1927);
and U2007 (N_2007,N_1925,N_1938);
nand U2008 (N_2008,N_1940,N_1928);
nand U2009 (N_2009,N_1900,N_1991);
and U2010 (N_2010,N_1944,N_1985);
nand U2011 (N_2011,N_1974,N_1977);
or U2012 (N_2012,N_1936,N_1968);
nand U2013 (N_2013,N_1932,N_1969);
or U2014 (N_2014,N_1973,N_1995);
or U2015 (N_2015,N_1910,N_1931);
nand U2016 (N_2016,N_1963,N_1978);
and U2017 (N_2017,N_1920,N_1996);
and U2018 (N_2018,N_1946,N_1939);
nand U2019 (N_2019,N_1952,N_1955);
and U2020 (N_2020,N_1913,N_1984);
nor U2021 (N_2021,N_1960,N_1904);
or U2022 (N_2022,N_1901,N_1957);
nor U2023 (N_2023,N_1989,N_1917);
and U2024 (N_2024,N_1980,N_1914);
and U2025 (N_2025,N_1924,N_1971);
and U2026 (N_2026,N_1976,N_1956);
nand U2027 (N_2027,N_1949,N_1923);
or U2028 (N_2028,N_1981,N_1993);
or U2029 (N_2029,N_1903,N_1967);
nor U2030 (N_2030,N_1966,N_1954);
and U2031 (N_2031,N_1992,N_1943);
or U2032 (N_2032,N_1937,N_1986);
and U2033 (N_2033,N_1948,N_1958);
or U2034 (N_2034,N_1970,N_1998);
nand U2035 (N_2035,N_1926,N_1983);
or U2036 (N_2036,N_1964,N_1951);
and U2037 (N_2037,N_1999,N_1921);
and U2038 (N_2038,N_1962,N_1959);
nor U2039 (N_2039,N_1994,N_1950);
or U2040 (N_2040,N_1905,N_1945);
or U2041 (N_2041,N_1929,N_1979);
nand U2042 (N_2042,N_1961,N_1908);
nor U2043 (N_2043,N_1916,N_1988);
and U2044 (N_2044,N_1972,N_1982);
nor U2045 (N_2045,N_1987,N_1933);
nand U2046 (N_2046,N_1902,N_1918);
nand U2047 (N_2047,N_1907,N_1911);
and U2048 (N_2048,N_1942,N_1934);
nand U2049 (N_2049,N_1919,N_1941);
and U2050 (N_2050,N_1951,N_1923);
and U2051 (N_2051,N_1928,N_1955);
nor U2052 (N_2052,N_1947,N_1988);
nor U2053 (N_2053,N_1941,N_1930);
nand U2054 (N_2054,N_1963,N_1942);
or U2055 (N_2055,N_1951,N_1919);
nor U2056 (N_2056,N_1980,N_1939);
nor U2057 (N_2057,N_1906,N_1967);
and U2058 (N_2058,N_1978,N_1923);
nor U2059 (N_2059,N_1980,N_1954);
xnor U2060 (N_2060,N_1977,N_1930);
or U2061 (N_2061,N_1948,N_1921);
nor U2062 (N_2062,N_1918,N_1988);
and U2063 (N_2063,N_1941,N_1905);
nand U2064 (N_2064,N_1938,N_1987);
nor U2065 (N_2065,N_1987,N_1929);
nor U2066 (N_2066,N_1931,N_1988);
nand U2067 (N_2067,N_1918,N_1906);
or U2068 (N_2068,N_1919,N_1961);
or U2069 (N_2069,N_1903,N_1995);
nor U2070 (N_2070,N_1950,N_1914);
nor U2071 (N_2071,N_1904,N_1990);
or U2072 (N_2072,N_1960,N_1948);
and U2073 (N_2073,N_1919,N_1939);
xnor U2074 (N_2074,N_1942,N_1993);
or U2075 (N_2075,N_1920,N_1955);
or U2076 (N_2076,N_1935,N_1968);
or U2077 (N_2077,N_1920,N_1987);
or U2078 (N_2078,N_1911,N_1988);
and U2079 (N_2079,N_1918,N_1929);
nor U2080 (N_2080,N_1987,N_1954);
and U2081 (N_2081,N_1994,N_1957);
nor U2082 (N_2082,N_1927,N_1905);
or U2083 (N_2083,N_1962,N_1906);
and U2084 (N_2084,N_1967,N_1932);
or U2085 (N_2085,N_1901,N_1942);
nor U2086 (N_2086,N_1929,N_1973);
and U2087 (N_2087,N_1976,N_1915);
or U2088 (N_2088,N_1923,N_1932);
or U2089 (N_2089,N_1973,N_1972);
and U2090 (N_2090,N_1969,N_1920);
nand U2091 (N_2091,N_1963,N_1980);
nand U2092 (N_2092,N_1941,N_1995);
or U2093 (N_2093,N_1934,N_1970);
nand U2094 (N_2094,N_1962,N_1914);
nand U2095 (N_2095,N_1951,N_1986);
nor U2096 (N_2096,N_1916,N_1917);
or U2097 (N_2097,N_1957,N_1979);
and U2098 (N_2098,N_1957,N_1982);
nand U2099 (N_2099,N_1975,N_1946);
and U2100 (N_2100,N_2016,N_2094);
or U2101 (N_2101,N_2009,N_2048);
nor U2102 (N_2102,N_2095,N_2057);
and U2103 (N_2103,N_2033,N_2015);
and U2104 (N_2104,N_2055,N_2061);
and U2105 (N_2105,N_2064,N_2082);
or U2106 (N_2106,N_2000,N_2078);
or U2107 (N_2107,N_2014,N_2020);
or U2108 (N_2108,N_2066,N_2012);
or U2109 (N_2109,N_2073,N_2038);
or U2110 (N_2110,N_2005,N_2096);
or U2111 (N_2111,N_2086,N_2004);
nor U2112 (N_2112,N_2056,N_2010);
and U2113 (N_2113,N_2068,N_2027);
and U2114 (N_2114,N_2025,N_2062);
xnor U2115 (N_2115,N_2051,N_2060);
nand U2116 (N_2116,N_2070,N_2074);
nor U2117 (N_2117,N_2002,N_2099);
and U2118 (N_2118,N_2089,N_2067);
and U2119 (N_2119,N_2030,N_2008);
nand U2120 (N_2120,N_2052,N_2037);
or U2121 (N_2121,N_2084,N_2026);
and U2122 (N_2122,N_2080,N_2053);
nand U2123 (N_2123,N_2085,N_2072);
and U2124 (N_2124,N_2079,N_2097);
nor U2125 (N_2125,N_2003,N_2077);
nor U2126 (N_2126,N_2045,N_2034);
and U2127 (N_2127,N_2071,N_2087);
nand U2128 (N_2128,N_2031,N_2023);
nand U2129 (N_2129,N_2040,N_2006);
or U2130 (N_2130,N_2001,N_2090);
and U2131 (N_2131,N_2039,N_2019);
or U2132 (N_2132,N_2024,N_2044);
nand U2133 (N_2133,N_2065,N_2063);
nor U2134 (N_2134,N_2083,N_2098);
nand U2135 (N_2135,N_2028,N_2050);
or U2136 (N_2136,N_2088,N_2054);
and U2137 (N_2137,N_2093,N_2081);
and U2138 (N_2138,N_2022,N_2018);
nor U2139 (N_2139,N_2076,N_2091);
or U2140 (N_2140,N_2011,N_2092);
nor U2141 (N_2141,N_2035,N_2013);
or U2142 (N_2142,N_2017,N_2047);
and U2143 (N_2143,N_2049,N_2041);
nor U2144 (N_2144,N_2042,N_2021);
or U2145 (N_2145,N_2046,N_2059);
nor U2146 (N_2146,N_2069,N_2036);
nor U2147 (N_2147,N_2043,N_2058);
nand U2148 (N_2148,N_2029,N_2007);
nand U2149 (N_2149,N_2032,N_2075);
nand U2150 (N_2150,N_2078,N_2003);
or U2151 (N_2151,N_2097,N_2065);
and U2152 (N_2152,N_2061,N_2076);
nand U2153 (N_2153,N_2095,N_2084);
nand U2154 (N_2154,N_2035,N_2089);
and U2155 (N_2155,N_2044,N_2089);
and U2156 (N_2156,N_2052,N_2057);
and U2157 (N_2157,N_2046,N_2038);
and U2158 (N_2158,N_2071,N_2068);
nor U2159 (N_2159,N_2085,N_2082);
or U2160 (N_2160,N_2084,N_2061);
nand U2161 (N_2161,N_2013,N_2096);
and U2162 (N_2162,N_2091,N_2044);
nor U2163 (N_2163,N_2090,N_2048);
or U2164 (N_2164,N_2061,N_2092);
nand U2165 (N_2165,N_2081,N_2038);
and U2166 (N_2166,N_2066,N_2092);
nor U2167 (N_2167,N_2081,N_2011);
or U2168 (N_2168,N_2056,N_2099);
and U2169 (N_2169,N_2058,N_2086);
or U2170 (N_2170,N_2087,N_2091);
nor U2171 (N_2171,N_2088,N_2085);
nand U2172 (N_2172,N_2072,N_2015);
or U2173 (N_2173,N_2093,N_2023);
or U2174 (N_2174,N_2049,N_2083);
or U2175 (N_2175,N_2086,N_2036);
or U2176 (N_2176,N_2097,N_2024);
and U2177 (N_2177,N_2033,N_2077);
or U2178 (N_2178,N_2066,N_2097);
or U2179 (N_2179,N_2065,N_2042);
nand U2180 (N_2180,N_2002,N_2035);
nand U2181 (N_2181,N_2073,N_2015);
nor U2182 (N_2182,N_2092,N_2024);
or U2183 (N_2183,N_2079,N_2022);
nor U2184 (N_2184,N_2095,N_2047);
or U2185 (N_2185,N_2060,N_2028);
nor U2186 (N_2186,N_2009,N_2064);
nand U2187 (N_2187,N_2038,N_2035);
nand U2188 (N_2188,N_2044,N_2096);
nor U2189 (N_2189,N_2040,N_2093);
nor U2190 (N_2190,N_2078,N_2085);
nand U2191 (N_2191,N_2060,N_2013);
and U2192 (N_2192,N_2069,N_2006);
nor U2193 (N_2193,N_2046,N_2057);
nand U2194 (N_2194,N_2073,N_2025);
nand U2195 (N_2195,N_2005,N_2091);
nor U2196 (N_2196,N_2082,N_2029);
nand U2197 (N_2197,N_2062,N_2031);
and U2198 (N_2198,N_2023,N_2043);
nor U2199 (N_2199,N_2098,N_2024);
nand U2200 (N_2200,N_2140,N_2174);
nand U2201 (N_2201,N_2194,N_2164);
nor U2202 (N_2202,N_2185,N_2195);
or U2203 (N_2203,N_2112,N_2139);
nand U2204 (N_2204,N_2134,N_2110);
nand U2205 (N_2205,N_2127,N_2189);
nand U2206 (N_2206,N_2183,N_2177);
nor U2207 (N_2207,N_2151,N_2113);
nor U2208 (N_2208,N_2136,N_2150);
nor U2209 (N_2209,N_2104,N_2111);
nand U2210 (N_2210,N_2123,N_2148);
nor U2211 (N_2211,N_2184,N_2199);
nand U2212 (N_2212,N_2105,N_2130);
nand U2213 (N_2213,N_2131,N_2168);
nor U2214 (N_2214,N_2192,N_2107);
and U2215 (N_2215,N_2138,N_2157);
nand U2216 (N_2216,N_2182,N_2135);
nand U2217 (N_2217,N_2114,N_2142);
nand U2218 (N_2218,N_2162,N_2197);
and U2219 (N_2219,N_2149,N_2180);
or U2220 (N_2220,N_2143,N_2120);
nand U2221 (N_2221,N_2145,N_2124);
nor U2222 (N_2222,N_2158,N_2161);
nand U2223 (N_2223,N_2196,N_2193);
or U2224 (N_2224,N_2159,N_2115);
nand U2225 (N_2225,N_2163,N_2137);
nor U2226 (N_2226,N_2147,N_2106);
nand U2227 (N_2227,N_2165,N_2128);
and U2228 (N_2228,N_2198,N_2155);
or U2229 (N_2229,N_2103,N_2172);
or U2230 (N_2230,N_2191,N_2176);
nand U2231 (N_2231,N_2119,N_2133);
nor U2232 (N_2232,N_2146,N_2160);
and U2233 (N_2233,N_2125,N_2188);
or U2234 (N_2234,N_2186,N_2171);
and U2235 (N_2235,N_2175,N_2156);
or U2236 (N_2236,N_2102,N_2178);
nand U2237 (N_2237,N_2132,N_2169);
or U2238 (N_2238,N_2181,N_2121);
and U2239 (N_2239,N_2100,N_2167);
nor U2240 (N_2240,N_2101,N_2118);
nand U2241 (N_2241,N_2152,N_2153);
nor U2242 (N_2242,N_2109,N_2108);
nand U2243 (N_2243,N_2129,N_2126);
and U2244 (N_2244,N_2170,N_2117);
and U2245 (N_2245,N_2154,N_2122);
nand U2246 (N_2246,N_2187,N_2173);
and U2247 (N_2247,N_2179,N_2166);
and U2248 (N_2248,N_2144,N_2190);
and U2249 (N_2249,N_2116,N_2141);
or U2250 (N_2250,N_2192,N_2178);
nand U2251 (N_2251,N_2148,N_2146);
or U2252 (N_2252,N_2191,N_2167);
nand U2253 (N_2253,N_2103,N_2190);
nand U2254 (N_2254,N_2122,N_2141);
and U2255 (N_2255,N_2143,N_2111);
nor U2256 (N_2256,N_2177,N_2175);
nand U2257 (N_2257,N_2105,N_2172);
and U2258 (N_2258,N_2187,N_2167);
nor U2259 (N_2259,N_2179,N_2113);
nor U2260 (N_2260,N_2122,N_2162);
or U2261 (N_2261,N_2165,N_2198);
nand U2262 (N_2262,N_2138,N_2127);
nand U2263 (N_2263,N_2137,N_2132);
or U2264 (N_2264,N_2183,N_2188);
nand U2265 (N_2265,N_2186,N_2137);
nor U2266 (N_2266,N_2109,N_2168);
xor U2267 (N_2267,N_2115,N_2176);
and U2268 (N_2268,N_2100,N_2148);
or U2269 (N_2269,N_2146,N_2159);
and U2270 (N_2270,N_2126,N_2102);
or U2271 (N_2271,N_2141,N_2188);
or U2272 (N_2272,N_2141,N_2112);
and U2273 (N_2273,N_2162,N_2195);
or U2274 (N_2274,N_2192,N_2113);
xnor U2275 (N_2275,N_2105,N_2147);
nor U2276 (N_2276,N_2104,N_2183);
nor U2277 (N_2277,N_2141,N_2173);
or U2278 (N_2278,N_2103,N_2108);
nor U2279 (N_2279,N_2164,N_2181);
and U2280 (N_2280,N_2156,N_2167);
nand U2281 (N_2281,N_2131,N_2143);
nand U2282 (N_2282,N_2156,N_2177);
or U2283 (N_2283,N_2133,N_2154);
or U2284 (N_2284,N_2196,N_2122);
and U2285 (N_2285,N_2186,N_2177);
or U2286 (N_2286,N_2175,N_2166);
or U2287 (N_2287,N_2115,N_2134);
nand U2288 (N_2288,N_2165,N_2105);
nand U2289 (N_2289,N_2143,N_2166);
and U2290 (N_2290,N_2120,N_2164);
nor U2291 (N_2291,N_2129,N_2168);
or U2292 (N_2292,N_2116,N_2158);
or U2293 (N_2293,N_2137,N_2181);
nand U2294 (N_2294,N_2180,N_2143);
or U2295 (N_2295,N_2147,N_2151);
or U2296 (N_2296,N_2168,N_2171);
and U2297 (N_2297,N_2121,N_2109);
nor U2298 (N_2298,N_2109,N_2179);
nand U2299 (N_2299,N_2182,N_2137);
and U2300 (N_2300,N_2248,N_2269);
nor U2301 (N_2301,N_2247,N_2256);
nor U2302 (N_2302,N_2284,N_2278);
nor U2303 (N_2303,N_2208,N_2283);
or U2304 (N_2304,N_2280,N_2219);
nand U2305 (N_2305,N_2209,N_2220);
nand U2306 (N_2306,N_2287,N_2265);
xnor U2307 (N_2307,N_2236,N_2207);
or U2308 (N_2308,N_2254,N_2275);
nand U2309 (N_2309,N_2279,N_2217);
nand U2310 (N_2310,N_2292,N_2218);
nor U2311 (N_2311,N_2250,N_2221);
and U2312 (N_2312,N_2224,N_2252);
nor U2313 (N_2313,N_2214,N_2237);
nand U2314 (N_2314,N_2274,N_2238);
nor U2315 (N_2315,N_2294,N_2210);
nand U2316 (N_2316,N_2233,N_2249);
nand U2317 (N_2317,N_2272,N_2228);
and U2318 (N_2318,N_2293,N_2245);
nor U2319 (N_2319,N_2216,N_2258);
xnor U2320 (N_2320,N_2268,N_2277);
nor U2321 (N_2321,N_2215,N_2282);
nor U2322 (N_2322,N_2295,N_2200);
nor U2323 (N_2323,N_2227,N_2232);
nor U2324 (N_2324,N_2264,N_2203);
or U2325 (N_2325,N_2212,N_2235);
and U2326 (N_2326,N_2225,N_2204);
or U2327 (N_2327,N_2226,N_2260);
and U2328 (N_2328,N_2262,N_2271);
nand U2329 (N_2329,N_2298,N_2261);
nand U2330 (N_2330,N_2273,N_2299);
nor U2331 (N_2331,N_2296,N_2206);
nand U2332 (N_2332,N_2297,N_2255);
nand U2333 (N_2333,N_2263,N_2288);
nand U2334 (N_2334,N_2201,N_2257);
and U2335 (N_2335,N_2285,N_2239);
nand U2336 (N_2336,N_2289,N_2222);
or U2337 (N_2337,N_2259,N_2281);
or U2338 (N_2338,N_2223,N_2246);
and U2339 (N_2339,N_2242,N_2234);
xnor U2340 (N_2340,N_2290,N_2266);
nand U2341 (N_2341,N_2244,N_2251);
or U2342 (N_2342,N_2202,N_2211);
xnor U2343 (N_2343,N_2229,N_2230);
nand U2344 (N_2344,N_2231,N_2243);
or U2345 (N_2345,N_2267,N_2205);
nor U2346 (N_2346,N_2213,N_2276);
or U2347 (N_2347,N_2240,N_2291);
nand U2348 (N_2348,N_2253,N_2286);
xnor U2349 (N_2349,N_2270,N_2241);
or U2350 (N_2350,N_2201,N_2253);
and U2351 (N_2351,N_2253,N_2217);
or U2352 (N_2352,N_2215,N_2294);
or U2353 (N_2353,N_2227,N_2203);
or U2354 (N_2354,N_2204,N_2236);
and U2355 (N_2355,N_2251,N_2289);
and U2356 (N_2356,N_2231,N_2296);
nor U2357 (N_2357,N_2275,N_2201);
nand U2358 (N_2358,N_2231,N_2221);
xnor U2359 (N_2359,N_2295,N_2219);
nor U2360 (N_2360,N_2226,N_2280);
and U2361 (N_2361,N_2265,N_2214);
or U2362 (N_2362,N_2295,N_2278);
nor U2363 (N_2363,N_2201,N_2263);
or U2364 (N_2364,N_2297,N_2248);
nand U2365 (N_2365,N_2212,N_2243);
and U2366 (N_2366,N_2236,N_2237);
and U2367 (N_2367,N_2200,N_2210);
nand U2368 (N_2368,N_2284,N_2253);
nor U2369 (N_2369,N_2281,N_2235);
nand U2370 (N_2370,N_2274,N_2295);
nand U2371 (N_2371,N_2203,N_2212);
nor U2372 (N_2372,N_2283,N_2292);
or U2373 (N_2373,N_2282,N_2247);
or U2374 (N_2374,N_2289,N_2202);
and U2375 (N_2375,N_2221,N_2217);
and U2376 (N_2376,N_2206,N_2243);
nand U2377 (N_2377,N_2299,N_2230);
nand U2378 (N_2378,N_2289,N_2223);
nor U2379 (N_2379,N_2280,N_2288);
and U2380 (N_2380,N_2294,N_2217);
nand U2381 (N_2381,N_2243,N_2259);
and U2382 (N_2382,N_2295,N_2221);
and U2383 (N_2383,N_2249,N_2268);
and U2384 (N_2384,N_2232,N_2286);
or U2385 (N_2385,N_2227,N_2216);
nand U2386 (N_2386,N_2256,N_2217);
nor U2387 (N_2387,N_2213,N_2273);
or U2388 (N_2388,N_2226,N_2219);
and U2389 (N_2389,N_2283,N_2224);
or U2390 (N_2390,N_2217,N_2297);
and U2391 (N_2391,N_2241,N_2225);
and U2392 (N_2392,N_2242,N_2278);
nor U2393 (N_2393,N_2212,N_2214);
or U2394 (N_2394,N_2251,N_2236);
and U2395 (N_2395,N_2285,N_2291);
nand U2396 (N_2396,N_2211,N_2212);
or U2397 (N_2397,N_2208,N_2205);
nand U2398 (N_2398,N_2201,N_2255);
and U2399 (N_2399,N_2243,N_2201);
nor U2400 (N_2400,N_2301,N_2307);
or U2401 (N_2401,N_2329,N_2386);
xnor U2402 (N_2402,N_2357,N_2385);
nand U2403 (N_2403,N_2393,N_2394);
nand U2404 (N_2404,N_2303,N_2358);
and U2405 (N_2405,N_2323,N_2353);
nand U2406 (N_2406,N_2354,N_2343);
and U2407 (N_2407,N_2372,N_2352);
or U2408 (N_2408,N_2334,N_2336);
or U2409 (N_2409,N_2317,N_2362);
nand U2410 (N_2410,N_2322,N_2383);
nand U2411 (N_2411,N_2346,N_2309);
or U2412 (N_2412,N_2369,N_2398);
or U2413 (N_2413,N_2318,N_2375);
and U2414 (N_2414,N_2349,N_2345);
and U2415 (N_2415,N_2364,N_2304);
and U2416 (N_2416,N_2337,N_2340);
and U2417 (N_2417,N_2348,N_2305);
nor U2418 (N_2418,N_2397,N_2373);
nand U2419 (N_2419,N_2377,N_2300);
or U2420 (N_2420,N_2399,N_2368);
nand U2421 (N_2421,N_2321,N_2366);
nor U2422 (N_2422,N_2351,N_2382);
nor U2423 (N_2423,N_2314,N_2316);
and U2424 (N_2424,N_2396,N_2313);
or U2425 (N_2425,N_2356,N_2389);
nor U2426 (N_2426,N_2361,N_2315);
nor U2427 (N_2427,N_2302,N_2319);
nand U2428 (N_2428,N_2387,N_2331);
and U2429 (N_2429,N_2350,N_2376);
or U2430 (N_2430,N_2347,N_2371);
nand U2431 (N_2431,N_2360,N_2311);
or U2432 (N_2432,N_2355,N_2379);
and U2433 (N_2433,N_2365,N_2330);
and U2434 (N_2434,N_2339,N_2328);
and U2435 (N_2435,N_2370,N_2312);
nor U2436 (N_2436,N_2335,N_2326);
or U2437 (N_2437,N_2388,N_2324);
nand U2438 (N_2438,N_2320,N_2367);
nor U2439 (N_2439,N_2378,N_2308);
nor U2440 (N_2440,N_2327,N_2381);
or U2441 (N_2441,N_2338,N_2380);
nand U2442 (N_2442,N_2333,N_2359);
nor U2443 (N_2443,N_2374,N_2392);
or U2444 (N_2444,N_2344,N_2306);
and U2445 (N_2445,N_2384,N_2390);
nand U2446 (N_2446,N_2332,N_2363);
and U2447 (N_2447,N_2391,N_2342);
and U2448 (N_2448,N_2325,N_2341);
and U2449 (N_2449,N_2310,N_2395);
or U2450 (N_2450,N_2319,N_2390);
nor U2451 (N_2451,N_2347,N_2399);
or U2452 (N_2452,N_2373,N_2300);
nand U2453 (N_2453,N_2308,N_2377);
or U2454 (N_2454,N_2318,N_2378);
or U2455 (N_2455,N_2321,N_2313);
nor U2456 (N_2456,N_2388,N_2319);
and U2457 (N_2457,N_2307,N_2321);
nor U2458 (N_2458,N_2377,N_2321);
nor U2459 (N_2459,N_2317,N_2324);
nand U2460 (N_2460,N_2359,N_2301);
or U2461 (N_2461,N_2399,N_2363);
or U2462 (N_2462,N_2315,N_2345);
or U2463 (N_2463,N_2360,N_2344);
xor U2464 (N_2464,N_2345,N_2320);
nor U2465 (N_2465,N_2359,N_2386);
nand U2466 (N_2466,N_2367,N_2354);
nand U2467 (N_2467,N_2391,N_2340);
nand U2468 (N_2468,N_2318,N_2379);
nor U2469 (N_2469,N_2339,N_2389);
and U2470 (N_2470,N_2350,N_2371);
nor U2471 (N_2471,N_2399,N_2359);
or U2472 (N_2472,N_2383,N_2389);
nor U2473 (N_2473,N_2320,N_2366);
nor U2474 (N_2474,N_2361,N_2340);
nand U2475 (N_2475,N_2334,N_2321);
nor U2476 (N_2476,N_2306,N_2373);
nand U2477 (N_2477,N_2381,N_2331);
and U2478 (N_2478,N_2300,N_2369);
or U2479 (N_2479,N_2322,N_2374);
nand U2480 (N_2480,N_2334,N_2302);
or U2481 (N_2481,N_2381,N_2391);
nand U2482 (N_2482,N_2304,N_2305);
or U2483 (N_2483,N_2307,N_2308);
or U2484 (N_2484,N_2327,N_2324);
nand U2485 (N_2485,N_2300,N_2374);
nor U2486 (N_2486,N_2326,N_2384);
or U2487 (N_2487,N_2370,N_2377);
or U2488 (N_2488,N_2310,N_2384);
or U2489 (N_2489,N_2308,N_2364);
nor U2490 (N_2490,N_2314,N_2346);
nor U2491 (N_2491,N_2362,N_2312);
nand U2492 (N_2492,N_2311,N_2367);
nor U2493 (N_2493,N_2324,N_2350);
or U2494 (N_2494,N_2355,N_2350);
nor U2495 (N_2495,N_2316,N_2389);
nand U2496 (N_2496,N_2314,N_2332);
and U2497 (N_2497,N_2307,N_2375);
or U2498 (N_2498,N_2307,N_2360);
nand U2499 (N_2499,N_2323,N_2365);
and U2500 (N_2500,N_2454,N_2457);
nand U2501 (N_2501,N_2402,N_2436);
nor U2502 (N_2502,N_2491,N_2428);
nor U2503 (N_2503,N_2403,N_2440);
nand U2504 (N_2504,N_2483,N_2479);
nand U2505 (N_2505,N_2486,N_2473);
nand U2506 (N_2506,N_2418,N_2496);
and U2507 (N_2507,N_2492,N_2443);
or U2508 (N_2508,N_2467,N_2476);
nor U2509 (N_2509,N_2499,N_2448);
or U2510 (N_2510,N_2433,N_2409);
and U2511 (N_2511,N_2485,N_2438);
nor U2512 (N_2512,N_2480,N_2431);
nor U2513 (N_2513,N_2465,N_2498);
nor U2514 (N_2514,N_2422,N_2429);
or U2515 (N_2515,N_2416,N_2413);
nor U2516 (N_2516,N_2463,N_2456);
or U2517 (N_2517,N_2453,N_2468);
or U2518 (N_2518,N_2478,N_2464);
or U2519 (N_2519,N_2441,N_2445);
or U2520 (N_2520,N_2414,N_2482);
nor U2521 (N_2521,N_2420,N_2439);
and U2522 (N_2522,N_2458,N_2462);
nor U2523 (N_2523,N_2430,N_2469);
or U2524 (N_2524,N_2407,N_2446);
nor U2525 (N_2525,N_2427,N_2444);
nor U2526 (N_2526,N_2424,N_2461);
or U2527 (N_2527,N_2406,N_2459);
and U2528 (N_2528,N_2415,N_2447);
and U2529 (N_2529,N_2472,N_2497);
nor U2530 (N_2530,N_2425,N_2450);
or U2531 (N_2531,N_2452,N_2495);
or U2532 (N_2532,N_2451,N_2419);
nor U2533 (N_2533,N_2404,N_2437);
or U2534 (N_2534,N_2449,N_2426);
or U2535 (N_2535,N_2408,N_2410);
nor U2536 (N_2536,N_2417,N_2494);
or U2537 (N_2537,N_2477,N_2484);
or U2538 (N_2538,N_2432,N_2442);
nand U2539 (N_2539,N_2466,N_2470);
nand U2540 (N_2540,N_2489,N_2412);
or U2541 (N_2541,N_2400,N_2488);
or U2542 (N_2542,N_2471,N_2401);
nand U2543 (N_2543,N_2435,N_2460);
nand U2544 (N_2544,N_2434,N_2481);
or U2545 (N_2545,N_2490,N_2411);
and U2546 (N_2546,N_2421,N_2455);
nor U2547 (N_2547,N_2474,N_2475);
or U2548 (N_2548,N_2405,N_2423);
or U2549 (N_2549,N_2493,N_2487);
or U2550 (N_2550,N_2436,N_2460);
nand U2551 (N_2551,N_2496,N_2454);
nor U2552 (N_2552,N_2431,N_2432);
nand U2553 (N_2553,N_2402,N_2497);
nand U2554 (N_2554,N_2455,N_2401);
nor U2555 (N_2555,N_2434,N_2429);
or U2556 (N_2556,N_2413,N_2498);
or U2557 (N_2557,N_2400,N_2426);
or U2558 (N_2558,N_2492,N_2483);
or U2559 (N_2559,N_2461,N_2492);
nor U2560 (N_2560,N_2420,N_2434);
and U2561 (N_2561,N_2438,N_2469);
or U2562 (N_2562,N_2468,N_2487);
and U2563 (N_2563,N_2460,N_2433);
nand U2564 (N_2564,N_2464,N_2413);
and U2565 (N_2565,N_2400,N_2419);
nand U2566 (N_2566,N_2405,N_2457);
and U2567 (N_2567,N_2453,N_2444);
or U2568 (N_2568,N_2415,N_2484);
and U2569 (N_2569,N_2482,N_2481);
or U2570 (N_2570,N_2419,N_2424);
and U2571 (N_2571,N_2445,N_2434);
nor U2572 (N_2572,N_2457,N_2497);
nand U2573 (N_2573,N_2407,N_2400);
or U2574 (N_2574,N_2452,N_2449);
or U2575 (N_2575,N_2482,N_2499);
and U2576 (N_2576,N_2465,N_2416);
nor U2577 (N_2577,N_2470,N_2442);
nand U2578 (N_2578,N_2440,N_2428);
or U2579 (N_2579,N_2417,N_2426);
nor U2580 (N_2580,N_2482,N_2456);
and U2581 (N_2581,N_2401,N_2472);
nand U2582 (N_2582,N_2484,N_2461);
nand U2583 (N_2583,N_2432,N_2490);
or U2584 (N_2584,N_2493,N_2475);
and U2585 (N_2585,N_2437,N_2469);
nand U2586 (N_2586,N_2499,N_2445);
nand U2587 (N_2587,N_2455,N_2429);
nand U2588 (N_2588,N_2466,N_2437);
nor U2589 (N_2589,N_2446,N_2423);
nand U2590 (N_2590,N_2474,N_2478);
or U2591 (N_2591,N_2458,N_2489);
nor U2592 (N_2592,N_2485,N_2465);
and U2593 (N_2593,N_2434,N_2428);
and U2594 (N_2594,N_2404,N_2493);
or U2595 (N_2595,N_2426,N_2405);
and U2596 (N_2596,N_2438,N_2426);
and U2597 (N_2597,N_2430,N_2496);
or U2598 (N_2598,N_2486,N_2437);
nor U2599 (N_2599,N_2455,N_2466);
nor U2600 (N_2600,N_2583,N_2544);
or U2601 (N_2601,N_2536,N_2592);
nand U2602 (N_2602,N_2512,N_2567);
nand U2603 (N_2603,N_2515,N_2550);
or U2604 (N_2604,N_2557,N_2559);
and U2605 (N_2605,N_2537,N_2587);
and U2606 (N_2606,N_2520,N_2576);
nor U2607 (N_2607,N_2566,N_2581);
nor U2608 (N_2608,N_2500,N_2516);
or U2609 (N_2609,N_2530,N_2598);
or U2610 (N_2610,N_2506,N_2570);
nor U2611 (N_2611,N_2585,N_2586);
and U2612 (N_2612,N_2501,N_2563);
and U2613 (N_2613,N_2556,N_2577);
nor U2614 (N_2614,N_2525,N_2528);
nor U2615 (N_2615,N_2521,N_2564);
and U2616 (N_2616,N_2542,N_2555);
nor U2617 (N_2617,N_2582,N_2578);
nor U2618 (N_2618,N_2539,N_2510);
and U2619 (N_2619,N_2560,N_2543);
or U2620 (N_2620,N_2511,N_2514);
nand U2621 (N_2621,N_2519,N_2548);
nor U2622 (N_2622,N_2546,N_2529);
nand U2623 (N_2623,N_2505,N_2554);
nor U2624 (N_2624,N_2523,N_2595);
and U2625 (N_2625,N_2562,N_2502);
and U2626 (N_2626,N_2545,N_2534);
nand U2627 (N_2627,N_2517,N_2551);
and U2628 (N_2628,N_2531,N_2599);
nor U2629 (N_2629,N_2532,N_2574);
nor U2630 (N_2630,N_2558,N_2571);
nor U2631 (N_2631,N_2527,N_2573);
or U2632 (N_2632,N_2572,N_2569);
nand U2633 (N_2633,N_2594,N_2580);
and U2634 (N_2634,N_2509,N_2568);
nand U2635 (N_2635,N_2518,N_2524);
and U2636 (N_2636,N_2553,N_2575);
and U2637 (N_2637,N_2547,N_2590);
nor U2638 (N_2638,N_2596,N_2504);
nor U2639 (N_2639,N_2579,N_2584);
nor U2640 (N_2640,N_2503,N_2522);
or U2641 (N_2641,N_2526,N_2541);
or U2642 (N_2642,N_2597,N_2588);
nand U2643 (N_2643,N_2538,N_2507);
nand U2644 (N_2644,N_2513,N_2591);
nor U2645 (N_2645,N_2552,N_2535);
and U2646 (N_2646,N_2589,N_2561);
or U2647 (N_2647,N_2533,N_2549);
nand U2648 (N_2648,N_2565,N_2593);
nor U2649 (N_2649,N_2508,N_2540);
or U2650 (N_2650,N_2530,N_2555);
and U2651 (N_2651,N_2551,N_2577);
nor U2652 (N_2652,N_2518,N_2508);
or U2653 (N_2653,N_2584,N_2557);
and U2654 (N_2654,N_2577,N_2550);
nor U2655 (N_2655,N_2512,N_2504);
and U2656 (N_2656,N_2512,N_2590);
or U2657 (N_2657,N_2502,N_2595);
nand U2658 (N_2658,N_2542,N_2583);
or U2659 (N_2659,N_2595,N_2508);
nor U2660 (N_2660,N_2527,N_2591);
or U2661 (N_2661,N_2545,N_2521);
and U2662 (N_2662,N_2531,N_2538);
nand U2663 (N_2663,N_2532,N_2579);
and U2664 (N_2664,N_2589,N_2534);
nand U2665 (N_2665,N_2501,N_2530);
nor U2666 (N_2666,N_2586,N_2572);
nor U2667 (N_2667,N_2594,N_2592);
and U2668 (N_2668,N_2563,N_2586);
nor U2669 (N_2669,N_2530,N_2517);
nand U2670 (N_2670,N_2540,N_2577);
or U2671 (N_2671,N_2537,N_2590);
nand U2672 (N_2672,N_2548,N_2596);
nor U2673 (N_2673,N_2599,N_2572);
and U2674 (N_2674,N_2593,N_2516);
nand U2675 (N_2675,N_2522,N_2507);
nand U2676 (N_2676,N_2597,N_2568);
and U2677 (N_2677,N_2594,N_2565);
and U2678 (N_2678,N_2559,N_2581);
or U2679 (N_2679,N_2530,N_2584);
nor U2680 (N_2680,N_2557,N_2549);
nor U2681 (N_2681,N_2583,N_2589);
and U2682 (N_2682,N_2550,N_2534);
and U2683 (N_2683,N_2584,N_2535);
or U2684 (N_2684,N_2526,N_2552);
nand U2685 (N_2685,N_2500,N_2557);
nand U2686 (N_2686,N_2519,N_2552);
nor U2687 (N_2687,N_2549,N_2582);
nor U2688 (N_2688,N_2524,N_2508);
nand U2689 (N_2689,N_2542,N_2500);
nand U2690 (N_2690,N_2583,N_2560);
or U2691 (N_2691,N_2587,N_2589);
nor U2692 (N_2692,N_2519,N_2520);
xor U2693 (N_2693,N_2526,N_2597);
or U2694 (N_2694,N_2585,N_2543);
nor U2695 (N_2695,N_2574,N_2592);
nor U2696 (N_2696,N_2534,N_2580);
nor U2697 (N_2697,N_2532,N_2598);
and U2698 (N_2698,N_2565,N_2560);
nor U2699 (N_2699,N_2536,N_2562);
nand U2700 (N_2700,N_2600,N_2691);
or U2701 (N_2701,N_2654,N_2606);
nand U2702 (N_2702,N_2682,N_2672);
and U2703 (N_2703,N_2633,N_2684);
nor U2704 (N_2704,N_2621,N_2693);
or U2705 (N_2705,N_2699,N_2623);
and U2706 (N_2706,N_2686,N_2648);
nor U2707 (N_2707,N_2678,N_2662);
nor U2708 (N_2708,N_2663,N_2629);
nor U2709 (N_2709,N_2624,N_2698);
or U2710 (N_2710,N_2632,N_2634);
and U2711 (N_2711,N_2645,N_2615);
or U2712 (N_2712,N_2692,N_2659);
nand U2713 (N_2713,N_2636,N_2638);
nand U2714 (N_2714,N_2671,N_2697);
nand U2715 (N_2715,N_2655,N_2658);
nand U2716 (N_2716,N_2681,N_2637);
or U2717 (N_2717,N_2687,N_2607);
nor U2718 (N_2718,N_2656,N_2608);
nand U2719 (N_2719,N_2643,N_2685);
nor U2720 (N_2720,N_2676,N_2625);
and U2721 (N_2721,N_2669,N_2642);
or U2722 (N_2722,N_2605,N_2652);
or U2723 (N_2723,N_2666,N_2616);
and U2724 (N_2724,N_2683,N_2626);
nand U2725 (N_2725,N_2618,N_2679);
nor U2726 (N_2726,N_2651,N_2612);
nor U2727 (N_2727,N_2601,N_2639);
or U2728 (N_2728,N_2611,N_2617);
nor U2729 (N_2729,N_2628,N_2604);
nor U2730 (N_2730,N_2640,N_2613);
or U2731 (N_2731,N_2635,N_2664);
nor U2732 (N_2732,N_2647,N_2695);
and U2733 (N_2733,N_2603,N_2630);
nor U2734 (N_2734,N_2631,N_2689);
and U2735 (N_2735,N_2674,N_2649);
nand U2736 (N_2736,N_2602,N_2668);
nand U2737 (N_2737,N_2667,N_2688);
nand U2738 (N_2738,N_2665,N_2653);
nor U2739 (N_2739,N_2660,N_2620);
or U2740 (N_2740,N_2675,N_2609);
and U2741 (N_2741,N_2657,N_2673);
nand U2742 (N_2742,N_2622,N_2650);
nor U2743 (N_2743,N_2619,N_2646);
and U2744 (N_2744,N_2644,N_2614);
nand U2745 (N_2745,N_2696,N_2641);
or U2746 (N_2746,N_2690,N_2627);
nor U2747 (N_2747,N_2610,N_2680);
nand U2748 (N_2748,N_2677,N_2661);
nand U2749 (N_2749,N_2694,N_2670);
nand U2750 (N_2750,N_2646,N_2602);
nand U2751 (N_2751,N_2609,N_2699);
and U2752 (N_2752,N_2689,N_2648);
and U2753 (N_2753,N_2642,N_2601);
nand U2754 (N_2754,N_2644,N_2623);
nand U2755 (N_2755,N_2643,N_2604);
nand U2756 (N_2756,N_2625,N_2615);
nor U2757 (N_2757,N_2652,N_2684);
nand U2758 (N_2758,N_2693,N_2685);
and U2759 (N_2759,N_2642,N_2619);
nand U2760 (N_2760,N_2649,N_2610);
or U2761 (N_2761,N_2694,N_2682);
nand U2762 (N_2762,N_2648,N_2664);
nand U2763 (N_2763,N_2606,N_2634);
or U2764 (N_2764,N_2628,N_2646);
nand U2765 (N_2765,N_2630,N_2619);
nand U2766 (N_2766,N_2607,N_2668);
nand U2767 (N_2767,N_2665,N_2680);
nand U2768 (N_2768,N_2671,N_2610);
and U2769 (N_2769,N_2603,N_2600);
or U2770 (N_2770,N_2648,N_2647);
and U2771 (N_2771,N_2632,N_2683);
or U2772 (N_2772,N_2678,N_2690);
or U2773 (N_2773,N_2650,N_2631);
nor U2774 (N_2774,N_2690,N_2600);
nand U2775 (N_2775,N_2686,N_2636);
nor U2776 (N_2776,N_2693,N_2635);
or U2777 (N_2777,N_2681,N_2610);
and U2778 (N_2778,N_2608,N_2690);
nor U2779 (N_2779,N_2634,N_2642);
nor U2780 (N_2780,N_2680,N_2614);
nand U2781 (N_2781,N_2630,N_2629);
or U2782 (N_2782,N_2692,N_2602);
nor U2783 (N_2783,N_2630,N_2625);
nor U2784 (N_2784,N_2668,N_2640);
nor U2785 (N_2785,N_2635,N_2600);
nor U2786 (N_2786,N_2669,N_2694);
nand U2787 (N_2787,N_2637,N_2624);
nor U2788 (N_2788,N_2650,N_2674);
nor U2789 (N_2789,N_2698,N_2649);
nor U2790 (N_2790,N_2695,N_2676);
nor U2791 (N_2791,N_2621,N_2685);
and U2792 (N_2792,N_2669,N_2689);
nand U2793 (N_2793,N_2611,N_2621);
nand U2794 (N_2794,N_2690,N_2630);
and U2795 (N_2795,N_2678,N_2649);
nor U2796 (N_2796,N_2666,N_2644);
or U2797 (N_2797,N_2644,N_2621);
and U2798 (N_2798,N_2629,N_2604);
nor U2799 (N_2799,N_2633,N_2672);
or U2800 (N_2800,N_2762,N_2739);
xor U2801 (N_2801,N_2759,N_2710);
and U2802 (N_2802,N_2717,N_2789);
and U2803 (N_2803,N_2777,N_2723);
nor U2804 (N_2804,N_2749,N_2796);
nand U2805 (N_2805,N_2728,N_2792);
nand U2806 (N_2806,N_2711,N_2774);
or U2807 (N_2807,N_2736,N_2768);
nand U2808 (N_2808,N_2754,N_2757);
nor U2809 (N_2809,N_2764,N_2729);
nor U2810 (N_2810,N_2761,N_2790);
and U2811 (N_2811,N_2718,N_2779);
nor U2812 (N_2812,N_2724,N_2704);
nand U2813 (N_2813,N_2709,N_2763);
nor U2814 (N_2814,N_2798,N_2776);
nand U2815 (N_2815,N_2791,N_2719);
nor U2816 (N_2816,N_2769,N_2726);
nand U2817 (N_2817,N_2713,N_2773);
nand U2818 (N_2818,N_2738,N_2786);
or U2819 (N_2819,N_2794,N_2727);
and U2820 (N_2820,N_2747,N_2760);
and U2821 (N_2821,N_2756,N_2737);
nor U2822 (N_2822,N_2725,N_2721);
and U2823 (N_2823,N_2788,N_2752);
or U2824 (N_2824,N_2740,N_2782);
nand U2825 (N_2825,N_2732,N_2775);
nand U2826 (N_2826,N_2706,N_2784);
nand U2827 (N_2827,N_2753,N_2778);
and U2828 (N_2828,N_2751,N_2745);
or U2829 (N_2829,N_2731,N_2741);
or U2830 (N_2830,N_2712,N_2730);
nand U2831 (N_2831,N_2714,N_2766);
or U2832 (N_2832,N_2780,N_2702);
nor U2833 (N_2833,N_2748,N_2722);
or U2834 (N_2834,N_2793,N_2771);
and U2835 (N_2835,N_2707,N_2781);
or U2836 (N_2836,N_2705,N_2708);
or U2837 (N_2837,N_2750,N_2772);
and U2838 (N_2838,N_2799,N_2758);
and U2839 (N_2839,N_2795,N_2720);
nor U2840 (N_2840,N_2755,N_2744);
nand U2841 (N_2841,N_2715,N_2770);
or U2842 (N_2842,N_2767,N_2765);
or U2843 (N_2843,N_2785,N_2746);
and U2844 (N_2844,N_2734,N_2701);
nand U2845 (N_2845,N_2743,N_2787);
or U2846 (N_2846,N_2700,N_2742);
nor U2847 (N_2847,N_2797,N_2733);
or U2848 (N_2848,N_2716,N_2735);
nor U2849 (N_2849,N_2783,N_2703);
or U2850 (N_2850,N_2776,N_2706);
or U2851 (N_2851,N_2776,N_2701);
or U2852 (N_2852,N_2787,N_2719);
and U2853 (N_2853,N_2769,N_2780);
or U2854 (N_2854,N_2747,N_2712);
or U2855 (N_2855,N_2767,N_2780);
nor U2856 (N_2856,N_2763,N_2799);
and U2857 (N_2857,N_2785,N_2716);
or U2858 (N_2858,N_2730,N_2722);
or U2859 (N_2859,N_2784,N_2744);
or U2860 (N_2860,N_2781,N_2754);
nor U2861 (N_2861,N_2790,N_2746);
nor U2862 (N_2862,N_2779,N_2790);
nor U2863 (N_2863,N_2716,N_2746);
nand U2864 (N_2864,N_2737,N_2795);
nand U2865 (N_2865,N_2763,N_2732);
or U2866 (N_2866,N_2782,N_2739);
or U2867 (N_2867,N_2731,N_2746);
and U2868 (N_2868,N_2751,N_2795);
nor U2869 (N_2869,N_2726,N_2780);
nand U2870 (N_2870,N_2788,N_2777);
nor U2871 (N_2871,N_2763,N_2736);
and U2872 (N_2872,N_2771,N_2755);
or U2873 (N_2873,N_2790,N_2706);
nand U2874 (N_2874,N_2723,N_2767);
or U2875 (N_2875,N_2700,N_2790);
nor U2876 (N_2876,N_2779,N_2760);
and U2877 (N_2877,N_2736,N_2757);
nand U2878 (N_2878,N_2777,N_2712);
nor U2879 (N_2879,N_2768,N_2785);
nor U2880 (N_2880,N_2789,N_2776);
and U2881 (N_2881,N_2780,N_2732);
nor U2882 (N_2882,N_2794,N_2773);
nand U2883 (N_2883,N_2723,N_2732);
xor U2884 (N_2884,N_2712,N_2711);
and U2885 (N_2885,N_2780,N_2785);
and U2886 (N_2886,N_2767,N_2709);
nor U2887 (N_2887,N_2748,N_2701);
nor U2888 (N_2888,N_2790,N_2718);
nand U2889 (N_2889,N_2791,N_2797);
and U2890 (N_2890,N_2754,N_2733);
or U2891 (N_2891,N_2785,N_2778);
or U2892 (N_2892,N_2712,N_2727);
nor U2893 (N_2893,N_2740,N_2773);
and U2894 (N_2894,N_2762,N_2736);
or U2895 (N_2895,N_2762,N_2748);
nand U2896 (N_2896,N_2706,N_2724);
nor U2897 (N_2897,N_2712,N_2795);
nand U2898 (N_2898,N_2733,N_2709);
nor U2899 (N_2899,N_2760,N_2755);
and U2900 (N_2900,N_2878,N_2815);
and U2901 (N_2901,N_2869,N_2885);
nand U2902 (N_2902,N_2856,N_2814);
nand U2903 (N_2903,N_2887,N_2882);
or U2904 (N_2904,N_2858,N_2894);
nand U2905 (N_2905,N_2861,N_2818);
nand U2906 (N_2906,N_2824,N_2852);
nand U2907 (N_2907,N_2854,N_2823);
nor U2908 (N_2908,N_2893,N_2828);
or U2909 (N_2909,N_2857,N_2866);
nor U2910 (N_2910,N_2889,N_2808);
nand U2911 (N_2911,N_2839,N_2868);
nor U2912 (N_2912,N_2835,N_2846);
or U2913 (N_2913,N_2816,N_2810);
nor U2914 (N_2914,N_2813,N_2825);
or U2915 (N_2915,N_2805,N_2863);
and U2916 (N_2916,N_2832,N_2801);
nor U2917 (N_2917,N_2817,N_2850);
nor U2918 (N_2918,N_2873,N_2862);
nor U2919 (N_2919,N_2870,N_2837);
and U2920 (N_2920,N_2888,N_2822);
nand U2921 (N_2921,N_2860,N_2892);
or U2922 (N_2922,N_2849,N_2895);
and U2923 (N_2923,N_2800,N_2851);
nand U2924 (N_2924,N_2819,N_2836);
or U2925 (N_2925,N_2845,N_2843);
nand U2926 (N_2926,N_2897,N_2871);
nor U2927 (N_2927,N_2834,N_2867);
nor U2928 (N_2928,N_2830,N_2827);
and U2929 (N_2929,N_2886,N_2876);
nand U2930 (N_2930,N_2803,N_2874);
or U2931 (N_2931,N_2865,N_2802);
and U2932 (N_2932,N_2872,N_2807);
nor U2933 (N_2933,N_2821,N_2877);
nand U2934 (N_2934,N_2842,N_2833);
or U2935 (N_2935,N_2855,N_2890);
or U2936 (N_2936,N_2840,N_2881);
and U2937 (N_2937,N_2891,N_2831);
and U2938 (N_2938,N_2811,N_2853);
nand U2939 (N_2939,N_2875,N_2826);
and U2940 (N_2940,N_2844,N_2841);
or U2941 (N_2941,N_2899,N_2838);
nand U2942 (N_2942,N_2809,N_2812);
nor U2943 (N_2943,N_2898,N_2804);
nand U2944 (N_2944,N_2848,N_2859);
nor U2945 (N_2945,N_2820,N_2896);
or U2946 (N_2946,N_2864,N_2879);
and U2947 (N_2947,N_2884,N_2880);
nand U2948 (N_2948,N_2829,N_2883);
and U2949 (N_2949,N_2806,N_2847);
nor U2950 (N_2950,N_2866,N_2854);
and U2951 (N_2951,N_2887,N_2875);
nand U2952 (N_2952,N_2817,N_2811);
nand U2953 (N_2953,N_2812,N_2807);
nor U2954 (N_2954,N_2857,N_2819);
nor U2955 (N_2955,N_2854,N_2819);
and U2956 (N_2956,N_2879,N_2875);
nor U2957 (N_2957,N_2838,N_2885);
nand U2958 (N_2958,N_2870,N_2824);
nor U2959 (N_2959,N_2812,N_2853);
and U2960 (N_2960,N_2889,N_2881);
nand U2961 (N_2961,N_2847,N_2898);
nand U2962 (N_2962,N_2894,N_2803);
and U2963 (N_2963,N_2888,N_2821);
nand U2964 (N_2964,N_2857,N_2862);
and U2965 (N_2965,N_2878,N_2843);
nand U2966 (N_2966,N_2872,N_2817);
nor U2967 (N_2967,N_2849,N_2854);
or U2968 (N_2968,N_2812,N_2838);
or U2969 (N_2969,N_2833,N_2846);
and U2970 (N_2970,N_2870,N_2826);
nand U2971 (N_2971,N_2839,N_2899);
and U2972 (N_2972,N_2885,N_2867);
or U2973 (N_2973,N_2808,N_2847);
nor U2974 (N_2974,N_2814,N_2884);
or U2975 (N_2975,N_2832,N_2893);
and U2976 (N_2976,N_2884,N_2877);
xnor U2977 (N_2977,N_2854,N_2878);
nand U2978 (N_2978,N_2843,N_2899);
nand U2979 (N_2979,N_2846,N_2850);
or U2980 (N_2980,N_2825,N_2856);
or U2981 (N_2981,N_2845,N_2846);
or U2982 (N_2982,N_2854,N_2862);
nor U2983 (N_2983,N_2899,N_2810);
nand U2984 (N_2984,N_2877,N_2880);
nor U2985 (N_2985,N_2848,N_2863);
or U2986 (N_2986,N_2873,N_2838);
nor U2987 (N_2987,N_2824,N_2801);
nand U2988 (N_2988,N_2875,N_2894);
nor U2989 (N_2989,N_2810,N_2884);
nor U2990 (N_2990,N_2875,N_2857);
and U2991 (N_2991,N_2833,N_2847);
nand U2992 (N_2992,N_2877,N_2863);
and U2993 (N_2993,N_2884,N_2893);
or U2994 (N_2994,N_2828,N_2873);
and U2995 (N_2995,N_2896,N_2861);
nor U2996 (N_2996,N_2870,N_2854);
or U2997 (N_2997,N_2867,N_2813);
nand U2998 (N_2998,N_2810,N_2873);
and U2999 (N_2999,N_2831,N_2860);
nand UO_0 (O_0,N_2901,N_2915);
nand UO_1 (O_1,N_2987,N_2977);
nand UO_2 (O_2,N_2902,N_2971);
nor UO_3 (O_3,N_2988,N_2943);
nor UO_4 (O_4,N_2986,N_2990);
nor UO_5 (O_5,N_2912,N_2913);
nand UO_6 (O_6,N_2965,N_2940);
or UO_7 (O_7,N_2951,N_2934);
or UO_8 (O_8,N_2945,N_2952);
nand UO_9 (O_9,N_2947,N_2938);
nor UO_10 (O_10,N_2976,N_2968);
and UO_11 (O_11,N_2981,N_2933);
or UO_12 (O_12,N_2909,N_2979);
nor UO_13 (O_13,N_2972,N_2925);
and UO_14 (O_14,N_2963,N_2926);
nor UO_15 (O_15,N_2959,N_2982);
and UO_16 (O_16,N_2905,N_2932);
nor UO_17 (O_17,N_2962,N_2999);
nor UO_18 (O_18,N_2978,N_2920);
and UO_19 (O_19,N_2991,N_2974);
nand UO_20 (O_20,N_2966,N_2907);
and UO_21 (O_21,N_2914,N_2946);
or UO_22 (O_22,N_2983,N_2930);
or UO_23 (O_23,N_2904,N_2969);
and UO_24 (O_24,N_2906,N_2942);
or UO_25 (O_25,N_2997,N_2924);
xnor UO_26 (O_26,N_2980,N_2957);
nand UO_27 (O_27,N_2948,N_2929);
or UO_28 (O_28,N_2949,N_2960);
nand UO_29 (O_29,N_2916,N_2919);
nor UO_30 (O_30,N_2910,N_2944);
or UO_31 (O_31,N_2975,N_2992);
nor UO_32 (O_32,N_2922,N_2998);
nor UO_33 (O_33,N_2967,N_2918);
nand UO_34 (O_34,N_2927,N_2900);
and UO_35 (O_35,N_2984,N_2936);
nor UO_36 (O_36,N_2950,N_2989);
nor UO_37 (O_37,N_2994,N_2911);
nor UO_38 (O_38,N_2939,N_2956);
nand UO_39 (O_39,N_2970,N_2958);
and UO_40 (O_40,N_2935,N_2917);
nand UO_41 (O_41,N_2903,N_2954);
or UO_42 (O_42,N_2908,N_2985);
nand UO_43 (O_43,N_2928,N_2955);
xnor UO_44 (O_44,N_2961,N_2964);
nand UO_45 (O_45,N_2953,N_2941);
nor UO_46 (O_46,N_2921,N_2996);
or UO_47 (O_47,N_2931,N_2993);
and UO_48 (O_48,N_2937,N_2923);
nand UO_49 (O_49,N_2995,N_2973);
or UO_50 (O_50,N_2924,N_2955);
and UO_51 (O_51,N_2950,N_2978);
nor UO_52 (O_52,N_2949,N_2954);
and UO_53 (O_53,N_2921,N_2984);
nand UO_54 (O_54,N_2987,N_2999);
or UO_55 (O_55,N_2923,N_2922);
nand UO_56 (O_56,N_2975,N_2953);
and UO_57 (O_57,N_2988,N_2944);
or UO_58 (O_58,N_2928,N_2922);
or UO_59 (O_59,N_2961,N_2900);
or UO_60 (O_60,N_2958,N_2955);
and UO_61 (O_61,N_2967,N_2984);
and UO_62 (O_62,N_2996,N_2930);
nor UO_63 (O_63,N_2990,N_2996);
nand UO_64 (O_64,N_2970,N_2952);
and UO_65 (O_65,N_2935,N_2957);
nor UO_66 (O_66,N_2992,N_2985);
and UO_67 (O_67,N_2989,N_2990);
nor UO_68 (O_68,N_2955,N_2900);
or UO_69 (O_69,N_2933,N_2974);
and UO_70 (O_70,N_2926,N_2992);
or UO_71 (O_71,N_2984,N_2945);
or UO_72 (O_72,N_2917,N_2949);
and UO_73 (O_73,N_2943,N_2910);
nor UO_74 (O_74,N_2965,N_2976);
or UO_75 (O_75,N_2959,N_2976);
and UO_76 (O_76,N_2924,N_2962);
or UO_77 (O_77,N_2915,N_2981);
nor UO_78 (O_78,N_2978,N_2901);
or UO_79 (O_79,N_2911,N_2917);
or UO_80 (O_80,N_2952,N_2965);
or UO_81 (O_81,N_2928,N_2947);
nand UO_82 (O_82,N_2943,N_2923);
or UO_83 (O_83,N_2953,N_2936);
and UO_84 (O_84,N_2932,N_2941);
xor UO_85 (O_85,N_2964,N_2932);
or UO_86 (O_86,N_2969,N_2999);
or UO_87 (O_87,N_2983,N_2973);
nand UO_88 (O_88,N_2925,N_2950);
or UO_89 (O_89,N_2949,N_2923);
nor UO_90 (O_90,N_2925,N_2922);
nand UO_91 (O_91,N_2943,N_2914);
nand UO_92 (O_92,N_2900,N_2938);
or UO_93 (O_93,N_2974,N_2967);
nor UO_94 (O_94,N_2997,N_2910);
and UO_95 (O_95,N_2968,N_2943);
and UO_96 (O_96,N_2994,N_2964);
nor UO_97 (O_97,N_2906,N_2970);
nand UO_98 (O_98,N_2971,N_2966);
or UO_99 (O_99,N_2998,N_2957);
nor UO_100 (O_100,N_2907,N_2987);
or UO_101 (O_101,N_2940,N_2915);
and UO_102 (O_102,N_2938,N_2913);
nor UO_103 (O_103,N_2976,N_2963);
or UO_104 (O_104,N_2978,N_2966);
and UO_105 (O_105,N_2949,N_2911);
nand UO_106 (O_106,N_2958,N_2905);
nor UO_107 (O_107,N_2906,N_2930);
nand UO_108 (O_108,N_2989,N_2965);
nand UO_109 (O_109,N_2966,N_2936);
nand UO_110 (O_110,N_2933,N_2946);
nand UO_111 (O_111,N_2937,N_2918);
or UO_112 (O_112,N_2931,N_2995);
nor UO_113 (O_113,N_2903,N_2909);
or UO_114 (O_114,N_2902,N_2931);
xnor UO_115 (O_115,N_2997,N_2939);
nor UO_116 (O_116,N_2989,N_2932);
nor UO_117 (O_117,N_2926,N_2974);
nor UO_118 (O_118,N_2911,N_2950);
nor UO_119 (O_119,N_2963,N_2989);
nor UO_120 (O_120,N_2988,N_2908);
and UO_121 (O_121,N_2922,N_2912);
or UO_122 (O_122,N_2973,N_2912);
and UO_123 (O_123,N_2939,N_2964);
or UO_124 (O_124,N_2945,N_2946);
nor UO_125 (O_125,N_2949,N_2988);
nor UO_126 (O_126,N_2974,N_2916);
and UO_127 (O_127,N_2964,N_2992);
nor UO_128 (O_128,N_2991,N_2996);
or UO_129 (O_129,N_2933,N_2941);
nor UO_130 (O_130,N_2944,N_2938);
nor UO_131 (O_131,N_2920,N_2937);
or UO_132 (O_132,N_2932,N_2953);
or UO_133 (O_133,N_2908,N_2954);
nor UO_134 (O_134,N_2931,N_2969);
nor UO_135 (O_135,N_2976,N_2900);
and UO_136 (O_136,N_2920,N_2960);
nor UO_137 (O_137,N_2915,N_2943);
nor UO_138 (O_138,N_2917,N_2930);
or UO_139 (O_139,N_2911,N_2929);
or UO_140 (O_140,N_2951,N_2941);
or UO_141 (O_141,N_2930,N_2960);
nor UO_142 (O_142,N_2957,N_2977);
or UO_143 (O_143,N_2909,N_2949);
and UO_144 (O_144,N_2963,N_2966);
nand UO_145 (O_145,N_2963,N_2927);
or UO_146 (O_146,N_2904,N_2927);
and UO_147 (O_147,N_2942,N_2930);
and UO_148 (O_148,N_2923,N_2911);
nand UO_149 (O_149,N_2991,N_2990);
nor UO_150 (O_150,N_2922,N_2921);
or UO_151 (O_151,N_2988,N_2924);
and UO_152 (O_152,N_2990,N_2944);
and UO_153 (O_153,N_2950,N_2972);
nand UO_154 (O_154,N_2950,N_2981);
nand UO_155 (O_155,N_2963,N_2982);
and UO_156 (O_156,N_2944,N_2936);
xor UO_157 (O_157,N_2976,N_2948);
nand UO_158 (O_158,N_2920,N_2931);
nand UO_159 (O_159,N_2972,N_2995);
or UO_160 (O_160,N_2981,N_2975);
nor UO_161 (O_161,N_2914,N_2950);
or UO_162 (O_162,N_2985,N_2989);
nor UO_163 (O_163,N_2918,N_2964);
or UO_164 (O_164,N_2906,N_2900);
or UO_165 (O_165,N_2971,N_2925);
xor UO_166 (O_166,N_2980,N_2972);
or UO_167 (O_167,N_2927,N_2987);
nand UO_168 (O_168,N_2990,N_2950);
and UO_169 (O_169,N_2970,N_2932);
nor UO_170 (O_170,N_2908,N_2907);
or UO_171 (O_171,N_2969,N_2980);
nand UO_172 (O_172,N_2941,N_2950);
nand UO_173 (O_173,N_2973,N_2977);
nor UO_174 (O_174,N_2989,N_2961);
nand UO_175 (O_175,N_2901,N_2936);
and UO_176 (O_176,N_2971,N_2987);
or UO_177 (O_177,N_2909,N_2942);
or UO_178 (O_178,N_2914,N_2989);
or UO_179 (O_179,N_2949,N_2958);
nor UO_180 (O_180,N_2934,N_2948);
and UO_181 (O_181,N_2962,N_2915);
nor UO_182 (O_182,N_2953,N_2994);
and UO_183 (O_183,N_2996,N_2959);
and UO_184 (O_184,N_2917,N_2987);
nand UO_185 (O_185,N_2934,N_2913);
and UO_186 (O_186,N_2970,N_2967);
nand UO_187 (O_187,N_2974,N_2943);
or UO_188 (O_188,N_2949,N_2978);
or UO_189 (O_189,N_2925,N_2912);
nand UO_190 (O_190,N_2960,N_2952);
and UO_191 (O_191,N_2950,N_2940);
nor UO_192 (O_192,N_2932,N_2985);
or UO_193 (O_193,N_2956,N_2987);
nand UO_194 (O_194,N_2959,N_2998);
nor UO_195 (O_195,N_2905,N_2937);
or UO_196 (O_196,N_2954,N_2904);
nor UO_197 (O_197,N_2920,N_2973);
and UO_198 (O_198,N_2975,N_2977);
or UO_199 (O_199,N_2900,N_2936);
or UO_200 (O_200,N_2945,N_2932);
nand UO_201 (O_201,N_2961,N_2979);
and UO_202 (O_202,N_2952,N_2972);
xor UO_203 (O_203,N_2999,N_2980);
nor UO_204 (O_204,N_2991,N_2901);
or UO_205 (O_205,N_2982,N_2933);
nor UO_206 (O_206,N_2922,N_2980);
nor UO_207 (O_207,N_2903,N_2994);
and UO_208 (O_208,N_2921,N_2999);
nand UO_209 (O_209,N_2962,N_2912);
or UO_210 (O_210,N_2970,N_2904);
and UO_211 (O_211,N_2931,N_2945);
and UO_212 (O_212,N_2962,N_2916);
and UO_213 (O_213,N_2915,N_2988);
nand UO_214 (O_214,N_2942,N_2970);
or UO_215 (O_215,N_2998,N_2955);
nor UO_216 (O_216,N_2900,N_2963);
or UO_217 (O_217,N_2977,N_2971);
and UO_218 (O_218,N_2921,N_2934);
nand UO_219 (O_219,N_2936,N_2970);
and UO_220 (O_220,N_2907,N_2949);
nand UO_221 (O_221,N_2915,N_2975);
and UO_222 (O_222,N_2963,N_2977);
and UO_223 (O_223,N_2917,N_2924);
or UO_224 (O_224,N_2954,N_2944);
nand UO_225 (O_225,N_2918,N_2984);
nor UO_226 (O_226,N_2965,N_2945);
nand UO_227 (O_227,N_2957,N_2991);
nand UO_228 (O_228,N_2961,N_2938);
nor UO_229 (O_229,N_2998,N_2973);
nor UO_230 (O_230,N_2960,N_2957);
or UO_231 (O_231,N_2964,N_2973);
nand UO_232 (O_232,N_2963,N_2912);
or UO_233 (O_233,N_2952,N_2958);
nor UO_234 (O_234,N_2926,N_2930);
nor UO_235 (O_235,N_2959,N_2983);
nor UO_236 (O_236,N_2907,N_2942);
nor UO_237 (O_237,N_2961,N_2905);
nor UO_238 (O_238,N_2919,N_2944);
and UO_239 (O_239,N_2959,N_2974);
and UO_240 (O_240,N_2918,N_2963);
or UO_241 (O_241,N_2951,N_2927);
nand UO_242 (O_242,N_2905,N_2936);
or UO_243 (O_243,N_2992,N_2910);
and UO_244 (O_244,N_2917,N_2992);
and UO_245 (O_245,N_2901,N_2951);
or UO_246 (O_246,N_2928,N_2913);
and UO_247 (O_247,N_2902,N_2954);
nand UO_248 (O_248,N_2933,N_2940);
and UO_249 (O_249,N_2973,N_2941);
or UO_250 (O_250,N_2998,N_2938);
and UO_251 (O_251,N_2911,N_2942);
nand UO_252 (O_252,N_2904,N_2972);
or UO_253 (O_253,N_2963,N_2931);
or UO_254 (O_254,N_2960,N_2953);
nor UO_255 (O_255,N_2971,N_2937);
or UO_256 (O_256,N_2965,N_2917);
or UO_257 (O_257,N_2909,N_2984);
and UO_258 (O_258,N_2957,N_2941);
or UO_259 (O_259,N_2992,N_2903);
nor UO_260 (O_260,N_2913,N_2930);
and UO_261 (O_261,N_2969,N_2910);
nor UO_262 (O_262,N_2918,N_2954);
and UO_263 (O_263,N_2946,N_2952);
or UO_264 (O_264,N_2963,N_2941);
or UO_265 (O_265,N_2908,N_2987);
or UO_266 (O_266,N_2954,N_2979);
or UO_267 (O_267,N_2959,N_2975);
nor UO_268 (O_268,N_2950,N_2962);
nand UO_269 (O_269,N_2984,N_2953);
or UO_270 (O_270,N_2916,N_2973);
nor UO_271 (O_271,N_2947,N_2956);
nor UO_272 (O_272,N_2994,N_2950);
or UO_273 (O_273,N_2934,N_2906);
nor UO_274 (O_274,N_2963,N_2958);
and UO_275 (O_275,N_2908,N_2946);
nand UO_276 (O_276,N_2941,N_2904);
nor UO_277 (O_277,N_2907,N_2902);
or UO_278 (O_278,N_2994,N_2937);
and UO_279 (O_279,N_2996,N_2910);
nor UO_280 (O_280,N_2934,N_2966);
and UO_281 (O_281,N_2975,N_2997);
nand UO_282 (O_282,N_2908,N_2969);
and UO_283 (O_283,N_2925,N_2953);
nor UO_284 (O_284,N_2951,N_2975);
or UO_285 (O_285,N_2926,N_2931);
nor UO_286 (O_286,N_2981,N_2911);
or UO_287 (O_287,N_2903,N_2930);
nand UO_288 (O_288,N_2949,N_2914);
nor UO_289 (O_289,N_2974,N_2961);
or UO_290 (O_290,N_2987,N_2995);
nand UO_291 (O_291,N_2920,N_2972);
nand UO_292 (O_292,N_2927,N_2913);
nand UO_293 (O_293,N_2943,N_2978);
nand UO_294 (O_294,N_2922,N_2903);
or UO_295 (O_295,N_2938,N_2925);
or UO_296 (O_296,N_2919,N_2952);
nand UO_297 (O_297,N_2922,N_2977);
and UO_298 (O_298,N_2926,N_2985);
and UO_299 (O_299,N_2958,N_2937);
nand UO_300 (O_300,N_2938,N_2967);
nand UO_301 (O_301,N_2934,N_2943);
or UO_302 (O_302,N_2983,N_2991);
or UO_303 (O_303,N_2919,N_2945);
and UO_304 (O_304,N_2971,N_2910);
or UO_305 (O_305,N_2989,N_2948);
nor UO_306 (O_306,N_2978,N_2906);
and UO_307 (O_307,N_2987,N_2960);
and UO_308 (O_308,N_2979,N_2919);
nand UO_309 (O_309,N_2998,N_2920);
or UO_310 (O_310,N_2908,N_2900);
nand UO_311 (O_311,N_2907,N_2926);
and UO_312 (O_312,N_2938,N_2989);
and UO_313 (O_313,N_2924,N_2977);
or UO_314 (O_314,N_2992,N_2934);
nand UO_315 (O_315,N_2900,N_2923);
or UO_316 (O_316,N_2979,N_2999);
nor UO_317 (O_317,N_2929,N_2970);
nor UO_318 (O_318,N_2940,N_2958);
nand UO_319 (O_319,N_2969,N_2944);
or UO_320 (O_320,N_2994,N_2902);
nor UO_321 (O_321,N_2929,N_2983);
nand UO_322 (O_322,N_2966,N_2956);
and UO_323 (O_323,N_2942,N_2985);
and UO_324 (O_324,N_2997,N_2973);
nor UO_325 (O_325,N_2981,N_2997);
and UO_326 (O_326,N_2926,N_2988);
and UO_327 (O_327,N_2963,N_2979);
nor UO_328 (O_328,N_2952,N_2982);
nor UO_329 (O_329,N_2907,N_2978);
nor UO_330 (O_330,N_2980,N_2931);
or UO_331 (O_331,N_2905,N_2944);
nor UO_332 (O_332,N_2939,N_2982);
nor UO_333 (O_333,N_2916,N_2915);
and UO_334 (O_334,N_2981,N_2932);
and UO_335 (O_335,N_2902,N_2936);
and UO_336 (O_336,N_2926,N_2910);
or UO_337 (O_337,N_2981,N_2992);
nor UO_338 (O_338,N_2979,N_2932);
nand UO_339 (O_339,N_2965,N_2972);
and UO_340 (O_340,N_2969,N_2972);
nor UO_341 (O_341,N_2988,N_2920);
and UO_342 (O_342,N_2961,N_2949);
nor UO_343 (O_343,N_2993,N_2903);
nand UO_344 (O_344,N_2920,N_2951);
and UO_345 (O_345,N_2960,N_2974);
nand UO_346 (O_346,N_2938,N_2911);
nor UO_347 (O_347,N_2903,N_2975);
and UO_348 (O_348,N_2903,N_2913);
nand UO_349 (O_349,N_2920,N_2995);
nor UO_350 (O_350,N_2910,N_2950);
or UO_351 (O_351,N_2980,N_2930);
and UO_352 (O_352,N_2987,N_2962);
or UO_353 (O_353,N_2992,N_2958);
and UO_354 (O_354,N_2921,N_2977);
and UO_355 (O_355,N_2973,N_2936);
or UO_356 (O_356,N_2914,N_2986);
nor UO_357 (O_357,N_2934,N_2980);
nor UO_358 (O_358,N_2968,N_2989);
nor UO_359 (O_359,N_2961,N_2998);
nor UO_360 (O_360,N_2993,N_2915);
or UO_361 (O_361,N_2956,N_2969);
or UO_362 (O_362,N_2999,N_2970);
and UO_363 (O_363,N_2950,N_2974);
nor UO_364 (O_364,N_2951,N_2949);
and UO_365 (O_365,N_2965,N_2901);
nor UO_366 (O_366,N_2972,N_2941);
nand UO_367 (O_367,N_2904,N_2986);
nand UO_368 (O_368,N_2934,N_2972);
or UO_369 (O_369,N_2939,N_2955);
and UO_370 (O_370,N_2919,N_2911);
nor UO_371 (O_371,N_2981,N_2948);
nand UO_372 (O_372,N_2946,N_2996);
nand UO_373 (O_373,N_2958,N_2956);
or UO_374 (O_374,N_2999,N_2988);
nand UO_375 (O_375,N_2942,N_2950);
and UO_376 (O_376,N_2958,N_2944);
nand UO_377 (O_377,N_2983,N_2995);
or UO_378 (O_378,N_2900,N_2974);
nor UO_379 (O_379,N_2966,N_2980);
nand UO_380 (O_380,N_2955,N_2959);
nand UO_381 (O_381,N_2974,N_2909);
or UO_382 (O_382,N_2962,N_2971);
or UO_383 (O_383,N_2903,N_2978);
nor UO_384 (O_384,N_2900,N_2954);
nand UO_385 (O_385,N_2970,N_2901);
nor UO_386 (O_386,N_2940,N_2966);
or UO_387 (O_387,N_2950,N_2957);
nor UO_388 (O_388,N_2951,N_2917);
or UO_389 (O_389,N_2973,N_2930);
xnor UO_390 (O_390,N_2917,N_2962);
and UO_391 (O_391,N_2909,N_2960);
nand UO_392 (O_392,N_2931,N_2978);
and UO_393 (O_393,N_2913,N_2950);
or UO_394 (O_394,N_2973,N_2940);
and UO_395 (O_395,N_2942,N_2908);
or UO_396 (O_396,N_2942,N_2989);
nand UO_397 (O_397,N_2975,N_2904);
or UO_398 (O_398,N_2994,N_2958);
nor UO_399 (O_399,N_2903,N_2928);
nand UO_400 (O_400,N_2939,N_2932);
or UO_401 (O_401,N_2954,N_2957);
nand UO_402 (O_402,N_2906,N_2953);
and UO_403 (O_403,N_2900,N_2995);
nor UO_404 (O_404,N_2947,N_2926);
nand UO_405 (O_405,N_2993,N_2990);
and UO_406 (O_406,N_2952,N_2975);
nand UO_407 (O_407,N_2999,N_2911);
and UO_408 (O_408,N_2989,N_2905);
or UO_409 (O_409,N_2970,N_2984);
xnor UO_410 (O_410,N_2915,N_2938);
nand UO_411 (O_411,N_2952,N_2904);
nand UO_412 (O_412,N_2994,N_2959);
or UO_413 (O_413,N_2939,N_2933);
or UO_414 (O_414,N_2908,N_2922);
and UO_415 (O_415,N_2975,N_2933);
and UO_416 (O_416,N_2995,N_2971);
or UO_417 (O_417,N_2986,N_2985);
nand UO_418 (O_418,N_2913,N_2988);
and UO_419 (O_419,N_2971,N_2921);
nor UO_420 (O_420,N_2950,N_2904);
or UO_421 (O_421,N_2981,N_2965);
nor UO_422 (O_422,N_2931,N_2988);
and UO_423 (O_423,N_2980,N_2918);
nand UO_424 (O_424,N_2923,N_2903);
nor UO_425 (O_425,N_2924,N_2981);
nand UO_426 (O_426,N_2922,N_2969);
nor UO_427 (O_427,N_2992,N_2951);
and UO_428 (O_428,N_2931,N_2939);
nand UO_429 (O_429,N_2968,N_2925);
or UO_430 (O_430,N_2939,N_2994);
and UO_431 (O_431,N_2927,N_2977);
nor UO_432 (O_432,N_2996,N_2992);
or UO_433 (O_433,N_2957,N_2915);
nor UO_434 (O_434,N_2918,N_2950);
or UO_435 (O_435,N_2982,N_2951);
or UO_436 (O_436,N_2925,N_2966);
and UO_437 (O_437,N_2988,N_2921);
or UO_438 (O_438,N_2996,N_2968);
and UO_439 (O_439,N_2984,N_2991);
nand UO_440 (O_440,N_2967,N_2986);
nand UO_441 (O_441,N_2967,N_2915);
nand UO_442 (O_442,N_2993,N_2943);
or UO_443 (O_443,N_2922,N_2937);
nand UO_444 (O_444,N_2975,N_2954);
nor UO_445 (O_445,N_2983,N_2984);
nand UO_446 (O_446,N_2907,N_2922);
nand UO_447 (O_447,N_2954,N_2988);
and UO_448 (O_448,N_2931,N_2944);
nand UO_449 (O_449,N_2924,N_2938);
and UO_450 (O_450,N_2901,N_2907);
or UO_451 (O_451,N_2995,N_2941);
nor UO_452 (O_452,N_2973,N_2919);
or UO_453 (O_453,N_2977,N_2918);
and UO_454 (O_454,N_2947,N_2974);
nor UO_455 (O_455,N_2981,N_2961);
nor UO_456 (O_456,N_2964,N_2976);
nand UO_457 (O_457,N_2900,N_2911);
nand UO_458 (O_458,N_2916,N_2996);
nand UO_459 (O_459,N_2950,N_2999);
nor UO_460 (O_460,N_2915,N_2931);
or UO_461 (O_461,N_2928,N_2988);
xnor UO_462 (O_462,N_2970,N_2972);
nor UO_463 (O_463,N_2949,N_2934);
and UO_464 (O_464,N_2965,N_2957);
or UO_465 (O_465,N_2979,N_2966);
and UO_466 (O_466,N_2970,N_2996);
nor UO_467 (O_467,N_2919,N_2903);
and UO_468 (O_468,N_2900,N_2967);
and UO_469 (O_469,N_2900,N_2943);
nor UO_470 (O_470,N_2995,N_2905);
and UO_471 (O_471,N_2970,N_2931);
nand UO_472 (O_472,N_2917,N_2953);
nand UO_473 (O_473,N_2976,N_2907);
nand UO_474 (O_474,N_2989,N_2971);
or UO_475 (O_475,N_2963,N_2945);
and UO_476 (O_476,N_2903,N_2949);
or UO_477 (O_477,N_2944,N_2963);
nor UO_478 (O_478,N_2902,N_2975);
or UO_479 (O_479,N_2955,N_2946);
nor UO_480 (O_480,N_2907,N_2900);
and UO_481 (O_481,N_2908,N_2972);
nand UO_482 (O_482,N_2906,N_2946);
nand UO_483 (O_483,N_2984,N_2933);
nand UO_484 (O_484,N_2994,N_2912);
nor UO_485 (O_485,N_2987,N_2914);
nor UO_486 (O_486,N_2981,N_2958);
nand UO_487 (O_487,N_2952,N_2997);
nand UO_488 (O_488,N_2920,N_2986);
and UO_489 (O_489,N_2907,N_2939);
nor UO_490 (O_490,N_2921,N_2938);
and UO_491 (O_491,N_2982,N_2919);
nand UO_492 (O_492,N_2961,N_2944);
xnor UO_493 (O_493,N_2909,N_2956);
or UO_494 (O_494,N_2959,N_2946);
nand UO_495 (O_495,N_2968,N_2902);
nand UO_496 (O_496,N_2989,N_2935);
and UO_497 (O_497,N_2961,N_2953);
nand UO_498 (O_498,N_2949,N_2962);
or UO_499 (O_499,N_2996,N_2994);
endmodule