module basic_1000_10000_1500_5_levels_2xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nand U0 (N_0,In_947,In_840);
and U1 (N_1,In_208,In_170);
nand U2 (N_2,In_710,In_106);
nor U3 (N_3,In_19,In_724);
and U4 (N_4,In_108,In_163);
or U5 (N_5,In_490,In_30);
nand U6 (N_6,In_593,In_68);
nor U7 (N_7,In_914,In_948);
nand U8 (N_8,In_830,In_267);
nor U9 (N_9,In_354,In_725);
or U10 (N_10,In_944,In_447);
nor U11 (N_11,In_920,In_425);
and U12 (N_12,In_618,In_649);
nor U13 (N_13,In_276,In_270);
or U14 (N_14,In_980,In_321);
or U15 (N_15,In_959,In_856);
and U16 (N_16,In_364,In_320);
or U17 (N_17,In_694,In_774);
and U18 (N_18,In_778,In_214);
nor U19 (N_19,In_40,In_84);
or U20 (N_20,In_49,In_719);
or U21 (N_21,In_446,In_736);
and U22 (N_22,In_288,In_240);
or U23 (N_23,In_32,In_620);
or U24 (N_24,In_556,In_723);
nand U25 (N_25,In_135,In_137);
nor U26 (N_26,In_881,In_924);
or U27 (N_27,In_118,In_528);
nand U28 (N_28,In_103,In_659);
or U29 (N_29,In_931,In_297);
or U30 (N_30,In_493,In_484);
nand U31 (N_31,In_245,In_526);
and U32 (N_32,In_677,In_460);
xor U33 (N_33,In_353,In_48);
nor U34 (N_34,In_94,In_396);
nand U35 (N_35,In_901,In_956);
nand U36 (N_36,In_949,In_718);
nand U37 (N_37,In_278,In_394);
nand U38 (N_38,In_735,In_603);
or U39 (N_39,In_745,In_442);
nor U40 (N_40,In_189,In_992);
and U41 (N_41,In_524,In_699);
nand U42 (N_42,In_144,In_669);
nor U43 (N_43,In_344,In_995);
nor U44 (N_44,In_294,In_802);
nor U45 (N_45,In_177,In_104);
xnor U46 (N_46,In_762,In_158);
or U47 (N_47,In_525,In_702);
nand U48 (N_48,In_129,In_458);
nor U49 (N_49,In_617,In_8);
nor U50 (N_50,In_266,In_18);
nor U51 (N_51,In_293,In_4);
and U52 (N_52,In_349,In_113);
xor U53 (N_53,In_749,In_209);
nor U54 (N_54,In_188,In_565);
and U55 (N_55,In_65,In_913);
nor U56 (N_56,In_87,In_591);
and U57 (N_57,In_898,In_822);
nand U58 (N_58,In_433,In_835);
nor U59 (N_59,In_503,In_336);
or U60 (N_60,In_777,In_863);
nand U61 (N_61,In_417,In_77);
nand U62 (N_62,In_849,In_95);
or U63 (N_63,In_839,In_81);
and U64 (N_64,In_27,In_615);
or U65 (N_65,In_207,In_585);
nor U66 (N_66,In_916,In_476);
nand U67 (N_67,In_482,In_776);
nor U68 (N_68,In_641,In_707);
and U69 (N_69,In_690,In_346);
nand U70 (N_70,In_993,In_559);
nand U71 (N_71,In_979,In_411);
and U72 (N_72,In_632,In_226);
nand U73 (N_73,In_60,In_653);
nand U74 (N_74,In_703,In_444);
nand U75 (N_75,In_800,In_287);
and U76 (N_76,In_536,In_594);
or U77 (N_77,In_773,In_866);
nand U78 (N_78,In_637,In_187);
or U79 (N_79,In_974,In_408);
or U80 (N_80,In_58,In_90);
or U81 (N_81,In_644,In_789);
and U82 (N_82,In_483,In_631);
or U83 (N_83,In_879,In_414);
nor U84 (N_84,In_784,In_100);
or U85 (N_85,In_125,In_627);
and U86 (N_86,In_398,In_613);
nor U87 (N_87,In_96,In_260);
nand U88 (N_88,In_728,In_117);
nand U89 (N_89,In_497,In_661);
or U90 (N_90,In_315,In_343);
nor U91 (N_91,In_56,In_792);
or U92 (N_92,In_431,In_574);
xor U93 (N_93,In_853,In_421);
and U94 (N_94,In_922,In_133);
nand U95 (N_95,In_679,In_160);
nand U96 (N_96,In_57,In_811);
nor U97 (N_97,In_737,In_656);
or U98 (N_98,In_572,In_558);
and U99 (N_99,In_561,In_392);
and U100 (N_100,In_934,In_584);
and U101 (N_101,In_608,In_872);
or U102 (N_102,In_846,In_801);
nor U103 (N_103,In_227,In_376);
nand U104 (N_104,In_804,In_410);
and U105 (N_105,In_206,In_341);
or U106 (N_106,In_616,In_467);
or U107 (N_107,In_324,In_305);
nor U108 (N_108,In_642,In_262);
nor U109 (N_109,In_850,In_127);
xor U110 (N_110,In_420,In_571);
xnor U111 (N_111,In_440,In_242);
or U112 (N_112,In_501,In_966);
nand U113 (N_113,In_579,In_468);
or U114 (N_114,In_666,In_734);
nand U115 (N_115,In_475,In_53);
and U116 (N_116,In_510,In_906);
nor U117 (N_117,In_314,In_93);
nor U118 (N_118,In_530,In_887);
xor U119 (N_119,In_542,In_697);
nand U120 (N_120,In_456,In_121);
nor U121 (N_121,In_80,In_692);
or U122 (N_122,In_828,In_652);
nor U123 (N_123,In_428,In_643);
or U124 (N_124,In_843,In_798);
or U125 (N_125,In_63,In_325);
nor U126 (N_126,In_858,In_409);
and U127 (N_127,In_857,In_547);
xnor U128 (N_128,In_646,In_676);
xor U129 (N_129,In_997,In_854);
nor U130 (N_130,In_888,In_356);
nor U131 (N_131,In_79,In_740);
nand U132 (N_132,In_836,In_996);
or U133 (N_133,In_391,In_464);
nand U134 (N_134,In_670,In_377);
and U135 (N_135,In_123,In_481);
and U136 (N_136,In_965,In_167);
nor U137 (N_137,In_303,In_371);
nor U138 (N_138,In_46,In_359);
and U139 (N_139,In_280,In_301);
nand U140 (N_140,In_806,In_969);
nand U141 (N_141,In_671,In_805);
nor U142 (N_142,In_415,In_779);
nor U143 (N_143,In_50,In_673);
and U144 (N_144,In_861,In_252);
nor U145 (N_145,In_900,In_488);
nor U146 (N_146,In_648,In_213);
nand U147 (N_147,In_557,In_578);
nor U148 (N_148,In_115,In_833);
and U149 (N_149,In_386,In_384);
or U150 (N_150,In_363,In_210);
nand U151 (N_151,In_935,In_165);
nor U152 (N_152,In_701,In_59);
or U153 (N_153,In_533,In_687);
nor U154 (N_154,In_471,In_139);
nand U155 (N_155,In_326,In_516);
nand U156 (N_156,In_991,In_246);
nand U157 (N_157,In_549,In_662);
nor U158 (N_158,In_712,In_66);
nor U159 (N_159,In_829,In_522);
and U160 (N_160,In_874,In_793);
xnor U161 (N_161,In_852,In_588);
nor U162 (N_162,In_215,In_132);
or U163 (N_163,In_519,In_17);
nor U164 (N_164,In_926,In_757);
or U165 (N_165,In_834,In_799);
nor U166 (N_166,In_824,In_611);
and U167 (N_167,In_672,In_248);
nand U168 (N_168,In_332,In_682);
nand U169 (N_169,In_105,In_954);
and U170 (N_170,In_292,In_282);
or U171 (N_171,In_201,In_284);
and U172 (N_172,In_31,In_604);
nor U173 (N_173,In_927,In_638);
or U174 (N_174,In_112,In_154);
and U175 (N_175,In_795,In_668);
or U176 (N_176,In_131,In_576);
nand U177 (N_177,In_52,In_496);
and U178 (N_178,In_936,In_469);
nand U179 (N_179,In_984,In_485);
nand U180 (N_180,In_10,In_610);
nand U181 (N_181,In_511,In_192);
nand U182 (N_182,In_752,In_381);
or U183 (N_183,In_827,In_686);
nor U184 (N_184,In_271,In_904);
nor U185 (N_185,In_491,In_554);
nand U186 (N_186,In_832,In_564);
nand U187 (N_187,In_352,In_894);
nor U188 (N_188,In_395,In_76);
or U189 (N_189,In_38,In_300);
or U190 (N_190,In_423,In_318);
nand U191 (N_191,In_771,In_575);
nor U192 (N_192,In_21,In_590);
or U193 (N_193,In_514,In_29);
xnor U194 (N_194,In_272,In_943);
and U195 (N_195,In_28,In_24);
and U196 (N_196,In_950,In_205);
nor U197 (N_197,In_930,In_438);
and U198 (N_198,In_917,In_595);
and U199 (N_199,In_876,In_534);
nand U200 (N_200,In_678,In_42);
or U201 (N_201,In_727,In_309);
and U202 (N_202,In_153,In_259);
nand U203 (N_203,In_709,In_597);
nor U204 (N_204,In_26,In_358);
nor U205 (N_205,In_383,In_439);
nor U206 (N_206,In_929,In_85);
nand U207 (N_207,In_472,In_498);
and U208 (N_208,In_255,In_71);
and U209 (N_209,In_838,In_961);
xnor U210 (N_210,In_987,In_3);
and U211 (N_211,In_212,In_580);
nand U212 (N_212,In_751,In_808);
nand U213 (N_213,In_122,In_903);
nand U214 (N_214,In_243,In_290);
nor U215 (N_215,In_454,In_495);
nand U216 (N_216,In_819,In_814);
nor U217 (N_217,In_116,In_543);
or U218 (N_218,In_817,In_770);
or U219 (N_219,In_860,In_161);
and U220 (N_220,In_695,In_126);
nor U221 (N_221,In_286,In_750);
nand U222 (N_222,In_261,In_787);
nor U223 (N_223,In_655,In_462);
or U224 (N_224,In_810,In_147);
nand U225 (N_225,In_385,In_298);
nor U226 (N_226,In_387,In_855);
nand U227 (N_227,In_990,In_92);
nor U228 (N_228,In_680,In_761);
and U229 (N_229,In_64,In_775);
or U230 (N_230,In_660,In_635);
nand U231 (N_231,In_291,In_923);
nor U232 (N_232,In_971,In_279);
nand U233 (N_233,In_114,In_361);
or U234 (N_234,In_848,In_527);
nor U235 (N_235,In_622,In_625);
and U236 (N_236,In_782,In_548);
nand U237 (N_237,In_143,In_487);
and U238 (N_238,In_202,In_864);
and U239 (N_239,In_263,In_818);
xnor U240 (N_240,In_859,In_746);
and U241 (N_241,In_577,In_871);
and U242 (N_242,In_128,In_470);
xor U243 (N_243,In_599,In_658);
nand U244 (N_244,In_945,In_541);
nand U245 (N_245,In_902,In_12);
nand U246 (N_246,In_319,In_765);
nor U247 (N_247,In_870,In_601);
or U248 (N_248,In_329,In_582);
nor U249 (N_249,In_311,In_551);
or U250 (N_250,In_140,In_5);
and U251 (N_251,In_960,In_639);
or U252 (N_252,In_862,In_696);
and U253 (N_253,In_907,In_111);
or U254 (N_254,In_119,In_407);
nor U255 (N_255,In_698,In_463);
or U256 (N_256,In_508,In_480);
and U257 (N_257,In_918,In_754);
nor U258 (N_258,In_758,In_239);
and U259 (N_259,In_891,In_217);
xnor U260 (N_260,In_986,In_928);
nor U261 (N_261,In_756,In_589);
or U262 (N_262,In_193,In_342);
xnor U263 (N_263,In_11,In_507);
and U264 (N_264,In_505,In_178);
nor U265 (N_265,In_457,In_640);
and U266 (N_266,In_550,In_667);
nor U267 (N_267,In_184,In_517);
nand U268 (N_268,In_389,In_970);
xnor U269 (N_269,In_772,In_844);
nor U270 (N_270,In_544,In_932);
nand U271 (N_271,In_403,In_847);
xnor U272 (N_272,In_759,In_665);
or U273 (N_273,In_841,In_99);
nand U274 (N_274,In_919,In_78);
nand U275 (N_275,In_72,In_809);
nand U276 (N_276,In_452,In_748);
nand U277 (N_277,In_355,In_351);
and U278 (N_278,In_22,In_739);
and U279 (N_279,In_450,In_166);
nor U280 (N_280,In_722,In_717);
nand U281 (N_281,In_138,In_573);
nand U282 (N_282,In_247,In_397);
nand U283 (N_283,In_837,In_897);
nand U284 (N_284,In_747,In_957);
and U285 (N_285,In_174,In_313);
or U286 (N_286,In_231,In_474);
and U287 (N_287,In_674,In_241);
nor U288 (N_288,In_769,In_538);
nand U289 (N_289,In_162,In_333);
and U290 (N_290,In_883,In_275);
nand U291 (N_291,In_952,In_268);
nor U292 (N_292,In_235,In_317);
nor U293 (N_293,In_994,In_13);
xnor U294 (N_294,In_513,In_0);
and U295 (N_295,In_607,In_865);
or U296 (N_296,In_647,In_726);
nand U297 (N_297,In_264,In_869);
or U298 (N_298,In_316,In_441);
or U299 (N_299,In_940,In_337);
or U300 (N_300,In_197,In_486);
or U301 (N_301,In_448,In_426);
or U302 (N_302,In_732,In_289);
or U303 (N_303,In_975,In_370);
xnor U304 (N_304,In_195,In_626);
or U305 (N_305,In_569,In_962);
or U306 (N_306,In_186,In_895);
or U307 (N_307,In_729,In_281);
or U308 (N_308,In_339,In_714);
or U309 (N_309,In_552,In_393);
and U310 (N_310,In_148,In_515);
nor U311 (N_311,In_37,In_418);
or U312 (N_312,In_741,In_560);
and U313 (N_313,In_390,In_156);
nor U314 (N_314,In_61,In_296);
nor U315 (N_315,In_405,In_803);
nor U316 (N_316,In_546,In_708);
or U317 (N_317,In_509,In_786);
nand U318 (N_318,In_624,In_198);
nand U319 (N_319,In_763,In_159);
or U320 (N_320,In_283,In_964);
and U321 (N_321,In_98,In_823);
nand U322 (N_322,In_365,In_941);
and U323 (N_323,In_629,In_842);
or U324 (N_324,In_338,In_285);
and U325 (N_325,In_743,In_731);
nand U326 (N_326,In_937,In_882);
nor U327 (N_327,In_766,In_15);
and U328 (N_328,In_130,In_650);
nand U329 (N_329,In_738,In_312);
xnor U330 (N_330,In_764,In_684);
nand U331 (N_331,In_911,In_374);
or U332 (N_332,In_436,In_89);
and U333 (N_333,In_753,In_372);
nand U334 (N_334,In_477,In_688);
nand U335 (N_335,In_568,In_185);
or U336 (N_336,In_54,In_523);
nor U337 (N_337,In_499,In_258);
nand U338 (N_338,In_150,In_586);
or U339 (N_339,In_369,In_890);
nand U340 (N_340,In_357,In_437);
and U341 (N_341,In_401,In_142);
nand U342 (N_342,In_400,In_691);
and U343 (N_343,In_47,In_304);
nand U344 (N_344,In_831,In_225);
or U345 (N_345,In_815,In_999);
or U346 (N_346,In_151,In_788);
or U347 (N_347,In_373,In_783);
and U348 (N_348,In_102,In_120);
and U349 (N_349,In_36,In_466);
nand U350 (N_350,In_2,In_628);
or U351 (N_351,In_73,In_478);
nand U352 (N_352,In_380,In_97);
and U353 (N_353,In_350,In_567);
and U354 (N_354,In_716,In_274);
nor U355 (N_355,In_465,In_877);
or U356 (N_356,In_33,In_257);
nor U357 (N_357,In_681,In_172);
nor U358 (N_358,In_715,In_479);
or U359 (N_359,In_981,In_175);
and U360 (N_360,In_500,In_330);
and U361 (N_361,In_875,In_938);
nand U362 (N_362,In_711,In_196);
or U363 (N_363,In_553,In_755);
and U364 (N_364,In_55,In_449);
nand U365 (N_365,In_190,In_596);
nor U366 (N_366,In_14,In_880);
or U367 (N_367,In_972,In_933);
or U368 (N_368,In_953,In_88);
or U369 (N_369,In_563,In_367);
nor U370 (N_370,In_328,In_265);
nand U371 (N_371,In_512,In_989);
nand U372 (N_372,In_909,In_583);
nand U373 (N_373,In_908,In_39);
or U374 (N_374,In_6,In_230);
nand U375 (N_375,In_306,In_253);
nand U376 (N_376,In_155,In_223);
nor U377 (N_377,In_958,In_461);
and U378 (N_378,In_70,In_51);
nand U379 (N_379,In_375,In_221);
and U380 (N_380,In_413,In_234);
nand U381 (N_381,In_445,In_110);
and U382 (N_382,In_16,In_915);
xor U383 (N_383,In_796,In_200);
and U384 (N_384,In_562,In_685);
nand U385 (N_385,In_899,In_45);
nand U386 (N_386,In_169,In_539);
and U387 (N_387,In_893,In_606);
and U388 (N_388,In_249,In_299);
nand U389 (N_389,In_494,In_360);
or U390 (N_390,In_744,In_345);
and U391 (N_391,In_402,In_220);
nand U392 (N_392,In_566,In_705);
and U393 (N_393,In_785,In_335);
and U394 (N_394,In_302,In_182);
nor U395 (N_395,In_905,In_236);
and U396 (N_396,In_250,In_75);
nand U397 (N_397,In_435,In_967);
and U398 (N_398,In_978,In_636);
and U399 (N_399,In_910,In_422);
nand U400 (N_400,In_233,In_107);
xnor U401 (N_401,In_645,In_224);
xnor U402 (N_402,In_362,In_327);
or U403 (N_403,In_794,In_378);
and U404 (N_404,In_134,In_430);
nand U405 (N_405,In_531,In_868);
and U406 (N_406,In_609,In_307);
and U407 (N_407,In_521,In_20);
or U408 (N_408,In_191,In_168);
and U409 (N_409,In_219,In_985);
nand U410 (N_410,In_942,In_540);
nor U411 (N_411,In_295,In_145);
nor U412 (N_412,In_878,In_973);
nand U413 (N_413,In_149,In_529);
nor U414 (N_414,In_323,In_797);
or U415 (N_415,In_340,In_700);
and U416 (N_416,In_41,In_675);
nand U417 (N_417,In_216,In_25);
or U418 (N_418,In_532,In_251);
nand U419 (N_419,In_713,In_331);
and U420 (N_420,In_555,In_74);
nor U421 (N_421,In_605,In_152);
and U422 (N_422,In_388,In_489);
nor U423 (N_423,In_845,In_1);
or U424 (N_424,In_504,In_101);
and U425 (N_425,In_612,In_619);
nand U426 (N_426,In_683,In_614);
and U427 (N_427,In_767,In_976);
nand U428 (N_428,In_379,In_238);
nand U429 (N_429,In_651,In_171);
and U430 (N_430,In_816,In_419);
nand U431 (N_431,In_760,In_781);
nand U432 (N_432,In_780,In_334);
nor U433 (N_433,In_183,In_109);
nand U434 (N_434,In_199,In_518);
or U435 (N_435,In_998,In_141);
nor U436 (N_436,In_406,In_256);
or U437 (N_437,In_194,In_742);
or U438 (N_438,In_768,In_244);
nor U439 (N_439,In_623,In_813);
or U440 (N_440,In_912,In_9);
and U441 (N_441,In_693,In_269);
nand U442 (N_442,In_136,In_412);
nand U443 (N_443,In_124,In_654);
nand U444 (N_444,In_404,In_164);
and U445 (N_445,In_432,In_825);
and U446 (N_446,In_229,In_416);
or U447 (N_447,In_939,In_277);
nor U448 (N_448,In_157,In_67);
or U449 (N_449,In_443,In_308);
and U450 (N_450,In_322,In_873);
nand U451 (N_451,In_537,In_473);
nand U452 (N_452,In_982,In_570);
and U453 (N_453,In_535,In_146);
or U454 (N_454,In_427,In_598);
or U455 (N_455,In_892,In_884);
or U456 (N_456,In_176,In_520);
nor U457 (N_457,In_502,In_983);
nor U458 (N_458,In_211,In_602);
or U459 (N_459,In_232,In_721);
and U460 (N_460,In_946,In_704);
nand U461 (N_461,In_977,In_925);
and U462 (N_462,In_506,In_807);
nand U463 (N_463,In_399,In_273);
or U464 (N_464,In_968,In_228);
xor U465 (N_465,In_23,In_459);
and U466 (N_466,In_91,In_826);
nand U467 (N_467,In_730,In_218);
xnor U468 (N_468,In_44,In_254);
and U469 (N_469,In_867,In_587);
and U470 (N_470,In_791,In_851);
nor U471 (N_471,In_434,In_821);
nand U472 (N_472,In_348,In_366);
or U473 (N_473,In_347,In_86);
nor U474 (N_474,In_222,In_988);
nor U475 (N_475,In_545,In_886);
nand U476 (N_476,In_453,In_689);
and U477 (N_477,In_664,In_592);
nor U478 (N_478,In_7,In_889);
or U479 (N_479,In_657,In_600);
and U480 (N_480,In_429,In_173);
nor U481 (N_481,In_69,In_237);
nand U482 (N_482,In_951,In_492);
nor U483 (N_483,In_790,In_310);
or U484 (N_484,In_83,In_181);
xor U485 (N_485,In_634,In_382);
and U486 (N_486,In_812,In_963);
nand U487 (N_487,In_35,In_630);
and U488 (N_488,In_733,In_179);
or U489 (N_489,In_368,In_621);
nor U490 (N_490,In_82,In_706);
nor U491 (N_491,In_424,In_203);
and U492 (N_492,In_43,In_663);
and U493 (N_493,In_204,In_451);
nand U494 (N_494,In_955,In_885);
nor U495 (N_495,In_180,In_62);
xor U496 (N_496,In_921,In_896);
or U497 (N_497,In_633,In_820);
and U498 (N_498,In_455,In_720);
nor U499 (N_499,In_581,In_34);
or U500 (N_500,In_992,In_259);
nor U501 (N_501,In_546,In_878);
nor U502 (N_502,In_461,In_816);
and U503 (N_503,In_811,In_847);
nor U504 (N_504,In_284,In_360);
or U505 (N_505,In_819,In_831);
or U506 (N_506,In_603,In_636);
nand U507 (N_507,In_406,In_339);
or U508 (N_508,In_302,In_333);
nand U509 (N_509,In_170,In_494);
or U510 (N_510,In_377,In_541);
nor U511 (N_511,In_309,In_726);
xnor U512 (N_512,In_229,In_769);
nor U513 (N_513,In_119,In_958);
and U514 (N_514,In_630,In_762);
nand U515 (N_515,In_53,In_295);
and U516 (N_516,In_330,In_941);
and U517 (N_517,In_246,In_601);
or U518 (N_518,In_473,In_160);
or U519 (N_519,In_588,In_285);
and U520 (N_520,In_93,In_812);
and U521 (N_521,In_805,In_528);
nor U522 (N_522,In_350,In_953);
nor U523 (N_523,In_118,In_370);
nor U524 (N_524,In_549,In_427);
and U525 (N_525,In_521,In_418);
and U526 (N_526,In_702,In_519);
nand U527 (N_527,In_53,In_784);
nor U528 (N_528,In_310,In_120);
nand U529 (N_529,In_331,In_222);
and U530 (N_530,In_736,In_329);
or U531 (N_531,In_762,In_742);
and U532 (N_532,In_418,In_112);
and U533 (N_533,In_579,In_454);
and U534 (N_534,In_297,In_281);
and U535 (N_535,In_193,In_991);
and U536 (N_536,In_746,In_264);
and U537 (N_537,In_224,In_637);
and U538 (N_538,In_366,In_880);
and U539 (N_539,In_503,In_99);
nor U540 (N_540,In_263,In_334);
or U541 (N_541,In_334,In_234);
nand U542 (N_542,In_382,In_68);
and U543 (N_543,In_734,In_877);
and U544 (N_544,In_563,In_466);
nor U545 (N_545,In_776,In_470);
and U546 (N_546,In_259,In_34);
or U547 (N_547,In_359,In_461);
nor U548 (N_548,In_538,In_16);
nand U549 (N_549,In_529,In_341);
nor U550 (N_550,In_771,In_465);
nor U551 (N_551,In_661,In_181);
or U552 (N_552,In_615,In_318);
nand U553 (N_553,In_14,In_1);
or U554 (N_554,In_484,In_368);
or U555 (N_555,In_177,In_64);
xor U556 (N_556,In_564,In_385);
nor U557 (N_557,In_104,In_166);
nor U558 (N_558,In_766,In_967);
nor U559 (N_559,In_50,In_907);
nand U560 (N_560,In_425,In_706);
or U561 (N_561,In_66,In_913);
nand U562 (N_562,In_489,In_365);
or U563 (N_563,In_392,In_362);
nor U564 (N_564,In_401,In_3);
nand U565 (N_565,In_529,In_573);
nor U566 (N_566,In_785,In_313);
nor U567 (N_567,In_191,In_213);
and U568 (N_568,In_394,In_344);
nand U569 (N_569,In_248,In_65);
nor U570 (N_570,In_228,In_761);
or U571 (N_571,In_446,In_480);
or U572 (N_572,In_824,In_798);
nand U573 (N_573,In_135,In_678);
or U574 (N_574,In_846,In_792);
nor U575 (N_575,In_647,In_990);
nand U576 (N_576,In_237,In_969);
nand U577 (N_577,In_633,In_700);
xor U578 (N_578,In_312,In_8);
nand U579 (N_579,In_143,In_20);
and U580 (N_580,In_159,In_608);
or U581 (N_581,In_394,In_322);
or U582 (N_582,In_20,In_538);
or U583 (N_583,In_835,In_100);
nand U584 (N_584,In_659,In_141);
or U585 (N_585,In_845,In_377);
or U586 (N_586,In_528,In_175);
nand U587 (N_587,In_899,In_558);
nor U588 (N_588,In_498,In_911);
or U589 (N_589,In_194,In_914);
or U590 (N_590,In_565,In_115);
nand U591 (N_591,In_826,In_655);
nand U592 (N_592,In_963,In_445);
or U593 (N_593,In_247,In_64);
and U594 (N_594,In_891,In_430);
nand U595 (N_595,In_392,In_384);
nand U596 (N_596,In_843,In_656);
nand U597 (N_597,In_98,In_167);
or U598 (N_598,In_270,In_339);
nand U599 (N_599,In_238,In_295);
or U600 (N_600,In_150,In_932);
or U601 (N_601,In_770,In_352);
nand U602 (N_602,In_596,In_487);
xor U603 (N_603,In_150,In_537);
nor U604 (N_604,In_397,In_602);
and U605 (N_605,In_45,In_502);
nor U606 (N_606,In_284,In_471);
nand U607 (N_607,In_867,In_451);
and U608 (N_608,In_326,In_321);
or U609 (N_609,In_936,In_304);
nand U610 (N_610,In_332,In_914);
nor U611 (N_611,In_298,In_409);
nand U612 (N_612,In_959,In_99);
or U613 (N_613,In_42,In_677);
xor U614 (N_614,In_634,In_496);
and U615 (N_615,In_878,In_693);
nor U616 (N_616,In_412,In_782);
nor U617 (N_617,In_53,In_950);
and U618 (N_618,In_224,In_348);
and U619 (N_619,In_17,In_163);
and U620 (N_620,In_633,In_354);
nor U621 (N_621,In_239,In_148);
or U622 (N_622,In_609,In_562);
nand U623 (N_623,In_7,In_208);
or U624 (N_624,In_47,In_802);
and U625 (N_625,In_470,In_240);
nor U626 (N_626,In_712,In_639);
nand U627 (N_627,In_7,In_257);
nand U628 (N_628,In_983,In_542);
nand U629 (N_629,In_896,In_706);
and U630 (N_630,In_397,In_762);
nand U631 (N_631,In_539,In_505);
nor U632 (N_632,In_55,In_903);
nand U633 (N_633,In_10,In_298);
nor U634 (N_634,In_73,In_34);
nand U635 (N_635,In_100,In_951);
and U636 (N_636,In_684,In_206);
nand U637 (N_637,In_956,In_252);
xor U638 (N_638,In_977,In_522);
or U639 (N_639,In_188,In_173);
nor U640 (N_640,In_757,In_576);
or U641 (N_641,In_890,In_302);
or U642 (N_642,In_720,In_151);
and U643 (N_643,In_611,In_938);
and U644 (N_644,In_582,In_305);
nand U645 (N_645,In_473,In_936);
nand U646 (N_646,In_390,In_442);
nand U647 (N_647,In_895,In_220);
nand U648 (N_648,In_183,In_693);
and U649 (N_649,In_702,In_798);
and U650 (N_650,In_342,In_11);
or U651 (N_651,In_671,In_677);
nor U652 (N_652,In_550,In_903);
nand U653 (N_653,In_423,In_301);
nand U654 (N_654,In_627,In_72);
or U655 (N_655,In_560,In_346);
nand U656 (N_656,In_523,In_855);
nand U657 (N_657,In_456,In_157);
nand U658 (N_658,In_184,In_52);
or U659 (N_659,In_556,In_450);
or U660 (N_660,In_497,In_268);
or U661 (N_661,In_545,In_243);
or U662 (N_662,In_563,In_825);
or U663 (N_663,In_617,In_690);
and U664 (N_664,In_923,In_283);
and U665 (N_665,In_260,In_314);
nor U666 (N_666,In_186,In_182);
nand U667 (N_667,In_30,In_430);
nor U668 (N_668,In_187,In_962);
nand U669 (N_669,In_323,In_110);
nor U670 (N_670,In_813,In_0);
and U671 (N_671,In_417,In_767);
or U672 (N_672,In_11,In_509);
nand U673 (N_673,In_322,In_400);
and U674 (N_674,In_968,In_288);
and U675 (N_675,In_98,In_213);
xor U676 (N_676,In_633,In_799);
or U677 (N_677,In_977,In_394);
and U678 (N_678,In_466,In_148);
nand U679 (N_679,In_825,In_258);
and U680 (N_680,In_801,In_603);
nor U681 (N_681,In_98,In_186);
and U682 (N_682,In_578,In_664);
or U683 (N_683,In_39,In_25);
nand U684 (N_684,In_169,In_318);
or U685 (N_685,In_195,In_42);
xnor U686 (N_686,In_388,In_951);
xnor U687 (N_687,In_784,In_413);
or U688 (N_688,In_973,In_763);
or U689 (N_689,In_144,In_897);
nor U690 (N_690,In_193,In_462);
nand U691 (N_691,In_356,In_720);
and U692 (N_692,In_797,In_431);
nand U693 (N_693,In_983,In_431);
nor U694 (N_694,In_24,In_496);
nor U695 (N_695,In_4,In_877);
and U696 (N_696,In_821,In_679);
nor U697 (N_697,In_755,In_822);
and U698 (N_698,In_247,In_887);
nand U699 (N_699,In_149,In_436);
xnor U700 (N_700,In_881,In_183);
and U701 (N_701,In_459,In_287);
nand U702 (N_702,In_976,In_961);
nor U703 (N_703,In_764,In_314);
or U704 (N_704,In_444,In_91);
or U705 (N_705,In_822,In_348);
and U706 (N_706,In_407,In_828);
and U707 (N_707,In_888,In_16);
or U708 (N_708,In_62,In_768);
nor U709 (N_709,In_372,In_483);
or U710 (N_710,In_268,In_96);
nand U711 (N_711,In_137,In_56);
nor U712 (N_712,In_991,In_199);
and U713 (N_713,In_992,In_467);
nand U714 (N_714,In_989,In_821);
nand U715 (N_715,In_447,In_355);
or U716 (N_716,In_749,In_766);
and U717 (N_717,In_759,In_1);
nor U718 (N_718,In_677,In_712);
and U719 (N_719,In_865,In_653);
nor U720 (N_720,In_491,In_879);
nand U721 (N_721,In_757,In_431);
and U722 (N_722,In_507,In_863);
or U723 (N_723,In_402,In_8);
nand U724 (N_724,In_767,In_497);
nor U725 (N_725,In_674,In_522);
or U726 (N_726,In_387,In_580);
and U727 (N_727,In_146,In_516);
nand U728 (N_728,In_148,In_589);
or U729 (N_729,In_871,In_824);
xnor U730 (N_730,In_407,In_873);
nand U731 (N_731,In_930,In_622);
and U732 (N_732,In_648,In_692);
nor U733 (N_733,In_771,In_535);
nand U734 (N_734,In_965,In_407);
or U735 (N_735,In_507,In_786);
and U736 (N_736,In_529,In_13);
or U737 (N_737,In_246,In_831);
nor U738 (N_738,In_483,In_147);
and U739 (N_739,In_196,In_296);
nor U740 (N_740,In_297,In_790);
or U741 (N_741,In_595,In_506);
nand U742 (N_742,In_211,In_942);
or U743 (N_743,In_178,In_439);
nand U744 (N_744,In_634,In_11);
nor U745 (N_745,In_575,In_373);
xor U746 (N_746,In_825,In_118);
or U747 (N_747,In_73,In_848);
or U748 (N_748,In_281,In_880);
nand U749 (N_749,In_511,In_252);
or U750 (N_750,In_385,In_624);
and U751 (N_751,In_755,In_907);
and U752 (N_752,In_649,In_14);
nand U753 (N_753,In_263,In_138);
or U754 (N_754,In_489,In_829);
nor U755 (N_755,In_74,In_735);
xor U756 (N_756,In_851,In_787);
nand U757 (N_757,In_380,In_182);
nor U758 (N_758,In_544,In_438);
or U759 (N_759,In_120,In_801);
xor U760 (N_760,In_985,In_39);
nor U761 (N_761,In_331,In_948);
nand U762 (N_762,In_610,In_768);
and U763 (N_763,In_821,In_692);
nand U764 (N_764,In_83,In_333);
or U765 (N_765,In_404,In_194);
and U766 (N_766,In_321,In_349);
and U767 (N_767,In_652,In_133);
or U768 (N_768,In_695,In_856);
or U769 (N_769,In_595,In_308);
nor U770 (N_770,In_657,In_583);
and U771 (N_771,In_89,In_798);
and U772 (N_772,In_6,In_535);
nor U773 (N_773,In_251,In_207);
and U774 (N_774,In_637,In_913);
nor U775 (N_775,In_518,In_990);
nor U776 (N_776,In_913,In_118);
and U777 (N_777,In_790,In_140);
and U778 (N_778,In_591,In_908);
nand U779 (N_779,In_396,In_327);
nand U780 (N_780,In_950,In_621);
xnor U781 (N_781,In_871,In_796);
or U782 (N_782,In_65,In_954);
or U783 (N_783,In_725,In_562);
nor U784 (N_784,In_461,In_658);
or U785 (N_785,In_102,In_368);
nor U786 (N_786,In_562,In_699);
nand U787 (N_787,In_686,In_38);
or U788 (N_788,In_450,In_127);
and U789 (N_789,In_710,In_757);
nor U790 (N_790,In_509,In_308);
or U791 (N_791,In_740,In_815);
nor U792 (N_792,In_536,In_600);
or U793 (N_793,In_63,In_654);
and U794 (N_794,In_553,In_526);
or U795 (N_795,In_182,In_171);
or U796 (N_796,In_293,In_318);
or U797 (N_797,In_141,In_886);
nand U798 (N_798,In_541,In_560);
xor U799 (N_799,In_538,In_986);
nand U800 (N_800,In_720,In_848);
or U801 (N_801,In_24,In_904);
nand U802 (N_802,In_172,In_807);
nor U803 (N_803,In_533,In_628);
nor U804 (N_804,In_634,In_925);
nor U805 (N_805,In_998,In_901);
or U806 (N_806,In_418,In_62);
xor U807 (N_807,In_39,In_256);
nor U808 (N_808,In_803,In_936);
nand U809 (N_809,In_96,In_62);
or U810 (N_810,In_718,In_729);
nor U811 (N_811,In_990,In_205);
nor U812 (N_812,In_945,In_263);
nand U813 (N_813,In_702,In_220);
and U814 (N_814,In_799,In_467);
nand U815 (N_815,In_416,In_737);
or U816 (N_816,In_314,In_189);
nor U817 (N_817,In_358,In_101);
or U818 (N_818,In_553,In_232);
nand U819 (N_819,In_149,In_664);
and U820 (N_820,In_444,In_396);
nand U821 (N_821,In_625,In_39);
or U822 (N_822,In_821,In_289);
and U823 (N_823,In_290,In_637);
or U824 (N_824,In_410,In_333);
or U825 (N_825,In_971,In_508);
and U826 (N_826,In_823,In_274);
nor U827 (N_827,In_458,In_786);
or U828 (N_828,In_876,In_123);
and U829 (N_829,In_661,In_573);
nand U830 (N_830,In_947,In_448);
or U831 (N_831,In_730,In_603);
and U832 (N_832,In_414,In_867);
nor U833 (N_833,In_259,In_359);
and U834 (N_834,In_479,In_665);
or U835 (N_835,In_331,In_468);
nor U836 (N_836,In_623,In_622);
nand U837 (N_837,In_389,In_601);
xor U838 (N_838,In_431,In_338);
and U839 (N_839,In_990,In_530);
nand U840 (N_840,In_51,In_372);
and U841 (N_841,In_942,In_725);
and U842 (N_842,In_53,In_291);
or U843 (N_843,In_363,In_883);
xor U844 (N_844,In_564,In_410);
nor U845 (N_845,In_961,In_325);
or U846 (N_846,In_443,In_320);
nor U847 (N_847,In_458,In_733);
nand U848 (N_848,In_536,In_718);
nand U849 (N_849,In_415,In_656);
nand U850 (N_850,In_818,In_861);
or U851 (N_851,In_202,In_988);
or U852 (N_852,In_353,In_205);
nor U853 (N_853,In_167,In_806);
and U854 (N_854,In_540,In_58);
or U855 (N_855,In_626,In_465);
and U856 (N_856,In_275,In_566);
nand U857 (N_857,In_408,In_865);
nor U858 (N_858,In_740,In_549);
and U859 (N_859,In_141,In_613);
nor U860 (N_860,In_110,In_353);
or U861 (N_861,In_874,In_424);
nand U862 (N_862,In_113,In_529);
and U863 (N_863,In_144,In_222);
or U864 (N_864,In_928,In_56);
nor U865 (N_865,In_455,In_430);
and U866 (N_866,In_657,In_414);
nor U867 (N_867,In_480,In_681);
nor U868 (N_868,In_36,In_275);
and U869 (N_869,In_703,In_555);
nand U870 (N_870,In_901,In_927);
and U871 (N_871,In_95,In_554);
or U872 (N_872,In_54,In_356);
and U873 (N_873,In_364,In_773);
or U874 (N_874,In_38,In_850);
nor U875 (N_875,In_171,In_106);
and U876 (N_876,In_835,In_545);
and U877 (N_877,In_802,In_126);
and U878 (N_878,In_737,In_729);
and U879 (N_879,In_907,In_196);
and U880 (N_880,In_839,In_827);
and U881 (N_881,In_939,In_448);
nor U882 (N_882,In_630,In_984);
or U883 (N_883,In_5,In_951);
or U884 (N_884,In_333,In_642);
nor U885 (N_885,In_221,In_882);
nand U886 (N_886,In_60,In_751);
nor U887 (N_887,In_361,In_944);
nor U888 (N_888,In_47,In_131);
or U889 (N_889,In_312,In_260);
nor U890 (N_890,In_221,In_800);
or U891 (N_891,In_799,In_934);
nand U892 (N_892,In_28,In_481);
or U893 (N_893,In_276,In_498);
and U894 (N_894,In_171,In_993);
nor U895 (N_895,In_835,In_792);
and U896 (N_896,In_143,In_16);
and U897 (N_897,In_57,In_740);
and U898 (N_898,In_184,In_828);
nor U899 (N_899,In_296,In_717);
nor U900 (N_900,In_84,In_519);
nand U901 (N_901,In_532,In_572);
nand U902 (N_902,In_654,In_154);
and U903 (N_903,In_580,In_845);
nor U904 (N_904,In_879,In_589);
nand U905 (N_905,In_84,In_215);
nand U906 (N_906,In_855,In_598);
or U907 (N_907,In_172,In_43);
or U908 (N_908,In_63,In_694);
xnor U909 (N_909,In_408,In_872);
and U910 (N_910,In_463,In_353);
nor U911 (N_911,In_220,In_741);
nor U912 (N_912,In_32,In_271);
nor U913 (N_913,In_905,In_580);
nand U914 (N_914,In_715,In_838);
nor U915 (N_915,In_817,In_692);
nand U916 (N_916,In_692,In_311);
or U917 (N_917,In_580,In_479);
nand U918 (N_918,In_624,In_928);
nand U919 (N_919,In_415,In_215);
and U920 (N_920,In_403,In_283);
nor U921 (N_921,In_181,In_828);
nor U922 (N_922,In_798,In_795);
xor U923 (N_923,In_427,In_728);
or U924 (N_924,In_460,In_184);
or U925 (N_925,In_399,In_118);
nor U926 (N_926,In_556,In_275);
or U927 (N_927,In_999,In_23);
xnor U928 (N_928,In_753,In_213);
xnor U929 (N_929,In_882,In_659);
or U930 (N_930,In_837,In_997);
or U931 (N_931,In_196,In_313);
nand U932 (N_932,In_609,In_892);
or U933 (N_933,In_117,In_829);
nor U934 (N_934,In_145,In_665);
nand U935 (N_935,In_880,In_769);
nor U936 (N_936,In_31,In_999);
nand U937 (N_937,In_522,In_612);
nand U938 (N_938,In_725,In_390);
nand U939 (N_939,In_894,In_681);
or U940 (N_940,In_682,In_263);
nor U941 (N_941,In_429,In_251);
or U942 (N_942,In_752,In_630);
nand U943 (N_943,In_49,In_395);
nand U944 (N_944,In_617,In_318);
and U945 (N_945,In_783,In_215);
and U946 (N_946,In_715,In_880);
xnor U947 (N_947,In_252,In_310);
nand U948 (N_948,In_180,In_582);
xor U949 (N_949,In_106,In_213);
nand U950 (N_950,In_614,In_684);
nand U951 (N_951,In_150,In_51);
xor U952 (N_952,In_657,In_395);
nor U953 (N_953,In_165,In_796);
or U954 (N_954,In_719,In_480);
nor U955 (N_955,In_91,In_539);
nor U956 (N_956,In_221,In_179);
xor U957 (N_957,In_876,In_411);
or U958 (N_958,In_874,In_360);
and U959 (N_959,In_872,In_579);
nand U960 (N_960,In_750,In_889);
or U961 (N_961,In_591,In_572);
and U962 (N_962,In_277,In_464);
and U963 (N_963,In_236,In_446);
and U964 (N_964,In_790,In_860);
or U965 (N_965,In_995,In_356);
nor U966 (N_966,In_325,In_320);
and U967 (N_967,In_591,In_506);
nor U968 (N_968,In_303,In_912);
and U969 (N_969,In_596,In_261);
and U970 (N_970,In_479,In_324);
nand U971 (N_971,In_570,In_523);
or U972 (N_972,In_949,In_749);
nand U973 (N_973,In_715,In_716);
and U974 (N_974,In_298,In_364);
nand U975 (N_975,In_467,In_29);
nor U976 (N_976,In_105,In_20);
or U977 (N_977,In_73,In_716);
nor U978 (N_978,In_705,In_91);
nor U979 (N_979,In_998,In_428);
or U980 (N_980,In_621,In_16);
or U981 (N_981,In_461,In_260);
or U982 (N_982,In_937,In_319);
nor U983 (N_983,In_938,In_388);
nor U984 (N_984,In_33,In_989);
or U985 (N_985,In_744,In_36);
nand U986 (N_986,In_548,In_204);
or U987 (N_987,In_858,In_54);
and U988 (N_988,In_602,In_277);
and U989 (N_989,In_847,In_95);
nor U990 (N_990,In_476,In_948);
nor U991 (N_991,In_612,In_165);
or U992 (N_992,In_344,In_860);
or U993 (N_993,In_55,In_474);
or U994 (N_994,In_58,In_507);
or U995 (N_995,In_952,In_658);
and U996 (N_996,In_383,In_881);
nand U997 (N_997,In_345,In_652);
or U998 (N_998,In_25,In_588);
nor U999 (N_999,In_871,In_23);
nand U1000 (N_1000,In_972,In_542);
and U1001 (N_1001,In_785,In_377);
and U1002 (N_1002,In_16,In_132);
nor U1003 (N_1003,In_26,In_34);
nor U1004 (N_1004,In_566,In_782);
nor U1005 (N_1005,In_168,In_931);
or U1006 (N_1006,In_194,In_953);
nand U1007 (N_1007,In_729,In_931);
and U1008 (N_1008,In_674,In_690);
or U1009 (N_1009,In_514,In_672);
nand U1010 (N_1010,In_583,In_658);
nor U1011 (N_1011,In_955,In_914);
nor U1012 (N_1012,In_271,In_976);
and U1013 (N_1013,In_270,In_671);
nand U1014 (N_1014,In_820,In_212);
nand U1015 (N_1015,In_175,In_49);
nand U1016 (N_1016,In_992,In_479);
nand U1017 (N_1017,In_795,In_579);
nand U1018 (N_1018,In_223,In_373);
nor U1019 (N_1019,In_551,In_932);
nor U1020 (N_1020,In_255,In_349);
nor U1021 (N_1021,In_321,In_103);
or U1022 (N_1022,In_977,In_581);
nand U1023 (N_1023,In_494,In_821);
and U1024 (N_1024,In_725,In_288);
nand U1025 (N_1025,In_334,In_861);
and U1026 (N_1026,In_258,In_454);
and U1027 (N_1027,In_504,In_383);
nand U1028 (N_1028,In_381,In_114);
and U1029 (N_1029,In_26,In_585);
nor U1030 (N_1030,In_891,In_375);
nand U1031 (N_1031,In_741,In_594);
and U1032 (N_1032,In_171,In_455);
nand U1033 (N_1033,In_842,In_228);
nand U1034 (N_1034,In_867,In_331);
and U1035 (N_1035,In_164,In_854);
nand U1036 (N_1036,In_834,In_6);
and U1037 (N_1037,In_798,In_417);
or U1038 (N_1038,In_881,In_581);
or U1039 (N_1039,In_802,In_923);
nor U1040 (N_1040,In_447,In_737);
and U1041 (N_1041,In_992,In_553);
nand U1042 (N_1042,In_975,In_366);
or U1043 (N_1043,In_270,In_531);
nand U1044 (N_1044,In_966,In_45);
nand U1045 (N_1045,In_604,In_48);
and U1046 (N_1046,In_588,In_182);
or U1047 (N_1047,In_625,In_24);
nor U1048 (N_1048,In_310,In_210);
nand U1049 (N_1049,In_130,In_465);
or U1050 (N_1050,In_19,In_820);
nor U1051 (N_1051,In_333,In_377);
nand U1052 (N_1052,In_339,In_348);
nor U1053 (N_1053,In_817,In_489);
and U1054 (N_1054,In_70,In_775);
nand U1055 (N_1055,In_175,In_707);
and U1056 (N_1056,In_315,In_454);
nand U1057 (N_1057,In_556,In_381);
and U1058 (N_1058,In_409,In_922);
and U1059 (N_1059,In_643,In_614);
and U1060 (N_1060,In_542,In_507);
nor U1061 (N_1061,In_584,In_622);
nor U1062 (N_1062,In_94,In_583);
nor U1063 (N_1063,In_919,In_406);
xnor U1064 (N_1064,In_621,In_441);
and U1065 (N_1065,In_766,In_817);
or U1066 (N_1066,In_721,In_39);
and U1067 (N_1067,In_870,In_610);
nor U1068 (N_1068,In_385,In_658);
or U1069 (N_1069,In_81,In_874);
nor U1070 (N_1070,In_889,In_262);
or U1071 (N_1071,In_616,In_189);
nor U1072 (N_1072,In_413,In_462);
or U1073 (N_1073,In_747,In_994);
and U1074 (N_1074,In_839,In_684);
nor U1075 (N_1075,In_388,In_323);
nor U1076 (N_1076,In_96,In_613);
nand U1077 (N_1077,In_360,In_702);
or U1078 (N_1078,In_113,In_586);
nand U1079 (N_1079,In_476,In_846);
nand U1080 (N_1080,In_426,In_221);
and U1081 (N_1081,In_475,In_346);
nand U1082 (N_1082,In_12,In_611);
nand U1083 (N_1083,In_663,In_950);
or U1084 (N_1084,In_578,In_672);
and U1085 (N_1085,In_286,In_266);
or U1086 (N_1086,In_498,In_398);
nand U1087 (N_1087,In_892,In_153);
nand U1088 (N_1088,In_186,In_54);
nand U1089 (N_1089,In_692,In_445);
nor U1090 (N_1090,In_0,In_249);
or U1091 (N_1091,In_958,In_136);
nor U1092 (N_1092,In_146,In_598);
or U1093 (N_1093,In_895,In_876);
and U1094 (N_1094,In_473,In_899);
nand U1095 (N_1095,In_176,In_284);
or U1096 (N_1096,In_358,In_213);
nor U1097 (N_1097,In_59,In_291);
or U1098 (N_1098,In_265,In_936);
nand U1099 (N_1099,In_997,In_638);
and U1100 (N_1100,In_842,In_958);
nor U1101 (N_1101,In_874,In_207);
nand U1102 (N_1102,In_271,In_593);
nor U1103 (N_1103,In_122,In_843);
or U1104 (N_1104,In_337,In_469);
xnor U1105 (N_1105,In_663,In_703);
or U1106 (N_1106,In_540,In_881);
and U1107 (N_1107,In_18,In_540);
nand U1108 (N_1108,In_230,In_490);
or U1109 (N_1109,In_229,In_476);
nor U1110 (N_1110,In_638,In_740);
or U1111 (N_1111,In_648,In_952);
nor U1112 (N_1112,In_849,In_732);
nor U1113 (N_1113,In_112,In_251);
and U1114 (N_1114,In_282,In_422);
nor U1115 (N_1115,In_106,In_100);
nor U1116 (N_1116,In_982,In_65);
nor U1117 (N_1117,In_721,In_133);
or U1118 (N_1118,In_148,In_943);
nor U1119 (N_1119,In_140,In_751);
nand U1120 (N_1120,In_802,In_999);
and U1121 (N_1121,In_545,In_346);
or U1122 (N_1122,In_601,In_355);
nand U1123 (N_1123,In_316,In_477);
nand U1124 (N_1124,In_466,In_520);
nand U1125 (N_1125,In_223,In_527);
or U1126 (N_1126,In_572,In_103);
or U1127 (N_1127,In_163,In_362);
xor U1128 (N_1128,In_750,In_188);
nand U1129 (N_1129,In_153,In_307);
or U1130 (N_1130,In_235,In_547);
nand U1131 (N_1131,In_850,In_389);
or U1132 (N_1132,In_796,In_738);
or U1133 (N_1133,In_147,In_922);
nand U1134 (N_1134,In_613,In_358);
or U1135 (N_1135,In_437,In_683);
or U1136 (N_1136,In_105,In_233);
nor U1137 (N_1137,In_629,In_55);
or U1138 (N_1138,In_733,In_448);
or U1139 (N_1139,In_986,In_85);
or U1140 (N_1140,In_959,In_634);
or U1141 (N_1141,In_893,In_228);
nand U1142 (N_1142,In_623,In_503);
nand U1143 (N_1143,In_954,In_490);
or U1144 (N_1144,In_742,In_588);
nor U1145 (N_1145,In_976,In_973);
nand U1146 (N_1146,In_587,In_891);
nand U1147 (N_1147,In_465,In_640);
nand U1148 (N_1148,In_264,In_137);
and U1149 (N_1149,In_196,In_383);
nor U1150 (N_1150,In_555,In_325);
nor U1151 (N_1151,In_355,In_237);
nor U1152 (N_1152,In_404,In_344);
and U1153 (N_1153,In_176,In_738);
nor U1154 (N_1154,In_73,In_382);
nand U1155 (N_1155,In_478,In_776);
and U1156 (N_1156,In_49,In_896);
nand U1157 (N_1157,In_861,In_735);
or U1158 (N_1158,In_277,In_392);
and U1159 (N_1159,In_58,In_768);
nand U1160 (N_1160,In_205,In_926);
or U1161 (N_1161,In_993,In_79);
nor U1162 (N_1162,In_504,In_698);
and U1163 (N_1163,In_784,In_773);
nor U1164 (N_1164,In_973,In_659);
nor U1165 (N_1165,In_441,In_808);
or U1166 (N_1166,In_822,In_32);
and U1167 (N_1167,In_409,In_823);
or U1168 (N_1168,In_537,In_493);
or U1169 (N_1169,In_548,In_886);
or U1170 (N_1170,In_762,In_306);
nor U1171 (N_1171,In_347,In_363);
nor U1172 (N_1172,In_971,In_942);
and U1173 (N_1173,In_401,In_612);
or U1174 (N_1174,In_150,In_914);
nor U1175 (N_1175,In_215,In_942);
nor U1176 (N_1176,In_291,In_862);
nor U1177 (N_1177,In_909,In_678);
nor U1178 (N_1178,In_729,In_944);
or U1179 (N_1179,In_891,In_827);
and U1180 (N_1180,In_937,In_236);
nand U1181 (N_1181,In_207,In_783);
or U1182 (N_1182,In_460,In_828);
and U1183 (N_1183,In_896,In_738);
nor U1184 (N_1184,In_571,In_673);
or U1185 (N_1185,In_687,In_403);
or U1186 (N_1186,In_89,In_91);
or U1187 (N_1187,In_924,In_466);
or U1188 (N_1188,In_402,In_894);
xnor U1189 (N_1189,In_750,In_513);
or U1190 (N_1190,In_950,In_336);
and U1191 (N_1191,In_261,In_741);
and U1192 (N_1192,In_756,In_439);
or U1193 (N_1193,In_465,In_276);
and U1194 (N_1194,In_280,In_808);
nor U1195 (N_1195,In_595,In_729);
and U1196 (N_1196,In_223,In_576);
and U1197 (N_1197,In_763,In_837);
and U1198 (N_1198,In_312,In_503);
or U1199 (N_1199,In_458,In_959);
and U1200 (N_1200,In_903,In_815);
and U1201 (N_1201,In_146,In_172);
and U1202 (N_1202,In_406,In_39);
nand U1203 (N_1203,In_512,In_441);
nand U1204 (N_1204,In_961,In_361);
or U1205 (N_1205,In_509,In_950);
and U1206 (N_1206,In_556,In_768);
and U1207 (N_1207,In_318,In_686);
or U1208 (N_1208,In_19,In_9);
and U1209 (N_1209,In_349,In_837);
and U1210 (N_1210,In_824,In_636);
nor U1211 (N_1211,In_76,In_541);
or U1212 (N_1212,In_864,In_897);
xnor U1213 (N_1213,In_690,In_983);
and U1214 (N_1214,In_45,In_82);
nand U1215 (N_1215,In_315,In_520);
or U1216 (N_1216,In_273,In_629);
or U1217 (N_1217,In_858,In_978);
nor U1218 (N_1218,In_58,In_555);
or U1219 (N_1219,In_375,In_146);
or U1220 (N_1220,In_564,In_489);
nand U1221 (N_1221,In_537,In_354);
nand U1222 (N_1222,In_493,In_729);
xor U1223 (N_1223,In_647,In_568);
or U1224 (N_1224,In_169,In_613);
nand U1225 (N_1225,In_839,In_237);
nor U1226 (N_1226,In_762,In_687);
nand U1227 (N_1227,In_415,In_296);
or U1228 (N_1228,In_576,In_183);
nor U1229 (N_1229,In_397,In_507);
or U1230 (N_1230,In_319,In_673);
nand U1231 (N_1231,In_93,In_211);
and U1232 (N_1232,In_697,In_126);
xor U1233 (N_1233,In_814,In_928);
or U1234 (N_1234,In_962,In_834);
nor U1235 (N_1235,In_834,In_474);
or U1236 (N_1236,In_849,In_857);
nor U1237 (N_1237,In_317,In_910);
nor U1238 (N_1238,In_115,In_739);
nand U1239 (N_1239,In_22,In_244);
and U1240 (N_1240,In_433,In_485);
nor U1241 (N_1241,In_681,In_523);
and U1242 (N_1242,In_334,In_289);
and U1243 (N_1243,In_519,In_71);
and U1244 (N_1244,In_473,In_975);
and U1245 (N_1245,In_655,In_193);
and U1246 (N_1246,In_825,In_805);
or U1247 (N_1247,In_388,In_779);
nand U1248 (N_1248,In_775,In_784);
or U1249 (N_1249,In_742,In_748);
or U1250 (N_1250,In_126,In_139);
nor U1251 (N_1251,In_55,In_344);
nor U1252 (N_1252,In_414,In_164);
nor U1253 (N_1253,In_84,In_707);
nor U1254 (N_1254,In_972,In_119);
nor U1255 (N_1255,In_104,In_321);
xnor U1256 (N_1256,In_941,In_580);
and U1257 (N_1257,In_840,In_819);
and U1258 (N_1258,In_641,In_900);
or U1259 (N_1259,In_158,In_17);
nor U1260 (N_1260,In_898,In_747);
nand U1261 (N_1261,In_208,In_301);
and U1262 (N_1262,In_986,In_981);
or U1263 (N_1263,In_13,In_585);
nand U1264 (N_1264,In_944,In_95);
nor U1265 (N_1265,In_585,In_903);
nor U1266 (N_1266,In_544,In_381);
or U1267 (N_1267,In_311,In_4);
or U1268 (N_1268,In_194,In_245);
nand U1269 (N_1269,In_300,In_960);
or U1270 (N_1270,In_990,In_352);
nand U1271 (N_1271,In_168,In_296);
nor U1272 (N_1272,In_618,In_205);
and U1273 (N_1273,In_365,In_604);
or U1274 (N_1274,In_425,In_70);
nor U1275 (N_1275,In_629,In_758);
and U1276 (N_1276,In_584,In_669);
nor U1277 (N_1277,In_378,In_157);
xor U1278 (N_1278,In_358,In_233);
and U1279 (N_1279,In_788,In_910);
or U1280 (N_1280,In_967,In_791);
nand U1281 (N_1281,In_525,In_889);
nor U1282 (N_1282,In_406,In_22);
nor U1283 (N_1283,In_280,In_142);
or U1284 (N_1284,In_85,In_325);
nand U1285 (N_1285,In_100,In_463);
and U1286 (N_1286,In_882,In_479);
and U1287 (N_1287,In_454,In_590);
nor U1288 (N_1288,In_942,In_200);
or U1289 (N_1289,In_409,In_561);
and U1290 (N_1290,In_880,In_781);
and U1291 (N_1291,In_474,In_117);
and U1292 (N_1292,In_768,In_100);
nand U1293 (N_1293,In_786,In_933);
and U1294 (N_1294,In_135,In_422);
nor U1295 (N_1295,In_691,In_293);
xor U1296 (N_1296,In_35,In_841);
nor U1297 (N_1297,In_488,In_119);
nor U1298 (N_1298,In_906,In_580);
and U1299 (N_1299,In_157,In_502);
and U1300 (N_1300,In_157,In_539);
or U1301 (N_1301,In_424,In_559);
and U1302 (N_1302,In_629,In_605);
nand U1303 (N_1303,In_393,In_897);
and U1304 (N_1304,In_99,In_203);
nand U1305 (N_1305,In_595,In_357);
or U1306 (N_1306,In_519,In_305);
nor U1307 (N_1307,In_420,In_186);
nor U1308 (N_1308,In_557,In_308);
nand U1309 (N_1309,In_14,In_973);
and U1310 (N_1310,In_292,In_565);
and U1311 (N_1311,In_181,In_696);
or U1312 (N_1312,In_727,In_577);
or U1313 (N_1313,In_676,In_586);
or U1314 (N_1314,In_0,In_972);
and U1315 (N_1315,In_660,In_112);
or U1316 (N_1316,In_437,In_622);
and U1317 (N_1317,In_945,In_749);
xor U1318 (N_1318,In_272,In_415);
or U1319 (N_1319,In_240,In_462);
nor U1320 (N_1320,In_26,In_292);
and U1321 (N_1321,In_992,In_632);
nand U1322 (N_1322,In_675,In_558);
or U1323 (N_1323,In_946,In_306);
nand U1324 (N_1324,In_988,In_809);
nand U1325 (N_1325,In_705,In_439);
xnor U1326 (N_1326,In_714,In_9);
nor U1327 (N_1327,In_322,In_692);
nand U1328 (N_1328,In_637,In_398);
nand U1329 (N_1329,In_252,In_179);
nor U1330 (N_1330,In_813,In_882);
xor U1331 (N_1331,In_522,In_339);
nand U1332 (N_1332,In_101,In_370);
or U1333 (N_1333,In_682,In_542);
and U1334 (N_1334,In_520,In_958);
nand U1335 (N_1335,In_507,In_580);
nor U1336 (N_1336,In_841,In_199);
and U1337 (N_1337,In_1,In_517);
or U1338 (N_1338,In_437,In_419);
nor U1339 (N_1339,In_862,In_471);
nand U1340 (N_1340,In_216,In_76);
nand U1341 (N_1341,In_451,In_61);
or U1342 (N_1342,In_855,In_998);
and U1343 (N_1343,In_72,In_234);
and U1344 (N_1344,In_99,In_197);
and U1345 (N_1345,In_24,In_431);
nor U1346 (N_1346,In_858,In_194);
or U1347 (N_1347,In_781,In_196);
nand U1348 (N_1348,In_670,In_948);
xor U1349 (N_1349,In_592,In_385);
or U1350 (N_1350,In_53,In_347);
nor U1351 (N_1351,In_998,In_621);
and U1352 (N_1352,In_967,In_645);
nor U1353 (N_1353,In_1,In_946);
nand U1354 (N_1354,In_777,In_72);
and U1355 (N_1355,In_414,In_415);
and U1356 (N_1356,In_94,In_952);
and U1357 (N_1357,In_628,In_374);
nand U1358 (N_1358,In_417,In_750);
nor U1359 (N_1359,In_571,In_525);
nor U1360 (N_1360,In_769,In_964);
or U1361 (N_1361,In_293,In_913);
xnor U1362 (N_1362,In_214,In_681);
or U1363 (N_1363,In_272,In_527);
nor U1364 (N_1364,In_576,In_730);
nor U1365 (N_1365,In_648,In_600);
nand U1366 (N_1366,In_756,In_904);
and U1367 (N_1367,In_917,In_624);
or U1368 (N_1368,In_181,In_488);
or U1369 (N_1369,In_947,In_944);
and U1370 (N_1370,In_602,In_481);
and U1371 (N_1371,In_155,In_89);
nand U1372 (N_1372,In_309,In_986);
and U1373 (N_1373,In_312,In_980);
and U1374 (N_1374,In_257,In_824);
or U1375 (N_1375,In_751,In_8);
nor U1376 (N_1376,In_234,In_73);
and U1377 (N_1377,In_932,In_692);
nand U1378 (N_1378,In_201,In_386);
or U1379 (N_1379,In_606,In_883);
or U1380 (N_1380,In_267,In_175);
and U1381 (N_1381,In_306,In_516);
and U1382 (N_1382,In_596,In_404);
nand U1383 (N_1383,In_801,In_562);
nor U1384 (N_1384,In_374,In_156);
and U1385 (N_1385,In_573,In_903);
xnor U1386 (N_1386,In_336,In_533);
or U1387 (N_1387,In_455,In_591);
and U1388 (N_1388,In_977,In_849);
and U1389 (N_1389,In_243,In_944);
nand U1390 (N_1390,In_678,In_140);
and U1391 (N_1391,In_479,In_768);
nor U1392 (N_1392,In_468,In_190);
nand U1393 (N_1393,In_952,In_61);
and U1394 (N_1394,In_74,In_429);
or U1395 (N_1395,In_312,In_680);
nand U1396 (N_1396,In_296,In_731);
or U1397 (N_1397,In_99,In_193);
nand U1398 (N_1398,In_355,In_478);
nor U1399 (N_1399,In_914,In_403);
nand U1400 (N_1400,In_757,In_383);
and U1401 (N_1401,In_174,In_572);
nand U1402 (N_1402,In_369,In_269);
nor U1403 (N_1403,In_233,In_415);
and U1404 (N_1404,In_614,In_427);
and U1405 (N_1405,In_492,In_673);
and U1406 (N_1406,In_703,In_330);
and U1407 (N_1407,In_496,In_934);
nand U1408 (N_1408,In_734,In_283);
nor U1409 (N_1409,In_764,In_734);
nor U1410 (N_1410,In_606,In_29);
nor U1411 (N_1411,In_612,In_814);
nor U1412 (N_1412,In_470,In_498);
and U1413 (N_1413,In_827,In_647);
and U1414 (N_1414,In_510,In_431);
nand U1415 (N_1415,In_426,In_192);
nand U1416 (N_1416,In_275,In_735);
nand U1417 (N_1417,In_164,In_981);
nor U1418 (N_1418,In_580,In_583);
or U1419 (N_1419,In_940,In_341);
or U1420 (N_1420,In_387,In_694);
and U1421 (N_1421,In_481,In_486);
nand U1422 (N_1422,In_109,In_697);
nor U1423 (N_1423,In_854,In_267);
nand U1424 (N_1424,In_714,In_982);
and U1425 (N_1425,In_731,In_396);
or U1426 (N_1426,In_47,In_376);
and U1427 (N_1427,In_904,In_169);
nor U1428 (N_1428,In_303,In_909);
nor U1429 (N_1429,In_120,In_645);
or U1430 (N_1430,In_355,In_406);
and U1431 (N_1431,In_196,In_773);
or U1432 (N_1432,In_485,In_161);
and U1433 (N_1433,In_673,In_525);
nor U1434 (N_1434,In_835,In_254);
nor U1435 (N_1435,In_282,In_794);
and U1436 (N_1436,In_27,In_308);
nand U1437 (N_1437,In_639,In_566);
or U1438 (N_1438,In_254,In_969);
or U1439 (N_1439,In_786,In_789);
nor U1440 (N_1440,In_896,In_82);
or U1441 (N_1441,In_457,In_620);
or U1442 (N_1442,In_382,In_446);
and U1443 (N_1443,In_801,In_699);
and U1444 (N_1444,In_451,In_5);
nor U1445 (N_1445,In_50,In_869);
or U1446 (N_1446,In_945,In_152);
nand U1447 (N_1447,In_584,In_589);
or U1448 (N_1448,In_470,In_952);
nand U1449 (N_1449,In_353,In_207);
nor U1450 (N_1450,In_53,In_885);
nor U1451 (N_1451,In_708,In_402);
or U1452 (N_1452,In_340,In_678);
nor U1453 (N_1453,In_671,In_668);
nand U1454 (N_1454,In_737,In_309);
nor U1455 (N_1455,In_86,In_221);
and U1456 (N_1456,In_149,In_604);
or U1457 (N_1457,In_587,In_43);
and U1458 (N_1458,In_909,In_396);
or U1459 (N_1459,In_28,In_818);
or U1460 (N_1460,In_818,In_239);
or U1461 (N_1461,In_440,In_73);
or U1462 (N_1462,In_503,In_31);
nor U1463 (N_1463,In_148,In_812);
nand U1464 (N_1464,In_423,In_284);
or U1465 (N_1465,In_996,In_37);
and U1466 (N_1466,In_172,In_526);
nand U1467 (N_1467,In_163,In_912);
and U1468 (N_1468,In_706,In_71);
nand U1469 (N_1469,In_990,In_417);
nor U1470 (N_1470,In_29,In_517);
or U1471 (N_1471,In_639,In_798);
nand U1472 (N_1472,In_537,In_61);
nand U1473 (N_1473,In_353,In_200);
nand U1474 (N_1474,In_21,In_470);
nor U1475 (N_1475,In_234,In_177);
nor U1476 (N_1476,In_592,In_740);
and U1477 (N_1477,In_126,In_538);
and U1478 (N_1478,In_807,In_624);
or U1479 (N_1479,In_146,In_24);
and U1480 (N_1480,In_972,In_743);
nand U1481 (N_1481,In_191,In_12);
or U1482 (N_1482,In_534,In_619);
or U1483 (N_1483,In_97,In_350);
nor U1484 (N_1484,In_396,In_35);
nor U1485 (N_1485,In_611,In_187);
and U1486 (N_1486,In_219,In_431);
nor U1487 (N_1487,In_524,In_835);
or U1488 (N_1488,In_615,In_908);
and U1489 (N_1489,In_929,In_794);
nand U1490 (N_1490,In_507,In_555);
nand U1491 (N_1491,In_990,In_634);
nor U1492 (N_1492,In_474,In_163);
nand U1493 (N_1493,In_588,In_460);
nor U1494 (N_1494,In_280,In_286);
or U1495 (N_1495,In_191,In_265);
or U1496 (N_1496,In_704,In_491);
xnor U1497 (N_1497,In_429,In_761);
nand U1498 (N_1498,In_754,In_113);
nor U1499 (N_1499,In_429,In_755);
and U1500 (N_1500,In_610,In_892);
nor U1501 (N_1501,In_53,In_393);
nor U1502 (N_1502,In_759,In_112);
and U1503 (N_1503,In_348,In_901);
or U1504 (N_1504,In_93,In_491);
and U1505 (N_1505,In_794,In_849);
and U1506 (N_1506,In_234,In_548);
or U1507 (N_1507,In_798,In_700);
or U1508 (N_1508,In_398,In_808);
nor U1509 (N_1509,In_97,In_142);
and U1510 (N_1510,In_97,In_226);
nor U1511 (N_1511,In_541,In_238);
or U1512 (N_1512,In_381,In_605);
nor U1513 (N_1513,In_836,In_41);
nand U1514 (N_1514,In_215,In_989);
nor U1515 (N_1515,In_474,In_83);
nand U1516 (N_1516,In_568,In_698);
or U1517 (N_1517,In_474,In_823);
nor U1518 (N_1518,In_410,In_54);
nand U1519 (N_1519,In_967,In_316);
nor U1520 (N_1520,In_860,In_432);
and U1521 (N_1521,In_711,In_287);
xnor U1522 (N_1522,In_259,In_980);
or U1523 (N_1523,In_712,In_359);
and U1524 (N_1524,In_921,In_93);
and U1525 (N_1525,In_718,In_253);
nor U1526 (N_1526,In_800,In_865);
or U1527 (N_1527,In_455,In_260);
nor U1528 (N_1528,In_319,In_419);
nand U1529 (N_1529,In_929,In_386);
or U1530 (N_1530,In_948,In_448);
and U1531 (N_1531,In_710,In_681);
and U1532 (N_1532,In_165,In_671);
nor U1533 (N_1533,In_542,In_219);
nor U1534 (N_1534,In_620,In_173);
and U1535 (N_1535,In_814,In_570);
or U1536 (N_1536,In_56,In_868);
nor U1537 (N_1537,In_339,In_164);
or U1538 (N_1538,In_433,In_16);
and U1539 (N_1539,In_980,In_6);
nand U1540 (N_1540,In_872,In_697);
or U1541 (N_1541,In_558,In_888);
nor U1542 (N_1542,In_363,In_86);
or U1543 (N_1543,In_355,In_52);
and U1544 (N_1544,In_60,In_510);
or U1545 (N_1545,In_518,In_54);
nand U1546 (N_1546,In_185,In_29);
nand U1547 (N_1547,In_663,In_212);
nor U1548 (N_1548,In_42,In_375);
and U1549 (N_1549,In_323,In_377);
nand U1550 (N_1550,In_121,In_937);
and U1551 (N_1551,In_497,In_768);
nor U1552 (N_1552,In_250,In_453);
nor U1553 (N_1553,In_965,In_719);
and U1554 (N_1554,In_780,In_756);
and U1555 (N_1555,In_155,In_413);
or U1556 (N_1556,In_581,In_704);
or U1557 (N_1557,In_364,In_787);
and U1558 (N_1558,In_234,In_973);
nor U1559 (N_1559,In_2,In_977);
and U1560 (N_1560,In_608,In_260);
nor U1561 (N_1561,In_895,In_576);
nor U1562 (N_1562,In_533,In_110);
nor U1563 (N_1563,In_510,In_806);
or U1564 (N_1564,In_529,In_569);
or U1565 (N_1565,In_785,In_994);
and U1566 (N_1566,In_168,In_895);
nor U1567 (N_1567,In_461,In_687);
or U1568 (N_1568,In_43,In_97);
nor U1569 (N_1569,In_318,In_602);
nor U1570 (N_1570,In_11,In_546);
and U1571 (N_1571,In_196,In_730);
and U1572 (N_1572,In_45,In_873);
nand U1573 (N_1573,In_530,In_73);
nor U1574 (N_1574,In_671,In_139);
and U1575 (N_1575,In_609,In_56);
nand U1576 (N_1576,In_30,In_843);
nor U1577 (N_1577,In_536,In_298);
or U1578 (N_1578,In_618,In_656);
or U1579 (N_1579,In_752,In_243);
and U1580 (N_1580,In_455,In_661);
or U1581 (N_1581,In_46,In_347);
and U1582 (N_1582,In_870,In_287);
and U1583 (N_1583,In_568,In_929);
nand U1584 (N_1584,In_931,In_456);
and U1585 (N_1585,In_348,In_479);
nand U1586 (N_1586,In_436,In_540);
and U1587 (N_1587,In_218,In_434);
nor U1588 (N_1588,In_411,In_456);
nand U1589 (N_1589,In_551,In_187);
nand U1590 (N_1590,In_793,In_225);
and U1591 (N_1591,In_132,In_761);
xor U1592 (N_1592,In_28,In_21);
xnor U1593 (N_1593,In_303,In_486);
or U1594 (N_1594,In_710,In_790);
nor U1595 (N_1595,In_424,In_533);
and U1596 (N_1596,In_994,In_837);
and U1597 (N_1597,In_133,In_962);
nand U1598 (N_1598,In_947,In_641);
and U1599 (N_1599,In_591,In_145);
or U1600 (N_1600,In_284,In_326);
and U1601 (N_1601,In_354,In_120);
nand U1602 (N_1602,In_253,In_797);
nor U1603 (N_1603,In_122,In_825);
and U1604 (N_1604,In_255,In_826);
xor U1605 (N_1605,In_541,In_874);
nor U1606 (N_1606,In_525,In_699);
nor U1607 (N_1607,In_848,In_187);
or U1608 (N_1608,In_737,In_164);
nand U1609 (N_1609,In_747,In_612);
and U1610 (N_1610,In_640,In_542);
and U1611 (N_1611,In_222,In_296);
xnor U1612 (N_1612,In_326,In_436);
and U1613 (N_1613,In_163,In_443);
nor U1614 (N_1614,In_115,In_478);
nor U1615 (N_1615,In_370,In_431);
or U1616 (N_1616,In_383,In_411);
nand U1617 (N_1617,In_369,In_360);
or U1618 (N_1618,In_451,In_796);
or U1619 (N_1619,In_116,In_160);
and U1620 (N_1620,In_996,In_339);
nand U1621 (N_1621,In_129,In_447);
nand U1622 (N_1622,In_920,In_420);
xor U1623 (N_1623,In_553,In_970);
nand U1624 (N_1624,In_189,In_483);
and U1625 (N_1625,In_775,In_815);
nand U1626 (N_1626,In_468,In_250);
nand U1627 (N_1627,In_940,In_711);
or U1628 (N_1628,In_679,In_740);
and U1629 (N_1629,In_897,In_690);
nand U1630 (N_1630,In_404,In_539);
or U1631 (N_1631,In_843,In_369);
and U1632 (N_1632,In_276,In_94);
or U1633 (N_1633,In_599,In_406);
or U1634 (N_1634,In_504,In_279);
or U1635 (N_1635,In_833,In_49);
and U1636 (N_1636,In_596,In_175);
nor U1637 (N_1637,In_438,In_860);
nand U1638 (N_1638,In_614,In_498);
or U1639 (N_1639,In_411,In_391);
nor U1640 (N_1640,In_817,In_402);
nand U1641 (N_1641,In_423,In_375);
nand U1642 (N_1642,In_227,In_938);
nand U1643 (N_1643,In_162,In_395);
or U1644 (N_1644,In_182,In_122);
nand U1645 (N_1645,In_539,In_181);
and U1646 (N_1646,In_719,In_813);
nand U1647 (N_1647,In_57,In_792);
nor U1648 (N_1648,In_837,In_186);
and U1649 (N_1649,In_428,In_523);
nor U1650 (N_1650,In_760,In_372);
nand U1651 (N_1651,In_282,In_893);
and U1652 (N_1652,In_425,In_5);
nand U1653 (N_1653,In_126,In_327);
or U1654 (N_1654,In_940,In_694);
xnor U1655 (N_1655,In_327,In_566);
nand U1656 (N_1656,In_963,In_663);
nand U1657 (N_1657,In_345,In_419);
nor U1658 (N_1658,In_388,In_326);
nor U1659 (N_1659,In_878,In_671);
and U1660 (N_1660,In_921,In_640);
or U1661 (N_1661,In_178,In_537);
nand U1662 (N_1662,In_538,In_145);
nor U1663 (N_1663,In_315,In_958);
and U1664 (N_1664,In_564,In_846);
nor U1665 (N_1665,In_651,In_258);
or U1666 (N_1666,In_169,In_516);
and U1667 (N_1667,In_874,In_550);
or U1668 (N_1668,In_574,In_249);
nand U1669 (N_1669,In_590,In_507);
and U1670 (N_1670,In_337,In_107);
nand U1671 (N_1671,In_869,In_590);
nor U1672 (N_1672,In_982,In_981);
nand U1673 (N_1673,In_756,In_532);
nand U1674 (N_1674,In_797,In_980);
nor U1675 (N_1675,In_718,In_703);
and U1676 (N_1676,In_369,In_565);
and U1677 (N_1677,In_578,In_851);
nand U1678 (N_1678,In_928,In_314);
or U1679 (N_1679,In_71,In_107);
nor U1680 (N_1680,In_664,In_728);
nor U1681 (N_1681,In_744,In_401);
nand U1682 (N_1682,In_758,In_928);
and U1683 (N_1683,In_73,In_892);
and U1684 (N_1684,In_176,In_10);
or U1685 (N_1685,In_437,In_861);
and U1686 (N_1686,In_927,In_677);
and U1687 (N_1687,In_543,In_477);
nor U1688 (N_1688,In_504,In_447);
or U1689 (N_1689,In_414,In_57);
nand U1690 (N_1690,In_899,In_444);
and U1691 (N_1691,In_473,In_928);
nand U1692 (N_1692,In_72,In_557);
nand U1693 (N_1693,In_506,In_462);
nand U1694 (N_1694,In_602,In_157);
nand U1695 (N_1695,In_889,In_287);
nand U1696 (N_1696,In_175,In_950);
nand U1697 (N_1697,In_807,In_627);
nand U1698 (N_1698,In_151,In_10);
nand U1699 (N_1699,In_556,In_859);
or U1700 (N_1700,In_271,In_992);
nor U1701 (N_1701,In_10,In_537);
nand U1702 (N_1702,In_17,In_84);
nor U1703 (N_1703,In_779,In_698);
and U1704 (N_1704,In_686,In_775);
and U1705 (N_1705,In_41,In_558);
nor U1706 (N_1706,In_172,In_946);
and U1707 (N_1707,In_893,In_911);
nand U1708 (N_1708,In_993,In_383);
nand U1709 (N_1709,In_346,In_501);
nor U1710 (N_1710,In_178,In_662);
nand U1711 (N_1711,In_893,In_980);
nor U1712 (N_1712,In_572,In_965);
and U1713 (N_1713,In_355,In_155);
and U1714 (N_1714,In_708,In_304);
or U1715 (N_1715,In_813,In_796);
nand U1716 (N_1716,In_972,In_915);
and U1717 (N_1717,In_883,In_140);
or U1718 (N_1718,In_228,In_288);
nor U1719 (N_1719,In_682,In_560);
nor U1720 (N_1720,In_792,In_590);
or U1721 (N_1721,In_348,In_809);
and U1722 (N_1722,In_902,In_241);
nor U1723 (N_1723,In_129,In_546);
nand U1724 (N_1724,In_569,In_311);
and U1725 (N_1725,In_143,In_283);
nand U1726 (N_1726,In_779,In_441);
and U1727 (N_1727,In_244,In_586);
nor U1728 (N_1728,In_138,In_533);
nor U1729 (N_1729,In_534,In_875);
nor U1730 (N_1730,In_66,In_183);
nor U1731 (N_1731,In_118,In_341);
nor U1732 (N_1732,In_36,In_685);
nand U1733 (N_1733,In_298,In_907);
or U1734 (N_1734,In_190,In_748);
nand U1735 (N_1735,In_46,In_514);
and U1736 (N_1736,In_22,In_401);
or U1737 (N_1737,In_273,In_994);
and U1738 (N_1738,In_929,In_221);
nand U1739 (N_1739,In_317,In_760);
nor U1740 (N_1740,In_433,In_738);
or U1741 (N_1741,In_592,In_483);
nand U1742 (N_1742,In_403,In_355);
nand U1743 (N_1743,In_727,In_988);
nand U1744 (N_1744,In_824,In_839);
nor U1745 (N_1745,In_512,In_922);
or U1746 (N_1746,In_142,In_56);
and U1747 (N_1747,In_204,In_734);
xnor U1748 (N_1748,In_33,In_942);
nor U1749 (N_1749,In_990,In_611);
nand U1750 (N_1750,In_922,In_90);
or U1751 (N_1751,In_553,In_642);
nor U1752 (N_1752,In_348,In_746);
nor U1753 (N_1753,In_672,In_420);
nor U1754 (N_1754,In_353,In_814);
nor U1755 (N_1755,In_215,In_830);
nor U1756 (N_1756,In_436,In_771);
nand U1757 (N_1757,In_501,In_224);
nand U1758 (N_1758,In_123,In_665);
or U1759 (N_1759,In_581,In_61);
nand U1760 (N_1760,In_753,In_464);
and U1761 (N_1761,In_132,In_209);
or U1762 (N_1762,In_989,In_240);
xor U1763 (N_1763,In_890,In_727);
xor U1764 (N_1764,In_775,In_207);
nand U1765 (N_1765,In_856,In_309);
or U1766 (N_1766,In_574,In_165);
or U1767 (N_1767,In_403,In_112);
nor U1768 (N_1768,In_116,In_228);
or U1769 (N_1769,In_736,In_989);
or U1770 (N_1770,In_453,In_326);
or U1771 (N_1771,In_531,In_480);
and U1772 (N_1772,In_490,In_142);
and U1773 (N_1773,In_339,In_307);
or U1774 (N_1774,In_349,In_256);
and U1775 (N_1775,In_43,In_999);
and U1776 (N_1776,In_967,In_576);
nor U1777 (N_1777,In_13,In_574);
nand U1778 (N_1778,In_80,In_376);
nand U1779 (N_1779,In_65,In_28);
and U1780 (N_1780,In_55,In_921);
or U1781 (N_1781,In_824,In_676);
or U1782 (N_1782,In_425,In_818);
nand U1783 (N_1783,In_92,In_33);
and U1784 (N_1784,In_660,In_947);
and U1785 (N_1785,In_397,In_784);
nor U1786 (N_1786,In_611,In_181);
nor U1787 (N_1787,In_300,In_522);
nor U1788 (N_1788,In_813,In_231);
nor U1789 (N_1789,In_652,In_987);
nor U1790 (N_1790,In_893,In_918);
nor U1791 (N_1791,In_944,In_140);
nor U1792 (N_1792,In_924,In_189);
or U1793 (N_1793,In_919,In_761);
or U1794 (N_1794,In_461,In_734);
or U1795 (N_1795,In_511,In_953);
nand U1796 (N_1796,In_921,In_104);
nor U1797 (N_1797,In_127,In_620);
nor U1798 (N_1798,In_673,In_811);
or U1799 (N_1799,In_828,In_611);
nand U1800 (N_1800,In_15,In_686);
nand U1801 (N_1801,In_350,In_305);
or U1802 (N_1802,In_921,In_58);
nor U1803 (N_1803,In_668,In_660);
nor U1804 (N_1804,In_452,In_43);
nand U1805 (N_1805,In_439,In_122);
or U1806 (N_1806,In_313,In_535);
and U1807 (N_1807,In_410,In_240);
nand U1808 (N_1808,In_111,In_96);
or U1809 (N_1809,In_767,In_713);
or U1810 (N_1810,In_389,In_159);
nor U1811 (N_1811,In_521,In_936);
and U1812 (N_1812,In_882,In_284);
and U1813 (N_1813,In_743,In_362);
nor U1814 (N_1814,In_330,In_0);
nor U1815 (N_1815,In_483,In_801);
and U1816 (N_1816,In_735,In_909);
nand U1817 (N_1817,In_557,In_40);
and U1818 (N_1818,In_989,In_271);
nor U1819 (N_1819,In_549,In_982);
nand U1820 (N_1820,In_607,In_114);
nand U1821 (N_1821,In_892,In_729);
or U1822 (N_1822,In_624,In_674);
nor U1823 (N_1823,In_344,In_285);
nand U1824 (N_1824,In_740,In_993);
nand U1825 (N_1825,In_167,In_586);
nor U1826 (N_1826,In_764,In_319);
nand U1827 (N_1827,In_960,In_735);
or U1828 (N_1828,In_586,In_200);
nor U1829 (N_1829,In_123,In_503);
or U1830 (N_1830,In_535,In_253);
nand U1831 (N_1831,In_919,In_91);
nand U1832 (N_1832,In_301,In_109);
xor U1833 (N_1833,In_132,In_679);
or U1834 (N_1834,In_242,In_210);
or U1835 (N_1835,In_789,In_863);
nand U1836 (N_1836,In_501,In_457);
nor U1837 (N_1837,In_264,In_969);
and U1838 (N_1838,In_635,In_230);
and U1839 (N_1839,In_377,In_792);
and U1840 (N_1840,In_36,In_702);
or U1841 (N_1841,In_649,In_734);
and U1842 (N_1842,In_500,In_356);
nand U1843 (N_1843,In_209,In_441);
nor U1844 (N_1844,In_280,In_107);
nor U1845 (N_1845,In_864,In_676);
nand U1846 (N_1846,In_507,In_214);
and U1847 (N_1847,In_256,In_947);
and U1848 (N_1848,In_386,In_207);
or U1849 (N_1849,In_605,In_799);
and U1850 (N_1850,In_248,In_916);
nand U1851 (N_1851,In_434,In_161);
and U1852 (N_1852,In_756,In_486);
nand U1853 (N_1853,In_252,In_433);
and U1854 (N_1854,In_262,In_29);
nand U1855 (N_1855,In_368,In_263);
and U1856 (N_1856,In_668,In_54);
nand U1857 (N_1857,In_138,In_381);
nand U1858 (N_1858,In_900,In_187);
and U1859 (N_1859,In_260,In_620);
nand U1860 (N_1860,In_338,In_412);
and U1861 (N_1861,In_405,In_96);
or U1862 (N_1862,In_314,In_5);
nand U1863 (N_1863,In_165,In_199);
and U1864 (N_1864,In_351,In_362);
and U1865 (N_1865,In_119,In_713);
nand U1866 (N_1866,In_436,In_468);
nand U1867 (N_1867,In_19,In_188);
nand U1868 (N_1868,In_42,In_978);
or U1869 (N_1869,In_873,In_59);
and U1870 (N_1870,In_789,In_885);
nor U1871 (N_1871,In_517,In_480);
nor U1872 (N_1872,In_651,In_907);
or U1873 (N_1873,In_316,In_199);
and U1874 (N_1874,In_712,In_240);
nor U1875 (N_1875,In_948,In_423);
and U1876 (N_1876,In_492,In_220);
nor U1877 (N_1877,In_205,In_777);
nor U1878 (N_1878,In_35,In_139);
nor U1879 (N_1879,In_971,In_114);
nand U1880 (N_1880,In_870,In_549);
or U1881 (N_1881,In_923,In_863);
nand U1882 (N_1882,In_830,In_781);
and U1883 (N_1883,In_652,In_98);
and U1884 (N_1884,In_827,In_943);
nor U1885 (N_1885,In_315,In_231);
nand U1886 (N_1886,In_77,In_236);
or U1887 (N_1887,In_26,In_822);
and U1888 (N_1888,In_530,In_558);
or U1889 (N_1889,In_317,In_152);
nor U1890 (N_1890,In_202,In_549);
nor U1891 (N_1891,In_143,In_938);
and U1892 (N_1892,In_584,In_131);
nand U1893 (N_1893,In_575,In_740);
and U1894 (N_1894,In_407,In_916);
or U1895 (N_1895,In_782,In_980);
or U1896 (N_1896,In_974,In_179);
or U1897 (N_1897,In_41,In_486);
nor U1898 (N_1898,In_133,In_457);
or U1899 (N_1899,In_45,In_615);
and U1900 (N_1900,In_5,In_432);
nor U1901 (N_1901,In_535,In_608);
and U1902 (N_1902,In_95,In_237);
nor U1903 (N_1903,In_506,In_935);
nand U1904 (N_1904,In_375,In_495);
nor U1905 (N_1905,In_892,In_512);
and U1906 (N_1906,In_953,In_305);
nor U1907 (N_1907,In_563,In_114);
nor U1908 (N_1908,In_882,In_697);
nor U1909 (N_1909,In_382,In_244);
and U1910 (N_1910,In_686,In_369);
or U1911 (N_1911,In_702,In_181);
or U1912 (N_1912,In_451,In_518);
nand U1913 (N_1913,In_102,In_631);
nand U1914 (N_1914,In_503,In_291);
nor U1915 (N_1915,In_481,In_970);
or U1916 (N_1916,In_598,In_982);
nand U1917 (N_1917,In_974,In_349);
and U1918 (N_1918,In_9,In_45);
nand U1919 (N_1919,In_139,In_791);
or U1920 (N_1920,In_181,In_233);
and U1921 (N_1921,In_212,In_821);
and U1922 (N_1922,In_565,In_584);
nand U1923 (N_1923,In_265,In_316);
and U1924 (N_1924,In_617,In_864);
and U1925 (N_1925,In_594,In_9);
or U1926 (N_1926,In_864,In_946);
and U1927 (N_1927,In_281,In_679);
nand U1928 (N_1928,In_458,In_528);
and U1929 (N_1929,In_664,In_470);
nand U1930 (N_1930,In_602,In_978);
nand U1931 (N_1931,In_843,In_973);
nand U1932 (N_1932,In_270,In_485);
and U1933 (N_1933,In_512,In_902);
or U1934 (N_1934,In_561,In_474);
nand U1935 (N_1935,In_828,In_434);
and U1936 (N_1936,In_891,In_49);
nand U1937 (N_1937,In_460,In_716);
nor U1938 (N_1938,In_319,In_664);
xor U1939 (N_1939,In_851,In_575);
or U1940 (N_1940,In_664,In_613);
or U1941 (N_1941,In_938,In_3);
nand U1942 (N_1942,In_151,In_770);
and U1943 (N_1943,In_452,In_631);
or U1944 (N_1944,In_501,In_343);
nor U1945 (N_1945,In_980,In_946);
and U1946 (N_1946,In_796,In_802);
and U1947 (N_1947,In_607,In_213);
xor U1948 (N_1948,In_176,In_64);
and U1949 (N_1949,In_495,In_224);
nand U1950 (N_1950,In_594,In_172);
and U1951 (N_1951,In_705,In_243);
or U1952 (N_1952,In_354,In_351);
nand U1953 (N_1953,In_324,In_127);
nor U1954 (N_1954,In_540,In_421);
or U1955 (N_1955,In_466,In_127);
and U1956 (N_1956,In_870,In_501);
nor U1957 (N_1957,In_18,In_41);
or U1958 (N_1958,In_806,In_329);
or U1959 (N_1959,In_306,In_632);
and U1960 (N_1960,In_280,In_153);
nor U1961 (N_1961,In_222,In_182);
and U1962 (N_1962,In_557,In_906);
xnor U1963 (N_1963,In_271,In_293);
nor U1964 (N_1964,In_244,In_898);
nand U1965 (N_1965,In_579,In_424);
nand U1966 (N_1966,In_318,In_161);
nand U1967 (N_1967,In_903,In_279);
and U1968 (N_1968,In_608,In_197);
or U1969 (N_1969,In_616,In_262);
nand U1970 (N_1970,In_321,In_694);
or U1971 (N_1971,In_274,In_827);
and U1972 (N_1972,In_654,In_970);
nand U1973 (N_1973,In_698,In_985);
nand U1974 (N_1974,In_53,In_39);
nand U1975 (N_1975,In_863,In_919);
nand U1976 (N_1976,In_298,In_280);
nor U1977 (N_1977,In_621,In_956);
nor U1978 (N_1978,In_878,In_12);
xor U1979 (N_1979,In_960,In_809);
nor U1980 (N_1980,In_298,In_312);
nor U1981 (N_1981,In_550,In_404);
or U1982 (N_1982,In_255,In_344);
nand U1983 (N_1983,In_173,In_16);
nor U1984 (N_1984,In_251,In_192);
nor U1985 (N_1985,In_297,In_929);
and U1986 (N_1986,In_161,In_406);
and U1987 (N_1987,In_606,In_966);
nand U1988 (N_1988,In_822,In_928);
nand U1989 (N_1989,In_199,In_980);
nand U1990 (N_1990,In_544,In_568);
or U1991 (N_1991,In_40,In_34);
or U1992 (N_1992,In_495,In_936);
nor U1993 (N_1993,In_731,In_690);
and U1994 (N_1994,In_813,In_209);
and U1995 (N_1995,In_825,In_623);
nand U1996 (N_1996,In_558,In_14);
nor U1997 (N_1997,In_808,In_259);
nand U1998 (N_1998,In_800,In_316);
and U1999 (N_1999,In_572,In_579);
nor U2000 (N_2000,N_54,N_1418);
nand U2001 (N_2001,N_270,N_210);
nor U2002 (N_2002,N_1073,N_1715);
nor U2003 (N_2003,N_1026,N_985);
nand U2004 (N_2004,N_1947,N_900);
nand U2005 (N_2005,N_330,N_1732);
or U2006 (N_2006,N_676,N_1712);
nand U2007 (N_2007,N_1781,N_995);
nor U2008 (N_2008,N_1237,N_1893);
or U2009 (N_2009,N_471,N_1508);
or U2010 (N_2010,N_1555,N_384);
nor U2011 (N_2011,N_527,N_784);
and U2012 (N_2012,N_969,N_1081);
and U2013 (N_2013,N_66,N_1637);
or U2014 (N_2014,N_709,N_670);
xnor U2015 (N_2015,N_491,N_1869);
nand U2016 (N_2016,N_566,N_851);
nor U2017 (N_2017,N_1266,N_961);
nor U2018 (N_2018,N_142,N_1965);
and U2019 (N_2019,N_1413,N_612);
nor U2020 (N_2020,N_1742,N_1853);
nand U2021 (N_2021,N_1557,N_117);
or U2022 (N_2022,N_138,N_1000);
xnor U2023 (N_2023,N_1954,N_1888);
and U2024 (N_2024,N_1638,N_1569);
nor U2025 (N_2025,N_737,N_810);
nand U2026 (N_2026,N_899,N_1390);
nor U2027 (N_2027,N_72,N_257);
nor U2028 (N_2028,N_608,N_1835);
nor U2029 (N_2029,N_1323,N_852);
nand U2030 (N_2030,N_31,N_1622);
nand U2031 (N_2031,N_1783,N_1377);
nor U2032 (N_2032,N_118,N_1868);
nor U2033 (N_2033,N_1375,N_1141);
or U2034 (N_2034,N_76,N_521);
nand U2035 (N_2035,N_254,N_228);
nand U2036 (N_2036,N_227,N_1654);
nand U2037 (N_2037,N_1604,N_1850);
nand U2038 (N_2038,N_753,N_157);
and U2039 (N_2039,N_372,N_1215);
and U2040 (N_2040,N_181,N_1762);
and U2041 (N_2041,N_989,N_263);
and U2042 (N_2042,N_686,N_1428);
nor U2043 (N_2043,N_1169,N_1095);
and U2044 (N_2044,N_1928,N_1220);
and U2045 (N_2045,N_124,N_1972);
nand U2046 (N_2046,N_291,N_1738);
or U2047 (N_2047,N_1499,N_399);
and U2048 (N_2048,N_708,N_1013);
and U2049 (N_2049,N_417,N_943);
or U2050 (N_2050,N_1686,N_189);
and U2051 (N_2051,N_29,N_159);
or U2052 (N_2052,N_238,N_1149);
nor U2053 (N_2053,N_744,N_963);
and U2054 (N_2054,N_1550,N_204);
nand U2055 (N_2055,N_277,N_693);
nand U2056 (N_2056,N_1474,N_508);
or U2057 (N_2057,N_947,N_146);
and U2058 (N_2058,N_822,N_1626);
xor U2059 (N_2059,N_519,N_973);
and U2060 (N_2060,N_1245,N_1528);
or U2061 (N_2061,N_554,N_721);
or U2062 (N_2062,N_1203,N_997);
nor U2063 (N_2063,N_1834,N_1238);
and U2064 (N_2064,N_671,N_1416);
xnor U2065 (N_2065,N_1564,N_928);
and U2066 (N_2066,N_1651,N_1523);
and U2067 (N_2067,N_588,N_774);
nor U2068 (N_2068,N_958,N_1748);
nand U2069 (N_2069,N_833,N_1405);
nor U2070 (N_2070,N_1709,N_550);
nor U2071 (N_2071,N_324,N_1098);
nor U2072 (N_2072,N_1484,N_1806);
and U2073 (N_2073,N_1792,N_451);
nand U2074 (N_2074,N_874,N_1349);
nand U2075 (N_2075,N_617,N_1194);
nand U2076 (N_2076,N_1312,N_1317);
and U2077 (N_2077,N_1678,N_1258);
and U2078 (N_2078,N_295,N_1348);
nand U2079 (N_2079,N_1771,N_338);
and U2080 (N_2080,N_678,N_871);
nor U2081 (N_2081,N_164,N_107);
or U2082 (N_2082,N_1219,N_727);
or U2083 (N_2083,N_1468,N_109);
or U2084 (N_2084,N_1874,N_1330);
or U2085 (N_2085,N_877,N_1608);
nand U2086 (N_2086,N_1520,N_901);
and U2087 (N_2087,N_1764,N_1155);
nor U2088 (N_2088,N_1267,N_1045);
and U2089 (N_2089,N_1364,N_1964);
xnor U2090 (N_2090,N_667,N_925);
nand U2091 (N_2091,N_252,N_461);
nand U2092 (N_2092,N_1036,N_5);
nor U2093 (N_2093,N_1690,N_377);
nor U2094 (N_2094,N_309,N_917);
or U2095 (N_2095,N_91,N_694);
nand U2096 (N_2096,N_1674,N_1136);
nor U2097 (N_2097,N_652,N_647);
and U2098 (N_2098,N_485,N_19);
nor U2099 (N_2099,N_1286,N_1586);
nor U2100 (N_2100,N_1675,N_1503);
or U2101 (N_2101,N_55,N_597);
and U2102 (N_2102,N_1163,N_1516);
nor U2103 (N_2103,N_746,N_1042);
nor U2104 (N_2104,N_1204,N_1437);
nand U2105 (N_2105,N_1251,N_1280);
and U2106 (N_2106,N_77,N_1560);
or U2107 (N_2107,N_1525,N_1090);
nand U2108 (N_2108,N_459,N_442);
and U2109 (N_2109,N_283,N_440);
and U2110 (N_2110,N_466,N_1059);
or U2111 (N_2111,N_885,N_365);
nor U2112 (N_2112,N_1359,N_75);
and U2113 (N_2113,N_980,N_960);
nand U2114 (N_2114,N_241,N_386);
and U2115 (N_2115,N_366,N_396);
or U2116 (N_2116,N_1154,N_1668);
nand U2117 (N_2117,N_1322,N_1049);
nand U2118 (N_2118,N_12,N_1249);
and U2119 (N_2119,N_1363,N_427);
and U2120 (N_2120,N_977,N_489);
nand U2121 (N_2121,N_1183,N_1378);
and U2122 (N_2122,N_119,N_533);
and U2123 (N_2123,N_574,N_1534);
and U2124 (N_2124,N_994,N_1092);
nor U2125 (N_2125,N_1898,N_1787);
nor U2126 (N_2126,N_1729,N_540);
nand U2127 (N_2127,N_331,N_1053);
nor U2128 (N_2128,N_363,N_93);
nand U2129 (N_2129,N_1327,N_1289);
and U2130 (N_2130,N_1447,N_239);
and U2131 (N_2131,N_1189,N_1467);
nand U2132 (N_2132,N_1663,N_1386);
and U2133 (N_2133,N_475,N_1234);
and U2134 (N_2134,N_1684,N_1096);
nand U2135 (N_2135,N_498,N_756);
or U2136 (N_2136,N_1782,N_1362);
nand U2137 (N_2137,N_457,N_1909);
xnor U2138 (N_2138,N_1271,N_1126);
and U2139 (N_2139,N_1372,N_1291);
and U2140 (N_2140,N_256,N_329);
nand U2141 (N_2141,N_1607,N_1841);
and U2142 (N_2142,N_594,N_615);
and U2143 (N_2143,N_73,N_1681);
nor U2144 (N_2144,N_1262,N_101);
xor U2145 (N_2145,N_1776,N_783);
and U2146 (N_2146,N_481,N_25);
nor U2147 (N_2147,N_750,N_1978);
or U2148 (N_2148,N_1578,N_1821);
and U2149 (N_2149,N_1700,N_545);
or U2150 (N_2150,N_1677,N_401);
nand U2151 (N_2151,N_41,N_201);
nand U2152 (N_2152,N_1120,N_1211);
or U2153 (N_2153,N_1736,N_362);
nand U2154 (N_2154,N_409,N_1643);
and U2155 (N_2155,N_1477,N_406);
nand U2156 (N_2156,N_1545,N_1759);
and U2157 (N_2157,N_1639,N_1165);
or U2158 (N_2158,N_356,N_1240);
nor U2159 (N_2159,N_416,N_130);
and U2160 (N_2160,N_1340,N_831);
and U2161 (N_2161,N_1839,N_939);
or U2162 (N_2162,N_133,N_870);
or U2163 (N_2163,N_891,N_1043);
and U2164 (N_2164,N_1366,N_182);
xor U2165 (N_2165,N_905,N_982);
nand U2166 (N_2166,N_1209,N_813);
nor U2167 (N_2167,N_1187,N_44);
or U2168 (N_2168,N_592,N_1975);
or U2169 (N_2169,N_663,N_1987);
nand U2170 (N_2170,N_328,N_1048);
or U2171 (N_2171,N_711,N_206);
nor U2172 (N_2172,N_1827,N_805);
nor U2173 (N_2173,N_613,N_1110);
and U2174 (N_2174,N_1921,N_873);
or U2175 (N_2175,N_1253,N_1966);
or U2176 (N_2176,N_589,N_896);
and U2177 (N_2177,N_1318,N_1730);
and U2178 (N_2178,N_1007,N_830);
nand U2179 (N_2179,N_776,N_669);
nor U2180 (N_2180,N_100,N_762);
and U2181 (N_2181,N_520,N_1296);
nand U2182 (N_2182,N_314,N_1683);
and U2183 (N_2183,N_734,N_21);
nor U2184 (N_2184,N_1460,N_1275);
or U2185 (N_2185,N_1172,N_1283);
nand U2186 (N_2186,N_430,N_707);
xor U2187 (N_2187,N_1876,N_1763);
or U2188 (N_2188,N_675,N_846);
nor U2189 (N_2189,N_549,N_469);
and U2190 (N_2190,N_1509,N_1808);
nand U2191 (N_2191,N_1846,N_70);
nand U2192 (N_2192,N_1800,N_1004);
nand U2193 (N_2193,N_1645,N_1252);
or U2194 (N_2194,N_562,N_1383);
or U2195 (N_2195,N_1804,N_1913);
xnor U2196 (N_2196,N_1582,N_1515);
and U2197 (N_2197,N_169,N_957);
nor U2198 (N_2198,N_438,N_1469);
and U2199 (N_2199,N_966,N_1157);
and U2200 (N_2200,N_651,N_983);
nor U2201 (N_2201,N_258,N_487);
nor U2202 (N_2202,N_1463,N_1670);
and U2203 (N_2203,N_546,N_1100);
nor U2204 (N_2204,N_301,N_567);
and U2205 (N_2205,N_649,N_1990);
nor U2206 (N_2206,N_832,N_1522);
nand U2207 (N_2207,N_111,N_271);
nor U2208 (N_2208,N_1478,N_1935);
nor U2209 (N_2209,N_420,N_1412);
nor U2210 (N_2210,N_856,N_251);
nor U2211 (N_2211,N_701,N_796);
nor U2212 (N_2212,N_765,N_246);
nand U2213 (N_2213,N_682,N_785);
and U2214 (N_2214,N_139,N_209);
and U2215 (N_2215,N_339,N_1139);
and U2216 (N_2216,N_1572,N_674);
or U2217 (N_2217,N_1077,N_655);
or U2218 (N_2218,N_658,N_447);
and U2219 (N_2219,N_1506,N_1803);
nand U2220 (N_2220,N_351,N_374);
nand U2221 (N_2221,N_979,N_360);
nand U2222 (N_2222,N_1823,N_732);
nand U2223 (N_2223,N_1033,N_300);
nand U2224 (N_2224,N_1153,N_883);
nand U2225 (N_2225,N_818,N_484);
and U2226 (N_2226,N_382,N_627);
nor U2227 (N_2227,N_1281,N_1968);
nor U2228 (N_2228,N_1174,N_1476);
and U2229 (N_2229,N_849,N_869);
and U2230 (N_2230,N_920,N_1959);
nand U2231 (N_2231,N_794,N_897);
nor U2232 (N_2232,N_630,N_65);
or U2233 (N_2233,N_286,N_316);
nand U2234 (N_2234,N_628,N_1754);
nor U2235 (N_2235,N_103,N_691);
and U2236 (N_2236,N_911,N_660);
or U2237 (N_2237,N_1575,N_174);
nor U2238 (N_2238,N_1339,N_448);
and U2239 (N_2239,N_778,N_1728);
nor U2240 (N_2240,N_940,N_786);
or U2241 (N_2241,N_751,N_1415);
nor U2242 (N_2242,N_1230,N_170);
nor U2243 (N_2243,N_1940,N_1186);
nor U2244 (N_2244,N_1926,N_1162);
and U2245 (N_2245,N_1963,N_1887);
nor U2246 (N_2246,N_1309,N_334);
xnor U2247 (N_2247,N_1649,N_58);
or U2248 (N_2248,N_1722,N_370);
or U2249 (N_2249,N_1111,N_1884);
and U2250 (N_2250,N_1093,N_1999);
nor U2251 (N_2251,N_1831,N_1099);
and U2252 (N_2252,N_1828,N_1878);
and U2253 (N_2253,N_1544,N_993);
and U2254 (N_2254,N_801,N_1551);
nor U2255 (N_2255,N_198,N_565);
and U2256 (N_2256,N_1871,N_1830);
nand U2257 (N_2257,N_90,N_1672);
nand U2258 (N_2258,N_1798,N_60);
nand U2259 (N_2259,N_444,N_972);
and U2260 (N_2260,N_1190,N_571);
nand U2261 (N_2261,N_1952,N_1369);
nor U2262 (N_2262,N_320,N_261);
nand U2263 (N_2263,N_1864,N_1440);
nor U2264 (N_2264,N_494,N_1837);
or U2265 (N_2265,N_1570,N_560);
and U2266 (N_2266,N_772,N_1064);
and U2267 (N_2267,N_656,N_1385);
nand U2268 (N_2268,N_698,N_1373);
nand U2269 (N_2269,N_575,N_975);
or U2270 (N_2270,N_1041,N_1051);
nand U2271 (N_2271,N_1886,N_74);
nand U2272 (N_2272,N_1411,N_821);
and U2273 (N_2273,N_1094,N_464);
and U2274 (N_2274,N_140,N_352);
nor U2275 (N_2275,N_177,N_614);
nor U2276 (N_2276,N_1780,N_1001);
or U2277 (N_2277,N_1350,N_1900);
and U2278 (N_2278,N_1005,N_81);
and U2279 (N_2279,N_1795,N_1480);
nand U2280 (N_2280,N_1290,N_1845);
or U2281 (N_2281,N_1388,N_910);
and U2282 (N_2282,N_563,N_872);
nand U2283 (N_2283,N_231,N_153);
and U2284 (N_2284,N_265,N_604);
nand U2285 (N_2285,N_322,N_1333);
nor U2286 (N_2286,N_1374,N_150);
or U2287 (N_2287,N_886,N_454);
nor U2288 (N_2288,N_505,N_1140);
or U2289 (N_2289,N_1593,N_172);
and U2290 (N_2290,N_529,N_455);
or U2291 (N_2291,N_1740,N_512);
or U2292 (N_2292,N_373,N_690);
nand U2293 (N_2293,N_912,N_1218);
xor U2294 (N_2294,N_1679,N_260);
nor U2295 (N_2295,N_213,N_586);
nor U2296 (N_2296,N_197,N_358);
nor U2297 (N_2297,N_141,N_535);
nand U2298 (N_2298,N_1427,N_720);
and U2299 (N_2299,N_1791,N_1533);
or U2300 (N_2300,N_1482,N_1257);
nand U2301 (N_2301,N_1807,N_1458);
nand U2302 (N_2302,N_1441,N_95);
nor U2303 (N_2303,N_407,N_446);
nand U2304 (N_2304,N_954,N_1671);
and U2305 (N_2305,N_1595,N_1518);
and U2306 (N_2306,N_930,N_1453);
nand U2307 (N_2307,N_1116,N_1076);
and U2308 (N_2308,N_421,N_525);
nand U2309 (N_2309,N_1535,N_841);
and U2310 (N_2310,N_923,N_828);
nor U2311 (N_2311,N_1083,N_1725);
or U2312 (N_2312,N_1983,N_978);
nor U2313 (N_2313,N_1897,N_1711);
and U2314 (N_2314,N_26,N_1387);
nor U2315 (N_2315,N_287,N_1347);
and U2316 (N_2316,N_1775,N_176);
or U2317 (N_2317,N_837,N_1487);
and U2318 (N_2318,N_1571,N_607);
or U2319 (N_2319,N_1250,N_230);
or U2320 (N_2320,N_3,N_340);
nand U2321 (N_2321,N_424,N_203);
nand U2322 (N_2322,N_815,N_1699);
nand U2323 (N_2323,N_276,N_1);
or U2324 (N_2324,N_1682,N_1851);
nand U2325 (N_2325,N_840,N_51);
nor U2326 (N_2326,N_1490,N_1532);
and U2327 (N_2327,N_183,N_1423);
and U2328 (N_2328,N_754,N_845);
nor U2329 (N_2329,N_405,N_517);
nor U2330 (N_2330,N_761,N_1634);
nand U2331 (N_2331,N_63,N_1495);
nand U2332 (N_2332,N_740,N_1695);
and U2333 (N_2333,N_890,N_1720);
and U2334 (N_2334,N_452,N_1816);
nor U2335 (N_2335,N_477,N_272);
nor U2336 (N_2336,N_53,N_561);
and U2337 (N_2337,N_1734,N_1242);
nand U2338 (N_2338,N_282,N_1135);
nand U2339 (N_2339,N_1256,N_1142);
and U2340 (N_2340,N_35,N_278);
nor U2341 (N_2341,N_1820,N_1777);
nand U2342 (N_2342,N_1168,N_1927);
and U2343 (N_2343,N_934,N_1319);
nor U2344 (N_2344,N_1310,N_804);
and U2345 (N_2345,N_1946,N_486);
or U2346 (N_2346,N_245,N_1201);
or U2347 (N_2347,N_555,N_1881);
nor U2348 (N_2348,N_1301,N_16);
or U2349 (N_2349,N_1217,N_1822);
nor U2350 (N_2350,N_564,N_522);
nand U2351 (N_2351,N_999,N_236);
and U2352 (N_2352,N_611,N_341);
nand U2353 (N_2353,N_312,N_689);
nand U2354 (N_2354,N_1594,N_394);
and U2355 (N_2355,N_110,N_1615);
and U2356 (N_2356,N_62,N_1994);
nand U2357 (N_2357,N_1693,N_1114);
or U2358 (N_2358,N_166,N_88);
or U2359 (N_2359,N_391,N_294);
and U2360 (N_2360,N_1833,N_1658);
nor U2361 (N_2361,N_1439,N_456);
or U2362 (N_2362,N_749,N_492);
nor U2363 (N_2363,N_470,N_1433);
nor U2364 (N_2364,N_1656,N_1879);
xor U2365 (N_2365,N_1475,N_1743);
nand U2366 (N_2366,N_290,N_593);
nand U2367 (N_2367,N_1911,N_1143);
nand U2368 (N_2368,N_114,N_1344);
or U2369 (N_2369,N_304,N_1832);
and U2370 (N_2370,N_1062,N_20);
and U2371 (N_2371,N_449,N_1829);
or U2372 (N_2372,N_847,N_1751);
and U2373 (N_2373,N_413,N_854);
nand U2374 (N_2374,N_1951,N_1971);
nand U2375 (N_2375,N_1993,N_573);
nor U2376 (N_2376,N_1737,N_666);
nand U2377 (N_2377,N_1337,N_1118);
nand U2378 (N_2378,N_1063,N_237);
nand U2379 (N_2379,N_938,N_1496);
or U2380 (N_2380,N_1089,N_702);
nand U2381 (N_2381,N_1510,N_1160);
nand U2382 (N_2382,N_359,N_1773);
or U2383 (N_2383,N_1769,N_878);
or U2384 (N_2384,N_1538,N_264);
and U2385 (N_2385,N_1723,N_87);
nor U2386 (N_2386,N_1727,N_1040);
or U2387 (N_2387,N_82,N_207);
and U2388 (N_2388,N_161,N_1321);
nor U2389 (N_2389,N_713,N_1922);
nor U2390 (N_2390,N_1580,N_1450);
or U2391 (N_2391,N_926,N_1577);
and U2392 (N_2392,N_1664,N_515);
nand U2393 (N_2393,N_1397,N_375);
nand U2394 (N_2394,N_249,N_1070);
or U2395 (N_2395,N_1548,N_1357);
or U2396 (N_2396,N_715,N_184);
and U2397 (N_2397,N_18,N_538);
and U2398 (N_2398,N_518,N_802);
nor U2399 (N_2399,N_970,N_346);
or U2400 (N_2400,N_557,N_1314);
and U2401 (N_2401,N_1273,N_1311);
nor U2402 (N_2402,N_1793,N_1524);
and U2403 (N_2403,N_321,N_1843);
nand U2404 (N_2404,N_1650,N_1497);
or U2405 (N_2405,N_281,N_867);
nand U2406 (N_2406,N_23,N_1904);
and U2407 (N_2407,N_462,N_817);
and U2408 (N_2408,N_606,N_1810);
nand U2409 (N_2409,N_1818,N_1356);
nand U2410 (N_2410,N_1653,N_149);
or U2411 (N_2411,N_218,N_1912);
and U2412 (N_2412,N_1284,N_136);
nor U2413 (N_2413,N_1840,N_1576);
nand U2414 (N_2414,N_1891,N_367);
and U2415 (N_2415,N_1179,N_868);
nor U2416 (N_2416,N_1766,N_1502);
or U2417 (N_2417,N_534,N_1752);
or U2418 (N_2418,N_1003,N_583);
and U2419 (N_2419,N_1091,N_1421);
or U2420 (N_2420,N_225,N_1161);
nor U2421 (N_2421,N_148,N_1589);
and U2422 (N_2422,N_992,N_1844);
nand U2423 (N_2423,N_1047,N_1080);
or U2424 (N_2424,N_638,N_326);
nand U2425 (N_2425,N_1687,N_1995);
and U2426 (N_2426,N_724,N_156);
nand U2427 (N_2427,N_0,N_1859);
and U2428 (N_2428,N_909,N_116);
nand U2429 (N_2429,N_57,N_1029);
nand U2430 (N_2430,N_104,N_490);
nor U2431 (N_2431,N_1491,N_1949);
nand U2432 (N_2432,N_1652,N_1768);
and U2433 (N_2433,N_1863,N_1899);
nor U2434 (N_2434,N_1075,N_706);
nor U2435 (N_2435,N_123,N_1233);
nor U2436 (N_2436,N_755,N_855);
nand U2437 (N_2437,N_547,N_1379);
and U2438 (N_2438,N_1527,N_1566);
nand U2439 (N_2439,N_493,N_1113);
nor U2440 (N_2440,N_1236,N_1613);
nor U2441 (N_2441,N_1420,N_1431);
nor U2442 (N_2442,N_1903,N_1747);
and U2443 (N_2443,N_1156,N_1500);
nand U2444 (N_2444,N_1996,N_1819);
or U2445 (N_2445,N_552,N_820);
nor U2446 (N_2446,N_650,N_719);
nor U2447 (N_2447,N_1028,N_279);
and U2448 (N_2448,N_1498,N_812);
and U2449 (N_2449,N_319,N_1929);
nand U2450 (N_2450,N_1010,N_1192);
and U2451 (N_2451,N_298,N_537);
and U2452 (N_2452,N_1483,N_1609);
or U2453 (N_2453,N_307,N_662);
nand U2454 (N_2454,N_325,N_79);
nand U2455 (N_2455,N_819,N_1210);
nor U2456 (N_2456,N_1907,N_1459);
nor U2457 (N_2457,N_1540,N_1244);
or U2458 (N_2458,N_1241,N_696);
nor U2459 (N_2459,N_1817,N_7);
nor U2460 (N_2460,N_881,N_1958);
nand U2461 (N_2461,N_46,N_1661);
or U2462 (N_2462,N_600,N_964);
nand U2463 (N_2463,N_480,N_345);
nor U2464 (N_2464,N_1274,N_191);
and U2465 (N_2465,N_904,N_1746);
nor U2466 (N_2466,N_1719,N_9);
and U2467 (N_2467,N_528,N_779);
and U2468 (N_2468,N_543,N_1293);
nor U2469 (N_2469,N_1813,N_1568);
or U2470 (N_2470,N_1127,N_797);
and U2471 (N_2471,N_305,N_903);
and U2472 (N_2472,N_137,N_922);
or U2473 (N_2473,N_598,N_731);
or U2474 (N_2474,N_387,N_631);
and U2475 (N_2475,N_299,N_463);
and U2476 (N_2476,N_1443,N_507);
nand U2477 (N_2477,N_1625,N_383);
nor U2478 (N_2478,N_1936,N_1930);
and U2479 (N_2479,N_1646,N_1150);
nor U2480 (N_2480,N_267,N_781);
or U2481 (N_2481,N_1772,N_1848);
or U2482 (N_2482,N_6,N_1470);
nor U2483 (N_2483,N_1731,N_1015);
nor U2484 (N_2484,N_1021,N_800);
and U2485 (N_2485,N_835,N_1429);
nand U2486 (N_2486,N_653,N_1852);
or U2487 (N_2487,N_996,N_1079);
or U2488 (N_2488,N_27,N_1246);
or U2489 (N_2489,N_1406,N_1438);
nor U2490 (N_2490,N_1805,N_1104);
nor U2491 (N_2491,N_1263,N_1425);
nand U2492 (N_2492,N_1148,N_906);
nor U2493 (N_2493,N_1235,N_411);
xnor U2494 (N_2494,N_1370,N_1485);
nand U2495 (N_2495,N_32,N_10);
and U2496 (N_2496,N_1603,N_500);
nand U2497 (N_2497,N_718,N_728);
or U2498 (N_2498,N_1741,N_450);
nor U2499 (N_2499,N_714,N_1130);
nand U2500 (N_2500,N_1889,N_1501);
and U2501 (N_2501,N_8,N_988);
nor U2502 (N_2502,N_769,N_1584);
nor U2503 (N_2503,N_541,N_668);
nor U2504 (N_2504,N_1982,N_932);
nor U2505 (N_2505,N_624,N_247);
and U2506 (N_2506,N_192,N_243);
and U2507 (N_2507,N_43,N_1991);
nand U2508 (N_2508,N_398,N_211);
nor U2509 (N_2509,N_1567,N_1022);
nand U2510 (N_2510,N_255,N_799);
nor U2511 (N_2511,N_1012,N_536);
nand U2512 (N_2512,N_866,N_748);
or U2513 (N_2513,N_14,N_1824);
nor U2514 (N_2514,N_950,N_1313);
nor U2515 (N_2515,N_39,N_1692);
and U2516 (N_2516,N_1380,N_1016);
or U2517 (N_2517,N_1336,N_986);
nand U2518 (N_2518,N_987,N_376);
nand U2519 (N_2519,N_128,N_1442);
and U2520 (N_2520,N_875,N_824);
or U2521 (N_2521,N_1472,N_1872);
nand U2522 (N_2522,N_1786,N_429);
nand U2523 (N_2523,N_268,N_1191);
and U2524 (N_2524,N_839,N_654);
nand U2525 (N_2525,N_343,N_1471);
nand U2526 (N_2526,N_1825,N_895);
nand U2527 (N_2527,N_842,N_1706);
and U2528 (N_2528,N_1173,N_395);
and U2529 (N_2529,N_465,N_1596);
or U2530 (N_2530,N_403,N_224);
nand U2531 (N_2531,N_214,N_423);
and U2532 (N_2532,N_2,N_50);
nand U2533 (N_2533,N_302,N_1796);
nor U2534 (N_2534,N_921,N_1802);
nand U2535 (N_2535,N_226,N_1109);
or U2536 (N_2536,N_1811,N_1176);
nor U2537 (N_2537,N_1197,N_98);
nand U2538 (N_2538,N_553,N_68);
nor U2539 (N_2539,N_297,N_1629);
or U2540 (N_2540,N_193,N_1328);
and U2541 (N_2541,N_1320,N_609);
or U2542 (N_2542,N_1108,N_1688);
nand U2543 (N_2543,N_1512,N_86);
and U2544 (N_2544,N_212,N_233);
nor U2545 (N_2545,N_898,N_1602);
nand U2546 (N_2546,N_1225,N_1151);
or U2547 (N_2547,N_478,N_1159);
or U2548 (N_2548,N_293,N_1721);
xor U2549 (N_2549,N_1224,N_1144);
nor U2550 (N_2550,N_1733,N_1689);
nor U2551 (N_2551,N_1300,N_1125);
or U2552 (N_2552,N_1950,N_1466);
nand U2553 (N_2553,N_1106,N_687);
nand U2554 (N_2554,N_1617,N_1526);
nand U2555 (N_2555,N_1132,N_11);
nor U2556 (N_2556,N_1493,N_1269);
or U2557 (N_2557,N_344,N_332);
nand U2558 (N_2558,N_1628,N_222);
and U2559 (N_2559,N_1785,N_1896);
nand U2560 (N_2560,N_1685,N_1346);
nor U2561 (N_2561,N_738,N_289);
or U2562 (N_2562,N_1750,N_1854);
nor U2563 (N_2563,N_1601,N_1640);
or U2564 (N_2564,N_793,N_1957);
nand U2565 (N_2565,N_1914,N_931);
xnor U2566 (N_2566,N_115,N_1365);
nor U2567 (N_2567,N_848,N_431);
nand U2568 (N_2568,N_1178,N_1992);
and U2569 (N_2569,N_151,N_180);
and U2570 (N_2570,N_1943,N_1647);
and U2571 (N_2571,N_38,N_1367);
and U2572 (N_2572,N_551,N_1559);
and U2573 (N_2573,N_834,N_390);
nand U2574 (N_2574,N_1057,N_1038);
nor U2575 (N_2575,N_232,N_388);
nor U2576 (N_2576,N_991,N_1395);
nand U2577 (N_2577,N_1065,N_1521);
nand U2578 (N_2578,N_342,N_1788);
nand U2579 (N_2579,N_791,N_1445);
nor U2580 (N_2580,N_1633,N_1917);
or U2581 (N_2581,N_1765,N_1606);
nand U2582 (N_2582,N_1087,N_688);
nand U2583 (N_2583,N_825,N_1836);
nand U2584 (N_2584,N_1648,N_145);
and U2585 (N_2585,N_705,N_1027);
and U2586 (N_2586,N_378,N_1146);
nor U2587 (N_2587,N_590,N_1718);
nand U2588 (N_2588,N_894,N_1454);
nor U2589 (N_2589,N_672,N_1667);
and U2590 (N_2590,N_595,N_1272);
or U2591 (N_2591,N_1017,N_864);
and U2592 (N_2592,N_1895,N_556);
nor U2593 (N_2593,N_790,N_108);
and U2594 (N_2594,N_1315,N_179);
nor U2595 (N_2595,N_1123,N_1196);
nand U2596 (N_2596,N_861,N_646);
nand U2597 (N_2597,N_1212,N_717);
or U2598 (N_2598,N_1341,N_1306);
nand U2599 (N_2599,N_1243,N_1228);
or U2600 (N_2600,N_1055,N_1944);
nand U2601 (N_2601,N_914,N_347);
and U2602 (N_2602,N_368,N_712);
xor U2603 (N_2603,N_397,N_1794);
nor U2604 (N_2604,N_134,N_1873);
or U2605 (N_2605,N_634,N_1464);
nor U2606 (N_2606,N_1451,N_1770);
and U2607 (N_2607,N_1345,N_974);
and U2608 (N_2608,N_1790,N_1117);
nor U2609 (N_2609,N_1214,N_15);
or U2610 (N_2610,N_432,N_1882);
or U2611 (N_2611,N_379,N_1060);
nand U2612 (N_2612,N_415,N_1488);
and U2613 (N_2613,N_971,N_681);
nor U2614 (N_2614,N_1666,N_188);
or U2615 (N_2615,N_1396,N_1403);
nor U2616 (N_2616,N_1184,N_1133);
nand U2617 (N_2617,N_336,N_635);
and U2618 (N_2618,N_131,N_610);
nand U2619 (N_2619,N_497,N_1513);
and U2620 (N_2620,N_1050,N_1014);
or U2621 (N_2621,N_1351,N_1444);
nor U2622 (N_2622,N_726,N_949);
or U2623 (N_2623,N_223,N_730);
nand U2624 (N_2624,N_1761,N_404);
nand U2625 (N_2625,N_1934,N_402);
and U2626 (N_2626,N_1973,N_219);
nand U2627 (N_2627,N_962,N_1708);
nor U2628 (N_2628,N_1409,N_1862);
and U2629 (N_2629,N_1724,N_1393);
nand U2630 (N_2630,N_187,N_1180);
or U2631 (N_2631,N_274,N_163);
or U2632 (N_2632,N_1910,N_496);
or U2633 (N_2633,N_526,N_460);
nor U2634 (N_2634,N_641,N_946);
nand U2635 (N_2635,N_1918,N_1767);
nand U2636 (N_2636,N_916,N_1546);
nand U2637 (N_2637,N_1565,N_677);
nand U2638 (N_2638,N_1414,N_1084);
xor U2639 (N_2639,N_1901,N_1962);
nor U2640 (N_2640,N_1164,N_1419);
xnor U2641 (N_2641,N_280,N_1221);
nor U2642 (N_2642,N_1955,N_1326);
nand U2643 (N_2643,N_1072,N_1299);
or U2644 (N_2644,N_1866,N_1206);
nand U2645 (N_2645,N_1591,N_643);
nor U2646 (N_2646,N_1967,N_1227);
nor U2647 (N_2647,N_474,N_1749);
or U2648 (N_2648,N_741,N_1703);
and U2649 (N_2649,N_745,N_1335);
nor U2650 (N_2650,N_1984,N_126);
nand U2651 (N_2651,N_918,N_303);
or U2652 (N_2652,N_242,N_826);
or U2653 (N_2653,N_235,N_1101);
nand U2654 (N_2654,N_333,N_1303);
nand U2655 (N_2655,N_619,N_1641);
or U2656 (N_2656,N_1614,N_657);
nand U2657 (N_2657,N_803,N_1507);
nor U2658 (N_2658,N_853,N_499);
or U2659 (N_2659,N_1288,N_1799);
nor U2660 (N_2660,N_1616,N_1147);
nor U2661 (N_2661,N_860,N_767);
nor U2662 (N_2662,N_1465,N_629);
nand U2663 (N_2663,N_503,N_1031);
or U2664 (N_2664,N_284,N_929);
nand U2665 (N_2665,N_1541,N_36);
or U2666 (N_2666,N_1068,N_1008);
nand U2667 (N_2667,N_171,N_273);
nand U2668 (N_2668,N_695,N_458);
or U2669 (N_2669,N_1107,N_809);
and U2670 (N_2670,N_22,N_1553);
and U2671 (N_2671,N_435,N_516);
and U2672 (N_2672,N_1600,N_106);
or U2673 (N_2673,N_1563,N_952);
nand U2674 (N_2674,N_1937,N_244);
and U2675 (N_2675,N_729,N_679);
nand U2676 (N_2676,N_1755,N_1814);
nor U2677 (N_2677,N_787,N_1986);
and U2678 (N_2678,N_544,N_1494);
or U2679 (N_2679,N_1890,N_355);
nor U2680 (N_2680,N_1278,N_1302);
and U2681 (N_2681,N_1583,N_1473);
nor U2682 (N_2682,N_736,N_1138);
and U2683 (N_2683,N_843,N_479);
nand U2684 (N_2684,N_937,N_120);
or U2685 (N_2685,N_1152,N_692);
or U2686 (N_2686,N_699,N_1426);
and U2687 (N_2687,N_350,N_948);
or U2688 (N_2688,N_1325,N_1137);
nand U2689 (N_2689,N_618,N_1195);
nor U2690 (N_2690,N_596,N_1558);
and U2691 (N_2691,N_1892,N_1924);
nor U2692 (N_2692,N_524,N_48);
and U2693 (N_2693,N_1757,N_1960);
nor U2694 (N_2694,N_437,N_1338);
nor U2695 (N_2695,N_381,N_838);
and U2696 (N_2696,N_768,N_648);
nor U2697 (N_2697,N_757,N_1856);
nor U2698 (N_2698,N_154,N_1011);
xor U2699 (N_2699,N_94,N_1023);
and U2700 (N_2700,N_472,N_829);
and U2701 (N_2701,N_967,N_1376);
or U2702 (N_2702,N_1655,N_1270);
and U2703 (N_2703,N_1556,N_661);
or U2704 (N_2704,N_1618,N_1979);
and U2705 (N_2705,N_585,N_173);
nand U2706 (N_2706,N_1297,N_789);
or U2707 (N_2707,N_64,N_1175);
or U2708 (N_2708,N_568,N_639);
nand U2709 (N_2709,N_445,N_250);
nor U2710 (N_2710,N_1660,N_1434);
nor U2711 (N_2711,N_371,N_410);
and U2712 (N_2712,N_1920,N_591);
nor U2713 (N_2713,N_1268,N_1452);
nand U2714 (N_2714,N_1121,N_626);
or U2715 (N_2715,N_1481,N_220);
nand U2716 (N_2716,N_764,N_1254);
or U2717 (N_2717,N_1815,N_1061);
and U2718 (N_2718,N_836,N_1974);
nor U2719 (N_2719,N_195,N_1669);
and U2720 (N_2720,N_959,N_915);
and U2721 (N_2721,N_1248,N_1875);
and U2722 (N_2722,N_1019,N_1739);
nand U2723 (N_2723,N_40,N_945);
nand U2724 (N_2724,N_569,N_49);
nor U2725 (N_2725,N_758,N_1056);
nor U2726 (N_2726,N_1970,N_1018);
or U2727 (N_2727,N_59,N_927);
and U2728 (N_2728,N_1371,N_105);
nand U2729 (N_2729,N_1145,N_434);
or U2730 (N_2730,N_1399,N_511);
nand U2731 (N_2731,N_807,N_580);
or U2732 (N_2732,N_1885,N_876);
nor U2733 (N_2733,N_582,N_733);
nand U2734 (N_2734,N_1105,N_514);
or U2735 (N_2735,N_1620,N_1124);
and U2736 (N_2736,N_882,N_642);
or U2737 (N_2737,N_288,N_976);
or U2738 (N_2738,N_433,N_1205);
or U2739 (N_2739,N_28,N_1255);
or U2740 (N_2740,N_531,N_129);
or U2741 (N_2741,N_354,N_823);
and U2742 (N_2742,N_1066,N_69);
or U2743 (N_2743,N_1710,N_1448);
or U2744 (N_2744,N_1329,N_308);
nor U2745 (N_2745,N_1277,N_380);
nor U2746 (N_2746,N_121,N_1294);
or U2747 (N_2747,N_30,N_97);
nor U2748 (N_2748,N_1809,N_412);
and U2749 (N_2749,N_84,N_933);
and U2750 (N_2750,N_1461,N_704);
and U2751 (N_2751,N_1360,N_788);
and U2752 (N_2752,N_1085,N_965);
and U2753 (N_2753,N_1753,N_1778);
and U2754 (N_2754,N_858,N_1536);
and U2755 (N_2755,N_1193,N_1213);
or U2756 (N_2756,N_941,N_393);
or U2757 (N_2757,N_1436,N_622);
or U2758 (N_2758,N_892,N_1554);
nor U2759 (N_2759,N_178,N_1745);
or U2760 (N_2760,N_441,N_735);
and U2761 (N_2761,N_1758,N_102);
or U2762 (N_2762,N_559,N_1636);
and U2763 (N_2763,N_1261,N_782);
nand U2764 (N_2764,N_78,N_935);
or U2765 (N_2765,N_862,N_1102);
or U2766 (N_2766,N_1547,N_889);
nand U2767 (N_2767,N_1697,N_147);
nand U2768 (N_2768,N_1635,N_1694);
xor U2769 (N_2769,N_1308,N_318);
and U2770 (N_2770,N_1981,N_488);
nor U2771 (N_2771,N_1826,N_275);
nand U2772 (N_2772,N_1037,N_1430);
nand U2773 (N_2773,N_908,N_221);
nor U2774 (N_2774,N_1932,N_1177);
or U2775 (N_2775,N_1292,N_1579);
nand U2776 (N_2776,N_884,N_759);
nand U2777 (N_2777,N_262,N_1479);
or U2778 (N_2778,N_1857,N_760);
or U2779 (N_2779,N_200,N_453);
xor U2780 (N_2780,N_644,N_1208);
or U2781 (N_2781,N_919,N_1539);
and U2782 (N_2782,N_723,N_414);
and U2783 (N_2783,N_1382,N_532);
and U2784 (N_2784,N_408,N_1103);
and U2785 (N_2785,N_888,N_752);
or U2786 (N_2786,N_601,N_353);
xor U2787 (N_2787,N_1519,N_1449);
nor U2788 (N_2788,N_419,N_1529);
or U2789 (N_2789,N_1082,N_1119);
or U2790 (N_2790,N_253,N_1122);
nor U2791 (N_2791,N_1456,N_827);
nor U2792 (N_2792,N_80,N_581);
and U2793 (N_2793,N_1941,N_1726);
nor U2794 (N_2794,N_578,N_1665);
and U2795 (N_2795,N_1039,N_944);
and U2796 (N_2796,N_306,N_956);
nor U2797 (N_2797,N_1202,N_621);
nor U2798 (N_2798,N_773,N_659);
or U2799 (N_2799,N_636,N_1052);
and U2800 (N_2800,N_863,N_792);
or U2801 (N_2801,N_502,N_426);
and U2802 (N_2802,N_4,N_348);
xor U2803 (N_2803,N_1129,N_645);
nand U2804 (N_2804,N_1279,N_47);
nor U2805 (N_2805,N_1486,N_1953);
nand U2806 (N_2806,N_1232,N_1673);
and U2807 (N_2807,N_34,N_968);
and U2808 (N_2808,N_71,N_1705);
and U2809 (N_2809,N_603,N_504);
or U2810 (N_2810,N_887,N_196);
nor U2811 (N_2811,N_1631,N_202);
and U2812 (N_2812,N_473,N_311);
or U2813 (N_2813,N_509,N_125);
or U2814 (N_2814,N_495,N_664);
nor U2815 (N_2815,N_1078,N_1398);
or U2816 (N_2816,N_1181,N_1530);
nor U2817 (N_2817,N_364,N_924);
and U2818 (N_2818,N_1167,N_710);
and U2819 (N_2819,N_1997,N_913);
and U2820 (N_2820,N_1961,N_1034);
nor U2821 (N_2821,N_89,N_1355);
and U2822 (N_2822,N_771,N_798);
and U2823 (N_2823,N_770,N_808);
and U2824 (N_2824,N_1915,N_37);
nor U2825 (N_2825,N_1969,N_248);
and U2826 (N_2826,N_240,N_96);
or U2827 (N_2827,N_1691,N_1158);
nand U2828 (N_2828,N_1353,N_510);
xnor U2829 (N_2829,N_1621,N_357);
or U2830 (N_2830,N_640,N_1998);
nor U2831 (N_2831,N_392,N_122);
nand U2832 (N_2832,N_337,N_327);
and U2833 (N_2833,N_716,N_1334);
nor U2834 (N_2834,N_1046,N_1032);
and U2835 (N_2835,N_143,N_1343);
or U2836 (N_2836,N_1410,N_13);
nand U2837 (N_2837,N_742,N_1166);
or U2838 (N_2838,N_780,N_936);
nand U2839 (N_2839,N_1587,N_542);
nor U2840 (N_2840,N_777,N_700);
nand U2841 (N_2841,N_1391,N_1331);
or U2842 (N_2842,N_45,N_1354);
or U2843 (N_2843,N_1260,N_61);
or U2844 (N_2844,N_335,N_1131);
nand U2845 (N_2845,N_17,N_1642);
or U2846 (N_2846,N_1009,N_1401);
nand U2847 (N_2847,N_1735,N_1067);
nor U2848 (N_2848,N_1514,N_990);
or U2849 (N_2849,N_190,N_1492);
nand U2850 (N_2850,N_266,N_158);
nor U2851 (N_2851,N_1424,N_1925);
or U2852 (N_2852,N_1455,N_775);
nand U2853 (N_2853,N_1342,N_1054);
and U2854 (N_2854,N_1368,N_317);
nor U2855 (N_2855,N_548,N_1352);
nand U2856 (N_2856,N_1985,N_501);
nand U2857 (N_2857,N_1200,N_1222);
or U2858 (N_2858,N_865,N_1432);
and U2859 (N_2859,N_1599,N_56);
or U2860 (N_2860,N_1304,N_1945);
nor U2861 (N_2861,N_1573,N_1933);
or U2862 (N_2862,N_1170,N_1552);
nand U2863 (N_2863,N_879,N_1610);
and U2864 (N_2864,N_572,N_52);
and U2865 (N_2865,N_42,N_587);
xor U2866 (N_2866,N_92,N_1717);
nor U2867 (N_2867,N_1858,N_1619);
or U2868 (N_2868,N_523,N_1389);
nand U2869 (N_2869,N_605,N_763);
and U2870 (N_2870,N_1744,N_439);
nand U2871 (N_2871,N_1207,N_1295);
or U2872 (N_2872,N_1381,N_483);
nand U2873 (N_2873,N_616,N_1543);
nand U2874 (N_2874,N_1562,N_1435);
nand U2875 (N_2875,N_1938,N_1128);
nor U2876 (N_2876,N_1115,N_747);
and U2877 (N_2877,N_1657,N_1231);
nand U2878 (N_2878,N_127,N_1676);
nor U2879 (N_2879,N_680,N_1659);
nor U2880 (N_2880,N_1024,N_33);
xor U2881 (N_2881,N_135,N_310);
or U2882 (N_2882,N_323,N_186);
and U2883 (N_2883,N_1462,N_113);
and U2884 (N_2884,N_577,N_1716);
xnor U2885 (N_2885,N_1702,N_296);
or U2886 (N_2886,N_665,N_506);
nand U2887 (N_2887,N_1006,N_1865);
and U2888 (N_2888,N_400,N_811);
nor U2889 (N_2889,N_1307,N_637);
nand U2890 (N_2890,N_633,N_814);
or U2891 (N_2891,N_349,N_1714);
or U2892 (N_2892,N_1384,N_112);
or U2893 (N_2893,N_1071,N_132);
nor U2894 (N_2894,N_194,N_880);
nand U2895 (N_2895,N_389,N_1988);
and U2896 (N_2896,N_1623,N_1894);
nor U2897 (N_2897,N_981,N_725);
nor U2898 (N_2898,N_1361,N_1074);
nand U2899 (N_2899,N_1058,N_1581);
and U2900 (N_2900,N_722,N_83);
nor U2901 (N_2901,N_576,N_1517);
or U2902 (N_2902,N_217,N_1916);
nand U2903 (N_2903,N_476,N_1774);
and U2904 (N_2904,N_1612,N_24);
and U2905 (N_2905,N_418,N_1956);
nor U2906 (N_2906,N_907,N_1779);
xor U2907 (N_2907,N_1097,N_216);
nor U2908 (N_2908,N_1976,N_1229);
nand U2909 (N_2909,N_1756,N_1264);
or U2910 (N_2910,N_1939,N_1408);
or U2911 (N_2911,N_1906,N_259);
or U2912 (N_2912,N_1417,N_1394);
nand U2913 (N_2913,N_99,N_175);
and U2914 (N_2914,N_285,N_234);
nand U2915 (N_2915,N_1134,N_984);
nand U2916 (N_2916,N_1611,N_1182);
or U2917 (N_2917,N_1265,N_467);
and U2918 (N_2918,N_685,N_144);
or U2919 (N_2919,N_683,N_361);
xor U2920 (N_2920,N_1849,N_795);
nor U2921 (N_2921,N_1035,N_893);
and U2922 (N_2922,N_1002,N_1698);
nand U2923 (N_2923,N_1332,N_168);
and U2924 (N_2924,N_1276,N_1632);
nor U2925 (N_2925,N_292,N_844);
xnor U2926 (N_2926,N_1942,N_1400);
nor U2927 (N_2927,N_1188,N_1561);
or U2928 (N_2928,N_1324,N_1511);
nor U2929 (N_2929,N_1592,N_902);
nand U2930 (N_2930,N_625,N_570);
nor U2931 (N_2931,N_67,N_1316);
nor U2932 (N_2932,N_1842,N_1044);
and U2933 (N_2933,N_1422,N_1877);
nor U2934 (N_2934,N_1358,N_859);
nand U2935 (N_2935,N_1605,N_1760);
or U2936 (N_2936,N_1030,N_1590);
nand U2937 (N_2937,N_1784,N_816);
and U2938 (N_2938,N_1931,N_436);
or U2939 (N_2939,N_1838,N_1585);
nor U2940 (N_2940,N_1402,N_162);
or U2941 (N_2941,N_1977,N_1287);
nand U2942 (N_2942,N_1088,N_1537);
nor U2943 (N_2943,N_1198,N_165);
or U2944 (N_2944,N_602,N_155);
nor U2945 (N_2945,N_1226,N_1069);
xor U2946 (N_2946,N_530,N_1305);
nor U2947 (N_2947,N_1185,N_468);
nand U2948 (N_2948,N_1112,N_215);
or U2949 (N_2949,N_269,N_1282);
and U2950 (N_2950,N_152,N_1239);
and U2951 (N_2951,N_673,N_1574);
and U2952 (N_2952,N_443,N_1847);
and U2953 (N_2953,N_1505,N_167);
or U2954 (N_2954,N_160,N_428);
or U2955 (N_2955,N_953,N_1171);
nor U2956 (N_2956,N_806,N_539);
and U2957 (N_2957,N_1908,N_584);
or U2958 (N_2958,N_1407,N_1701);
nand U2959 (N_2959,N_1392,N_1880);
nor U2960 (N_2960,N_1624,N_199);
nor U2961 (N_2961,N_1489,N_1597);
nor U2962 (N_2962,N_998,N_703);
nor U2963 (N_2963,N_1797,N_1588);
or U2964 (N_2964,N_1531,N_850);
and U2965 (N_2965,N_1457,N_1707);
nand U2966 (N_2966,N_1644,N_684);
nand U2967 (N_2967,N_313,N_1404);
nand U2968 (N_2968,N_1989,N_1812);
and U2969 (N_2969,N_1446,N_620);
and U2970 (N_2970,N_1905,N_1199);
or U2971 (N_2971,N_1662,N_1216);
and U2972 (N_2972,N_208,N_1801);
nor U2973 (N_2973,N_697,N_1860);
or U2974 (N_2974,N_513,N_229);
or U2975 (N_2975,N_1223,N_1627);
nand U2976 (N_2976,N_632,N_1902);
nand U2977 (N_2977,N_1630,N_1025);
or U2978 (N_2978,N_1919,N_739);
nor U2979 (N_2979,N_1086,N_1867);
nand U2980 (N_2980,N_558,N_1870);
nor U2981 (N_2981,N_385,N_1504);
nand U2982 (N_2982,N_1542,N_1948);
xnor U2983 (N_2983,N_1247,N_205);
nand U2984 (N_2984,N_1883,N_766);
and U2985 (N_2985,N_1980,N_1855);
or U2986 (N_2986,N_1549,N_579);
nor U2987 (N_2987,N_743,N_1020);
nand U2988 (N_2988,N_951,N_955);
or U2989 (N_2989,N_942,N_315);
or U2990 (N_2990,N_1696,N_185);
nor U2991 (N_2991,N_1861,N_369);
and U2992 (N_2992,N_857,N_623);
or U2993 (N_2993,N_1259,N_85);
xor U2994 (N_2994,N_422,N_1923);
nand U2995 (N_2995,N_482,N_599);
or U2996 (N_2996,N_1704,N_1285);
xnor U2997 (N_2997,N_1598,N_1298);
nand U2998 (N_2998,N_1789,N_1713);
nand U2999 (N_2999,N_1680,N_425);
or U3000 (N_3000,N_1845,N_1325);
nand U3001 (N_3001,N_307,N_48);
nor U3002 (N_3002,N_127,N_1053);
and U3003 (N_3003,N_1670,N_352);
nor U3004 (N_3004,N_63,N_698);
or U3005 (N_3005,N_655,N_1512);
and U3006 (N_3006,N_173,N_729);
nand U3007 (N_3007,N_673,N_1299);
nand U3008 (N_3008,N_1765,N_1508);
or U3009 (N_3009,N_59,N_288);
nand U3010 (N_3010,N_1043,N_1934);
or U3011 (N_3011,N_1165,N_1545);
and U3012 (N_3012,N_1964,N_351);
nand U3013 (N_3013,N_372,N_1629);
and U3014 (N_3014,N_1966,N_967);
nor U3015 (N_3015,N_251,N_1651);
nor U3016 (N_3016,N_834,N_1214);
and U3017 (N_3017,N_798,N_721);
or U3018 (N_3018,N_55,N_1617);
nor U3019 (N_3019,N_1122,N_678);
or U3020 (N_3020,N_390,N_1937);
nand U3021 (N_3021,N_1740,N_963);
and U3022 (N_3022,N_1563,N_886);
nand U3023 (N_3023,N_540,N_1358);
or U3024 (N_3024,N_1220,N_802);
nor U3025 (N_3025,N_1406,N_579);
nor U3026 (N_3026,N_272,N_1141);
or U3027 (N_3027,N_1713,N_1037);
nand U3028 (N_3028,N_55,N_409);
nand U3029 (N_3029,N_1242,N_1463);
nor U3030 (N_3030,N_695,N_780);
nand U3031 (N_3031,N_1091,N_122);
and U3032 (N_3032,N_1021,N_1683);
nor U3033 (N_3033,N_1358,N_1254);
or U3034 (N_3034,N_1612,N_1197);
xnor U3035 (N_3035,N_523,N_1052);
or U3036 (N_3036,N_1442,N_1148);
and U3037 (N_3037,N_1153,N_870);
nor U3038 (N_3038,N_444,N_1049);
nand U3039 (N_3039,N_492,N_1105);
nand U3040 (N_3040,N_1325,N_710);
and U3041 (N_3041,N_681,N_220);
nor U3042 (N_3042,N_707,N_711);
and U3043 (N_3043,N_1852,N_1233);
or U3044 (N_3044,N_1683,N_1014);
or U3045 (N_3045,N_1400,N_566);
nor U3046 (N_3046,N_217,N_1893);
or U3047 (N_3047,N_817,N_1205);
or U3048 (N_3048,N_1109,N_1704);
or U3049 (N_3049,N_302,N_562);
nand U3050 (N_3050,N_876,N_560);
nand U3051 (N_3051,N_298,N_235);
and U3052 (N_3052,N_378,N_339);
nor U3053 (N_3053,N_64,N_1511);
nand U3054 (N_3054,N_16,N_1529);
nor U3055 (N_3055,N_33,N_1058);
nor U3056 (N_3056,N_1872,N_917);
nand U3057 (N_3057,N_602,N_821);
nand U3058 (N_3058,N_1466,N_1291);
nand U3059 (N_3059,N_235,N_353);
and U3060 (N_3060,N_147,N_227);
nand U3061 (N_3061,N_1876,N_532);
or U3062 (N_3062,N_1836,N_985);
xnor U3063 (N_3063,N_1444,N_526);
nor U3064 (N_3064,N_1066,N_1028);
and U3065 (N_3065,N_594,N_940);
and U3066 (N_3066,N_159,N_633);
or U3067 (N_3067,N_418,N_1778);
xnor U3068 (N_3068,N_1936,N_1991);
and U3069 (N_3069,N_1914,N_725);
nand U3070 (N_3070,N_243,N_1018);
nand U3071 (N_3071,N_24,N_1859);
nand U3072 (N_3072,N_664,N_1148);
or U3073 (N_3073,N_149,N_737);
nand U3074 (N_3074,N_402,N_1563);
nor U3075 (N_3075,N_645,N_67);
nor U3076 (N_3076,N_1409,N_573);
nand U3077 (N_3077,N_417,N_146);
nand U3078 (N_3078,N_1826,N_1886);
nand U3079 (N_3079,N_650,N_383);
or U3080 (N_3080,N_1312,N_706);
nand U3081 (N_3081,N_319,N_701);
nor U3082 (N_3082,N_1204,N_1511);
nor U3083 (N_3083,N_1031,N_1930);
or U3084 (N_3084,N_754,N_138);
and U3085 (N_3085,N_1236,N_1933);
or U3086 (N_3086,N_787,N_1021);
nand U3087 (N_3087,N_1254,N_317);
nor U3088 (N_3088,N_1826,N_1459);
and U3089 (N_3089,N_1018,N_1199);
nand U3090 (N_3090,N_1217,N_1780);
and U3091 (N_3091,N_300,N_1114);
and U3092 (N_3092,N_1916,N_1949);
nor U3093 (N_3093,N_3,N_1504);
nor U3094 (N_3094,N_264,N_1238);
and U3095 (N_3095,N_1648,N_922);
nor U3096 (N_3096,N_1811,N_705);
and U3097 (N_3097,N_784,N_288);
and U3098 (N_3098,N_509,N_699);
and U3099 (N_3099,N_969,N_186);
or U3100 (N_3100,N_1938,N_1959);
nor U3101 (N_3101,N_206,N_1682);
nor U3102 (N_3102,N_86,N_1796);
or U3103 (N_3103,N_1545,N_1686);
and U3104 (N_3104,N_140,N_1305);
or U3105 (N_3105,N_662,N_1458);
or U3106 (N_3106,N_1027,N_1655);
or U3107 (N_3107,N_1619,N_548);
or U3108 (N_3108,N_750,N_1766);
or U3109 (N_3109,N_1735,N_1545);
or U3110 (N_3110,N_231,N_232);
nor U3111 (N_3111,N_1297,N_1711);
nor U3112 (N_3112,N_1231,N_719);
or U3113 (N_3113,N_1097,N_70);
or U3114 (N_3114,N_1969,N_54);
nand U3115 (N_3115,N_326,N_642);
nor U3116 (N_3116,N_922,N_847);
nor U3117 (N_3117,N_486,N_1388);
xor U3118 (N_3118,N_410,N_1673);
or U3119 (N_3119,N_105,N_847);
nand U3120 (N_3120,N_845,N_52);
xor U3121 (N_3121,N_568,N_77);
nor U3122 (N_3122,N_1383,N_1660);
nor U3123 (N_3123,N_639,N_715);
nor U3124 (N_3124,N_1802,N_418);
nand U3125 (N_3125,N_1504,N_1574);
nor U3126 (N_3126,N_130,N_655);
nor U3127 (N_3127,N_225,N_678);
xnor U3128 (N_3128,N_1696,N_683);
xnor U3129 (N_3129,N_643,N_1351);
or U3130 (N_3130,N_1250,N_492);
or U3131 (N_3131,N_1914,N_139);
and U3132 (N_3132,N_1940,N_790);
nand U3133 (N_3133,N_4,N_13);
or U3134 (N_3134,N_994,N_56);
nor U3135 (N_3135,N_1526,N_82);
nor U3136 (N_3136,N_1247,N_347);
nor U3137 (N_3137,N_158,N_898);
or U3138 (N_3138,N_557,N_113);
or U3139 (N_3139,N_1715,N_1666);
or U3140 (N_3140,N_934,N_219);
or U3141 (N_3141,N_1862,N_269);
nand U3142 (N_3142,N_1539,N_1656);
nand U3143 (N_3143,N_1684,N_327);
or U3144 (N_3144,N_226,N_1595);
or U3145 (N_3145,N_1808,N_632);
or U3146 (N_3146,N_1755,N_1756);
or U3147 (N_3147,N_375,N_1657);
or U3148 (N_3148,N_1553,N_1988);
nor U3149 (N_3149,N_904,N_439);
and U3150 (N_3150,N_1477,N_1266);
and U3151 (N_3151,N_294,N_909);
nand U3152 (N_3152,N_449,N_640);
and U3153 (N_3153,N_630,N_832);
or U3154 (N_3154,N_575,N_581);
nor U3155 (N_3155,N_1454,N_1620);
or U3156 (N_3156,N_443,N_437);
or U3157 (N_3157,N_1525,N_130);
or U3158 (N_3158,N_677,N_1676);
and U3159 (N_3159,N_631,N_1765);
nor U3160 (N_3160,N_361,N_1910);
or U3161 (N_3161,N_1403,N_1013);
nor U3162 (N_3162,N_1806,N_1235);
or U3163 (N_3163,N_450,N_1647);
nor U3164 (N_3164,N_1357,N_612);
xnor U3165 (N_3165,N_1793,N_353);
and U3166 (N_3166,N_1538,N_158);
nor U3167 (N_3167,N_1064,N_1815);
and U3168 (N_3168,N_385,N_1728);
nand U3169 (N_3169,N_1487,N_1617);
or U3170 (N_3170,N_350,N_1047);
nand U3171 (N_3171,N_1140,N_479);
nand U3172 (N_3172,N_1703,N_1919);
and U3173 (N_3173,N_1949,N_863);
nand U3174 (N_3174,N_1344,N_1136);
nor U3175 (N_3175,N_1938,N_1361);
nand U3176 (N_3176,N_25,N_1930);
or U3177 (N_3177,N_1182,N_253);
or U3178 (N_3178,N_521,N_1577);
nor U3179 (N_3179,N_116,N_42);
nand U3180 (N_3180,N_510,N_928);
nand U3181 (N_3181,N_848,N_1953);
nor U3182 (N_3182,N_483,N_1688);
nor U3183 (N_3183,N_1985,N_1064);
xor U3184 (N_3184,N_1382,N_889);
nor U3185 (N_3185,N_1645,N_369);
and U3186 (N_3186,N_1061,N_1179);
nor U3187 (N_3187,N_1252,N_1965);
nand U3188 (N_3188,N_1,N_1385);
and U3189 (N_3189,N_238,N_715);
nor U3190 (N_3190,N_1522,N_677);
nor U3191 (N_3191,N_1037,N_280);
nor U3192 (N_3192,N_1097,N_42);
and U3193 (N_3193,N_494,N_822);
nor U3194 (N_3194,N_244,N_1524);
and U3195 (N_3195,N_1507,N_279);
nand U3196 (N_3196,N_1601,N_635);
and U3197 (N_3197,N_1265,N_431);
or U3198 (N_3198,N_309,N_648);
or U3199 (N_3199,N_773,N_614);
or U3200 (N_3200,N_1609,N_1147);
nand U3201 (N_3201,N_1443,N_307);
or U3202 (N_3202,N_968,N_458);
and U3203 (N_3203,N_980,N_121);
nor U3204 (N_3204,N_1832,N_1694);
or U3205 (N_3205,N_1028,N_1722);
nor U3206 (N_3206,N_632,N_1598);
nor U3207 (N_3207,N_261,N_1027);
nand U3208 (N_3208,N_197,N_1741);
nor U3209 (N_3209,N_1784,N_1207);
nor U3210 (N_3210,N_704,N_7);
and U3211 (N_3211,N_1836,N_547);
nor U3212 (N_3212,N_544,N_1152);
nand U3213 (N_3213,N_271,N_1305);
or U3214 (N_3214,N_202,N_854);
and U3215 (N_3215,N_1411,N_689);
or U3216 (N_3216,N_1841,N_685);
nand U3217 (N_3217,N_1372,N_1993);
or U3218 (N_3218,N_760,N_921);
nor U3219 (N_3219,N_1988,N_541);
or U3220 (N_3220,N_858,N_372);
nor U3221 (N_3221,N_1363,N_1399);
nand U3222 (N_3222,N_1359,N_992);
or U3223 (N_3223,N_403,N_1560);
nand U3224 (N_3224,N_1519,N_545);
nor U3225 (N_3225,N_518,N_1722);
or U3226 (N_3226,N_280,N_546);
or U3227 (N_3227,N_849,N_1263);
and U3228 (N_3228,N_1920,N_597);
and U3229 (N_3229,N_538,N_1300);
and U3230 (N_3230,N_502,N_990);
nand U3231 (N_3231,N_1881,N_1146);
and U3232 (N_3232,N_376,N_1920);
or U3233 (N_3233,N_855,N_1348);
or U3234 (N_3234,N_224,N_586);
nand U3235 (N_3235,N_1268,N_265);
nand U3236 (N_3236,N_1866,N_956);
nor U3237 (N_3237,N_1528,N_715);
or U3238 (N_3238,N_232,N_1253);
or U3239 (N_3239,N_1949,N_87);
or U3240 (N_3240,N_816,N_1763);
nor U3241 (N_3241,N_1614,N_455);
or U3242 (N_3242,N_241,N_354);
and U3243 (N_3243,N_280,N_548);
nor U3244 (N_3244,N_1819,N_433);
nand U3245 (N_3245,N_965,N_680);
nor U3246 (N_3246,N_61,N_453);
nand U3247 (N_3247,N_45,N_484);
or U3248 (N_3248,N_401,N_130);
or U3249 (N_3249,N_1779,N_111);
nand U3250 (N_3250,N_725,N_1975);
or U3251 (N_3251,N_785,N_349);
nor U3252 (N_3252,N_1416,N_1047);
nand U3253 (N_3253,N_250,N_386);
and U3254 (N_3254,N_1733,N_1573);
or U3255 (N_3255,N_143,N_155);
nor U3256 (N_3256,N_660,N_818);
nand U3257 (N_3257,N_1350,N_73);
nand U3258 (N_3258,N_1917,N_460);
and U3259 (N_3259,N_1181,N_193);
nor U3260 (N_3260,N_913,N_625);
or U3261 (N_3261,N_1646,N_556);
nand U3262 (N_3262,N_804,N_1371);
and U3263 (N_3263,N_464,N_953);
nand U3264 (N_3264,N_971,N_1870);
nand U3265 (N_3265,N_957,N_1142);
nand U3266 (N_3266,N_1272,N_1284);
and U3267 (N_3267,N_1242,N_674);
nor U3268 (N_3268,N_1506,N_930);
and U3269 (N_3269,N_1140,N_432);
nand U3270 (N_3270,N_645,N_1050);
nand U3271 (N_3271,N_277,N_598);
and U3272 (N_3272,N_90,N_1732);
nor U3273 (N_3273,N_511,N_849);
nor U3274 (N_3274,N_1456,N_1164);
or U3275 (N_3275,N_551,N_1933);
or U3276 (N_3276,N_1609,N_1295);
nor U3277 (N_3277,N_1149,N_1863);
nor U3278 (N_3278,N_792,N_1663);
and U3279 (N_3279,N_1489,N_1958);
xnor U3280 (N_3280,N_1118,N_205);
nand U3281 (N_3281,N_1499,N_1610);
nor U3282 (N_3282,N_1057,N_711);
nor U3283 (N_3283,N_1134,N_1109);
and U3284 (N_3284,N_1848,N_788);
or U3285 (N_3285,N_213,N_1338);
nor U3286 (N_3286,N_258,N_997);
xnor U3287 (N_3287,N_1419,N_1951);
and U3288 (N_3288,N_816,N_847);
or U3289 (N_3289,N_692,N_1695);
or U3290 (N_3290,N_628,N_1299);
nand U3291 (N_3291,N_1305,N_1213);
and U3292 (N_3292,N_478,N_1783);
nand U3293 (N_3293,N_1260,N_1310);
or U3294 (N_3294,N_1271,N_854);
and U3295 (N_3295,N_111,N_179);
nand U3296 (N_3296,N_1219,N_176);
or U3297 (N_3297,N_1930,N_851);
and U3298 (N_3298,N_1568,N_1660);
nor U3299 (N_3299,N_1207,N_290);
nor U3300 (N_3300,N_1735,N_511);
nand U3301 (N_3301,N_1033,N_1600);
nand U3302 (N_3302,N_1898,N_800);
nand U3303 (N_3303,N_1530,N_1911);
and U3304 (N_3304,N_1807,N_1821);
or U3305 (N_3305,N_1539,N_658);
or U3306 (N_3306,N_238,N_1388);
or U3307 (N_3307,N_1485,N_1216);
and U3308 (N_3308,N_1811,N_1705);
nor U3309 (N_3309,N_150,N_208);
nor U3310 (N_3310,N_750,N_34);
or U3311 (N_3311,N_1267,N_1162);
nor U3312 (N_3312,N_1661,N_675);
or U3313 (N_3313,N_1568,N_1852);
and U3314 (N_3314,N_502,N_627);
nand U3315 (N_3315,N_192,N_1221);
xnor U3316 (N_3316,N_929,N_420);
or U3317 (N_3317,N_153,N_18);
and U3318 (N_3318,N_1946,N_1858);
nor U3319 (N_3319,N_1732,N_357);
and U3320 (N_3320,N_423,N_86);
or U3321 (N_3321,N_866,N_1289);
or U3322 (N_3322,N_1274,N_764);
nor U3323 (N_3323,N_202,N_1470);
or U3324 (N_3324,N_1303,N_1606);
nor U3325 (N_3325,N_1975,N_783);
nand U3326 (N_3326,N_335,N_772);
nor U3327 (N_3327,N_1034,N_994);
or U3328 (N_3328,N_379,N_1907);
and U3329 (N_3329,N_1584,N_1612);
or U3330 (N_3330,N_1095,N_721);
or U3331 (N_3331,N_1279,N_920);
and U3332 (N_3332,N_677,N_323);
and U3333 (N_3333,N_551,N_1543);
and U3334 (N_3334,N_1520,N_1193);
and U3335 (N_3335,N_1652,N_1684);
and U3336 (N_3336,N_294,N_1547);
nand U3337 (N_3337,N_1083,N_1600);
or U3338 (N_3338,N_535,N_482);
or U3339 (N_3339,N_1486,N_1110);
or U3340 (N_3340,N_249,N_503);
nor U3341 (N_3341,N_797,N_1536);
and U3342 (N_3342,N_276,N_248);
or U3343 (N_3343,N_3,N_1921);
and U3344 (N_3344,N_779,N_1945);
nand U3345 (N_3345,N_151,N_486);
nand U3346 (N_3346,N_1100,N_477);
and U3347 (N_3347,N_412,N_304);
and U3348 (N_3348,N_782,N_1654);
and U3349 (N_3349,N_1324,N_547);
nor U3350 (N_3350,N_400,N_1621);
nor U3351 (N_3351,N_607,N_764);
nand U3352 (N_3352,N_576,N_236);
or U3353 (N_3353,N_1092,N_1810);
nor U3354 (N_3354,N_65,N_391);
and U3355 (N_3355,N_919,N_1457);
nor U3356 (N_3356,N_754,N_1919);
and U3357 (N_3357,N_1011,N_264);
nor U3358 (N_3358,N_1425,N_21);
nand U3359 (N_3359,N_32,N_937);
or U3360 (N_3360,N_1543,N_792);
and U3361 (N_3361,N_759,N_671);
nand U3362 (N_3362,N_1989,N_1758);
nand U3363 (N_3363,N_1901,N_810);
and U3364 (N_3364,N_860,N_770);
nand U3365 (N_3365,N_856,N_423);
and U3366 (N_3366,N_617,N_837);
nand U3367 (N_3367,N_441,N_607);
nand U3368 (N_3368,N_1622,N_1836);
nor U3369 (N_3369,N_734,N_29);
or U3370 (N_3370,N_123,N_906);
nand U3371 (N_3371,N_484,N_1682);
nor U3372 (N_3372,N_1329,N_1417);
or U3373 (N_3373,N_1503,N_1023);
or U3374 (N_3374,N_405,N_1042);
or U3375 (N_3375,N_1209,N_677);
nor U3376 (N_3376,N_526,N_1778);
and U3377 (N_3377,N_957,N_1563);
or U3378 (N_3378,N_1438,N_454);
nor U3379 (N_3379,N_1012,N_1662);
nand U3380 (N_3380,N_850,N_192);
or U3381 (N_3381,N_1923,N_1741);
and U3382 (N_3382,N_107,N_879);
and U3383 (N_3383,N_683,N_498);
nand U3384 (N_3384,N_1996,N_1721);
nand U3385 (N_3385,N_1099,N_1827);
nor U3386 (N_3386,N_400,N_519);
and U3387 (N_3387,N_1255,N_1629);
nand U3388 (N_3388,N_1834,N_972);
or U3389 (N_3389,N_439,N_1388);
nand U3390 (N_3390,N_912,N_596);
and U3391 (N_3391,N_1890,N_1903);
and U3392 (N_3392,N_1366,N_598);
or U3393 (N_3393,N_1445,N_849);
nand U3394 (N_3394,N_384,N_1715);
or U3395 (N_3395,N_1874,N_1180);
or U3396 (N_3396,N_1742,N_1707);
and U3397 (N_3397,N_652,N_600);
and U3398 (N_3398,N_1681,N_688);
or U3399 (N_3399,N_954,N_142);
or U3400 (N_3400,N_1568,N_841);
and U3401 (N_3401,N_1309,N_71);
nor U3402 (N_3402,N_306,N_1838);
and U3403 (N_3403,N_576,N_778);
nor U3404 (N_3404,N_863,N_1193);
nor U3405 (N_3405,N_1432,N_1474);
xor U3406 (N_3406,N_1331,N_1168);
and U3407 (N_3407,N_770,N_1245);
or U3408 (N_3408,N_13,N_62);
or U3409 (N_3409,N_79,N_681);
or U3410 (N_3410,N_1415,N_15);
or U3411 (N_3411,N_827,N_986);
nor U3412 (N_3412,N_149,N_1278);
and U3413 (N_3413,N_1875,N_1491);
and U3414 (N_3414,N_1775,N_1364);
and U3415 (N_3415,N_517,N_267);
and U3416 (N_3416,N_348,N_279);
nor U3417 (N_3417,N_577,N_684);
and U3418 (N_3418,N_551,N_894);
nor U3419 (N_3419,N_740,N_405);
and U3420 (N_3420,N_1595,N_1601);
nand U3421 (N_3421,N_1740,N_997);
xnor U3422 (N_3422,N_784,N_1550);
or U3423 (N_3423,N_397,N_407);
or U3424 (N_3424,N_564,N_166);
nor U3425 (N_3425,N_572,N_995);
or U3426 (N_3426,N_1963,N_757);
and U3427 (N_3427,N_1113,N_1525);
or U3428 (N_3428,N_1783,N_1315);
nand U3429 (N_3429,N_1874,N_1794);
nand U3430 (N_3430,N_494,N_1821);
nand U3431 (N_3431,N_1824,N_1172);
or U3432 (N_3432,N_1009,N_1953);
nand U3433 (N_3433,N_1634,N_312);
xor U3434 (N_3434,N_7,N_26);
nor U3435 (N_3435,N_1242,N_820);
or U3436 (N_3436,N_471,N_1248);
nor U3437 (N_3437,N_182,N_351);
xor U3438 (N_3438,N_614,N_725);
or U3439 (N_3439,N_548,N_23);
or U3440 (N_3440,N_21,N_1494);
nor U3441 (N_3441,N_148,N_347);
nor U3442 (N_3442,N_1501,N_1404);
xnor U3443 (N_3443,N_1844,N_393);
nor U3444 (N_3444,N_1727,N_847);
nor U3445 (N_3445,N_629,N_1754);
or U3446 (N_3446,N_1055,N_926);
and U3447 (N_3447,N_318,N_1399);
nand U3448 (N_3448,N_722,N_863);
nand U3449 (N_3449,N_1133,N_1453);
and U3450 (N_3450,N_1958,N_424);
and U3451 (N_3451,N_140,N_456);
and U3452 (N_3452,N_706,N_1331);
nor U3453 (N_3453,N_854,N_767);
nor U3454 (N_3454,N_1315,N_1946);
or U3455 (N_3455,N_1217,N_990);
xor U3456 (N_3456,N_1074,N_1391);
nor U3457 (N_3457,N_340,N_1422);
nor U3458 (N_3458,N_1735,N_228);
nand U3459 (N_3459,N_382,N_619);
nand U3460 (N_3460,N_309,N_32);
and U3461 (N_3461,N_573,N_1044);
and U3462 (N_3462,N_1193,N_814);
or U3463 (N_3463,N_1195,N_669);
nor U3464 (N_3464,N_491,N_103);
and U3465 (N_3465,N_1857,N_147);
nor U3466 (N_3466,N_49,N_338);
or U3467 (N_3467,N_903,N_1712);
nand U3468 (N_3468,N_1009,N_134);
and U3469 (N_3469,N_847,N_719);
nand U3470 (N_3470,N_1140,N_1409);
and U3471 (N_3471,N_1648,N_233);
and U3472 (N_3472,N_1194,N_1671);
nor U3473 (N_3473,N_1763,N_887);
and U3474 (N_3474,N_1114,N_1894);
nand U3475 (N_3475,N_1221,N_479);
nor U3476 (N_3476,N_134,N_1781);
or U3477 (N_3477,N_1127,N_1833);
and U3478 (N_3478,N_1978,N_37);
nor U3479 (N_3479,N_1894,N_501);
nor U3480 (N_3480,N_525,N_1994);
nand U3481 (N_3481,N_1433,N_1639);
and U3482 (N_3482,N_448,N_1807);
nand U3483 (N_3483,N_1381,N_1726);
nand U3484 (N_3484,N_511,N_1472);
and U3485 (N_3485,N_884,N_1694);
nand U3486 (N_3486,N_1161,N_1098);
or U3487 (N_3487,N_25,N_1020);
nand U3488 (N_3488,N_1677,N_314);
and U3489 (N_3489,N_1760,N_859);
and U3490 (N_3490,N_1362,N_114);
and U3491 (N_3491,N_627,N_541);
nand U3492 (N_3492,N_1064,N_1344);
or U3493 (N_3493,N_425,N_613);
or U3494 (N_3494,N_1230,N_965);
nor U3495 (N_3495,N_77,N_921);
nand U3496 (N_3496,N_1015,N_284);
and U3497 (N_3497,N_952,N_957);
xnor U3498 (N_3498,N_272,N_1111);
nand U3499 (N_3499,N_1222,N_1235);
nor U3500 (N_3500,N_1649,N_525);
and U3501 (N_3501,N_154,N_1913);
nor U3502 (N_3502,N_535,N_1727);
nand U3503 (N_3503,N_233,N_1695);
nand U3504 (N_3504,N_500,N_242);
and U3505 (N_3505,N_1031,N_1195);
nor U3506 (N_3506,N_502,N_1348);
nor U3507 (N_3507,N_1924,N_1523);
nor U3508 (N_3508,N_689,N_944);
nand U3509 (N_3509,N_228,N_1587);
nor U3510 (N_3510,N_788,N_1409);
or U3511 (N_3511,N_141,N_1061);
nor U3512 (N_3512,N_980,N_89);
nor U3513 (N_3513,N_1459,N_1264);
nand U3514 (N_3514,N_1072,N_1168);
and U3515 (N_3515,N_1186,N_120);
nand U3516 (N_3516,N_1840,N_407);
or U3517 (N_3517,N_1019,N_1474);
or U3518 (N_3518,N_1481,N_1658);
nor U3519 (N_3519,N_718,N_66);
nand U3520 (N_3520,N_646,N_1756);
nand U3521 (N_3521,N_1306,N_1657);
and U3522 (N_3522,N_757,N_1153);
and U3523 (N_3523,N_100,N_793);
and U3524 (N_3524,N_140,N_703);
and U3525 (N_3525,N_997,N_689);
and U3526 (N_3526,N_30,N_811);
nand U3527 (N_3527,N_808,N_1691);
nor U3528 (N_3528,N_714,N_496);
or U3529 (N_3529,N_1059,N_1798);
nor U3530 (N_3530,N_1149,N_570);
and U3531 (N_3531,N_63,N_650);
xnor U3532 (N_3532,N_842,N_825);
or U3533 (N_3533,N_402,N_1800);
xnor U3534 (N_3534,N_1817,N_650);
nand U3535 (N_3535,N_72,N_1050);
nand U3536 (N_3536,N_508,N_734);
nor U3537 (N_3537,N_1933,N_1757);
or U3538 (N_3538,N_1595,N_861);
or U3539 (N_3539,N_1579,N_395);
or U3540 (N_3540,N_280,N_1826);
and U3541 (N_3541,N_1412,N_1637);
nor U3542 (N_3542,N_133,N_1666);
or U3543 (N_3543,N_1462,N_294);
xnor U3544 (N_3544,N_1433,N_1895);
and U3545 (N_3545,N_390,N_1844);
or U3546 (N_3546,N_738,N_20);
nand U3547 (N_3547,N_1848,N_1962);
or U3548 (N_3548,N_1072,N_1091);
nand U3549 (N_3549,N_1890,N_1295);
nand U3550 (N_3550,N_638,N_234);
nor U3551 (N_3551,N_1667,N_720);
nor U3552 (N_3552,N_1724,N_559);
nor U3553 (N_3553,N_753,N_1147);
or U3554 (N_3554,N_43,N_1645);
nand U3555 (N_3555,N_675,N_1398);
or U3556 (N_3556,N_813,N_607);
or U3557 (N_3557,N_1615,N_1005);
nand U3558 (N_3558,N_368,N_1480);
nor U3559 (N_3559,N_1689,N_451);
nand U3560 (N_3560,N_1088,N_307);
nand U3561 (N_3561,N_1249,N_1773);
and U3562 (N_3562,N_997,N_768);
and U3563 (N_3563,N_1256,N_1833);
nand U3564 (N_3564,N_537,N_1391);
nand U3565 (N_3565,N_392,N_958);
nand U3566 (N_3566,N_1059,N_1866);
nand U3567 (N_3567,N_823,N_1868);
nor U3568 (N_3568,N_1305,N_1751);
nand U3569 (N_3569,N_1427,N_1330);
and U3570 (N_3570,N_623,N_1570);
and U3571 (N_3571,N_44,N_1551);
nor U3572 (N_3572,N_1554,N_853);
nor U3573 (N_3573,N_683,N_368);
and U3574 (N_3574,N_641,N_374);
nor U3575 (N_3575,N_1493,N_693);
nor U3576 (N_3576,N_166,N_1454);
or U3577 (N_3577,N_1588,N_767);
or U3578 (N_3578,N_670,N_1056);
nor U3579 (N_3579,N_1191,N_309);
nor U3580 (N_3580,N_409,N_1635);
or U3581 (N_3581,N_768,N_82);
or U3582 (N_3582,N_647,N_1992);
nand U3583 (N_3583,N_1132,N_799);
xor U3584 (N_3584,N_1792,N_200);
and U3585 (N_3585,N_521,N_99);
or U3586 (N_3586,N_1787,N_669);
or U3587 (N_3587,N_560,N_1984);
and U3588 (N_3588,N_1819,N_495);
nand U3589 (N_3589,N_806,N_998);
nor U3590 (N_3590,N_691,N_1959);
nor U3591 (N_3591,N_432,N_1577);
nand U3592 (N_3592,N_1023,N_1257);
or U3593 (N_3593,N_592,N_1714);
or U3594 (N_3594,N_599,N_1304);
nor U3595 (N_3595,N_599,N_534);
nor U3596 (N_3596,N_855,N_1847);
nand U3597 (N_3597,N_383,N_775);
or U3598 (N_3598,N_286,N_1517);
and U3599 (N_3599,N_828,N_1788);
and U3600 (N_3600,N_1015,N_1830);
nand U3601 (N_3601,N_1669,N_1735);
nor U3602 (N_3602,N_737,N_1027);
and U3603 (N_3603,N_1561,N_1646);
or U3604 (N_3604,N_398,N_1404);
and U3605 (N_3605,N_1143,N_980);
and U3606 (N_3606,N_822,N_219);
or U3607 (N_3607,N_1304,N_1467);
nor U3608 (N_3608,N_750,N_1612);
nor U3609 (N_3609,N_109,N_53);
and U3610 (N_3610,N_1819,N_1493);
or U3611 (N_3611,N_300,N_1466);
and U3612 (N_3612,N_52,N_112);
nor U3613 (N_3613,N_246,N_1055);
and U3614 (N_3614,N_539,N_1827);
nand U3615 (N_3615,N_1102,N_648);
nand U3616 (N_3616,N_320,N_117);
and U3617 (N_3617,N_1861,N_1530);
or U3618 (N_3618,N_1928,N_619);
or U3619 (N_3619,N_891,N_1255);
nor U3620 (N_3620,N_1162,N_1338);
or U3621 (N_3621,N_121,N_351);
and U3622 (N_3622,N_1615,N_743);
or U3623 (N_3623,N_466,N_726);
or U3624 (N_3624,N_418,N_318);
nand U3625 (N_3625,N_1180,N_1167);
and U3626 (N_3626,N_733,N_487);
or U3627 (N_3627,N_1442,N_369);
and U3628 (N_3628,N_1131,N_630);
nor U3629 (N_3629,N_1253,N_1004);
and U3630 (N_3630,N_37,N_769);
or U3631 (N_3631,N_53,N_1490);
or U3632 (N_3632,N_1837,N_57);
or U3633 (N_3633,N_244,N_1178);
nand U3634 (N_3634,N_878,N_1702);
nand U3635 (N_3635,N_184,N_60);
nor U3636 (N_3636,N_177,N_3);
or U3637 (N_3637,N_542,N_516);
or U3638 (N_3638,N_1926,N_715);
nor U3639 (N_3639,N_39,N_568);
nor U3640 (N_3640,N_1931,N_856);
nor U3641 (N_3641,N_1691,N_848);
and U3642 (N_3642,N_696,N_825);
nor U3643 (N_3643,N_1698,N_1827);
and U3644 (N_3644,N_1809,N_816);
or U3645 (N_3645,N_141,N_708);
or U3646 (N_3646,N_1877,N_394);
nor U3647 (N_3647,N_1750,N_2);
xor U3648 (N_3648,N_633,N_1313);
nor U3649 (N_3649,N_128,N_1809);
nor U3650 (N_3650,N_784,N_911);
or U3651 (N_3651,N_409,N_1118);
nand U3652 (N_3652,N_1664,N_1805);
and U3653 (N_3653,N_1700,N_438);
nor U3654 (N_3654,N_1382,N_799);
and U3655 (N_3655,N_628,N_1654);
nor U3656 (N_3656,N_865,N_66);
or U3657 (N_3657,N_1604,N_244);
nor U3658 (N_3658,N_1817,N_1055);
xor U3659 (N_3659,N_880,N_627);
or U3660 (N_3660,N_53,N_1829);
or U3661 (N_3661,N_939,N_1327);
nand U3662 (N_3662,N_1408,N_1414);
nor U3663 (N_3663,N_460,N_407);
or U3664 (N_3664,N_1694,N_1161);
nor U3665 (N_3665,N_59,N_1873);
and U3666 (N_3666,N_331,N_1398);
xor U3667 (N_3667,N_1856,N_1920);
or U3668 (N_3668,N_785,N_1092);
or U3669 (N_3669,N_1679,N_1971);
and U3670 (N_3670,N_289,N_315);
and U3671 (N_3671,N_1778,N_503);
nand U3672 (N_3672,N_1590,N_951);
xnor U3673 (N_3673,N_59,N_364);
nor U3674 (N_3674,N_1287,N_501);
nand U3675 (N_3675,N_1537,N_167);
or U3676 (N_3676,N_1423,N_1226);
and U3677 (N_3677,N_661,N_517);
nand U3678 (N_3678,N_1016,N_1439);
or U3679 (N_3679,N_677,N_1767);
and U3680 (N_3680,N_309,N_831);
or U3681 (N_3681,N_396,N_1379);
nand U3682 (N_3682,N_313,N_256);
or U3683 (N_3683,N_1600,N_190);
and U3684 (N_3684,N_1643,N_500);
nor U3685 (N_3685,N_531,N_235);
or U3686 (N_3686,N_1198,N_1708);
nand U3687 (N_3687,N_806,N_394);
or U3688 (N_3688,N_763,N_807);
nand U3689 (N_3689,N_984,N_1021);
xnor U3690 (N_3690,N_703,N_1556);
nand U3691 (N_3691,N_1090,N_1842);
and U3692 (N_3692,N_1587,N_587);
and U3693 (N_3693,N_970,N_776);
nand U3694 (N_3694,N_163,N_1115);
and U3695 (N_3695,N_1243,N_788);
nand U3696 (N_3696,N_1587,N_596);
and U3697 (N_3697,N_1065,N_725);
nor U3698 (N_3698,N_462,N_1067);
or U3699 (N_3699,N_577,N_1568);
nor U3700 (N_3700,N_1673,N_1125);
nand U3701 (N_3701,N_273,N_526);
or U3702 (N_3702,N_1656,N_1320);
and U3703 (N_3703,N_508,N_424);
and U3704 (N_3704,N_1918,N_1072);
or U3705 (N_3705,N_293,N_1848);
and U3706 (N_3706,N_85,N_0);
nor U3707 (N_3707,N_1854,N_1176);
and U3708 (N_3708,N_1555,N_1086);
and U3709 (N_3709,N_550,N_1187);
nand U3710 (N_3710,N_1197,N_1116);
xor U3711 (N_3711,N_779,N_91);
nand U3712 (N_3712,N_1800,N_242);
or U3713 (N_3713,N_1126,N_1911);
and U3714 (N_3714,N_1538,N_612);
nor U3715 (N_3715,N_792,N_848);
nor U3716 (N_3716,N_961,N_1293);
or U3717 (N_3717,N_1801,N_255);
or U3718 (N_3718,N_1338,N_1557);
nand U3719 (N_3719,N_952,N_534);
nand U3720 (N_3720,N_1972,N_253);
nor U3721 (N_3721,N_1525,N_77);
xor U3722 (N_3722,N_601,N_557);
nand U3723 (N_3723,N_383,N_1258);
nor U3724 (N_3724,N_1971,N_742);
nor U3725 (N_3725,N_1807,N_1703);
and U3726 (N_3726,N_1454,N_383);
or U3727 (N_3727,N_1693,N_906);
nor U3728 (N_3728,N_1347,N_421);
and U3729 (N_3729,N_455,N_866);
nand U3730 (N_3730,N_51,N_671);
nand U3731 (N_3731,N_1723,N_1019);
nor U3732 (N_3732,N_1685,N_869);
and U3733 (N_3733,N_322,N_1186);
nor U3734 (N_3734,N_1652,N_1576);
xnor U3735 (N_3735,N_259,N_1872);
nor U3736 (N_3736,N_1981,N_374);
nand U3737 (N_3737,N_515,N_1771);
or U3738 (N_3738,N_353,N_53);
nor U3739 (N_3739,N_1762,N_1776);
nor U3740 (N_3740,N_1920,N_1268);
or U3741 (N_3741,N_655,N_477);
nor U3742 (N_3742,N_835,N_1828);
nand U3743 (N_3743,N_180,N_724);
nor U3744 (N_3744,N_289,N_461);
or U3745 (N_3745,N_1845,N_76);
or U3746 (N_3746,N_1065,N_1351);
and U3747 (N_3747,N_164,N_551);
xnor U3748 (N_3748,N_1174,N_1100);
nor U3749 (N_3749,N_1645,N_1445);
or U3750 (N_3750,N_1199,N_604);
or U3751 (N_3751,N_30,N_290);
nor U3752 (N_3752,N_1965,N_1637);
nor U3753 (N_3753,N_1465,N_507);
nand U3754 (N_3754,N_180,N_709);
and U3755 (N_3755,N_1802,N_1486);
nand U3756 (N_3756,N_1690,N_1414);
nand U3757 (N_3757,N_1071,N_1370);
nor U3758 (N_3758,N_1476,N_184);
or U3759 (N_3759,N_1478,N_265);
or U3760 (N_3760,N_1630,N_710);
or U3761 (N_3761,N_419,N_758);
or U3762 (N_3762,N_964,N_815);
nor U3763 (N_3763,N_518,N_45);
or U3764 (N_3764,N_1457,N_808);
and U3765 (N_3765,N_319,N_1494);
and U3766 (N_3766,N_1181,N_89);
or U3767 (N_3767,N_515,N_1897);
nor U3768 (N_3768,N_1947,N_1943);
nor U3769 (N_3769,N_326,N_1229);
and U3770 (N_3770,N_1584,N_1519);
nand U3771 (N_3771,N_371,N_1355);
nor U3772 (N_3772,N_700,N_667);
nor U3773 (N_3773,N_289,N_1473);
nand U3774 (N_3774,N_68,N_475);
nor U3775 (N_3775,N_1157,N_244);
nand U3776 (N_3776,N_1047,N_1212);
or U3777 (N_3777,N_555,N_671);
or U3778 (N_3778,N_1289,N_469);
and U3779 (N_3779,N_1753,N_287);
nand U3780 (N_3780,N_373,N_496);
nor U3781 (N_3781,N_1214,N_1729);
and U3782 (N_3782,N_1971,N_854);
or U3783 (N_3783,N_1189,N_538);
nor U3784 (N_3784,N_302,N_177);
nor U3785 (N_3785,N_378,N_818);
and U3786 (N_3786,N_1971,N_1081);
nand U3787 (N_3787,N_1445,N_919);
nor U3788 (N_3788,N_1376,N_1362);
nor U3789 (N_3789,N_1866,N_1929);
nand U3790 (N_3790,N_1952,N_1394);
nand U3791 (N_3791,N_889,N_912);
nand U3792 (N_3792,N_1361,N_1787);
nand U3793 (N_3793,N_1572,N_1916);
nand U3794 (N_3794,N_1504,N_1629);
or U3795 (N_3795,N_1182,N_1347);
nand U3796 (N_3796,N_623,N_82);
nand U3797 (N_3797,N_1065,N_1534);
nand U3798 (N_3798,N_1335,N_1593);
nand U3799 (N_3799,N_1866,N_792);
or U3800 (N_3800,N_215,N_1257);
or U3801 (N_3801,N_342,N_1407);
nand U3802 (N_3802,N_19,N_575);
nand U3803 (N_3803,N_1364,N_1482);
and U3804 (N_3804,N_5,N_1148);
or U3805 (N_3805,N_1383,N_595);
nand U3806 (N_3806,N_1212,N_697);
nor U3807 (N_3807,N_224,N_1703);
and U3808 (N_3808,N_542,N_336);
nor U3809 (N_3809,N_199,N_21);
and U3810 (N_3810,N_1459,N_1017);
nand U3811 (N_3811,N_1818,N_579);
nand U3812 (N_3812,N_1031,N_895);
nor U3813 (N_3813,N_947,N_623);
or U3814 (N_3814,N_40,N_765);
and U3815 (N_3815,N_915,N_1533);
and U3816 (N_3816,N_590,N_1319);
xnor U3817 (N_3817,N_1624,N_1342);
and U3818 (N_3818,N_1545,N_1910);
xor U3819 (N_3819,N_145,N_1556);
nand U3820 (N_3820,N_1850,N_1337);
nand U3821 (N_3821,N_1118,N_1534);
and U3822 (N_3822,N_1307,N_106);
nand U3823 (N_3823,N_851,N_750);
nand U3824 (N_3824,N_758,N_1594);
nor U3825 (N_3825,N_1774,N_1707);
nor U3826 (N_3826,N_188,N_1641);
or U3827 (N_3827,N_1942,N_819);
or U3828 (N_3828,N_1634,N_678);
nor U3829 (N_3829,N_1873,N_1791);
nor U3830 (N_3830,N_220,N_1564);
and U3831 (N_3831,N_887,N_1265);
nand U3832 (N_3832,N_1191,N_1842);
and U3833 (N_3833,N_1349,N_722);
and U3834 (N_3834,N_1230,N_1557);
nor U3835 (N_3835,N_466,N_598);
or U3836 (N_3836,N_1596,N_1370);
or U3837 (N_3837,N_1130,N_1688);
or U3838 (N_3838,N_1033,N_1585);
or U3839 (N_3839,N_851,N_1034);
nor U3840 (N_3840,N_921,N_870);
or U3841 (N_3841,N_261,N_537);
nor U3842 (N_3842,N_288,N_813);
nand U3843 (N_3843,N_279,N_953);
nand U3844 (N_3844,N_744,N_1655);
nor U3845 (N_3845,N_1599,N_1207);
and U3846 (N_3846,N_961,N_1922);
nor U3847 (N_3847,N_699,N_1433);
nor U3848 (N_3848,N_675,N_492);
nand U3849 (N_3849,N_1360,N_1024);
or U3850 (N_3850,N_898,N_1187);
nand U3851 (N_3851,N_897,N_16);
or U3852 (N_3852,N_1711,N_842);
nor U3853 (N_3853,N_209,N_1600);
nor U3854 (N_3854,N_482,N_860);
or U3855 (N_3855,N_108,N_741);
nand U3856 (N_3856,N_789,N_587);
or U3857 (N_3857,N_367,N_395);
and U3858 (N_3858,N_1558,N_1237);
nor U3859 (N_3859,N_590,N_226);
nor U3860 (N_3860,N_664,N_1767);
or U3861 (N_3861,N_1167,N_427);
nor U3862 (N_3862,N_1177,N_411);
or U3863 (N_3863,N_1134,N_1673);
and U3864 (N_3864,N_1702,N_1436);
or U3865 (N_3865,N_419,N_1950);
nand U3866 (N_3866,N_445,N_702);
or U3867 (N_3867,N_397,N_1132);
xor U3868 (N_3868,N_919,N_1846);
or U3869 (N_3869,N_1543,N_1311);
and U3870 (N_3870,N_1845,N_115);
and U3871 (N_3871,N_621,N_1851);
nand U3872 (N_3872,N_1475,N_1765);
nand U3873 (N_3873,N_526,N_1465);
nor U3874 (N_3874,N_166,N_737);
nand U3875 (N_3875,N_1916,N_1273);
and U3876 (N_3876,N_574,N_767);
nand U3877 (N_3877,N_1915,N_1549);
or U3878 (N_3878,N_940,N_1200);
nor U3879 (N_3879,N_128,N_1674);
or U3880 (N_3880,N_614,N_1274);
nor U3881 (N_3881,N_37,N_302);
nor U3882 (N_3882,N_1600,N_1817);
nor U3883 (N_3883,N_1101,N_1211);
and U3884 (N_3884,N_1705,N_1304);
or U3885 (N_3885,N_239,N_1947);
and U3886 (N_3886,N_49,N_1751);
or U3887 (N_3887,N_464,N_915);
xnor U3888 (N_3888,N_1989,N_977);
and U3889 (N_3889,N_1834,N_930);
nand U3890 (N_3890,N_876,N_1214);
nor U3891 (N_3891,N_454,N_1099);
nand U3892 (N_3892,N_721,N_466);
nand U3893 (N_3893,N_1220,N_145);
and U3894 (N_3894,N_1251,N_367);
nand U3895 (N_3895,N_73,N_355);
nand U3896 (N_3896,N_492,N_1053);
or U3897 (N_3897,N_795,N_364);
nor U3898 (N_3898,N_1629,N_1077);
or U3899 (N_3899,N_632,N_1178);
nand U3900 (N_3900,N_1833,N_198);
nand U3901 (N_3901,N_398,N_561);
and U3902 (N_3902,N_352,N_1856);
or U3903 (N_3903,N_1581,N_852);
xnor U3904 (N_3904,N_1776,N_1459);
nor U3905 (N_3905,N_1608,N_498);
or U3906 (N_3906,N_1184,N_19);
nand U3907 (N_3907,N_473,N_422);
nor U3908 (N_3908,N_659,N_771);
and U3909 (N_3909,N_1721,N_964);
xor U3910 (N_3910,N_1598,N_1590);
nand U3911 (N_3911,N_1806,N_1199);
or U3912 (N_3912,N_1949,N_221);
nand U3913 (N_3913,N_1943,N_1505);
or U3914 (N_3914,N_1328,N_552);
nand U3915 (N_3915,N_1930,N_1985);
or U3916 (N_3916,N_1902,N_327);
nor U3917 (N_3917,N_1469,N_1792);
nand U3918 (N_3918,N_1393,N_1483);
and U3919 (N_3919,N_156,N_928);
nor U3920 (N_3920,N_350,N_225);
nor U3921 (N_3921,N_1001,N_514);
or U3922 (N_3922,N_1381,N_902);
or U3923 (N_3923,N_936,N_1772);
or U3924 (N_3924,N_1715,N_139);
or U3925 (N_3925,N_663,N_1295);
and U3926 (N_3926,N_60,N_1571);
xnor U3927 (N_3927,N_1980,N_1258);
and U3928 (N_3928,N_864,N_939);
and U3929 (N_3929,N_1965,N_1065);
or U3930 (N_3930,N_1413,N_1407);
nand U3931 (N_3931,N_795,N_393);
or U3932 (N_3932,N_1732,N_398);
and U3933 (N_3933,N_1789,N_1667);
xor U3934 (N_3934,N_1098,N_210);
nor U3935 (N_3935,N_1842,N_33);
nand U3936 (N_3936,N_1077,N_228);
nor U3937 (N_3937,N_321,N_1603);
and U3938 (N_3938,N_695,N_86);
and U3939 (N_3939,N_68,N_1960);
nor U3940 (N_3940,N_999,N_417);
nand U3941 (N_3941,N_957,N_1345);
nand U3942 (N_3942,N_1704,N_954);
nand U3943 (N_3943,N_686,N_717);
nand U3944 (N_3944,N_1323,N_193);
or U3945 (N_3945,N_1635,N_786);
and U3946 (N_3946,N_1832,N_944);
nand U3947 (N_3947,N_407,N_1887);
or U3948 (N_3948,N_857,N_823);
or U3949 (N_3949,N_93,N_186);
and U3950 (N_3950,N_1231,N_740);
or U3951 (N_3951,N_1153,N_1030);
nand U3952 (N_3952,N_1046,N_1914);
or U3953 (N_3953,N_591,N_697);
or U3954 (N_3954,N_1025,N_76);
or U3955 (N_3955,N_18,N_986);
and U3956 (N_3956,N_1437,N_304);
nand U3957 (N_3957,N_706,N_412);
nor U3958 (N_3958,N_1651,N_1684);
nand U3959 (N_3959,N_441,N_313);
or U3960 (N_3960,N_1310,N_1169);
nand U3961 (N_3961,N_1024,N_993);
and U3962 (N_3962,N_360,N_1223);
or U3963 (N_3963,N_278,N_1469);
nor U3964 (N_3964,N_177,N_1214);
and U3965 (N_3965,N_1971,N_760);
and U3966 (N_3966,N_1858,N_682);
nand U3967 (N_3967,N_1272,N_76);
nand U3968 (N_3968,N_25,N_1643);
nand U3969 (N_3969,N_1084,N_1688);
or U3970 (N_3970,N_509,N_1375);
nand U3971 (N_3971,N_1152,N_456);
nor U3972 (N_3972,N_1622,N_1830);
nor U3973 (N_3973,N_1293,N_835);
and U3974 (N_3974,N_1542,N_628);
nand U3975 (N_3975,N_1272,N_1747);
and U3976 (N_3976,N_1228,N_279);
or U3977 (N_3977,N_481,N_358);
and U3978 (N_3978,N_150,N_1630);
nor U3979 (N_3979,N_606,N_237);
nand U3980 (N_3980,N_1372,N_591);
nor U3981 (N_3981,N_1708,N_1150);
nand U3982 (N_3982,N_122,N_1947);
nand U3983 (N_3983,N_391,N_805);
nor U3984 (N_3984,N_1096,N_729);
and U3985 (N_3985,N_583,N_687);
nand U3986 (N_3986,N_488,N_1592);
nand U3987 (N_3987,N_601,N_673);
nand U3988 (N_3988,N_461,N_1293);
nand U3989 (N_3989,N_1642,N_716);
nor U3990 (N_3990,N_516,N_56);
or U3991 (N_3991,N_1909,N_1784);
nand U3992 (N_3992,N_1910,N_864);
nor U3993 (N_3993,N_1005,N_497);
xor U3994 (N_3994,N_1440,N_1329);
nor U3995 (N_3995,N_1524,N_1093);
or U3996 (N_3996,N_689,N_661);
or U3997 (N_3997,N_1970,N_286);
nand U3998 (N_3998,N_1814,N_1089);
or U3999 (N_3999,N_1630,N_825);
nand U4000 (N_4000,N_2698,N_3776);
and U4001 (N_4001,N_3238,N_2472);
nand U4002 (N_4002,N_2893,N_2358);
nand U4003 (N_4003,N_2627,N_3895);
nor U4004 (N_4004,N_3837,N_2444);
nor U4005 (N_4005,N_2142,N_3102);
nand U4006 (N_4006,N_3143,N_3642);
nand U4007 (N_4007,N_3487,N_3987);
nor U4008 (N_4008,N_2239,N_3902);
nor U4009 (N_4009,N_2240,N_2006);
or U4010 (N_4010,N_3964,N_3896);
nand U4011 (N_4011,N_2703,N_2987);
or U4012 (N_4012,N_2648,N_2201);
nand U4013 (N_4013,N_2646,N_2799);
and U4014 (N_4014,N_3121,N_3971);
and U4015 (N_4015,N_3009,N_2876);
nor U4016 (N_4016,N_2496,N_3353);
nand U4017 (N_4017,N_2293,N_3537);
and U4018 (N_4018,N_2013,N_3655);
nand U4019 (N_4019,N_2965,N_2680);
or U4020 (N_4020,N_3171,N_3311);
nand U4021 (N_4021,N_3893,N_2125);
and U4022 (N_4022,N_2165,N_2296);
or U4023 (N_4023,N_3578,N_3381);
or U4024 (N_4024,N_3147,N_2722);
nor U4025 (N_4025,N_2523,N_3141);
and U4026 (N_4026,N_2575,N_2489);
nand U4027 (N_4027,N_3799,N_2018);
and U4028 (N_4028,N_3069,N_3038);
or U4029 (N_4029,N_2728,N_2994);
nor U4030 (N_4030,N_3188,N_2830);
nand U4031 (N_4031,N_2288,N_2289);
or U4032 (N_4032,N_3013,N_3476);
and U4033 (N_4033,N_2481,N_3074);
or U4034 (N_4034,N_2363,N_2498);
or U4035 (N_4035,N_2669,N_3425);
xor U4036 (N_4036,N_2063,N_2615);
or U4037 (N_4037,N_3145,N_2137);
or U4038 (N_4038,N_2280,N_2075);
nand U4039 (N_4039,N_2490,N_2268);
nand U4040 (N_4040,N_2393,N_3260);
nor U4041 (N_4041,N_2053,N_2727);
and U4042 (N_4042,N_2607,N_2145);
nand U4043 (N_4043,N_3870,N_3072);
nor U4044 (N_4044,N_3990,N_2902);
and U4045 (N_4045,N_3054,N_2353);
or U4046 (N_4046,N_2130,N_3667);
and U4047 (N_4047,N_2894,N_2598);
nand U4048 (N_4048,N_2959,N_2046);
nor U4049 (N_4049,N_2157,N_3111);
nand U4050 (N_4050,N_3394,N_3498);
nor U4051 (N_4051,N_2072,N_3191);
or U4052 (N_4052,N_2205,N_3092);
nand U4053 (N_4053,N_2820,N_3917);
or U4054 (N_4054,N_3478,N_2433);
nor U4055 (N_4055,N_2847,N_2022);
and U4056 (N_4056,N_2789,N_2525);
nand U4057 (N_4057,N_2333,N_3692);
and U4058 (N_4058,N_2313,N_2181);
nand U4059 (N_4059,N_3854,N_3649);
or U4060 (N_4060,N_3749,N_3753);
and U4061 (N_4061,N_3900,N_3445);
nand U4062 (N_4062,N_2981,N_3631);
xnor U4063 (N_4063,N_3670,N_3572);
nor U4064 (N_4064,N_2792,N_2485);
and U4065 (N_4065,N_2687,N_3493);
nor U4066 (N_4066,N_2582,N_2086);
xor U4067 (N_4067,N_2527,N_3265);
nand U4068 (N_4068,N_3391,N_3177);
or U4069 (N_4069,N_3120,N_3993);
nor U4070 (N_4070,N_2016,N_3582);
or U4071 (N_4071,N_2635,N_3880);
and U4072 (N_4072,N_3082,N_3182);
nor U4073 (N_4073,N_3660,N_3587);
or U4074 (N_4074,N_2070,N_3291);
nor U4075 (N_4075,N_2911,N_3939);
nor U4076 (N_4076,N_3978,N_2983);
nand U4077 (N_4077,N_2609,N_3563);
or U4078 (N_4078,N_3404,N_2448);
nor U4079 (N_4079,N_3058,N_2032);
nor U4080 (N_4080,N_2816,N_3833);
nor U4081 (N_4081,N_3746,N_3328);
and U4082 (N_4082,N_2973,N_2369);
or U4083 (N_4083,N_2144,N_2291);
nand U4084 (N_4084,N_2504,N_2860);
nor U4085 (N_4085,N_3108,N_2715);
nor U4086 (N_4086,N_3152,N_3702);
nand U4087 (N_4087,N_3161,N_3383);
or U4088 (N_4088,N_2019,N_2478);
nor U4089 (N_4089,N_3050,N_3230);
nor U4090 (N_4090,N_3947,N_2991);
nand U4091 (N_4091,N_3458,N_3264);
xnor U4092 (N_4092,N_3714,N_2337);
or U4093 (N_4093,N_3836,N_3122);
nand U4094 (N_4094,N_2865,N_3806);
nor U4095 (N_4095,N_3609,N_3675);
nor U4096 (N_4096,N_3332,N_2743);
nor U4097 (N_4097,N_3247,N_3929);
or U4098 (N_4098,N_3342,N_3178);
and U4099 (N_4099,N_3674,N_2899);
and U4100 (N_4100,N_2350,N_3000);
or U4101 (N_4101,N_3850,N_2770);
or U4102 (N_4102,N_2050,N_2348);
and U4103 (N_4103,N_2397,N_2682);
xnor U4104 (N_4104,N_3056,N_2202);
nand U4105 (N_4105,N_3731,N_3555);
and U4106 (N_4106,N_3873,N_3792);
nor U4107 (N_4107,N_3401,N_2193);
and U4108 (N_4108,N_3010,N_3744);
and U4109 (N_4109,N_2749,N_2331);
or U4110 (N_4110,N_3948,N_3514);
and U4111 (N_4111,N_3403,N_3349);
or U4112 (N_4112,N_3208,N_2888);
and U4113 (N_4113,N_3979,N_3775);
nor U4114 (N_4114,N_3489,N_3912);
and U4115 (N_4115,N_2930,N_2473);
and U4116 (N_4116,N_2735,N_3067);
and U4117 (N_4117,N_2737,N_3008);
nand U4118 (N_4118,N_2631,N_3685);
nor U4119 (N_4119,N_3384,N_3767);
and U4120 (N_4120,N_2681,N_2626);
or U4121 (N_4121,N_3452,N_2361);
nand U4122 (N_4122,N_2804,N_3524);
or U4123 (N_4123,N_2967,N_2778);
or U4124 (N_4124,N_2282,N_3876);
and U4125 (N_4125,N_3310,N_2920);
or U4126 (N_4126,N_2560,N_3765);
nand U4127 (N_4127,N_3626,N_3881);
nor U4128 (N_4128,N_2510,N_2219);
and U4129 (N_4129,N_3913,N_3818);
and U4130 (N_4130,N_3512,N_3925);
nor U4131 (N_4131,N_3550,N_2807);
nand U4132 (N_4132,N_2691,N_3614);
and U4133 (N_4133,N_3859,N_3878);
nand U4134 (N_4134,N_3025,N_2952);
and U4135 (N_4135,N_3337,N_3099);
or U4136 (N_4136,N_3073,N_3831);
nand U4137 (N_4137,N_2080,N_3457);
or U4138 (N_4138,N_3138,N_2442);
and U4139 (N_4139,N_2660,N_3576);
nor U4140 (N_4140,N_2175,N_2622);
and U4141 (N_4141,N_2121,N_3505);
and U4142 (N_4142,N_3322,N_2827);
xor U4143 (N_4143,N_2771,N_2007);
nand U4144 (N_4144,N_3522,N_2301);
and U4145 (N_4145,N_2927,N_2136);
nand U4146 (N_4146,N_2003,N_3999);
nor U4147 (N_4147,N_3421,N_3211);
or U4148 (N_4148,N_2307,N_2755);
and U4149 (N_4149,N_3222,N_2924);
and U4150 (N_4150,N_3981,N_2859);
or U4151 (N_4151,N_3521,N_2047);
and U4152 (N_4152,N_3419,N_2066);
and U4153 (N_4153,N_3237,N_2717);
nand U4154 (N_4154,N_2445,N_3742);
nor U4155 (N_4155,N_2537,N_2354);
and U4156 (N_4156,N_2320,N_3816);
nand U4157 (N_4157,N_3169,N_2197);
or U4158 (N_4158,N_2059,N_3661);
nand U4159 (N_4159,N_2813,N_3543);
nor U4160 (N_4160,N_2535,N_2399);
nand U4161 (N_4161,N_3351,N_3144);
nand U4162 (N_4162,N_3965,N_3723);
xor U4163 (N_4163,N_2336,N_3276);
nand U4164 (N_4164,N_3640,N_3860);
or U4165 (N_4165,N_2094,N_3619);
or U4166 (N_4166,N_2932,N_3068);
and U4167 (N_4167,N_2150,N_2487);
nand U4168 (N_4168,N_3719,N_3579);
and U4169 (N_4169,N_3195,N_2836);
xor U4170 (N_4170,N_2443,N_3710);
nand U4171 (N_4171,N_2324,N_2432);
or U4172 (N_4172,N_2383,N_3345);
or U4173 (N_4173,N_2896,N_3275);
or U4174 (N_4174,N_2795,N_3908);
or U4175 (N_4175,N_2613,N_2664);
nor U4176 (N_4176,N_2095,N_3059);
or U4177 (N_4177,N_2592,N_3185);
or U4178 (N_4178,N_2985,N_3812);
or U4179 (N_4179,N_3199,N_2229);
nor U4180 (N_4180,N_2149,N_3471);
nor U4181 (N_4181,N_3474,N_2848);
nor U4182 (N_4182,N_3807,N_3743);
or U4183 (N_4183,N_2583,N_2449);
or U4184 (N_4184,N_3029,N_2968);
nor U4185 (N_4185,N_3584,N_2367);
or U4186 (N_4186,N_2321,N_3148);
or U4187 (N_4187,N_2076,N_3805);
and U4188 (N_4188,N_3604,N_2111);
nand U4189 (N_4189,N_2849,N_2990);
nor U4190 (N_4190,N_3654,N_2242);
or U4191 (N_4191,N_3671,N_3861);
nor U4192 (N_4192,N_2460,N_3201);
nor U4193 (N_4193,N_2906,N_2707);
or U4194 (N_4194,N_3282,N_3508);
nand U4195 (N_4195,N_2665,N_3110);
and U4196 (N_4196,N_2532,N_3115);
and U4197 (N_4197,N_2312,N_3545);
or U4198 (N_4198,N_3669,N_3216);
and U4199 (N_4199,N_2656,N_3323);
nor U4200 (N_4200,N_3872,N_3826);
nor U4201 (N_4201,N_3440,N_3963);
or U4202 (N_4202,N_2274,N_2343);
or U4203 (N_4203,N_3296,N_2394);
and U4204 (N_4204,N_2103,N_2886);
nor U4205 (N_4205,N_3683,N_2414);
nor U4206 (N_4206,N_3408,N_3162);
nand U4207 (N_4207,N_2087,N_2342);
nor U4208 (N_4208,N_2567,N_3035);
nor U4209 (N_4209,N_2738,N_3104);
nand U4210 (N_4210,N_2261,N_3319);
and U4211 (N_4211,N_3490,N_3789);
nand U4212 (N_4212,N_3766,N_2116);
or U4213 (N_4213,N_3151,N_3610);
or U4214 (N_4214,N_3266,N_3561);
or U4215 (N_4215,N_3300,N_2328);
or U4216 (N_4216,N_2135,N_3361);
or U4217 (N_4217,N_2823,N_2513);
nor U4218 (N_4218,N_2793,N_3858);
nand U4219 (N_4219,N_2765,N_2556);
and U4220 (N_4220,N_3270,N_3730);
nor U4221 (N_4221,N_3814,N_2416);
nor U4222 (N_4222,N_3303,N_2156);
nand U4223 (N_4223,N_2637,N_2387);
or U4224 (N_4224,N_3109,N_2554);
nand U4225 (N_4225,N_3663,N_2247);
nand U4226 (N_4226,N_3580,N_2015);
and U4227 (N_4227,N_2690,N_2419);
and U4228 (N_4228,N_2571,N_2420);
and U4229 (N_4229,N_2199,N_2127);
nand U4230 (N_4230,N_3701,N_3435);
nor U4231 (N_4231,N_3028,N_3468);
and U4232 (N_4232,N_3679,N_3224);
and U4233 (N_4233,N_3616,N_2624);
nor U4234 (N_4234,N_3732,N_2625);
nand U4235 (N_4235,N_2054,N_3290);
and U4236 (N_4236,N_2641,N_3772);
xnor U4237 (N_4237,N_2340,N_2862);
nand U4238 (N_4238,N_2503,N_2235);
or U4239 (N_4239,N_3849,N_2051);
nor U4240 (N_4240,N_2346,N_3063);
or U4241 (N_4241,N_3784,N_2064);
and U4242 (N_4242,N_2905,N_3336);
nand U4243 (N_4243,N_3373,N_3206);
and U4244 (N_4244,N_3758,N_3358);
or U4245 (N_4245,N_3020,N_2226);
and U4246 (N_4246,N_2725,N_3738);
xnor U4247 (N_4247,N_3242,N_2177);
or U4248 (N_4248,N_2225,N_2605);
and U4249 (N_4249,N_3533,N_3463);
nand U4250 (N_4250,N_3856,N_2109);
nor U4251 (N_4251,N_3874,N_3485);
or U4252 (N_4252,N_2082,N_2559);
and U4253 (N_4253,N_3084,N_2421);
and U4254 (N_4254,N_3910,N_2060);
or U4255 (N_4255,N_2269,N_2227);
xnor U4256 (N_4256,N_2833,N_2904);
or U4257 (N_4257,N_3790,N_2106);
and U4258 (N_4258,N_3601,N_2424);
or U4259 (N_4259,N_3871,N_3156);
nand U4260 (N_4260,N_3124,N_3372);
or U4261 (N_4261,N_3711,N_3693);
nor U4262 (N_4262,N_2480,N_2801);
and U4263 (N_4263,N_3538,N_2056);
or U4264 (N_4264,N_2907,N_2946);
nand U4265 (N_4265,N_2612,N_2285);
nor U4266 (N_4266,N_2702,N_2538);
xnor U4267 (N_4267,N_2835,N_3431);
nor U4268 (N_4268,N_2146,N_2376);
or U4269 (N_4269,N_2601,N_3262);
and U4270 (N_4270,N_2689,N_2325);
nor U4271 (N_4271,N_3748,N_2871);
nor U4272 (N_4272,N_2295,N_2775);
nor U4273 (N_4273,N_3131,N_2079);
nor U4274 (N_4274,N_3426,N_3308);
xnor U4275 (N_4275,N_3348,N_3956);
and U4276 (N_4276,N_3221,N_3518);
and U4277 (N_4277,N_3479,N_3664);
nand U4278 (N_4278,N_3477,N_3941);
xnor U4279 (N_4279,N_2132,N_2566);
nand U4280 (N_4280,N_3497,N_3243);
nor U4281 (N_4281,N_3657,N_3223);
nand U4282 (N_4282,N_2163,N_2852);
or U4283 (N_4283,N_2676,N_2238);
and U4284 (N_4284,N_2417,N_3439);
and U4285 (N_4285,N_3396,N_2644);
nor U4286 (N_4286,N_3924,N_2492);
or U4287 (N_4287,N_3571,N_3321);
or U4288 (N_4288,N_2814,N_2761);
or U4289 (N_4289,N_2319,N_2610);
or U4290 (N_4290,N_2469,N_2491);
nor U4291 (N_4291,N_2314,N_3274);
nand U4292 (N_4292,N_3975,N_2391);
nand U4293 (N_4293,N_2275,N_2895);
nor U4294 (N_4294,N_2172,N_3135);
nor U4295 (N_4295,N_3921,N_3170);
nor U4296 (N_4296,N_3509,N_3249);
nand U4297 (N_4297,N_2042,N_3036);
nand U4298 (N_4298,N_3958,N_2953);
nand U4299 (N_4299,N_2948,N_2372);
nand U4300 (N_4300,N_2774,N_2956);
and U4301 (N_4301,N_3718,N_3811);
and U4302 (N_4302,N_3491,N_3954);
and U4303 (N_4303,N_3053,N_2962);
nand U4304 (N_4304,N_3644,N_3039);
or U4305 (N_4305,N_2740,N_2458);
or U4306 (N_4306,N_2550,N_2547);
nor U4307 (N_4307,N_2365,N_3184);
nand U4308 (N_4308,N_3150,N_2476);
nand U4309 (N_4309,N_3196,N_2021);
or U4310 (N_4310,N_2237,N_2746);
or U4311 (N_4311,N_2263,N_2159);
nand U4312 (N_4312,N_3694,N_3153);
or U4313 (N_4313,N_2884,N_3339);
or U4314 (N_4314,N_2450,N_2029);
nand U4315 (N_4315,N_2705,N_3139);
nand U4316 (N_4316,N_3297,N_2944);
and U4317 (N_4317,N_3622,N_3842);
or U4318 (N_4318,N_3852,N_3155);
nor U4319 (N_4319,N_2655,N_3233);
nand U4320 (N_4320,N_3728,N_3335);
or U4321 (N_4321,N_3133,N_3295);
nand U4322 (N_4322,N_3386,N_3783);
and U4323 (N_4323,N_3919,N_3160);
and U4324 (N_4324,N_3785,N_3472);
or U4325 (N_4325,N_3369,N_2260);
or U4326 (N_4326,N_2283,N_3005);
or U4327 (N_4327,N_3639,N_2744);
or U4328 (N_4328,N_3653,N_2506);
or U4329 (N_4329,N_2180,N_3217);
nor U4330 (N_4330,N_2539,N_2874);
and U4331 (N_4331,N_3447,N_3847);
nor U4332 (N_4332,N_3251,N_3539);
nor U4333 (N_4333,N_2597,N_2477);
and U4334 (N_4334,N_3415,N_3496);
and U4335 (N_4335,N_3080,N_3344);
and U4336 (N_4336,N_3374,N_3095);
nor U4337 (N_4337,N_3729,N_2494);
or U4338 (N_4338,N_2045,N_2658);
and U4339 (N_4339,N_2522,N_2166);
and U4340 (N_4340,N_3562,N_3484);
and U4341 (N_4341,N_3492,N_2067);
or U4342 (N_4342,N_2327,N_2590);
or U4343 (N_4343,N_3354,N_2454);
or U4344 (N_4344,N_3536,N_3988);
nand U4345 (N_4345,N_3090,N_3717);
nor U4346 (N_4346,N_3163,N_3098);
and U4347 (N_4347,N_3959,N_3031);
nand U4348 (N_4348,N_3434,N_3123);
nor U4349 (N_4349,N_2138,N_3112);
or U4350 (N_4350,N_2380,N_3835);
and U4351 (N_4351,N_3280,N_3846);
nand U4352 (N_4352,N_2604,N_2666);
nand U4353 (N_4353,N_3984,N_2182);
or U4354 (N_4354,N_3281,N_3828);
nor U4355 (N_4355,N_3630,N_3957);
nand U4356 (N_4356,N_3455,N_3933);
or U4357 (N_4357,N_2951,N_3596);
or U4358 (N_4358,N_3564,N_3172);
nand U4359 (N_4359,N_2553,N_3051);
and U4360 (N_4360,N_3695,N_2910);
and U4361 (N_4361,N_2357,N_3991);
and U4362 (N_4362,N_3802,N_3441);
and U4363 (N_4363,N_3607,N_3130);
nand U4364 (N_4364,N_2418,N_3643);
nor U4365 (N_4365,N_2360,N_2617);
nor U4366 (N_4366,N_3175,N_3094);
nor U4367 (N_4367,N_3218,N_3909);
nand U4368 (N_4368,N_3226,N_2670);
nand U4369 (N_4369,N_2782,N_2534);
and U4370 (N_4370,N_2008,N_3375);
nand U4371 (N_4371,N_3357,N_2435);
or U4372 (N_4372,N_3613,N_2499);
or U4373 (N_4373,N_3684,N_2389);
nor U4374 (N_4374,N_3840,N_2170);
nand U4375 (N_4375,N_3107,N_3867);
or U4376 (N_4376,N_3911,N_3884);
nand U4377 (N_4377,N_2118,N_2208);
xor U4378 (N_4378,N_2362,N_3313);
nand U4379 (N_4379,N_2084,N_3532);
nand U4380 (N_4380,N_3405,N_3327);
nor U4381 (N_4381,N_3691,N_3119);
or U4382 (N_4382,N_3324,N_2751);
nor U4383 (N_4383,N_2262,N_2993);
nand U4384 (N_4384,N_2196,N_2721);
xor U4385 (N_4385,N_3307,N_2286);
nor U4386 (N_4386,N_2341,N_3089);
nand U4387 (N_4387,N_2908,N_3416);
nand U4388 (N_4388,N_2844,N_2471);
and U4389 (N_4389,N_3168,N_3598);
nor U4390 (N_4390,N_3583,N_3869);
and U4391 (N_4391,N_3034,N_2564);
or U4392 (N_4392,N_2011,N_3590);
nor U4393 (N_4393,N_3727,N_3915);
nand U4394 (N_4394,N_3213,N_2516);
or U4395 (N_4395,N_2733,N_2997);
xor U4396 (N_4396,N_2495,N_2950);
nand U4397 (N_4397,N_2290,N_2468);
nor U4398 (N_4398,N_2384,N_3202);
nand U4399 (N_4399,N_3838,N_2700);
xnor U4400 (N_4400,N_2398,N_3972);
and U4401 (N_4401,N_2565,N_3597);
nor U4402 (N_4402,N_2937,N_2014);
and U4403 (N_4403,N_3889,N_3877);
and U4404 (N_4404,N_2378,N_2359);
or U4405 (N_4405,N_3863,N_3682);
nor U4406 (N_4406,N_2482,N_2633);
nor U4407 (N_4407,N_2147,N_2043);
and U4408 (N_4408,N_2843,N_2171);
and U4409 (N_4409,N_3331,N_2811);
and U4410 (N_4410,N_2031,N_2334);
nand U4411 (N_4411,N_2368,N_2834);
xnor U4412 (N_4412,N_2921,N_2329);
nor U4413 (N_4413,N_2206,N_3707);
xnor U4414 (N_4414,N_2912,N_2570);
and U4415 (N_4415,N_3848,N_3210);
nor U4416 (N_4416,N_3791,N_2992);
or U4417 (N_4417,N_2264,N_3057);
nor U4418 (N_4418,N_2241,N_2732);
nand U4419 (N_4419,N_3239,N_3637);
nor U4420 (N_4420,N_3475,N_2736);
and U4421 (N_4421,N_2922,N_3116);
or U4422 (N_4422,N_2374,N_3207);
nor U4423 (N_4423,N_3501,N_2228);
or U4424 (N_4424,N_3347,N_2839);
nand U4425 (N_4425,N_2758,N_2821);
nand U4426 (N_4426,N_3267,N_2276);
and U4427 (N_4427,N_2892,N_2875);
nand U4428 (N_4428,N_2752,N_3568);
or U4429 (N_4429,N_3427,N_3482);
nand U4430 (N_4430,N_2999,N_2415);
or U4431 (N_4431,N_3822,N_3885);
and U4432 (N_4432,N_2713,N_2585);
xnor U4433 (N_4433,N_2791,N_2568);
or U4434 (N_4434,N_3253,N_3658);
or U4435 (N_4435,N_3605,N_3012);
or U4436 (N_4436,N_2521,N_2940);
nor U4437 (N_4437,N_3469,N_3857);
nand U4438 (N_4438,N_3819,N_2863);
and U4439 (N_4439,N_2542,N_3367);
or U4440 (N_4440,N_3411,N_2438);
and U4441 (N_4441,N_2187,N_3943);
and U4442 (N_4442,N_2697,N_3510);
nand U4443 (N_4443,N_2618,N_3608);
and U4444 (N_4444,N_2270,N_2716);
and U4445 (N_4445,N_2794,N_3892);
or U4446 (N_4446,N_2509,N_3462);
nand U4447 (N_4447,N_3436,N_2284);
or U4448 (N_4448,N_3989,N_3952);
xnor U4449 (N_4449,N_2957,N_3739);
nor U4450 (N_4450,N_2057,N_2654);
or U4451 (N_4451,N_2798,N_3944);
nor U4452 (N_4452,N_2867,N_2379);
nor U4453 (N_4453,N_2796,N_3378);
or U4454 (N_4454,N_3454,N_3759);
and U4455 (N_4455,N_2302,N_3986);
nor U4456 (N_4456,N_2198,N_3879);
nand U4457 (N_4457,N_3528,N_3527);
nor U4458 (N_4458,N_2077,N_3985);
nor U4459 (N_4459,N_3370,N_2528);
nor U4460 (N_4460,N_3777,N_2561);
xnor U4461 (N_4461,N_2139,N_2153);
nand U4462 (N_4462,N_2204,N_3798);
or U4463 (N_4463,N_3645,N_2838);
and U4464 (N_4464,N_3382,N_3966);
nor U4465 (N_4465,N_2955,N_3641);
and U4466 (N_4466,N_2524,N_3395);
or U4467 (N_4467,N_3097,N_3423);
and U4468 (N_4468,N_2686,N_3726);
nand U4469 (N_4469,N_3390,N_2864);
nand U4470 (N_4470,N_2882,N_3190);
and U4471 (N_4471,N_3624,N_2304);
nor U4472 (N_4472,N_2594,N_2479);
or U4473 (N_4473,N_2779,N_2310);
nand U4474 (N_4474,N_3023,N_2577);
and U4475 (N_4475,N_2164,N_2396);
or U4476 (N_4476,N_3517,N_2298);
nor U4477 (N_4477,N_2272,N_2373);
or U4478 (N_4478,N_2299,N_3839);
nor U4479 (N_4479,N_2104,N_2712);
xnor U4480 (N_4480,N_3566,N_3021);
and U4481 (N_4481,N_3735,N_2459);
nand U4482 (N_4482,N_3315,N_3646);
xnor U4483 (N_4483,N_2949,N_3531);
nor U4484 (N_4484,N_3134,N_3618);
nor U4485 (N_4485,N_2230,N_2897);
nor U4486 (N_4486,N_3953,N_2024);
nor U4487 (N_4487,N_3071,N_2335);
and U4488 (N_4488,N_3855,N_3903);
and U4489 (N_4489,N_3551,N_2776);
nand U4490 (N_4490,N_3887,N_2638);
nand U4491 (N_4491,N_3801,N_3453);
xor U4492 (N_4492,N_2085,N_3398);
or U4493 (N_4493,N_3935,N_3793);
nor U4494 (N_4494,N_3540,N_3920);
and U4495 (N_4495,N_3142,N_3376);
and U4496 (N_4496,N_2366,N_3681);
and U4497 (N_4497,N_2787,N_3570);
nand U4498 (N_4498,N_3588,N_2271);
and U4499 (N_4499,N_2388,N_3938);
and U4500 (N_4500,N_2578,N_3166);
nor U4501 (N_4501,N_3060,N_3813);
and U4502 (N_4502,N_2381,N_3236);
and U4503 (N_4503,N_2192,N_2777);
and U4504 (N_4504,N_2579,N_3350);
nor U4505 (N_4505,N_2975,N_2603);
nor U4506 (N_4506,N_2939,N_2195);
nand U4507 (N_4507,N_3554,N_3585);
and U4508 (N_4508,N_3140,N_3033);
and U4509 (N_4509,N_3215,N_2475);
nand U4510 (N_4510,N_3574,N_3968);
and U4511 (N_4511,N_2012,N_3556);
xnor U4512 (N_4512,N_2760,N_3377);
and U4513 (N_4513,N_3136,N_3232);
nor U4514 (N_4514,N_3678,N_2552);
nor U4515 (N_4515,N_2718,N_2675);
and U4516 (N_4516,N_2441,N_3269);
nor U4517 (N_4517,N_3413,N_3715);
and U4518 (N_4518,N_2209,N_2548);
nor U4519 (N_4519,N_3897,N_2212);
nand U4520 (N_4520,N_3385,N_2861);
and U4521 (N_4521,N_2653,N_2339);
nand U4522 (N_4522,N_3794,N_2002);
and U4523 (N_4523,N_2000,N_3076);
nand U4524 (N_4524,N_2898,N_3697);
or U4525 (N_4525,N_3722,N_3334);
and U4526 (N_4526,N_2706,N_2356);
nand U4527 (N_4527,N_2158,N_2315);
or U4528 (N_4528,N_2255,N_2501);
nor U4529 (N_4529,N_3830,N_3901);
and U4530 (N_4530,N_3557,N_3338);
nand U4531 (N_4531,N_2463,N_2591);
and U4532 (N_4532,N_2619,N_3559);
nor U4533 (N_4533,N_3399,N_2243);
nand U4534 (N_4534,N_2245,N_3078);
nand U4535 (N_4535,N_2266,N_3511);
and U4536 (N_4536,N_2426,N_3341);
or U4537 (N_4537,N_3922,N_3875);
or U4538 (N_4538,N_3212,N_2969);
and U4539 (N_4539,N_3737,N_3443);
nand U4540 (N_4540,N_2780,N_2620);
or U4541 (N_4541,N_2858,N_2623);
nand U4542 (N_4542,N_3567,N_3093);
and U4543 (N_4543,N_3768,N_3937);
nand U4544 (N_4544,N_2663,N_2599);
or U4545 (N_4545,N_3397,N_3918);
or U4546 (N_4546,N_2120,N_2117);
nand U4547 (N_4547,N_3293,N_2797);
nand U4548 (N_4548,N_2580,N_2410);
nand U4549 (N_4549,N_3091,N_2058);
or U4550 (N_4550,N_2828,N_2647);
nor U4551 (N_4551,N_3575,N_3634);
or U4552 (N_4552,N_3449,N_2674);
or U4553 (N_4553,N_3248,N_2330);
nor U4554 (N_4554,N_3810,N_2071);
and U4555 (N_4555,N_3360,N_2107);
nor U4556 (N_4556,N_2541,N_2403);
nand U4557 (N_4557,N_2593,N_3259);
nor U4558 (N_4558,N_3200,N_3733);
xnor U4559 (N_4559,N_3229,N_3503);
and U4560 (N_4560,N_3481,N_2141);
and U4561 (N_4561,N_2114,N_3594);
nor U4562 (N_4562,N_3316,N_3278);
and U4563 (N_4563,N_3502,N_3553);
and U4564 (N_4564,N_3523,N_2933);
or U4565 (N_4565,N_2370,N_3302);
and U4566 (N_4566,N_2409,N_3114);
nand U4567 (N_4567,N_2110,N_2035);
nor U4568 (N_4568,N_2105,N_3101);
and U4569 (N_4569,N_3882,N_2996);
nand U4570 (N_4570,N_3287,N_2023);
and U4571 (N_4571,N_2406,N_2434);
nand U4572 (N_4572,N_2526,N_3680);
nand U4573 (N_4573,N_2978,N_2514);
nor U4574 (N_4574,N_3906,N_3309);
nand U4575 (N_4575,N_2694,N_2092);
nand U4576 (N_4576,N_2044,N_2854);
or U4577 (N_4577,N_3343,N_3652);
nor U4578 (N_4578,N_2316,N_3603);
nor U4579 (N_4579,N_2089,N_3055);
and U4580 (N_4580,N_2639,N_2989);
nand U4581 (N_4581,N_2879,N_3393);
nand U4582 (N_4582,N_2128,N_3778);
or U4583 (N_4583,N_3326,N_2634);
or U4584 (N_4584,N_2600,N_3183);
or U4585 (N_4585,N_3894,N_2562);
or U4586 (N_4586,N_2065,N_3928);
and U4587 (N_4587,N_2649,N_2581);
and U4588 (N_4588,N_3832,N_3032);
nand U4589 (N_4589,N_2505,N_2842);
or U4590 (N_4590,N_2588,N_3829);
or U4591 (N_4591,N_2611,N_3030);
and U4592 (N_4592,N_2788,N_2651);
and U4593 (N_4593,N_2630,N_2190);
or U4594 (N_4594,N_2688,N_2033);
or U4595 (N_4595,N_2869,N_3250);
nor U4596 (N_4596,N_3193,N_3209);
xor U4597 (N_4597,N_2711,N_2347);
and U4598 (N_4598,N_2753,N_2464);
or U4599 (N_4599,N_2220,N_2693);
nand U4600 (N_4600,N_2306,N_3227);
nor U4601 (N_4601,N_3362,N_2868);
nand U4602 (N_4602,N_3494,N_2119);
or U4603 (N_4603,N_3480,N_2277);
nor U4604 (N_4604,N_3364,N_3581);
nor U4605 (N_4605,N_3003,N_3659);
and U4606 (N_4606,N_3004,N_3438);
nand U4607 (N_4607,N_2068,N_2083);
nor U4608 (N_4608,N_2456,N_3014);
nand U4609 (N_4609,N_3636,N_3180);
and U4610 (N_4610,N_2451,N_3796);
and U4611 (N_4611,N_3277,N_3506);
and U4612 (N_4612,N_2880,N_2081);
nor U4613 (N_4613,N_3725,N_2576);
nor U4614 (N_4614,N_3542,N_3973);
or U4615 (N_4615,N_2231,N_3252);
nor U4616 (N_4616,N_2739,N_2037);
nor U4617 (N_4617,N_2587,N_2877);
xor U4618 (N_4618,N_3980,N_3930);
or U4619 (N_4619,N_3734,N_3516);
and U4620 (N_4620,N_3591,N_2901);
nand U4621 (N_4621,N_3061,N_3611);
and U4622 (N_4622,N_2377,N_2161);
nand U4623 (N_4623,N_2203,N_2140);
nand U4624 (N_4624,N_2822,N_2160);
or U4625 (N_4625,N_2520,N_3432);
or U4626 (N_4626,N_3617,N_2439);
and U4627 (N_4627,N_3235,N_2850);
or U4628 (N_4628,N_2026,N_2185);
or U4629 (N_4629,N_3632,N_3706);
or U4630 (N_4630,N_2355,N_3352);
nor U4631 (N_4631,N_3845,N_2112);
and U4632 (N_4632,N_2786,N_3736);
nand U4633 (N_4633,N_2152,N_2726);
or U4634 (N_4634,N_3041,N_3994);
or U4635 (N_4635,N_2825,N_2945);
and U4636 (N_4636,N_3273,N_2941);
nand U4637 (N_4637,N_2866,N_3504);
or U4638 (N_4638,N_2536,N_3716);
and U4639 (N_4639,N_3507,N_2769);
nor U4640 (N_4640,N_2980,N_3638);
nor U4641 (N_4641,N_2891,N_2401);
nand U4642 (N_4642,N_3625,N_3244);
or U4643 (N_4643,N_2436,N_2683);
or U4644 (N_4644,N_3220,N_3547);
and U4645 (N_4645,N_3633,N_3330);
or U4646 (N_4646,N_2371,N_3752);
nor U4647 (N_4647,N_3573,N_2098);
nand U4648 (N_4648,N_2048,N_2966);
or U4649 (N_4649,N_3773,N_3703);
nand U4650 (N_4650,N_2803,N_3665);
and U4651 (N_4651,N_2317,N_2466);
xnor U4652 (N_4652,N_2052,N_3197);
and U4653 (N_4653,N_3650,N_2824);
or U4654 (N_4654,N_2574,N_3081);
xnor U4655 (N_4655,N_2972,N_3841);
or U4656 (N_4656,N_3666,N_3126);
and U4657 (N_4657,N_3245,N_3620);
nand U4658 (N_4658,N_2101,N_3825);
nor U4659 (N_4659,N_2584,N_3677);
and U4660 (N_4660,N_2546,N_3368);
nor U4661 (N_4661,N_3967,N_3525);
nand U4662 (N_4662,N_3467,N_2061);
nand U4663 (N_4663,N_2375,N_3129);
nor U4664 (N_4664,N_3755,N_3001);
nand U4665 (N_4665,N_3668,N_2621);
nor U4666 (N_4666,N_3125,N_2252);
or U4667 (N_4667,N_3446,N_2278);
nand U4668 (N_4668,N_2964,N_3754);
or U4669 (N_4669,N_3165,N_3779);
nand U4670 (N_4670,N_2684,N_2916);
nor U4671 (N_4671,N_2982,N_2614);
or U4672 (N_4672,N_2429,N_3083);
and U4673 (N_4673,N_2890,N_2977);
and U4674 (N_4674,N_2741,N_3194);
and U4675 (N_4675,N_2872,N_3621);
nand U4676 (N_4676,N_2596,N_2332);
nand U4677 (N_4677,N_3079,N_2256);
xor U4678 (N_4678,N_3612,N_2529);
nand U4679 (N_4679,N_3414,N_3127);
nor U4680 (N_4680,N_2055,N_3932);
nor U4681 (N_4681,N_2947,N_3945);
nand U4682 (N_4682,N_3868,N_2486);
or U4683 (N_4683,N_3306,N_3936);
or U4684 (N_4684,N_2040,N_2213);
or U4685 (N_4685,N_3782,N_2233);
or U4686 (N_4686,N_3299,N_2772);
or U4687 (N_4687,N_3192,N_2352);
nand U4688 (N_4688,N_2249,N_2595);
nand U4689 (N_4689,N_2540,N_3461);
nand U4690 (N_4690,N_2914,N_3356);
and U4691 (N_4691,N_3007,N_2696);
and U4692 (N_4692,N_3907,N_3955);
nand U4693 (N_4693,N_3676,N_3257);
nor U4694 (N_4694,N_2483,N_2129);
nor U4695 (N_4695,N_2232,N_3495);
nand U4696 (N_4696,N_2709,N_2467);
xnor U4697 (N_4697,N_3272,N_3771);
nand U4698 (N_4698,N_3747,N_2457);
nor U4699 (N_4699,N_2091,N_2708);
and U4700 (N_4700,N_3781,N_3628);
nor U4701 (N_4701,N_2958,N_3998);
nor U4702 (N_4702,N_3164,N_2078);
or U4703 (N_4703,N_2926,N_3289);
nor U4704 (N_4704,N_2124,N_2672);
nor U4705 (N_4705,N_2531,N_2411);
and U4706 (N_4706,N_3433,N_2960);
xor U4707 (N_4707,N_3176,N_2632);
or U4708 (N_4708,N_3803,N_3969);
and U4709 (N_4709,N_2134,N_2971);
and U4710 (N_4710,N_2508,N_3241);
nor U4711 (N_4711,N_3075,N_2628);
nor U4712 (N_4712,N_2507,N_3750);
or U4713 (N_4713,N_3077,N_2878);
or U4714 (N_4714,N_3318,N_2217);
nand U4715 (N_4715,N_2723,N_3179);
or U4716 (N_4716,N_2073,N_2194);
or U4717 (N_4717,N_3708,N_2659);
or U4718 (N_4718,N_3214,N_3904);
or U4719 (N_4719,N_2747,N_3821);
nand U4720 (N_4720,N_3602,N_2025);
or U4721 (N_4721,N_3365,N_2074);
nand U4722 (N_4722,N_3704,N_3815);
nand U4723 (N_4723,N_2812,N_2273);
nor U4724 (N_4724,N_3118,N_2258);
and U4725 (N_4725,N_3699,N_2748);
or U4726 (N_4726,N_2515,N_3255);
and U4727 (N_4727,N_3048,N_2251);
or U4728 (N_4728,N_3040,N_3488);
nand U4729 (N_4729,N_3926,N_2963);
or U4730 (N_4730,N_3062,N_2294);
and U4731 (N_4731,N_2287,N_3256);
and U4732 (N_4732,N_2207,N_2385);
or U4733 (N_4733,N_3088,N_2188);
or U4734 (N_4734,N_3764,N_3442);
or U4735 (N_4735,N_2422,N_2234);
nor U4736 (N_4736,N_2155,N_2349);
nand U4737 (N_4737,N_2096,N_3285);
or U4738 (N_4738,N_2323,N_2935);
or U4739 (N_4739,N_2248,N_2853);
or U4740 (N_4740,N_2189,N_3246);
and U4741 (N_4741,N_3465,N_3371);
and U4742 (N_4742,N_2168,N_3268);
or U4743 (N_4743,N_2754,N_3096);
nor U4744 (N_4744,N_2802,N_2167);
and U4745 (N_4745,N_3851,N_3052);
and U4746 (N_4746,N_2502,N_2176);
nor U4747 (N_4747,N_2036,N_2533);
nand U4748 (N_4748,N_3558,N_2034);
nor U4749 (N_4749,N_3914,N_3146);
or U4750 (N_4750,N_3788,N_2216);
and U4751 (N_4751,N_3689,N_3486);
or U4752 (N_4752,N_2279,N_2001);
and U4753 (N_4753,N_2257,N_2326);
nand U4754 (N_4754,N_3043,N_2530);
nor U4755 (N_4755,N_2773,N_2913);
and U4756 (N_4756,N_2870,N_3464);
nand U4757 (N_4757,N_3234,N_2855);
nor U4758 (N_4758,N_3515,N_2673);
nor U4759 (N_4759,N_3132,N_3760);
and U4760 (N_4760,N_2009,N_3429);
or U4761 (N_4761,N_2629,N_3263);
or U4762 (N_4762,N_2470,N_3231);
nor U4763 (N_4763,N_2020,N_3891);
nand U4764 (N_4764,N_2984,N_3117);
and U4765 (N_4765,N_2885,N_3346);
and U4766 (N_4766,N_3519,N_2724);
and U4767 (N_4767,N_3672,N_3698);
nand U4768 (N_4768,N_3128,N_3712);
or U4769 (N_4769,N_2731,N_2408);
and U4770 (N_4770,N_2244,N_3024);
nand U4771 (N_4771,N_2841,N_3820);
and U4772 (N_4772,N_2636,N_2186);
nand U4773 (N_4773,N_2809,N_3934);
nand U4774 (N_4774,N_3424,N_3015);
nand U4775 (N_4775,N_2184,N_3763);
nand U4776 (N_4776,N_3459,N_2344);
or U4777 (N_4777,N_2768,N_3187);
nor U4778 (N_4778,N_3586,N_3283);
and U4779 (N_4779,N_3599,N_2543);
nor U4780 (N_4780,N_2123,N_2062);
nor U4781 (N_4781,N_2267,N_2437);
nand U4782 (N_4782,N_2742,N_3623);
and U4783 (N_4783,N_3279,N_2090);
or U4784 (N_4784,N_2750,N_2174);
nand U4785 (N_4785,N_2122,N_2250);
nor U4786 (N_4786,N_2390,N_2917);
nor U4787 (N_4787,N_3544,N_2453);
or U4788 (N_4788,N_2762,N_2589);
nor U4789 (N_4789,N_3314,N_3923);
nor U4790 (N_4790,N_3898,N_3333);
and U4791 (N_4791,N_3770,N_2640);
or U4792 (N_4792,N_2936,N_2309);
and U4793 (N_4793,N_3740,N_3086);
and U4794 (N_4794,N_2856,N_2661);
and U4795 (N_4795,N_3977,N_2281);
nor U4796 (N_4796,N_2224,N_2845);
nor U4797 (N_4797,N_3890,N_2455);
and U4798 (N_4798,N_3049,N_2846);
and U4799 (N_4799,N_2766,N_2017);
xor U4800 (N_4800,N_2382,N_3627);
nand U4801 (N_4801,N_2692,N_3466);
and U4802 (N_4802,N_2484,N_3106);
nor U4803 (N_4803,N_2093,N_3189);
and U4804 (N_4804,N_2815,N_3931);
nor U4805 (N_4805,N_2428,N_2452);
or U4806 (N_4806,N_3499,N_2918);
nand U4807 (N_4807,N_2785,N_2925);
and U4808 (N_4808,N_3687,N_2246);
or U4809 (N_4809,N_2826,N_3982);
nand U4810 (N_4810,N_3843,N_3363);
and U4811 (N_4811,N_3606,N_2211);
nand U4812 (N_4812,N_2805,N_3817);
and U4813 (N_4813,N_2404,N_3400);
nand U4814 (N_4814,N_2818,N_3615);
or U4815 (N_4815,N_3388,N_2677);
nor U4816 (N_4816,N_2986,N_2763);
or U4817 (N_4817,N_2678,N_3006);
and U4818 (N_4818,N_3549,N_3541);
and U4819 (N_4819,N_2039,N_2364);
nand U4820 (N_4820,N_2934,N_2545);
nand U4821 (N_4821,N_2500,N_3995);
xor U4822 (N_4822,N_3087,N_3085);
xor U4823 (N_4823,N_3159,N_3546);
and U4824 (N_4824,N_3500,N_2407);
or U4825 (N_4825,N_3787,N_3927);
or U4826 (N_4826,N_2671,N_2699);
xnor U4827 (N_4827,N_2942,N_3011);
nand U4828 (N_4828,N_2808,N_2215);
xnor U4829 (N_4829,N_3569,N_3407);
nand U4830 (N_4830,N_2745,N_3780);
nand U4831 (N_4831,N_3595,N_3651);
or U4832 (N_4832,N_3905,N_3254);
or U4833 (N_4833,N_2151,N_3662);
and U4834 (N_4834,N_2832,N_3534);
nand U4835 (N_4835,N_2100,N_3552);
and U4836 (N_4836,N_3795,N_2446);
and U4837 (N_4837,N_2701,N_2028);
or U4838 (N_4838,N_2465,N_2425);
or U4839 (N_4839,N_2704,N_2143);
nor U4840 (N_4840,N_3420,N_2102);
nor U4841 (N_4841,N_3705,N_2800);
and U4842 (N_4842,N_3713,N_2179);
and U4843 (N_4843,N_3673,N_2004);
and U4844 (N_4844,N_3298,N_3996);
and U4845 (N_4845,N_2200,N_3864);
and U4846 (N_4846,N_3899,N_2126);
or U4847 (N_4847,N_3940,N_3430);
and U4848 (N_4848,N_3301,N_3100);
xnor U4849 (N_4849,N_2511,N_2297);
nand U4850 (N_4850,N_3951,N_3960);
or U4851 (N_4851,N_2558,N_2679);
and U4852 (N_4852,N_2608,N_3417);
nand U4853 (N_4853,N_2431,N_3045);
and U4854 (N_4854,N_2430,N_2318);
nand U4855 (N_4855,N_2943,N_2097);
nand U4856 (N_4856,N_2041,N_2108);
nor U4857 (N_4857,N_2643,N_3992);
nor U4858 (N_4858,N_2183,N_3271);
nand U4859 (N_4859,N_3800,N_2069);
and U4860 (N_4860,N_3866,N_3997);
nand U4861 (N_4861,N_2191,N_3970);
and U4862 (N_4862,N_3412,N_3824);
nand U4863 (N_4863,N_2572,N_3809);
xnor U4864 (N_4864,N_2929,N_3629);
nor U4865 (N_4865,N_3317,N_2154);
or U4866 (N_4866,N_2900,N_2685);
nor U4867 (N_4867,N_2810,N_3022);
nor U4868 (N_4868,N_3070,N_2764);
nand U4869 (N_4869,N_2938,N_3304);
or U4870 (N_4870,N_3686,N_3520);
or U4871 (N_4871,N_2616,N_3422);
nor U4872 (N_4872,N_3325,N_3294);
nand U4873 (N_4873,N_2923,N_3387);
and U4874 (N_4874,N_3366,N_2311);
or U4875 (N_4875,N_3392,N_3406);
and U4876 (N_4876,N_3018,N_2338);
nand U4877 (N_4877,N_2038,N_3047);
and U4878 (N_4878,N_3066,N_2657);
nor U4879 (N_4879,N_2259,N_3786);
nor U4880 (N_4880,N_2005,N_3853);
and U4881 (N_4881,N_3359,N_3974);
and U4882 (N_4882,N_2214,N_2474);
and U4883 (N_4883,N_2027,N_3225);
nor U4884 (N_4884,N_3113,N_2405);
and U4885 (N_4885,N_2569,N_3448);
nor U4886 (N_4886,N_3946,N_3690);
nand U4887 (N_4887,N_3451,N_3823);
nor U4888 (N_4888,N_3548,N_3976);
nor U4889 (N_4889,N_2767,N_2493);
nand U4890 (N_4890,N_3721,N_2974);
xnor U4891 (N_4891,N_2322,N_2650);
and U4892 (N_4892,N_3962,N_2919);
nand U4893 (N_4893,N_2667,N_3883);
nor U4894 (N_4894,N_2178,N_2423);
nor U4895 (N_4895,N_3808,N_3174);
and U4896 (N_4896,N_3709,N_2730);
nor U4897 (N_4897,N_3312,N_2756);
and U4898 (N_4898,N_2915,N_3064);
nor U4899 (N_4899,N_3409,N_2254);
and U4900 (N_4900,N_2851,N_2784);
nor U4901 (N_4901,N_2544,N_2030);
xor U4902 (N_4902,N_3560,N_2857);
nor U4903 (N_4903,N_3042,N_2169);
or U4904 (N_4904,N_2979,N_3720);
nand U4905 (N_4905,N_2606,N_2887);
nand U4906 (N_4906,N_2995,N_2903);
nand U4907 (N_4907,N_2976,N_2462);
nand U4908 (N_4908,N_3592,N_3916);
or U4909 (N_4909,N_2345,N_2440);
and U4910 (N_4910,N_3741,N_3228);
or U4911 (N_4911,N_2386,N_3167);
nor U4912 (N_4912,N_3757,N_3456);
nor U4913 (N_4913,N_2873,N_2402);
and U4914 (N_4914,N_2551,N_3428);
nand U4915 (N_4915,N_2447,N_3483);
nand U4916 (N_4916,N_2222,N_3844);
and U4917 (N_4917,N_3600,N_3774);
or U4918 (N_4918,N_3198,N_3288);
nand U4919 (N_4919,N_2305,N_2602);
and U4920 (N_4920,N_2148,N_3157);
nand U4921 (N_4921,N_2889,N_3949);
nand U4922 (N_4922,N_3204,N_2162);
or U4923 (N_4923,N_2714,N_3724);
or U4924 (N_4924,N_2734,N_3002);
or U4925 (N_4925,N_2088,N_3286);
or U4926 (N_4926,N_2720,N_3186);
and U4927 (N_4927,N_3019,N_3261);
or U4928 (N_4928,N_3513,N_2099);
nand U4929 (N_4929,N_2781,N_2218);
and U4930 (N_4930,N_2133,N_2662);
or U4931 (N_4931,N_3149,N_2519);
nand U4932 (N_4932,N_3284,N_3983);
nor U4933 (N_4933,N_2395,N_3444);
nand U4934 (N_4934,N_2783,N_2555);
and U4935 (N_4935,N_2292,N_3804);
nor U4936 (N_4936,N_3240,N_2512);
nand U4937 (N_4937,N_3258,N_2488);
or U4938 (N_4938,N_2883,N_3942);
nor U4939 (N_4939,N_2010,N_3389);
nand U4940 (N_4940,N_3700,N_3340);
xnor U4941 (N_4941,N_3203,N_2695);
and U4942 (N_4942,N_3026,N_2173);
and U4943 (N_4943,N_2517,N_3696);
or U4944 (N_4944,N_2881,N_2400);
nor U4945 (N_4945,N_3745,N_3205);
or U4946 (N_4946,N_2729,N_3329);
nand U4947 (N_4947,N_2413,N_2645);
nor U4948 (N_4948,N_2223,N_3647);
nor U4949 (N_4949,N_3450,N_3016);
nor U4950 (N_4950,N_2928,N_3418);
and U4951 (N_4951,N_3530,N_3762);
nor U4952 (N_4952,N_3027,N_3865);
nor U4953 (N_4953,N_3173,N_2427);
xnor U4954 (N_4954,N_3635,N_2829);
nand U4955 (N_4955,N_2557,N_2303);
nor U4956 (N_4956,N_2265,N_2837);
nor U4957 (N_4957,N_3158,N_3751);
nand U4958 (N_4958,N_3037,N_3105);
or U4959 (N_4959,N_2113,N_2253);
nor U4960 (N_4960,N_2563,N_3756);
or U4961 (N_4961,N_3355,N_2351);
nand U4962 (N_4962,N_3379,N_2412);
or U4963 (N_4963,N_2757,N_3950);
nand U4964 (N_4964,N_3535,N_3827);
and U4965 (N_4965,N_3437,N_2308);
and U4966 (N_4966,N_2909,N_2719);
nand U4967 (N_4967,N_3219,N_3648);
nand U4968 (N_4968,N_3103,N_3589);
and U4969 (N_4969,N_3834,N_3017);
and U4970 (N_4970,N_3761,N_2954);
and U4971 (N_4971,N_2497,N_2300);
nor U4972 (N_4972,N_2392,N_3473);
nor U4973 (N_4973,N_2831,N_2840);
or U4974 (N_4974,N_3529,N_3181);
or U4975 (N_4975,N_2759,N_2573);
nand U4976 (N_4976,N_3862,N_2461);
and U4977 (N_4977,N_3688,N_3460);
or U4978 (N_4978,N_2817,N_3044);
nor U4979 (N_4979,N_3526,N_3565);
nor U4980 (N_4980,N_2710,N_3470);
nor U4981 (N_4981,N_2961,N_2668);
nor U4982 (N_4982,N_3797,N_3593);
nand U4983 (N_4983,N_3888,N_3656);
nor U4984 (N_4984,N_3886,N_2049);
nand U4985 (N_4985,N_2131,N_2970);
nor U4986 (N_4986,N_3961,N_3305);
nand U4987 (N_4987,N_2652,N_3046);
nand U4988 (N_4988,N_2790,N_2518);
nor U4989 (N_4989,N_2236,N_2221);
nand U4990 (N_4990,N_3769,N_3154);
or U4991 (N_4991,N_2931,N_3320);
and U4992 (N_4992,N_3402,N_2819);
or U4993 (N_4993,N_2115,N_2210);
nand U4994 (N_4994,N_3292,N_2988);
or U4995 (N_4995,N_2642,N_3065);
or U4996 (N_4996,N_2549,N_3137);
and U4997 (N_4997,N_2586,N_3577);
and U4998 (N_4998,N_2806,N_3410);
nor U4999 (N_4999,N_2998,N_3380);
or U5000 (N_5000,N_3810,N_2318);
and U5001 (N_5001,N_3052,N_3622);
nand U5002 (N_5002,N_2126,N_3482);
nand U5003 (N_5003,N_2383,N_3188);
nand U5004 (N_5004,N_3265,N_3380);
or U5005 (N_5005,N_2084,N_2049);
nand U5006 (N_5006,N_2192,N_2218);
xor U5007 (N_5007,N_3613,N_2131);
xor U5008 (N_5008,N_2075,N_3480);
nor U5009 (N_5009,N_3633,N_2109);
or U5010 (N_5010,N_3921,N_2742);
and U5011 (N_5011,N_2989,N_2586);
or U5012 (N_5012,N_2876,N_3141);
and U5013 (N_5013,N_3746,N_3049);
nor U5014 (N_5014,N_3207,N_2267);
and U5015 (N_5015,N_3134,N_3675);
and U5016 (N_5016,N_2467,N_3847);
and U5017 (N_5017,N_3795,N_3794);
and U5018 (N_5018,N_3679,N_3782);
nor U5019 (N_5019,N_2687,N_2424);
nand U5020 (N_5020,N_3821,N_3482);
or U5021 (N_5021,N_3229,N_2335);
nand U5022 (N_5022,N_2684,N_3142);
nor U5023 (N_5023,N_2585,N_3818);
nor U5024 (N_5024,N_3000,N_3013);
nand U5025 (N_5025,N_3500,N_2371);
nor U5026 (N_5026,N_2726,N_2033);
nand U5027 (N_5027,N_3121,N_3525);
nand U5028 (N_5028,N_2309,N_2988);
nor U5029 (N_5029,N_2465,N_3519);
and U5030 (N_5030,N_2475,N_3903);
or U5031 (N_5031,N_3259,N_2398);
nand U5032 (N_5032,N_2985,N_3588);
and U5033 (N_5033,N_2712,N_2510);
nand U5034 (N_5034,N_2421,N_3320);
and U5035 (N_5035,N_2487,N_2139);
nand U5036 (N_5036,N_3570,N_2690);
and U5037 (N_5037,N_3609,N_2583);
nand U5038 (N_5038,N_2055,N_3320);
nor U5039 (N_5039,N_3778,N_3273);
xnor U5040 (N_5040,N_3235,N_3556);
nor U5041 (N_5041,N_3821,N_2497);
nand U5042 (N_5042,N_2096,N_3056);
nand U5043 (N_5043,N_3567,N_3481);
or U5044 (N_5044,N_3962,N_3662);
or U5045 (N_5045,N_3381,N_2791);
and U5046 (N_5046,N_3391,N_3029);
nand U5047 (N_5047,N_2974,N_2464);
or U5048 (N_5048,N_2401,N_2392);
nor U5049 (N_5049,N_3546,N_2501);
nand U5050 (N_5050,N_3787,N_3709);
nor U5051 (N_5051,N_3047,N_3650);
nor U5052 (N_5052,N_2698,N_3227);
nor U5053 (N_5053,N_2166,N_2948);
nand U5054 (N_5054,N_2681,N_2908);
nand U5055 (N_5055,N_2567,N_3716);
or U5056 (N_5056,N_3978,N_3448);
nand U5057 (N_5057,N_2145,N_3537);
or U5058 (N_5058,N_3427,N_2727);
and U5059 (N_5059,N_2833,N_3808);
and U5060 (N_5060,N_2330,N_2637);
nor U5061 (N_5061,N_2881,N_3436);
nor U5062 (N_5062,N_2125,N_3817);
xnor U5063 (N_5063,N_3704,N_3250);
or U5064 (N_5064,N_3149,N_3384);
and U5065 (N_5065,N_2467,N_3131);
or U5066 (N_5066,N_3729,N_3177);
or U5067 (N_5067,N_3434,N_2143);
nand U5068 (N_5068,N_3350,N_2347);
nand U5069 (N_5069,N_3081,N_3137);
or U5070 (N_5070,N_3239,N_3739);
nand U5071 (N_5071,N_2982,N_3212);
or U5072 (N_5072,N_3898,N_3872);
or U5073 (N_5073,N_3812,N_2751);
or U5074 (N_5074,N_3649,N_3761);
nand U5075 (N_5075,N_3510,N_2907);
nand U5076 (N_5076,N_3086,N_2568);
nand U5077 (N_5077,N_2345,N_3102);
or U5078 (N_5078,N_2577,N_3735);
nand U5079 (N_5079,N_3033,N_2759);
nor U5080 (N_5080,N_2523,N_3641);
or U5081 (N_5081,N_3979,N_2267);
nor U5082 (N_5082,N_3305,N_2949);
nand U5083 (N_5083,N_3380,N_3713);
nor U5084 (N_5084,N_3117,N_3412);
and U5085 (N_5085,N_2371,N_3747);
and U5086 (N_5086,N_3316,N_2107);
nand U5087 (N_5087,N_2607,N_3074);
nor U5088 (N_5088,N_2402,N_3509);
nor U5089 (N_5089,N_3766,N_3704);
and U5090 (N_5090,N_3441,N_3740);
nand U5091 (N_5091,N_2079,N_3367);
xnor U5092 (N_5092,N_3593,N_2534);
and U5093 (N_5093,N_2884,N_2516);
nor U5094 (N_5094,N_2655,N_2543);
nand U5095 (N_5095,N_3282,N_3549);
and U5096 (N_5096,N_2716,N_2705);
nor U5097 (N_5097,N_3556,N_2370);
or U5098 (N_5098,N_2995,N_2338);
and U5099 (N_5099,N_3878,N_3497);
nor U5100 (N_5100,N_3371,N_2787);
and U5101 (N_5101,N_3761,N_3602);
nor U5102 (N_5102,N_3740,N_3057);
or U5103 (N_5103,N_2499,N_3356);
nor U5104 (N_5104,N_2474,N_2030);
or U5105 (N_5105,N_3644,N_3541);
nand U5106 (N_5106,N_3676,N_3859);
or U5107 (N_5107,N_3111,N_3499);
nor U5108 (N_5108,N_3968,N_2804);
nor U5109 (N_5109,N_2335,N_2135);
nand U5110 (N_5110,N_2879,N_3349);
and U5111 (N_5111,N_3124,N_2654);
or U5112 (N_5112,N_3155,N_2213);
and U5113 (N_5113,N_2810,N_2478);
or U5114 (N_5114,N_3123,N_2430);
and U5115 (N_5115,N_3812,N_3511);
or U5116 (N_5116,N_2009,N_2540);
nand U5117 (N_5117,N_3631,N_3735);
nand U5118 (N_5118,N_3912,N_2265);
or U5119 (N_5119,N_3647,N_3165);
nand U5120 (N_5120,N_2196,N_2512);
or U5121 (N_5121,N_3085,N_3955);
or U5122 (N_5122,N_2543,N_3969);
and U5123 (N_5123,N_3457,N_2702);
nand U5124 (N_5124,N_3401,N_2579);
and U5125 (N_5125,N_2323,N_3029);
and U5126 (N_5126,N_2465,N_3320);
nand U5127 (N_5127,N_2839,N_2427);
and U5128 (N_5128,N_3407,N_3447);
nor U5129 (N_5129,N_2055,N_2458);
nor U5130 (N_5130,N_3622,N_2043);
nand U5131 (N_5131,N_2357,N_3963);
nand U5132 (N_5132,N_2501,N_2469);
and U5133 (N_5133,N_2052,N_3221);
nand U5134 (N_5134,N_2020,N_2057);
nand U5135 (N_5135,N_2858,N_2636);
and U5136 (N_5136,N_2548,N_3656);
nor U5137 (N_5137,N_3938,N_3058);
or U5138 (N_5138,N_3425,N_3892);
nand U5139 (N_5139,N_3801,N_2810);
and U5140 (N_5140,N_3860,N_2157);
nor U5141 (N_5141,N_2394,N_2194);
and U5142 (N_5142,N_3584,N_3307);
nand U5143 (N_5143,N_2059,N_2997);
xor U5144 (N_5144,N_2293,N_2500);
or U5145 (N_5145,N_2156,N_2155);
or U5146 (N_5146,N_2938,N_3832);
nand U5147 (N_5147,N_2334,N_2668);
xor U5148 (N_5148,N_2528,N_3285);
and U5149 (N_5149,N_3513,N_2103);
and U5150 (N_5150,N_2309,N_3460);
nand U5151 (N_5151,N_2557,N_2449);
or U5152 (N_5152,N_2291,N_3915);
and U5153 (N_5153,N_3059,N_2027);
or U5154 (N_5154,N_3480,N_2749);
and U5155 (N_5155,N_2056,N_2280);
or U5156 (N_5156,N_3422,N_3341);
or U5157 (N_5157,N_2617,N_2426);
and U5158 (N_5158,N_2394,N_2819);
and U5159 (N_5159,N_2675,N_3854);
xnor U5160 (N_5160,N_3014,N_2596);
nand U5161 (N_5161,N_2840,N_3851);
nand U5162 (N_5162,N_3070,N_2076);
or U5163 (N_5163,N_3779,N_3242);
nor U5164 (N_5164,N_2949,N_2244);
and U5165 (N_5165,N_2787,N_3727);
nand U5166 (N_5166,N_3649,N_3043);
nand U5167 (N_5167,N_3470,N_3119);
and U5168 (N_5168,N_3045,N_2291);
nor U5169 (N_5169,N_2813,N_2080);
nand U5170 (N_5170,N_2417,N_2337);
nor U5171 (N_5171,N_2661,N_2813);
and U5172 (N_5172,N_2958,N_3027);
or U5173 (N_5173,N_2537,N_2952);
nand U5174 (N_5174,N_2141,N_2037);
nand U5175 (N_5175,N_2822,N_2042);
and U5176 (N_5176,N_2932,N_2919);
nand U5177 (N_5177,N_3694,N_2136);
nor U5178 (N_5178,N_2774,N_2644);
and U5179 (N_5179,N_2507,N_2989);
nor U5180 (N_5180,N_2105,N_2963);
nand U5181 (N_5181,N_2652,N_2087);
or U5182 (N_5182,N_2853,N_3687);
or U5183 (N_5183,N_3905,N_3924);
and U5184 (N_5184,N_2634,N_3633);
nor U5185 (N_5185,N_3436,N_3616);
nand U5186 (N_5186,N_3214,N_3892);
and U5187 (N_5187,N_2779,N_3618);
and U5188 (N_5188,N_2636,N_2988);
or U5189 (N_5189,N_3388,N_2251);
nor U5190 (N_5190,N_2043,N_3675);
and U5191 (N_5191,N_3401,N_3415);
or U5192 (N_5192,N_2802,N_3457);
and U5193 (N_5193,N_3939,N_2032);
nor U5194 (N_5194,N_2831,N_3454);
nor U5195 (N_5195,N_2970,N_2601);
nand U5196 (N_5196,N_3083,N_2717);
nor U5197 (N_5197,N_3035,N_2898);
or U5198 (N_5198,N_2065,N_3544);
nand U5199 (N_5199,N_2879,N_3621);
xor U5200 (N_5200,N_2393,N_2507);
or U5201 (N_5201,N_2730,N_3924);
nand U5202 (N_5202,N_2754,N_2151);
nor U5203 (N_5203,N_2391,N_2775);
nor U5204 (N_5204,N_3918,N_2299);
and U5205 (N_5205,N_3917,N_3253);
nor U5206 (N_5206,N_3068,N_3891);
nand U5207 (N_5207,N_3859,N_2358);
or U5208 (N_5208,N_2673,N_2207);
or U5209 (N_5209,N_2420,N_3893);
and U5210 (N_5210,N_2433,N_3088);
nand U5211 (N_5211,N_2825,N_2854);
nor U5212 (N_5212,N_2219,N_2369);
nand U5213 (N_5213,N_3803,N_3729);
nand U5214 (N_5214,N_3194,N_2657);
and U5215 (N_5215,N_3889,N_2140);
and U5216 (N_5216,N_2890,N_2758);
nor U5217 (N_5217,N_2075,N_3628);
or U5218 (N_5218,N_2650,N_2898);
nor U5219 (N_5219,N_3058,N_3928);
nand U5220 (N_5220,N_2238,N_3081);
nor U5221 (N_5221,N_2149,N_2538);
and U5222 (N_5222,N_2081,N_2278);
nand U5223 (N_5223,N_2229,N_2759);
or U5224 (N_5224,N_2951,N_3006);
nor U5225 (N_5225,N_3025,N_2672);
and U5226 (N_5226,N_2068,N_2459);
nor U5227 (N_5227,N_2849,N_3354);
or U5228 (N_5228,N_3818,N_3997);
or U5229 (N_5229,N_3889,N_3990);
or U5230 (N_5230,N_3853,N_3673);
nor U5231 (N_5231,N_2341,N_3303);
nand U5232 (N_5232,N_2403,N_3788);
nand U5233 (N_5233,N_2455,N_3223);
nor U5234 (N_5234,N_3796,N_3341);
xor U5235 (N_5235,N_3759,N_2067);
and U5236 (N_5236,N_3834,N_2694);
or U5237 (N_5237,N_2593,N_3227);
nand U5238 (N_5238,N_2403,N_3683);
nor U5239 (N_5239,N_2271,N_3935);
nand U5240 (N_5240,N_2099,N_3537);
or U5241 (N_5241,N_3744,N_3799);
nand U5242 (N_5242,N_3506,N_2502);
nand U5243 (N_5243,N_3236,N_2354);
nand U5244 (N_5244,N_3344,N_2097);
and U5245 (N_5245,N_2276,N_2948);
or U5246 (N_5246,N_3927,N_3568);
and U5247 (N_5247,N_3319,N_3627);
nand U5248 (N_5248,N_2379,N_3840);
nand U5249 (N_5249,N_3226,N_3535);
or U5250 (N_5250,N_2528,N_3358);
nand U5251 (N_5251,N_2282,N_3311);
nor U5252 (N_5252,N_3794,N_3011);
nor U5253 (N_5253,N_3102,N_2430);
and U5254 (N_5254,N_3050,N_3203);
nor U5255 (N_5255,N_3228,N_3198);
and U5256 (N_5256,N_3375,N_3013);
nor U5257 (N_5257,N_3684,N_3408);
nand U5258 (N_5258,N_3811,N_3504);
nand U5259 (N_5259,N_3450,N_3559);
nor U5260 (N_5260,N_2817,N_3655);
or U5261 (N_5261,N_2914,N_2807);
nand U5262 (N_5262,N_2292,N_3169);
and U5263 (N_5263,N_2446,N_2161);
or U5264 (N_5264,N_2848,N_2534);
and U5265 (N_5265,N_2515,N_3899);
or U5266 (N_5266,N_2250,N_3679);
and U5267 (N_5267,N_3257,N_3159);
or U5268 (N_5268,N_3819,N_3291);
xor U5269 (N_5269,N_3299,N_3636);
or U5270 (N_5270,N_3304,N_3362);
nor U5271 (N_5271,N_2224,N_3377);
and U5272 (N_5272,N_3910,N_2268);
nand U5273 (N_5273,N_3062,N_2815);
or U5274 (N_5274,N_3843,N_2037);
or U5275 (N_5275,N_3659,N_3765);
nor U5276 (N_5276,N_2207,N_3504);
and U5277 (N_5277,N_3305,N_3174);
or U5278 (N_5278,N_2361,N_2933);
nand U5279 (N_5279,N_3868,N_2963);
and U5280 (N_5280,N_2205,N_3335);
or U5281 (N_5281,N_2085,N_3551);
and U5282 (N_5282,N_3241,N_2643);
and U5283 (N_5283,N_2974,N_3372);
nand U5284 (N_5284,N_3140,N_3143);
nor U5285 (N_5285,N_3036,N_3727);
and U5286 (N_5286,N_2553,N_2065);
nor U5287 (N_5287,N_3646,N_2039);
nand U5288 (N_5288,N_3444,N_3112);
and U5289 (N_5289,N_3844,N_2356);
and U5290 (N_5290,N_2721,N_2789);
or U5291 (N_5291,N_2541,N_3494);
nand U5292 (N_5292,N_3720,N_3225);
and U5293 (N_5293,N_3103,N_3718);
nand U5294 (N_5294,N_3777,N_3212);
nand U5295 (N_5295,N_3934,N_3077);
and U5296 (N_5296,N_3413,N_2444);
and U5297 (N_5297,N_2138,N_3735);
nand U5298 (N_5298,N_2409,N_3346);
xnor U5299 (N_5299,N_2262,N_2152);
xor U5300 (N_5300,N_3964,N_2535);
nand U5301 (N_5301,N_2555,N_3781);
nand U5302 (N_5302,N_3915,N_2404);
and U5303 (N_5303,N_3966,N_3402);
nor U5304 (N_5304,N_3950,N_2883);
and U5305 (N_5305,N_3901,N_3930);
or U5306 (N_5306,N_2512,N_3485);
or U5307 (N_5307,N_2777,N_2012);
and U5308 (N_5308,N_3294,N_2395);
nand U5309 (N_5309,N_2123,N_2335);
nor U5310 (N_5310,N_3701,N_2381);
nand U5311 (N_5311,N_3309,N_2836);
nor U5312 (N_5312,N_2857,N_2701);
nand U5313 (N_5313,N_3432,N_3523);
or U5314 (N_5314,N_2927,N_3359);
nand U5315 (N_5315,N_3467,N_2604);
nand U5316 (N_5316,N_2336,N_3908);
and U5317 (N_5317,N_2419,N_2401);
xor U5318 (N_5318,N_2943,N_3953);
nor U5319 (N_5319,N_3632,N_2845);
nor U5320 (N_5320,N_3615,N_2753);
nor U5321 (N_5321,N_2510,N_2795);
nor U5322 (N_5322,N_2482,N_2982);
nor U5323 (N_5323,N_3567,N_3811);
nand U5324 (N_5324,N_3917,N_2508);
or U5325 (N_5325,N_2530,N_2417);
or U5326 (N_5326,N_3333,N_2956);
nor U5327 (N_5327,N_3712,N_3064);
nor U5328 (N_5328,N_3245,N_2153);
or U5329 (N_5329,N_3175,N_2161);
nor U5330 (N_5330,N_2952,N_2810);
nand U5331 (N_5331,N_2070,N_3831);
and U5332 (N_5332,N_3452,N_3135);
nand U5333 (N_5333,N_2358,N_3063);
nor U5334 (N_5334,N_2223,N_3993);
nor U5335 (N_5335,N_3691,N_2996);
nand U5336 (N_5336,N_2958,N_3719);
nand U5337 (N_5337,N_3082,N_3775);
and U5338 (N_5338,N_2845,N_2905);
and U5339 (N_5339,N_3081,N_3420);
and U5340 (N_5340,N_2029,N_3895);
or U5341 (N_5341,N_2337,N_3691);
nor U5342 (N_5342,N_3415,N_3249);
nand U5343 (N_5343,N_2691,N_2690);
or U5344 (N_5344,N_2796,N_2920);
or U5345 (N_5345,N_2316,N_3546);
nor U5346 (N_5346,N_3586,N_3680);
and U5347 (N_5347,N_3604,N_2056);
or U5348 (N_5348,N_2574,N_2076);
nor U5349 (N_5349,N_2609,N_2883);
nand U5350 (N_5350,N_2961,N_2763);
nand U5351 (N_5351,N_2807,N_2159);
and U5352 (N_5352,N_3048,N_3750);
or U5353 (N_5353,N_3109,N_2825);
xnor U5354 (N_5354,N_3396,N_2693);
or U5355 (N_5355,N_2391,N_2854);
or U5356 (N_5356,N_3995,N_2955);
and U5357 (N_5357,N_3415,N_2417);
nor U5358 (N_5358,N_3868,N_3934);
or U5359 (N_5359,N_2520,N_2168);
or U5360 (N_5360,N_2381,N_2866);
xnor U5361 (N_5361,N_3813,N_3596);
and U5362 (N_5362,N_2064,N_2288);
nand U5363 (N_5363,N_3977,N_3921);
and U5364 (N_5364,N_2335,N_2131);
or U5365 (N_5365,N_3254,N_3669);
and U5366 (N_5366,N_3216,N_3467);
and U5367 (N_5367,N_3122,N_2917);
or U5368 (N_5368,N_3578,N_3119);
nor U5369 (N_5369,N_3033,N_3876);
or U5370 (N_5370,N_2201,N_3857);
nor U5371 (N_5371,N_3627,N_3877);
and U5372 (N_5372,N_2292,N_3319);
nor U5373 (N_5373,N_3805,N_3817);
nand U5374 (N_5374,N_2385,N_3691);
nand U5375 (N_5375,N_2755,N_3298);
nor U5376 (N_5376,N_2927,N_2849);
and U5377 (N_5377,N_3377,N_2529);
and U5378 (N_5378,N_3331,N_2346);
and U5379 (N_5379,N_2799,N_2759);
nand U5380 (N_5380,N_3005,N_3146);
nor U5381 (N_5381,N_3707,N_3768);
or U5382 (N_5382,N_3746,N_2977);
and U5383 (N_5383,N_3505,N_3602);
or U5384 (N_5384,N_3373,N_3685);
nand U5385 (N_5385,N_2945,N_2142);
or U5386 (N_5386,N_2138,N_2985);
and U5387 (N_5387,N_3931,N_3204);
nor U5388 (N_5388,N_3603,N_2020);
nor U5389 (N_5389,N_3914,N_3530);
or U5390 (N_5390,N_3659,N_3893);
nor U5391 (N_5391,N_2015,N_3842);
xor U5392 (N_5392,N_3717,N_3624);
or U5393 (N_5393,N_3131,N_3810);
or U5394 (N_5394,N_2370,N_3924);
and U5395 (N_5395,N_2572,N_2892);
nand U5396 (N_5396,N_3994,N_3275);
or U5397 (N_5397,N_2480,N_2066);
or U5398 (N_5398,N_2692,N_3965);
and U5399 (N_5399,N_2018,N_2852);
nand U5400 (N_5400,N_3444,N_2432);
nand U5401 (N_5401,N_2657,N_3692);
or U5402 (N_5402,N_3661,N_2704);
nand U5403 (N_5403,N_2971,N_2142);
and U5404 (N_5404,N_3173,N_3294);
and U5405 (N_5405,N_2144,N_3505);
and U5406 (N_5406,N_3661,N_2238);
nand U5407 (N_5407,N_3121,N_3035);
nand U5408 (N_5408,N_2660,N_3783);
nand U5409 (N_5409,N_3329,N_2386);
nor U5410 (N_5410,N_2266,N_3894);
nor U5411 (N_5411,N_2077,N_3927);
and U5412 (N_5412,N_2065,N_3608);
and U5413 (N_5413,N_2143,N_3141);
nand U5414 (N_5414,N_3117,N_3649);
nor U5415 (N_5415,N_3173,N_3907);
and U5416 (N_5416,N_3573,N_3256);
or U5417 (N_5417,N_2406,N_3190);
nor U5418 (N_5418,N_3236,N_2127);
nor U5419 (N_5419,N_2596,N_2854);
nand U5420 (N_5420,N_3726,N_2230);
nand U5421 (N_5421,N_3980,N_2134);
nor U5422 (N_5422,N_3035,N_3178);
nor U5423 (N_5423,N_2236,N_3672);
xor U5424 (N_5424,N_3353,N_2415);
nand U5425 (N_5425,N_2400,N_2982);
or U5426 (N_5426,N_3663,N_3449);
and U5427 (N_5427,N_2921,N_2154);
nor U5428 (N_5428,N_2959,N_2565);
nand U5429 (N_5429,N_2499,N_2808);
or U5430 (N_5430,N_3229,N_3705);
and U5431 (N_5431,N_2199,N_2817);
nand U5432 (N_5432,N_3253,N_3024);
nor U5433 (N_5433,N_3445,N_3492);
and U5434 (N_5434,N_2353,N_3134);
and U5435 (N_5435,N_2812,N_2115);
nor U5436 (N_5436,N_2188,N_2200);
and U5437 (N_5437,N_2046,N_3373);
and U5438 (N_5438,N_3234,N_2489);
or U5439 (N_5439,N_2091,N_3486);
and U5440 (N_5440,N_2882,N_2463);
and U5441 (N_5441,N_3278,N_3589);
nor U5442 (N_5442,N_3670,N_2315);
and U5443 (N_5443,N_3285,N_2236);
nand U5444 (N_5444,N_3050,N_3706);
nand U5445 (N_5445,N_2679,N_3825);
and U5446 (N_5446,N_2443,N_3626);
nor U5447 (N_5447,N_3936,N_3447);
or U5448 (N_5448,N_2370,N_2111);
nor U5449 (N_5449,N_2028,N_3712);
nor U5450 (N_5450,N_2452,N_3882);
nor U5451 (N_5451,N_3181,N_2569);
or U5452 (N_5452,N_2024,N_2277);
nor U5453 (N_5453,N_3742,N_3560);
and U5454 (N_5454,N_3903,N_3521);
nor U5455 (N_5455,N_3883,N_3793);
or U5456 (N_5456,N_3733,N_3233);
nand U5457 (N_5457,N_3455,N_3425);
nand U5458 (N_5458,N_3713,N_2149);
or U5459 (N_5459,N_2704,N_2053);
or U5460 (N_5460,N_2125,N_3244);
nand U5461 (N_5461,N_2754,N_2270);
nor U5462 (N_5462,N_3338,N_2806);
nand U5463 (N_5463,N_3009,N_2234);
nor U5464 (N_5464,N_2045,N_2474);
and U5465 (N_5465,N_2449,N_3688);
and U5466 (N_5466,N_3218,N_2099);
nand U5467 (N_5467,N_2375,N_3184);
or U5468 (N_5468,N_2130,N_3449);
nor U5469 (N_5469,N_3107,N_3383);
and U5470 (N_5470,N_2993,N_2194);
nand U5471 (N_5471,N_3240,N_2328);
nand U5472 (N_5472,N_2683,N_3536);
or U5473 (N_5473,N_3464,N_2862);
and U5474 (N_5474,N_3347,N_3529);
or U5475 (N_5475,N_3392,N_3917);
nor U5476 (N_5476,N_2876,N_2395);
or U5477 (N_5477,N_3950,N_2753);
nor U5478 (N_5478,N_3287,N_3452);
or U5479 (N_5479,N_3856,N_2101);
xor U5480 (N_5480,N_3854,N_2768);
nand U5481 (N_5481,N_3893,N_2207);
nand U5482 (N_5482,N_2330,N_3830);
and U5483 (N_5483,N_2710,N_2949);
nor U5484 (N_5484,N_3180,N_2206);
nor U5485 (N_5485,N_3689,N_2890);
and U5486 (N_5486,N_3217,N_2906);
or U5487 (N_5487,N_3582,N_3494);
nor U5488 (N_5488,N_2403,N_2157);
or U5489 (N_5489,N_2756,N_3708);
nor U5490 (N_5490,N_2771,N_2174);
and U5491 (N_5491,N_3357,N_3870);
nand U5492 (N_5492,N_2634,N_3168);
and U5493 (N_5493,N_2504,N_2020);
nor U5494 (N_5494,N_3736,N_2254);
and U5495 (N_5495,N_3812,N_2016);
or U5496 (N_5496,N_3716,N_3730);
or U5497 (N_5497,N_3296,N_3924);
and U5498 (N_5498,N_2999,N_3819);
or U5499 (N_5499,N_2055,N_3813);
xor U5500 (N_5500,N_2401,N_2028);
or U5501 (N_5501,N_2960,N_2012);
and U5502 (N_5502,N_2136,N_3273);
nor U5503 (N_5503,N_2141,N_2984);
nand U5504 (N_5504,N_2114,N_3179);
or U5505 (N_5505,N_3239,N_2020);
and U5506 (N_5506,N_2338,N_2585);
nand U5507 (N_5507,N_2811,N_2936);
nor U5508 (N_5508,N_2441,N_3197);
nor U5509 (N_5509,N_2072,N_2261);
or U5510 (N_5510,N_3968,N_3524);
nor U5511 (N_5511,N_2279,N_3695);
xnor U5512 (N_5512,N_2663,N_2351);
or U5513 (N_5513,N_2860,N_3872);
nand U5514 (N_5514,N_3480,N_3468);
nor U5515 (N_5515,N_3463,N_3943);
and U5516 (N_5516,N_3245,N_2803);
or U5517 (N_5517,N_3353,N_2905);
nor U5518 (N_5518,N_3325,N_3646);
or U5519 (N_5519,N_3560,N_2353);
or U5520 (N_5520,N_2754,N_2453);
nor U5521 (N_5521,N_3443,N_3672);
nor U5522 (N_5522,N_3456,N_2993);
and U5523 (N_5523,N_2840,N_3842);
and U5524 (N_5524,N_3716,N_2073);
and U5525 (N_5525,N_2353,N_2827);
nand U5526 (N_5526,N_2343,N_2816);
or U5527 (N_5527,N_2058,N_2542);
nand U5528 (N_5528,N_2176,N_2567);
or U5529 (N_5529,N_3090,N_3161);
nand U5530 (N_5530,N_3038,N_3072);
xnor U5531 (N_5531,N_3098,N_3042);
or U5532 (N_5532,N_2205,N_2845);
nor U5533 (N_5533,N_2874,N_3971);
nand U5534 (N_5534,N_2314,N_3643);
nor U5535 (N_5535,N_3929,N_2790);
nand U5536 (N_5536,N_2704,N_2547);
nand U5537 (N_5537,N_3200,N_3986);
or U5538 (N_5538,N_2292,N_2356);
nor U5539 (N_5539,N_3716,N_3214);
or U5540 (N_5540,N_2499,N_3735);
or U5541 (N_5541,N_2566,N_3607);
and U5542 (N_5542,N_3500,N_2560);
nand U5543 (N_5543,N_3528,N_3726);
nand U5544 (N_5544,N_3930,N_2389);
and U5545 (N_5545,N_2334,N_2346);
and U5546 (N_5546,N_3867,N_3744);
nand U5547 (N_5547,N_3515,N_2747);
and U5548 (N_5548,N_2265,N_3778);
nand U5549 (N_5549,N_3653,N_2824);
nand U5550 (N_5550,N_2075,N_3678);
and U5551 (N_5551,N_2885,N_3159);
nor U5552 (N_5552,N_3493,N_3935);
and U5553 (N_5553,N_3082,N_2169);
nand U5554 (N_5554,N_2335,N_3195);
nor U5555 (N_5555,N_3744,N_2931);
or U5556 (N_5556,N_3218,N_2796);
nand U5557 (N_5557,N_2290,N_2968);
nor U5558 (N_5558,N_3563,N_3840);
nand U5559 (N_5559,N_2069,N_2496);
or U5560 (N_5560,N_2778,N_3202);
and U5561 (N_5561,N_2971,N_3083);
nand U5562 (N_5562,N_2809,N_2306);
and U5563 (N_5563,N_3778,N_3304);
nor U5564 (N_5564,N_2180,N_2867);
or U5565 (N_5565,N_2605,N_2010);
and U5566 (N_5566,N_2680,N_3745);
nand U5567 (N_5567,N_2644,N_2360);
or U5568 (N_5568,N_2977,N_3373);
or U5569 (N_5569,N_3971,N_3335);
nand U5570 (N_5570,N_3123,N_3609);
and U5571 (N_5571,N_3025,N_2566);
nand U5572 (N_5572,N_3730,N_2991);
and U5573 (N_5573,N_3474,N_3368);
and U5574 (N_5574,N_3297,N_2646);
nor U5575 (N_5575,N_3764,N_3431);
or U5576 (N_5576,N_2284,N_3128);
nor U5577 (N_5577,N_3988,N_2830);
or U5578 (N_5578,N_2041,N_3579);
nand U5579 (N_5579,N_3955,N_3626);
or U5580 (N_5580,N_2798,N_3866);
and U5581 (N_5581,N_2739,N_3301);
and U5582 (N_5582,N_2794,N_3306);
nor U5583 (N_5583,N_3514,N_3977);
or U5584 (N_5584,N_3967,N_3786);
nand U5585 (N_5585,N_2725,N_2134);
and U5586 (N_5586,N_2430,N_2767);
nand U5587 (N_5587,N_3478,N_2090);
nand U5588 (N_5588,N_2023,N_3425);
nand U5589 (N_5589,N_2297,N_3809);
nor U5590 (N_5590,N_3164,N_2868);
nor U5591 (N_5591,N_3601,N_2139);
or U5592 (N_5592,N_2016,N_3305);
nor U5593 (N_5593,N_3416,N_3036);
xnor U5594 (N_5594,N_3436,N_3535);
nand U5595 (N_5595,N_3064,N_2261);
or U5596 (N_5596,N_2760,N_2019);
nor U5597 (N_5597,N_2961,N_2943);
nor U5598 (N_5598,N_3965,N_2405);
and U5599 (N_5599,N_3100,N_3661);
and U5600 (N_5600,N_3839,N_2881);
xnor U5601 (N_5601,N_2219,N_2817);
and U5602 (N_5602,N_3845,N_3043);
and U5603 (N_5603,N_2811,N_3975);
nor U5604 (N_5604,N_2932,N_2937);
nand U5605 (N_5605,N_3944,N_3767);
or U5606 (N_5606,N_3259,N_2088);
nor U5607 (N_5607,N_2674,N_3583);
or U5608 (N_5608,N_3387,N_2610);
nand U5609 (N_5609,N_3522,N_3179);
and U5610 (N_5610,N_2403,N_3649);
nand U5611 (N_5611,N_3653,N_2964);
or U5612 (N_5612,N_3681,N_2948);
nor U5613 (N_5613,N_2206,N_2975);
or U5614 (N_5614,N_3594,N_3406);
or U5615 (N_5615,N_2655,N_2579);
and U5616 (N_5616,N_3254,N_3670);
and U5617 (N_5617,N_2619,N_3448);
nand U5618 (N_5618,N_2363,N_2160);
and U5619 (N_5619,N_3050,N_3088);
nand U5620 (N_5620,N_2537,N_3431);
or U5621 (N_5621,N_3207,N_3184);
nand U5622 (N_5622,N_2279,N_3084);
nor U5623 (N_5623,N_3535,N_3231);
nand U5624 (N_5624,N_2549,N_2987);
or U5625 (N_5625,N_3629,N_2845);
nor U5626 (N_5626,N_3529,N_3116);
or U5627 (N_5627,N_3998,N_3118);
nor U5628 (N_5628,N_2438,N_2376);
nand U5629 (N_5629,N_2238,N_2179);
nor U5630 (N_5630,N_2798,N_3576);
and U5631 (N_5631,N_2591,N_2718);
or U5632 (N_5632,N_3617,N_2893);
nand U5633 (N_5633,N_3127,N_3374);
nor U5634 (N_5634,N_2175,N_3466);
xor U5635 (N_5635,N_3348,N_3456);
and U5636 (N_5636,N_3011,N_3322);
nor U5637 (N_5637,N_3341,N_2181);
xor U5638 (N_5638,N_3594,N_2954);
nand U5639 (N_5639,N_3101,N_2489);
nand U5640 (N_5640,N_2590,N_2886);
or U5641 (N_5641,N_3480,N_2468);
nor U5642 (N_5642,N_3379,N_3266);
nor U5643 (N_5643,N_2929,N_3858);
and U5644 (N_5644,N_2750,N_3765);
or U5645 (N_5645,N_2852,N_3112);
and U5646 (N_5646,N_3128,N_3974);
and U5647 (N_5647,N_2250,N_3446);
nand U5648 (N_5648,N_3691,N_2560);
nand U5649 (N_5649,N_3117,N_3545);
or U5650 (N_5650,N_2867,N_2794);
and U5651 (N_5651,N_2410,N_2133);
nand U5652 (N_5652,N_2964,N_2072);
or U5653 (N_5653,N_3242,N_2158);
nand U5654 (N_5654,N_2927,N_2263);
nand U5655 (N_5655,N_2444,N_3218);
nand U5656 (N_5656,N_3645,N_2706);
nor U5657 (N_5657,N_3090,N_3184);
or U5658 (N_5658,N_3548,N_3946);
or U5659 (N_5659,N_3959,N_3908);
or U5660 (N_5660,N_3580,N_2035);
nor U5661 (N_5661,N_2078,N_2455);
and U5662 (N_5662,N_2761,N_3777);
and U5663 (N_5663,N_2907,N_3239);
nor U5664 (N_5664,N_3511,N_3125);
nand U5665 (N_5665,N_2049,N_3586);
nor U5666 (N_5666,N_3483,N_3157);
or U5667 (N_5667,N_3144,N_3357);
nor U5668 (N_5668,N_2652,N_3700);
nand U5669 (N_5669,N_3974,N_3451);
or U5670 (N_5670,N_3343,N_3706);
nand U5671 (N_5671,N_3536,N_2517);
or U5672 (N_5672,N_2159,N_3252);
nor U5673 (N_5673,N_3823,N_2099);
nor U5674 (N_5674,N_2399,N_3648);
nand U5675 (N_5675,N_2172,N_3349);
and U5676 (N_5676,N_3649,N_2525);
or U5677 (N_5677,N_2327,N_2751);
nor U5678 (N_5678,N_2975,N_3912);
nor U5679 (N_5679,N_3509,N_3916);
nand U5680 (N_5680,N_2500,N_2201);
nand U5681 (N_5681,N_2657,N_3520);
and U5682 (N_5682,N_3113,N_3171);
or U5683 (N_5683,N_3823,N_3247);
nor U5684 (N_5684,N_3414,N_3012);
nand U5685 (N_5685,N_3007,N_2459);
or U5686 (N_5686,N_3217,N_2373);
or U5687 (N_5687,N_2549,N_2911);
or U5688 (N_5688,N_3964,N_2815);
nor U5689 (N_5689,N_3444,N_2091);
and U5690 (N_5690,N_3729,N_2425);
nor U5691 (N_5691,N_3066,N_3491);
or U5692 (N_5692,N_2937,N_3786);
or U5693 (N_5693,N_3444,N_3482);
nand U5694 (N_5694,N_3198,N_3506);
nand U5695 (N_5695,N_3122,N_3219);
or U5696 (N_5696,N_2908,N_3148);
and U5697 (N_5697,N_3865,N_3148);
and U5698 (N_5698,N_3388,N_3532);
nand U5699 (N_5699,N_3084,N_3732);
nand U5700 (N_5700,N_2975,N_3280);
or U5701 (N_5701,N_2027,N_3926);
nor U5702 (N_5702,N_3039,N_3569);
nand U5703 (N_5703,N_3019,N_2651);
or U5704 (N_5704,N_2021,N_3797);
nor U5705 (N_5705,N_3750,N_3592);
and U5706 (N_5706,N_3134,N_2576);
nand U5707 (N_5707,N_2836,N_3349);
nor U5708 (N_5708,N_3123,N_2933);
or U5709 (N_5709,N_3288,N_2121);
nor U5710 (N_5710,N_3667,N_3999);
nor U5711 (N_5711,N_2777,N_2621);
or U5712 (N_5712,N_2405,N_3806);
nand U5713 (N_5713,N_2156,N_2176);
nand U5714 (N_5714,N_2991,N_2317);
nor U5715 (N_5715,N_3719,N_3688);
or U5716 (N_5716,N_2801,N_3293);
nand U5717 (N_5717,N_2158,N_3364);
nor U5718 (N_5718,N_3209,N_3761);
or U5719 (N_5719,N_2546,N_2522);
nor U5720 (N_5720,N_3637,N_2634);
nor U5721 (N_5721,N_3225,N_2790);
or U5722 (N_5722,N_3288,N_3933);
nor U5723 (N_5723,N_3665,N_2392);
or U5724 (N_5724,N_3844,N_3750);
nor U5725 (N_5725,N_2519,N_2617);
nor U5726 (N_5726,N_3021,N_3539);
nor U5727 (N_5727,N_2783,N_2219);
xor U5728 (N_5728,N_3956,N_3469);
xor U5729 (N_5729,N_3061,N_3769);
nand U5730 (N_5730,N_2447,N_2587);
nand U5731 (N_5731,N_3254,N_3697);
nor U5732 (N_5732,N_2908,N_3243);
nand U5733 (N_5733,N_3722,N_3442);
or U5734 (N_5734,N_2068,N_3715);
or U5735 (N_5735,N_2036,N_2185);
nor U5736 (N_5736,N_2426,N_2649);
and U5737 (N_5737,N_3971,N_2506);
or U5738 (N_5738,N_2540,N_3895);
xor U5739 (N_5739,N_2287,N_2570);
nor U5740 (N_5740,N_2118,N_3988);
or U5741 (N_5741,N_2939,N_3970);
nand U5742 (N_5742,N_3503,N_2680);
and U5743 (N_5743,N_3482,N_3408);
nor U5744 (N_5744,N_2020,N_3920);
nor U5745 (N_5745,N_2627,N_3062);
or U5746 (N_5746,N_3396,N_2797);
nor U5747 (N_5747,N_2489,N_2940);
nor U5748 (N_5748,N_3798,N_2519);
and U5749 (N_5749,N_3240,N_3574);
and U5750 (N_5750,N_3033,N_2368);
and U5751 (N_5751,N_3301,N_3798);
nand U5752 (N_5752,N_3090,N_2104);
nand U5753 (N_5753,N_2673,N_2306);
nand U5754 (N_5754,N_3607,N_2535);
nand U5755 (N_5755,N_3364,N_2815);
and U5756 (N_5756,N_2889,N_2532);
nor U5757 (N_5757,N_3475,N_2974);
nand U5758 (N_5758,N_2563,N_2181);
and U5759 (N_5759,N_3803,N_3348);
or U5760 (N_5760,N_2681,N_2631);
or U5761 (N_5761,N_2360,N_3643);
and U5762 (N_5762,N_2366,N_3864);
or U5763 (N_5763,N_2396,N_2525);
xnor U5764 (N_5764,N_2733,N_3025);
nand U5765 (N_5765,N_3291,N_2033);
xor U5766 (N_5766,N_3713,N_3030);
nand U5767 (N_5767,N_3504,N_2950);
nor U5768 (N_5768,N_2445,N_2737);
nor U5769 (N_5769,N_3861,N_2879);
and U5770 (N_5770,N_3847,N_2383);
nor U5771 (N_5771,N_2417,N_3954);
or U5772 (N_5772,N_2497,N_3691);
or U5773 (N_5773,N_3366,N_2666);
or U5774 (N_5774,N_2853,N_2147);
and U5775 (N_5775,N_3019,N_2184);
and U5776 (N_5776,N_2472,N_2724);
nor U5777 (N_5777,N_2787,N_2856);
and U5778 (N_5778,N_2905,N_3766);
nand U5779 (N_5779,N_2796,N_3987);
nor U5780 (N_5780,N_2104,N_3793);
and U5781 (N_5781,N_3400,N_2442);
and U5782 (N_5782,N_2069,N_2030);
or U5783 (N_5783,N_3151,N_2604);
and U5784 (N_5784,N_3497,N_2728);
or U5785 (N_5785,N_3575,N_3262);
or U5786 (N_5786,N_2424,N_2101);
nand U5787 (N_5787,N_2498,N_2580);
or U5788 (N_5788,N_2824,N_2592);
nor U5789 (N_5789,N_3186,N_2669);
nor U5790 (N_5790,N_3623,N_3597);
or U5791 (N_5791,N_2299,N_2463);
nor U5792 (N_5792,N_3851,N_2189);
nand U5793 (N_5793,N_3586,N_2889);
nand U5794 (N_5794,N_3199,N_2899);
xor U5795 (N_5795,N_2883,N_2586);
or U5796 (N_5796,N_2227,N_3432);
and U5797 (N_5797,N_3588,N_3252);
nand U5798 (N_5798,N_3237,N_3507);
or U5799 (N_5799,N_3284,N_3473);
nor U5800 (N_5800,N_2948,N_3856);
nand U5801 (N_5801,N_2932,N_3529);
nor U5802 (N_5802,N_2566,N_2575);
nand U5803 (N_5803,N_3411,N_2602);
nor U5804 (N_5804,N_3056,N_2780);
or U5805 (N_5805,N_3807,N_2705);
nand U5806 (N_5806,N_2079,N_2153);
or U5807 (N_5807,N_2233,N_3846);
nor U5808 (N_5808,N_2892,N_3141);
nand U5809 (N_5809,N_2096,N_2730);
and U5810 (N_5810,N_3540,N_3624);
nand U5811 (N_5811,N_2249,N_3050);
or U5812 (N_5812,N_2147,N_2782);
nor U5813 (N_5813,N_2936,N_2226);
nand U5814 (N_5814,N_2514,N_2622);
and U5815 (N_5815,N_3392,N_2032);
and U5816 (N_5816,N_2380,N_3768);
and U5817 (N_5817,N_2002,N_2193);
and U5818 (N_5818,N_3252,N_3228);
and U5819 (N_5819,N_2576,N_2986);
nand U5820 (N_5820,N_3056,N_3005);
nor U5821 (N_5821,N_2375,N_3661);
nand U5822 (N_5822,N_3026,N_3198);
or U5823 (N_5823,N_2867,N_3794);
nand U5824 (N_5824,N_3385,N_3216);
or U5825 (N_5825,N_2084,N_3096);
nand U5826 (N_5826,N_3208,N_2188);
and U5827 (N_5827,N_2305,N_3826);
nand U5828 (N_5828,N_2778,N_2307);
or U5829 (N_5829,N_2638,N_2017);
and U5830 (N_5830,N_3263,N_3604);
or U5831 (N_5831,N_3826,N_3979);
nand U5832 (N_5832,N_2415,N_3825);
nor U5833 (N_5833,N_2876,N_2008);
nand U5834 (N_5834,N_2072,N_2422);
xor U5835 (N_5835,N_2567,N_3752);
or U5836 (N_5836,N_3315,N_3441);
or U5837 (N_5837,N_2547,N_3048);
and U5838 (N_5838,N_3074,N_2076);
nand U5839 (N_5839,N_3713,N_3267);
nand U5840 (N_5840,N_2359,N_2519);
or U5841 (N_5841,N_2059,N_3071);
nand U5842 (N_5842,N_2367,N_3600);
and U5843 (N_5843,N_3128,N_3666);
and U5844 (N_5844,N_3723,N_3061);
nand U5845 (N_5845,N_2111,N_3891);
or U5846 (N_5846,N_2108,N_3452);
nand U5847 (N_5847,N_3024,N_3667);
or U5848 (N_5848,N_3664,N_2676);
nand U5849 (N_5849,N_3664,N_3099);
or U5850 (N_5850,N_2183,N_3590);
nor U5851 (N_5851,N_3023,N_3155);
nand U5852 (N_5852,N_2509,N_2415);
and U5853 (N_5853,N_3612,N_2518);
nand U5854 (N_5854,N_3606,N_2126);
or U5855 (N_5855,N_3152,N_2701);
or U5856 (N_5856,N_3235,N_3858);
xnor U5857 (N_5857,N_3610,N_2505);
or U5858 (N_5858,N_3715,N_3362);
or U5859 (N_5859,N_3989,N_3010);
nor U5860 (N_5860,N_3489,N_3845);
or U5861 (N_5861,N_3253,N_3428);
and U5862 (N_5862,N_2077,N_3637);
or U5863 (N_5863,N_3688,N_3437);
nor U5864 (N_5864,N_2865,N_3663);
nor U5865 (N_5865,N_3372,N_2017);
nand U5866 (N_5866,N_2372,N_2999);
or U5867 (N_5867,N_3474,N_2287);
nand U5868 (N_5868,N_2725,N_2708);
nand U5869 (N_5869,N_2067,N_2946);
and U5870 (N_5870,N_2844,N_3565);
or U5871 (N_5871,N_3703,N_3367);
or U5872 (N_5872,N_3063,N_3324);
or U5873 (N_5873,N_2171,N_2291);
or U5874 (N_5874,N_2785,N_3351);
and U5875 (N_5875,N_2435,N_2098);
xnor U5876 (N_5876,N_2324,N_2337);
or U5877 (N_5877,N_2198,N_3709);
nor U5878 (N_5878,N_2730,N_2552);
or U5879 (N_5879,N_2306,N_2321);
nand U5880 (N_5880,N_2035,N_3729);
or U5881 (N_5881,N_3365,N_2476);
nand U5882 (N_5882,N_2467,N_2166);
nor U5883 (N_5883,N_3428,N_3529);
or U5884 (N_5884,N_3965,N_2225);
nor U5885 (N_5885,N_2265,N_2757);
or U5886 (N_5886,N_3986,N_2859);
and U5887 (N_5887,N_3602,N_2192);
nand U5888 (N_5888,N_3789,N_2134);
and U5889 (N_5889,N_3995,N_3823);
or U5890 (N_5890,N_3960,N_3378);
and U5891 (N_5891,N_3782,N_3006);
and U5892 (N_5892,N_3022,N_2046);
or U5893 (N_5893,N_3492,N_2718);
or U5894 (N_5894,N_2538,N_3348);
and U5895 (N_5895,N_3028,N_2755);
and U5896 (N_5896,N_3764,N_3620);
or U5897 (N_5897,N_3510,N_3749);
nor U5898 (N_5898,N_3654,N_2388);
nand U5899 (N_5899,N_3903,N_2087);
nor U5900 (N_5900,N_3448,N_2787);
or U5901 (N_5901,N_3305,N_2950);
or U5902 (N_5902,N_3191,N_3158);
and U5903 (N_5903,N_2305,N_2267);
and U5904 (N_5904,N_2555,N_3451);
xor U5905 (N_5905,N_2241,N_2246);
and U5906 (N_5906,N_2256,N_3729);
or U5907 (N_5907,N_2704,N_3727);
or U5908 (N_5908,N_3729,N_2037);
and U5909 (N_5909,N_3943,N_3782);
nor U5910 (N_5910,N_2831,N_3468);
nand U5911 (N_5911,N_2536,N_3012);
nand U5912 (N_5912,N_2477,N_3664);
nor U5913 (N_5913,N_3872,N_2390);
or U5914 (N_5914,N_3713,N_3994);
nor U5915 (N_5915,N_2718,N_3674);
nor U5916 (N_5916,N_2590,N_2339);
or U5917 (N_5917,N_2021,N_3624);
or U5918 (N_5918,N_3401,N_3178);
or U5919 (N_5919,N_3647,N_3979);
or U5920 (N_5920,N_3548,N_3002);
xnor U5921 (N_5921,N_2173,N_2193);
nand U5922 (N_5922,N_2169,N_3688);
nand U5923 (N_5923,N_3242,N_3116);
xor U5924 (N_5924,N_2573,N_3654);
or U5925 (N_5925,N_2899,N_2518);
nand U5926 (N_5926,N_3351,N_3538);
or U5927 (N_5927,N_2440,N_3944);
nand U5928 (N_5928,N_3515,N_3290);
and U5929 (N_5929,N_3201,N_2786);
nor U5930 (N_5930,N_3786,N_2686);
nand U5931 (N_5931,N_2217,N_2229);
and U5932 (N_5932,N_2659,N_3702);
xnor U5933 (N_5933,N_2245,N_2517);
nand U5934 (N_5934,N_3136,N_3121);
nor U5935 (N_5935,N_3457,N_2962);
nor U5936 (N_5936,N_3728,N_2579);
or U5937 (N_5937,N_2606,N_2881);
and U5938 (N_5938,N_2155,N_2620);
or U5939 (N_5939,N_2183,N_2523);
nand U5940 (N_5940,N_3313,N_2148);
and U5941 (N_5941,N_2139,N_2746);
xor U5942 (N_5942,N_3548,N_2853);
nor U5943 (N_5943,N_2935,N_2803);
or U5944 (N_5944,N_2043,N_2810);
and U5945 (N_5945,N_2930,N_3440);
and U5946 (N_5946,N_2517,N_2569);
nand U5947 (N_5947,N_3323,N_3713);
nor U5948 (N_5948,N_2977,N_2878);
nor U5949 (N_5949,N_3623,N_3780);
or U5950 (N_5950,N_3175,N_2383);
nor U5951 (N_5951,N_2526,N_3661);
and U5952 (N_5952,N_3650,N_3192);
or U5953 (N_5953,N_2176,N_2934);
nand U5954 (N_5954,N_2633,N_2715);
nand U5955 (N_5955,N_3067,N_3220);
nor U5956 (N_5956,N_2087,N_2416);
or U5957 (N_5957,N_2119,N_3062);
nor U5958 (N_5958,N_3338,N_2682);
nand U5959 (N_5959,N_3800,N_2527);
nand U5960 (N_5960,N_3487,N_2344);
or U5961 (N_5961,N_2526,N_2722);
nor U5962 (N_5962,N_3171,N_3234);
and U5963 (N_5963,N_2834,N_2511);
or U5964 (N_5964,N_2958,N_2652);
nand U5965 (N_5965,N_3074,N_2179);
nor U5966 (N_5966,N_2848,N_2790);
or U5967 (N_5967,N_3941,N_3755);
or U5968 (N_5968,N_2259,N_3202);
or U5969 (N_5969,N_3142,N_3998);
nand U5970 (N_5970,N_3256,N_3448);
and U5971 (N_5971,N_2179,N_2565);
or U5972 (N_5972,N_3739,N_2164);
or U5973 (N_5973,N_2012,N_2019);
and U5974 (N_5974,N_2606,N_2415);
or U5975 (N_5975,N_3703,N_3479);
and U5976 (N_5976,N_3046,N_3219);
nand U5977 (N_5977,N_3701,N_3268);
nand U5978 (N_5978,N_2210,N_2951);
and U5979 (N_5979,N_3211,N_2074);
and U5980 (N_5980,N_2411,N_3507);
and U5981 (N_5981,N_3843,N_2141);
nand U5982 (N_5982,N_2861,N_3657);
nor U5983 (N_5983,N_2668,N_3399);
nor U5984 (N_5984,N_3178,N_2291);
nor U5985 (N_5985,N_2137,N_3936);
nor U5986 (N_5986,N_3851,N_2814);
or U5987 (N_5987,N_2286,N_2400);
nand U5988 (N_5988,N_2876,N_2110);
and U5989 (N_5989,N_2062,N_3521);
nand U5990 (N_5990,N_3914,N_2445);
or U5991 (N_5991,N_3114,N_2595);
or U5992 (N_5992,N_3928,N_3046);
or U5993 (N_5993,N_3824,N_3032);
nor U5994 (N_5994,N_3372,N_3543);
nand U5995 (N_5995,N_3993,N_2890);
nand U5996 (N_5996,N_3344,N_3504);
or U5997 (N_5997,N_2364,N_3565);
or U5998 (N_5998,N_2118,N_2602);
nor U5999 (N_5999,N_2411,N_2227);
or U6000 (N_6000,N_4714,N_5430);
and U6001 (N_6001,N_4785,N_4839);
nor U6002 (N_6002,N_4347,N_4343);
and U6003 (N_6003,N_5707,N_4331);
nand U6004 (N_6004,N_5719,N_5669);
nand U6005 (N_6005,N_4588,N_4288);
nor U6006 (N_6006,N_5378,N_5713);
and U6007 (N_6007,N_4648,N_4652);
nor U6008 (N_6008,N_5164,N_5167);
and U6009 (N_6009,N_4927,N_5860);
or U6010 (N_6010,N_4622,N_5774);
nand U6011 (N_6011,N_5037,N_4938);
nand U6012 (N_6012,N_5304,N_5036);
or U6013 (N_6013,N_5629,N_4110);
or U6014 (N_6014,N_4464,N_5355);
nand U6015 (N_6015,N_5313,N_4923);
nand U6016 (N_6016,N_4607,N_4140);
or U6017 (N_6017,N_4612,N_5300);
or U6018 (N_6018,N_4339,N_5877);
or U6019 (N_6019,N_4273,N_4935);
and U6020 (N_6020,N_4005,N_5203);
and U6021 (N_6021,N_5471,N_5958);
nand U6022 (N_6022,N_5820,N_5563);
and U6023 (N_6023,N_5485,N_4354);
and U6024 (N_6024,N_5571,N_4081);
xnor U6025 (N_6025,N_5648,N_5805);
and U6026 (N_6026,N_5269,N_5800);
nand U6027 (N_6027,N_5038,N_4779);
and U6028 (N_6028,N_5978,N_5219);
or U6029 (N_6029,N_5930,N_4497);
nand U6030 (N_6030,N_4346,N_5489);
or U6031 (N_6031,N_4492,N_4344);
or U6032 (N_6032,N_4787,N_4133);
nand U6033 (N_6033,N_4155,N_4127);
nand U6034 (N_6034,N_5929,N_4739);
or U6035 (N_6035,N_4585,N_4771);
or U6036 (N_6036,N_5284,N_5566);
nand U6037 (N_6037,N_4016,N_5866);
or U6038 (N_6038,N_5375,N_4035);
nand U6039 (N_6039,N_5808,N_4809);
and U6040 (N_6040,N_4191,N_5701);
nand U6041 (N_6041,N_5690,N_4039);
or U6042 (N_6042,N_5322,N_5951);
nand U6043 (N_6043,N_4093,N_4091);
nand U6044 (N_6044,N_5308,N_5888);
nand U6045 (N_6045,N_5714,N_4798);
and U6046 (N_6046,N_5814,N_5840);
or U6047 (N_6047,N_4524,N_4724);
or U6048 (N_6048,N_5613,N_5370);
nor U6049 (N_6049,N_5383,N_5542);
nor U6050 (N_6050,N_5658,N_5672);
or U6051 (N_6051,N_4842,N_4527);
nand U6052 (N_6052,N_5551,N_4246);
nand U6053 (N_6053,N_5768,N_5532);
nor U6054 (N_6054,N_4028,N_5356);
or U6055 (N_6055,N_4706,N_5041);
nand U6056 (N_6056,N_5557,N_4632);
nor U6057 (N_6057,N_4022,N_4726);
and U6058 (N_6058,N_5806,N_4117);
nand U6059 (N_6059,N_4529,N_5108);
nand U6060 (N_6060,N_5664,N_5520);
nand U6061 (N_6061,N_4708,N_4631);
nand U6062 (N_6062,N_4310,N_5169);
nor U6063 (N_6063,N_4330,N_4767);
nand U6064 (N_6064,N_4291,N_5140);
or U6065 (N_6065,N_4534,N_5055);
or U6066 (N_6066,N_5801,N_5425);
or U6067 (N_6067,N_5926,N_4223);
nor U6068 (N_6068,N_4718,N_5955);
and U6069 (N_6069,N_4009,N_5757);
or U6070 (N_6070,N_5773,N_4912);
nand U6071 (N_6071,N_4734,N_4198);
or U6072 (N_6072,N_5883,N_5467);
nor U6073 (N_6073,N_4851,N_4523);
and U6074 (N_6074,N_5004,N_4104);
or U6075 (N_6075,N_5908,N_5072);
or U6076 (N_6076,N_4516,N_4882);
nand U6077 (N_6077,N_5096,N_5528);
or U6078 (N_6078,N_4214,N_4545);
nand U6079 (N_6079,N_5366,N_5755);
and U6080 (N_6080,N_4557,N_4922);
nor U6081 (N_6081,N_5770,N_5101);
or U6082 (N_6082,N_4669,N_4797);
nand U6083 (N_6083,N_4159,N_4293);
and U6084 (N_6084,N_4551,N_4967);
or U6085 (N_6085,N_4504,N_5438);
nand U6086 (N_6086,N_4975,N_4627);
nor U6087 (N_6087,N_4898,N_4827);
nand U6088 (N_6088,N_4889,N_4287);
nand U6089 (N_6089,N_4532,N_4619);
and U6090 (N_6090,N_4074,N_4983);
and U6091 (N_6091,N_4556,N_4378);
nor U6092 (N_6092,N_5148,N_5406);
xor U6093 (N_6093,N_4752,N_4602);
or U6094 (N_6094,N_4984,N_5711);
and U6095 (N_6095,N_4618,N_5367);
nand U6096 (N_6096,N_5069,N_5143);
and U6097 (N_6097,N_5116,N_4033);
and U6098 (N_6098,N_5689,N_5364);
or U6099 (N_6099,N_5581,N_4704);
nand U6100 (N_6100,N_5631,N_4826);
and U6101 (N_6101,N_4371,N_5585);
nand U6102 (N_6102,N_4232,N_5600);
nand U6103 (N_6103,N_4899,N_5057);
nor U6104 (N_6104,N_4375,N_4334);
xnor U6105 (N_6105,N_5330,N_5226);
nor U6106 (N_6106,N_5099,N_5081);
nor U6107 (N_6107,N_5392,N_4462);
nor U6108 (N_6108,N_5750,N_4494);
nand U6109 (N_6109,N_5797,N_4693);
nor U6110 (N_6110,N_5190,N_5744);
nor U6111 (N_6111,N_5176,N_5098);
or U6112 (N_6112,N_5128,N_4073);
and U6113 (N_6113,N_5079,N_4628);
nand U6114 (N_6114,N_4459,N_5174);
and U6115 (N_6115,N_4136,N_4289);
or U6116 (N_6116,N_5545,N_5197);
and U6117 (N_6117,N_4226,N_5454);
nor U6118 (N_6118,N_5513,N_5087);
nand U6119 (N_6119,N_5863,N_4461);
or U6120 (N_6120,N_5060,N_4397);
nand U6121 (N_6121,N_5256,N_5379);
or U6122 (N_6122,N_5646,N_4380);
nor U6123 (N_6123,N_5158,N_5180);
and U6124 (N_6124,N_4796,N_4634);
nor U6125 (N_6125,N_5712,N_4626);
nor U6126 (N_6126,N_5018,N_4653);
nor U6127 (N_6127,N_5335,N_5246);
nand U6128 (N_6128,N_4003,N_4940);
or U6129 (N_6129,N_4629,N_5997);
nor U6130 (N_6130,N_5278,N_5595);
nand U6131 (N_6131,N_4620,N_5780);
nand U6132 (N_6132,N_5334,N_5062);
and U6133 (N_6133,N_4259,N_5977);
nand U6134 (N_6134,N_5051,N_4871);
xor U6135 (N_6135,N_4408,N_5804);
nor U6136 (N_6136,N_4055,N_5608);
nand U6137 (N_6137,N_4624,N_4054);
nand U6138 (N_6138,N_4472,N_5100);
nand U6139 (N_6139,N_5695,N_4132);
and U6140 (N_6140,N_4245,N_4357);
nand U6141 (N_6141,N_5259,N_4107);
and U6142 (N_6142,N_5498,N_4500);
and U6143 (N_6143,N_4373,N_4743);
and U6144 (N_6144,N_5594,N_4420);
nand U6145 (N_6145,N_5746,N_4828);
nor U6146 (N_6146,N_4543,N_5500);
nor U6147 (N_6147,N_4526,N_4006);
nand U6148 (N_6148,N_5045,N_5453);
or U6149 (N_6149,N_4419,N_5654);
nand U6150 (N_6150,N_5042,N_4998);
nor U6151 (N_6151,N_5716,N_5272);
and U6152 (N_6152,N_5136,N_5227);
and U6153 (N_6153,N_4309,N_4803);
nor U6154 (N_6154,N_5832,N_5775);
and U6155 (N_6155,N_5647,N_5080);
and U6156 (N_6156,N_4192,N_5418);
xnor U6157 (N_6157,N_5010,N_5767);
or U6158 (N_6158,N_4158,N_5465);
nor U6159 (N_6159,N_5861,N_4587);
nand U6160 (N_6160,N_4429,N_4021);
nor U6161 (N_6161,N_4699,N_4918);
and U6162 (N_6162,N_4163,N_4831);
or U6163 (N_6163,N_4732,N_4646);
nand U6164 (N_6164,N_5276,N_5828);
or U6165 (N_6165,N_5992,N_4834);
and U6166 (N_6166,N_4453,N_4616);
nor U6167 (N_6167,N_4554,N_4980);
and U6168 (N_6168,N_5573,N_4134);
and U6169 (N_6169,N_4097,N_4987);
nand U6170 (N_6170,N_4361,N_5807);
and U6171 (N_6171,N_5986,N_4057);
or U6172 (N_6172,N_4592,N_5535);
nand U6173 (N_6173,N_5466,N_4236);
or U6174 (N_6174,N_5231,N_5293);
and U6175 (N_6175,N_4234,N_5050);
nand U6176 (N_6176,N_5688,N_4954);
and U6177 (N_6177,N_4180,N_5907);
and U6178 (N_6178,N_4445,N_5415);
and U6179 (N_6179,N_5939,N_4594);
nand U6180 (N_6180,N_5961,N_5186);
nor U6181 (N_6181,N_5771,N_5184);
or U6182 (N_6182,N_4308,N_4555);
nand U6183 (N_6183,N_5589,N_5312);
and U6184 (N_6184,N_5914,N_4352);
nand U6185 (N_6185,N_5615,N_5870);
and U6186 (N_6186,N_4569,N_4893);
or U6187 (N_6187,N_5338,N_5554);
nor U6188 (N_6188,N_5374,N_4399);
or U6189 (N_6189,N_4559,N_4151);
or U6190 (N_6190,N_4738,N_5550);
nand U6191 (N_6191,N_4270,N_4836);
and U6192 (N_6192,N_4422,N_4640);
nor U6193 (N_6193,N_5680,N_4683);
nand U6194 (N_6194,N_5791,N_5628);
and U6195 (N_6195,N_5816,N_4274);
or U6196 (N_6196,N_5792,N_5074);
nor U6197 (N_6197,N_5603,N_5657);
nor U6198 (N_6198,N_5909,N_5781);
nand U6199 (N_6199,N_5030,N_5213);
nand U6200 (N_6200,N_4802,N_4471);
xor U6201 (N_6201,N_5091,N_5985);
nor U6202 (N_6202,N_4338,N_5687);
and U6203 (N_6203,N_5604,N_4013);
nand U6204 (N_6204,N_4099,N_4239);
nor U6205 (N_6205,N_5922,N_4024);
nor U6206 (N_6206,N_5845,N_5844);
nor U6207 (N_6207,N_4290,N_5145);
or U6208 (N_6208,N_5023,N_5422);
and U6209 (N_6209,N_4037,N_5071);
or U6210 (N_6210,N_5541,N_5154);
and U6211 (N_6211,N_5731,N_4892);
nand U6212 (N_6212,N_5979,N_5280);
or U6213 (N_6213,N_4835,N_4867);
or U6214 (N_6214,N_4038,N_5857);
and U6215 (N_6215,N_5084,N_5409);
or U6216 (N_6216,N_4657,N_4218);
nor U6217 (N_6217,N_5377,N_4415);
and U6218 (N_6218,N_5590,N_5878);
nand U6219 (N_6219,N_4586,N_4979);
and U6220 (N_6220,N_4335,N_5987);
nor U6221 (N_6221,N_5682,N_5401);
nor U6222 (N_6222,N_5956,N_4482);
or U6223 (N_6223,N_5141,N_4508);
and U6224 (N_6224,N_4926,N_4207);
and U6225 (N_6225,N_5205,N_4790);
and U6226 (N_6226,N_4368,N_4515);
nor U6227 (N_6227,N_5691,N_5325);
nor U6228 (N_6228,N_5812,N_4059);
and U6229 (N_6229,N_4072,N_5214);
and U6230 (N_6230,N_5880,N_4930);
and U6231 (N_6231,N_4649,N_4799);
and U6232 (N_6232,N_5747,N_5763);
and U6233 (N_6233,N_4503,N_4105);
nor U6234 (N_6234,N_5830,N_5717);
or U6235 (N_6235,N_5009,N_5484);
or U6236 (N_6236,N_4235,N_4436);
nand U6237 (N_6237,N_4682,N_4131);
nand U6238 (N_6238,N_5028,N_5432);
nor U6239 (N_6239,N_4934,N_4004);
or U6240 (N_6240,N_5522,N_4014);
and U6241 (N_6241,N_4553,N_5292);
or U6242 (N_6242,N_4574,N_4604);
and U6243 (N_6243,N_5821,N_5361);
nand U6244 (N_6244,N_4919,N_5833);
nand U6245 (N_6245,N_5501,N_5889);
or U6246 (N_6246,N_5358,N_5097);
nor U6247 (N_6247,N_5988,N_4583);
and U6248 (N_6248,N_5078,N_4880);
or U6249 (N_6249,N_4801,N_4036);
or U6250 (N_6250,N_5105,N_4905);
or U6251 (N_6251,N_5633,N_4100);
nor U6252 (N_6252,N_5734,N_5350);
xor U6253 (N_6253,N_5753,N_4027);
nor U6254 (N_6254,N_5049,N_4617);
nor U6255 (N_6255,N_4056,N_5480);
and U6256 (N_6256,N_5663,N_4550);
nor U6257 (N_6257,N_5412,N_5061);
nand U6258 (N_6258,N_4053,N_5200);
nor U6259 (N_6259,N_4991,N_4098);
nor U6260 (N_6260,N_4625,N_5346);
and U6261 (N_6261,N_4662,N_5918);
and U6262 (N_6262,N_4161,N_5574);
nand U6263 (N_6263,N_5721,N_5188);
nand U6264 (N_6264,N_4818,N_4731);
and U6265 (N_6265,N_4176,N_5965);
and U6266 (N_6266,N_4552,N_5611);
nand U6267 (N_6267,N_5443,N_5228);
nor U6268 (N_6268,N_4753,N_4479);
xor U6269 (N_6269,N_4026,N_5900);
or U6270 (N_6270,N_5189,N_5389);
nand U6271 (N_6271,N_5423,N_4489);
and U6272 (N_6272,N_4391,N_5811);
or U6273 (N_6273,N_5504,N_5211);
and U6274 (N_6274,N_5351,N_4392);
or U6275 (N_6275,N_5268,N_5578);
and U6276 (N_6276,N_4965,N_5540);
nor U6277 (N_6277,N_4725,N_4389);
nor U6278 (N_6278,N_4883,N_5207);
nor U6279 (N_6279,N_4441,N_4242);
and U6280 (N_6280,N_4763,N_5488);
nor U6281 (N_6281,N_5014,N_5619);
nand U6282 (N_6282,N_4456,N_4447);
and U6283 (N_6283,N_4253,N_5279);
or U6284 (N_6284,N_5469,N_5923);
nand U6285 (N_6285,N_4486,N_5837);
or U6286 (N_6286,N_5984,N_5602);
and U6287 (N_6287,N_4457,N_5076);
or U6288 (N_6288,N_5368,N_5156);
nand U6289 (N_6289,N_4491,N_5973);
nor U6290 (N_6290,N_5130,N_4008);
nand U6291 (N_6291,N_4558,N_5614);
nor U6292 (N_6292,N_5135,N_5494);
or U6293 (N_6293,N_5790,N_5427);
xor U6294 (N_6294,N_5170,N_5435);
nor U6295 (N_6295,N_5990,N_4316);
or U6296 (N_6296,N_4638,N_4584);
nor U6297 (N_6297,N_5847,N_5348);
nand U6298 (N_6298,N_4359,N_4194);
nor U6299 (N_6299,N_4473,N_5727);
nand U6300 (N_6300,N_4852,N_5303);
nand U6301 (N_6301,N_4804,N_5787);
nor U6302 (N_6302,N_4139,N_4522);
nor U6303 (N_6303,N_5904,N_4034);
nand U6304 (N_6304,N_5343,N_4351);
nor U6305 (N_6305,N_4814,N_5548);
and U6306 (N_6306,N_4512,N_5886);
or U6307 (N_6307,N_5618,N_4830);
and U6308 (N_6308,N_4737,N_5575);
nor U6309 (N_6309,N_4147,N_4668);
and U6310 (N_6310,N_5533,N_4568);
nor U6311 (N_6311,N_5458,N_4513);
nor U6312 (N_6312,N_4044,N_4854);
and U6313 (N_6313,N_4149,N_5094);
and U6314 (N_6314,N_5996,N_5569);
and U6315 (N_6315,N_4621,N_4789);
nor U6316 (N_6316,N_4781,N_5623);
or U6317 (N_6317,N_4298,N_4000);
nor U6318 (N_6318,N_5796,N_5950);
nand U6319 (N_6319,N_4172,N_4805);
nand U6320 (N_6320,N_4539,N_5117);
and U6321 (N_6321,N_4845,N_4786);
or U6322 (N_6322,N_5802,N_4299);
or U6323 (N_6323,N_5066,N_5035);
or U6324 (N_6324,N_5952,N_5649);
nand U6325 (N_6325,N_5307,N_4944);
nor U6326 (N_6326,N_4863,N_4483);
or U6327 (N_6327,N_5674,N_5249);
xnor U6328 (N_6328,N_4681,N_4976);
xnor U6329 (N_6329,N_4521,N_4700);
nand U6330 (N_6330,N_4564,N_5560);
nand U6331 (N_6331,N_4571,N_4302);
or U6332 (N_6332,N_5456,N_4085);
nand U6333 (N_6333,N_4510,N_4988);
and U6334 (N_6334,N_5749,N_5123);
and U6335 (N_6335,N_4937,N_5895);
or U6336 (N_6336,N_5932,N_4329);
and U6337 (N_6337,N_5034,N_4914);
and U6338 (N_6338,N_5017,N_5349);
and U6339 (N_6339,N_4156,N_5901);
nand U6340 (N_6340,N_4661,N_4455);
or U6341 (N_6341,N_5621,N_4506);
or U6342 (N_6342,N_5172,N_4600);
nand U6343 (N_6343,N_4451,N_4300);
nand U6344 (N_6344,N_4715,N_4742);
and U6345 (N_6345,N_4324,N_4285);
nor U6346 (N_6346,N_5263,N_5114);
or U6347 (N_6347,N_5181,N_4868);
and U6348 (N_6348,N_4215,N_5320);
and U6349 (N_6349,N_4679,N_5175);
nor U6350 (N_6350,N_4325,N_5580);
nor U6351 (N_6351,N_4650,N_5417);
nand U6352 (N_6352,N_4237,N_5885);
nor U6353 (N_6353,N_5162,N_4001);
xnor U6354 (N_6354,N_4754,N_5291);
or U6355 (N_6355,N_5110,N_5391);
xor U6356 (N_6356,N_5710,N_4130);
nor U6357 (N_6357,N_4760,N_5974);
nand U6358 (N_6358,N_4659,N_5760);
nand U6359 (N_6359,N_5819,N_5779);
or U6360 (N_6360,N_5893,N_4671);
nor U6361 (N_6361,N_5544,N_4773);
nor U6362 (N_6362,N_4087,N_4171);
nand U6363 (N_6363,N_5577,N_5419);
nor U6364 (N_6364,N_5113,N_5464);
nor U6365 (N_6365,N_4046,N_4520);
and U6366 (N_6366,N_4203,N_5362);
nor U6367 (N_6367,N_4644,N_5702);
or U6368 (N_6368,N_4162,N_4222);
nand U6369 (N_6369,N_5549,N_4881);
nor U6370 (N_6370,N_4264,N_5586);
and U6371 (N_6371,N_4165,N_5896);
or U6372 (N_6372,N_4387,N_5319);
and U6373 (N_6373,N_5739,N_4090);
and U6374 (N_6374,N_4744,N_5206);
nand U6375 (N_6375,N_5875,N_4258);
nand U6376 (N_6376,N_5124,N_4903);
or U6377 (N_6377,N_4480,N_5261);
or U6378 (N_6378,N_4950,N_4123);
or U6379 (N_6379,N_4311,N_5290);
or U6380 (N_6380,N_4705,N_4017);
nor U6381 (N_6381,N_5720,N_4665);
or U6382 (N_6382,N_4860,N_4953);
nor U6383 (N_6383,N_5981,N_4577);
and U6384 (N_6384,N_5122,N_5244);
or U6385 (N_6385,N_4374,N_4250);
and U6386 (N_6386,N_4048,N_5386);
or U6387 (N_6387,N_5000,N_4332);
nor U6388 (N_6388,N_5125,N_5953);
and U6389 (N_6389,N_4141,N_4676);
and U6390 (N_6390,N_5022,N_5697);
and U6391 (N_6391,N_5083,N_5152);
and U6392 (N_6392,N_4116,N_5698);
nor U6393 (N_6393,N_5474,N_5596);
nand U6394 (N_6394,N_5460,N_5872);
nand U6395 (N_6395,N_5972,N_4169);
or U6396 (N_6396,N_5675,N_5835);
nand U6397 (N_6397,N_4326,N_4794);
nand U6398 (N_6398,N_5518,N_4249);
or U6399 (N_6399,N_5309,N_5229);
nor U6400 (N_6400,N_4204,N_5891);
nor U6401 (N_6401,N_4769,N_4808);
and U6402 (N_6402,N_5182,N_4611);
nand U6403 (N_6403,N_5352,N_4740);
or U6404 (N_6404,N_4989,N_4960);
or U6405 (N_6405,N_4637,N_4260);
nor U6406 (N_6406,N_5638,N_5137);
nand U6407 (N_6407,N_4921,N_4697);
or U6408 (N_6408,N_5483,N_4286);
and U6409 (N_6409,N_4365,N_5931);
nand U6410 (N_6410,N_5311,N_4319);
and U6411 (N_6411,N_5917,N_4800);
and U6412 (N_6412,N_5341,N_5743);
nand U6413 (N_6413,N_4677,N_5598);
nand U6414 (N_6414,N_5902,N_4108);
nand U6415 (N_6415,N_5413,N_5506);
nor U6416 (N_6416,N_4115,N_4859);
and U6417 (N_6417,N_5039,N_4342);
nand U6418 (N_6418,N_5521,N_5270);
nand U6419 (N_6419,N_4674,N_5241);
and U6420 (N_6420,N_4128,N_4728);
and U6421 (N_6421,N_5601,N_5397);
and U6422 (N_6422,N_4995,N_5473);
and U6423 (N_6423,N_5394,N_4590);
nor U6424 (N_6424,N_4507,N_4405);
or U6425 (N_6425,N_5555,N_4358);
nor U6426 (N_6426,N_5525,N_5511);
nor U6427 (N_6427,N_5193,N_5884);
and U6428 (N_6428,N_5287,N_5218);
nor U6429 (N_6429,N_5232,N_5850);
or U6430 (N_6430,N_5758,N_4255);
xor U6431 (N_6431,N_5584,N_4792);
nor U6432 (N_6432,N_5553,N_4759);
nand U6433 (N_6433,N_4446,N_4184);
nor U6434 (N_6434,N_5421,N_5390);
or U6435 (N_6435,N_4848,N_4615);
nand U6436 (N_6436,N_4297,N_4933);
and U6437 (N_6437,N_4762,N_5450);
or U6438 (N_6438,N_5199,N_5250);
nand U6439 (N_6439,N_5626,N_5046);
and U6440 (N_6440,N_5963,N_4846);
or U6441 (N_6441,N_4873,N_4932);
and U6442 (N_6442,N_5795,N_4748);
and U6443 (N_6443,N_5147,N_4416);
and U6444 (N_6444,N_5587,N_4470);
and U6445 (N_6445,N_4481,N_5946);
or U6446 (N_6446,N_5620,N_5195);
nand U6447 (N_6447,N_4541,N_5892);
nor U6448 (N_6448,N_4498,N_5915);
and U6449 (N_6449,N_5699,N_4047);
or U6450 (N_6450,N_4511,N_5191);
or U6451 (N_6451,N_4467,N_5678);
and U6452 (N_6452,N_4148,N_4888);
or U6453 (N_6453,N_5998,N_5765);
or U6454 (N_6454,N_4102,N_4411);
or U6455 (N_6455,N_4684,N_4112);
nand U6456 (N_6456,N_4598,N_5472);
xnor U6457 (N_6457,N_5593,N_4663);
or U6458 (N_6458,N_5693,N_4439);
nand U6459 (N_6459,N_5134,N_5927);
nor U6460 (N_6460,N_5643,N_5538);
or U6461 (N_6461,N_4908,N_5849);
and U6462 (N_6462,N_5433,N_4296);
and U6463 (N_6463,N_5273,N_4948);
or U6464 (N_6464,N_4701,N_5371);
and U6465 (N_6465,N_4832,N_4660);
and U6466 (N_6466,N_4042,N_5995);
nand U6467 (N_6467,N_5139,N_5971);
or U6468 (N_6468,N_4061,N_4126);
nor U6469 (N_6469,N_5026,N_4064);
nor U6470 (N_6470,N_4114,N_5337);
and U6471 (N_6471,N_4186,N_5357);
or U6472 (N_6472,N_4197,N_5869);
or U6473 (N_6473,N_5067,N_5111);
nor U6474 (N_6474,N_4853,N_5434);
nor U6475 (N_6475,N_5298,N_4573);
and U6476 (N_6476,N_4040,N_5911);
nand U6477 (N_6477,N_4857,N_5033);
and U6478 (N_6478,N_4060,N_5165);
or U6479 (N_6479,N_4071,N_4572);
nand U6480 (N_6480,N_4518,N_4261);
and U6481 (N_6481,N_4187,N_5376);
and U6482 (N_6482,N_5913,N_5395);
and U6483 (N_6483,N_5021,N_5715);
or U6484 (N_6484,N_5428,N_4069);
and U6485 (N_6485,N_5700,N_4596);
or U6486 (N_6486,N_4363,N_5133);
nor U6487 (N_6487,N_4431,N_4897);
nand U6488 (N_6488,N_5463,N_4484);
nor U6489 (N_6489,N_5238,N_4709);
nor U6490 (N_6490,N_4078,N_4206);
nor U6491 (N_6491,N_5120,N_4355);
nor U6492 (N_6492,N_4143,N_4228);
and U6493 (N_6493,N_4578,N_4837);
and U6494 (N_6494,N_4010,N_5668);
and U6495 (N_6495,N_4613,N_5616);
and U6496 (N_6496,N_5980,N_5517);
and U6497 (N_6497,N_4639,N_5556);
nand U6498 (N_6498,N_5329,N_4900);
nor U6499 (N_6499,N_4997,N_4576);
and U6500 (N_6500,N_5336,N_4777);
nor U6501 (N_6501,N_4381,N_5381);
and U6502 (N_6502,N_5810,N_4719);
nand U6503 (N_6503,N_5834,N_4788);
nand U6504 (N_6504,N_4396,N_4764);
or U6505 (N_6505,N_4694,N_4711);
nor U6506 (N_6506,N_5202,N_5360);
or U6507 (N_6507,N_5059,N_5185);
nor U6508 (N_6508,N_5732,N_5161);
nand U6509 (N_6509,N_4393,N_4702);
nor U6510 (N_6510,N_5764,N_5073);
nor U6511 (N_6511,N_5933,N_5297);
or U6512 (N_6512,N_4911,N_4774);
nand U6513 (N_6513,N_4723,N_4667);
nand U6514 (N_6514,N_5728,N_4537);
nand U6515 (N_6515,N_4376,N_4275);
or U6516 (N_6516,N_4689,N_4806);
or U6517 (N_6517,N_5007,N_4086);
nor U6518 (N_6518,N_4982,N_5373);
and U6519 (N_6519,N_5969,N_4733);
nand U6520 (N_6520,N_4179,N_4720);
and U6521 (N_6521,N_4154,N_5568);
and U6522 (N_6522,N_4372,N_5031);
nor U6523 (N_6523,N_4812,N_5671);
nor U6524 (N_6524,N_4122,N_5920);
nand U6525 (N_6525,N_4083,N_5064);
nor U6526 (N_6526,N_4328,N_4025);
or U6527 (N_6527,N_5653,N_5959);
nor U6528 (N_6528,N_4525,N_5679);
nand U6529 (N_6529,N_4443,N_5324);
nand U6530 (N_6530,N_4418,N_4438);
and U6531 (N_6531,N_4783,N_4051);
nor U6532 (N_6532,N_4582,N_5102);
nand U6533 (N_6533,N_4043,N_4018);
nand U6534 (N_6534,N_4279,N_5151);
or U6535 (N_6535,N_5253,N_5868);
and U6536 (N_6536,N_5503,N_4066);
or U6537 (N_6537,N_4210,N_4929);
nor U6538 (N_6538,N_4872,N_4780);
and U6539 (N_6539,N_5119,N_4219);
and U6540 (N_6540,N_4542,N_5393);
xor U6541 (N_6541,N_5709,N_5784);
nand U6542 (N_6542,N_4741,N_4698);
xnor U6543 (N_6543,N_4382,N_5854);
nor U6544 (N_6544,N_4349,N_4896);
or U6545 (N_6545,N_5776,N_5605);
or U6546 (N_6546,N_5048,N_4195);
nand U6547 (N_6547,N_5677,N_5286);
nor U6548 (N_6548,N_4595,N_5597);
and U6549 (N_6549,N_4548,N_4142);
or U6550 (N_6550,N_5382,N_4496);
nand U6551 (N_6551,N_5314,N_5194);
nand U6552 (N_6552,N_5916,N_5242);
nand U6553 (N_6553,N_5331,N_5887);
and U6554 (N_6554,N_5726,N_4323);
and U6555 (N_6555,N_5630,N_4295);
or U6556 (N_6556,N_4211,N_4757);
nand U6557 (N_6557,N_5476,N_4217);
or U6558 (N_6558,N_5786,N_4791);
nand U6559 (N_6559,N_4540,N_4425);
nand U6560 (N_6560,N_4019,N_4247);
nor U6561 (N_6561,N_5032,N_5722);
or U6562 (N_6562,N_5534,N_5372);
or U6563 (N_6563,N_4233,N_5457);
or U6564 (N_6564,N_5741,N_4973);
or U6565 (N_6565,N_5941,N_4829);
nand U6566 (N_6566,N_5642,N_5442);
xnor U6567 (N_6567,N_4442,N_4412);
nand U6568 (N_6568,N_4717,N_5737);
nor U6569 (N_6569,N_5983,N_4713);
nor U6570 (N_6570,N_5612,N_4749);
and U6571 (N_6571,N_4850,N_5874);
nand U6572 (N_6572,N_4065,N_5239);
or U6573 (N_6573,N_4838,N_4417);
nand U6574 (N_6574,N_4928,N_4593);
and U6575 (N_6575,N_4306,N_4784);
and U6576 (N_6576,N_4340,N_4193);
and U6577 (N_6577,N_5281,N_4862);
nand U6578 (N_6578,N_4020,N_5267);
nand U6579 (N_6579,N_4474,N_5536);
nor U6580 (N_6580,N_4913,N_5670);
nor U6581 (N_6581,N_4007,N_4902);
and U6582 (N_6582,N_5043,N_4395);
or U6583 (N_6583,N_4341,N_5644);
nand U6584 (N_6584,N_4795,N_5935);
nand U6585 (N_6585,N_5570,N_5815);
nand U6586 (N_6586,N_5447,N_5736);
and U6587 (N_6587,N_5340,N_5431);
or U6588 (N_6588,N_5966,N_4936);
nand U6589 (N_6589,N_4570,N_4248);
nand U6590 (N_6590,N_5662,N_5565);
xor U6591 (N_6591,N_5429,N_5011);
or U6592 (N_6592,N_5512,N_4068);
or U6593 (N_6593,N_5492,N_5407);
or U6594 (N_6594,N_4645,N_5609);
nand U6595 (N_6595,N_4360,N_5163);
or U6596 (N_6596,N_5127,N_5742);
nand U6597 (N_6597,N_4609,N_4050);
xnor U6598 (N_6598,N_4722,N_5153);
nand U6599 (N_6599,N_4895,N_5683);
or U6600 (N_6600,N_5063,N_5315);
nand U6601 (N_6601,N_5991,N_5339);
nor U6602 (N_6602,N_4450,N_4710);
nand U6603 (N_6603,N_4978,N_5384);
nor U6604 (N_6604,N_5944,N_4894);
nand U6605 (N_6605,N_5862,N_4691);
nand U6606 (N_6606,N_4844,N_5510);
and U6607 (N_6607,N_5260,N_4002);
nor U6608 (N_6608,N_5058,N_4610);
nor U6609 (N_6609,N_5879,N_5858);
or U6610 (N_6610,N_5859,N_4736);
and U6611 (N_6611,N_5962,N_5333);
and U6612 (N_6612,N_4178,N_4307);
and U6613 (N_6613,N_5344,N_4992);
and U6614 (N_6614,N_4642,N_5890);
xor U6615 (N_6615,N_4843,N_5166);
nor U6616 (N_6616,N_5065,N_5424);
nand U6617 (N_6617,N_5696,N_4167);
nand U6618 (N_6618,N_5579,N_4129);
or U6619 (N_6619,N_5572,N_5029);
or U6620 (N_6620,N_4125,N_5234);
and U6621 (N_6621,N_5543,N_4314);
or U6622 (N_6622,N_4943,N_4466);
or U6623 (N_6623,N_4729,N_4655);
or U6624 (N_6624,N_4770,N_5665);
nand U6625 (N_6625,N_5756,N_4756);
nor U6626 (N_6626,N_4089,N_4949);
nor U6627 (N_6627,N_4212,N_4477);
or U6628 (N_6628,N_5523,N_5426);
nor U6629 (N_6629,N_5326,N_4608);
nand U6630 (N_6630,N_4623,N_5144);
and U6631 (N_6631,N_5082,N_5725);
nor U6632 (N_6632,N_5198,N_5903);
and U6633 (N_6633,N_4561,N_5651);
nand U6634 (N_6634,N_4413,N_5481);
nor U6635 (N_6635,N_5531,N_4269);
or U6636 (N_6636,N_5332,N_5236);
and U6637 (N_6637,N_5999,N_4312);
nand U6638 (N_6638,N_4106,N_5639);
or U6639 (N_6639,N_5441,N_4244);
nand U6640 (N_6640,N_4082,N_4964);
nand U6641 (N_6641,N_5968,N_5686);
or U6642 (N_6642,N_5685,N_4658);
nand U6643 (N_6643,N_5044,N_5856);
nand U6644 (N_6644,N_5173,N_4121);
nand U6645 (N_6645,N_5772,N_5851);
and U6646 (N_6646,N_4202,N_4278);
nand U6647 (N_6647,N_4687,N_5524);
nor U6648 (N_6648,N_5095,N_5826);
nor U6649 (N_6649,N_5225,N_4535);
or U6650 (N_6650,N_5809,N_4996);
nand U6651 (N_6651,N_5388,N_4750);
nand U6652 (N_6652,N_4580,N_5836);
nand U6653 (N_6653,N_4916,N_5655);
nor U6654 (N_6654,N_4636,N_4560);
and U6655 (N_6655,N_5841,N_5881);
nand U6656 (N_6656,N_5131,N_5252);
or U6657 (N_6657,N_5321,N_5898);
or U6658 (N_6658,N_5947,N_5539);
and U6659 (N_6659,N_4394,N_4252);
nand U6660 (N_6660,N_5666,N_4271);
and U6661 (N_6661,N_5223,N_5905);
or U6662 (N_6662,N_4282,N_5274);
or U6663 (N_6663,N_5562,N_4414);
nor U6664 (N_6664,N_5509,N_5086);
and U6665 (N_6665,N_5196,N_4957);
or U6666 (N_6666,N_5328,N_4972);
and U6667 (N_6667,N_4985,N_5558);
nor U6668 (N_6668,N_4495,N_5006);
or U6669 (N_6669,N_4320,N_5192);
and U6670 (N_6670,N_5960,N_5112);
nand U6671 (N_6671,N_5237,N_4675);
or U6672 (N_6672,N_5954,N_5793);
or U6673 (N_6673,N_4782,N_4468);
nand U6674 (N_6674,N_5451,N_5634);
and U6675 (N_6675,N_5001,N_5491);
and U6676 (N_6676,N_4432,N_5622);
nand U6677 (N_6677,N_5694,N_5410);
nand U6678 (N_6678,N_4303,N_5730);
nand U6679 (N_6679,N_5479,N_4350);
nand U6680 (N_6680,N_5945,N_4761);
nand U6681 (N_6681,N_4597,N_5477);
nand U6682 (N_6682,N_5706,N_5455);
and U6683 (N_6683,N_5762,N_5839);
and U6684 (N_6684,N_4067,N_5865);
or U6685 (N_6685,N_4031,N_4968);
nor U6686 (N_6686,N_4591,N_4063);
nand U6687 (N_6687,N_4403,N_5365);
nor U6688 (N_6688,N_4712,N_5146);
nand U6689 (N_6689,N_4493,N_5938);
nand U6690 (N_6690,N_4433,N_4811);
and U6691 (N_6691,N_5783,N_5437);
nand U6692 (N_6692,N_5359,N_4076);
nand U6693 (N_6693,N_4348,N_4406);
nor U6694 (N_6694,N_5867,N_5529);
or U6695 (N_6695,N_4847,N_5459);
or U6696 (N_6696,N_4094,N_4875);
nor U6697 (N_6697,N_5761,N_4864);
nand U6698 (N_6698,N_5497,N_5882);
and U6699 (N_6699,N_4011,N_5310);
and U6700 (N_6700,N_5233,N_5015);
xnor U6701 (N_6701,N_5846,N_4603);
or U6702 (N_6702,N_4196,N_5132);
nand U6703 (N_6703,N_5754,N_4401);
and U6704 (N_6704,N_5288,N_4181);
or U6705 (N_6705,N_5275,N_4485);
and U6706 (N_6706,N_4961,N_4058);
and U6707 (N_6707,N_5940,N_4183);
nor U6708 (N_6708,N_4213,N_4907);
and U6709 (N_6709,N_4703,N_5289);
and U6710 (N_6710,N_4549,N_4735);
nor U6711 (N_6711,N_4221,N_4336);
nor U6712 (N_6712,N_4955,N_5210);
nand U6713 (N_6713,N_5486,N_5676);
and U6714 (N_6714,N_4890,N_4925);
and U6715 (N_6715,N_5264,N_4776);
nand U6716 (N_6716,N_4029,N_5301);
nor U6717 (N_6717,N_5519,N_4268);
or U6718 (N_6718,N_4209,N_5003);
nor U6719 (N_6719,N_5345,N_5040);
nand U6720 (N_6720,N_4566,N_4887);
nand U6721 (N_6721,N_4807,N_5254);
nand U6722 (N_6722,N_4437,N_4254);
or U6723 (N_6723,N_4849,N_4909);
nand U6724 (N_6724,N_5777,N_4160);
or U6725 (N_6725,N_5129,N_5475);
nor U6726 (N_6726,N_4817,N_5502);
nor U6727 (N_6727,N_5013,N_5266);
nor U6728 (N_6728,N_4793,N_4692);
nor U6729 (N_6729,N_4530,N_4190);
nor U6730 (N_6730,N_5316,N_4379);
nor U6731 (N_6731,N_4546,N_4265);
or U6732 (N_6732,N_5047,N_4092);
or U6733 (N_6733,N_4225,N_5323);
or U6734 (N_6734,N_5027,N_4981);
and U6735 (N_6735,N_5296,N_4430);
nand U6736 (N_6736,N_5561,N_4962);
xor U6737 (N_6737,N_5149,N_5118);
or U6738 (N_6738,N_5445,N_4277);
nor U6739 (N_6739,N_5088,N_5056);
or U6740 (N_6740,N_5993,N_4821);
or U6741 (N_6741,N_5748,N_5733);
and U6742 (N_6742,N_4855,N_4400);
nor U6743 (N_6743,N_4153,N_5089);
nand U6744 (N_6744,N_5610,N_5752);
nand U6745 (N_6745,N_4118,N_4075);
nor U6746 (N_6746,N_5012,N_5824);
nor U6747 (N_6747,N_5627,N_4220);
nand U6748 (N_6748,N_5782,N_4502);
nand U6749 (N_6749,N_5871,N_4294);
nand U6750 (N_6750,N_4538,N_5703);
nand U6751 (N_6751,N_4901,N_5625);
nor U6752 (N_6752,N_4490,N_4651);
nor U6753 (N_6753,N_4643,N_5240);
and U6754 (N_6754,N_4012,N_5967);
or U6755 (N_6755,N_5155,N_4390);
xnor U6756 (N_6756,N_4096,N_5363);
or U6757 (N_6757,N_4428,N_5295);
nand U6758 (N_6758,N_4318,N_4727);
nand U6759 (N_6759,N_4426,N_5843);
and U6760 (N_6760,N_5369,N_5583);
nand U6761 (N_6761,N_4707,N_4276);
nor U6762 (N_6762,N_5910,N_4721);
nor U6763 (N_6763,N_5515,N_4501);
nor U6764 (N_6764,N_4562,N_5090);
nor U6765 (N_6765,N_5735,N_4182);
nand U6766 (N_6766,N_5617,N_4321);
and U6767 (N_6767,N_4878,N_4861);
nand U6768 (N_6768,N_5599,N_4856);
nand U6769 (N_6769,N_5449,N_4440);
and U6770 (N_6770,N_4292,N_5400);
or U6771 (N_6771,N_4281,N_5212);
and U6772 (N_6772,N_4301,N_5964);
or U6773 (N_6773,N_4150,N_4766);
nor U6774 (N_6774,N_5404,N_5853);
nor U6775 (N_6775,N_5948,N_4476);
or U6776 (N_6776,N_5729,N_4383);
xnor U6777 (N_6777,N_5738,N_4230);
nand U6778 (N_6778,N_5104,N_5224);
nor U6779 (N_6779,N_4262,N_5302);
nand U6780 (N_6780,N_5008,N_4145);
nor U6781 (N_6781,N_4963,N_4041);
nand U6782 (N_6782,N_5659,N_5085);
nand U6783 (N_6783,N_5652,N_5478);
or U6784 (N_6784,N_4280,N_4168);
nor U6785 (N_6785,N_4810,N_4478);
and U6786 (N_6786,N_5527,N_5052);
or U6787 (N_6787,N_4970,N_4144);
and U6788 (N_6788,N_4283,N_5505);
nor U6789 (N_6789,N_4458,N_4084);
or U6790 (N_6790,N_5271,N_4680);
and U6791 (N_6791,N_5452,N_5183);
or U6792 (N_6792,N_5107,N_5306);
nand U6793 (N_6793,N_4547,N_4820);
or U6794 (N_6794,N_4263,N_5005);
or U6795 (N_6795,N_4755,N_5115);
nor U6796 (N_6796,N_4974,N_5592);
nand U6797 (N_6797,N_5751,N_5177);
nand U6798 (N_6798,N_5482,N_4103);
xnor U6799 (N_6799,N_5150,N_5103);
nand U6800 (N_6800,N_4869,N_4730);
nand U6801 (N_6801,N_5342,N_5864);
or U6802 (N_6802,N_5408,N_5187);
and U6803 (N_6803,N_5106,N_5546);
or U6804 (N_6804,N_4364,N_5645);
or U6805 (N_6805,N_4124,N_5684);
and U6806 (N_6806,N_4402,N_5994);
xor U6807 (N_6807,N_5949,N_5740);
nand U6808 (N_6808,N_5020,N_4959);
nor U6809 (N_6809,N_5215,N_5681);
or U6810 (N_6810,N_4969,N_4080);
or U6811 (N_6811,N_4958,N_4915);
xnor U6812 (N_6812,N_5283,N_4641);
nand U6813 (N_6813,N_4266,N_5789);
or U6814 (N_6814,N_4672,N_5402);
nand U6815 (N_6815,N_4454,N_4877);
nor U6816 (N_6816,N_5822,N_4778);
nor U6817 (N_6817,N_5635,N_5440);
nor U6818 (N_6818,N_5171,N_4421);
or U6819 (N_6819,N_5444,N_4452);
and U6820 (N_6820,N_4906,N_4424);
nand U6821 (N_6821,N_5157,N_5692);
nor U6822 (N_6822,N_5705,N_4079);
or U6823 (N_6823,N_5468,N_5436);
nand U6824 (N_6824,N_5251,N_4238);
nand U6825 (N_6825,N_5002,N_5396);
and U6826 (N_6826,N_4243,N_5924);
or U6827 (N_6827,N_4751,N_4544);
nor U6828 (N_6828,N_5928,N_4840);
nand U6829 (N_6829,N_4146,N_4956);
and U6830 (N_6830,N_4745,N_5912);
nand U6831 (N_6831,N_5204,N_4188);
and U6832 (N_6832,N_5217,N_5660);
and U6833 (N_6833,N_4579,N_4666);
or U6834 (N_6834,N_5724,N_4205);
nor U6835 (N_6835,N_5201,N_5255);
nand U6836 (N_6836,N_5723,N_5817);
nand U6837 (N_6837,N_5353,N_5842);
nand U6838 (N_6838,N_5495,N_4575);
or U6839 (N_6839,N_4816,N_5399);
nor U6840 (N_6840,N_4815,N_4966);
or U6841 (N_6841,N_4999,N_5019);
nand U6842 (N_6842,N_5848,N_5564);
nand U6843 (N_6843,N_4630,N_4327);
or U6844 (N_6844,N_5838,N_5420);
and U6845 (N_6845,N_5831,N_5347);
and U6846 (N_6846,N_5552,N_4823);
nor U6847 (N_6847,N_5894,N_5398);
xor U6848 (N_6848,N_4865,N_4986);
and U6849 (N_6849,N_5208,N_5818);
nor U6850 (N_6850,N_5937,N_5673);
and U6851 (N_6851,N_5507,N_5220);
and U6852 (N_6852,N_4924,N_5514);
or U6853 (N_6853,N_5855,N_4448);
or U6854 (N_6854,N_4654,N_4201);
or U6855 (N_6855,N_5559,N_4879);
nand U6856 (N_6856,N_4670,N_4947);
or U6857 (N_6857,N_4231,N_5222);
nor U6858 (N_6858,N_4353,N_5934);
or U6859 (N_6859,N_5025,N_4509);
xnor U6860 (N_6860,N_4256,N_4356);
and U6861 (N_6861,N_4407,N_5637);
or U6862 (N_6862,N_4994,N_5667);
nor U6863 (N_6863,N_5282,N_5650);
and U6864 (N_6864,N_5258,N_5446);
nor U6865 (N_6865,N_5788,N_5380);
and U6866 (N_6866,N_4045,N_5414);
and U6867 (N_6867,N_4049,N_4514);
and U6868 (N_6868,N_4993,N_5265);
nor U6869 (N_6869,N_5230,N_4565);
xor U6870 (N_6870,N_4664,N_4686);
and U6871 (N_6871,N_4920,N_5957);
and U6872 (N_6872,N_4874,N_5982);
nor U6873 (N_6873,N_5708,N_4251);
and U6874 (N_6874,N_5235,N_4157);
and U6875 (N_6875,N_4173,N_5327);
and U6876 (N_6876,N_5803,N_4531);
or U6877 (N_6877,N_5461,N_5641);
nor U6878 (N_6878,N_5582,N_4678);
and U6879 (N_6879,N_4931,N_4015);
nor U6880 (N_6880,N_5109,N_4813);
nand U6881 (N_6881,N_5799,N_5262);
or U6882 (N_6882,N_5829,N_5277);
nor U6883 (N_6883,N_4267,N_4946);
nand U6884 (N_6884,N_4635,N_4465);
or U6885 (N_6885,N_5285,N_4435);
nor U6886 (N_6886,N_4052,N_5247);
nor U6887 (N_6887,N_4990,N_5852);
nor U6888 (N_6888,N_5024,N_4647);
and U6889 (N_6889,N_4951,N_4345);
and U6890 (N_6890,N_4475,N_4362);
or U6891 (N_6891,N_4313,N_5068);
and U6892 (N_6892,N_4533,N_4870);
nor U6893 (N_6893,N_4866,N_5567);
or U6894 (N_6894,N_4185,N_5490);
and U6895 (N_6895,N_4088,N_5138);
or U6896 (N_6896,N_4070,N_4135);
nand U6897 (N_6897,N_5318,N_4199);
nand U6898 (N_6898,N_4599,N_4942);
or U6899 (N_6899,N_4758,N_4101);
nand U6900 (N_6900,N_5823,N_4858);
nand U6901 (N_6901,N_5016,N_5925);
or U6902 (N_6902,N_5257,N_5576);
nand U6903 (N_6903,N_5656,N_5159);
nor U6904 (N_6904,N_5588,N_4216);
or U6905 (N_6905,N_5636,N_5448);
nand U6906 (N_6906,N_4696,N_4939);
and U6907 (N_6907,N_5245,N_4952);
or U6908 (N_6908,N_5591,N_5462);
or U6909 (N_6909,N_4589,N_4605);
nor U6910 (N_6910,N_4449,N_5718);
or U6911 (N_6911,N_4606,N_4772);
or U6912 (N_6912,N_5243,N_5305);
or U6913 (N_6913,N_4370,N_4398);
nand U6914 (N_6914,N_4517,N_4910);
or U6915 (N_6915,N_5526,N_5778);
nor U6916 (N_6916,N_4633,N_4410);
or U6917 (N_6917,N_4032,N_4765);
or U6918 (N_6918,N_5516,N_4119);
and U6919 (N_6919,N_4366,N_4427);
and U6920 (N_6920,N_5496,N_5906);
nand U6921 (N_6921,N_5121,N_5508);
and U6922 (N_6922,N_4200,N_5248);
nor U6923 (N_6923,N_5936,N_4488);
and U6924 (N_6924,N_5142,N_5209);
nor U6925 (N_6925,N_4434,N_4062);
nand U6926 (N_6926,N_4208,N_4886);
or U6927 (N_6927,N_5093,N_5387);
and U6928 (N_6928,N_5766,N_4824);
nand U6929 (N_6929,N_5798,N_4388);
nand U6930 (N_6930,N_4716,N_4177);
nand U6931 (N_6931,N_4166,N_4833);
xor U6932 (N_6932,N_4499,N_5873);
and U6933 (N_6933,N_4876,N_5989);
and U6934 (N_6934,N_4227,N_4257);
and U6935 (N_6935,N_4384,N_5607);
and U6936 (N_6936,N_4614,N_5825);
or U6937 (N_6937,N_5299,N_4528);
nand U6938 (N_6938,N_4941,N_5975);
or U6939 (N_6939,N_5179,N_5813);
nand U6940 (N_6940,N_5403,N_4152);
and U6941 (N_6941,N_5077,N_4113);
nand U6942 (N_6942,N_5092,N_4095);
xor U6943 (N_6943,N_4284,N_5704);
nor U6944 (N_6944,N_5921,N_5640);
and U6945 (N_6945,N_4337,N_4164);
nor U6946 (N_6946,N_4409,N_5794);
nand U6947 (N_6947,N_4120,N_5632);
and U6948 (N_6948,N_4305,N_5897);
nor U6949 (N_6949,N_4825,N_4174);
and U6950 (N_6950,N_4272,N_4322);
nand U6951 (N_6951,N_5160,N_4404);
nor U6952 (N_6952,N_4367,N_5294);
or U6953 (N_6953,N_5126,N_4077);
or U6954 (N_6954,N_5745,N_5385);
nand U6955 (N_6955,N_4746,N_5942);
and U6956 (N_6956,N_4673,N_4563);
nand U6957 (N_6957,N_5075,N_4567);
nand U6958 (N_6958,N_5168,N_4423);
and U6959 (N_6959,N_4385,N_5411);
nand U6960 (N_6960,N_5054,N_4891);
and U6961 (N_6961,N_4175,N_4685);
or U6962 (N_6962,N_4229,N_5769);
nor U6963 (N_6963,N_5537,N_5053);
and U6964 (N_6964,N_5943,N_4971);
xnor U6965 (N_6965,N_4904,N_5487);
and U6966 (N_6966,N_5547,N_5354);
and U6967 (N_6967,N_5919,N_5317);
nand U6968 (N_6968,N_4601,N_4189);
or U6969 (N_6969,N_5827,N_5499);
or U6970 (N_6970,N_4688,N_5216);
nor U6971 (N_6971,N_4695,N_4240);
or U6972 (N_6972,N_5070,N_4519);
nand U6973 (N_6973,N_5416,N_4241);
nand U6974 (N_6974,N_4333,N_4690);
and U6975 (N_6975,N_4444,N_5470);
and U6976 (N_6976,N_4030,N_4884);
or U6977 (N_6977,N_5624,N_4460);
and U6978 (N_6978,N_5759,N_5405);
and U6979 (N_6979,N_4819,N_4487);
and U6980 (N_6980,N_4885,N_5493);
nor U6981 (N_6981,N_4775,N_5899);
or U6982 (N_6982,N_5661,N_4768);
and U6983 (N_6983,N_4917,N_4822);
nand U6984 (N_6984,N_4369,N_4841);
nor U6985 (N_6985,N_4109,N_5178);
or U6986 (N_6986,N_5221,N_5530);
nand U6987 (N_6987,N_4386,N_4656);
nor U6988 (N_6988,N_4463,N_5439);
and U6989 (N_6989,N_4111,N_4170);
nor U6990 (N_6990,N_4315,N_4304);
or U6991 (N_6991,N_5785,N_4137);
nor U6992 (N_6992,N_4945,N_4138);
nor U6993 (N_6993,N_4023,N_4747);
and U6994 (N_6994,N_4317,N_4224);
nand U6995 (N_6995,N_5606,N_5970);
xor U6996 (N_6996,N_4377,N_5976);
nor U6997 (N_6997,N_5876,N_4581);
nor U6998 (N_6998,N_4536,N_4977);
and U6999 (N_6999,N_4469,N_4505);
or U7000 (N_7000,N_4477,N_5929);
nand U7001 (N_7001,N_5396,N_5814);
nor U7002 (N_7002,N_4465,N_4193);
nand U7003 (N_7003,N_5365,N_5169);
or U7004 (N_7004,N_4647,N_5378);
nand U7005 (N_7005,N_5446,N_4639);
and U7006 (N_7006,N_5460,N_4345);
or U7007 (N_7007,N_4567,N_5420);
nand U7008 (N_7008,N_5572,N_4979);
nand U7009 (N_7009,N_4543,N_4332);
or U7010 (N_7010,N_4974,N_4233);
or U7011 (N_7011,N_4498,N_4055);
or U7012 (N_7012,N_4859,N_4969);
and U7013 (N_7013,N_4357,N_4915);
nand U7014 (N_7014,N_4001,N_5003);
or U7015 (N_7015,N_4308,N_5598);
or U7016 (N_7016,N_5392,N_4256);
and U7017 (N_7017,N_4495,N_4250);
nor U7018 (N_7018,N_4723,N_5087);
xor U7019 (N_7019,N_5591,N_4946);
and U7020 (N_7020,N_5064,N_4262);
nor U7021 (N_7021,N_5292,N_5406);
nand U7022 (N_7022,N_4368,N_5214);
nand U7023 (N_7023,N_5700,N_5410);
or U7024 (N_7024,N_4397,N_4408);
or U7025 (N_7025,N_5696,N_4184);
and U7026 (N_7026,N_4845,N_5344);
nor U7027 (N_7027,N_4295,N_4013);
nor U7028 (N_7028,N_5232,N_4153);
nor U7029 (N_7029,N_5762,N_4333);
and U7030 (N_7030,N_5892,N_5224);
xor U7031 (N_7031,N_4852,N_4091);
or U7032 (N_7032,N_4724,N_4984);
nor U7033 (N_7033,N_4756,N_4791);
nor U7034 (N_7034,N_4347,N_4222);
nand U7035 (N_7035,N_4386,N_4832);
or U7036 (N_7036,N_5129,N_4918);
nor U7037 (N_7037,N_5974,N_5743);
nand U7038 (N_7038,N_5307,N_4082);
and U7039 (N_7039,N_4735,N_4425);
or U7040 (N_7040,N_5496,N_4970);
nor U7041 (N_7041,N_4179,N_4103);
nand U7042 (N_7042,N_4386,N_5483);
nor U7043 (N_7043,N_4117,N_4334);
and U7044 (N_7044,N_4615,N_5548);
nor U7045 (N_7045,N_4380,N_4059);
nand U7046 (N_7046,N_4820,N_5539);
nor U7047 (N_7047,N_5584,N_5979);
nand U7048 (N_7048,N_4973,N_4639);
nor U7049 (N_7049,N_5822,N_4524);
and U7050 (N_7050,N_4803,N_5316);
nand U7051 (N_7051,N_4034,N_4359);
or U7052 (N_7052,N_5789,N_5007);
or U7053 (N_7053,N_5505,N_5329);
or U7054 (N_7054,N_4661,N_4682);
and U7055 (N_7055,N_4930,N_5413);
nor U7056 (N_7056,N_4465,N_4634);
or U7057 (N_7057,N_4303,N_5043);
or U7058 (N_7058,N_4808,N_4039);
or U7059 (N_7059,N_5264,N_4414);
or U7060 (N_7060,N_4839,N_5244);
xor U7061 (N_7061,N_4829,N_4491);
nor U7062 (N_7062,N_5203,N_4186);
or U7063 (N_7063,N_4851,N_4485);
nor U7064 (N_7064,N_5919,N_5272);
nand U7065 (N_7065,N_5151,N_4337);
or U7066 (N_7066,N_5572,N_4067);
or U7067 (N_7067,N_4682,N_4301);
and U7068 (N_7068,N_5819,N_5312);
nand U7069 (N_7069,N_5904,N_5372);
nand U7070 (N_7070,N_4041,N_4254);
or U7071 (N_7071,N_5108,N_4335);
or U7072 (N_7072,N_4099,N_4628);
and U7073 (N_7073,N_5260,N_4309);
or U7074 (N_7074,N_4934,N_4956);
and U7075 (N_7075,N_4072,N_4734);
and U7076 (N_7076,N_4416,N_4114);
and U7077 (N_7077,N_4983,N_5417);
nand U7078 (N_7078,N_4322,N_4499);
and U7079 (N_7079,N_5526,N_5084);
nor U7080 (N_7080,N_4181,N_4405);
nor U7081 (N_7081,N_4567,N_5479);
or U7082 (N_7082,N_4166,N_5867);
and U7083 (N_7083,N_5866,N_5690);
nor U7084 (N_7084,N_5496,N_4934);
or U7085 (N_7085,N_5631,N_5792);
and U7086 (N_7086,N_5745,N_4472);
nor U7087 (N_7087,N_4427,N_5845);
and U7088 (N_7088,N_4139,N_5539);
and U7089 (N_7089,N_4765,N_4784);
and U7090 (N_7090,N_5829,N_4385);
and U7091 (N_7091,N_4232,N_5542);
nand U7092 (N_7092,N_4632,N_4487);
and U7093 (N_7093,N_4145,N_5140);
and U7094 (N_7094,N_5303,N_4501);
or U7095 (N_7095,N_5682,N_5518);
nand U7096 (N_7096,N_4658,N_4787);
nor U7097 (N_7097,N_5031,N_4715);
and U7098 (N_7098,N_4510,N_4664);
nand U7099 (N_7099,N_5574,N_5855);
nor U7100 (N_7100,N_5321,N_4118);
nor U7101 (N_7101,N_4007,N_4743);
and U7102 (N_7102,N_5084,N_4736);
nand U7103 (N_7103,N_5758,N_5297);
or U7104 (N_7104,N_4508,N_4237);
or U7105 (N_7105,N_4405,N_4461);
or U7106 (N_7106,N_4419,N_4954);
or U7107 (N_7107,N_4582,N_4592);
xor U7108 (N_7108,N_4622,N_4671);
and U7109 (N_7109,N_4069,N_5828);
xor U7110 (N_7110,N_4073,N_4854);
or U7111 (N_7111,N_5942,N_4061);
nand U7112 (N_7112,N_5634,N_4825);
or U7113 (N_7113,N_5460,N_4093);
and U7114 (N_7114,N_5574,N_5546);
or U7115 (N_7115,N_5868,N_5495);
nor U7116 (N_7116,N_5217,N_5686);
or U7117 (N_7117,N_5099,N_5348);
nand U7118 (N_7118,N_5123,N_4913);
nor U7119 (N_7119,N_4975,N_4634);
nand U7120 (N_7120,N_4635,N_4195);
or U7121 (N_7121,N_5842,N_4934);
or U7122 (N_7122,N_4659,N_5972);
or U7123 (N_7123,N_4031,N_5023);
nor U7124 (N_7124,N_5830,N_4491);
and U7125 (N_7125,N_4936,N_5124);
nor U7126 (N_7126,N_5551,N_4807);
and U7127 (N_7127,N_5637,N_5040);
and U7128 (N_7128,N_4927,N_4879);
xnor U7129 (N_7129,N_5493,N_5150);
or U7130 (N_7130,N_5479,N_5905);
or U7131 (N_7131,N_4525,N_5822);
nor U7132 (N_7132,N_5724,N_5983);
nand U7133 (N_7133,N_4765,N_4356);
nand U7134 (N_7134,N_4967,N_5194);
or U7135 (N_7135,N_4379,N_4650);
nor U7136 (N_7136,N_4783,N_5036);
nor U7137 (N_7137,N_5388,N_4977);
or U7138 (N_7138,N_4042,N_5815);
or U7139 (N_7139,N_4072,N_4375);
and U7140 (N_7140,N_5396,N_5610);
or U7141 (N_7141,N_5144,N_5363);
xnor U7142 (N_7142,N_5696,N_5529);
and U7143 (N_7143,N_5291,N_5643);
nor U7144 (N_7144,N_4877,N_5220);
nor U7145 (N_7145,N_4362,N_5697);
xor U7146 (N_7146,N_5785,N_5450);
or U7147 (N_7147,N_4664,N_5566);
nor U7148 (N_7148,N_5348,N_5791);
nand U7149 (N_7149,N_5255,N_5831);
and U7150 (N_7150,N_4466,N_5279);
nor U7151 (N_7151,N_5751,N_4035);
nor U7152 (N_7152,N_4554,N_5559);
nor U7153 (N_7153,N_4874,N_4263);
nand U7154 (N_7154,N_4398,N_4695);
nor U7155 (N_7155,N_4133,N_5829);
nor U7156 (N_7156,N_4048,N_5509);
nor U7157 (N_7157,N_5807,N_4230);
nor U7158 (N_7158,N_5071,N_4788);
and U7159 (N_7159,N_4255,N_5949);
nand U7160 (N_7160,N_5287,N_5796);
or U7161 (N_7161,N_4618,N_5672);
nand U7162 (N_7162,N_4910,N_4800);
or U7163 (N_7163,N_4953,N_4868);
nand U7164 (N_7164,N_4627,N_4432);
and U7165 (N_7165,N_5365,N_5355);
and U7166 (N_7166,N_5641,N_4992);
nor U7167 (N_7167,N_4272,N_5504);
or U7168 (N_7168,N_4460,N_4491);
or U7169 (N_7169,N_4856,N_5683);
nand U7170 (N_7170,N_5145,N_5860);
and U7171 (N_7171,N_4198,N_4098);
or U7172 (N_7172,N_4018,N_4160);
nand U7173 (N_7173,N_4572,N_5986);
or U7174 (N_7174,N_5717,N_5637);
or U7175 (N_7175,N_4952,N_4090);
or U7176 (N_7176,N_5204,N_5048);
nand U7177 (N_7177,N_5481,N_5958);
or U7178 (N_7178,N_5530,N_4631);
or U7179 (N_7179,N_5824,N_4083);
or U7180 (N_7180,N_5663,N_4178);
nand U7181 (N_7181,N_4908,N_5834);
nor U7182 (N_7182,N_5424,N_5542);
or U7183 (N_7183,N_4925,N_4122);
nor U7184 (N_7184,N_4763,N_5726);
nand U7185 (N_7185,N_5064,N_4497);
nor U7186 (N_7186,N_4273,N_5624);
and U7187 (N_7187,N_4526,N_5815);
and U7188 (N_7188,N_4073,N_4308);
nor U7189 (N_7189,N_5991,N_5085);
or U7190 (N_7190,N_4811,N_4621);
nor U7191 (N_7191,N_5204,N_5069);
or U7192 (N_7192,N_5878,N_5049);
and U7193 (N_7193,N_5591,N_4075);
nor U7194 (N_7194,N_4415,N_4127);
or U7195 (N_7195,N_5512,N_5007);
xor U7196 (N_7196,N_4510,N_5462);
or U7197 (N_7197,N_5651,N_4213);
and U7198 (N_7198,N_5499,N_4927);
nand U7199 (N_7199,N_5372,N_5352);
or U7200 (N_7200,N_4411,N_5439);
nor U7201 (N_7201,N_4390,N_4598);
nor U7202 (N_7202,N_4402,N_4570);
and U7203 (N_7203,N_4644,N_4075);
nor U7204 (N_7204,N_4712,N_5921);
nor U7205 (N_7205,N_4902,N_5862);
nor U7206 (N_7206,N_5933,N_4475);
nor U7207 (N_7207,N_4070,N_5977);
and U7208 (N_7208,N_5171,N_5837);
or U7209 (N_7209,N_5287,N_4842);
nand U7210 (N_7210,N_4741,N_5460);
nand U7211 (N_7211,N_5394,N_5220);
nor U7212 (N_7212,N_4383,N_5081);
nor U7213 (N_7213,N_5805,N_4897);
or U7214 (N_7214,N_4956,N_4571);
nor U7215 (N_7215,N_4533,N_5729);
and U7216 (N_7216,N_5644,N_4967);
and U7217 (N_7217,N_4916,N_5983);
and U7218 (N_7218,N_5490,N_5225);
and U7219 (N_7219,N_4882,N_4440);
or U7220 (N_7220,N_4400,N_5266);
nand U7221 (N_7221,N_5665,N_4663);
xor U7222 (N_7222,N_5183,N_5951);
nor U7223 (N_7223,N_5290,N_4584);
or U7224 (N_7224,N_5014,N_4337);
and U7225 (N_7225,N_4543,N_4321);
nand U7226 (N_7226,N_4168,N_5516);
nor U7227 (N_7227,N_5383,N_5280);
and U7228 (N_7228,N_4551,N_5637);
and U7229 (N_7229,N_5673,N_4614);
and U7230 (N_7230,N_5352,N_5371);
nor U7231 (N_7231,N_5598,N_4091);
nor U7232 (N_7232,N_5789,N_5198);
nor U7233 (N_7233,N_4982,N_5982);
nor U7234 (N_7234,N_4487,N_5642);
nor U7235 (N_7235,N_4071,N_5668);
or U7236 (N_7236,N_5714,N_4772);
nor U7237 (N_7237,N_5616,N_4048);
or U7238 (N_7238,N_4096,N_4369);
nor U7239 (N_7239,N_4617,N_4874);
or U7240 (N_7240,N_4597,N_4783);
or U7241 (N_7241,N_4786,N_5736);
nor U7242 (N_7242,N_4283,N_5804);
or U7243 (N_7243,N_5356,N_5582);
nor U7244 (N_7244,N_4322,N_5476);
nor U7245 (N_7245,N_5014,N_4146);
nand U7246 (N_7246,N_5307,N_5005);
nor U7247 (N_7247,N_5020,N_5265);
nor U7248 (N_7248,N_5854,N_4774);
nor U7249 (N_7249,N_5241,N_4793);
nor U7250 (N_7250,N_5378,N_5074);
nand U7251 (N_7251,N_5153,N_4090);
or U7252 (N_7252,N_4340,N_5905);
and U7253 (N_7253,N_5276,N_4941);
nor U7254 (N_7254,N_4326,N_5358);
and U7255 (N_7255,N_4621,N_5544);
and U7256 (N_7256,N_4297,N_4402);
and U7257 (N_7257,N_4915,N_4018);
nor U7258 (N_7258,N_5692,N_5498);
nor U7259 (N_7259,N_4574,N_4025);
nand U7260 (N_7260,N_4031,N_5574);
nand U7261 (N_7261,N_4533,N_4589);
nor U7262 (N_7262,N_5698,N_4489);
and U7263 (N_7263,N_5105,N_5009);
or U7264 (N_7264,N_5656,N_4451);
or U7265 (N_7265,N_4227,N_5539);
or U7266 (N_7266,N_4200,N_5544);
and U7267 (N_7267,N_4124,N_4286);
and U7268 (N_7268,N_5557,N_4051);
or U7269 (N_7269,N_4135,N_5985);
nor U7270 (N_7270,N_4620,N_4604);
xor U7271 (N_7271,N_4994,N_5371);
nor U7272 (N_7272,N_5259,N_4636);
nor U7273 (N_7273,N_5807,N_5998);
or U7274 (N_7274,N_5751,N_5943);
and U7275 (N_7275,N_5881,N_5187);
and U7276 (N_7276,N_5867,N_5036);
and U7277 (N_7277,N_4459,N_5608);
nor U7278 (N_7278,N_4458,N_4863);
and U7279 (N_7279,N_5349,N_5054);
nand U7280 (N_7280,N_4149,N_4320);
nor U7281 (N_7281,N_5490,N_4751);
nand U7282 (N_7282,N_4306,N_4213);
or U7283 (N_7283,N_4198,N_5702);
xnor U7284 (N_7284,N_5922,N_5342);
and U7285 (N_7285,N_4469,N_4269);
and U7286 (N_7286,N_5805,N_5281);
nand U7287 (N_7287,N_4109,N_5451);
xnor U7288 (N_7288,N_5321,N_5906);
or U7289 (N_7289,N_5487,N_4848);
nor U7290 (N_7290,N_5836,N_4999);
or U7291 (N_7291,N_5238,N_4842);
and U7292 (N_7292,N_5127,N_5124);
or U7293 (N_7293,N_4762,N_5439);
and U7294 (N_7294,N_4735,N_5803);
and U7295 (N_7295,N_4555,N_4024);
and U7296 (N_7296,N_5814,N_5195);
and U7297 (N_7297,N_5122,N_4706);
nand U7298 (N_7298,N_5412,N_4445);
or U7299 (N_7299,N_5611,N_5511);
xor U7300 (N_7300,N_4041,N_4709);
nand U7301 (N_7301,N_5891,N_4076);
and U7302 (N_7302,N_4441,N_5401);
and U7303 (N_7303,N_4473,N_4484);
nor U7304 (N_7304,N_4805,N_4845);
and U7305 (N_7305,N_4866,N_4244);
nand U7306 (N_7306,N_4317,N_5708);
or U7307 (N_7307,N_4996,N_5210);
and U7308 (N_7308,N_4753,N_4945);
nor U7309 (N_7309,N_4437,N_4680);
nand U7310 (N_7310,N_5591,N_5920);
or U7311 (N_7311,N_5591,N_5380);
nor U7312 (N_7312,N_4807,N_5439);
or U7313 (N_7313,N_4672,N_4561);
nand U7314 (N_7314,N_4500,N_5071);
nor U7315 (N_7315,N_5073,N_4583);
and U7316 (N_7316,N_5215,N_4473);
and U7317 (N_7317,N_5077,N_5835);
or U7318 (N_7318,N_5119,N_4616);
and U7319 (N_7319,N_5180,N_4249);
nand U7320 (N_7320,N_4101,N_4270);
nor U7321 (N_7321,N_4175,N_5528);
and U7322 (N_7322,N_5438,N_4897);
nand U7323 (N_7323,N_5363,N_5972);
nor U7324 (N_7324,N_4635,N_5722);
nor U7325 (N_7325,N_5878,N_5862);
nor U7326 (N_7326,N_4516,N_4992);
nor U7327 (N_7327,N_5532,N_4301);
or U7328 (N_7328,N_5668,N_4128);
or U7329 (N_7329,N_5503,N_5393);
nor U7330 (N_7330,N_5290,N_4843);
or U7331 (N_7331,N_5024,N_5305);
nor U7332 (N_7332,N_5900,N_5049);
nor U7333 (N_7333,N_4026,N_5794);
nor U7334 (N_7334,N_4598,N_4445);
nand U7335 (N_7335,N_5714,N_4536);
nand U7336 (N_7336,N_4934,N_4170);
nand U7337 (N_7337,N_4487,N_5319);
nand U7338 (N_7338,N_4955,N_5545);
nand U7339 (N_7339,N_4660,N_4469);
or U7340 (N_7340,N_5028,N_5786);
nor U7341 (N_7341,N_4658,N_4031);
and U7342 (N_7342,N_5648,N_5300);
and U7343 (N_7343,N_5955,N_4348);
nor U7344 (N_7344,N_4179,N_4987);
nor U7345 (N_7345,N_5742,N_4105);
or U7346 (N_7346,N_4298,N_4764);
or U7347 (N_7347,N_4483,N_5750);
and U7348 (N_7348,N_5676,N_5119);
nor U7349 (N_7349,N_5378,N_5843);
nor U7350 (N_7350,N_4311,N_5535);
nand U7351 (N_7351,N_4710,N_4852);
or U7352 (N_7352,N_4256,N_5728);
and U7353 (N_7353,N_4208,N_5025);
nand U7354 (N_7354,N_5851,N_5439);
nand U7355 (N_7355,N_5824,N_4574);
and U7356 (N_7356,N_5997,N_5218);
and U7357 (N_7357,N_4690,N_4833);
nor U7358 (N_7358,N_5851,N_5608);
and U7359 (N_7359,N_4549,N_5391);
and U7360 (N_7360,N_5018,N_4589);
and U7361 (N_7361,N_4428,N_5211);
nand U7362 (N_7362,N_5280,N_5361);
or U7363 (N_7363,N_4894,N_5817);
and U7364 (N_7364,N_5149,N_5684);
nor U7365 (N_7365,N_4559,N_5942);
nor U7366 (N_7366,N_4081,N_4555);
nor U7367 (N_7367,N_4416,N_5240);
or U7368 (N_7368,N_4544,N_4004);
or U7369 (N_7369,N_4376,N_5368);
or U7370 (N_7370,N_5434,N_4495);
nor U7371 (N_7371,N_5048,N_5494);
or U7372 (N_7372,N_4650,N_5758);
or U7373 (N_7373,N_4093,N_5464);
nand U7374 (N_7374,N_5117,N_4249);
nor U7375 (N_7375,N_5591,N_4714);
or U7376 (N_7376,N_4738,N_4661);
nand U7377 (N_7377,N_5120,N_4952);
or U7378 (N_7378,N_4666,N_4646);
or U7379 (N_7379,N_4987,N_4762);
nor U7380 (N_7380,N_5156,N_4241);
nor U7381 (N_7381,N_5790,N_4667);
and U7382 (N_7382,N_5062,N_4578);
nor U7383 (N_7383,N_4623,N_4844);
and U7384 (N_7384,N_4494,N_5300);
nor U7385 (N_7385,N_4994,N_5122);
nor U7386 (N_7386,N_5557,N_5608);
or U7387 (N_7387,N_5407,N_5321);
nor U7388 (N_7388,N_5703,N_5896);
nor U7389 (N_7389,N_5342,N_4479);
nor U7390 (N_7390,N_5397,N_5248);
nand U7391 (N_7391,N_4097,N_4250);
nand U7392 (N_7392,N_5710,N_5050);
and U7393 (N_7393,N_5434,N_4941);
nor U7394 (N_7394,N_5466,N_4398);
nand U7395 (N_7395,N_4230,N_5312);
nor U7396 (N_7396,N_4799,N_5868);
nand U7397 (N_7397,N_4774,N_5036);
nor U7398 (N_7398,N_4718,N_4300);
or U7399 (N_7399,N_4772,N_5910);
and U7400 (N_7400,N_5465,N_4378);
nand U7401 (N_7401,N_4121,N_5037);
and U7402 (N_7402,N_4144,N_5671);
nor U7403 (N_7403,N_4445,N_5944);
xnor U7404 (N_7404,N_5787,N_4188);
nor U7405 (N_7405,N_5621,N_4686);
or U7406 (N_7406,N_4885,N_4942);
xor U7407 (N_7407,N_4316,N_5392);
nand U7408 (N_7408,N_5553,N_5171);
nand U7409 (N_7409,N_4412,N_5168);
or U7410 (N_7410,N_4827,N_4814);
nand U7411 (N_7411,N_5975,N_4303);
and U7412 (N_7412,N_4849,N_4065);
nor U7413 (N_7413,N_5719,N_4979);
and U7414 (N_7414,N_4745,N_5045);
and U7415 (N_7415,N_5428,N_5687);
or U7416 (N_7416,N_4057,N_5349);
nand U7417 (N_7417,N_5479,N_5061);
nand U7418 (N_7418,N_5046,N_4031);
and U7419 (N_7419,N_4240,N_5281);
nor U7420 (N_7420,N_4289,N_4272);
nand U7421 (N_7421,N_4588,N_5947);
and U7422 (N_7422,N_4100,N_5918);
nor U7423 (N_7423,N_4707,N_5172);
nor U7424 (N_7424,N_5820,N_5086);
or U7425 (N_7425,N_4190,N_5669);
xnor U7426 (N_7426,N_4806,N_4030);
nor U7427 (N_7427,N_5721,N_5251);
nor U7428 (N_7428,N_4710,N_4577);
or U7429 (N_7429,N_5577,N_4350);
or U7430 (N_7430,N_5229,N_4742);
nand U7431 (N_7431,N_5779,N_5405);
and U7432 (N_7432,N_4527,N_5076);
nand U7433 (N_7433,N_5463,N_4311);
nand U7434 (N_7434,N_5331,N_4105);
or U7435 (N_7435,N_5904,N_5475);
xnor U7436 (N_7436,N_5636,N_4573);
or U7437 (N_7437,N_5472,N_4305);
nand U7438 (N_7438,N_5649,N_4233);
nor U7439 (N_7439,N_4649,N_5941);
and U7440 (N_7440,N_5739,N_4649);
nor U7441 (N_7441,N_5531,N_4073);
and U7442 (N_7442,N_4845,N_4372);
nor U7443 (N_7443,N_5961,N_5081);
or U7444 (N_7444,N_5435,N_5452);
nor U7445 (N_7445,N_4701,N_4371);
nand U7446 (N_7446,N_4018,N_5105);
xor U7447 (N_7447,N_5735,N_5216);
and U7448 (N_7448,N_4435,N_4909);
or U7449 (N_7449,N_4925,N_5899);
nor U7450 (N_7450,N_4639,N_5075);
nand U7451 (N_7451,N_4999,N_5670);
or U7452 (N_7452,N_4334,N_4862);
nor U7453 (N_7453,N_5677,N_4330);
and U7454 (N_7454,N_5394,N_4447);
nand U7455 (N_7455,N_4669,N_5682);
or U7456 (N_7456,N_4096,N_5953);
or U7457 (N_7457,N_4231,N_4687);
nor U7458 (N_7458,N_5574,N_4934);
nand U7459 (N_7459,N_5493,N_5840);
nor U7460 (N_7460,N_5027,N_4393);
nor U7461 (N_7461,N_5109,N_4772);
nor U7462 (N_7462,N_4939,N_4249);
nor U7463 (N_7463,N_5489,N_5826);
and U7464 (N_7464,N_5426,N_4077);
and U7465 (N_7465,N_4386,N_5382);
nor U7466 (N_7466,N_5651,N_4436);
nand U7467 (N_7467,N_5284,N_4147);
and U7468 (N_7468,N_4419,N_5571);
nand U7469 (N_7469,N_4754,N_4067);
or U7470 (N_7470,N_5650,N_4791);
or U7471 (N_7471,N_5929,N_5561);
nor U7472 (N_7472,N_4295,N_4024);
xnor U7473 (N_7473,N_4933,N_5947);
nand U7474 (N_7474,N_5154,N_5453);
nand U7475 (N_7475,N_5501,N_5794);
and U7476 (N_7476,N_5187,N_5804);
nand U7477 (N_7477,N_4599,N_5810);
or U7478 (N_7478,N_4484,N_5596);
or U7479 (N_7479,N_5392,N_4456);
and U7480 (N_7480,N_5410,N_5339);
or U7481 (N_7481,N_5199,N_5348);
and U7482 (N_7482,N_4274,N_5105);
or U7483 (N_7483,N_4166,N_5605);
and U7484 (N_7484,N_4599,N_5578);
nor U7485 (N_7485,N_4944,N_5708);
or U7486 (N_7486,N_5318,N_5210);
or U7487 (N_7487,N_5135,N_4031);
nand U7488 (N_7488,N_5871,N_5590);
nand U7489 (N_7489,N_4002,N_5491);
or U7490 (N_7490,N_5003,N_5326);
or U7491 (N_7491,N_5284,N_5140);
or U7492 (N_7492,N_5280,N_5967);
and U7493 (N_7493,N_4274,N_4987);
nand U7494 (N_7494,N_5027,N_4459);
or U7495 (N_7495,N_5772,N_4696);
or U7496 (N_7496,N_5335,N_4043);
or U7497 (N_7497,N_4080,N_4709);
nand U7498 (N_7498,N_5629,N_4325);
and U7499 (N_7499,N_4691,N_5603);
or U7500 (N_7500,N_4534,N_5564);
nor U7501 (N_7501,N_4801,N_4108);
nand U7502 (N_7502,N_5196,N_5025);
nand U7503 (N_7503,N_5809,N_4268);
nor U7504 (N_7504,N_4882,N_4366);
nand U7505 (N_7505,N_5175,N_4003);
and U7506 (N_7506,N_5116,N_5626);
nor U7507 (N_7507,N_5957,N_5383);
nor U7508 (N_7508,N_5064,N_4797);
nand U7509 (N_7509,N_4311,N_5326);
nor U7510 (N_7510,N_5900,N_5848);
and U7511 (N_7511,N_4833,N_5549);
xnor U7512 (N_7512,N_5213,N_4875);
nand U7513 (N_7513,N_5523,N_4465);
nor U7514 (N_7514,N_4843,N_5816);
and U7515 (N_7515,N_4232,N_5645);
and U7516 (N_7516,N_4339,N_5201);
or U7517 (N_7517,N_4279,N_4516);
and U7518 (N_7518,N_5541,N_5841);
nand U7519 (N_7519,N_5642,N_5699);
nor U7520 (N_7520,N_4562,N_4130);
nand U7521 (N_7521,N_5460,N_5908);
nand U7522 (N_7522,N_4090,N_5654);
or U7523 (N_7523,N_5383,N_5478);
xor U7524 (N_7524,N_4908,N_4292);
nand U7525 (N_7525,N_4234,N_5762);
nor U7526 (N_7526,N_5146,N_5295);
and U7527 (N_7527,N_4971,N_5068);
nor U7528 (N_7528,N_5084,N_5317);
or U7529 (N_7529,N_4959,N_5736);
or U7530 (N_7530,N_4642,N_4223);
or U7531 (N_7531,N_5511,N_4608);
xor U7532 (N_7532,N_4234,N_5100);
nand U7533 (N_7533,N_4296,N_4350);
nor U7534 (N_7534,N_5843,N_5189);
nor U7535 (N_7535,N_4081,N_5250);
nand U7536 (N_7536,N_5445,N_4721);
and U7537 (N_7537,N_4740,N_4372);
or U7538 (N_7538,N_5555,N_5049);
nand U7539 (N_7539,N_4304,N_4383);
or U7540 (N_7540,N_5975,N_5780);
or U7541 (N_7541,N_5168,N_4891);
nor U7542 (N_7542,N_5665,N_5921);
nand U7543 (N_7543,N_5960,N_5096);
and U7544 (N_7544,N_5115,N_5450);
nor U7545 (N_7545,N_4031,N_5157);
or U7546 (N_7546,N_5466,N_5253);
nand U7547 (N_7547,N_4701,N_4282);
and U7548 (N_7548,N_5314,N_5067);
nand U7549 (N_7549,N_5387,N_5242);
or U7550 (N_7550,N_5811,N_4505);
nand U7551 (N_7551,N_4031,N_5494);
nand U7552 (N_7552,N_4030,N_4155);
nand U7553 (N_7553,N_4870,N_4979);
nor U7554 (N_7554,N_5713,N_5340);
nor U7555 (N_7555,N_4085,N_4252);
and U7556 (N_7556,N_5989,N_5193);
and U7557 (N_7557,N_5868,N_4965);
nand U7558 (N_7558,N_4600,N_5424);
xor U7559 (N_7559,N_4385,N_5921);
nand U7560 (N_7560,N_4690,N_5247);
or U7561 (N_7561,N_5238,N_5763);
or U7562 (N_7562,N_5614,N_4984);
and U7563 (N_7563,N_5305,N_4463);
nor U7564 (N_7564,N_5033,N_5321);
or U7565 (N_7565,N_5862,N_5554);
nand U7566 (N_7566,N_4125,N_5606);
or U7567 (N_7567,N_4695,N_5321);
and U7568 (N_7568,N_5043,N_5317);
nand U7569 (N_7569,N_5413,N_5972);
nor U7570 (N_7570,N_4899,N_5300);
nand U7571 (N_7571,N_4417,N_4695);
and U7572 (N_7572,N_4408,N_5760);
or U7573 (N_7573,N_4399,N_5628);
nand U7574 (N_7574,N_5417,N_5409);
nor U7575 (N_7575,N_5475,N_4958);
nor U7576 (N_7576,N_4557,N_5879);
and U7577 (N_7577,N_4983,N_4126);
and U7578 (N_7578,N_5917,N_5043);
nand U7579 (N_7579,N_5461,N_4086);
or U7580 (N_7580,N_4578,N_4305);
nand U7581 (N_7581,N_5493,N_4121);
nand U7582 (N_7582,N_4985,N_4711);
nand U7583 (N_7583,N_4826,N_4449);
and U7584 (N_7584,N_4942,N_5569);
nand U7585 (N_7585,N_4668,N_4667);
xnor U7586 (N_7586,N_5341,N_4006);
and U7587 (N_7587,N_4185,N_4112);
nor U7588 (N_7588,N_4673,N_4335);
nor U7589 (N_7589,N_4417,N_5623);
and U7590 (N_7590,N_4713,N_4139);
or U7591 (N_7591,N_5081,N_4772);
nor U7592 (N_7592,N_4234,N_4564);
nor U7593 (N_7593,N_5104,N_5373);
or U7594 (N_7594,N_5713,N_4888);
nand U7595 (N_7595,N_5453,N_5941);
nor U7596 (N_7596,N_4042,N_4750);
or U7597 (N_7597,N_5568,N_5204);
nor U7598 (N_7598,N_4661,N_5106);
and U7599 (N_7599,N_4612,N_4355);
nor U7600 (N_7600,N_5535,N_5264);
nand U7601 (N_7601,N_5688,N_4218);
nor U7602 (N_7602,N_5523,N_5859);
nor U7603 (N_7603,N_4816,N_5171);
and U7604 (N_7604,N_4070,N_5011);
or U7605 (N_7605,N_5573,N_5319);
nand U7606 (N_7606,N_5532,N_4559);
nand U7607 (N_7607,N_5760,N_4706);
nand U7608 (N_7608,N_5235,N_4117);
or U7609 (N_7609,N_4967,N_5839);
xnor U7610 (N_7610,N_4894,N_5642);
nor U7611 (N_7611,N_5751,N_5552);
nand U7612 (N_7612,N_5765,N_4784);
nand U7613 (N_7613,N_4782,N_5828);
and U7614 (N_7614,N_4214,N_4003);
nand U7615 (N_7615,N_4546,N_5310);
xor U7616 (N_7616,N_5882,N_4872);
nand U7617 (N_7617,N_4124,N_4502);
nor U7618 (N_7618,N_4720,N_5741);
or U7619 (N_7619,N_4915,N_4397);
or U7620 (N_7620,N_4522,N_5693);
nor U7621 (N_7621,N_4073,N_5934);
and U7622 (N_7622,N_5158,N_4023);
nor U7623 (N_7623,N_5010,N_5067);
and U7624 (N_7624,N_4781,N_4598);
nand U7625 (N_7625,N_5815,N_5503);
nand U7626 (N_7626,N_5037,N_5098);
nand U7627 (N_7627,N_5517,N_4625);
and U7628 (N_7628,N_5404,N_4692);
nand U7629 (N_7629,N_5403,N_5742);
and U7630 (N_7630,N_4128,N_5250);
nand U7631 (N_7631,N_4651,N_4672);
nand U7632 (N_7632,N_4139,N_5083);
nor U7633 (N_7633,N_4161,N_4528);
nor U7634 (N_7634,N_4342,N_4188);
or U7635 (N_7635,N_5615,N_4463);
or U7636 (N_7636,N_4605,N_4518);
nand U7637 (N_7637,N_5876,N_4067);
nor U7638 (N_7638,N_4121,N_4161);
nor U7639 (N_7639,N_4230,N_4821);
or U7640 (N_7640,N_4847,N_5493);
and U7641 (N_7641,N_5808,N_4944);
or U7642 (N_7642,N_5545,N_4257);
nor U7643 (N_7643,N_4904,N_5230);
nor U7644 (N_7644,N_4392,N_5116);
and U7645 (N_7645,N_4843,N_5631);
and U7646 (N_7646,N_4548,N_4066);
nor U7647 (N_7647,N_4172,N_5618);
nand U7648 (N_7648,N_4146,N_5961);
and U7649 (N_7649,N_5088,N_4714);
and U7650 (N_7650,N_5601,N_4463);
nand U7651 (N_7651,N_5103,N_5163);
nand U7652 (N_7652,N_5243,N_4868);
or U7653 (N_7653,N_4863,N_4429);
and U7654 (N_7654,N_5419,N_4933);
xnor U7655 (N_7655,N_4621,N_4743);
nor U7656 (N_7656,N_5439,N_5077);
nand U7657 (N_7657,N_4584,N_4277);
or U7658 (N_7658,N_5499,N_5916);
and U7659 (N_7659,N_5041,N_5351);
or U7660 (N_7660,N_4737,N_4760);
and U7661 (N_7661,N_5578,N_4414);
or U7662 (N_7662,N_5896,N_5695);
or U7663 (N_7663,N_4981,N_5290);
and U7664 (N_7664,N_4573,N_4516);
or U7665 (N_7665,N_5642,N_4324);
or U7666 (N_7666,N_5932,N_5336);
and U7667 (N_7667,N_4169,N_5736);
nand U7668 (N_7668,N_5929,N_5896);
and U7669 (N_7669,N_5214,N_4155);
and U7670 (N_7670,N_5373,N_4235);
nand U7671 (N_7671,N_5356,N_5282);
nand U7672 (N_7672,N_4577,N_4386);
nand U7673 (N_7673,N_5888,N_5395);
nand U7674 (N_7674,N_5646,N_4085);
and U7675 (N_7675,N_5522,N_4701);
nor U7676 (N_7676,N_4028,N_5700);
nand U7677 (N_7677,N_4188,N_5717);
nand U7678 (N_7678,N_5590,N_4962);
and U7679 (N_7679,N_5713,N_4307);
nor U7680 (N_7680,N_4838,N_4241);
or U7681 (N_7681,N_5540,N_5416);
nand U7682 (N_7682,N_5501,N_4648);
xnor U7683 (N_7683,N_4170,N_5053);
or U7684 (N_7684,N_5834,N_5932);
nand U7685 (N_7685,N_4742,N_4649);
or U7686 (N_7686,N_5526,N_5872);
nor U7687 (N_7687,N_5378,N_4273);
nand U7688 (N_7688,N_4795,N_4778);
nand U7689 (N_7689,N_4602,N_5565);
and U7690 (N_7690,N_5106,N_4458);
xor U7691 (N_7691,N_4137,N_4428);
and U7692 (N_7692,N_5974,N_5330);
nand U7693 (N_7693,N_5950,N_5708);
or U7694 (N_7694,N_5880,N_4260);
nand U7695 (N_7695,N_5544,N_4714);
nand U7696 (N_7696,N_5705,N_4460);
nand U7697 (N_7697,N_5026,N_4825);
or U7698 (N_7698,N_5419,N_5165);
xnor U7699 (N_7699,N_5014,N_4795);
nand U7700 (N_7700,N_5453,N_5172);
or U7701 (N_7701,N_5762,N_4029);
xor U7702 (N_7702,N_5661,N_4541);
nand U7703 (N_7703,N_4212,N_5202);
nor U7704 (N_7704,N_5517,N_4031);
nand U7705 (N_7705,N_5437,N_5460);
nand U7706 (N_7706,N_5195,N_5762);
nand U7707 (N_7707,N_4589,N_5527);
nor U7708 (N_7708,N_4560,N_4775);
nand U7709 (N_7709,N_4109,N_4918);
and U7710 (N_7710,N_5348,N_4964);
or U7711 (N_7711,N_5640,N_5668);
nor U7712 (N_7712,N_4935,N_4129);
nand U7713 (N_7713,N_5496,N_5034);
and U7714 (N_7714,N_4598,N_4086);
and U7715 (N_7715,N_5759,N_4519);
nor U7716 (N_7716,N_5437,N_5085);
and U7717 (N_7717,N_4717,N_5456);
nand U7718 (N_7718,N_5233,N_5170);
nand U7719 (N_7719,N_5090,N_4839);
nand U7720 (N_7720,N_5570,N_4967);
or U7721 (N_7721,N_5165,N_5959);
or U7722 (N_7722,N_4903,N_5910);
nor U7723 (N_7723,N_5084,N_4137);
nor U7724 (N_7724,N_4824,N_5276);
nor U7725 (N_7725,N_5529,N_5264);
or U7726 (N_7726,N_5026,N_5709);
and U7727 (N_7727,N_4310,N_4406);
and U7728 (N_7728,N_4762,N_4861);
nor U7729 (N_7729,N_5498,N_4771);
nor U7730 (N_7730,N_5547,N_5709);
nor U7731 (N_7731,N_5532,N_4905);
nand U7732 (N_7732,N_5822,N_5566);
nand U7733 (N_7733,N_5200,N_4735);
nor U7734 (N_7734,N_5112,N_4095);
nor U7735 (N_7735,N_4300,N_5248);
nand U7736 (N_7736,N_5553,N_5948);
nor U7737 (N_7737,N_5731,N_5962);
and U7738 (N_7738,N_5629,N_5280);
nor U7739 (N_7739,N_4917,N_4431);
nand U7740 (N_7740,N_4833,N_5979);
and U7741 (N_7741,N_4797,N_5870);
nor U7742 (N_7742,N_5193,N_5941);
nand U7743 (N_7743,N_4346,N_5715);
or U7744 (N_7744,N_4025,N_5550);
and U7745 (N_7745,N_5861,N_4445);
and U7746 (N_7746,N_5723,N_5794);
xor U7747 (N_7747,N_4111,N_4028);
nor U7748 (N_7748,N_5794,N_4728);
and U7749 (N_7749,N_5317,N_4659);
nand U7750 (N_7750,N_4310,N_4364);
or U7751 (N_7751,N_5891,N_4847);
and U7752 (N_7752,N_5784,N_5689);
nand U7753 (N_7753,N_4212,N_5974);
and U7754 (N_7754,N_5273,N_5137);
and U7755 (N_7755,N_4438,N_5326);
or U7756 (N_7756,N_5877,N_4425);
or U7757 (N_7757,N_5718,N_4764);
nand U7758 (N_7758,N_4281,N_4766);
and U7759 (N_7759,N_4897,N_4639);
nand U7760 (N_7760,N_4404,N_5228);
nand U7761 (N_7761,N_5670,N_4116);
and U7762 (N_7762,N_5353,N_4060);
and U7763 (N_7763,N_4703,N_5623);
and U7764 (N_7764,N_4748,N_4500);
and U7765 (N_7765,N_4312,N_5692);
nor U7766 (N_7766,N_4794,N_4988);
and U7767 (N_7767,N_4047,N_4341);
and U7768 (N_7768,N_5380,N_4702);
and U7769 (N_7769,N_5415,N_5237);
or U7770 (N_7770,N_4734,N_5411);
and U7771 (N_7771,N_4686,N_4644);
and U7772 (N_7772,N_5813,N_5123);
or U7773 (N_7773,N_5261,N_5822);
nor U7774 (N_7774,N_4274,N_5351);
and U7775 (N_7775,N_4926,N_5173);
nor U7776 (N_7776,N_4166,N_5187);
and U7777 (N_7777,N_5087,N_5230);
nand U7778 (N_7778,N_4876,N_5117);
or U7779 (N_7779,N_4654,N_5841);
or U7780 (N_7780,N_5109,N_4626);
and U7781 (N_7781,N_4833,N_5889);
nand U7782 (N_7782,N_4094,N_5831);
nand U7783 (N_7783,N_4266,N_4662);
and U7784 (N_7784,N_4731,N_5998);
or U7785 (N_7785,N_4971,N_5205);
nand U7786 (N_7786,N_5031,N_4878);
or U7787 (N_7787,N_4075,N_5086);
nor U7788 (N_7788,N_5158,N_4305);
or U7789 (N_7789,N_4497,N_4291);
and U7790 (N_7790,N_4545,N_5727);
nor U7791 (N_7791,N_4881,N_4108);
and U7792 (N_7792,N_5754,N_4534);
and U7793 (N_7793,N_5386,N_5273);
nand U7794 (N_7794,N_4055,N_5522);
or U7795 (N_7795,N_4557,N_4342);
or U7796 (N_7796,N_4556,N_4571);
nand U7797 (N_7797,N_4105,N_5836);
and U7798 (N_7798,N_4639,N_5003);
or U7799 (N_7799,N_5378,N_5050);
nor U7800 (N_7800,N_4437,N_4317);
nor U7801 (N_7801,N_5088,N_4760);
nand U7802 (N_7802,N_5245,N_4470);
nand U7803 (N_7803,N_5387,N_4053);
xnor U7804 (N_7804,N_5150,N_5571);
nand U7805 (N_7805,N_4944,N_5145);
nor U7806 (N_7806,N_5754,N_5206);
nand U7807 (N_7807,N_4655,N_5473);
nor U7808 (N_7808,N_5306,N_5723);
or U7809 (N_7809,N_4494,N_4400);
nand U7810 (N_7810,N_5534,N_5346);
or U7811 (N_7811,N_4368,N_5792);
or U7812 (N_7812,N_5442,N_5563);
nor U7813 (N_7813,N_4127,N_5547);
xnor U7814 (N_7814,N_5791,N_5117);
or U7815 (N_7815,N_4598,N_4945);
nand U7816 (N_7816,N_4263,N_5624);
or U7817 (N_7817,N_4281,N_4618);
or U7818 (N_7818,N_5627,N_5156);
or U7819 (N_7819,N_4788,N_4087);
or U7820 (N_7820,N_4100,N_4867);
nor U7821 (N_7821,N_5619,N_4755);
nand U7822 (N_7822,N_5442,N_4959);
nand U7823 (N_7823,N_5058,N_5761);
nand U7824 (N_7824,N_5896,N_4058);
nor U7825 (N_7825,N_5557,N_5425);
nand U7826 (N_7826,N_5434,N_4884);
nor U7827 (N_7827,N_4819,N_5310);
or U7828 (N_7828,N_4219,N_4044);
and U7829 (N_7829,N_5185,N_5794);
or U7830 (N_7830,N_5792,N_5029);
nor U7831 (N_7831,N_4942,N_5421);
or U7832 (N_7832,N_5231,N_5012);
xor U7833 (N_7833,N_5829,N_4588);
nor U7834 (N_7834,N_4473,N_5287);
nor U7835 (N_7835,N_5576,N_5942);
or U7836 (N_7836,N_4504,N_4649);
nor U7837 (N_7837,N_5112,N_5039);
nor U7838 (N_7838,N_5336,N_5860);
and U7839 (N_7839,N_4549,N_5059);
or U7840 (N_7840,N_5354,N_4292);
and U7841 (N_7841,N_4315,N_5139);
nor U7842 (N_7842,N_5927,N_5279);
nor U7843 (N_7843,N_4451,N_4622);
or U7844 (N_7844,N_4150,N_5284);
or U7845 (N_7845,N_5334,N_5342);
nor U7846 (N_7846,N_5476,N_5816);
and U7847 (N_7847,N_5277,N_5191);
nor U7848 (N_7848,N_4767,N_5427);
and U7849 (N_7849,N_4183,N_5948);
nor U7850 (N_7850,N_5272,N_4486);
or U7851 (N_7851,N_4508,N_5790);
nand U7852 (N_7852,N_4700,N_4980);
or U7853 (N_7853,N_4042,N_4825);
and U7854 (N_7854,N_5985,N_4003);
and U7855 (N_7855,N_4687,N_4576);
nand U7856 (N_7856,N_4862,N_4450);
or U7857 (N_7857,N_4779,N_4517);
or U7858 (N_7858,N_4334,N_5245);
and U7859 (N_7859,N_4334,N_4679);
or U7860 (N_7860,N_4509,N_5122);
nor U7861 (N_7861,N_5910,N_5630);
or U7862 (N_7862,N_5333,N_4305);
or U7863 (N_7863,N_4211,N_5278);
nor U7864 (N_7864,N_5362,N_5450);
or U7865 (N_7865,N_4394,N_4110);
or U7866 (N_7866,N_4074,N_5655);
xnor U7867 (N_7867,N_4409,N_5499);
nor U7868 (N_7868,N_4270,N_5900);
nor U7869 (N_7869,N_5418,N_4162);
nand U7870 (N_7870,N_5062,N_5668);
nand U7871 (N_7871,N_5026,N_4886);
nand U7872 (N_7872,N_5405,N_4194);
and U7873 (N_7873,N_5385,N_5736);
and U7874 (N_7874,N_4390,N_5558);
or U7875 (N_7875,N_5780,N_4775);
and U7876 (N_7876,N_5814,N_5523);
or U7877 (N_7877,N_5288,N_4617);
nor U7878 (N_7878,N_4261,N_5545);
or U7879 (N_7879,N_5100,N_4785);
or U7880 (N_7880,N_4188,N_5502);
and U7881 (N_7881,N_4840,N_5470);
nor U7882 (N_7882,N_5595,N_5369);
nor U7883 (N_7883,N_5815,N_5719);
and U7884 (N_7884,N_4550,N_4872);
nor U7885 (N_7885,N_5566,N_4394);
and U7886 (N_7886,N_4401,N_5887);
nor U7887 (N_7887,N_5337,N_4502);
and U7888 (N_7888,N_4331,N_4071);
or U7889 (N_7889,N_4129,N_5588);
nor U7890 (N_7890,N_5340,N_4606);
nand U7891 (N_7891,N_5344,N_4411);
and U7892 (N_7892,N_4301,N_5997);
or U7893 (N_7893,N_4586,N_5317);
and U7894 (N_7894,N_4467,N_5632);
nor U7895 (N_7895,N_4877,N_5993);
xor U7896 (N_7896,N_4852,N_5001);
nand U7897 (N_7897,N_4651,N_5075);
nor U7898 (N_7898,N_4890,N_5152);
or U7899 (N_7899,N_5718,N_5271);
or U7900 (N_7900,N_4413,N_4165);
xor U7901 (N_7901,N_4030,N_4477);
nor U7902 (N_7902,N_5245,N_4929);
nor U7903 (N_7903,N_4624,N_4376);
and U7904 (N_7904,N_5818,N_5601);
xor U7905 (N_7905,N_5915,N_5327);
nand U7906 (N_7906,N_4284,N_4544);
nand U7907 (N_7907,N_4760,N_4437);
nor U7908 (N_7908,N_5724,N_4264);
nand U7909 (N_7909,N_5112,N_4679);
or U7910 (N_7910,N_4441,N_5476);
or U7911 (N_7911,N_4023,N_5737);
or U7912 (N_7912,N_5261,N_5208);
nor U7913 (N_7913,N_4779,N_4926);
nor U7914 (N_7914,N_4901,N_4680);
and U7915 (N_7915,N_4291,N_5939);
nor U7916 (N_7916,N_4381,N_4273);
or U7917 (N_7917,N_4927,N_4889);
nand U7918 (N_7918,N_4901,N_4187);
nand U7919 (N_7919,N_5413,N_4964);
nand U7920 (N_7920,N_5178,N_4596);
and U7921 (N_7921,N_4884,N_5633);
nand U7922 (N_7922,N_4135,N_5651);
or U7923 (N_7923,N_4657,N_5009);
nor U7924 (N_7924,N_5880,N_5631);
and U7925 (N_7925,N_5821,N_5017);
xnor U7926 (N_7926,N_4139,N_4060);
nand U7927 (N_7927,N_5284,N_4657);
nand U7928 (N_7928,N_5088,N_4688);
nor U7929 (N_7929,N_4676,N_5285);
and U7930 (N_7930,N_5838,N_5832);
nand U7931 (N_7931,N_4216,N_5060);
nand U7932 (N_7932,N_5685,N_5572);
xor U7933 (N_7933,N_5273,N_5445);
or U7934 (N_7934,N_5805,N_5304);
nand U7935 (N_7935,N_4890,N_4847);
nor U7936 (N_7936,N_4314,N_4605);
nor U7937 (N_7937,N_5799,N_4220);
and U7938 (N_7938,N_4305,N_4563);
nor U7939 (N_7939,N_5921,N_4562);
nor U7940 (N_7940,N_4801,N_4644);
and U7941 (N_7941,N_5041,N_4881);
nor U7942 (N_7942,N_5809,N_5781);
or U7943 (N_7943,N_4562,N_4620);
nand U7944 (N_7944,N_4208,N_4619);
nand U7945 (N_7945,N_5883,N_5867);
and U7946 (N_7946,N_4425,N_5846);
and U7947 (N_7947,N_5347,N_4971);
and U7948 (N_7948,N_5813,N_4296);
nand U7949 (N_7949,N_4310,N_5227);
nand U7950 (N_7950,N_5836,N_5095);
nand U7951 (N_7951,N_5745,N_5310);
or U7952 (N_7952,N_5705,N_4110);
nand U7953 (N_7953,N_4212,N_4219);
and U7954 (N_7954,N_4302,N_5512);
nor U7955 (N_7955,N_4075,N_4895);
nor U7956 (N_7956,N_4830,N_4325);
nor U7957 (N_7957,N_5823,N_5474);
nand U7958 (N_7958,N_5308,N_4797);
nor U7959 (N_7959,N_5833,N_4435);
nand U7960 (N_7960,N_5457,N_4415);
nand U7961 (N_7961,N_4642,N_4730);
nor U7962 (N_7962,N_5607,N_5816);
or U7963 (N_7963,N_5364,N_4227);
nand U7964 (N_7964,N_4900,N_5338);
and U7965 (N_7965,N_4774,N_4080);
nand U7966 (N_7966,N_4326,N_5965);
or U7967 (N_7967,N_4784,N_5746);
or U7968 (N_7968,N_5792,N_5437);
nor U7969 (N_7969,N_4027,N_5726);
nand U7970 (N_7970,N_5786,N_5644);
and U7971 (N_7971,N_5879,N_5567);
nand U7972 (N_7972,N_4474,N_4513);
and U7973 (N_7973,N_5245,N_4261);
or U7974 (N_7974,N_4460,N_4864);
nor U7975 (N_7975,N_4871,N_4831);
or U7976 (N_7976,N_5147,N_4109);
nor U7977 (N_7977,N_4405,N_5994);
nor U7978 (N_7978,N_5510,N_4537);
nand U7979 (N_7979,N_5917,N_4442);
nand U7980 (N_7980,N_5157,N_4091);
nor U7981 (N_7981,N_5693,N_5896);
and U7982 (N_7982,N_5782,N_5310);
nand U7983 (N_7983,N_4206,N_4345);
and U7984 (N_7984,N_5352,N_5460);
nor U7985 (N_7985,N_5044,N_5995);
nor U7986 (N_7986,N_5833,N_4784);
or U7987 (N_7987,N_5399,N_4435);
or U7988 (N_7988,N_4336,N_4500);
or U7989 (N_7989,N_5239,N_5902);
nand U7990 (N_7990,N_4909,N_5678);
or U7991 (N_7991,N_4459,N_4402);
nor U7992 (N_7992,N_4484,N_4800);
and U7993 (N_7993,N_4010,N_5748);
and U7994 (N_7994,N_5188,N_5402);
nand U7995 (N_7995,N_4952,N_4953);
nor U7996 (N_7996,N_4319,N_4366);
nand U7997 (N_7997,N_4932,N_4323);
and U7998 (N_7998,N_4180,N_5145);
nand U7999 (N_7999,N_4469,N_5016);
nor U8000 (N_8000,N_6259,N_6200);
or U8001 (N_8001,N_7567,N_6250);
nand U8002 (N_8002,N_7147,N_6266);
xor U8003 (N_8003,N_6613,N_6540);
and U8004 (N_8004,N_7592,N_6794);
and U8005 (N_8005,N_6461,N_6251);
and U8006 (N_8006,N_6054,N_6309);
nand U8007 (N_8007,N_7859,N_7530);
or U8008 (N_8008,N_7435,N_6811);
and U8009 (N_8009,N_7512,N_6393);
nor U8010 (N_8010,N_7845,N_6357);
and U8011 (N_8011,N_7935,N_6733);
nor U8012 (N_8012,N_6735,N_6053);
and U8013 (N_8013,N_6503,N_6090);
or U8014 (N_8014,N_6809,N_6414);
nor U8015 (N_8015,N_6877,N_6185);
or U8016 (N_8016,N_7714,N_6376);
nand U8017 (N_8017,N_6425,N_7151);
nand U8018 (N_8018,N_7885,N_7405);
nor U8019 (N_8019,N_7084,N_6700);
and U8020 (N_8020,N_6355,N_6391);
and U8021 (N_8021,N_7760,N_6550);
or U8022 (N_8022,N_7924,N_7934);
and U8023 (N_8023,N_6782,N_7825);
nand U8024 (N_8024,N_6037,N_6896);
nand U8025 (N_8025,N_7360,N_7014);
nor U8026 (N_8026,N_6319,N_6203);
nand U8027 (N_8027,N_7977,N_6839);
or U8028 (N_8028,N_6953,N_6799);
or U8029 (N_8029,N_6658,N_6876);
nand U8030 (N_8030,N_7895,N_6863);
or U8031 (N_8031,N_7287,N_6124);
nor U8032 (N_8032,N_7695,N_6846);
nor U8033 (N_8033,N_7400,N_7093);
and U8034 (N_8034,N_7545,N_6862);
nand U8035 (N_8035,N_7890,N_7737);
nand U8036 (N_8036,N_6349,N_7039);
or U8037 (N_8037,N_7773,N_7336);
nor U8038 (N_8038,N_6383,N_7976);
and U8039 (N_8039,N_6107,N_6034);
and U8040 (N_8040,N_6458,N_6462);
nor U8041 (N_8041,N_6298,N_6209);
or U8042 (N_8042,N_6138,N_6365);
nor U8043 (N_8043,N_7484,N_6036);
and U8044 (N_8044,N_7578,N_7502);
and U8045 (N_8045,N_7791,N_7826);
and U8046 (N_8046,N_6316,N_6871);
nor U8047 (N_8047,N_7543,N_6883);
and U8048 (N_8048,N_7096,N_6895);
and U8049 (N_8049,N_7036,N_6438);
nor U8050 (N_8050,N_6274,N_6022);
and U8051 (N_8051,N_7755,N_7271);
nand U8052 (N_8052,N_6720,N_6318);
and U8053 (N_8053,N_7769,N_7029);
nor U8054 (N_8054,N_7541,N_6143);
nand U8055 (N_8055,N_7944,N_7647);
nand U8056 (N_8056,N_6556,N_6601);
nand U8057 (N_8057,N_6120,N_6164);
nand U8058 (N_8058,N_7315,N_6586);
nand U8059 (N_8059,N_7079,N_6031);
nor U8060 (N_8060,N_6715,N_7836);
or U8061 (N_8061,N_6753,N_7062);
or U8062 (N_8062,N_7320,N_6845);
nand U8063 (N_8063,N_6078,N_6016);
or U8064 (N_8064,N_7197,N_6160);
or U8065 (N_8065,N_6714,N_6562);
nand U8066 (N_8066,N_7101,N_6331);
nor U8067 (N_8067,N_6084,N_7408);
or U8068 (N_8068,N_7645,N_6244);
nand U8069 (N_8069,N_6872,N_6171);
nor U8070 (N_8070,N_6935,N_7120);
nor U8071 (N_8071,N_6342,N_7879);
nor U8072 (N_8072,N_7259,N_7945);
or U8073 (N_8073,N_7019,N_6749);
and U8074 (N_8074,N_7429,N_7478);
or U8075 (N_8075,N_7385,N_7839);
and U8076 (N_8076,N_7889,N_6701);
or U8077 (N_8077,N_7196,N_7696);
or U8078 (N_8078,N_7169,N_7787);
or U8079 (N_8079,N_6284,N_7431);
or U8080 (N_8080,N_7805,N_6707);
nor U8081 (N_8081,N_6727,N_7739);
nand U8082 (N_8082,N_7437,N_6282);
and U8083 (N_8083,N_7177,N_7402);
and U8084 (N_8084,N_6335,N_6841);
nor U8085 (N_8085,N_6098,N_7453);
nand U8086 (N_8086,N_7003,N_7579);
or U8087 (N_8087,N_7919,N_7970);
nand U8088 (N_8088,N_6385,N_7966);
and U8089 (N_8089,N_7964,N_6111);
or U8090 (N_8090,N_6497,N_7951);
nor U8091 (N_8091,N_6297,N_6804);
nand U8092 (N_8092,N_6673,N_7247);
nor U8093 (N_8093,N_6265,N_6829);
or U8094 (N_8094,N_7662,N_6437);
or U8095 (N_8095,N_6415,N_6954);
or U8096 (N_8096,N_6228,N_6636);
nand U8097 (N_8097,N_6469,N_6231);
nand U8098 (N_8098,N_7312,N_6330);
nor U8099 (N_8099,N_7493,N_7359);
or U8100 (N_8100,N_7877,N_6956);
nand U8101 (N_8101,N_6010,N_6494);
and U8102 (N_8102,N_6240,N_7228);
and U8103 (N_8103,N_6970,N_7793);
and U8104 (N_8104,N_6370,N_6763);
nor U8105 (N_8105,N_6945,N_7927);
nand U8106 (N_8106,N_6396,N_6739);
nor U8107 (N_8107,N_7290,N_6600);
xnor U8108 (N_8108,N_6071,N_7221);
or U8109 (N_8109,N_7346,N_6802);
nor U8110 (N_8110,N_6592,N_7099);
and U8111 (N_8111,N_6192,N_7911);
nand U8112 (N_8112,N_6619,N_7384);
or U8113 (N_8113,N_6993,N_7412);
and U8114 (N_8114,N_7644,N_7165);
nand U8115 (N_8115,N_7560,N_7089);
or U8116 (N_8116,N_6175,N_6374);
and U8117 (N_8117,N_6201,N_7204);
nand U8118 (N_8118,N_7978,N_7018);
nor U8119 (N_8119,N_6836,N_6598);
nor U8120 (N_8120,N_6405,N_6565);
and U8121 (N_8121,N_6774,N_7713);
or U8122 (N_8122,N_6280,N_6857);
nand U8123 (N_8123,N_6091,N_6410);
nand U8124 (N_8124,N_7032,N_6906);
or U8125 (N_8125,N_6639,N_6198);
and U8126 (N_8126,N_7518,N_6190);
nand U8127 (N_8127,N_6867,N_6239);
nor U8128 (N_8128,N_6610,N_7137);
nor U8129 (N_8129,N_6212,N_7648);
nand U8130 (N_8130,N_6974,N_6074);
nor U8131 (N_8131,N_6798,N_7562);
or U8132 (N_8132,N_7997,N_6483);
nor U8133 (N_8133,N_6449,N_6125);
nor U8134 (N_8134,N_6995,N_7017);
nor U8135 (N_8135,N_7979,N_7707);
and U8136 (N_8136,N_6771,N_7548);
nand U8137 (N_8137,N_6059,N_7738);
nand U8138 (N_8138,N_6402,N_7956);
nor U8139 (N_8139,N_7426,N_6176);
and U8140 (N_8140,N_6165,N_6810);
nor U8141 (N_8141,N_7237,N_6545);
nand U8142 (N_8142,N_7571,N_7637);
nand U8143 (N_8143,N_7386,N_7712);
or U8144 (N_8144,N_7771,N_7328);
and U8145 (N_8145,N_6830,N_7223);
nand U8146 (N_8146,N_6388,N_6267);
xnor U8147 (N_8147,N_7534,N_6672);
and U8148 (N_8148,N_7163,N_7598);
and U8149 (N_8149,N_6434,N_6568);
and U8150 (N_8150,N_6346,N_7702);
and U8151 (N_8151,N_6843,N_7396);
and U8152 (N_8152,N_6641,N_6020);
nor U8153 (N_8153,N_6777,N_7500);
and U8154 (N_8154,N_6805,N_6778);
nor U8155 (N_8155,N_7060,N_7476);
xor U8156 (N_8156,N_7987,N_7333);
and U8157 (N_8157,N_7851,N_6987);
nand U8158 (N_8158,N_6959,N_7296);
and U8159 (N_8159,N_6423,N_6307);
and U8160 (N_8160,N_6129,N_7536);
or U8161 (N_8161,N_7238,N_7471);
nor U8162 (N_8162,N_7378,N_6068);
or U8163 (N_8163,N_6585,N_7905);
or U8164 (N_8164,N_6271,N_6647);
or U8165 (N_8165,N_6910,N_6485);
or U8166 (N_8166,N_6630,N_6989);
nor U8167 (N_8167,N_7557,N_7461);
nor U8168 (N_8168,N_6716,N_7656);
nor U8169 (N_8169,N_6622,N_7337);
and U8170 (N_8170,N_7217,N_6606);
nor U8171 (N_8171,N_6229,N_6013);
and U8172 (N_8172,N_7130,N_7257);
and U8173 (N_8173,N_7861,N_6327);
or U8174 (N_8174,N_7240,N_7600);
and U8175 (N_8175,N_6587,N_6279);
or U8176 (N_8176,N_7837,N_6116);
nand U8177 (N_8177,N_6957,N_6089);
nand U8178 (N_8178,N_7703,N_7954);
and U8179 (N_8179,N_6884,N_6555);
and U8180 (N_8180,N_7466,N_6324);
nand U8181 (N_8181,N_6287,N_6464);
and U8182 (N_8182,N_7377,N_6269);
or U8183 (N_8183,N_6387,N_7743);
nand U8184 (N_8184,N_6696,N_7006);
and U8185 (N_8185,N_6703,N_7225);
or U8186 (N_8186,N_6828,N_7349);
nand U8187 (N_8187,N_7943,N_6960);
nor U8188 (N_8188,N_7065,N_6687);
nor U8189 (N_8189,N_6508,N_7128);
nand U8190 (N_8190,N_7380,N_7303);
nor U8191 (N_8191,N_7416,N_6926);
or U8192 (N_8192,N_6050,N_6303);
nor U8193 (N_8193,N_6534,N_7661);
or U8194 (N_8194,N_7636,N_7201);
and U8195 (N_8195,N_7780,N_6631);
nand U8196 (N_8196,N_6787,N_7794);
nor U8197 (N_8197,N_6167,N_7432);
nand U8198 (N_8198,N_7558,N_6473);
and U8199 (N_8199,N_7799,N_6885);
and U8200 (N_8200,N_6080,N_6024);
and U8201 (N_8201,N_6982,N_6312);
or U8202 (N_8202,N_6332,N_6021);
nor U8203 (N_8203,N_6182,N_7666);
or U8204 (N_8204,N_7125,N_6134);
nand U8205 (N_8205,N_6886,N_7144);
nor U8206 (N_8206,N_6163,N_6547);
and U8207 (N_8207,N_7081,N_6361);
or U8208 (N_8208,N_7403,N_6934);
nor U8209 (N_8209,N_6684,N_7043);
or U8210 (N_8210,N_6242,N_7803);
and U8211 (N_8211,N_6966,N_6903);
nor U8212 (N_8212,N_7941,N_6916);
nand U8213 (N_8213,N_7449,N_7485);
nand U8214 (N_8214,N_7732,N_7507);
and U8215 (N_8215,N_7191,N_7807);
xnor U8216 (N_8216,N_7095,N_6121);
or U8217 (N_8217,N_6853,N_7948);
nand U8218 (N_8218,N_6699,N_6723);
and U8219 (N_8219,N_6975,N_6408);
nand U8220 (N_8220,N_6820,N_7317);
nand U8221 (N_8221,N_6257,N_7835);
nand U8222 (N_8222,N_7782,N_7189);
or U8223 (N_8223,N_7064,N_6215);
nand U8224 (N_8224,N_6310,N_7862);
nor U8225 (N_8225,N_7041,N_7309);
or U8226 (N_8226,N_6133,N_7961);
and U8227 (N_8227,N_7352,N_7857);
and U8228 (N_8228,N_7234,N_7959);
nand U8229 (N_8229,N_7716,N_7646);
nor U8230 (N_8230,N_6911,N_6079);
nor U8231 (N_8231,N_7588,N_6409);
nor U8232 (N_8232,N_7776,N_7602);
and U8233 (N_8233,N_7947,N_7786);
nor U8234 (N_8234,N_7030,N_6301);
and U8235 (N_8235,N_6112,N_7906);
and U8236 (N_8236,N_7143,N_6808);
or U8237 (N_8237,N_7741,N_7054);
and U8238 (N_8238,N_7832,N_7627);
nor U8239 (N_8239,N_6292,N_6999);
or U8240 (N_8240,N_6236,N_7464);
nor U8241 (N_8241,N_7470,N_7730);
xnor U8242 (N_8242,N_7488,N_6130);
nand U8243 (N_8243,N_6218,N_7902);
xor U8244 (N_8244,N_7136,N_6609);
or U8245 (N_8245,N_7338,N_6627);
and U8246 (N_8246,N_6847,N_6375);
nor U8247 (N_8247,N_7838,N_6923);
and U8248 (N_8248,N_7884,N_7563);
nand U8249 (N_8249,N_6145,N_6444);
xnor U8250 (N_8250,N_6214,N_7483);
nand U8251 (N_8251,N_6529,N_6363);
nor U8252 (N_8252,N_7823,N_7972);
or U8253 (N_8253,N_7601,N_7901);
nor U8254 (N_8254,N_7281,N_7181);
or U8255 (N_8255,N_7692,N_7445);
and U8256 (N_8256,N_7671,N_7697);
nor U8257 (N_8257,N_7762,N_7635);
or U8258 (N_8258,N_6360,N_7494);
nand U8259 (N_8259,N_7300,N_7605);
nand U8260 (N_8260,N_7167,N_7407);
nand U8261 (N_8261,N_6936,N_7023);
and U8262 (N_8262,N_7993,N_6043);
nand U8263 (N_8263,N_7842,N_7055);
or U8264 (N_8264,N_6142,N_7314);
nor U8265 (N_8265,N_6887,N_7058);
or U8266 (N_8266,N_7569,N_6477);
or U8267 (N_8267,N_7072,N_6148);
nor U8268 (N_8268,N_6732,N_7157);
nand U8269 (N_8269,N_6191,N_6245);
or U8270 (N_8270,N_7392,N_6261);
or U8271 (N_8271,N_6674,N_6102);
or U8272 (N_8272,N_7001,N_6649);
nand U8273 (N_8273,N_7747,N_6317);
nand U8274 (N_8274,N_7176,N_7731);
and U8275 (N_8275,N_6412,N_6073);
and U8276 (N_8276,N_7971,N_7555);
nor U8277 (N_8277,N_6315,N_7580);
or U8278 (N_8278,N_6168,N_6457);
nand U8279 (N_8279,N_7654,N_6762);
nand U8280 (N_8280,N_7658,N_6334);
nand U8281 (N_8281,N_7524,N_6573);
and U8282 (N_8282,N_6058,N_6984);
and U8283 (N_8283,N_7016,N_7694);
nor U8284 (N_8284,N_7698,N_7491);
and U8285 (N_8285,N_7874,N_7508);
and U8286 (N_8286,N_7946,N_6217);
or U8287 (N_8287,N_7200,N_7620);
and U8288 (N_8288,N_6042,N_7870);
nand U8289 (N_8289,N_7438,N_7634);
or U8290 (N_8290,N_7751,N_7450);
or U8291 (N_8291,N_6669,N_7289);
or U8292 (N_8292,N_7677,N_6117);
nand U8293 (N_8293,N_6602,N_7374);
nor U8294 (N_8294,N_6431,N_6670);
and U8295 (N_8295,N_6407,N_6634);
or U8296 (N_8296,N_7574,N_6660);
nand U8297 (N_8297,N_7275,N_6776);
and U8298 (N_8298,N_6104,N_6256);
nand U8299 (N_8299,N_7267,N_6305);
and U8300 (N_8300,N_6166,N_7659);
or U8301 (N_8301,N_7958,N_7998);
or U8302 (N_8302,N_6759,N_7324);
or U8303 (N_8303,N_7570,N_6411);
or U8304 (N_8304,N_7112,N_7622);
nor U8305 (N_8305,N_6174,N_7778);
nor U8306 (N_8306,N_7241,N_7930);
and U8307 (N_8307,N_6482,N_6768);
nor U8308 (N_8308,N_7080,N_6950);
or U8309 (N_8309,N_7564,N_6183);
and U8310 (N_8310,N_6389,N_6290);
nor U8311 (N_8311,N_7231,N_7710);
and U8312 (N_8312,N_7091,N_7067);
or U8313 (N_8313,N_7085,N_6521);
nand U8314 (N_8314,N_6326,N_7295);
nor U8315 (N_8315,N_6439,N_7355);
and U8316 (N_8316,N_7261,N_7288);
nand U8317 (N_8317,N_6765,N_7783);
or U8318 (N_8318,N_6859,N_6651);
or U8319 (N_8319,N_7367,N_7322);
xor U8320 (N_8320,N_6426,N_7283);
and U8321 (N_8321,N_7307,N_6030);
and U8322 (N_8322,N_7424,N_7316);
nand U8323 (N_8323,N_6403,N_6452);
xnor U8324 (N_8324,N_7373,N_6195);
nand U8325 (N_8325,N_7891,N_6679);
nand U8326 (N_8326,N_6468,N_7013);
nor U8327 (N_8327,N_6527,N_7969);
nand U8328 (N_8328,N_7653,N_7076);
and U8329 (N_8329,N_7918,N_6087);
and U8330 (N_8330,N_7684,N_7596);
or U8331 (N_8331,N_6029,N_6793);
nor U8332 (N_8332,N_6546,N_7599);
and U8333 (N_8333,N_6572,N_7764);
or U8334 (N_8334,N_6996,N_7625);
and U8335 (N_8335,N_6785,N_6943);
nor U8336 (N_8336,N_7606,N_6688);
nor U8337 (N_8337,N_7527,N_7912);
or U8338 (N_8338,N_7452,N_7790);
and U8339 (N_8339,N_7556,N_7904);
and U8340 (N_8340,N_6027,N_7253);
or U8341 (N_8341,N_7418,N_6795);
nor U8342 (N_8342,N_7734,N_6986);
nand U8343 (N_8343,N_6947,N_6907);
or U8344 (N_8344,N_7633,N_7893);
nor U8345 (N_8345,N_6077,N_7528);
nand U8346 (N_8346,N_7473,N_6502);
or U8347 (N_8347,N_6476,N_7156);
nand U8348 (N_8348,N_6211,N_7111);
or U8349 (N_8349,N_7430,N_7990);
and U8350 (N_8350,N_6341,N_6156);
nand U8351 (N_8351,N_6644,N_7973);
nor U8352 (N_8352,N_7066,N_7505);
and U8353 (N_8353,N_7414,N_7342);
nand U8354 (N_8354,N_7004,N_6837);
or U8355 (N_8355,N_7075,N_7434);
and U8356 (N_8356,N_6543,N_6874);
nor U8357 (N_8357,N_6386,N_7999);
or U8358 (N_8358,N_6969,N_6379);
or U8359 (N_8359,N_7428,N_7362);
and U8360 (N_8360,N_7593,N_7985);
and U8361 (N_8361,N_7846,N_7802);
and U8362 (N_8362,N_6158,N_6614);
and U8363 (N_8363,N_7304,N_7767);
and U8364 (N_8364,N_7103,N_7929);
or U8365 (N_8365,N_7607,N_6377);
or U8366 (N_8366,N_6973,N_7327);
nand U8367 (N_8367,N_6942,N_6322);
nor U8368 (N_8368,N_7398,N_7537);
nand U8369 (N_8369,N_6161,N_7753);
and U8370 (N_8370,N_7046,N_7719);
nand U8371 (N_8371,N_6583,N_7375);
nor U8372 (N_8372,N_7497,N_6247);
nand U8373 (N_8373,N_7952,N_7808);
nor U8374 (N_8374,N_7256,N_7159);
and U8375 (N_8375,N_6815,N_7708);
nor U8376 (N_8376,N_6248,N_6559);
and U8377 (N_8377,N_6345,N_6603);
nor U8378 (N_8378,N_7172,N_7132);
xor U8379 (N_8379,N_6803,N_6306);
nor U8380 (N_8380,N_7009,N_6283);
or U8381 (N_8381,N_7082,N_6490);
nor U8382 (N_8382,N_6662,N_7243);
nor U8383 (N_8383,N_6738,N_7109);
nor U8384 (N_8384,N_7989,N_6308);
nand U8385 (N_8385,N_7609,N_6033);
nand U8386 (N_8386,N_7729,N_6786);
and U8387 (N_8387,N_7899,N_7504);
and U8388 (N_8388,N_7192,N_7190);
nand U8389 (N_8389,N_7850,N_6620);
nand U8390 (N_8390,N_6371,N_6766);
xnor U8391 (N_8391,N_6492,N_7628);
or U8392 (N_8392,N_7614,N_6018);
nand U8393 (N_8393,N_7759,N_6612);
or U8394 (N_8394,N_7554,N_6530);
or U8395 (N_8395,N_6390,N_7589);
nor U8396 (N_8396,N_7916,N_7439);
nand U8397 (N_8397,N_7012,N_6047);
nor U8398 (N_8398,N_7404,N_6235);
nand U8399 (N_8399,N_6552,N_7994);
nand U8400 (N_8400,N_6571,N_6009);
or U8401 (N_8401,N_7672,N_7335);
nand U8402 (N_8402,N_7108,N_7361);
or U8403 (N_8403,N_7331,N_6671);
nor U8404 (N_8404,N_7489,N_6510);
nand U8405 (N_8405,N_7178,N_7756);
and U8406 (N_8406,N_6210,N_6584);
and U8407 (N_8407,N_7638,N_7110);
nand U8408 (N_8408,N_7800,N_6232);
or U8409 (N_8409,N_6155,N_6475);
or U8410 (N_8410,N_7549,N_6048);
and U8411 (N_8411,N_7199,N_6243);
nand U8412 (N_8412,N_6575,N_7369);
nand U8413 (N_8413,N_7002,N_7551);
or U8414 (N_8414,N_6618,N_7682);
nor U8415 (N_8415,N_6276,N_7056);
and U8416 (N_8416,N_6536,N_7925);
nand U8417 (N_8417,N_7115,N_6004);
nor U8418 (N_8418,N_7031,N_6237);
nor U8419 (N_8419,N_6702,N_6698);
and U8420 (N_8420,N_7784,N_7297);
nor U8421 (N_8421,N_6840,N_6734);
and U8422 (N_8422,N_6372,N_6500);
or U8423 (N_8423,N_6173,N_6904);
xor U8424 (N_8424,N_6460,N_7198);
xor U8425 (N_8425,N_6105,N_6382);
and U8426 (N_8426,N_6478,N_7991);
and U8427 (N_8427,N_7219,N_7763);
nand U8428 (N_8428,N_7690,N_7853);
and U8429 (N_8429,N_6272,N_7683);
or U8430 (N_8430,N_6420,N_7010);
nor U8431 (N_8431,N_6992,N_6321);
or U8432 (N_8432,N_7873,N_7896);
nand U8433 (N_8433,N_6083,N_7063);
nand U8434 (N_8434,N_7441,N_7260);
or U8435 (N_8435,N_6724,N_6593);
nand U8436 (N_8436,N_6358,N_6806);
nand U8437 (N_8437,N_7718,N_7388);
and U8438 (N_8438,N_7594,N_7323);
nand U8439 (N_8439,N_6435,N_7581);
nand U8440 (N_8440,N_7926,N_7202);
and U8441 (N_8441,N_6685,N_6495);
nand U8442 (N_8442,N_7621,N_6920);
nand U8443 (N_8443,N_7117,N_6854);
nand U8444 (N_8444,N_6114,N_7915);
and U8445 (N_8445,N_6144,N_7344);
and U8446 (N_8446,N_6474,N_6351);
or U8447 (N_8447,N_6325,N_6921);
nand U8448 (N_8448,N_7576,N_6661);
nand U8449 (N_8449,N_7397,N_7291);
nor U8450 (N_8450,N_6560,N_7468);
and U8451 (N_8451,N_7406,N_7611);
nand U8452 (N_8452,N_7768,N_6380);
or U8453 (N_8453,N_6533,N_6711);
xor U8454 (N_8454,N_6226,N_6666);
nor U8455 (N_8455,N_6094,N_6710);
and U8456 (N_8456,N_7141,N_7538);
and U8457 (N_8457,N_6032,N_7106);
xor U8458 (N_8458,N_6101,N_6905);
and U8459 (N_8459,N_7894,N_6648);
and U8460 (N_8460,N_6384,N_6557);
nand U8461 (N_8461,N_7282,N_7427);
nand U8462 (N_8462,N_7306,N_7921);
nor U8463 (N_8463,N_6676,N_7519);
nor U8464 (N_8464,N_7715,N_6339);
and U8465 (N_8465,N_6898,N_7033);
nor U8466 (N_8466,N_7843,N_7211);
nand U8467 (N_8467,N_7852,N_7248);
or U8468 (N_8468,N_7587,N_6399);
nand U8469 (N_8469,N_7436,N_7669);
nor U8470 (N_8470,N_7631,N_7616);
or U8471 (N_8471,N_7539,N_7045);
nor U8472 (N_8472,N_6596,N_7900);
or U8473 (N_8473,N_7351,N_6750);
nor U8474 (N_8474,N_7280,N_6937);
and U8475 (N_8475,N_6890,N_7848);
nor U8476 (N_8476,N_7146,N_7678);
or U8477 (N_8477,N_6693,N_6189);
or U8478 (N_8478,N_6456,N_6624);
or U8479 (N_8479,N_7785,N_6281);
or U8480 (N_8480,N_6925,N_7313);
and U8481 (N_8481,N_7801,N_6747);
nand U8482 (N_8482,N_6962,N_7640);
and U8483 (N_8483,N_7821,N_7910);
xnor U8484 (N_8484,N_7815,N_7048);
and U8485 (N_8485,N_7552,N_6677);
nor U8486 (N_8486,N_6406,N_7829);
or U8487 (N_8487,N_7540,N_6913);
and U8488 (N_8488,N_6930,N_6899);
and U8489 (N_8489,N_7833,N_7639);
xor U8490 (N_8490,N_6875,N_7028);
and U8491 (N_8491,N_7114,N_6621);
nand U8492 (N_8492,N_7415,N_7856);
nand U8493 (N_8493,N_7590,N_6667);
nor U8494 (N_8494,N_7179,N_7481);
nor U8495 (N_8495,N_6635,N_6605);
and U8496 (N_8496,N_7263,N_6052);
nor U8497 (N_8497,N_7255,N_7026);
or U8498 (N_8498,N_7175,N_6574);
nor U8499 (N_8499,N_6721,N_6328);
nor U8500 (N_8500,N_6756,N_6816);
nor U8501 (N_8501,N_6352,N_7188);
or U8502 (N_8502,N_7139,N_7573);
and U8503 (N_8503,N_7419,N_6781);
or U8504 (N_8504,N_6775,N_6958);
and U8505 (N_8505,N_7332,N_6302);
nand U8506 (N_8506,N_7350,N_6499);
nand U8507 (N_8507,N_6553,N_6238);
nor U8508 (N_8508,N_7107,N_7897);
and U8509 (N_8509,N_7040,N_7044);
or U8510 (N_8510,N_7447,N_6817);
nor U8511 (N_8511,N_7725,N_6655);
nand U8512 (N_8512,N_7603,N_7939);
and U8513 (N_8513,N_6866,N_6481);
or U8514 (N_8514,N_6726,N_7207);
nor U8515 (N_8515,N_6169,N_7129);
nor U8516 (N_8516,N_7883,N_6860);
or U8517 (N_8517,N_7986,N_6440);
nand U8518 (N_8518,N_7499,N_7083);
nor U8519 (N_8519,N_7531,N_6580);
xor U8520 (N_8520,N_6162,N_6675);
nor U8521 (N_8521,N_6418,N_7462);
or U8522 (N_8522,N_6177,N_6295);
or U8523 (N_8523,N_6512,N_6814);
or U8524 (N_8524,N_6131,N_6792);
or U8525 (N_8525,N_6686,N_6951);
xor U8526 (N_8526,N_7864,N_6188);
or U8527 (N_8527,N_7868,N_7704);
and U8528 (N_8528,N_6758,N_7871);
or U8529 (N_8529,N_7142,N_7262);
or U8530 (N_8530,N_7727,N_7617);
nor U8531 (N_8531,N_6197,N_6304);
nor U8532 (N_8532,N_6366,N_7166);
nor U8533 (N_8533,N_7148,N_6065);
nor U8534 (N_8534,N_6813,N_7568);
or U8535 (N_8535,N_6746,N_7254);
or U8536 (N_8536,N_6541,N_7706);
and U8537 (N_8537,N_6730,N_7319);
nand U8538 (N_8538,N_6722,N_6848);
nand U8539 (N_8539,N_6472,N_7119);
nor U8540 (N_8540,N_7792,N_7457);
and U8541 (N_8541,N_7409,N_6773);
and U8542 (N_8542,N_7798,N_6196);
nor U8543 (N_8543,N_6858,N_7503);
xor U8544 (N_8544,N_7806,N_6524);
and U8545 (N_8545,N_7865,N_6788);
and U8546 (N_8546,N_7227,N_6977);
or U8547 (N_8547,N_6288,N_6136);
nand U8548 (N_8548,N_6400,N_7443);
nand U8549 (N_8549,N_7847,N_6336);
or U8550 (N_8550,N_7266,N_6908);
nand U8551 (N_8551,N_7047,N_6081);
or U8552 (N_8552,N_6745,N_7668);
or U8553 (N_8553,N_7265,N_7817);
nor U8554 (N_8554,N_7675,N_6404);
nor U8555 (N_8555,N_6865,N_7088);
and U8556 (N_8556,N_7218,N_7220);
and U8557 (N_8557,N_6972,N_6113);
nor U8558 (N_8558,N_7963,N_6216);
and U8559 (N_8559,N_7390,N_7474);
and U8560 (N_8560,N_7226,N_7909);
or U8561 (N_8561,N_7077,N_7250);
or U8562 (N_8562,N_6964,N_7391);
or U8563 (N_8563,N_6743,N_7463);
and U8564 (N_8564,N_6823,N_7748);
and U8565 (N_8565,N_6157,N_6713);
and U8566 (N_8566,N_7914,N_6889);
nand U8567 (N_8567,N_7813,N_7827);
nor U8568 (N_8568,N_6273,N_7618);
nor U8569 (N_8569,N_6147,N_6608);
nand U8570 (N_8570,N_7318,N_6570);
nand U8571 (N_8571,N_6653,N_6914);
nand U8572 (N_8572,N_6589,N_6023);
nand U8573 (N_8573,N_7442,N_6881);
or U8574 (N_8574,N_7357,N_7071);
or U8575 (N_8575,N_6432,N_6225);
nand U8576 (N_8576,N_6507,N_7425);
nand U8577 (N_8577,N_6213,N_6946);
or U8578 (N_8578,N_6539,N_6506);
and U8579 (N_8579,N_7366,N_7740);
nor U8580 (N_8580,N_7506,N_6931);
nor U8581 (N_8581,N_6737,N_6873);
nand U8582 (N_8582,N_6007,N_7863);
or U8583 (N_8583,N_7819,N_7532);
and U8584 (N_8584,N_7816,N_6241);
nand U8585 (N_8585,N_7667,N_6819);
and U8586 (N_8586,N_7135,N_7830);
and U8587 (N_8587,N_6718,N_6451);
or U8588 (N_8588,N_6172,N_7379);
and U8589 (N_8589,N_7610,N_6994);
nand U8590 (N_8590,N_7053,N_6123);
nand U8591 (N_8591,N_7529,N_7348);
nor U8592 (N_8592,N_7809,N_7688);
and U8593 (N_8593,N_6289,N_7957);
or U8594 (N_8594,N_6255,N_6002);
or U8595 (N_8595,N_6712,N_7170);
nor U8596 (N_8596,N_6353,N_6955);
and U8597 (N_8597,N_7649,N_7433);
nor U8598 (N_8598,N_7105,N_7643);
and U8599 (N_8599,N_6929,N_6800);
nor U8600 (N_8600,N_6924,N_6689);
nand U8601 (N_8601,N_6690,N_6126);
nor U8602 (N_8602,N_7232,N_6625);
nand U8603 (N_8603,N_7623,N_6607);
and U8604 (N_8604,N_6291,N_7521);
nor U8605 (N_8605,N_7305,N_6441);
or U8606 (N_8606,N_6135,N_7583);
nand U8607 (N_8607,N_7586,N_6487);
or U8608 (N_8608,N_7233,N_7572);
nand U8609 (N_8609,N_6264,N_7343);
nor U8610 (N_8610,N_6268,N_7490);
nand U8611 (N_8611,N_6918,N_7657);
nor U8612 (N_8612,N_6869,N_6039);
or U8613 (N_8613,N_7389,N_6070);
nor U8614 (N_8614,N_7394,N_6531);
nor U8615 (N_8615,N_7203,N_7122);
and U8616 (N_8616,N_6362,N_7584);
nor U8617 (N_8617,N_6061,N_6367);
nor U8618 (N_8618,N_7995,N_6394);
or U8619 (N_8619,N_6067,N_6719);
nand U8620 (N_8620,N_6465,N_7482);
nor U8621 (N_8621,N_7693,N_6137);
nor U8622 (N_8622,N_7301,N_7411);
and U8623 (N_8623,N_7651,N_7953);
or U8624 (N_8624,N_7050,N_6709);
nor U8625 (N_8625,N_6509,N_6343);
and U8626 (N_8626,N_6897,N_6752);
and U8627 (N_8627,N_6519,N_6678);
nand U8628 (N_8628,N_6528,N_7078);
or U8629 (N_8629,N_6208,N_7855);
nand U8630 (N_8630,N_6554,N_7582);
or U8631 (N_8631,N_6652,N_6150);
or U8632 (N_8632,N_6998,N_6447);
and U8633 (N_8633,N_6159,N_6230);
and U8634 (N_8634,N_7465,N_6180);
nand U8635 (N_8635,N_7709,N_7866);
nand U8636 (N_8636,N_7020,N_7514);
nor U8637 (N_8637,N_7150,N_6170);
or U8638 (N_8638,N_7691,N_7752);
or U8639 (N_8639,N_7721,N_7744);
or U8640 (N_8640,N_7933,N_7024);
or U8641 (N_8641,N_7401,N_6056);
and U8642 (N_8642,N_7113,N_7057);
xor U8643 (N_8643,N_7458,N_6416);
nor U8644 (N_8644,N_7937,N_7981);
or U8645 (N_8645,N_6003,N_6967);
nand U8646 (N_8646,N_7758,N_7229);
nor U8647 (N_8647,N_6430,N_6359);
nand U8648 (N_8648,N_6683,N_6825);
nor U8649 (N_8649,N_7286,N_7073);
and U8650 (N_8650,N_7936,N_6522);
or U8651 (N_8651,N_7585,N_7962);
xor U8652 (N_8652,N_6258,N_6278);
or U8653 (N_8653,N_6373,N_6413);
nor U8654 (N_8654,N_6069,N_6262);
and U8655 (N_8655,N_7070,N_6968);
nand U8656 (N_8656,N_7726,N_6152);
and U8657 (N_8657,N_6944,N_7173);
and U8658 (N_8658,N_6479,N_7974);
and U8659 (N_8659,N_7339,N_6293);
or U8660 (N_8660,N_6491,N_7027);
nor U8661 (N_8661,N_7334,N_7892);
and U8662 (N_8662,N_7277,N_7330);
nor U8663 (N_8663,N_6821,N_6442);
and U8664 (N_8664,N_6347,N_7345);
or U8665 (N_8665,N_6035,N_6204);
nor U8666 (N_8666,N_7460,N_7278);
nor U8667 (N_8667,N_7886,N_7069);
and U8668 (N_8668,N_7797,N_6154);
and U8669 (N_8669,N_6392,N_7216);
xor U8670 (N_8670,N_7968,N_6012);
nor U8671 (N_8671,N_6149,N_7511);
nor U8672 (N_8672,N_6395,N_6832);
nor U8673 (N_8673,N_7038,N_7448);
nand U8674 (N_8674,N_7965,N_6797);
and U8675 (N_8675,N_6471,N_6692);
or U8676 (N_8676,N_7422,N_6695);
and U8677 (N_8677,N_7236,N_6096);
or U8678 (N_8678,N_6852,N_6578);
or U8679 (N_8679,N_7898,N_7194);
or U8680 (N_8680,N_6294,N_6657);
or U8681 (N_8681,N_6764,N_7270);
nor U8682 (N_8682,N_7310,N_6591);
nor U8683 (N_8683,N_6997,N_7230);
nand U8684 (N_8684,N_7681,N_6014);
nand U8685 (N_8685,N_7456,N_7149);
nand U8686 (N_8686,N_7975,N_7268);
nand U8687 (N_8687,N_6221,N_6082);
and U8688 (N_8688,N_6827,N_6549);
and U8689 (N_8689,N_6397,N_7765);
and U8690 (N_8690,N_6501,N_7687);
or U8691 (N_8691,N_6900,N_7276);
nor U8692 (N_8692,N_7356,N_7124);
nor U8693 (N_8693,N_6643,N_6398);
or U8694 (N_8694,N_6901,N_7417);
and U8695 (N_8695,N_6665,N_7880);
nand U8696 (N_8696,N_7860,N_6329);
or U8697 (N_8697,N_6638,N_6663);
or U8698 (N_8698,N_7273,N_7795);
nand U8699 (N_8699,N_6518,N_7381);
and U8700 (N_8700,N_7796,N_6323);
nand U8701 (N_8701,N_7612,N_7547);
nand U8702 (N_8702,N_6939,N_6099);
and U8703 (N_8703,N_6933,N_6354);
nand U8704 (N_8704,N_6526,N_7878);
or U8705 (N_8705,N_7960,N_7996);
nand U8706 (N_8706,N_6949,N_7245);
nor U8707 (N_8707,N_6757,N_6015);
nor U8708 (N_8708,N_7365,N_7517);
nor U8709 (N_8709,N_6260,N_7724);
and U8710 (N_8710,N_7326,N_7098);
xnor U8711 (N_8711,N_7372,N_6005);
nand U8712 (N_8712,N_6588,N_6401);
nor U8713 (N_8713,N_7049,N_7475);
or U8714 (N_8714,N_7311,N_6337);
and U8715 (N_8715,N_7742,N_7745);
or U8716 (N_8716,N_6467,N_7467);
nor U8717 (N_8717,N_7811,N_7523);
nor U8718 (N_8718,N_6378,N_6616);
or U8719 (N_8719,N_6062,N_6705);
nand U8720 (N_8720,N_7224,N_7722);
and U8721 (N_8721,N_6971,N_7949);
nand U8722 (N_8722,N_7059,N_7092);
or U8723 (N_8723,N_7208,N_7535);
nor U8724 (N_8724,N_7510,N_7118);
and U8725 (N_8725,N_6731,N_6028);
nor U8726 (N_8726,N_6963,N_7387);
and U8727 (N_8727,N_7162,N_6041);
nand U8728 (N_8728,N_7206,N_6535);
nor U8729 (N_8729,N_7161,N_6122);
nor U8730 (N_8730,N_7655,N_6141);
xnor U8731 (N_8731,N_7051,N_6205);
nor U8732 (N_8732,N_6489,N_6537);
nor U8733 (N_8733,N_6263,N_7660);
and U8734 (N_8734,N_6311,N_7674);
xor U8735 (N_8735,N_7566,N_7477);
or U8736 (N_8736,N_6523,N_6744);
or U8737 (N_8737,N_7520,N_7154);
or U8738 (N_8738,N_7917,N_6466);
and U8739 (N_8739,N_6019,N_6801);
nor U8740 (N_8740,N_7750,N_7561);
nor U8741 (N_8741,N_7242,N_6045);
and U8742 (N_8742,N_6891,N_6017);
nand U8743 (N_8743,N_6691,N_7185);
and U8744 (N_8744,N_6076,N_6429);
nand U8745 (N_8745,N_6139,N_6085);
nand U8746 (N_8746,N_7486,N_6582);
or U8747 (N_8747,N_6044,N_6300);
nand U8748 (N_8748,N_7244,N_6193);
nor U8749 (N_8749,N_6517,N_7812);
nand U8750 (N_8750,N_7364,N_6564);
nand U8751 (N_8751,N_7025,N_7138);
nand U8752 (N_8752,N_6646,N_6520);
nor U8753 (N_8753,N_6991,N_6092);
or U8754 (N_8754,N_7544,N_7858);
nor U8755 (N_8755,N_6455,N_6850);
nor U8756 (N_8756,N_7775,N_7604);
nand U8757 (N_8757,N_7480,N_7824);
nand U8758 (N_8758,N_6706,N_7302);
and U8759 (N_8759,N_6178,N_7992);
nor U8760 (N_8760,N_7876,N_6493);
or U8761 (N_8761,N_6006,N_7516);
xor U8762 (N_8762,N_6222,N_7164);
nor U8763 (N_8763,N_7353,N_6577);
or U8764 (N_8764,N_6561,N_6941);
nand U8765 (N_8765,N_7498,N_6640);
or U8766 (N_8766,N_7676,N_6842);
xnor U8767 (N_8767,N_6548,N_6818);
and U8768 (N_8768,N_7086,N_6981);
and U8769 (N_8769,N_6807,N_7022);
nor U8770 (N_8770,N_6748,N_6594);
nor U8771 (N_8771,N_6253,N_6008);
nand U8772 (N_8772,N_6484,N_7293);
or U8773 (N_8773,N_7140,N_6772);
nor U8774 (N_8774,N_6207,N_6751);
or U8775 (N_8775,N_6988,N_7299);
or U8776 (N_8776,N_7222,N_7354);
nand U8777 (N_8777,N_7565,N_7341);
nor U8778 (N_8778,N_6454,N_6912);
or U8779 (N_8779,N_6421,N_7061);
nor U8780 (N_8780,N_6513,N_6849);
nor U8781 (N_8781,N_7272,N_6761);
and U8782 (N_8782,N_6604,N_6922);
nand U8783 (N_8783,N_7820,N_6313);
or U8784 (N_8784,N_6151,N_7284);
nor U8785 (N_8785,N_6851,N_6694);
or U8786 (N_8786,N_7575,N_6878);
nor U8787 (N_8787,N_7258,N_6369);
nand U8788 (N_8788,N_6450,N_7686);
or U8789 (N_8789,N_6179,N_6796);
and U8790 (N_8790,N_6350,N_6001);
nand U8791 (N_8791,N_7828,N_6436);
and U8792 (N_8792,N_6254,N_7212);
nand U8793 (N_8793,N_7650,N_6617);
nand U8794 (N_8794,N_6633,N_6340);
and U8795 (N_8795,N_6252,N_7087);
or U8796 (N_8796,N_7754,N_7550);
or U8797 (N_8797,N_6642,N_6046);
nor U8798 (N_8798,N_7308,N_6626);
nand U8799 (N_8799,N_7818,N_7717);
nor U8800 (N_8800,N_7766,N_6224);
or U8801 (N_8801,N_6654,N_7757);
and U8802 (N_8802,N_6049,N_7922);
and U8803 (N_8803,N_6515,N_7679);
or U8804 (N_8804,N_7728,N_6838);
nand U8805 (N_8805,N_6344,N_6127);
or U8806 (N_8806,N_7395,N_7423);
or U8807 (N_8807,N_6980,N_6234);
nand U8808 (N_8808,N_7455,N_7153);
or U8809 (N_8809,N_7102,N_7689);
nor U8810 (N_8810,N_7205,N_7074);
and U8811 (N_8811,N_6000,N_6769);
or U8812 (N_8812,N_7608,N_7983);
and U8813 (N_8813,N_7577,N_6567);
and U8814 (N_8814,N_7235,N_6729);
and U8815 (N_8815,N_7000,N_7881);
or U8816 (N_8816,N_7371,N_7814);
nand U8817 (N_8817,N_6563,N_6368);
nor U8818 (N_8818,N_7182,N_7875);
nand U8819 (N_8819,N_6754,N_7632);
nand U8820 (N_8820,N_6220,N_6880);
or U8821 (N_8821,N_6516,N_6894);
nor U8822 (N_8822,N_6051,N_7701);
nor U8823 (N_8823,N_6109,N_6659);
or U8824 (N_8824,N_7950,N_7869);
and U8825 (N_8825,N_6985,N_6128);
nand U8826 (N_8826,N_7967,N_7615);
nor U8827 (N_8827,N_7630,N_7746);
or U8828 (N_8828,N_6597,N_7376);
nand U8829 (N_8829,N_7187,N_6320);
or U8830 (N_8830,N_7673,N_6202);
nand U8831 (N_8831,N_7908,N_6831);
or U8832 (N_8832,N_6932,N_7214);
or U8833 (N_8833,N_7664,N_6864);
nor U8834 (N_8834,N_7887,N_6917);
nand U8835 (N_8835,N_6026,N_6976);
nand U8836 (N_8836,N_6055,N_7509);
nor U8837 (N_8837,N_6488,N_7822);
nand U8838 (N_8838,N_6011,N_7168);
or U8839 (N_8839,N_7068,N_7440);
and U8840 (N_8840,N_6270,N_6595);
nor U8841 (N_8841,N_6186,N_7269);
and U8842 (N_8842,N_6296,N_6199);
nor U8843 (N_8843,N_7492,N_6038);
xor U8844 (N_8844,N_7595,N_6656);
xnor U8845 (N_8845,N_7444,N_7772);
nor U8846 (N_8846,N_7652,N_7685);
or U8847 (N_8847,N_6856,N_7420);
nand U8848 (N_8848,N_7239,N_6422);
nor U8849 (N_8849,N_7008,N_7501);
and U8850 (N_8850,N_7104,N_7882);
nor U8851 (N_8851,N_6783,N_6095);
and U8852 (N_8852,N_7034,N_6664);
nand U8853 (N_8853,N_7383,N_6835);
or U8854 (N_8854,N_7184,N_7736);
and U8855 (N_8855,N_6443,N_6097);
nand U8856 (N_8856,N_6990,N_6532);
and U8857 (N_8857,N_6060,N_7393);
nor U8858 (N_8858,N_6459,N_6338);
or U8859 (N_8859,N_6504,N_7938);
or U8860 (N_8860,N_7735,N_7264);
nor U8861 (N_8861,N_7274,N_6505);
and U8862 (N_8862,N_6140,N_7294);
and U8863 (N_8863,N_7446,N_7252);
or U8864 (N_8864,N_6888,N_6611);
nor U8865 (N_8865,N_6704,N_7699);
and U8866 (N_8866,N_6146,N_6417);
or U8867 (N_8867,N_6486,N_7624);
or U8868 (N_8868,N_6364,N_7597);
nor U8869 (N_8869,N_6790,N_7940);
nand U8870 (N_8870,N_7546,N_6064);
nor U8871 (N_8871,N_6496,N_7711);
or U8872 (N_8872,N_6348,N_6187);
and U8873 (N_8873,N_7913,N_7663);
or U8874 (N_8874,N_7127,N_6632);
nand U8875 (N_8875,N_7988,N_6952);
or U8876 (N_8876,N_7788,N_7700);
and U8877 (N_8877,N_7923,N_7298);
nand U8878 (N_8878,N_7131,N_6668);
xor U8879 (N_8879,N_7021,N_7155);
or U8880 (N_8880,N_6299,N_7410);
nand U8881 (N_8881,N_6480,N_6767);
or U8882 (N_8882,N_7421,N_7145);
and U8883 (N_8883,N_7629,N_7370);
and U8884 (N_8884,N_7097,N_6181);
nor U8885 (N_8885,N_6736,N_6779);
nand U8886 (N_8886,N_6558,N_6542);
nor U8887 (N_8887,N_6855,N_6286);
nor U8888 (N_8888,N_6833,N_6086);
or U8889 (N_8889,N_7928,N_7591);
nor U8890 (N_8890,N_7641,N_7347);
nand U8891 (N_8891,N_7515,N_7779);
and U8892 (N_8892,N_7761,N_7626);
nand U8893 (N_8893,N_7292,N_6103);
and U8894 (N_8894,N_6433,N_7522);
xnor U8895 (N_8895,N_7613,N_7867);
nand U8896 (N_8896,N_6861,N_7513);
nand U8897 (N_8897,N_7723,N_6184);
and U8898 (N_8898,N_6979,N_6511);
and U8899 (N_8899,N_7872,N_7210);
or U8900 (N_8900,N_6826,N_6093);
nand U8901 (N_8901,N_6615,N_7249);
nand U8902 (N_8902,N_7495,N_7246);
and U8903 (N_8903,N_7559,N_7733);
nor U8904 (N_8904,N_7749,N_7542);
or U8905 (N_8905,N_6879,N_6576);
nor U8906 (N_8906,N_6928,N_6498);
and U8907 (N_8907,N_6742,N_6100);
nor U8908 (N_8908,N_6463,N_7042);
nor U8909 (N_8909,N_7888,N_6961);
or U8910 (N_8910,N_7171,N_6697);
and U8911 (N_8911,N_6381,N_6233);
nor U8912 (N_8912,N_6915,N_7526);
nand U8913 (N_8913,N_7496,N_7100);
and U8914 (N_8914,N_7183,N_6314);
nor U8915 (N_8915,N_6249,N_7358);
or U8916 (N_8916,N_7789,N_7854);
and U8917 (N_8917,N_6728,N_6740);
nand U8918 (N_8918,N_6581,N_7487);
or U8919 (N_8919,N_7705,N_7459);
and U8920 (N_8920,N_6025,N_7804);
and U8921 (N_8921,N_7015,N_7451);
and U8922 (N_8922,N_7094,N_7810);
nand U8923 (N_8923,N_7955,N_7126);
nor U8924 (N_8924,N_6682,N_6118);
nor U8925 (N_8925,N_7469,N_7831);
nand U8926 (N_8926,N_7553,N_7841);
or U8927 (N_8927,N_6599,N_7180);
or U8928 (N_8928,N_6824,N_7665);
and U8929 (N_8929,N_6909,N_6948);
nand U8930 (N_8930,N_7123,N_6356);
nor U8931 (N_8931,N_6978,N_7642);
and U8932 (N_8932,N_6965,N_7777);
or U8933 (N_8933,N_7195,N_6446);
and U8934 (N_8934,N_7399,N_7413);
nor U8935 (N_8935,N_6219,N_6927);
nand U8936 (N_8936,N_6902,N_6708);
or U8937 (N_8937,N_7770,N_7116);
or U8938 (N_8938,N_6275,N_6983);
nand U8939 (N_8939,N_6791,N_6770);
nand U8940 (N_8940,N_6246,N_6066);
or U8941 (N_8941,N_7619,N_7340);
nor U8942 (N_8942,N_7849,N_6453);
or U8943 (N_8943,N_7840,N_6206);
or U8944 (N_8944,N_6681,N_6629);
or U8945 (N_8945,N_6870,N_6822);
or U8946 (N_8946,N_7670,N_6893);
or U8947 (N_8947,N_6569,N_6590);
and U8948 (N_8948,N_7215,N_6834);
nand U8949 (N_8949,N_7454,N_6057);
and U8950 (N_8950,N_6637,N_6623);
and U8951 (N_8951,N_7007,N_7052);
and U8952 (N_8952,N_6544,N_6106);
nand U8953 (N_8953,N_7279,N_6063);
or U8954 (N_8954,N_6780,N_6812);
nand U8955 (N_8955,N_6333,N_7158);
or U8956 (N_8956,N_7931,N_7920);
nor U8957 (N_8957,N_7321,N_7479);
or U8958 (N_8958,N_6227,N_7363);
and U8959 (N_8959,N_6072,N_6110);
nand U8960 (N_8960,N_7980,N_6424);
nor U8961 (N_8961,N_6075,N_7720);
or U8962 (N_8962,N_6844,N_7133);
nor U8963 (N_8963,N_7984,N_7368);
nand U8964 (N_8964,N_6882,N_7193);
nor U8965 (N_8965,N_6115,N_6938);
or U8966 (N_8966,N_6194,N_7152);
or U8967 (N_8967,N_6153,N_7174);
nand U8968 (N_8968,N_6919,N_6566);
nor U8969 (N_8969,N_7942,N_7160);
nor U8970 (N_8970,N_6755,N_6445);
nand U8971 (N_8971,N_6784,N_7533);
nand U8972 (N_8972,N_6650,N_7382);
nand U8973 (N_8973,N_7472,N_7844);
nor U8974 (N_8974,N_6717,N_7932);
or U8975 (N_8975,N_6680,N_6428);
nor U8976 (N_8976,N_6628,N_7209);
xor U8977 (N_8977,N_7186,N_7834);
or U8978 (N_8978,N_6427,N_6132);
nor U8979 (N_8979,N_7121,N_7781);
nor U8980 (N_8980,N_6448,N_6514);
or U8981 (N_8981,N_6551,N_7680);
nand U8982 (N_8982,N_6040,N_6525);
nand U8983 (N_8983,N_6108,N_7774);
or U8984 (N_8984,N_6645,N_7213);
or U8985 (N_8985,N_7903,N_6223);
nor U8986 (N_8986,N_6538,N_6741);
or U8987 (N_8987,N_6760,N_6789);
xnor U8988 (N_8988,N_7325,N_6940);
nand U8989 (N_8989,N_6419,N_7251);
nor U8990 (N_8990,N_7005,N_6892);
or U8991 (N_8991,N_7907,N_7329);
or U8992 (N_8992,N_7982,N_6277);
nor U8993 (N_8993,N_6868,N_6119);
nand U8994 (N_8994,N_7285,N_6088);
nand U8995 (N_8995,N_6470,N_7035);
nor U8996 (N_8996,N_6725,N_7037);
nor U8997 (N_8997,N_7011,N_7525);
and U8998 (N_8998,N_7134,N_6579);
nor U8999 (N_8999,N_6285,N_7090);
xnor U9000 (N_9000,N_7334,N_7512);
nand U9001 (N_9001,N_6754,N_7601);
nand U9002 (N_9002,N_6289,N_6453);
nor U9003 (N_9003,N_7744,N_7600);
or U9004 (N_9004,N_7342,N_7006);
or U9005 (N_9005,N_6620,N_7066);
nand U9006 (N_9006,N_6775,N_7018);
nor U9007 (N_9007,N_7968,N_7053);
nor U9008 (N_9008,N_7590,N_7849);
xor U9009 (N_9009,N_6142,N_7764);
nor U9010 (N_9010,N_7096,N_6304);
or U9011 (N_9011,N_7880,N_7805);
nand U9012 (N_9012,N_6632,N_6792);
nand U9013 (N_9013,N_6944,N_7684);
nand U9014 (N_9014,N_7518,N_7158);
and U9015 (N_9015,N_6362,N_7365);
or U9016 (N_9016,N_7217,N_6502);
and U9017 (N_9017,N_7901,N_7381);
or U9018 (N_9018,N_6651,N_7451);
nor U9019 (N_9019,N_6668,N_6973);
or U9020 (N_9020,N_7934,N_7349);
nor U9021 (N_9021,N_7969,N_6220);
nor U9022 (N_9022,N_6878,N_7860);
nor U9023 (N_9023,N_6028,N_6721);
nand U9024 (N_9024,N_6450,N_7006);
and U9025 (N_9025,N_6354,N_7481);
nand U9026 (N_9026,N_7623,N_7181);
and U9027 (N_9027,N_6992,N_7893);
nor U9028 (N_9028,N_7509,N_6352);
xor U9029 (N_9029,N_6835,N_6566);
xor U9030 (N_9030,N_7409,N_6156);
and U9031 (N_9031,N_7310,N_6698);
nor U9032 (N_9032,N_7238,N_6150);
nand U9033 (N_9033,N_7897,N_7248);
nand U9034 (N_9034,N_7188,N_6541);
nor U9035 (N_9035,N_7063,N_6664);
nor U9036 (N_9036,N_7826,N_7724);
nand U9037 (N_9037,N_6567,N_6025);
or U9038 (N_9038,N_6042,N_7674);
nor U9039 (N_9039,N_6370,N_7853);
or U9040 (N_9040,N_7366,N_7056);
nor U9041 (N_9041,N_7311,N_7793);
or U9042 (N_9042,N_7111,N_7799);
and U9043 (N_9043,N_7036,N_6605);
and U9044 (N_9044,N_6351,N_6030);
or U9045 (N_9045,N_6662,N_7381);
nor U9046 (N_9046,N_7808,N_7663);
and U9047 (N_9047,N_6416,N_6151);
and U9048 (N_9048,N_7880,N_7312);
xnor U9049 (N_9049,N_6645,N_6759);
nor U9050 (N_9050,N_7856,N_6566);
nand U9051 (N_9051,N_7352,N_6827);
or U9052 (N_9052,N_6231,N_6822);
nor U9053 (N_9053,N_6484,N_6895);
and U9054 (N_9054,N_6725,N_7796);
nand U9055 (N_9055,N_6860,N_7782);
nand U9056 (N_9056,N_7169,N_7420);
nand U9057 (N_9057,N_6725,N_6812);
and U9058 (N_9058,N_6908,N_7837);
and U9059 (N_9059,N_6801,N_7109);
nand U9060 (N_9060,N_6434,N_7386);
nor U9061 (N_9061,N_6750,N_6703);
or U9062 (N_9062,N_7317,N_7720);
or U9063 (N_9063,N_6039,N_7389);
nor U9064 (N_9064,N_7065,N_6755);
and U9065 (N_9065,N_7404,N_6493);
or U9066 (N_9066,N_6473,N_6135);
nor U9067 (N_9067,N_7549,N_7710);
nand U9068 (N_9068,N_6386,N_6125);
nand U9069 (N_9069,N_7577,N_6003);
or U9070 (N_9070,N_6708,N_7072);
nand U9071 (N_9071,N_7008,N_7913);
and U9072 (N_9072,N_6962,N_7883);
nand U9073 (N_9073,N_6446,N_6411);
or U9074 (N_9074,N_7510,N_6033);
and U9075 (N_9075,N_7247,N_7444);
and U9076 (N_9076,N_6533,N_7131);
nand U9077 (N_9077,N_6050,N_6144);
or U9078 (N_9078,N_7258,N_6386);
and U9079 (N_9079,N_6791,N_6618);
nor U9080 (N_9080,N_6297,N_6844);
or U9081 (N_9081,N_6238,N_7664);
nor U9082 (N_9082,N_7827,N_7895);
nor U9083 (N_9083,N_7187,N_7701);
nor U9084 (N_9084,N_7434,N_6369);
or U9085 (N_9085,N_7711,N_6139);
and U9086 (N_9086,N_6404,N_7814);
and U9087 (N_9087,N_7330,N_6728);
nor U9088 (N_9088,N_6013,N_7943);
nor U9089 (N_9089,N_7438,N_7784);
and U9090 (N_9090,N_7803,N_6665);
or U9091 (N_9091,N_6621,N_6223);
xor U9092 (N_9092,N_6279,N_6194);
nand U9093 (N_9093,N_7901,N_7188);
and U9094 (N_9094,N_7416,N_7266);
nand U9095 (N_9095,N_6850,N_7847);
xor U9096 (N_9096,N_7736,N_6500);
and U9097 (N_9097,N_7616,N_6094);
nor U9098 (N_9098,N_6413,N_6149);
or U9099 (N_9099,N_6202,N_6970);
nand U9100 (N_9100,N_7008,N_7986);
nand U9101 (N_9101,N_7108,N_7187);
nor U9102 (N_9102,N_7728,N_6271);
nand U9103 (N_9103,N_6445,N_7308);
nor U9104 (N_9104,N_7927,N_7859);
and U9105 (N_9105,N_7418,N_7298);
nand U9106 (N_9106,N_6984,N_6206);
nand U9107 (N_9107,N_7201,N_7211);
or U9108 (N_9108,N_7973,N_7425);
or U9109 (N_9109,N_6329,N_7581);
or U9110 (N_9110,N_7455,N_7268);
or U9111 (N_9111,N_7497,N_6290);
and U9112 (N_9112,N_7454,N_6342);
nand U9113 (N_9113,N_6064,N_7616);
or U9114 (N_9114,N_6740,N_6882);
or U9115 (N_9115,N_6437,N_7707);
and U9116 (N_9116,N_6666,N_6384);
and U9117 (N_9117,N_6770,N_7944);
nor U9118 (N_9118,N_7570,N_6153);
or U9119 (N_9119,N_6416,N_7165);
nand U9120 (N_9120,N_7379,N_6578);
and U9121 (N_9121,N_6476,N_7573);
and U9122 (N_9122,N_6189,N_6082);
and U9123 (N_9123,N_7613,N_7295);
or U9124 (N_9124,N_7745,N_7587);
nor U9125 (N_9125,N_7145,N_7067);
and U9126 (N_9126,N_6834,N_7785);
and U9127 (N_9127,N_6111,N_7900);
or U9128 (N_9128,N_7712,N_7377);
and U9129 (N_9129,N_7192,N_6441);
or U9130 (N_9130,N_7372,N_6715);
or U9131 (N_9131,N_7770,N_7682);
nand U9132 (N_9132,N_7894,N_6303);
and U9133 (N_9133,N_7506,N_6470);
or U9134 (N_9134,N_6639,N_7737);
nor U9135 (N_9135,N_7351,N_7397);
and U9136 (N_9136,N_6416,N_6176);
nand U9137 (N_9137,N_7407,N_6184);
or U9138 (N_9138,N_6626,N_6886);
and U9139 (N_9139,N_7876,N_7121);
nor U9140 (N_9140,N_6423,N_6365);
and U9141 (N_9141,N_6879,N_7947);
nand U9142 (N_9142,N_6228,N_6906);
nor U9143 (N_9143,N_7316,N_6237);
nor U9144 (N_9144,N_7899,N_6207);
and U9145 (N_9145,N_7762,N_7790);
and U9146 (N_9146,N_6158,N_7762);
nand U9147 (N_9147,N_6505,N_7718);
and U9148 (N_9148,N_6208,N_6578);
and U9149 (N_9149,N_6054,N_6325);
and U9150 (N_9150,N_7405,N_6283);
nor U9151 (N_9151,N_6354,N_7241);
or U9152 (N_9152,N_6768,N_6615);
or U9153 (N_9153,N_7789,N_6647);
and U9154 (N_9154,N_6980,N_7015);
nor U9155 (N_9155,N_6833,N_6306);
or U9156 (N_9156,N_7155,N_7893);
or U9157 (N_9157,N_6265,N_7148);
nor U9158 (N_9158,N_7481,N_6034);
nor U9159 (N_9159,N_6718,N_6133);
and U9160 (N_9160,N_7239,N_6071);
xnor U9161 (N_9161,N_6726,N_6384);
and U9162 (N_9162,N_7630,N_7662);
and U9163 (N_9163,N_6414,N_6822);
nor U9164 (N_9164,N_6489,N_7703);
and U9165 (N_9165,N_6318,N_7084);
xnor U9166 (N_9166,N_6933,N_7316);
or U9167 (N_9167,N_6362,N_6448);
nand U9168 (N_9168,N_7623,N_7721);
nor U9169 (N_9169,N_7018,N_7795);
nand U9170 (N_9170,N_6438,N_7428);
nand U9171 (N_9171,N_7442,N_6596);
or U9172 (N_9172,N_6902,N_7164);
or U9173 (N_9173,N_6253,N_6692);
and U9174 (N_9174,N_7911,N_7883);
and U9175 (N_9175,N_6889,N_7776);
and U9176 (N_9176,N_7779,N_7570);
nand U9177 (N_9177,N_6116,N_6697);
nor U9178 (N_9178,N_6742,N_7592);
nand U9179 (N_9179,N_6045,N_6465);
and U9180 (N_9180,N_7945,N_7487);
or U9181 (N_9181,N_6538,N_6009);
nor U9182 (N_9182,N_6252,N_6894);
nor U9183 (N_9183,N_7637,N_7285);
or U9184 (N_9184,N_6183,N_6767);
nor U9185 (N_9185,N_6491,N_6526);
and U9186 (N_9186,N_6676,N_6108);
nand U9187 (N_9187,N_7142,N_7528);
nand U9188 (N_9188,N_6125,N_7794);
nand U9189 (N_9189,N_7936,N_7122);
nor U9190 (N_9190,N_6505,N_7620);
or U9191 (N_9191,N_7034,N_7713);
and U9192 (N_9192,N_7303,N_6395);
nor U9193 (N_9193,N_7569,N_7538);
nor U9194 (N_9194,N_6535,N_6921);
and U9195 (N_9195,N_6484,N_6055);
nor U9196 (N_9196,N_6288,N_7595);
and U9197 (N_9197,N_6337,N_6424);
nand U9198 (N_9198,N_6329,N_7782);
or U9199 (N_9199,N_6160,N_6326);
nand U9200 (N_9200,N_7731,N_7387);
nor U9201 (N_9201,N_7030,N_7511);
nor U9202 (N_9202,N_7964,N_6720);
nor U9203 (N_9203,N_7528,N_6483);
and U9204 (N_9204,N_7573,N_6295);
nor U9205 (N_9205,N_7585,N_6188);
nor U9206 (N_9206,N_7515,N_6908);
or U9207 (N_9207,N_7462,N_7568);
and U9208 (N_9208,N_7185,N_7211);
or U9209 (N_9209,N_6733,N_6034);
or U9210 (N_9210,N_6106,N_6728);
or U9211 (N_9211,N_6000,N_7188);
or U9212 (N_9212,N_6432,N_6894);
nor U9213 (N_9213,N_6421,N_7788);
nor U9214 (N_9214,N_7856,N_7075);
or U9215 (N_9215,N_6914,N_6046);
nor U9216 (N_9216,N_7622,N_6731);
nand U9217 (N_9217,N_6519,N_7992);
and U9218 (N_9218,N_6387,N_7539);
nor U9219 (N_9219,N_6619,N_7318);
nor U9220 (N_9220,N_6084,N_6712);
and U9221 (N_9221,N_6260,N_6486);
nor U9222 (N_9222,N_7566,N_7234);
and U9223 (N_9223,N_7070,N_6454);
and U9224 (N_9224,N_7706,N_7024);
and U9225 (N_9225,N_7230,N_7488);
and U9226 (N_9226,N_7725,N_6237);
and U9227 (N_9227,N_6807,N_7529);
or U9228 (N_9228,N_6059,N_6815);
and U9229 (N_9229,N_6832,N_7645);
or U9230 (N_9230,N_6478,N_7693);
nor U9231 (N_9231,N_7901,N_6071);
nand U9232 (N_9232,N_7698,N_6748);
nand U9233 (N_9233,N_6610,N_6646);
or U9234 (N_9234,N_6301,N_6176);
nor U9235 (N_9235,N_7595,N_6483);
and U9236 (N_9236,N_7946,N_6511);
and U9237 (N_9237,N_6756,N_6885);
nor U9238 (N_9238,N_6029,N_7509);
and U9239 (N_9239,N_7247,N_7367);
nor U9240 (N_9240,N_7587,N_7201);
nand U9241 (N_9241,N_6932,N_7829);
nor U9242 (N_9242,N_7985,N_6687);
nand U9243 (N_9243,N_6485,N_6255);
nor U9244 (N_9244,N_7832,N_7831);
nand U9245 (N_9245,N_7878,N_7410);
nor U9246 (N_9246,N_6453,N_7493);
nand U9247 (N_9247,N_6789,N_7651);
nand U9248 (N_9248,N_7233,N_6582);
nor U9249 (N_9249,N_6425,N_6847);
or U9250 (N_9250,N_6746,N_7280);
and U9251 (N_9251,N_7702,N_6545);
or U9252 (N_9252,N_6448,N_6467);
or U9253 (N_9253,N_7841,N_7566);
or U9254 (N_9254,N_7107,N_6042);
and U9255 (N_9255,N_6230,N_6878);
and U9256 (N_9256,N_6786,N_6088);
or U9257 (N_9257,N_7929,N_6096);
nor U9258 (N_9258,N_7077,N_6924);
nand U9259 (N_9259,N_6633,N_7178);
or U9260 (N_9260,N_7772,N_7743);
nand U9261 (N_9261,N_6561,N_6202);
and U9262 (N_9262,N_7861,N_6286);
or U9263 (N_9263,N_6240,N_6634);
and U9264 (N_9264,N_6233,N_6415);
nor U9265 (N_9265,N_6690,N_7409);
and U9266 (N_9266,N_6699,N_6880);
nor U9267 (N_9267,N_6542,N_7376);
xor U9268 (N_9268,N_7059,N_7555);
or U9269 (N_9269,N_6324,N_7770);
and U9270 (N_9270,N_6278,N_6570);
or U9271 (N_9271,N_6391,N_6708);
nand U9272 (N_9272,N_7551,N_6146);
nand U9273 (N_9273,N_6299,N_7377);
nand U9274 (N_9274,N_7250,N_7973);
or U9275 (N_9275,N_7815,N_7904);
or U9276 (N_9276,N_7960,N_7592);
or U9277 (N_9277,N_7955,N_7887);
and U9278 (N_9278,N_6292,N_7360);
nor U9279 (N_9279,N_7911,N_6880);
and U9280 (N_9280,N_7010,N_7784);
and U9281 (N_9281,N_7060,N_6740);
or U9282 (N_9282,N_6934,N_6001);
nand U9283 (N_9283,N_6101,N_6837);
nand U9284 (N_9284,N_6642,N_6712);
and U9285 (N_9285,N_7585,N_6693);
and U9286 (N_9286,N_7822,N_6075);
xor U9287 (N_9287,N_6288,N_7520);
or U9288 (N_9288,N_7122,N_6304);
nor U9289 (N_9289,N_7785,N_6984);
and U9290 (N_9290,N_7491,N_6403);
or U9291 (N_9291,N_7374,N_7013);
nand U9292 (N_9292,N_7536,N_7620);
and U9293 (N_9293,N_7551,N_7464);
nor U9294 (N_9294,N_6086,N_7849);
nor U9295 (N_9295,N_7662,N_6287);
or U9296 (N_9296,N_7627,N_6802);
nor U9297 (N_9297,N_7144,N_7867);
xnor U9298 (N_9298,N_7405,N_6361);
nor U9299 (N_9299,N_7176,N_6496);
xor U9300 (N_9300,N_7822,N_7860);
and U9301 (N_9301,N_7828,N_7722);
nand U9302 (N_9302,N_6166,N_7391);
xor U9303 (N_9303,N_7003,N_7045);
and U9304 (N_9304,N_6226,N_6707);
nor U9305 (N_9305,N_7633,N_6068);
xnor U9306 (N_9306,N_7658,N_6221);
or U9307 (N_9307,N_7745,N_6451);
nand U9308 (N_9308,N_6496,N_6916);
nor U9309 (N_9309,N_7848,N_7342);
nor U9310 (N_9310,N_6027,N_7143);
or U9311 (N_9311,N_7970,N_7295);
or U9312 (N_9312,N_7456,N_6871);
nor U9313 (N_9313,N_6367,N_7471);
nand U9314 (N_9314,N_7205,N_6198);
and U9315 (N_9315,N_7907,N_6303);
nand U9316 (N_9316,N_7923,N_7959);
nand U9317 (N_9317,N_6939,N_6284);
or U9318 (N_9318,N_6043,N_6285);
nand U9319 (N_9319,N_6415,N_6409);
and U9320 (N_9320,N_7323,N_7254);
nand U9321 (N_9321,N_7363,N_7203);
and U9322 (N_9322,N_7950,N_6461);
or U9323 (N_9323,N_7199,N_7854);
and U9324 (N_9324,N_7425,N_6878);
and U9325 (N_9325,N_6841,N_6929);
or U9326 (N_9326,N_7676,N_6620);
nor U9327 (N_9327,N_6357,N_7814);
and U9328 (N_9328,N_6675,N_6040);
and U9329 (N_9329,N_7369,N_7946);
nor U9330 (N_9330,N_6717,N_7916);
and U9331 (N_9331,N_6603,N_7787);
or U9332 (N_9332,N_6536,N_7013);
nor U9333 (N_9333,N_7310,N_6154);
and U9334 (N_9334,N_6788,N_7892);
or U9335 (N_9335,N_6834,N_6666);
nand U9336 (N_9336,N_7063,N_7292);
nand U9337 (N_9337,N_7466,N_6423);
nand U9338 (N_9338,N_6302,N_7365);
or U9339 (N_9339,N_6522,N_6434);
or U9340 (N_9340,N_6614,N_6292);
or U9341 (N_9341,N_6611,N_7751);
nor U9342 (N_9342,N_6240,N_7627);
nand U9343 (N_9343,N_6467,N_6965);
nor U9344 (N_9344,N_7586,N_7546);
and U9345 (N_9345,N_7533,N_7110);
nand U9346 (N_9346,N_6404,N_6737);
nor U9347 (N_9347,N_6303,N_7793);
nand U9348 (N_9348,N_6706,N_7174);
nand U9349 (N_9349,N_6828,N_6659);
nor U9350 (N_9350,N_6236,N_7326);
nor U9351 (N_9351,N_7791,N_7268);
and U9352 (N_9352,N_7177,N_7776);
or U9353 (N_9353,N_6816,N_6173);
xor U9354 (N_9354,N_7206,N_7981);
nand U9355 (N_9355,N_7542,N_6593);
or U9356 (N_9356,N_6794,N_6570);
nand U9357 (N_9357,N_6766,N_6712);
or U9358 (N_9358,N_6094,N_6511);
and U9359 (N_9359,N_7519,N_7868);
and U9360 (N_9360,N_7828,N_6666);
and U9361 (N_9361,N_6364,N_7468);
or U9362 (N_9362,N_7724,N_7593);
or U9363 (N_9363,N_6266,N_6277);
and U9364 (N_9364,N_7003,N_6876);
or U9365 (N_9365,N_6372,N_7215);
and U9366 (N_9366,N_7786,N_7524);
and U9367 (N_9367,N_6442,N_7071);
nor U9368 (N_9368,N_7172,N_7036);
nor U9369 (N_9369,N_7832,N_6591);
nand U9370 (N_9370,N_7196,N_7804);
nand U9371 (N_9371,N_7966,N_6545);
nand U9372 (N_9372,N_6121,N_6312);
nor U9373 (N_9373,N_7701,N_6536);
or U9374 (N_9374,N_6278,N_6329);
and U9375 (N_9375,N_7177,N_6698);
or U9376 (N_9376,N_6867,N_7242);
nor U9377 (N_9377,N_6441,N_6440);
nand U9378 (N_9378,N_6888,N_7183);
nand U9379 (N_9379,N_7342,N_7657);
and U9380 (N_9380,N_7061,N_7767);
and U9381 (N_9381,N_7035,N_6013);
nor U9382 (N_9382,N_6917,N_7559);
nand U9383 (N_9383,N_6124,N_6789);
nand U9384 (N_9384,N_7255,N_6839);
and U9385 (N_9385,N_7675,N_7849);
xnor U9386 (N_9386,N_6076,N_6922);
or U9387 (N_9387,N_7829,N_6038);
xor U9388 (N_9388,N_7766,N_6631);
nor U9389 (N_9389,N_7199,N_6682);
nand U9390 (N_9390,N_7845,N_7289);
nand U9391 (N_9391,N_7928,N_6069);
or U9392 (N_9392,N_6495,N_7141);
nor U9393 (N_9393,N_7835,N_7104);
nand U9394 (N_9394,N_7710,N_7895);
or U9395 (N_9395,N_6067,N_7735);
xor U9396 (N_9396,N_7903,N_6896);
or U9397 (N_9397,N_7612,N_7486);
nand U9398 (N_9398,N_7245,N_7349);
and U9399 (N_9399,N_7404,N_6537);
nand U9400 (N_9400,N_7360,N_7648);
and U9401 (N_9401,N_6068,N_6148);
nand U9402 (N_9402,N_6001,N_7088);
or U9403 (N_9403,N_6426,N_6785);
nor U9404 (N_9404,N_7293,N_7963);
and U9405 (N_9405,N_6513,N_6635);
xnor U9406 (N_9406,N_6635,N_6351);
nor U9407 (N_9407,N_7672,N_7638);
or U9408 (N_9408,N_7596,N_6603);
nor U9409 (N_9409,N_6365,N_6458);
nor U9410 (N_9410,N_7769,N_6554);
nor U9411 (N_9411,N_7915,N_6599);
or U9412 (N_9412,N_6166,N_6419);
nand U9413 (N_9413,N_7297,N_7204);
and U9414 (N_9414,N_7398,N_7622);
and U9415 (N_9415,N_7907,N_6326);
or U9416 (N_9416,N_7963,N_6145);
nor U9417 (N_9417,N_7396,N_7404);
and U9418 (N_9418,N_7905,N_7649);
nor U9419 (N_9419,N_7799,N_7753);
or U9420 (N_9420,N_6357,N_6946);
or U9421 (N_9421,N_7359,N_7198);
nor U9422 (N_9422,N_6394,N_7435);
nand U9423 (N_9423,N_6248,N_7326);
nand U9424 (N_9424,N_7039,N_7338);
or U9425 (N_9425,N_7274,N_7624);
nand U9426 (N_9426,N_7156,N_7851);
or U9427 (N_9427,N_7023,N_6913);
nor U9428 (N_9428,N_7132,N_6479);
nand U9429 (N_9429,N_7980,N_6233);
or U9430 (N_9430,N_6858,N_7172);
and U9431 (N_9431,N_7837,N_6476);
and U9432 (N_9432,N_7021,N_7475);
nor U9433 (N_9433,N_7781,N_6907);
or U9434 (N_9434,N_7330,N_6547);
nor U9435 (N_9435,N_7663,N_6383);
nand U9436 (N_9436,N_6713,N_6042);
nor U9437 (N_9437,N_6462,N_6194);
nor U9438 (N_9438,N_6822,N_7197);
or U9439 (N_9439,N_6949,N_7160);
or U9440 (N_9440,N_7168,N_6745);
nand U9441 (N_9441,N_6373,N_6071);
nand U9442 (N_9442,N_7441,N_6946);
xor U9443 (N_9443,N_7133,N_7726);
and U9444 (N_9444,N_6811,N_7469);
nor U9445 (N_9445,N_7867,N_6862);
nand U9446 (N_9446,N_7166,N_6055);
and U9447 (N_9447,N_7035,N_6284);
and U9448 (N_9448,N_6235,N_6302);
and U9449 (N_9449,N_7890,N_6418);
or U9450 (N_9450,N_6510,N_7642);
or U9451 (N_9451,N_7263,N_7401);
nor U9452 (N_9452,N_6061,N_6161);
nor U9453 (N_9453,N_6742,N_7122);
nor U9454 (N_9454,N_7372,N_7171);
nor U9455 (N_9455,N_6692,N_6257);
or U9456 (N_9456,N_6915,N_6452);
and U9457 (N_9457,N_7098,N_7172);
and U9458 (N_9458,N_7788,N_6098);
nor U9459 (N_9459,N_7250,N_6068);
or U9460 (N_9460,N_7665,N_6607);
nor U9461 (N_9461,N_6607,N_6228);
or U9462 (N_9462,N_7642,N_7491);
nor U9463 (N_9463,N_7812,N_7441);
nor U9464 (N_9464,N_6145,N_6053);
or U9465 (N_9465,N_6196,N_7575);
nand U9466 (N_9466,N_6902,N_6816);
nand U9467 (N_9467,N_7414,N_6035);
nand U9468 (N_9468,N_6468,N_7905);
nand U9469 (N_9469,N_6296,N_7884);
and U9470 (N_9470,N_6549,N_6849);
or U9471 (N_9471,N_6463,N_6271);
or U9472 (N_9472,N_6321,N_6252);
or U9473 (N_9473,N_6174,N_7227);
or U9474 (N_9474,N_7719,N_7268);
nand U9475 (N_9475,N_7077,N_7550);
nand U9476 (N_9476,N_7372,N_7476);
or U9477 (N_9477,N_6863,N_6017);
or U9478 (N_9478,N_6411,N_7908);
and U9479 (N_9479,N_7400,N_6569);
nor U9480 (N_9480,N_6540,N_6155);
and U9481 (N_9481,N_7221,N_7037);
or U9482 (N_9482,N_7210,N_7765);
and U9483 (N_9483,N_7564,N_7553);
or U9484 (N_9484,N_7211,N_6032);
and U9485 (N_9485,N_7670,N_7569);
and U9486 (N_9486,N_7028,N_6321);
nor U9487 (N_9487,N_6800,N_7418);
and U9488 (N_9488,N_6031,N_7583);
nand U9489 (N_9489,N_6356,N_6009);
and U9490 (N_9490,N_7883,N_6696);
nand U9491 (N_9491,N_7483,N_7190);
nand U9492 (N_9492,N_6296,N_6765);
and U9493 (N_9493,N_6386,N_6344);
nor U9494 (N_9494,N_7112,N_7243);
and U9495 (N_9495,N_6361,N_6916);
and U9496 (N_9496,N_7724,N_7380);
nand U9497 (N_9497,N_7512,N_6461);
and U9498 (N_9498,N_7826,N_6228);
or U9499 (N_9499,N_7058,N_6033);
nor U9500 (N_9500,N_7328,N_7186);
nor U9501 (N_9501,N_7257,N_7972);
nor U9502 (N_9502,N_6909,N_7345);
nand U9503 (N_9503,N_7838,N_7401);
or U9504 (N_9504,N_6787,N_6283);
and U9505 (N_9505,N_6051,N_7458);
nand U9506 (N_9506,N_6123,N_6577);
nand U9507 (N_9507,N_7159,N_6148);
nor U9508 (N_9508,N_6812,N_6607);
nand U9509 (N_9509,N_7738,N_7831);
nor U9510 (N_9510,N_6207,N_6916);
or U9511 (N_9511,N_6058,N_6143);
nor U9512 (N_9512,N_6789,N_6217);
and U9513 (N_9513,N_7487,N_7661);
nand U9514 (N_9514,N_6941,N_6705);
nor U9515 (N_9515,N_7398,N_6380);
and U9516 (N_9516,N_7847,N_7192);
nor U9517 (N_9517,N_7501,N_6355);
and U9518 (N_9518,N_6493,N_7791);
and U9519 (N_9519,N_6817,N_7837);
nor U9520 (N_9520,N_7775,N_6711);
and U9521 (N_9521,N_7721,N_7119);
and U9522 (N_9522,N_6351,N_7224);
nor U9523 (N_9523,N_6500,N_7717);
nand U9524 (N_9524,N_6788,N_6503);
and U9525 (N_9525,N_7451,N_6788);
nand U9526 (N_9526,N_6098,N_7242);
nand U9527 (N_9527,N_6275,N_7902);
and U9528 (N_9528,N_7719,N_7370);
and U9529 (N_9529,N_6490,N_7842);
nand U9530 (N_9530,N_6935,N_6637);
nor U9531 (N_9531,N_7444,N_7850);
and U9532 (N_9532,N_7388,N_6345);
nand U9533 (N_9533,N_6674,N_6172);
or U9534 (N_9534,N_6411,N_6616);
nand U9535 (N_9535,N_7316,N_6767);
nand U9536 (N_9536,N_6159,N_6632);
nor U9537 (N_9537,N_7955,N_7016);
or U9538 (N_9538,N_7686,N_6337);
nor U9539 (N_9539,N_6481,N_7985);
nand U9540 (N_9540,N_6116,N_7471);
nor U9541 (N_9541,N_7061,N_6606);
nor U9542 (N_9542,N_7461,N_7755);
nor U9543 (N_9543,N_6676,N_7029);
nor U9544 (N_9544,N_6420,N_7798);
nor U9545 (N_9545,N_7515,N_7410);
or U9546 (N_9546,N_7528,N_6087);
or U9547 (N_9547,N_6578,N_7625);
and U9548 (N_9548,N_6474,N_6790);
nand U9549 (N_9549,N_6335,N_7143);
nand U9550 (N_9550,N_6178,N_6575);
and U9551 (N_9551,N_6717,N_7040);
and U9552 (N_9552,N_6684,N_7759);
nor U9553 (N_9553,N_6384,N_7472);
nor U9554 (N_9554,N_6377,N_6445);
or U9555 (N_9555,N_7132,N_6626);
or U9556 (N_9556,N_7152,N_6807);
nor U9557 (N_9557,N_7892,N_7168);
or U9558 (N_9558,N_6537,N_6594);
or U9559 (N_9559,N_7397,N_7452);
xnor U9560 (N_9560,N_6357,N_6545);
nand U9561 (N_9561,N_7878,N_7078);
nor U9562 (N_9562,N_7876,N_7116);
nor U9563 (N_9563,N_7467,N_6816);
and U9564 (N_9564,N_6239,N_6076);
nor U9565 (N_9565,N_7600,N_6730);
nor U9566 (N_9566,N_7000,N_7505);
and U9567 (N_9567,N_7583,N_6417);
and U9568 (N_9568,N_7476,N_6960);
or U9569 (N_9569,N_6228,N_6224);
nand U9570 (N_9570,N_6950,N_7892);
and U9571 (N_9571,N_7388,N_6955);
or U9572 (N_9572,N_7459,N_7230);
nand U9573 (N_9573,N_6560,N_6937);
nor U9574 (N_9574,N_7530,N_7568);
and U9575 (N_9575,N_7145,N_6133);
or U9576 (N_9576,N_7199,N_6267);
xor U9577 (N_9577,N_6523,N_6997);
nor U9578 (N_9578,N_6386,N_6478);
nor U9579 (N_9579,N_7256,N_6575);
or U9580 (N_9580,N_6134,N_6040);
nor U9581 (N_9581,N_6304,N_7862);
nor U9582 (N_9582,N_7378,N_7693);
and U9583 (N_9583,N_7822,N_6122);
and U9584 (N_9584,N_6499,N_7096);
and U9585 (N_9585,N_6456,N_6920);
nand U9586 (N_9586,N_7108,N_7266);
nor U9587 (N_9587,N_7654,N_7963);
nand U9588 (N_9588,N_7944,N_6937);
and U9589 (N_9589,N_7492,N_6550);
nand U9590 (N_9590,N_7323,N_7400);
or U9591 (N_9591,N_7543,N_6669);
nand U9592 (N_9592,N_7684,N_6067);
nand U9593 (N_9593,N_7385,N_6129);
and U9594 (N_9594,N_7710,N_6696);
and U9595 (N_9595,N_7888,N_6460);
or U9596 (N_9596,N_6885,N_6732);
and U9597 (N_9597,N_7875,N_7301);
nand U9598 (N_9598,N_7275,N_6938);
nor U9599 (N_9599,N_6169,N_7116);
nor U9600 (N_9600,N_6875,N_6578);
nand U9601 (N_9601,N_7830,N_7013);
or U9602 (N_9602,N_7585,N_6199);
and U9603 (N_9603,N_6258,N_6606);
nand U9604 (N_9604,N_6560,N_6588);
nand U9605 (N_9605,N_7400,N_6502);
and U9606 (N_9606,N_7270,N_7787);
and U9607 (N_9607,N_6075,N_6273);
and U9608 (N_9608,N_6325,N_7218);
or U9609 (N_9609,N_7050,N_7973);
or U9610 (N_9610,N_6234,N_6976);
nand U9611 (N_9611,N_7097,N_7646);
nor U9612 (N_9612,N_7714,N_7723);
nor U9613 (N_9613,N_7272,N_7637);
or U9614 (N_9614,N_7992,N_6802);
and U9615 (N_9615,N_7992,N_6514);
or U9616 (N_9616,N_7606,N_6209);
and U9617 (N_9617,N_7077,N_6404);
nor U9618 (N_9618,N_6876,N_6846);
or U9619 (N_9619,N_6963,N_7994);
nand U9620 (N_9620,N_7805,N_7015);
nor U9621 (N_9621,N_6429,N_7032);
or U9622 (N_9622,N_7119,N_7704);
nand U9623 (N_9623,N_7953,N_6002);
nand U9624 (N_9624,N_7385,N_6514);
and U9625 (N_9625,N_7024,N_7450);
or U9626 (N_9626,N_6666,N_6601);
nand U9627 (N_9627,N_6910,N_7070);
or U9628 (N_9628,N_7860,N_7683);
nor U9629 (N_9629,N_7452,N_7840);
or U9630 (N_9630,N_6984,N_7513);
and U9631 (N_9631,N_7206,N_6938);
or U9632 (N_9632,N_6938,N_7309);
or U9633 (N_9633,N_7019,N_6706);
or U9634 (N_9634,N_7779,N_6769);
or U9635 (N_9635,N_7992,N_7234);
nand U9636 (N_9636,N_6284,N_6944);
nor U9637 (N_9637,N_6805,N_7182);
nor U9638 (N_9638,N_6451,N_6435);
nand U9639 (N_9639,N_7210,N_7345);
or U9640 (N_9640,N_7820,N_6721);
nand U9641 (N_9641,N_6616,N_6691);
or U9642 (N_9642,N_6935,N_6647);
nor U9643 (N_9643,N_6972,N_7519);
nand U9644 (N_9644,N_7769,N_7012);
nand U9645 (N_9645,N_7885,N_7008);
nor U9646 (N_9646,N_7677,N_6252);
and U9647 (N_9647,N_7846,N_7722);
and U9648 (N_9648,N_6265,N_6831);
and U9649 (N_9649,N_6989,N_6682);
or U9650 (N_9650,N_6563,N_7931);
or U9651 (N_9651,N_7295,N_6014);
nand U9652 (N_9652,N_7905,N_7468);
and U9653 (N_9653,N_6581,N_7464);
and U9654 (N_9654,N_7030,N_6940);
nand U9655 (N_9655,N_7690,N_7768);
nand U9656 (N_9656,N_7898,N_6040);
or U9657 (N_9657,N_7485,N_7210);
and U9658 (N_9658,N_7351,N_6288);
or U9659 (N_9659,N_6289,N_7496);
and U9660 (N_9660,N_7226,N_7268);
or U9661 (N_9661,N_7510,N_7589);
or U9662 (N_9662,N_6005,N_6014);
and U9663 (N_9663,N_6264,N_6077);
nand U9664 (N_9664,N_7573,N_6381);
nand U9665 (N_9665,N_6847,N_6915);
and U9666 (N_9666,N_6624,N_7266);
or U9667 (N_9667,N_7554,N_7183);
nor U9668 (N_9668,N_7721,N_7050);
and U9669 (N_9669,N_6220,N_6157);
or U9670 (N_9670,N_7327,N_6153);
or U9671 (N_9671,N_6683,N_7197);
xor U9672 (N_9672,N_6569,N_7924);
nor U9673 (N_9673,N_7704,N_6860);
nand U9674 (N_9674,N_7354,N_6000);
nor U9675 (N_9675,N_6591,N_7416);
or U9676 (N_9676,N_6722,N_6428);
nand U9677 (N_9677,N_6963,N_6481);
or U9678 (N_9678,N_6733,N_6818);
nor U9679 (N_9679,N_7386,N_7315);
or U9680 (N_9680,N_7883,N_6080);
nand U9681 (N_9681,N_6883,N_6046);
nand U9682 (N_9682,N_7669,N_6284);
nand U9683 (N_9683,N_7481,N_6585);
and U9684 (N_9684,N_6607,N_6507);
or U9685 (N_9685,N_6279,N_7265);
nor U9686 (N_9686,N_7603,N_6703);
nand U9687 (N_9687,N_6933,N_6959);
nand U9688 (N_9688,N_7148,N_7458);
nor U9689 (N_9689,N_6405,N_7470);
or U9690 (N_9690,N_6018,N_6908);
nor U9691 (N_9691,N_6708,N_6939);
xnor U9692 (N_9692,N_6466,N_7148);
nand U9693 (N_9693,N_6948,N_7363);
nand U9694 (N_9694,N_6349,N_7533);
xnor U9695 (N_9695,N_6906,N_6811);
or U9696 (N_9696,N_6565,N_6117);
or U9697 (N_9697,N_6266,N_6589);
nand U9698 (N_9698,N_6621,N_7314);
nand U9699 (N_9699,N_7220,N_7223);
and U9700 (N_9700,N_7264,N_7811);
nand U9701 (N_9701,N_7142,N_7205);
and U9702 (N_9702,N_6954,N_6309);
nor U9703 (N_9703,N_7896,N_6801);
or U9704 (N_9704,N_6451,N_7074);
or U9705 (N_9705,N_6189,N_6705);
nor U9706 (N_9706,N_6631,N_6949);
nand U9707 (N_9707,N_7910,N_7490);
and U9708 (N_9708,N_6615,N_6808);
or U9709 (N_9709,N_6561,N_6994);
xnor U9710 (N_9710,N_7560,N_7475);
nand U9711 (N_9711,N_7802,N_7250);
nand U9712 (N_9712,N_7051,N_7454);
and U9713 (N_9713,N_7670,N_6775);
nor U9714 (N_9714,N_6178,N_6631);
and U9715 (N_9715,N_7562,N_6192);
or U9716 (N_9716,N_6231,N_6937);
nor U9717 (N_9717,N_7127,N_7982);
and U9718 (N_9718,N_7996,N_6335);
or U9719 (N_9719,N_6937,N_7975);
nor U9720 (N_9720,N_6308,N_7853);
or U9721 (N_9721,N_6362,N_7812);
xor U9722 (N_9722,N_6983,N_6687);
and U9723 (N_9723,N_6193,N_7007);
or U9724 (N_9724,N_7549,N_7221);
or U9725 (N_9725,N_7047,N_6470);
or U9726 (N_9726,N_7404,N_7335);
or U9727 (N_9727,N_7892,N_6595);
and U9728 (N_9728,N_7049,N_7941);
nor U9729 (N_9729,N_7524,N_7514);
and U9730 (N_9730,N_7461,N_7299);
nor U9731 (N_9731,N_7060,N_6272);
nor U9732 (N_9732,N_7346,N_7570);
or U9733 (N_9733,N_6366,N_7734);
or U9734 (N_9734,N_7986,N_7487);
nor U9735 (N_9735,N_7173,N_6809);
or U9736 (N_9736,N_6249,N_6485);
and U9737 (N_9737,N_7930,N_6004);
nand U9738 (N_9738,N_6637,N_7300);
nand U9739 (N_9739,N_6622,N_7230);
nor U9740 (N_9740,N_6213,N_6058);
and U9741 (N_9741,N_7276,N_6011);
and U9742 (N_9742,N_7753,N_6970);
or U9743 (N_9743,N_6227,N_7322);
nor U9744 (N_9744,N_6664,N_7664);
xnor U9745 (N_9745,N_7394,N_6636);
nor U9746 (N_9746,N_6963,N_6168);
and U9747 (N_9747,N_6700,N_6192);
or U9748 (N_9748,N_7585,N_7281);
and U9749 (N_9749,N_6332,N_6643);
nor U9750 (N_9750,N_7075,N_7139);
and U9751 (N_9751,N_7107,N_7579);
nand U9752 (N_9752,N_6768,N_6984);
xnor U9753 (N_9753,N_6609,N_7836);
nand U9754 (N_9754,N_6323,N_6497);
and U9755 (N_9755,N_7386,N_7395);
nand U9756 (N_9756,N_6394,N_7525);
nor U9757 (N_9757,N_7243,N_7207);
nand U9758 (N_9758,N_7252,N_6986);
or U9759 (N_9759,N_6173,N_6241);
nor U9760 (N_9760,N_6325,N_7875);
nor U9761 (N_9761,N_6784,N_7327);
and U9762 (N_9762,N_7534,N_6304);
nand U9763 (N_9763,N_6933,N_7859);
nor U9764 (N_9764,N_6219,N_6017);
nand U9765 (N_9765,N_6606,N_6266);
and U9766 (N_9766,N_7470,N_6099);
nor U9767 (N_9767,N_7832,N_7932);
xor U9768 (N_9768,N_6219,N_7519);
nor U9769 (N_9769,N_6486,N_7886);
nor U9770 (N_9770,N_6630,N_7315);
nand U9771 (N_9771,N_6876,N_6238);
nor U9772 (N_9772,N_6637,N_7987);
nor U9773 (N_9773,N_7434,N_7780);
nand U9774 (N_9774,N_7822,N_7618);
or U9775 (N_9775,N_6216,N_7309);
nor U9776 (N_9776,N_6824,N_7948);
nand U9777 (N_9777,N_7460,N_7965);
nor U9778 (N_9778,N_6351,N_7171);
or U9779 (N_9779,N_6958,N_7768);
nand U9780 (N_9780,N_6449,N_6407);
and U9781 (N_9781,N_6695,N_6707);
nor U9782 (N_9782,N_7672,N_7729);
and U9783 (N_9783,N_6319,N_6981);
nand U9784 (N_9784,N_7176,N_6704);
nand U9785 (N_9785,N_7139,N_7254);
and U9786 (N_9786,N_7446,N_7725);
and U9787 (N_9787,N_6168,N_7355);
or U9788 (N_9788,N_7369,N_7786);
nor U9789 (N_9789,N_7582,N_7400);
nand U9790 (N_9790,N_6820,N_7488);
or U9791 (N_9791,N_7482,N_6359);
nor U9792 (N_9792,N_6742,N_6169);
nor U9793 (N_9793,N_6516,N_7202);
and U9794 (N_9794,N_7317,N_7243);
nor U9795 (N_9795,N_6425,N_7273);
nor U9796 (N_9796,N_6404,N_7900);
or U9797 (N_9797,N_6294,N_7430);
nor U9798 (N_9798,N_6471,N_6212);
nand U9799 (N_9799,N_6498,N_7697);
and U9800 (N_9800,N_6332,N_7905);
xor U9801 (N_9801,N_6168,N_6248);
nand U9802 (N_9802,N_6177,N_7583);
and U9803 (N_9803,N_7068,N_7664);
or U9804 (N_9804,N_7738,N_6929);
and U9805 (N_9805,N_7662,N_6121);
nand U9806 (N_9806,N_6975,N_7507);
nor U9807 (N_9807,N_6998,N_6629);
nand U9808 (N_9808,N_7386,N_7050);
nor U9809 (N_9809,N_7260,N_6845);
and U9810 (N_9810,N_6206,N_6875);
nand U9811 (N_9811,N_6831,N_7893);
and U9812 (N_9812,N_6576,N_6488);
xnor U9813 (N_9813,N_6136,N_6764);
nand U9814 (N_9814,N_6644,N_6786);
or U9815 (N_9815,N_7543,N_7909);
xor U9816 (N_9816,N_6516,N_7816);
nand U9817 (N_9817,N_6898,N_6127);
or U9818 (N_9818,N_6252,N_6707);
nor U9819 (N_9819,N_6001,N_6332);
xor U9820 (N_9820,N_6742,N_7403);
nand U9821 (N_9821,N_6350,N_6937);
and U9822 (N_9822,N_7106,N_6055);
nor U9823 (N_9823,N_6496,N_6210);
nor U9824 (N_9824,N_7739,N_6554);
and U9825 (N_9825,N_6997,N_6585);
and U9826 (N_9826,N_6857,N_6075);
or U9827 (N_9827,N_6901,N_6913);
or U9828 (N_9828,N_6097,N_6353);
nand U9829 (N_9829,N_7278,N_6170);
or U9830 (N_9830,N_7177,N_6423);
nor U9831 (N_9831,N_6251,N_6242);
xnor U9832 (N_9832,N_6745,N_7143);
or U9833 (N_9833,N_7860,N_6514);
or U9834 (N_9834,N_7978,N_6480);
and U9835 (N_9835,N_6805,N_7303);
nand U9836 (N_9836,N_6394,N_6090);
and U9837 (N_9837,N_7840,N_6422);
nand U9838 (N_9838,N_6423,N_7827);
and U9839 (N_9839,N_6488,N_7198);
nand U9840 (N_9840,N_7062,N_6698);
or U9841 (N_9841,N_7229,N_7020);
nand U9842 (N_9842,N_7181,N_7858);
or U9843 (N_9843,N_6389,N_6822);
nor U9844 (N_9844,N_7315,N_7793);
nand U9845 (N_9845,N_6769,N_6050);
nand U9846 (N_9846,N_6336,N_7351);
or U9847 (N_9847,N_7492,N_6359);
nor U9848 (N_9848,N_7209,N_7217);
nor U9849 (N_9849,N_6489,N_7505);
and U9850 (N_9850,N_7645,N_6931);
or U9851 (N_9851,N_6046,N_6387);
and U9852 (N_9852,N_6765,N_7986);
nor U9853 (N_9853,N_6976,N_7455);
nand U9854 (N_9854,N_7017,N_6734);
nor U9855 (N_9855,N_7682,N_7766);
and U9856 (N_9856,N_6885,N_6778);
nand U9857 (N_9857,N_6744,N_6557);
xnor U9858 (N_9858,N_7969,N_6995);
and U9859 (N_9859,N_7167,N_7754);
and U9860 (N_9860,N_6281,N_6474);
or U9861 (N_9861,N_7823,N_6823);
nor U9862 (N_9862,N_7570,N_6747);
or U9863 (N_9863,N_7281,N_6594);
or U9864 (N_9864,N_6868,N_7208);
or U9865 (N_9865,N_6763,N_6326);
nand U9866 (N_9866,N_7742,N_7245);
and U9867 (N_9867,N_7619,N_7642);
or U9868 (N_9868,N_7665,N_6141);
nor U9869 (N_9869,N_7310,N_6903);
nand U9870 (N_9870,N_6032,N_6426);
nor U9871 (N_9871,N_6666,N_7922);
and U9872 (N_9872,N_7030,N_7399);
nand U9873 (N_9873,N_7237,N_7021);
nand U9874 (N_9874,N_6891,N_7051);
nor U9875 (N_9875,N_7251,N_7666);
or U9876 (N_9876,N_6682,N_7738);
or U9877 (N_9877,N_7912,N_6029);
nor U9878 (N_9878,N_7389,N_7371);
and U9879 (N_9879,N_7694,N_6706);
nand U9880 (N_9880,N_7768,N_7893);
nor U9881 (N_9881,N_6007,N_6311);
or U9882 (N_9882,N_6666,N_7557);
nand U9883 (N_9883,N_6639,N_7025);
nor U9884 (N_9884,N_6054,N_6160);
or U9885 (N_9885,N_6247,N_6502);
and U9886 (N_9886,N_6057,N_6393);
nand U9887 (N_9887,N_7515,N_6749);
nand U9888 (N_9888,N_6430,N_7361);
nand U9889 (N_9889,N_7297,N_7377);
nand U9890 (N_9890,N_6783,N_7414);
nand U9891 (N_9891,N_7446,N_7889);
or U9892 (N_9892,N_7361,N_7903);
and U9893 (N_9893,N_7734,N_6444);
or U9894 (N_9894,N_7393,N_7721);
nor U9895 (N_9895,N_7818,N_6059);
and U9896 (N_9896,N_6896,N_7689);
nor U9897 (N_9897,N_7921,N_6555);
nand U9898 (N_9898,N_7151,N_7326);
nor U9899 (N_9899,N_6587,N_7920);
nand U9900 (N_9900,N_6908,N_6073);
and U9901 (N_9901,N_7030,N_7359);
nand U9902 (N_9902,N_7117,N_6324);
and U9903 (N_9903,N_6948,N_6209);
xnor U9904 (N_9904,N_7064,N_7022);
and U9905 (N_9905,N_6184,N_6670);
nor U9906 (N_9906,N_6649,N_6111);
nand U9907 (N_9907,N_6633,N_6972);
or U9908 (N_9908,N_6754,N_7917);
and U9909 (N_9909,N_6103,N_6340);
nand U9910 (N_9910,N_6403,N_6927);
or U9911 (N_9911,N_7224,N_6484);
and U9912 (N_9912,N_7088,N_7954);
nand U9913 (N_9913,N_6927,N_7692);
nor U9914 (N_9914,N_7613,N_6211);
nor U9915 (N_9915,N_7801,N_6622);
nor U9916 (N_9916,N_6055,N_7394);
nor U9917 (N_9917,N_6314,N_7682);
and U9918 (N_9918,N_6405,N_6676);
nand U9919 (N_9919,N_6217,N_6472);
nand U9920 (N_9920,N_7985,N_7766);
nand U9921 (N_9921,N_7386,N_7095);
nand U9922 (N_9922,N_7737,N_6966);
nand U9923 (N_9923,N_7262,N_7930);
nor U9924 (N_9924,N_7103,N_6419);
or U9925 (N_9925,N_7214,N_7058);
or U9926 (N_9926,N_7131,N_6710);
nor U9927 (N_9927,N_7258,N_6831);
or U9928 (N_9928,N_6053,N_6067);
nor U9929 (N_9929,N_7690,N_6644);
nand U9930 (N_9930,N_6701,N_7578);
nand U9931 (N_9931,N_7724,N_6883);
and U9932 (N_9932,N_6877,N_7250);
and U9933 (N_9933,N_6875,N_6016);
and U9934 (N_9934,N_6271,N_7329);
nand U9935 (N_9935,N_6900,N_7137);
or U9936 (N_9936,N_7927,N_6059);
nand U9937 (N_9937,N_6846,N_6972);
or U9938 (N_9938,N_6778,N_7730);
nand U9939 (N_9939,N_7520,N_7166);
or U9940 (N_9940,N_7357,N_7130);
or U9941 (N_9941,N_7911,N_7345);
or U9942 (N_9942,N_7170,N_6125);
and U9943 (N_9943,N_7486,N_6666);
xnor U9944 (N_9944,N_6086,N_7570);
and U9945 (N_9945,N_7480,N_7741);
and U9946 (N_9946,N_7855,N_7641);
or U9947 (N_9947,N_6511,N_6679);
nor U9948 (N_9948,N_7132,N_7880);
nor U9949 (N_9949,N_6114,N_7477);
nor U9950 (N_9950,N_7023,N_7803);
and U9951 (N_9951,N_7581,N_6494);
nand U9952 (N_9952,N_6433,N_7734);
or U9953 (N_9953,N_6602,N_6497);
nor U9954 (N_9954,N_7449,N_6040);
nor U9955 (N_9955,N_6127,N_6787);
nand U9956 (N_9956,N_7781,N_6558);
nand U9957 (N_9957,N_6648,N_6032);
nor U9958 (N_9958,N_7928,N_7006);
nor U9959 (N_9959,N_7040,N_7536);
and U9960 (N_9960,N_6157,N_6609);
or U9961 (N_9961,N_7001,N_7107);
nor U9962 (N_9962,N_7205,N_7269);
or U9963 (N_9963,N_7363,N_7897);
nand U9964 (N_9964,N_6912,N_6695);
and U9965 (N_9965,N_6378,N_6957);
and U9966 (N_9966,N_6135,N_7835);
or U9967 (N_9967,N_6558,N_7288);
or U9968 (N_9968,N_6183,N_7239);
nand U9969 (N_9969,N_7521,N_7171);
xor U9970 (N_9970,N_7096,N_7459);
nor U9971 (N_9971,N_6999,N_7287);
or U9972 (N_9972,N_7589,N_6256);
and U9973 (N_9973,N_6121,N_7692);
nor U9974 (N_9974,N_6757,N_7226);
nand U9975 (N_9975,N_7046,N_6544);
or U9976 (N_9976,N_7783,N_7697);
nor U9977 (N_9977,N_7528,N_7120);
nor U9978 (N_9978,N_7667,N_6746);
nand U9979 (N_9979,N_6809,N_6214);
or U9980 (N_9980,N_7888,N_6260);
nand U9981 (N_9981,N_6305,N_7812);
nand U9982 (N_9982,N_6983,N_6505);
or U9983 (N_9983,N_7029,N_6056);
nor U9984 (N_9984,N_7029,N_7841);
and U9985 (N_9985,N_6614,N_6351);
or U9986 (N_9986,N_7782,N_6639);
and U9987 (N_9987,N_6068,N_6434);
nor U9988 (N_9988,N_6447,N_7649);
nor U9989 (N_9989,N_6462,N_6324);
nand U9990 (N_9990,N_6645,N_6289);
or U9991 (N_9991,N_6483,N_6523);
and U9992 (N_9992,N_6009,N_7621);
or U9993 (N_9993,N_7248,N_6375);
and U9994 (N_9994,N_7604,N_7129);
nor U9995 (N_9995,N_7839,N_6721);
or U9996 (N_9996,N_6848,N_6422);
and U9997 (N_9997,N_7326,N_7139);
nand U9998 (N_9998,N_7730,N_7976);
and U9999 (N_9999,N_6681,N_6615);
nand UO_0 (O_0,N_9894,N_8776);
and UO_1 (O_1,N_8618,N_8649);
nand UO_2 (O_2,N_9933,N_8648);
and UO_3 (O_3,N_9799,N_9822);
nand UO_4 (O_4,N_9541,N_9774);
and UO_5 (O_5,N_9821,N_8152);
nor UO_6 (O_6,N_9651,N_8303);
and UO_7 (O_7,N_8269,N_8889);
or UO_8 (O_8,N_8996,N_9740);
nor UO_9 (O_9,N_8815,N_9996);
and UO_10 (O_10,N_9805,N_8172);
nor UO_11 (O_11,N_8698,N_8426);
nand UO_12 (O_12,N_9167,N_9274);
or UO_13 (O_13,N_9516,N_8007);
nor UO_14 (O_14,N_8543,N_9661);
or UO_15 (O_15,N_8507,N_8693);
nor UO_16 (O_16,N_9265,N_8765);
and UO_17 (O_17,N_8188,N_8340);
nand UO_18 (O_18,N_9536,N_9751);
and UO_19 (O_19,N_8042,N_9948);
or UO_20 (O_20,N_8612,N_8357);
and UO_21 (O_21,N_8533,N_9110);
or UO_22 (O_22,N_9625,N_9643);
nor UO_23 (O_23,N_9079,N_8165);
nor UO_24 (O_24,N_8561,N_9750);
and UO_25 (O_25,N_8314,N_8917);
nand UO_26 (O_26,N_9723,N_8305);
or UO_27 (O_27,N_8457,N_8619);
xor UO_28 (O_28,N_9061,N_8548);
and UO_29 (O_29,N_9424,N_8247);
or UO_30 (O_30,N_9904,N_8713);
nor UO_31 (O_31,N_9322,N_8341);
and UO_32 (O_32,N_9957,N_9486);
nand UO_33 (O_33,N_9871,N_8704);
or UO_34 (O_34,N_8692,N_8335);
and UO_35 (O_35,N_9150,N_8096);
and UO_36 (O_36,N_9888,N_8892);
and UO_37 (O_37,N_8034,N_9186);
nor UO_38 (O_38,N_8937,N_8216);
or UO_39 (O_39,N_9685,N_9830);
or UO_40 (O_40,N_9573,N_8367);
nand UO_41 (O_41,N_9914,N_8856);
xnor UO_42 (O_42,N_8381,N_9719);
xor UO_43 (O_43,N_9294,N_8928);
nor UO_44 (O_44,N_9381,N_8793);
nor UO_45 (O_45,N_9713,N_8631);
xnor UO_46 (O_46,N_8031,N_8998);
nand UO_47 (O_47,N_8444,N_8415);
or UO_48 (O_48,N_9977,N_9236);
or UO_49 (O_49,N_9959,N_8267);
nand UO_50 (O_50,N_8270,N_8600);
nand UO_51 (O_51,N_9578,N_8223);
nor UO_52 (O_52,N_9058,N_8769);
and UO_53 (O_53,N_8865,N_8604);
nand UO_54 (O_54,N_9641,N_8321);
or UO_55 (O_55,N_9581,N_9758);
nor UO_56 (O_56,N_9208,N_9846);
nand UO_57 (O_57,N_9817,N_8439);
and UO_58 (O_58,N_9820,N_9562);
and UO_59 (O_59,N_9847,N_9320);
nor UO_60 (O_60,N_8682,N_9158);
and UO_61 (O_61,N_9816,N_8753);
and UO_62 (O_62,N_8014,N_9577);
or UO_63 (O_63,N_8201,N_9863);
nor UO_64 (O_64,N_8602,N_9038);
or UO_65 (O_65,N_9304,N_8762);
nor UO_66 (O_66,N_9440,N_9442);
or UO_67 (O_67,N_8894,N_8897);
or UO_68 (O_68,N_8553,N_9289);
nor UO_69 (O_69,N_9133,N_9203);
nand UO_70 (O_70,N_9323,N_8028);
or UO_71 (O_71,N_8639,N_8151);
nor UO_72 (O_72,N_8912,N_8187);
nand UO_73 (O_73,N_8530,N_8154);
nand UO_74 (O_74,N_9912,N_9645);
or UO_75 (O_75,N_8491,N_8578);
and UO_76 (O_76,N_8641,N_8024);
nor UO_77 (O_77,N_9161,N_9270);
or UO_78 (O_78,N_8922,N_9238);
nor UO_79 (O_79,N_8646,N_9334);
nor UO_80 (O_80,N_9211,N_8809);
nor UO_81 (O_81,N_9946,N_9048);
or UO_82 (O_82,N_8326,N_9831);
xnor UO_83 (O_83,N_8951,N_9919);
nor UO_84 (O_84,N_8363,N_9547);
nand UO_85 (O_85,N_9934,N_9902);
nor UO_86 (O_86,N_9614,N_8003);
nand UO_87 (O_87,N_9200,N_8637);
nor UO_88 (O_88,N_9829,N_8675);
nand UO_89 (O_89,N_9098,N_8816);
or UO_90 (O_90,N_8958,N_8421);
or UO_91 (O_91,N_9170,N_8512);
or UO_92 (O_92,N_8244,N_8697);
nor UO_93 (O_93,N_9962,N_8760);
nor UO_94 (O_94,N_9070,N_9439);
nand UO_95 (O_95,N_9164,N_9035);
or UO_96 (O_96,N_9371,N_9088);
nand UO_97 (O_97,N_9319,N_8744);
or UO_98 (O_98,N_8943,N_8521);
or UO_99 (O_99,N_8198,N_8925);
or UO_100 (O_100,N_9195,N_9796);
or UO_101 (O_101,N_9353,N_8538);
or UO_102 (O_102,N_8685,N_9143);
nand UO_103 (O_103,N_8098,N_9107);
or UO_104 (O_104,N_8589,N_8354);
nand UO_105 (O_105,N_8857,N_9858);
and UO_106 (O_106,N_8866,N_9668);
or UO_107 (O_107,N_8399,N_8060);
nand UO_108 (O_108,N_8080,N_8268);
or UO_109 (O_109,N_9767,N_9501);
nor UO_110 (O_110,N_8683,N_8821);
and UO_111 (O_111,N_8924,N_9564);
or UO_112 (O_112,N_9795,N_8283);
or UO_113 (O_113,N_8715,N_9823);
and UO_114 (O_114,N_9332,N_9369);
nand UO_115 (O_115,N_9819,N_8380);
and UO_116 (O_116,N_9108,N_9835);
and UO_117 (O_117,N_9591,N_8699);
and UO_118 (O_118,N_9254,N_9706);
nor UO_119 (O_119,N_9695,N_8555);
nand UO_120 (O_120,N_9991,N_9433);
nand UO_121 (O_121,N_9908,N_9775);
and UO_122 (O_122,N_9394,N_9772);
or UO_123 (O_123,N_8624,N_8272);
nand UO_124 (O_124,N_8804,N_9530);
xor UO_125 (O_125,N_8869,N_9684);
or UO_126 (O_126,N_9647,N_8626);
nand UO_127 (O_127,N_8838,N_8174);
xnor UO_128 (O_128,N_9426,N_9415);
nand UO_129 (O_129,N_9184,N_9072);
and UO_130 (O_130,N_8472,N_9509);
nand UO_131 (O_131,N_8502,N_8064);
nor UO_132 (O_132,N_8938,N_9802);
or UO_133 (O_133,N_9295,N_9216);
nor UO_134 (O_134,N_9698,N_8617);
or UO_135 (O_135,N_8927,N_8807);
nand UO_136 (O_136,N_9901,N_8166);
nand UO_137 (O_137,N_8633,N_8228);
and UO_138 (O_138,N_8205,N_9284);
or UO_139 (O_139,N_9328,N_9436);
nand UO_140 (O_140,N_9636,N_8373);
nand UO_141 (O_141,N_9836,N_9720);
xor UO_142 (O_142,N_8070,N_9592);
or UO_143 (O_143,N_8375,N_8842);
nand UO_144 (O_144,N_8733,N_8241);
nor UO_145 (O_145,N_9642,N_9696);
or UO_146 (O_146,N_9811,N_8132);
and UO_147 (O_147,N_9518,N_8263);
and UO_148 (O_148,N_8450,N_8297);
nand UO_149 (O_149,N_9496,N_8689);
and UO_150 (O_150,N_9413,N_8351);
and UO_151 (O_151,N_8078,N_8386);
nor UO_152 (O_152,N_9543,N_9384);
or UO_153 (O_153,N_8443,N_8501);
nor UO_154 (O_154,N_8334,N_8904);
or UO_155 (O_155,N_9618,N_9937);
nand UO_156 (O_156,N_9055,N_9920);
or UO_157 (O_157,N_8480,N_8588);
or UO_158 (O_158,N_9165,N_9903);
or UO_159 (O_159,N_9271,N_9327);
nand UO_160 (O_160,N_9884,N_8503);
or UO_161 (O_161,N_9140,N_8182);
and UO_162 (O_162,N_9728,N_8707);
nor UO_163 (O_163,N_8248,N_8150);
or UO_164 (O_164,N_8886,N_8500);
or UO_165 (O_165,N_8611,N_9585);
nor UO_166 (O_166,N_8966,N_9374);
nor UO_167 (O_167,N_8104,N_9561);
nand UO_168 (O_168,N_9080,N_8318);
or UO_169 (O_169,N_9213,N_8515);
and UO_170 (O_170,N_8420,N_8668);
nor UO_171 (O_171,N_9860,N_9664);
nor UO_172 (O_172,N_8650,N_9659);
and UO_173 (O_173,N_8710,N_9030);
or UO_174 (O_174,N_8803,N_9454);
nand UO_175 (O_175,N_9141,N_8220);
and UO_176 (O_176,N_9168,N_8986);
nor UO_177 (O_177,N_8881,N_8116);
nor UO_178 (O_178,N_9670,N_9762);
or UO_179 (O_179,N_9301,N_9722);
nor UO_180 (O_180,N_9872,N_8948);
or UO_181 (O_181,N_8999,N_8526);
or UO_182 (O_182,N_8284,N_8011);
nand UO_183 (O_183,N_9050,N_8863);
xnor UO_184 (O_184,N_9565,N_9191);
nand UO_185 (O_185,N_9183,N_9125);
nand UO_186 (O_186,N_8254,N_8061);
nor UO_187 (O_187,N_8071,N_8581);
and UO_188 (O_188,N_9973,N_8738);
nor UO_189 (O_189,N_8979,N_9124);
nand UO_190 (O_190,N_9623,N_8067);
or UO_191 (O_191,N_9631,N_8723);
or UO_192 (O_192,N_9905,N_9113);
nor UO_193 (O_193,N_8901,N_8135);
xor UO_194 (O_194,N_8178,N_9635);
and UO_195 (O_195,N_8687,N_9155);
and UO_196 (O_196,N_8926,N_8320);
or UO_197 (O_197,N_9842,N_9026);
nor UO_198 (O_198,N_9593,N_8642);
nor UO_199 (O_199,N_8125,N_8885);
and UO_200 (O_200,N_8158,N_8211);
or UO_201 (O_201,N_8627,N_9961);
or UO_202 (O_202,N_9528,N_9730);
and UO_203 (O_203,N_8890,N_9727);
and UO_204 (O_204,N_9324,N_8566);
and UO_205 (O_205,N_8829,N_8414);
nor UO_206 (O_206,N_9103,N_9041);
nand UO_207 (O_207,N_8868,N_8562);
or UO_208 (O_208,N_8221,N_9489);
and UO_209 (O_209,N_8694,N_9257);
nor UO_210 (O_210,N_9575,N_8279);
nor UO_211 (O_211,N_8781,N_8814);
and UO_212 (O_212,N_8371,N_8280);
nand UO_213 (O_213,N_9985,N_9674);
nand UO_214 (O_214,N_9339,N_8576);
nand UO_215 (O_215,N_9313,N_8123);
nor UO_216 (O_216,N_8325,N_8477);
xor UO_217 (O_217,N_8240,N_8957);
nor UO_218 (O_218,N_8103,N_8458);
and UO_219 (O_219,N_8993,N_9465);
nand UO_220 (O_220,N_9747,N_8843);
and UO_221 (O_221,N_8117,N_8140);
nand UO_222 (O_222,N_8249,N_8790);
and UO_223 (O_223,N_9280,N_9428);
nor UO_224 (O_224,N_9016,N_9028);
nand UO_225 (O_225,N_9326,N_8218);
nor UO_226 (O_226,N_8967,N_8105);
or UO_227 (O_227,N_8556,N_9074);
nand UO_228 (O_228,N_9132,N_8171);
or UO_229 (O_229,N_9084,N_9924);
nor UO_230 (O_230,N_8913,N_8573);
nor UO_231 (O_231,N_9637,N_8233);
nor UO_232 (O_232,N_8590,N_8980);
nor UO_233 (O_233,N_8134,N_9979);
nor UO_234 (O_234,N_9330,N_9926);
and UO_235 (O_235,N_9307,N_8185);
and UO_236 (O_236,N_8819,N_9288);
nand UO_237 (O_237,N_9956,N_9073);
and UO_238 (O_238,N_8539,N_8408);
and UO_239 (O_239,N_9091,N_8782);
xor UO_240 (O_240,N_9130,N_9671);
or UO_241 (O_241,N_9019,N_8615);
or UO_242 (O_242,N_9492,N_9711);
or UO_243 (O_243,N_8382,N_8264);
nor UO_244 (O_244,N_8720,N_9552);
nand UO_245 (O_245,N_8564,N_9175);
nor UO_246 (O_246,N_9735,N_8518);
and UO_247 (O_247,N_9285,N_8989);
nand UO_248 (O_248,N_9567,N_8250);
nor UO_249 (O_249,N_9794,N_9502);
nand UO_250 (O_250,N_9752,N_9527);
nand UO_251 (O_251,N_8114,N_8106);
or UO_252 (O_252,N_8235,N_9954);
or UO_253 (O_253,N_8126,N_8160);
or UO_254 (O_254,N_9754,N_9586);
and UO_255 (O_255,N_8427,N_9356);
nor UO_256 (O_256,N_9405,N_9114);
nor UO_257 (O_257,N_8965,N_9421);
and UO_258 (O_258,N_8862,N_8570);
nor UO_259 (O_259,N_8919,N_9146);
nor UO_260 (O_260,N_9742,N_9721);
nand UO_261 (O_261,N_9785,N_9615);
and UO_262 (O_262,N_9344,N_8644);
nor UO_263 (O_263,N_9172,N_9495);
and UO_264 (O_264,N_9443,N_8121);
and UO_265 (O_265,N_9169,N_8794);
nand UO_266 (O_266,N_9065,N_9718);
nor UO_267 (O_267,N_9764,N_8497);
and UO_268 (O_268,N_9563,N_8025);
or UO_269 (O_269,N_9475,N_8473);
nor UO_270 (O_270,N_9966,N_9691);
nand UO_271 (O_271,N_9708,N_8832);
or UO_272 (O_272,N_8709,N_8545);
or UO_273 (O_273,N_9382,N_8008);
and UO_274 (O_274,N_8184,N_8137);
nor UO_275 (O_275,N_9112,N_9268);
nand UO_276 (O_276,N_9673,N_9628);
nand UO_277 (O_277,N_8625,N_9755);
or UO_278 (O_278,N_8461,N_9776);
or UO_279 (O_279,N_9990,N_8660);
or UO_280 (O_280,N_8859,N_9494);
or UO_281 (O_281,N_9629,N_9460);
or UO_282 (O_282,N_9089,N_8065);
nor UO_283 (O_283,N_9232,N_9147);
nand UO_284 (O_284,N_9781,N_9570);
or UO_285 (O_285,N_9459,N_9748);
nor UO_286 (O_286,N_8895,N_8860);
or UO_287 (O_287,N_9532,N_8558);
or UO_288 (O_288,N_8026,N_9619);
and UO_289 (O_289,N_9018,N_8778);
or UO_290 (O_290,N_9769,N_8990);
and UO_291 (O_291,N_9438,N_9710);
nor UO_292 (O_292,N_9553,N_9677);
nor UO_293 (O_293,N_9481,N_8976);
nand UO_294 (O_294,N_8879,N_8728);
nand UO_295 (O_295,N_9185,N_8058);
nand UO_296 (O_296,N_8510,N_8206);
nand UO_297 (O_297,N_9159,N_9950);
nor UO_298 (O_298,N_8173,N_8469);
nor UO_299 (O_299,N_9850,N_8679);
nor UO_300 (O_300,N_8099,N_9535);
nor UO_301 (O_301,N_9451,N_8735);
nand UO_302 (O_302,N_8483,N_8867);
nor UO_303 (O_303,N_8676,N_8584);
or UO_304 (O_304,N_9930,N_9972);
or UO_305 (O_305,N_8987,N_9649);
xor UO_306 (O_306,N_8508,N_9005);
or UO_307 (O_307,N_9505,N_9792);
nand UO_308 (O_308,N_9907,N_8056);
nor UO_309 (O_309,N_8253,N_8462);
nand UO_310 (O_310,N_8608,N_9978);
and UO_311 (O_311,N_8434,N_8000);
and UO_312 (O_312,N_9012,N_8470);
and UO_313 (O_313,N_9929,N_8955);
and UO_314 (O_314,N_8690,N_8906);
nor UO_315 (O_315,N_8516,N_8256);
nand UO_316 (O_316,N_8786,N_8830);
and UO_317 (O_317,N_8342,N_8485);
nand UO_318 (O_318,N_8995,N_9834);
or UO_319 (O_319,N_9062,N_8484);
nor UO_320 (O_320,N_8037,N_9539);
or UO_321 (O_321,N_8601,N_9782);
nand UO_322 (O_322,N_9109,N_9529);
nand UO_323 (O_323,N_8203,N_8899);
nand UO_324 (O_324,N_9941,N_8175);
and UO_325 (O_325,N_9408,N_9044);
nor UO_326 (O_326,N_9498,N_8294);
nor UO_327 (O_327,N_8826,N_9572);
or UO_328 (O_328,N_8953,N_8616);
nand UO_329 (O_329,N_9968,N_9855);
nor UO_330 (O_330,N_9947,N_9241);
and UO_331 (O_331,N_8847,N_9497);
and UO_332 (O_332,N_9360,N_9364);
nor UO_333 (O_333,N_9149,N_9583);
nor UO_334 (O_334,N_9514,N_8835);
nand UO_335 (O_335,N_9699,N_8308);
nand UO_336 (O_336,N_9264,N_9815);
and UO_337 (O_337,N_8640,N_8146);
and UO_338 (O_338,N_8232,N_8529);
or UO_339 (O_339,N_8419,N_9456);
or UO_340 (O_340,N_8143,N_9244);
or UO_341 (O_341,N_9476,N_8429);
nor UO_342 (O_342,N_8936,N_9461);
nor UO_343 (O_343,N_9190,N_9839);
nand UO_344 (O_344,N_8094,N_8898);
and UO_345 (O_345,N_8127,N_9546);
or UO_346 (O_346,N_8355,N_9129);
nor UO_347 (O_347,N_9471,N_8811);
xor UO_348 (O_348,N_8586,N_9305);
and UO_349 (O_349,N_8422,N_9283);
nor UO_350 (O_350,N_9602,N_8124);
nor UO_351 (O_351,N_8563,N_9142);
or UO_352 (O_352,N_8721,N_9337);
nor UO_353 (O_353,N_9542,N_9757);
or UO_354 (O_354,N_8651,N_8577);
nor UO_355 (O_355,N_8849,N_8102);
and UO_356 (O_356,N_9824,N_9134);
nor UO_357 (O_357,N_8672,N_8213);
nand UO_358 (O_358,N_9624,N_9916);
and UO_359 (O_359,N_9152,N_8686);
and UO_360 (O_360,N_9126,N_9228);
and UO_361 (O_361,N_9523,N_9653);
or UO_362 (O_362,N_8701,N_9444);
or UO_363 (O_363,N_9432,N_8932);
and UO_364 (O_364,N_8463,N_9911);
xnor UO_365 (O_365,N_9027,N_8571);
nor UO_366 (O_366,N_8086,N_8169);
xor UO_367 (O_367,N_9549,N_8368);
or UO_368 (O_368,N_9092,N_8441);
nand UO_369 (O_369,N_9975,N_9231);
or UO_370 (O_370,N_9144,N_8416);
nor UO_371 (O_371,N_8652,N_9100);
nor UO_372 (O_372,N_8306,N_8891);
nand UO_373 (O_373,N_9256,N_9226);
nor UO_374 (O_374,N_9046,N_8915);
nand UO_375 (O_375,N_8729,N_8082);
or UO_376 (O_376,N_9045,N_9998);
or UO_377 (O_377,N_8409,N_8930);
nor UO_378 (O_378,N_9809,N_8093);
or UO_379 (O_379,N_9511,N_8837);
or UO_380 (O_380,N_9212,N_8278);
nand UO_381 (O_381,N_8517,N_8179);
and UO_382 (O_382,N_9943,N_8896);
and UO_383 (O_383,N_8196,N_9652);
nand UO_384 (O_384,N_9009,N_8754);
and UO_385 (O_385,N_8120,N_8433);
nand UO_386 (O_386,N_8550,N_9876);
and UO_387 (O_387,N_9004,N_8275);
or UO_388 (O_388,N_9874,N_9841);
or UO_389 (O_389,N_8110,N_8850);
and UO_390 (O_390,N_9955,N_9679);
or UO_391 (O_391,N_9886,N_9189);
or UO_392 (O_392,N_9632,N_9810);
and UO_393 (O_393,N_8771,N_8909);
xor UO_394 (O_394,N_8488,N_9136);
or UO_395 (O_395,N_8168,N_8224);
and UO_396 (O_396,N_9033,N_9725);
and UO_397 (O_397,N_8313,N_8873);
and UO_398 (O_398,N_8317,N_9665);
nor UO_399 (O_399,N_8864,N_8593);
nand UO_400 (O_400,N_9617,N_8369);
nand UO_401 (O_401,N_8506,N_9524);
nand UO_402 (O_402,N_9621,N_8229);
or UO_403 (O_403,N_9176,N_8300);
or UO_404 (O_404,N_8487,N_9362);
nor UO_405 (O_405,N_9500,N_8509);
nand UO_406 (O_406,N_9951,N_9389);
and UO_407 (O_407,N_9927,N_8594);
nand UO_408 (O_408,N_9474,N_9559);
nor UO_409 (O_409,N_8663,N_8455);
or UO_410 (O_410,N_9391,N_9892);
or UO_411 (O_411,N_8519,N_8131);
nand UO_412 (O_412,N_8460,N_9897);
nor UO_413 (O_413,N_9517,N_9249);
nand UO_414 (O_414,N_9419,N_9230);
nor UO_415 (O_415,N_8645,N_8107);
and UO_416 (O_416,N_8424,N_8076);
or UO_417 (O_417,N_8875,N_8960);
or UO_418 (O_418,N_8481,N_8255);
nor UO_419 (O_419,N_8410,N_8083);
or UO_420 (O_420,N_8069,N_8021);
nor UO_421 (O_421,N_8020,N_9574);
nand UO_422 (O_422,N_9967,N_8315);
nand UO_423 (O_423,N_9272,N_9803);
nand UO_424 (O_424,N_9866,N_8671);
nor UO_425 (O_425,N_8430,N_8452);
nand UO_426 (O_426,N_8199,N_9101);
nand UO_427 (O_427,N_8716,N_8144);
and UO_428 (O_428,N_9569,N_8724);
nor UO_429 (O_429,N_9939,N_9379);
and UO_430 (O_430,N_9064,N_9844);
xnor UO_431 (O_431,N_9262,N_8226);
nand UO_432 (O_432,N_8607,N_9983);
or UO_433 (O_433,N_9034,N_8498);
nand UO_434 (O_434,N_9837,N_8741);
nand UO_435 (O_435,N_8392,N_9784);
xnor UO_436 (O_436,N_9398,N_8973);
and UO_437 (O_437,N_9281,N_8541);
nand UO_438 (O_438,N_8737,N_8394);
or UO_439 (O_439,N_8339,N_9499);
nor UO_440 (O_440,N_8494,N_9890);
and UO_441 (O_441,N_8183,N_9047);
and UO_442 (O_442,N_8393,N_9355);
nand UO_443 (O_443,N_8242,N_8582);
xor UO_444 (O_444,N_8634,N_9995);
nor UO_445 (O_445,N_9644,N_9007);
nor UO_446 (O_446,N_8757,N_8459);
nand UO_447 (O_447,N_8149,N_8779);
nor UO_448 (O_448,N_9013,N_9345);
nor UO_449 (O_449,N_8290,N_8527);
or UO_450 (O_450,N_9945,N_9906);
nor UO_451 (O_451,N_8759,N_9702);
and UO_452 (O_452,N_9411,N_9425);
and UO_453 (O_453,N_8537,N_8387);
or UO_454 (O_454,N_8052,N_9198);
or UO_455 (O_455,N_9331,N_9786);
and UO_456 (O_456,N_8916,N_8714);
nand UO_457 (O_457,N_8360,N_8330);
or UO_458 (O_458,N_9812,N_8664);
and UO_459 (O_459,N_8877,N_9071);
and UO_460 (O_460,N_9464,N_8920);
or UO_461 (O_461,N_8599,N_9446);
nand UO_462 (O_462,N_8111,N_9448);
nor UO_463 (O_463,N_8230,N_8364);
nor UO_464 (O_464,N_8446,N_8975);
or UO_465 (O_465,N_8490,N_8261);
nor UO_466 (O_466,N_9825,N_9707);
and UO_467 (O_467,N_9397,N_9031);
nor UO_468 (O_468,N_9215,N_8192);
nor UO_469 (O_469,N_9878,N_8827);
and UO_470 (O_470,N_9145,N_8170);
or UO_471 (O_471,N_9131,N_9544);
nand UO_472 (O_472,N_8595,N_9219);
nand UO_473 (O_473,N_9859,N_8972);
and UO_474 (O_474,N_8274,N_8788);
and UO_475 (O_475,N_9291,N_8115);
nand UO_476 (O_476,N_8479,N_8992);
nand UO_477 (O_477,N_8939,N_8888);
nand UO_478 (O_478,N_8981,N_8013);
nor UO_479 (O_479,N_9705,N_8567);
nor UO_480 (O_480,N_8468,N_8722);
nand UO_481 (O_481,N_8903,N_9453);
nor UO_482 (O_482,N_9714,N_9588);
nand UO_483 (O_483,N_8177,N_9733);
nor UO_484 (O_484,N_8400,N_9376);
nor UO_485 (O_485,N_9717,N_8820);
nor UO_486 (O_486,N_8756,N_9519);
nor UO_487 (O_487,N_9455,N_9808);
or UO_488 (O_488,N_9278,N_9885);
and UO_489 (O_489,N_9655,N_9377);
or UO_490 (O_490,N_8260,N_9506);
and UO_491 (O_491,N_9049,N_8840);
nor UO_492 (O_492,N_9255,N_8307);
nand UO_493 (O_493,N_9548,N_8823);
nor UO_494 (O_494,N_8622,N_8702);
nand UO_495 (O_495,N_8289,N_8466);
or UO_496 (O_496,N_9056,N_8141);
nand UO_497 (O_497,N_8551,N_8108);
and UO_498 (O_498,N_9227,N_8265);
or UO_499 (O_499,N_9763,N_8963);
or UO_500 (O_500,N_9760,N_9877);
and UO_501 (O_501,N_9650,N_9022);
nand UO_502 (O_502,N_9612,N_8323);
and UO_503 (O_503,N_9917,N_8258);
and UO_504 (O_504,N_9373,N_9944);
or UO_505 (O_505,N_8511,N_8041);
or UO_506 (O_506,N_9490,N_8449);
and UO_507 (O_507,N_8194,N_9918);
nand UO_508 (O_508,N_9037,N_9276);
or UO_509 (O_509,N_9335,N_8825);
nand UO_510 (O_510,N_9843,N_8465);
or UO_511 (O_511,N_9317,N_8101);
nor UO_512 (O_512,N_8332,N_8614);
nand UO_513 (O_513,N_8050,N_9250);
nor UO_514 (O_514,N_9923,N_9534);
nand UO_515 (O_515,N_9738,N_9982);
nor UO_516 (O_516,N_8384,N_8505);
and UO_517 (O_517,N_8969,N_8678);
nor UO_518 (O_518,N_8504,N_9017);
nor UO_519 (O_519,N_9880,N_9387);
nand UO_520 (O_520,N_8876,N_8952);
nand UO_521 (O_521,N_9590,N_9259);
and UO_522 (O_522,N_9512,N_9589);
and UO_523 (O_523,N_9090,N_9818);
nand UO_524 (O_524,N_8406,N_9683);
nand UO_525 (O_525,N_9607,N_8798);
nor UO_526 (O_526,N_8749,N_8040);
nand UO_527 (O_527,N_8090,N_9154);
and UO_528 (O_528,N_8910,N_8942);
and UO_529 (O_529,N_8810,N_8708);
and UO_530 (O_530,N_9309,N_8900);
nand UO_531 (O_531,N_8606,N_9378);
nand UO_532 (O_532,N_8775,N_9687);
or UO_533 (O_533,N_8659,N_9220);
and UO_534 (O_534,N_9953,N_9069);
nand UO_535 (O_535,N_9666,N_9582);
or UO_536 (O_536,N_8596,N_9971);
or UO_537 (O_537,N_8846,N_8680);
and UO_538 (O_538,N_9806,N_9551);
nor UO_539 (O_539,N_8251,N_8425);
or UO_540 (O_540,N_9210,N_8077);
nand UO_541 (O_541,N_8176,N_8657);
nand UO_542 (O_542,N_8880,N_8745);
and UO_543 (O_543,N_8319,N_9620);
or UO_544 (O_544,N_9095,N_8520);
nand UO_545 (O_545,N_9746,N_9392);
nand UO_546 (O_546,N_9025,N_8883);
or UO_547 (O_547,N_9225,N_9214);
nor UO_548 (O_548,N_9452,N_9217);
nor UO_549 (O_549,N_9840,N_9105);
xnor UO_550 (O_550,N_8136,N_9640);
or UO_551 (O_551,N_9002,N_8057);
nor UO_552 (O_552,N_8968,N_9416);
and UO_553 (O_553,N_9694,N_9568);
and UO_554 (O_554,N_9609,N_9522);
nand UO_555 (O_555,N_9209,N_9560);
and UO_556 (O_556,N_9300,N_8579);
nand UO_557 (O_557,N_8210,N_9052);
or UO_558 (O_558,N_9429,N_9119);
xnor UO_559 (O_559,N_8605,N_8238);
nor UO_560 (O_560,N_9660,N_9692);
nand UO_561 (O_561,N_8217,N_8163);
nor UO_562 (O_562,N_8066,N_9404);
xnor UO_563 (O_563,N_8806,N_8861);
or UO_564 (O_564,N_8941,N_8298);
nor UO_565 (O_565,N_9765,N_9610);
nor UO_566 (O_566,N_9006,N_9417);
and UO_567 (O_567,N_8544,N_9368);
or UO_568 (O_568,N_8271,N_9409);
nand UO_569 (O_569,N_8674,N_8751);
and UO_570 (O_570,N_8746,N_8286);
nand UO_571 (O_571,N_8528,N_9538);
or UO_572 (O_572,N_8492,N_9845);
nor UO_573 (O_573,N_8147,N_9097);
and UO_574 (O_574,N_9580,N_9743);
nand UO_575 (O_575,N_9960,N_9887);
and UO_576 (O_576,N_8081,N_9681);
and UO_577 (O_577,N_8747,N_9293);
and UO_578 (O_578,N_8331,N_9078);
nand UO_579 (O_579,N_9243,N_9437);
xor UO_580 (O_580,N_8397,N_9251);
nand UO_581 (O_581,N_8774,N_9634);
nand UO_582 (O_582,N_8666,N_9768);
nor UO_583 (O_583,N_8677,N_9359);
nand UO_584 (O_584,N_8391,N_9672);
or UO_585 (O_585,N_9658,N_9087);
or UO_586 (O_586,N_8621,N_8288);
nand UO_587 (O_587,N_9187,N_9701);
nor UO_588 (O_588,N_9478,N_9011);
or UO_589 (O_589,N_9601,N_9341);
or UO_590 (O_590,N_8726,N_9407);
nand UO_591 (O_591,N_8474,N_9800);
and UO_592 (O_592,N_9479,N_8456);
or UO_593 (O_593,N_9989,N_9282);
nor UO_594 (O_594,N_8112,N_9594);
nand UO_595 (O_595,N_8575,N_9510);
or UO_596 (O_596,N_9430,N_9032);
nand UO_597 (O_597,N_9788,N_8944);
and UO_598 (O_598,N_9992,N_9993);
nand UO_599 (O_599,N_8389,N_8353);
or UO_600 (O_600,N_8227,N_9662);
nand UO_601 (O_601,N_9739,N_9279);
and UO_602 (O_602,N_8155,N_9173);
nor UO_603 (O_603,N_9826,N_8428);
nor UO_604 (O_604,N_8792,N_9246);
nor UO_605 (O_605,N_8475,N_9412);
and UO_606 (O_606,N_8546,N_9540);
nand UO_607 (O_607,N_8662,N_9117);
nor UO_608 (O_608,N_9599,N_8167);
nand UO_609 (O_609,N_8647,N_9302);
nor UO_610 (O_610,N_9576,N_9361);
xor UO_611 (O_611,N_8592,N_9269);
nor UO_612 (O_612,N_8396,N_9414);
or UO_613 (O_613,N_9237,N_8390);
or UO_614 (O_614,N_9472,N_9777);
and UO_615 (O_615,N_9181,N_9224);
and UO_616 (O_616,N_9123,N_9613);
or UO_617 (O_617,N_9059,N_8212);
nand UO_618 (O_618,N_8717,N_8739);
nand UO_619 (O_619,N_9949,N_9352);
xor UO_620 (O_620,N_9121,N_8994);
nor UO_621 (O_621,N_8361,N_8598);
and UO_622 (O_622,N_9138,N_9441);
nor UO_623 (O_623,N_8379,N_9557);
or UO_624 (O_624,N_8328,N_8407);
and UO_625 (O_625,N_8044,N_9148);
or UO_626 (O_626,N_9520,N_8348);
or UO_627 (O_627,N_8934,N_9605);
or UO_628 (O_628,N_9616,N_9988);
or UO_629 (O_629,N_8853,N_9969);
and UO_630 (O_630,N_9235,N_8336);
nor UO_631 (O_631,N_8301,N_9375);
nand UO_632 (O_632,N_8752,N_9160);
nor UO_633 (O_633,N_8623,N_8552);
or UO_634 (O_634,N_8302,N_8736);
nor UO_635 (O_635,N_8761,N_9744);
and UO_636 (O_636,N_9366,N_8365);
nor UO_637 (O_637,N_8947,N_8281);
and UO_638 (O_638,N_8696,N_9724);
and UO_639 (O_639,N_8358,N_8467);
nor UO_640 (O_640,N_8985,N_9234);
nand UO_641 (O_641,N_9287,N_9940);
or UO_642 (O_642,N_9638,N_9932);
nand UO_643 (O_643,N_8376,N_8667);
or UO_644 (O_644,N_8542,N_8291);
nor UO_645 (O_645,N_8486,N_9895);
nor UO_646 (O_646,N_9218,N_8092);
or UO_647 (O_647,N_9253,N_8959);
and UO_648 (O_648,N_9606,N_8016);
nor UO_649 (O_649,N_9370,N_8565);
and UO_650 (O_650,N_8587,N_9804);
nand UO_651 (O_651,N_8695,N_8385);
and UO_652 (O_652,N_8964,N_8961);
nor UO_653 (O_653,N_9507,N_9057);
or UO_654 (O_654,N_9686,N_9054);
or UO_655 (O_655,N_9179,N_9199);
xnor UO_656 (O_656,N_8748,N_9365);
and UO_657 (O_657,N_8048,N_9690);
nand UO_658 (O_658,N_8673,N_8918);
nand UO_659 (O_659,N_9856,N_8493);
nand UO_660 (O_660,N_8554,N_9965);
or UO_661 (O_661,N_8157,N_9521);
or UO_662 (O_662,N_8654,N_9697);
nor UO_663 (O_663,N_8161,N_8204);
and UO_664 (O_664,N_8597,N_9075);
or UO_665 (O_665,N_9192,N_9303);
or UO_666 (O_666,N_9931,N_8130);
nor UO_667 (O_667,N_8656,N_8113);
or UO_668 (O_668,N_9388,N_8312);
nor UO_669 (O_669,N_9689,N_8091);
nor UO_670 (O_670,N_9166,N_8523);
and UO_671 (O_671,N_9654,N_9870);
nor UO_672 (O_672,N_8079,N_8085);
and UO_673 (O_673,N_9597,N_9700);
and UO_674 (O_674,N_8983,N_8404);
nor UO_675 (O_675,N_9290,N_9503);
and UO_676 (O_676,N_8068,N_9139);
and UO_677 (O_677,N_9537,N_9063);
or UO_678 (O_678,N_8725,N_9556);
or UO_679 (O_679,N_9174,N_9096);
or UO_680 (O_680,N_8214,N_8374);
nor UO_681 (O_681,N_9128,N_9458);
nand UO_682 (O_682,N_9766,N_9403);
nor UO_683 (O_683,N_8195,N_9197);
or UO_684 (O_684,N_8852,N_8276);
or UO_685 (O_685,N_9611,N_8496);
or UO_686 (O_686,N_9163,N_9367);
or UO_687 (O_687,N_8902,N_9584);
and UO_688 (O_688,N_9603,N_8190);
nor UO_689 (O_689,N_8764,N_9678);
nor UO_690 (O_690,N_8785,N_8036);
and UO_691 (O_691,N_8087,N_8997);
or UO_692 (O_692,N_9067,N_8700);
nor UO_693 (O_693,N_9889,N_8349);
or UO_694 (O_694,N_8128,N_9449);
nand UO_695 (O_695,N_9402,N_9891);
nand UO_696 (O_696,N_8129,N_9311);
and UO_697 (O_697,N_8824,N_9608);
or UO_698 (O_698,N_9463,N_9749);
nor UO_699 (O_699,N_8186,N_8447);
and UO_700 (O_700,N_9771,N_8841);
and UO_701 (O_701,N_9773,N_8072);
nor UO_702 (O_702,N_9162,N_9122);
or UO_703 (O_703,N_8295,N_8059);
nor UO_704 (O_704,N_9480,N_9182);
nor UO_705 (O_705,N_8164,N_9204);
or UO_706 (O_706,N_8732,N_9976);
or UO_707 (O_707,N_8665,N_8984);
nand UO_708 (O_708,N_9693,N_9477);
or UO_709 (O_709,N_9036,N_8200);
and UO_710 (O_710,N_9864,N_9928);
and UO_711 (O_711,N_8039,N_8954);
nand UO_712 (O_712,N_8783,N_8266);
xnor UO_713 (O_713,N_9111,N_8495);
nor UO_714 (O_714,N_8005,N_9223);
nor UO_715 (O_715,N_9066,N_8145);
or UO_716 (O_716,N_9709,N_8222);
or UO_717 (O_717,N_8243,N_9469);
and UO_718 (O_718,N_9487,N_9318);
and UO_719 (O_719,N_9896,N_9526);
nand UO_720 (O_720,N_8403,N_9447);
and UO_721 (O_721,N_9868,N_9260);
or UO_722 (O_722,N_9462,N_9883);
nor UO_723 (O_723,N_8629,N_9086);
and UO_724 (O_724,N_8844,N_8033);
nor UO_725 (O_725,N_9400,N_8310);
and UO_726 (O_726,N_8591,N_9734);
or UO_727 (O_727,N_9997,N_8032);
or UO_728 (O_728,N_9431,N_9485);
and UO_729 (O_729,N_9233,N_8632);
nor UO_730 (O_730,N_9239,N_9240);
nor UO_731 (O_731,N_8089,N_8019);
xnor UO_732 (O_732,N_9936,N_8580);
nor UO_733 (O_733,N_9024,N_9656);
nand UO_734 (O_734,N_8789,N_8181);
nor UO_735 (O_735,N_8202,N_9915);
nand UO_736 (O_736,N_8858,N_8755);
nor UO_737 (O_737,N_8043,N_8451);
or UO_738 (O_738,N_8345,N_9626);
nor UO_739 (O_739,N_9342,N_8719);
nor UO_740 (O_740,N_9395,N_8431);
or UO_741 (O_741,N_9221,N_8585);
nor UO_742 (O_742,N_8299,N_8388);
nand UO_743 (O_743,N_8002,N_9994);
and UO_744 (O_744,N_8740,N_9491);
and UO_745 (O_745,N_9467,N_9296);
and UO_746 (O_746,N_9358,N_8854);
or UO_747 (O_747,N_8812,N_8356);
nand UO_748 (O_748,N_8805,N_9306);
and UO_749 (O_749,N_8661,N_8855);
or UO_750 (O_750,N_9630,N_8075);
or UO_751 (O_751,N_8872,N_8568);
or UO_752 (O_752,N_9504,N_8362);
or UO_753 (O_753,N_9196,N_9222);
or UO_754 (O_754,N_8418,N_9704);
nand UO_755 (O_755,N_8442,N_9881);
nand UO_756 (O_756,N_8800,N_8991);
and UO_757 (O_757,N_8791,N_9321);
and UO_758 (O_758,N_8027,N_9854);
nor UO_759 (O_759,N_9020,N_9814);
or UO_760 (O_760,N_8818,N_8569);
or UO_761 (O_761,N_8239,N_9832);
or UO_762 (O_762,N_9420,N_9869);
and UO_763 (O_763,N_8119,N_9970);
or UO_764 (O_764,N_9484,N_8231);
nor UO_765 (O_765,N_8777,N_9266);
xor UO_766 (O_766,N_8423,N_8197);
and UO_767 (O_767,N_9171,N_9003);
and UO_768 (O_768,N_9383,N_9473);
nor UO_769 (O_769,N_8730,N_9862);
and UO_770 (O_770,N_9267,N_8945);
nand UO_771 (O_771,N_9263,N_9952);
or UO_772 (O_772,N_8574,N_8887);
nor UO_773 (O_773,N_8845,N_8001);
and UO_774 (O_774,N_9115,N_9910);
or UO_775 (O_775,N_9566,N_8929);
and UO_776 (O_776,N_8347,N_8402);
nor UO_777 (O_777,N_8638,N_9913);
or UO_778 (O_778,N_8905,N_9427);
or UO_779 (O_779,N_8706,N_8559);
and UO_780 (O_780,N_9571,N_9639);
or UO_781 (O_781,N_8988,N_9531);
xnor UO_782 (O_782,N_9275,N_8191);
or UO_783 (O_783,N_9043,N_8982);
and UO_784 (O_784,N_8015,N_8338);
nor UO_785 (O_785,N_9828,N_8049);
and UO_786 (O_786,N_8370,N_8549);
nand UO_787 (O_787,N_9791,N_8828);
nor UO_788 (O_788,N_8908,N_8246);
nor UO_789 (O_789,N_9732,N_8046);
nor UO_790 (O_790,N_9082,N_8822);
nor UO_791 (O_791,N_8884,N_8727);
or UO_792 (O_792,N_8282,N_8572);
and UO_793 (O_793,N_9349,N_8398);
nor UO_794 (O_794,N_8907,N_8023);
nor UO_795 (O_795,N_9399,N_8257);
nand UO_796 (O_796,N_8343,N_9648);
nand UO_797 (O_797,N_9093,N_8801);
and UO_798 (O_798,N_8304,N_8287);
nor UO_799 (O_799,N_8237,N_9346);
nor UO_800 (O_800,N_8703,N_9600);
nor UO_801 (O_801,N_8329,N_8534);
or UO_802 (O_802,N_8524,N_8731);
and UO_803 (O_803,N_9422,N_9604);
and UO_804 (O_804,N_8411,N_8471);
nor UO_805 (O_805,N_9981,N_9675);
nor UO_806 (O_806,N_8513,N_9258);
or UO_807 (O_807,N_9627,N_8522);
nand UO_808 (O_808,N_8802,N_8536);
nand UO_809 (O_809,N_9587,N_8609);
nand UO_810 (O_810,N_9867,N_8956);
and UO_811 (O_811,N_8344,N_9329);
nand UO_812 (O_812,N_9261,N_9410);
nand UO_813 (O_813,N_8742,N_8097);
and UO_814 (O_814,N_8547,N_8162);
or UO_815 (O_815,N_8133,N_8405);
nor UO_816 (O_816,N_9396,N_9882);
and UO_817 (O_817,N_8095,N_8743);
nand UO_818 (O_818,N_9974,N_9116);
and UO_819 (O_819,N_8560,N_9801);
and UO_820 (O_820,N_8327,N_9898);
and UO_821 (O_821,N_9357,N_8655);
and UO_822 (O_822,N_9180,N_8073);
nand UO_823 (O_823,N_9099,N_8540);
or UO_824 (O_824,N_9550,N_9515);
nand UO_825 (O_825,N_9482,N_8322);
and UO_826 (O_826,N_9778,N_9545);
nor UO_827 (O_827,N_8193,N_8871);
and UO_828 (O_828,N_8796,N_8445);
or UO_829 (O_829,N_8808,N_9900);
or UO_830 (O_830,N_9001,N_8525);
and UO_831 (O_831,N_8337,N_9853);
xnor UO_832 (O_832,N_9770,N_8603);
or UO_833 (O_833,N_8053,N_9316);
and UO_834 (O_834,N_8773,N_9385);
and UO_835 (O_835,N_9737,N_8799);
nor UO_836 (O_836,N_8139,N_8236);
or UO_837 (O_837,N_8118,N_8018);
and UO_838 (O_838,N_9297,N_9205);
or UO_839 (O_839,N_8464,N_8413);
or UO_840 (O_840,N_8401,N_9102);
nand UO_841 (O_841,N_8010,N_9229);
or UO_842 (O_842,N_9401,N_9053);
and UO_843 (O_843,N_9508,N_9875);
or UO_844 (O_844,N_9273,N_9347);
or UO_845 (O_845,N_8436,N_9354);
and UO_846 (O_846,N_9468,N_9298);
nand UO_847 (O_847,N_9789,N_8009);
and UO_848 (O_848,N_9340,N_8277);
nand UO_849 (O_849,N_8225,N_9942);
nor UO_850 (O_850,N_8395,N_8453);
nor UO_851 (O_851,N_8763,N_9731);
and UO_852 (O_852,N_9712,N_8378);
and UO_853 (O_853,N_8962,N_9807);
nand UO_854 (O_854,N_9798,N_9248);
nand UO_855 (O_855,N_8219,N_9780);
nand UO_856 (O_856,N_8153,N_8670);
or UO_857 (O_857,N_9202,N_9000);
nand UO_858 (O_858,N_9958,N_9466);
nor UO_859 (O_859,N_8004,N_9083);
nand UO_860 (O_860,N_8893,N_8734);
nor UO_861 (O_861,N_9676,N_8921);
nand UO_862 (O_862,N_8911,N_9470);
nand UO_863 (O_863,N_8180,N_8787);
or UO_864 (O_864,N_8412,N_9533);
or UO_865 (O_865,N_8262,N_8630);
or UO_866 (O_866,N_8817,N_9156);
nor UO_867 (O_867,N_8870,N_9633);
or UO_868 (O_868,N_8063,N_9104);
nand UO_869 (O_869,N_9299,N_8970);
or UO_870 (O_870,N_8383,N_9308);
and UO_871 (O_871,N_9120,N_8435);
nor UO_872 (O_872,N_9076,N_8029);
and UO_873 (O_873,N_9029,N_8931);
or UO_874 (O_874,N_8758,N_9137);
nor UO_875 (O_875,N_9980,N_9314);
or UO_876 (O_876,N_8372,N_8208);
or UO_877 (O_877,N_8359,N_8833);
and UO_878 (O_878,N_9857,N_8045);
nand UO_879 (O_879,N_8848,N_8273);
nor UO_880 (O_880,N_9177,N_9350);
nor UO_881 (O_881,N_8978,N_8628);
and UO_882 (O_882,N_9363,N_8839);
or UO_883 (O_883,N_8215,N_9865);
nand UO_884 (O_884,N_8417,N_8681);
nand UO_885 (O_885,N_8440,N_9999);
nor UO_886 (O_886,N_9935,N_9964);
nand UO_887 (O_887,N_8688,N_9206);
or UO_888 (O_888,N_8977,N_9688);
or UO_889 (O_889,N_9787,N_8971);
or UO_890 (O_890,N_9348,N_8055);
or UO_891 (O_891,N_8333,N_9068);
nand UO_892 (O_892,N_9094,N_8292);
or UO_893 (O_893,N_9445,N_9051);
nand UO_894 (O_894,N_8933,N_9386);
nand UO_895 (O_895,N_9393,N_9450);
or UO_896 (O_896,N_8813,N_9493);
nor UO_897 (O_897,N_9338,N_9106);
and UO_898 (O_898,N_8482,N_9986);
and UO_899 (O_899,N_9118,N_8643);
nand UO_900 (O_900,N_9813,N_9247);
and UO_901 (O_901,N_8234,N_8620);
nor UO_902 (O_902,N_8772,N_8293);
and UO_903 (O_903,N_9194,N_9286);
nor UO_904 (O_904,N_9756,N_8557);
or UO_905 (O_905,N_9418,N_8635);
nor UO_906 (O_906,N_9423,N_8038);
or UO_907 (O_907,N_9077,N_8035);
nand UO_908 (O_908,N_8874,N_9390);
and UO_909 (O_909,N_8946,N_9351);
nor UO_910 (O_910,N_8878,N_8012);
nor UO_911 (O_911,N_8532,N_9558);
and UO_912 (O_912,N_8084,N_9987);
and UO_913 (O_913,N_9015,N_9023);
nand UO_914 (O_914,N_9039,N_8245);
nand UO_915 (O_915,N_8074,N_8156);
and UO_916 (O_916,N_9852,N_9434);
nor UO_917 (O_917,N_8017,N_8311);
nand UO_918 (O_918,N_9178,N_8669);
or UO_919 (O_919,N_8437,N_9646);
nand UO_920 (O_920,N_9021,N_8705);
and UO_921 (O_921,N_9513,N_8366);
nor UO_922 (O_922,N_9554,N_8054);
nand UO_923 (O_923,N_9729,N_8949);
or UO_924 (O_924,N_9922,N_9435);
xnor UO_925 (O_925,N_8940,N_9372);
and UO_926 (O_926,N_9312,N_9741);
or UO_927 (O_927,N_8610,N_9242);
nor UO_928 (O_928,N_8252,N_9201);
or UO_929 (O_929,N_9193,N_8851);
nor UO_930 (O_930,N_9336,N_8352);
nor UO_931 (O_931,N_8784,N_9127);
or UO_932 (O_932,N_9333,N_8489);
and UO_933 (O_933,N_8766,N_9793);
nand UO_934 (O_934,N_8296,N_9325);
and UO_935 (O_935,N_9040,N_8712);
or UO_936 (O_936,N_9963,N_8882);
or UO_937 (O_937,N_8613,N_9081);
and UO_938 (O_938,N_8207,N_8768);
and UO_939 (O_939,N_9525,N_9682);
or UO_940 (O_940,N_9060,N_9759);
and UO_941 (O_941,N_9797,N_8285);
or UO_942 (O_942,N_8051,N_9555);
nand UO_943 (O_943,N_8324,N_8535);
nor UO_944 (O_944,N_8088,N_9716);
or UO_945 (O_945,N_9135,N_8795);
nor UO_946 (O_946,N_8138,N_9669);
and UO_947 (O_947,N_8448,N_9622);
nor UO_948 (O_948,N_9292,N_8531);
and UO_949 (O_949,N_9921,N_8159);
and UO_950 (O_950,N_9488,N_9207);
or UO_951 (O_951,N_9598,N_8834);
nor UO_952 (O_952,N_9483,N_8100);
nand UO_953 (O_953,N_8122,N_9893);
xnor UO_954 (O_954,N_8636,N_9667);
xnor UO_955 (O_955,N_9188,N_8309);
nand UO_956 (O_956,N_9315,N_9151);
or UO_957 (O_957,N_8684,N_9014);
nor UO_958 (O_958,N_9252,N_9873);
and UO_959 (O_959,N_8770,N_9380);
nor UO_960 (O_960,N_8148,N_9680);
nand UO_961 (O_961,N_9909,N_9085);
or UO_962 (O_962,N_9849,N_8377);
nor UO_963 (O_963,N_8316,N_9783);
and UO_964 (O_964,N_9042,N_8718);
and UO_965 (O_965,N_9736,N_8691);
nor UO_966 (O_966,N_8514,N_8750);
nor UO_967 (O_967,N_8142,N_9938);
nand UO_968 (O_968,N_9008,N_9984);
xnor UO_969 (O_969,N_9157,N_9310);
nor UO_970 (O_970,N_8711,N_9879);
and UO_971 (O_971,N_9925,N_9245);
nor UO_972 (O_972,N_8653,N_8189);
nand UO_973 (O_973,N_8499,N_8478);
nor UO_974 (O_974,N_9861,N_9790);
nor UO_975 (O_975,N_8935,N_9277);
and UO_976 (O_976,N_8209,N_8797);
nand UO_977 (O_977,N_8923,N_9833);
nand UO_978 (O_978,N_8914,N_9715);
nand UO_979 (O_979,N_8432,N_8476);
and UO_980 (O_980,N_8836,N_9657);
nor UO_981 (O_981,N_8022,N_9406);
nor UO_982 (O_982,N_9779,N_8583);
xor UO_983 (O_983,N_8259,N_8658);
nor UO_984 (O_984,N_9457,N_9761);
or UO_985 (O_985,N_8047,N_9703);
and UO_986 (O_986,N_9745,N_8109);
nand UO_987 (O_987,N_9851,N_9595);
nand UO_988 (O_988,N_9153,N_9596);
and UO_989 (O_989,N_9726,N_8454);
nor UO_990 (O_990,N_9838,N_9663);
or UO_991 (O_991,N_8006,N_9753);
and UO_992 (O_992,N_8062,N_9899);
or UO_993 (O_993,N_8350,N_9343);
nand UO_994 (O_994,N_8950,N_9579);
nand UO_995 (O_995,N_9848,N_8831);
or UO_996 (O_996,N_8346,N_8030);
nand UO_997 (O_997,N_9010,N_8780);
nand UO_998 (O_998,N_9827,N_8974);
and UO_999 (O_999,N_8767,N_8438);
and UO_1000 (O_1000,N_8364,N_8283);
and UO_1001 (O_1001,N_9310,N_9449);
and UO_1002 (O_1002,N_8808,N_8662);
or UO_1003 (O_1003,N_8517,N_9490);
or UO_1004 (O_1004,N_9079,N_9233);
and UO_1005 (O_1005,N_9485,N_9505);
nand UO_1006 (O_1006,N_8029,N_9508);
nor UO_1007 (O_1007,N_9705,N_8581);
nand UO_1008 (O_1008,N_9386,N_8930);
nand UO_1009 (O_1009,N_9433,N_8129);
nor UO_1010 (O_1010,N_9590,N_8177);
or UO_1011 (O_1011,N_9107,N_8787);
nand UO_1012 (O_1012,N_9256,N_8471);
and UO_1013 (O_1013,N_9812,N_9503);
nor UO_1014 (O_1014,N_9148,N_8256);
nand UO_1015 (O_1015,N_8820,N_9447);
or UO_1016 (O_1016,N_9345,N_9002);
and UO_1017 (O_1017,N_9958,N_9767);
nand UO_1018 (O_1018,N_9930,N_8118);
nand UO_1019 (O_1019,N_8740,N_9700);
and UO_1020 (O_1020,N_8934,N_8480);
and UO_1021 (O_1021,N_8076,N_9053);
nand UO_1022 (O_1022,N_9033,N_8629);
and UO_1023 (O_1023,N_9443,N_8098);
nand UO_1024 (O_1024,N_8705,N_9546);
nand UO_1025 (O_1025,N_9227,N_8102);
or UO_1026 (O_1026,N_9069,N_9676);
or UO_1027 (O_1027,N_8668,N_9807);
nand UO_1028 (O_1028,N_8407,N_9460);
or UO_1029 (O_1029,N_9523,N_9429);
and UO_1030 (O_1030,N_9533,N_8872);
or UO_1031 (O_1031,N_8389,N_9043);
nand UO_1032 (O_1032,N_8870,N_9356);
or UO_1033 (O_1033,N_8381,N_8646);
and UO_1034 (O_1034,N_8861,N_9895);
nand UO_1035 (O_1035,N_8850,N_8606);
nor UO_1036 (O_1036,N_8972,N_9125);
nand UO_1037 (O_1037,N_8499,N_9105);
and UO_1038 (O_1038,N_9834,N_8096);
nand UO_1039 (O_1039,N_9002,N_8925);
and UO_1040 (O_1040,N_8302,N_8198);
or UO_1041 (O_1041,N_9910,N_9197);
or UO_1042 (O_1042,N_9539,N_8937);
nand UO_1043 (O_1043,N_9717,N_9979);
nor UO_1044 (O_1044,N_9929,N_8448);
nor UO_1045 (O_1045,N_8478,N_8553);
or UO_1046 (O_1046,N_8101,N_9201);
nand UO_1047 (O_1047,N_8373,N_9482);
nor UO_1048 (O_1048,N_9308,N_8150);
nor UO_1049 (O_1049,N_9181,N_8668);
nand UO_1050 (O_1050,N_9605,N_9559);
nor UO_1051 (O_1051,N_8829,N_8380);
or UO_1052 (O_1052,N_8142,N_9067);
and UO_1053 (O_1053,N_8432,N_9895);
nand UO_1054 (O_1054,N_8363,N_9503);
and UO_1055 (O_1055,N_8963,N_9775);
or UO_1056 (O_1056,N_9500,N_8475);
and UO_1057 (O_1057,N_8134,N_9064);
nor UO_1058 (O_1058,N_9137,N_9171);
or UO_1059 (O_1059,N_9495,N_9486);
nor UO_1060 (O_1060,N_9800,N_8671);
or UO_1061 (O_1061,N_9043,N_9899);
and UO_1062 (O_1062,N_8844,N_8799);
nor UO_1063 (O_1063,N_8174,N_8887);
or UO_1064 (O_1064,N_9641,N_8765);
nor UO_1065 (O_1065,N_8056,N_9199);
nor UO_1066 (O_1066,N_9687,N_9126);
nor UO_1067 (O_1067,N_9060,N_8414);
nand UO_1068 (O_1068,N_9445,N_9749);
and UO_1069 (O_1069,N_8400,N_9051);
nand UO_1070 (O_1070,N_9641,N_9665);
nand UO_1071 (O_1071,N_8140,N_9851);
or UO_1072 (O_1072,N_8908,N_8552);
nand UO_1073 (O_1073,N_9695,N_8061);
or UO_1074 (O_1074,N_9033,N_9011);
or UO_1075 (O_1075,N_9760,N_8604);
and UO_1076 (O_1076,N_8608,N_9331);
and UO_1077 (O_1077,N_8004,N_8595);
or UO_1078 (O_1078,N_9538,N_8406);
nor UO_1079 (O_1079,N_8379,N_8860);
nand UO_1080 (O_1080,N_8381,N_8302);
nor UO_1081 (O_1081,N_8888,N_8246);
or UO_1082 (O_1082,N_8324,N_9292);
nor UO_1083 (O_1083,N_9468,N_8558);
and UO_1084 (O_1084,N_8079,N_9176);
nand UO_1085 (O_1085,N_8767,N_8248);
nor UO_1086 (O_1086,N_9972,N_9650);
nor UO_1087 (O_1087,N_8062,N_8737);
or UO_1088 (O_1088,N_9212,N_9159);
or UO_1089 (O_1089,N_8753,N_8248);
nand UO_1090 (O_1090,N_9628,N_8437);
and UO_1091 (O_1091,N_8017,N_8694);
or UO_1092 (O_1092,N_8679,N_8427);
nand UO_1093 (O_1093,N_9439,N_8875);
nor UO_1094 (O_1094,N_8956,N_9641);
nand UO_1095 (O_1095,N_9086,N_9526);
or UO_1096 (O_1096,N_8176,N_9683);
nor UO_1097 (O_1097,N_8349,N_9512);
nand UO_1098 (O_1098,N_9639,N_8659);
nand UO_1099 (O_1099,N_9974,N_8394);
or UO_1100 (O_1100,N_9194,N_9018);
nor UO_1101 (O_1101,N_8200,N_9628);
nand UO_1102 (O_1102,N_9001,N_9436);
nor UO_1103 (O_1103,N_8928,N_8475);
nand UO_1104 (O_1104,N_8262,N_8927);
nand UO_1105 (O_1105,N_8597,N_8376);
or UO_1106 (O_1106,N_9439,N_9885);
nand UO_1107 (O_1107,N_8793,N_9403);
or UO_1108 (O_1108,N_8514,N_8120);
or UO_1109 (O_1109,N_8337,N_8111);
nand UO_1110 (O_1110,N_9957,N_8682);
or UO_1111 (O_1111,N_9372,N_8371);
or UO_1112 (O_1112,N_8737,N_9453);
or UO_1113 (O_1113,N_8870,N_8727);
nor UO_1114 (O_1114,N_9105,N_9962);
nor UO_1115 (O_1115,N_9987,N_9028);
and UO_1116 (O_1116,N_8366,N_8517);
and UO_1117 (O_1117,N_8253,N_8928);
xor UO_1118 (O_1118,N_8466,N_9142);
or UO_1119 (O_1119,N_8922,N_8053);
nor UO_1120 (O_1120,N_9574,N_9685);
or UO_1121 (O_1121,N_8404,N_8862);
or UO_1122 (O_1122,N_8089,N_8744);
or UO_1123 (O_1123,N_8190,N_8570);
and UO_1124 (O_1124,N_9125,N_9902);
and UO_1125 (O_1125,N_8702,N_9162);
and UO_1126 (O_1126,N_8105,N_9354);
nor UO_1127 (O_1127,N_9675,N_8586);
and UO_1128 (O_1128,N_8755,N_9964);
or UO_1129 (O_1129,N_8858,N_8092);
or UO_1130 (O_1130,N_9620,N_9468);
nor UO_1131 (O_1131,N_9876,N_8321);
nor UO_1132 (O_1132,N_9730,N_9614);
or UO_1133 (O_1133,N_9660,N_9975);
nand UO_1134 (O_1134,N_9352,N_9915);
nor UO_1135 (O_1135,N_9847,N_9875);
nand UO_1136 (O_1136,N_9617,N_9099);
or UO_1137 (O_1137,N_8644,N_9465);
nand UO_1138 (O_1138,N_8767,N_9589);
nand UO_1139 (O_1139,N_9154,N_8658);
and UO_1140 (O_1140,N_8443,N_9304);
or UO_1141 (O_1141,N_8542,N_8656);
nor UO_1142 (O_1142,N_8012,N_8161);
and UO_1143 (O_1143,N_8989,N_8736);
nand UO_1144 (O_1144,N_8205,N_9820);
or UO_1145 (O_1145,N_8320,N_8800);
nand UO_1146 (O_1146,N_8760,N_9042);
nand UO_1147 (O_1147,N_9833,N_9616);
xor UO_1148 (O_1148,N_9222,N_9617);
or UO_1149 (O_1149,N_9359,N_8267);
nor UO_1150 (O_1150,N_9473,N_9568);
or UO_1151 (O_1151,N_9084,N_9787);
or UO_1152 (O_1152,N_8260,N_9563);
and UO_1153 (O_1153,N_8981,N_8313);
nand UO_1154 (O_1154,N_8482,N_9969);
nor UO_1155 (O_1155,N_9065,N_9308);
and UO_1156 (O_1156,N_8663,N_8379);
nand UO_1157 (O_1157,N_8581,N_8807);
nor UO_1158 (O_1158,N_8297,N_8738);
nand UO_1159 (O_1159,N_8716,N_8859);
and UO_1160 (O_1160,N_9440,N_8552);
and UO_1161 (O_1161,N_9020,N_9450);
nand UO_1162 (O_1162,N_8182,N_9420);
and UO_1163 (O_1163,N_9783,N_8242);
and UO_1164 (O_1164,N_9715,N_8887);
nand UO_1165 (O_1165,N_8351,N_9845);
nand UO_1166 (O_1166,N_9289,N_9362);
nor UO_1167 (O_1167,N_9560,N_8524);
nand UO_1168 (O_1168,N_8652,N_9174);
and UO_1169 (O_1169,N_9289,N_8593);
or UO_1170 (O_1170,N_9182,N_9881);
xnor UO_1171 (O_1171,N_8030,N_8492);
and UO_1172 (O_1172,N_9153,N_8495);
nor UO_1173 (O_1173,N_8418,N_8108);
and UO_1174 (O_1174,N_9033,N_8912);
and UO_1175 (O_1175,N_9979,N_9220);
nand UO_1176 (O_1176,N_8684,N_8076);
or UO_1177 (O_1177,N_9503,N_9884);
or UO_1178 (O_1178,N_8347,N_8301);
and UO_1179 (O_1179,N_8414,N_8106);
and UO_1180 (O_1180,N_9338,N_8010);
or UO_1181 (O_1181,N_8555,N_9045);
and UO_1182 (O_1182,N_8695,N_9911);
and UO_1183 (O_1183,N_9146,N_8648);
or UO_1184 (O_1184,N_9914,N_9808);
or UO_1185 (O_1185,N_8154,N_9895);
nand UO_1186 (O_1186,N_9975,N_8096);
and UO_1187 (O_1187,N_8896,N_9883);
nor UO_1188 (O_1188,N_8070,N_8749);
nor UO_1189 (O_1189,N_8614,N_8031);
nand UO_1190 (O_1190,N_9350,N_9884);
nand UO_1191 (O_1191,N_9480,N_8735);
nor UO_1192 (O_1192,N_8967,N_8060);
and UO_1193 (O_1193,N_9332,N_9397);
nand UO_1194 (O_1194,N_8601,N_9111);
nor UO_1195 (O_1195,N_8915,N_8080);
or UO_1196 (O_1196,N_8922,N_8949);
nor UO_1197 (O_1197,N_8437,N_8107);
or UO_1198 (O_1198,N_8111,N_8292);
and UO_1199 (O_1199,N_9265,N_9254);
and UO_1200 (O_1200,N_8609,N_9999);
nor UO_1201 (O_1201,N_9974,N_8613);
or UO_1202 (O_1202,N_8103,N_9900);
or UO_1203 (O_1203,N_9829,N_9492);
nand UO_1204 (O_1204,N_8065,N_9496);
nand UO_1205 (O_1205,N_9956,N_9479);
nand UO_1206 (O_1206,N_9408,N_8428);
nand UO_1207 (O_1207,N_9595,N_9823);
or UO_1208 (O_1208,N_8099,N_8704);
or UO_1209 (O_1209,N_9819,N_8189);
or UO_1210 (O_1210,N_8344,N_9563);
and UO_1211 (O_1211,N_8108,N_9533);
nor UO_1212 (O_1212,N_8047,N_8479);
or UO_1213 (O_1213,N_8511,N_8191);
nor UO_1214 (O_1214,N_8313,N_9080);
and UO_1215 (O_1215,N_8998,N_9092);
nor UO_1216 (O_1216,N_9862,N_9798);
and UO_1217 (O_1217,N_9875,N_8742);
nor UO_1218 (O_1218,N_8293,N_8132);
nor UO_1219 (O_1219,N_9867,N_9072);
nand UO_1220 (O_1220,N_8024,N_9824);
and UO_1221 (O_1221,N_8916,N_8053);
nand UO_1222 (O_1222,N_8724,N_8660);
and UO_1223 (O_1223,N_8930,N_8896);
or UO_1224 (O_1224,N_8638,N_9840);
and UO_1225 (O_1225,N_9040,N_9711);
xnor UO_1226 (O_1226,N_8514,N_9718);
or UO_1227 (O_1227,N_8654,N_9560);
nand UO_1228 (O_1228,N_9767,N_9745);
or UO_1229 (O_1229,N_9241,N_9134);
and UO_1230 (O_1230,N_9178,N_8857);
and UO_1231 (O_1231,N_8156,N_9653);
nor UO_1232 (O_1232,N_8485,N_8694);
nand UO_1233 (O_1233,N_9218,N_9981);
nand UO_1234 (O_1234,N_8977,N_8397);
and UO_1235 (O_1235,N_8282,N_9431);
and UO_1236 (O_1236,N_8026,N_8289);
or UO_1237 (O_1237,N_9863,N_8860);
and UO_1238 (O_1238,N_8113,N_8600);
and UO_1239 (O_1239,N_8402,N_9814);
and UO_1240 (O_1240,N_9979,N_9593);
and UO_1241 (O_1241,N_9072,N_9901);
and UO_1242 (O_1242,N_8201,N_8651);
nand UO_1243 (O_1243,N_8102,N_8448);
and UO_1244 (O_1244,N_8941,N_9718);
nand UO_1245 (O_1245,N_8696,N_8008);
nand UO_1246 (O_1246,N_9893,N_8152);
nor UO_1247 (O_1247,N_9009,N_9026);
nor UO_1248 (O_1248,N_9276,N_8646);
nand UO_1249 (O_1249,N_8110,N_9877);
nor UO_1250 (O_1250,N_9331,N_9308);
nor UO_1251 (O_1251,N_8965,N_9934);
and UO_1252 (O_1252,N_8666,N_8072);
and UO_1253 (O_1253,N_8206,N_9000);
nand UO_1254 (O_1254,N_8266,N_9719);
nand UO_1255 (O_1255,N_9902,N_9849);
and UO_1256 (O_1256,N_8914,N_8494);
nor UO_1257 (O_1257,N_8920,N_8884);
or UO_1258 (O_1258,N_8218,N_8432);
and UO_1259 (O_1259,N_8766,N_8968);
and UO_1260 (O_1260,N_9450,N_9982);
or UO_1261 (O_1261,N_9975,N_8293);
and UO_1262 (O_1262,N_9768,N_9628);
and UO_1263 (O_1263,N_9564,N_8084);
xnor UO_1264 (O_1264,N_8541,N_8784);
and UO_1265 (O_1265,N_9929,N_8907);
and UO_1266 (O_1266,N_9249,N_9740);
or UO_1267 (O_1267,N_8786,N_9538);
nand UO_1268 (O_1268,N_8068,N_9343);
nand UO_1269 (O_1269,N_8354,N_8389);
or UO_1270 (O_1270,N_8148,N_8370);
and UO_1271 (O_1271,N_8832,N_9528);
nor UO_1272 (O_1272,N_9997,N_8094);
or UO_1273 (O_1273,N_9798,N_9724);
nor UO_1274 (O_1274,N_8609,N_8255);
and UO_1275 (O_1275,N_9339,N_8673);
and UO_1276 (O_1276,N_8638,N_9924);
nor UO_1277 (O_1277,N_8385,N_9102);
or UO_1278 (O_1278,N_9746,N_8920);
nand UO_1279 (O_1279,N_9936,N_9750);
or UO_1280 (O_1280,N_9397,N_8798);
and UO_1281 (O_1281,N_9600,N_8327);
and UO_1282 (O_1282,N_9730,N_8847);
nand UO_1283 (O_1283,N_8187,N_9317);
and UO_1284 (O_1284,N_9435,N_9105);
nor UO_1285 (O_1285,N_8286,N_9095);
and UO_1286 (O_1286,N_8831,N_9542);
or UO_1287 (O_1287,N_9767,N_9693);
nor UO_1288 (O_1288,N_9902,N_9189);
nand UO_1289 (O_1289,N_8910,N_8900);
and UO_1290 (O_1290,N_9325,N_8518);
nor UO_1291 (O_1291,N_8178,N_8430);
or UO_1292 (O_1292,N_8133,N_9648);
and UO_1293 (O_1293,N_9677,N_8664);
nor UO_1294 (O_1294,N_8384,N_8889);
and UO_1295 (O_1295,N_9771,N_8996);
nor UO_1296 (O_1296,N_9926,N_9061);
nand UO_1297 (O_1297,N_9584,N_8414);
nand UO_1298 (O_1298,N_9052,N_9469);
or UO_1299 (O_1299,N_8981,N_8099);
nor UO_1300 (O_1300,N_8137,N_9366);
nor UO_1301 (O_1301,N_8627,N_9923);
or UO_1302 (O_1302,N_8097,N_9290);
nand UO_1303 (O_1303,N_9863,N_9214);
or UO_1304 (O_1304,N_8861,N_9532);
and UO_1305 (O_1305,N_8771,N_8129);
nor UO_1306 (O_1306,N_9214,N_8025);
or UO_1307 (O_1307,N_8794,N_8554);
nor UO_1308 (O_1308,N_8916,N_9167);
nand UO_1309 (O_1309,N_9311,N_9453);
or UO_1310 (O_1310,N_8144,N_8054);
xnor UO_1311 (O_1311,N_8834,N_9028);
or UO_1312 (O_1312,N_8982,N_8441);
nand UO_1313 (O_1313,N_9293,N_8824);
or UO_1314 (O_1314,N_9601,N_9730);
and UO_1315 (O_1315,N_9274,N_9327);
nor UO_1316 (O_1316,N_8044,N_8174);
and UO_1317 (O_1317,N_8368,N_9726);
or UO_1318 (O_1318,N_8494,N_8744);
nand UO_1319 (O_1319,N_8441,N_8406);
or UO_1320 (O_1320,N_9546,N_8947);
and UO_1321 (O_1321,N_8134,N_8827);
or UO_1322 (O_1322,N_9593,N_9373);
nor UO_1323 (O_1323,N_8277,N_9902);
nor UO_1324 (O_1324,N_9658,N_8426);
nor UO_1325 (O_1325,N_8789,N_8276);
nand UO_1326 (O_1326,N_9320,N_8836);
and UO_1327 (O_1327,N_8600,N_8140);
nand UO_1328 (O_1328,N_9052,N_9638);
nand UO_1329 (O_1329,N_9768,N_9338);
nor UO_1330 (O_1330,N_8358,N_8450);
or UO_1331 (O_1331,N_8282,N_8599);
nand UO_1332 (O_1332,N_9563,N_8783);
nand UO_1333 (O_1333,N_8061,N_9070);
nand UO_1334 (O_1334,N_9798,N_9267);
or UO_1335 (O_1335,N_9724,N_8766);
and UO_1336 (O_1336,N_9498,N_8945);
nor UO_1337 (O_1337,N_8384,N_9142);
nor UO_1338 (O_1338,N_8753,N_9943);
or UO_1339 (O_1339,N_9269,N_8132);
nand UO_1340 (O_1340,N_9860,N_9184);
or UO_1341 (O_1341,N_9221,N_9139);
nor UO_1342 (O_1342,N_9441,N_8031);
nand UO_1343 (O_1343,N_9409,N_9839);
or UO_1344 (O_1344,N_9649,N_8850);
nand UO_1345 (O_1345,N_9156,N_9484);
and UO_1346 (O_1346,N_8066,N_8383);
nor UO_1347 (O_1347,N_9619,N_8665);
or UO_1348 (O_1348,N_9226,N_8388);
and UO_1349 (O_1349,N_9879,N_8400);
nor UO_1350 (O_1350,N_9416,N_9764);
or UO_1351 (O_1351,N_8309,N_8662);
nand UO_1352 (O_1352,N_9965,N_8830);
nor UO_1353 (O_1353,N_8509,N_8499);
nand UO_1354 (O_1354,N_8971,N_9337);
nand UO_1355 (O_1355,N_9622,N_8585);
or UO_1356 (O_1356,N_8633,N_9327);
and UO_1357 (O_1357,N_9620,N_8732);
nor UO_1358 (O_1358,N_8515,N_8816);
and UO_1359 (O_1359,N_8897,N_9341);
or UO_1360 (O_1360,N_9263,N_9211);
nor UO_1361 (O_1361,N_8132,N_8502);
and UO_1362 (O_1362,N_9885,N_8105);
and UO_1363 (O_1363,N_8927,N_8212);
nand UO_1364 (O_1364,N_9109,N_9221);
nand UO_1365 (O_1365,N_9074,N_9399);
and UO_1366 (O_1366,N_9251,N_8601);
xnor UO_1367 (O_1367,N_9611,N_8809);
or UO_1368 (O_1368,N_8452,N_8658);
nor UO_1369 (O_1369,N_8711,N_9485);
nand UO_1370 (O_1370,N_9256,N_9999);
and UO_1371 (O_1371,N_9379,N_9197);
and UO_1372 (O_1372,N_9011,N_9139);
nor UO_1373 (O_1373,N_9623,N_9148);
or UO_1374 (O_1374,N_9123,N_9804);
and UO_1375 (O_1375,N_9148,N_9986);
and UO_1376 (O_1376,N_8662,N_9701);
and UO_1377 (O_1377,N_9896,N_9497);
nand UO_1378 (O_1378,N_9607,N_8646);
nor UO_1379 (O_1379,N_8435,N_8214);
nor UO_1380 (O_1380,N_8197,N_8061);
or UO_1381 (O_1381,N_8153,N_8345);
nor UO_1382 (O_1382,N_8509,N_8143);
or UO_1383 (O_1383,N_8563,N_8029);
nor UO_1384 (O_1384,N_9420,N_9272);
xnor UO_1385 (O_1385,N_8883,N_9654);
or UO_1386 (O_1386,N_9237,N_9483);
nand UO_1387 (O_1387,N_8435,N_8172);
nand UO_1388 (O_1388,N_9960,N_9667);
and UO_1389 (O_1389,N_9963,N_9229);
and UO_1390 (O_1390,N_8261,N_9443);
xnor UO_1391 (O_1391,N_9954,N_9991);
or UO_1392 (O_1392,N_8597,N_8079);
nor UO_1393 (O_1393,N_9682,N_9620);
and UO_1394 (O_1394,N_8273,N_9794);
nand UO_1395 (O_1395,N_8972,N_8569);
xnor UO_1396 (O_1396,N_8472,N_8093);
nand UO_1397 (O_1397,N_9025,N_9609);
nor UO_1398 (O_1398,N_9007,N_8354);
or UO_1399 (O_1399,N_8450,N_9326);
nand UO_1400 (O_1400,N_8163,N_9047);
or UO_1401 (O_1401,N_8324,N_9207);
nor UO_1402 (O_1402,N_8649,N_9232);
nand UO_1403 (O_1403,N_9289,N_9041);
nor UO_1404 (O_1404,N_9634,N_9971);
nor UO_1405 (O_1405,N_8035,N_9939);
and UO_1406 (O_1406,N_9894,N_8116);
and UO_1407 (O_1407,N_9826,N_8922);
xor UO_1408 (O_1408,N_8019,N_8376);
nor UO_1409 (O_1409,N_8208,N_8897);
or UO_1410 (O_1410,N_8660,N_9199);
nand UO_1411 (O_1411,N_9987,N_9523);
nor UO_1412 (O_1412,N_8216,N_9693);
nor UO_1413 (O_1413,N_8755,N_8081);
nand UO_1414 (O_1414,N_8161,N_9231);
nand UO_1415 (O_1415,N_9047,N_9590);
and UO_1416 (O_1416,N_9844,N_8011);
and UO_1417 (O_1417,N_9649,N_9820);
and UO_1418 (O_1418,N_8633,N_8330);
nor UO_1419 (O_1419,N_8961,N_9080);
or UO_1420 (O_1420,N_8229,N_8294);
and UO_1421 (O_1421,N_9716,N_8936);
nand UO_1422 (O_1422,N_8917,N_9071);
xor UO_1423 (O_1423,N_8629,N_9876);
and UO_1424 (O_1424,N_8296,N_8669);
and UO_1425 (O_1425,N_9036,N_8312);
or UO_1426 (O_1426,N_9724,N_9116);
nand UO_1427 (O_1427,N_8015,N_8672);
nand UO_1428 (O_1428,N_8445,N_8327);
nor UO_1429 (O_1429,N_9504,N_9138);
or UO_1430 (O_1430,N_8302,N_9854);
nor UO_1431 (O_1431,N_8085,N_8708);
nand UO_1432 (O_1432,N_9855,N_8055);
nor UO_1433 (O_1433,N_9513,N_9623);
nor UO_1434 (O_1434,N_9302,N_8503);
nand UO_1435 (O_1435,N_9284,N_9600);
or UO_1436 (O_1436,N_9964,N_8129);
nor UO_1437 (O_1437,N_8261,N_9664);
nor UO_1438 (O_1438,N_9307,N_8798);
nor UO_1439 (O_1439,N_8762,N_9821);
nor UO_1440 (O_1440,N_9101,N_9375);
or UO_1441 (O_1441,N_9767,N_9721);
or UO_1442 (O_1442,N_8310,N_9783);
nand UO_1443 (O_1443,N_9520,N_9459);
or UO_1444 (O_1444,N_8520,N_9990);
and UO_1445 (O_1445,N_8942,N_9375);
nor UO_1446 (O_1446,N_9484,N_8044);
and UO_1447 (O_1447,N_9856,N_9879);
or UO_1448 (O_1448,N_8596,N_9894);
and UO_1449 (O_1449,N_9819,N_8161);
nor UO_1450 (O_1450,N_9627,N_9811);
nor UO_1451 (O_1451,N_9528,N_8471);
nor UO_1452 (O_1452,N_9554,N_9323);
and UO_1453 (O_1453,N_8162,N_9686);
or UO_1454 (O_1454,N_8452,N_8061);
nand UO_1455 (O_1455,N_8183,N_9930);
and UO_1456 (O_1456,N_9844,N_9727);
or UO_1457 (O_1457,N_9283,N_8438);
or UO_1458 (O_1458,N_9374,N_9912);
nand UO_1459 (O_1459,N_9208,N_9277);
and UO_1460 (O_1460,N_9821,N_9674);
nor UO_1461 (O_1461,N_8992,N_9211);
nor UO_1462 (O_1462,N_8560,N_9449);
xor UO_1463 (O_1463,N_8568,N_9427);
or UO_1464 (O_1464,N_9538,N_8565);
xnor UO_1465 (O_1465,N_8759,N_8073);
or UO_1466 (O_1466,N_9759,N_8413);
nand UO_1467 (O_1467,N_9852,N_9299);
nor UO_1468 (O_1468,N_8921,N_9139);
and UO_1469 (O_1469,N_8844,N_8657);
or UO_1470 (O_1470,N_9092,N_9572);
nor UO_1471 (O_1471,N_8546,N_9014);
nand UO_1472 (O_1472,N_8113,N_8032);
nor UO_1473 (O_1473,N_8340,N_9977);
or UO_1474 (O_1474,N_8118,N_9873);
and UO_1475 (O_1475,N_9652,N_8032);
or UO_1476 (O_1476,N_9220,N_9692);
or UO_1477 (O_1477,N_8302,N_9183);
or UO_1478 (O_1478,N_8082,N_8831);
nor UO_1479 (O_1479,N_9169,N_8973);
or UO_1480 (O_1480,N_8672,N_8947);
or UO_1481 (O_1481,N_9690,N_9775);
nor UO_1482 (O_1482,N_9957,N_8821);
nor UO_1483 (O_1483,N_8777,N_9551);
nor UO_1484 (O_1484,N_9170,N_9289);
nand UO_1485 (O_1485,N_8413,N_8909);
nor UO_1486 (O_1486,N_8050,N_9962);
nor UO_1487 (O_1487,N_8365,N_9541);
or UO_1488 (O_1488,N_8898,N_9146);
nand UO_1489 (O_1489,N_8404,N_9744);
or UO_1490 (O_1490,N_8546,N_9784);
or UO_1491 (O_1491,N_9756,N_8171);
and UO_1492 (O_1492,N_8939,N_8438);
nor UO_1493 (O_1493,N_9533,N_8805);
nand UO_1494 (O_1494,N_9723,N_9987);
nand UO_1495 (O_1495,N_8173,N_9756);
or UO_1496 (O_1496,N_8961,N_9469);
nand UO_1497 (O_1497,N_8935,N_9296);
and UO_1498 (O_1498,N_9083,N_8338);
and UO_1499 (O_1499,N_9852,N_8351);
endmodule