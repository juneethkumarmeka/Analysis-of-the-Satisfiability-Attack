module basic_1000_10000_1500_10_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
or U0 (N_0,In_380,In_370);
nand U1 (N_1,In_546,In_795);
nor U2 (N_2,In_488,In_661);
xor U3 (N_3,In_772,In_324);
nand U4 (N_4,In_239,In_178);
or U5 (N_5,In_723,In_111);
or U6 (N_6,In_789,In_508);
and U7 (N_7,In_297,In_229);
and U8 (N_8,In_707,In_873);
and U9 (N_9,In_947,In_462);
nor U10 (N_10,In_376,In_425);
xor U11 (N_11,In_694,In_448);
and U12 (N_12,In_305,In_361);
and U13 (N_13,In_104,In_470);
nand U14 (N_14,In_279,In_575);
xnor U15 (N_15,In_583,In_536);
nand U16 (N_16,In_405,In_533);
xor U17 (N_17,In_341,In_650);
xor U18 (N_18,In_82,In_952);
and U19 (N_19,In_609,In_327);
nand U20 (N_20,In_474,In_782);
xnor U21 (N_21,In_643,In_957);
nand U22 (N_22,In_90,In_917);
nand U23 (N_23,In_636,In_978);
or U24 (N_24,In_298,In_70);
nor U25 (N_25,In_129,In_803);
nor U26 (N_26,In_688,In_95);
or U27 (N_27,In_904,In_318);
nor U28 (N_28,In_792,In_778);
xnor U29 (N_29,In_377,In_754);
and U30 (N_30,In_215,In_103);
or U31 (N_31,In_530,In_240);
nor U32 (N_32,In_163,In_971);
nor U33 (N_33,In_303,In_704);
or U34 (N_34,In_612,In_191);
nand U35 (N_35,In_185,In_976);
nor U36 (N_36,In_892,In_895);
nor U37 (N_37,In_597,In_130);
xor U38 (N_38,In_582,In_729);
and U39 (N_39,In_220,In_137);
xor U40 (N_40,In_426,In_316);
xnor U41 (N_41,In_871,In_801);
nor U42 (N_42,In_202,In_598);
and U43 (N_43,In_925,In_738);
or U44 (N_44,In_617,In_8);
nor U45 (N_45,In_392,In_315);
or U46 (N_46,In_711,In_944);
and U47 (N_47,In_601,In_352);
xor U48 (N_48,In_192,In_715);
and U49 (N_49,In_347,In_172);
or U50 (N_50,In_161,In_436);
xnor U51 (N_51,In_152,In_808);
xnor U52 (N_52,In_517,In_767);
nand U53 (N_53,In_541,In_639);
or U54 (N_54,In_557,In_840);
nor U55 (N_55,In_248,In_684);
nor U56 (N_56,In_817,In_32);
and U57 (N_57,In_22,In_948);
xor U58 (N_58,In_275,In_653);
or U59 (N_59,In_584,In_168);
and U60 (N_60,In_972,In_753);
nor U61 (N_61,In_856,In_476);
xnor U62 (N_62,In_791,In_926);
xnor U63 (N_63,In_264,In_397);
and U64 (N_64,In_673,In_903);
nand U65 (N_65,In_350,In_120);
xnor U66 (N_66,In_837,In_362);
xor U67 (N_67,In_799,In_709);
nand U68 (N_68,In_491,In_263);
nand U69 (N_69,In_402,In_831);
nor U70 (N_70,In_809,In_632);
nor U71 (N_71,In_189,In_681);
nor U72 (N_72,In_683,In_400);
nor U73 (N_73,In_459,In_260);
and U74 (N_74,In_314,In_919);
and U75 (N_75,In_527,In_146);
nand U76 (N_76,In_339,In_992);
and U77 (N_77,In_826,In_678);
nor U78 (N_78,In_660,In_593);
or U79 (N_79,In_542,In_473);
nor U80 (N_80,In_885,In_469);
and U81 (N_81,In_43,In_76);
and U82 (N_82,In_969,In_812);
and U83 (N_83,In_44,In_828);
or U84 (N_84,In_993,In_276);
nand U85 (N_85,In_68,In_890);
and U86 (N_86,In_594,In_272);
xor U87 (N_87,In_351,In_519);
nand U88 (N_88,In_1,In_113);
nor U89 (N_89,In_946,In_563);
and U90 (N_90,In_65,In_943);
and U91 (N_91,In_87,In_468);
and U92 (N_92,In_337,In_197);
nand U93 (N_93,In_289,In_356);
or U94 (N_94,In_934,In_706);
nand U95 (N_95,In_209,In_463);
xnor U96 (N_96,In_40,In_449);
nand U97 (N_97,In_518,In_453);
nand U98 (N_98,In_291,In_242);
nand U99 (N_99,In_633,In_184);
xnor U100 (N_100,In_52,In_97);
xnor U101 (N_101,In_713,In_63);
xnor U102 (N_102,In_876,In_243);
and U103 (N_103,In_91,In_731);
or U104 (N_104,In_482,In_514);
nor U105 (N_105,In_929,In_857);
nand U106 (N_106,In_283,In_825);
and U107 (N_107,In_319,In_638);
nor U108 (N_108,In_222,In_11);
xnor U109 (N_109,In_427,In_702);
nor U110 (N_110,In_342,In_665);
nand U111 (N_111,In_133,In_317);
and U112 (N_112,In_496,In_198);
xor U113 (N_113,In_628,In_552);
xnor U114 (N_114,In_572,In_896);
xnor U115 (N_115,In_625,In_33);
and U116 (N_116,In_768,In_680);
nand U117 (N_117,In_15,In_48);
nor U118 (N_118,In_607,In_596);
xnor U119 (N_119,In_570,In_101);
xnor U120 (N_120,In_378,In_728);
or U121 (N_121,In_889,In_730);
and U122 (N_122,In_559,In_320);
nand U123 (N_123,In_72,In_391);
and U124 (N_124,In_849,In_699);
xor U125 (N_125,In_188,In_679);
xnor U126 (N_126,In_281,In_868);
nor U127 (N_127,In_949,In_382);
nand U128 (N_128,In_458,In_287);
and U129 (N_129,In_696,In_656);
or U130 (N_130,In_935,In_50);
nand U131 (N_131,In_770,In_909);
nand U132 (N_132,In_591,In_842);
nor U133 (N_133,In_428,In_150);
and U134 (N_134,In_211,In_126);
nor U135 (N_135,In_30,In_798);
or U136 (N_136,In_410,In_567);
or U137 (N_137,In_877,In_525);
nand U138 (N_138,In_424,In_196);
nand U139 (N_139,In_647,In_936);
nor U140 (N_140,In_164,In_813);
xnor U141 (N_141,In_16,In_784);
xnor U142 (N_142,In_829,In_659);
nor U143 (N_143,In_708,In_760);
and U144 (N_144,In_59,In_838);
xor U145 (N_145,In_853,In_937);
nor U146 (N_146,In_367,In_25);
and U147 (N_147,In_345,In_726);
and U148 (N_148,In_45,In_86);
nand U149 (N_149,In_590,In_471);
or U150 (N_150,In_785,In_771);
xor U151 (N_151,In_920,In_983);
xor U152 (N_152,In_35,In_657);
xor U153 (N_153,In_233,In_64);
and U154 (N_154,In_266,In_802);
nand U155 (N_155,In_495,In_10);
xnor U156 (N_156,In_938,In_695);
or U157 (N_157,In_506,In_334);
and U158 (N_158,In_26,In_611);
and U159 (N_159,In_225,In_592);
nand U160 (N_160,In_237,In_2);
xnor U161 (N_161,In_143,In_381);
xor U162 (N_162,In_295,In_252);
or U163 (N_163,In_452,In_939);
nand U164 (N_164,In_832,In_522);
and U165 (N_165,In_756,In_136);
and U166 (N_166,In_984,In_973);
or U167 (N_167,In_918,In_39);
or U168 (N_168,In_433,In_996);
and U169 (N_169,In_526,In_787);
nand U170 (N_170,In_986,In_388);
nor U171 (N_171,In_109,In_304);
or U172 (N_172,In_29,In_790);
nor U173 (N_173,In_308,In_814);
nand U174 (N_174,In_475,In_486);
nor U175 (N_175,In_132,In_589);
or U176 (N_176,In_182,In_535);
xor U177 (N_177,In_556,In_338);
xnor U178 (N_178,In_565,In_851);
nand U179 (N_179,In_941,In_258);
nor U180 (N_180,In_775,In_764);
or U181 (N_181,In_953,In_416);
or U182 (N_182,In_667,In_614);
or U183 (N_183,In_293,In_824);
and U184 (N_184,In_127,In_698);
nand U185 (N_185,In_968,In_821);
nand U186 (N_186,In_478,In_302);
or U187 (N_187,In_558,In_883);
xor U188 (N_188,In_578,In_863);
nand U189 (N_189,In_834,In_691);
xor U190 (N_190,In_415,In_716);
nor U191 (N_191,In_623,In_550);
nand U192 (N_192,In_204,In_443);
and U193 (N_193,In_531,In_321);
and U194 (N_194,In_9,In_499);
or U195 (N_195,In_447,In_385);
nor U196 (N_196,In_634,In_245);
and U197 (N_197,In_646,In_555);
xnor U198 (N_198,In_199,In_24);
nor U199 (N_199,In_477,In_67);
nor U200 (N_200,In_924,In_580);
xor U201 (N_201,In_460,In_125);
and U202 (N_202,In_364,In_265);
nor U203 (N_203,In_124,In_835);
and U204 (N_204,In_395,In_176);
xor U205 (N_205,In_256,In_654);
or U206 (N_206,In_902,In_502);
nor U207 (N_207,In_931,In_340);
xor U208 (N_208,In_515,In_740);
and U209 (N_209,In_92,In_102);
xnor U210 (N_210,In_0,In_271);
nor U211 (N_211,In_100,In_174);
nor U212 (N_212,In_855,In_457);
xnor U213 (N_213,In_774,In_898);
or U214 (N_214,In_620,In_674);
nand U215 (N_215,In_879,In_537);
and U216 (N_216,In_444,In_344);
and U217 (N_217,In_445,In_93);
or U218 (N_218,In_843,In_326);
nand U219 (N_219,In_144,In_867);
and U220 (N_220,In_155,In_74);
xnor U221 (N_221,In_399,In_933);
xnor U222 (N_222,In_777,In_762);
or U223 (N_223,In_897,In_874);
or U224 (N_224,In_306,In_77);
xnor U225 (N_225,In_165,In_655);
xor U226 (N_226,In_769,In_761);
nand U227 (N_227,In_6,In_332);
xor U228 (N_228,In_438,In_142);
nor U229 (N_229,In_55,In_744);
nand U230 (N_230,In_751,In_869);
nand U231 (N_231,In_247,In_195);
or U232 (N_232,In_203,In_216);
nand U233 (N_233,In_489,In_865);
or U234 (N_234,In_417,In_547);
nand U235 (N_235,In_963,In_18);
nand U236 (N_236,In_278,In_300);
xor U237 (N_237,In_131,In_480);
nor U238 (N_238,In_280,In_907);
nand U239 (N_239,In_269,In_836);
nand U240 (N_240,In_915,In_355);
or U241 (N_241,In_732,In_750);
xor U242 (N_242,In_14,In_114);
xor U243 (N_243,In_466,In_157);
nor U244 (N_244,In_505,In_520);
and U245 (N_245,In_69,In_467);
xnor U246 (N_246,In_85,In_299);
xnor U247 (N_247,In_571,In_500);
nand U248 (N_248,In_807,In_493);
nor U249 (N_249,In_183,In_159);
or U250 (N_250,In_490,In_781);
nand U251 (N_251,In_440,In_21);
or U252 (N_252,In_720,In_312);
xor U253 (N_253,In_138,In_4);
nand U254 (N_254,In_618,In_587);
xnor U255 (N_255,In_734,In_238);
nand U256 (N_256,In_872,In_637);
nor U257 (N_257,In_145,In_179);
xnor U258 (N_258,In_573,In_3);
or U259 (N_259,In_359,In_412);
and U260 (N_260,In_685,In_509);
or U261 (N_261,In_742,In_227);
nand U262 (N_262,In_284,In_207);
xor U263 (N_263,In_83,In_576);
xor U264 (N_264,In_219,In_249);
and U265 (N_265,In_210,In_394);
and U266 (N_266,In_561,In_37);
or U267 (N_267,In_322,In_375);
nor U268 (N_268,In_672,In_434);
nand U269 (N_269,In_881,In_441);
and U270 (N_270,In_579,In_759);
or U271 (N_271,In_135,In_613);
or U272 (N_272,In_747,In_651);
and U273 (N_273,In_66,In_58);
xnor U274 (N_274,In_257,In_577);
nand U275 (N_275,In_171,In_822);
nor U276 (N_276,In_122,In_940);
nor U277 (N_277,In_360,In_259);
xnor U278 (N_278,In_47,In_420);
and U279 (N_279,In_290,In_481);
nand U280 (N_280,In_73,In_282);
nand U281 (N_281,In_998,In_878);
and U282 (N_282,In_927,In_419);
xor U283 (N_283,In_528,In_534);
xnor U284 (N_284,In_980,In_286);
and U285 (N_285,In_970,In_267);
or U286 (N_286,In_999,In_664);
xor U287 (N_287,In_98,In_20);
or U288 (N_288,In_390,In_560);
xnor U289 (N_289,In_529,In_372);
nand U290 (N_290,In_36,In_989);
and U291 (N_291,In_516,In_689);
xor U292 (N_292,In_358,In_173);
nand U293 (N_293,In_630,In_860);
or U294 (N_294,In_200,In_603);
and U295 (N_295,In_408,In_7);
nand U296 (N_296,In_619,In_450);
or U297 (N_297,In_773,In_682);
nand U298 (N_298,In_693,In_421);
or U299 (N_299,In_544,In_733);
nor U300 (N_300,In_991,In_507);
nand U301 (N_301,In_662,In_187);
nand U302 (N_302,In_46,In_635);
nand U303 (N_303,In_78,In_626);
and U304 (N_304,In_884,In_810);
nor U305 (N_305,In_749,In_686);
nand U306 (N_306,In_62,In_437);
nand U307 (N_307,In_748,In_900);
and U308 (N_308,In_224,In_128);
and U309 (N_309,In_96,In_629);
nor U310 (N_310,In_294,In_366);
or U311 (N_311,In_956,In_253);
xor U312 (N_312,In_217,In_581);
xnor U313 (N_313,In_671,In_994);
xor U314 (N_314,In_140,In_251);
nor U315 (N_315,In_154,In_735);
or U316 (N_316,In_553,In_353);
nor U317 (N_317,In_640,In_270);
or U318 (N_318,In_990,In_309);
or U319 (N_319,In_811,In_886);
nor U320 (N_320,In_13,In_866);
xor U321 (N_321,In_610,In_621);
nor U322 (N_322,In_89,In_487);
or U323 (N_323,In_277,In_422);
xor U324 (N_324,In_465,In_725);
nor U325 (N_325,In_739,In_776);
nor U326 (N_326,In_12,In_472);
xor U327 (N_327,In_911,In_170);
and U328 (N_328,In_899,In_737);
nor U329 (N_329,In_690,In_223);
nor U330 (N_330,In_23,In_543);
nand U331 (N_331,In_110,In_942);
nor U332 (N_332,In_532,In_371);
and U333 (N_333,In_977,In_307);
or U334 (N_334,In_962,In_88);
nor U335 (N_335,In_585,In_84);
nor U336 (N_336,In_741,In_830);
or U337 (N_337,In_244,In_602);
nand U338 (N_338,In_846,In_285);
or U339 (N_339,In_719,In_374);
or U340 (N_340,In_631,In_357);
xor U341 (N_341,In_888,In_523);
nand U342 (N_342,In_997,In_461);
xor U343 (N_343,In_94,In_139);
or U344 (N_344,In_439,In_982);
xnor U345 (N_345,In_464,In_819);
or U346 (N_346,In_411,In_724);
xnor U347 (N_347,In_369,In_687);
nor U348 (N_348,In_368,In_615);
nor U349 (N_349,In_141,In_914);
nand U350 (N_350,In_49,In_894);
nand U351 (N_351,In_714,In_107);
nand U352 (N_352,In_147,In_151);
xor U353 (N_353,In_804,In_669);
or U354 (N_354,In_823,In_880);
or U355 (N_355,In_336,In_166);
nor U356 (N_356,In_668,In_60);
nor U357 (N_357,In_181,In_346);
nor U358 (N_358,In_622,In_503);
nand U359 (N_359,In_670,In_847);
and U360 (N_360,In_692,In_213);
nand U361 (N_361,In_524,In_967);
and U362 (N_362,In_479,In_384);
and U363 (N_363,In_882,In_649);
xnor U364 (N_364,In_54,In_988);
or U365 (N_365,In_42,In_456);
nand U366 (N_366,In_348,In_906);
or U367 (N_367,In_588,In_288);
nand U368 (N_368,In_512,In_180);
or U369 (N_369,In_232,In_710);
and U370 (N_370,In_61,In_966);
nand U371 (N_371,In_833,In_859);
or U372 (N_372,In_118,In_964);
and U373 (N_373,In_794,In_254);
xor U374 (N_374,In_862,In_407);
xor U375 (N_375,In_349,In_912);
nor U376 (N_376,In_175,In_17);
nor U377 (N_377,In_301,In_910);
xor U378 (N_378,In_423,In_117);
nand U379 (N_379,In_404,In_800);
and U380 (N_380,In_162,In_945);
and U381 (N_381,In_454,In_53);
nor U382 (N_382,In_406,In_605);
and U383 (N_383,In_212,In_158);
nor U384 (N_384,In_975,In_648);
and U385 (N_385,In_595,In_160);
and U386 (N_386,In_844,In_743);
nand U387 (N_387,In_75,In_123);
or U388 (N_388,In_105,In_701);
or U389 (N_389,In_343,In_205);
and U390 (N_390,In_226,In_758);
xnor U391 (N_391,In_383,In_870);
nand U392 (N_392,In_922,In_841);
xnor U393 (N_393,In_951,In_446);
nand U394 (N_394,In_193,In_373);
and U395 (N_395,In_389,In_177);
or U396 (N_396,In_494,In_845);
xnor U397 (N_397,In_854,In_186);
or U398 (N_398,In_148,In_921);
and U399 (N_399,In_923,In_783);
xnor U400 (N_400,In_228,In_169);
or U401 (N_401,In_99,In_608);
nor U402 (N_402,In_797,In_566);
and U403 (N_403,In_116,In_231);
nand U404 (N_404,In_905,In_235);
and U405 (N_405,In_766,In_913);
nor U406 (N_406,In_396,In_752);
xor U407 (N_407,In_330,In_958);
xnor U408 (N_408,In_112,In_727);
nand U409 (N_409,In_57,In_658);
or U410 (N_410,In_354,In_663);
or U411 (N_411,In_786,In_757);
nor U412 (N_412,In_335,In_928);
or U413 (N_413,In_379,In_538);
or U414 (N_414,In_393,In_431);
nor U415 (N_415,In_31,In_413);
nand U416 (N_416,In_108,In_916);
xor U417 (N_417,In_214,In_642);
nor U418 (N_418,In_403,In_562);
and U419 (N_419,In_763,In_484);
or U420 (N_420,In_119,In_292);
nor U421 (N_421,In_483,In_959);
or U422 (N_422,In_246,In_765);
or U423 (N_423,In_624,In_549);
nor U424 (N_424,In_788,In_387);
nand U425 (N_425,In_296,In_310);
or U426 (N_426,In_755,In_329);
or U427 (N_427,In_208,In_818);
and U428 (N_428,In_569,In_331);
and U429 (N_429,In_156,In_262);
and U430 (N_430,In_796,In_194);
xnor U431 (N_431,In_28,In_234);
or U432 (N_432,In_5,In_600);
and U433 (N_433,In_599,In_930);
nor U434 (N_434,In_401,In_365);
xor U435 (N_435,In_981,In_606);
and U436 (N_436,In_793,In_51);
xor U437 (N_437,In_539,In_652);
and U438 (N_438,In_604,In_492);
or U439 (N_439,In_950,In_697);
or U440 (N_440,In_167,In_513);
and U441 (N_441,In_442,In_861);
nand U442 (N_442,In_722,In_34);
nor U443 (N_443,In_115,In_627);
nand U444 (N_444,In_409,In_134);
nand U445 (N_445,In_736,In_250);
nor U446 (N_446,In_328,In_79);
xnor U447 (N_447,In_398,In_891);
nand U448 (N_448,In_979,In_932);
and U449 (N_449,In_149,In_908);
or U450 (N_450,In_574,In_551);
nor U451 (N_451,In_816,In_893);
xor U452 (N_452,In_435,In_548);
nand U453 (N_453,In_954,In_779);
or U454 (N_454,In_564,In_641);
xor U455 (N_455,In_268,In_273);
or U456 (N_456,In_815,In_858);
nor U457 (N_457,In_718,In_255);
xor U458 (N_458,In_38,In_218);
xor U459 (N_459,In_41,In_121);
xnor U460 (N_460,In_504,In_206);
nand U461 (N_461,In_230,In_80);
or U462 (N_462,In_705,In_666);
xor U463 (N_463,In_676,In_864);
nand U464 (N_464,In_554,In_703);
or U465 (N_465,In_451,In_780);
or U466 (N_466,In_429,In_221);
nand U467 (N_467,In_521,In_677);
nand U468 (N_468,In_311,In_901);
nor U469 (N_469,In_827,In_511);
nand U470 (N_470,In_700,In_850);
or U471 (N_471,In_995,In_510);
nor U472 (N_472,In_241,In_839);
xor U473 (N_473,In_568,In_414);
nand U474 (N_474,In_323,In_806);
and U475 (N_475,In_201,In_586);
or U476 (N_476,In_497,In_545);
nand U477 (N_477,In_745,In_418);
nor U478 (N_478,In_153,In_485);
or U479 (N_479,In_106,In_325);
nand U480 (N_480,In_852,In_960);
nor U481 (N_481,In_887,In_805);
nand U482 (N_482,In_363,In_616);
and U483 (N_483,In_190,In_236);
or U484 (N_484,In_19,In_746);
or U485 (N_485,In_386,In_645);
nand U486 (N_486,In_81,In_501);
or U487 (N_487,In_432,In_875);
nand U488 (N_488,In_540,In_313);
nand U489 (N_489,In_261,In_71);
nor U490 (N_490,In_712,In_56);
nor U491 (N_491,In_985,In_717);
or U492 (N_492,In_820,In_965);
or U493 (N_493,In_675,In_27);
and U494 (N_494,In_974,In_498);
or U495 (N_495,In_644,In_274);
and U496 (N_496,In_955,In_961);
nand U497 (N_497,In_721,In_848);
xor U498 (N_498,In_430,In_987);
or U499 (N_499,In_333,In_455);
and U500 (N_500,In_78,In_212);
or U501 (N_501,In_800,In_439);
nor U502 (N_502,In_766,In_452);
nand U503 (N_503,In_918,In_666);
xor U504 (N_504,In_349,In_538);
or U505 (N_505,In_275,In_560);
xnor U506 (N_506,In_493,In_797);
xnor U507 (N_507,In_207,In_30);
nor U508 (N_508,In_129,In_943);
or U509 (N_509,In_36,In_51);
xnor U510 (N_510,In_701,In_30);
or U511 (N_511,In_892,In_705);
or U512 (N_512,In_336,In_797);
nor U513 (N_513,In_54,In_958);
and U514 (N_514,In_418,In_568);
or U515 (N_515,In_805,In_39);
xor U516 (N_516,In_773,In_883);
or U517 (N_517,In_287,In_181);
xnor U518 (N_518,In_512,In_1);
nor U519 (N_519,In_292,In_255);
nand U520 (N_520,In_476,In_805);
nor U521 (N_521,In_265,In_788);
nor U522 (N_522,In_159,In_72);
nor U523 (N_523,In_983,In_945);
or U524 (N_524,In_699,In_114);
nand U525 (N_525,In_474,In_288);
or U526 (N_526,In_587,In_887);
nand U527 (N_527,In_572,In_324);
xnor U528 (N_528,In_698,In_521);
nor U529 (N_529,In_619,In_775);
nand U530 (N_530,In_915,In_294);
nor U531 (N_531,In_82,In_265);
and U532 (N_532,In_973,In_966);
nor U533 (N_533,In_263,In_305);
and U534 (N_534,In_724,In_750);
xnor U535 (N_535,In_554,In_663);
xor U536 (N_536,In_691,In_115);
or U537 (N_537,In_430,In_15);
xnor U538 (N_538,In_757,In_232);
xnor U539 (N_539,In_450,In_340);
xnor U540 (N_540,In_112,In_801);
nor U541 (N_541,In_279,In_18);
or U542 (N_542,In_131,In_63);
and U543 (N_543,In_70,In_518);
or U544 (N_544,In_558,In_730);
or U545 (N_545,In_951,In_512);
or U546 (N_546,In_504,In_786);
or U547 (N_547,In_781,In_880);
or U548 (N_548,In_937,In_419);
nor U549 (N_549,In_593,In_596);
nand U550 (N_550,In_236,In_979);
nand U551 (N_551,In_477,In_221);
and U552 (N_552,In_358,In_564);
nand U553 (N_553,In_156,In_539);
and U554 (N_554,In_550,In_996);
or U555 (N_555,In_320,In_868);
xor U556 (N_556,In_772,In_132);
nand U557 (N_557,In_360,In_438);
or U558 (N_558,In_0,In_725);
nand U559 (N_559,In_80,In_654);
or U560 (N_560,In_502,In_649);
xnor U561 (N_561,In_988,In_223);
nor U562 (N_562,In_88,In_559);
or U563 (N_563,In_985,In_100);
xor U564 (N_564,In_518,In_367);
or U565 (N_565,In_762,In_823);
or U566 (N_566,In_954,In_443);
nor U567 (N_567,In_991,In_665);
or U568 (N_568,In_539,In_305);
and U569 (N_569,In_257,In_366);
nand U570 (N_570,In_442,In_933);
and U571 (N_571,In_424,In_805);
and U572 (N_572,In_788,In_771);
nor U573 (N_573,In_388,In_602);
and U574 (N_574,In_609,In_525);
and U575 (N_575,In_892,In_707);
and U576 (N_576,In_983,In_429);
or U577 (N_577,In_919,In_774);
nand U578 (N_578,In_570,In_203);
or U579 (N_579,In_940,In_778);
and U580 (N_580,In_152,In_730);
and U581 (N_581,In_887,In_616);
nand U582 (N_582,In_636,In_885);
and U583 (N_583,In_911,In_984);
and U584 (N_584,In_564,In_506);
and U585 (N_585,In_238,In_766);
and U586 (N_586,In_101,In_30);
xnor U587 (N_587,In_584,In_3);
xnor U588 (N_588,In_813,In_682);
nand U589 (N_589,In_468,In_810);
xnor U590 (N_590,In_723,In_879);
nor U591 (N_591,In_781,In_553);
xor U592 (N_592,In_361,In_464);
and U593 (N_593,In_120,In_950);
or U594 (N_594,In_559,In_205);
or U595 (N_595,In_219,In_188);
or U596 (N_596,In_877,In_405);
nand U597 (N_597,In_373,In_598);
nor U598 (N_598,In_653,In_726);
nor U599 (N_599,In_470,In_894);
and U600 (N_600,In_11,In_676);
nand U601 (N_601,In_567,In_346);
nand U602 (N_602,In_401,In_347);
and U603 (N_603,In_808,In_786);
or U604 (N_604,In_571,In_116);
or U605 (N_605,In_835,In_66);
or U606 (N_606,In_324,In_844);
and U607 (N_607,In_128,In_27);
xor U608 (N_608,In_59,In_609);
or U609 (N_609,In_322,In_636);
nand U610 (N_610,In_850,In_155);
nand U611 (N_611,In_570,In_781);
nor U612 (N_612,In_457,In_806);
or U613 (N_613,In_785,In_680);
nand U614 (N_614,In_312,In_22);
xor U615 (N_615,In_833,In_381);
xor U616 (N_616,In_265,In_535);
or U617 (N_617,In_93,In_295);
or U618 (N_618,In_802,In_875);
or U619 (N_619,In_82,In_53);
and U620 (N_620,In_262,In_566);
or U621 (N_621,In_668,In_747);
nand U622 (N_622,In_308,In_550);
xnor U623 (N_623,In_406,In_891);
nor U624 (N_624,In_392,In_575);
or U625 (N_625,In_261,In_892);
xor U626 (N_626,In_1,In_703);
nor U627 (N_627,In_580,In_827);
nor U628 (N_628,In_82,In_383);
xnor U629 (N_629,In_660,In_511);
nor U630 (N_630,In_370,In_363);
nor U631 (N_631,In_417,In_339);
xnor U632 (N_632,In_71,In_926);
nor U633 (N_633,In_134,In_525);
and U634 (N_634,In_534,In_588);
nand U635 (N_635,In_495,In_978);
and U636 (N_636,In_915,In_631);
nand U637 (N_637,In_998,In_425);
nand U638 (N_638,In_864,In_657);
xnor U639 (N_639,In_486,In_590);
xor U640 (N_640,In_970,In_747);
xor U641 (N_641,In_922,In_843);
and U642 (N_642,In_124,In_235);
nor U643 (N_643,In_125,In_536);
and U644 (N_644,In_384,In_574);
xor U645 (N_645,In_302,In_965);
or U646 (N_646,In_958,In_654);
or U647 (N_647,In_718,In_614);
and U648 (N_648,In_930,In_183);
xor U649 (N_649,In_47,In_2);
nor U650 (N_650,In_113,In_29);
or U651 (N_651,In_417,In_513);
and U652 (N_652,In_401,In_21);
xor U653 (N_653,In_2,In_551);
and U654 (N_654,In_553,In_225);
xor U655 (N_655,In_860,In_46);
xor U656 (N_656,In_867,In_367);
nor U657 (N_657,In_676,In_489);
xnor U658 (N_658,In_596,In_24);
and U659 (N_659,In_256,In_705);
or U660 (N_660,In_535,In_581);
or U661 (N_661,In_672,In_69);
nand U662 (N_662,In_471,In_979);
or U663 (N_663,In_386,In_908);
nand U664 (N_664,In_825,In_406);
xor U665 (N_665,In_465,In_918);
and U666 (N_666,In_424,In_97);
and U667 (N_667,In_398,In_82);
nor U668 (N_668,In_123,In_610);
nor U669 (N_669,In_682,In_757);
nand U670 (N_670,In_66,In_505);
nand U671 (N_671,In_169,In_651);
nand U672 (N_672,In_676,In_964);
xor U673 (N_673,In_382,In_65);
nand U674 (N_674,In_25,In_889);
and U675 (N_675,In_656,In_307);
nand U676 (N_676,In_969,In_731);
nand U677 (N_677,In_12,In_486);
and U678 (N_678,In_314,In_610);
and U679 (N_679,In_774,In_610);
xor U680 (N_680,In_376,In_358);
nand U681 (N_681,In_571,In_79);
nand U682 (N_682,In_54,In_370);
nand U683 (N_683,In_831,In_124);
and U684 (N_684,In_500,In_445);
and U685 (N_685,In_975,In_947);
nor U686 (N_686,In_124,In_41);
nor U687 (N_687,In_930,In_812);
or U688 (N_688,In_317,In_549);
nor U689 (N_689,In_626,In_781);
xor U690 (N_690,In_284,In_150);
nor U691 (N_691,In_460,In_684);
or U692 (N_692,In_226,In_830);
nor U693 (N_693,In_650,In_598);
nor U694 (N_694,In_264,In_601);
nand U695 (N_695,In_545,In_250);
and U696 (N_696,In_724,In_468);
xor U697 (N_697,In_897,In_995);
nor U698 (N_698,In_998,In_675);
xnor U699 (N_699,In_257,In_543);
and U700 (N_700,In_506,In_218);
and U701 (N_701,In_631,In_730);
and U702 (N_702,In_365,In_154);
xnor U703 (N_703,In_296,In_109);
nand U704 (N_704,In_219,In_555);
nor U705 (N_705,In_854,In_48);
and U706 (N_706,In_958,In_440);
nor U707 (N_707,In_50,In_586);
nor U708 (N_708,In_318,In_397);
nand U709 (N_709,In_200,In_974);
or U710 (N_710,In_684,In_672);
xor U711 (N_711,In_323,In_965);
or U712 (N_712,In_581,In_47);
and U713 (N_713,In_679,In_257);
and U714 (N_714,In_233,In_706);
nor U715 (N_715,In_6,In_708);
and U716 (N_716,In_839,In_240);
or U717 (N_717,In_47,In_752);
and U718 (N_718,In_565,In_420);
nand U719 (N_719,In_486,In_491);
and U720 (N_720,In_504,In_703);
or U721 (N_721,In_529,In_541);
nand U722 (N_722,In_127,In_44);
nor U723 (N_723,In_591,In_994);
xnor U724 (N_724,In_164,In_260);
nor U725 (N_725,In_879,In_860);
nand U726 (N_726,In_713,In_332);
and U727 (N_727,In_937,In_602);
nor U728 (N_728,In_87,In_959);
xnor U729 (N_729,In_388,In_368);
nand U730 (N_730,In_589,In_906);
or U731 (N_731,In_948,In_136);
and U732 (N_732,In_614,In_3);
nor U733 (N_733,In_728,In_12);
and U734 (N_734,In_965,In_141);
nand U735 (N_735,In_661,In_518);
and U736 (N_736,In_196,In_172);
xnor U737 (N_737,In_683,In_702);
or U738 (N_738,In_778,In_448);
or U739 (N_739,In_822,In_48);
xnor U740 (N_740,In_746,In_42);
or U741 (N_741,In_397,In_9);
and U742 (N_742,In_708,In_29);
xnor U743 (N_743,In_691,In_848);
nor U744 (N_744,In_657,In_347);
and U745 (N_745,In_979,In_771);
xnor U746 (N_746,In_22,In_722);
nor U747 (N_747,In_160,In_71);
or U748 (N_748,In_217,In_451);
nand U749 (N_749,In_386,In_227);
and U750 (N_750,In_566,In_330);
xnor U751 (N_751,In_430,In_976);
nand U752 (N_752,In_821,In_266);
xor U753 (N_753,In_251,In_143);
nand U754 (N_754,In_206,In_908);
and U755 (N_755,In_193,In_615);
nand U756 (N_756,In_293,In_718);
and U757 (N_757,In_735,In_848);
and U758 (N_758,In_559,In_380);
xnor U759 (N_759,In_673,In_335);
nand U760 (N_760,In_47,In_837);
nand U761 (N_761,In_178,In_626);
nor U762 (N_762,In_731,In_781);
nor U763 (N_763,In_135,In_409);
xnor U764 (N_764,In_667,In_530);
and U765 (N_765,In_32,In_106);
and U766 (N_766,In_165,In_430);
nand U767 (N_767,In_614,In_441);
nor U768 (N_768,In_37,In_630);
xor U769 (N_769,In_247,In_3);
nand U770 (N_770,In_373,In_79);
nor U771 (N_771,In_639,In_790);
nor U772 (N_772,In_606,In_371);
nor U773 (N_773,In_843,In_297);
and U774 (N_774,In_282,In_856);
and U775 (N_775,In_679,In_544);
or U776 (N_776,In_917,In_968);
xnor U777 (N_777,In_442,In_430);
xor U778 (N_778,In_734,In_272);
xor U779 (N_779,In_348,In_200);
or U780 (N_780,In_177,In_828);
xnor U781 (N_781,In_469,In_508);
xnor U782 (N_782,In_621,In_364);
or U783 (N_783,In_462,In_51);
xor U784 (N_784,In_125,In_875);
nor U785 (N_785,In_923,In_56);
nor U786 (N_786,In_535,In_324);
or U787 (N_787,In_704,In_938);
and U788 (N_788,In_152,In_435);
xor U789 (N_789,In_994,In_421);
nor U790 (N_790,In_378,In_590);
or U791 (N_791,In_407,In_975);
nand U792 (N_792,In_43,In_733);
xnor U793 (N_793,In_622,In_479);
nand U794 (N_794,In_661,In_84);
nor U795 (N_795,In_75,In_911);
xor U796 (N_796,In_56,In_473);
or U797 (N_797,In_366,In_718);
nor U798 (N_798,In_466,In_256);
and U799 (N_799,In_223,In_851);
nor U800 (N_800,In_792,In_215);
nand U801 (N_801,In_638,In_791);
nand U802 (N_802,In_16,In_665);
nand U803 (N_803,In_277,In_28);
xor U804 (N_804,In_769,In_516);
nand U805 (N_805,In_544,In_273);
or U806 (N_806,In_549,In_49);
nor U807 (N_807,In_562,In_578);
and U808 (N_808,In_969,In_682);
or U809 (N_809,In_799,In_345);
nor U810 (N_810,In_130,In_548);
and U811 (N_811,In_553,In_179);
nor U812 (N_812,In_605,In_203);
or U813 (N_813,In_106,In_531);
nand U814 (N_814,In_794,In_681);
or U815 (N_815,In_254,In_723);
and U816 (N_816,In_783,In_650);
nor U817 (N_817,In_220,In_655);
xor U818 (N_818,In_75,In_747);
nor U819 (N_819,In_791,In_682);
and U820 (N_820,In_764,In_914);
and U821 (N_821,In_877,In_819);
and U822 (N_822,In_854,In_931);
xnor U823 (N_823,In_901,In_396);
or U824 (N_824,In_390,In_325);
nor U825 (N_825,In_11,In_15);
nor U826 (N_826,In_933,In_228);
nor U827 (N_827,In_215,In_824);
or U828 (N_828,In_962,In_946);
xor U829 (N_829,In_794,In_140);
and U830 (N_830,In_725,In_875);
or U831 (N_831,In_35,In_82);
nor U832 (N_832,In_510,In_588);
and U833 (N_833,In_980,In_695);
or U834 (N_834,In_86,In_908);
nor U835 (N_835,In_560,In_451);
xnor U836 (N_836,In_961,In_782);
or U837 (N_837,In_796,In_116);
nor U838 (N_838,In_749,In_794);
xor U839 (N_839,In_898,In_56);
and U840 (N_840,In_522,In_224);
nor U841 (N_841,In_504,In_701);
xor U842 (N_842,In_507,In_405);
and U843 (N_843,In_475,In_97);
and U844 (N_844,In_292,In_401);
nor U845 (N_845,In_859,In_837);
or U846 (N_846,In_680,In_534);
or U847 (N_847,In_91,In_44);
or U848 (N_848,In_204,In_905);
nand U849 (N_849,In_610,In_442);
and U850 (N_850,In_500,In_351);
nor U851 (N_851,In_155,In_905);
nor U852 (N_852,In_457,In_598);
nand U853 (N_853,In_365,In_580);
nand U854 (N_854,In_35,In_436);
nand U855 (N_855,In_459,In_417);
or U856 (N_856,In_463,In_831);
and U857 (N_857,In_105,In_435);
or U858 (N_858,In_783,In_526);
or U859 (N_859,In_644,In_320);
xnor U860 (N_860,In_741,In_731);
nand U861 (N_861,In_558,In_444);
or U862 (N_862,In_920,In_222);
or U863 (N_863,In_342,In_227);
or U864 (N_864,In_330,In_793);
and U865 (N_865,In_845,In_187);
xnor U866 (N_866,In_930,In_802);
nor U867 (N_867,In_293,In_72);
nand U868 (N_868,In_238,In_331);
nand U869 (N_869,In_311,In_319);
and U870 (N_870,In_441,In_899);
or U871 (N_871,In_152,In_918);
and U872 (N_872,In_864,In_234);
and U873 (N_873,In_220,In_894);
and U874 (N_874,In_4,In_888);
or U875 (N_875,In_713,In_136);
nor U876 (N_876,In_91,In_237);
and U877 (N_877,In_575,In_636);
and U878 (N_878,In_155,In_108);
and U879 (N_879,In_222,In_135);
nor U880 (N_880,In_747,In_194);
nor U881 (N_881,In_727,In_375);
nand U882 (N_882,In_317,In_659);
xor U883 (N_883,In_431,In_275);
and U884 (N_884,In_561,In_569);
or U885 (N_885,In_88,In_647);
nand U886 (N_886,In_495,In_725);
nand U887 (N_887,In_282,In_833);
or U888 (N_888,In_790,In_526);
or U889 (N_889,In_577,In_876);
and U890 (N_890,In_979,In_632);
or U891 (N_891,In_457,In_28);
xor U892 (N_892,In_883,In_412);
nor U893 (N_893,In_337,In_277);
or U894 (N_894,In_289,In_260);
or U895 (N_895,In_304,In_298);
nor U896 (N_896,In_614,In_279);
and U897 (N_897,In_908,In_122);
xnor U898 (N_898,In_919,In_857);
nand U899 (N_899,In_493,In_435);
xor U900 (N_900,In_47,In_575);
nand U901 (N_901,In_498,In_9);
nand U902 (N_902,In_622,In_160);
and U903 (N_903,In_717,In_592);
nor U904 (N_904,In_627,In_512);
or U905 (N_905,In_883,In_462);
nor U906 (N_906,In_497,In_270);
nor U907 (N_907,In_918,In_470);
or U908 (N_908,In_761,In_785);
nand U909 (N_909,In_492,In_564);
and U910 (N_910,In_422,In_841);
nand U911 (N_911,In_912,In_872);
xnor U912 (N_912,In_77,In_510);
nor U913 (N_913,In_849,In_702);
xor U914 (N_914,In_370,In_122);
nor U915 (N_915,In_971,In_705);
or U916 (N_916,In_545,In_399);
xor U917 (N_917,In_24,In_768);
or U918 (N_918,In_620,In_819);
nand U919 (N_919,In_708,In_917);
nand U920 (N_920,In_765,In_822);
or U921 (N_921,In_560,In_909);
nand U922 (N_922,In_935,In_215);
xnor U923 (N_923,In_329,In_215);
xor U924 (N_924,In_112,In_892);
nand U925 (N_925,In_139,In_840);
or U926 (N_926,In_765,In_306);
nor U927 (N_927,In_519,In_37);
and U928 (N_928,In_562,In_458);
xor U929 (N_929,In_895,In_801);
or U930 (N_930,In_580,In_679);
nor U931 (N_931,In_974,In_46);
or U932 (N_932,In_466,In_199);
or U933 (N_933,In_873,In_66);
nand U934 (N_934,In_449,In_28);
nand U935 (N_935,In_523,In_884);
or U936 (N_936,In_505,In_901);
or U937 (N_937,In_272,In_860);
nand U938 (N_938,In_113,In_761);
xnor U939 (N_939,In_856,In_369);
xnor U940 (N_940,In_267,In_533);
nor U941 (N_941,In_191,In_269);
or U942 (N_942,In_764,In_88);
nand U943 (N_943,In_432,In_405);
nand U944 (N_944,In_818,In_557);
and U945 (N_945,In_594,In_810);
and U946 (N_946,In_84,In_253);
and U947 (N_947,In_347,In_219);
nand U948 (N_948,In_224,In_183);
nand U949 (N_949,In_775,In_251);
xnor U950 (N_950,In_950,In_125);
nor U951 (N_951,In_943,In_47);
nand U952 (N_952,In_588,In_284);
xor U953 (N_953,In_705,In_942);
or U954 (N_954,In_559,In_387);
nor U955 (N_955,In_952,In_80);
or U956 (N_956,In_139,In_911);
and U957 (N_957,In_426,In_763);
nand U958 (N_958,In_999,In_273);
xnor U959 (N_959,In_722,In_612);
nor U960 (N_960,In_298,In_875);
nand U961 (N_961,In_714,In_407);
and U962 (N_962,In_626,In_943);
and U963 (N_963,In_667,In_924);
and U964 (N_964,In_842,In_683);
nor U965 (N_965,In_854,In_133);
nor U966 (N_966,In_941,In_953);
nor U967 (N_967,In_476,In_785);
nand U968 (N_968,In_148,In_421);
xnor U969 (N_969,In_35,In_804);
nor U970 (N_970,In_123,In_347);
nor U971 (N_971,In_776,In_793);
nor U972 (N_972,In_630,In_730);
or U973 (N_973,In_625,In_891);
or U974 (N_974,In_546,In_769);
and U975 (N_975,In_5,In_908);
xnor U976 (N_976,In_512,In_214);
or U977 (N_977,In_139,In_864);
or U978 (N_978,In_323,In_353);
nor U979 (N_979,In_392,In_797);
and U980 (N_980,In_737,In_716);
nand U981 (N_981,In_228,In_757);
or U982 (N_982,In_538,In_171);
nor U983 (N_983,In_463,In_147);
and U984 (N_984,In_309,In_138);
and U985 (N_985,In_490,In_136);
xor U986 (N_986,In_691,In_36);
or U987 (N_987,In_475,In_854);
nand U988 (N_988,In_493,In_554);
nand U989 (N_989,In_583,In_87);
nand U990 (N_990,In_847,In_962);
nand U991 (N_991,In_908,In_949);
xor U992 (N_992,In_775,In_763);
nand U993 (N_993,In_23,In_814);
nor U994 (N_994,In_530,In_792);
xor U995 (N_995,In_344,In_38);
or U996 (N_996,In_534,In_479);
xnor U997 (N_997,In_978,In_226);
and U998 (N_998,In_773,In_37);
or U999 (N_999,In_736,In_289);
xnor U1000 (N_1000,N_70,N_424);
or U1001 (N_1001,N_733,N_590);
xnor U1002 (N_1002,N_444,N_218);
and U1003 (N_1003,N_32,N_489);
nor U1004 (N_1004,N_982,N_958);
nand U1005 (N_1005,N_41,N_110);
nor U1006 (N_1006,N_978,N_684);
nor U1007 (N_1007,N_674,N_563);
nor U1008 (N_1008,N_395,N_726);
or U1009 (N_1009,N_435,N_367);
nor U1010 (N_1010,N_48,N_589);
nand U1011 (N_1011,N_297,N_178);
xor U1012 (N_1012,N_704,N_644);
nor U1013 (N_1013,N_266,N_541);
nand U1014 (N_1014,N_856,N_912);
nor U1015 (N_1015,N_406,N_353);
xor U1016 (N_1016,N_467,N_604);
nor U1017 (N_1017,N_224,N_165);
xnor U1018 (N_1018,N_250,N_522);
xnor U1019 (N_1019,N_942,N_378);
nand U1020 (N_1020,N_261,N_865);
and U1021 (N_1021,N_331,N_140);
xnor U1022 (N_1022,N_791,N_764);
nand U1023 (N_1023,N_623,N_918);
xnor U1024 (N_1024,N_386,N_330);
and U1025 (N_1025,N_88,N_789);
nand U1026 (N_1026,N_356,N_818);
and U1027 (N_1027,N_280,N_102);
xnor U1028 (N_1028,N_638,N_392);
and U1029 (N_1029,N_549,N_333);
nand U1030 (N_1030,N_785,N_78);
nand U1031 (N_1031,N_230,N_658);
nor U1032 (N_1032,N_470,N_962);
and U1033 (N_1033,N_432,N_566);
and U1034 (N_1034,N_204,N_894);
or U1035 (N_1035,N_570,N_95);
and U1036 (N_1036,N_838,N_167);
nand U1037 (N_1037,N_234,N_253);
or U1038 (N_1038,N_402,N_488);
nor U1039 (N_1039,N_870,N_162);
nor U1040 (N_1040,N_502,N_538);
nand U1041 (N_1041,N_646,N_968);
nand U1042 (N_1042,N_565,N_405);
or U1043 (N_1043,N_672,N_582);
xor U1044 (N_1044,N_927,N_74);
or U1045 (N_1045,N_871,N_873);
and U1046 (N_1046,N_398,N_242);
nor U1047 (N_1047,N_374,N_564);
or U1048 (N_1048,N_525,N_967);
or U1049 (N_1049,N_686,N_259);
xnor U1050 (N_1050,N_680,N_437);
nand U1051 (N_1051,N_106,N_782);
nor U1052 (N_1052,N_143,N_752);
and U1053 (N_1053,N_372,N_248);
xor U1054 (N_1054,N_159,N_660);
nor U1055 (N_1055,N_338,N_177);
and U1056 (N_1056,N_120,N_6);
nor U1057 (N_1057,N_901,N_370);
and U1058 (N_1058,N_152,N_529);
nand U1059 (N_1059,N_805,N_238);
and U1060 (N_1060,N_27,N_548);
and U1061 (N_1061,N_233,N_126);
nand U1062 (N_1062,N_622,N_493);
and U1063 (N_1063,N_343,N_896);
xor U1064 (N_1064,N_699,N_216);
or U1065 (N_1065,N_592,N_54);
xnor U1066 (N_1066,N_568,N_419);
and U1067 (N_1067,N_947,N_948);
and U1068 (N_1068,N_768,N_943);
or U1069 (N_1069,N_933,N_545);
xor U1070 (N_1070,N_503,N_546);
or U1071 (N_1071,N_677,N_830);
and U1072 (N_1072,N_624,N_670);
xor U1073 (N_1073,N_202,N_841);
nand U1074 (N_1074,N_137,N_852);
nand U1075 (N_1075,N_985,N_595);
xnor U1076 (N_1076,N_891,N_341);
and U1077 (N_1077,N_829,N_758);
nor U1078 (N_1078,N_929,N_303);
nand U1079 (N_1079,N_937,N_39);
xor U1080 (N_1080,N_664,N_468);
xnor U1081 (N_1081,N_851,N_125);
or U1082 (N_1082,N_278,N_635);
xnor U1083 (N_1083,N_669,N_104);
nand U1084 (N_1084,N_240,N_119);
or U1085 (N_1085,N_799,N_360);
and U1086 (N_1086,N_505,N_802);
or U1087 (N_1087,N_875,N_209);
or U1088 (N_1088,N_792,N_25);
or U1089 (N_1089,N_410,N_394);
or U1090 (N_1090,N_915,N_243);
xnor U1091 (N_1091,N_507,N_232);
or U1092 (N_1092,N_399,N_313);
nor U1093 (N_1093,N_897,N_715);
and U1094 (N_1094,N_600,N_151);
and U1095 (N_1095,N_889,N_597);
and U1096 (N_1096,N_426,N_581);
or U1097 (N_1097,N_161,N_56);
nand U1098 (N_1098,N_314,N_214);
and U1099 (N_1099,N_690,N_652);
nand U1100 (N_1100,N_134,N_815);
and U1101 (N_1101,N_182,N_301);
nand U1102 (N_1102,N_626,N_509);
or U1103 (N_1103,N_979,N_989);
nor U1104 (N_1104,N_422,N_984);
or U1105 (N_1105,N_450,N_171);
and U1106 (N_1106,N_701,N_255);
xnor U1107 (N_1107,N_878,N_212);
and U1108 (N_1108,N_607,N_499);
or U1109 (N_1109,N_369,N_75);
nand U1110 (N_1110,N_380,N_970);
and U1111 (N_1111,N_874,N_459);
nand U1112 (N_1112,N_904,N_425);
nand U1113 (N_1113,N_659,N_973);
xnor U1114 (N_1114,N_971,N_390);
nand U1115 (N_1115,N_521,N_895);
xnor U1116 (N_1116,N_481,N_630);
nor U1117 (N_1117,N_634,N_431);
nand U1118 (N_1118,N_666,N_832);
or U1119 (N_1119,N_364,N_265);
xor U1120 (N_1120,N_544,N_37);
or U1121 (N_1121,N_717,N_617);
or U1122 (N_1122,N_2,N_835);
and U1123 (N_1123,N_17,N_418);
nor U1124 (N_1124,N_58,N_408);
xnor U1125 (N_1125,N_256,N_316);
nor U1126 (N_1126,N_696,N_480);
nor U1127 (N_1127,N_289,N_515);
nor U1128 (N_1128,N_187,N_584);
and U1129 (N_1129,N_291,N_737);
or U1130 (N_1130,N_326,N_89);
or U1131 (N_1131,N_391,N_287);
or U1132 (N_1132,N_649,N_713);
nor U1133 (N_1133,N_124,N_769);
and U1134 (N_1134,N_198,N_703);
xnor U1135 (N_1135,N_487,N_147);
or U1136 (N_1136,N_466,N_188);
or U1137 (N_1137,N_571,N_492);
nand U1138 (N_1138,N_7,N_477);
or U1139 (N_1139,N_801,N_67);
nand U1140 (N_1140,N_164,N_413);
xor U1141 (N_1141,N_504,N_235);
or U1142 (N_1142,N_864,N_194);
nor U1143 (N_1143,N_930,N_186);
xnor U1144 (N_1144,N_997,N_169);
and U1145 (N_1145,N_817,N_80);
and U1146 (N_1146,N_714,N_602);
xor U1147 (N_1147,N_578,N_803);
nor U1148 (N_1148,N_166,N_108);
and U1149 (N_1149,N_149,N_132);
xor U1150 (N_1150,N_441,N_440);
nor U1151 (N_1151,N_760,N_559);
xor U1152 (N_1152,N_561,N_741);
nor U1153 (N_1153,N_656,N_393);
xnor U1154 (N_1154,N_919,N_476);
nand U1155 (N_1155,N_757,N_553);
and U1156 (N_1156,N_71,N_532);
xnor U1157 (N_1157,N_511,N_576);
xor U1158 (N_1158,N_952,N_954);
nor U1159 (N_1159,N_993,N_325);
and U1160 (N_1160,N_695,N_923);
xnor U1161 (N_1161,N_562,N_770);
nand U1162 (N_1162,N_898,N_368);
and U1163 (N_1163,N_955,N_172);
xor U1164 (N_1164,N_739,N_61);
nand U1165 (N_1165,N_384,N_662);
or U1166 (N_1166,N_18,N_365);
nand U1167 (N_1167,N_647,N_429);
or U1168 (N_1168,N_26,N_258);
nand U1169 (N_1169,N_113,N_179);
or U1170 (N_1170,N_761,N_439);
nor U1171 (N_1171,N_846,N_254);
nor U1172 (N_1172,N_577,N_28);
and U1173 (N_1173,N_296,N_797);
xor U1174 (N_1174,N_358,N_362);
and U1175 (N_1175,N_987,N_344);
or U1176 (N_1176,N_618,N_270);
nand U1177 (N_1177,N_10,N_931);
nor U1178 (N_1178,N_133,N_909);
nand U1179 (N_1179,N_195,N_153);
and U1180 (N_1180,N_754,N_381);
xnor U1181 (N_1181,N_591,N_735);
or U1182 (N_1182,N_351,N_636);
and U1183 (N_1183,N_249,N_749);
nand U1184 (N_1184,N_244,N_535);
and U1185 (N_1185,N_292,N_691);
nor U1186 (N_1186,N_827,N_980);
nor U1187 (N_1187,N_808,N_252);
nor U1188 (N_1188,N_479,N_86);
or U1189 (N_1189,N_711,N_184);
xnor U1190 (N_1190,N_349,N_174);
nor U1191 (N_1191,N_210,N_53);
nor U1192 (N_1192,N_679,N_879);
nor U1193 (N_1193,N_543,N_700);
and U1194 (N_1194,N_778,N_523);
or U1195 (N_1195,N_632,N_199);
xor U1196 (N_1196,N_96,N_678);
xnor U1197 (N_1197,N_464,N_569);
nor U1198 (N_1198,N_453,N_998);
xnor U1199 (N_1199,N_47,N_887);
and U1200 (N_1200,N_920,N_773);
or U1201 (N_1201,N_196,N_375);
and U1202 (N_1202,N_825,N_60);
nor U1203 (N_1203,N_725,N_842);
or U1204 (N_1204,N_355,N_45);
or U1205 (N_1205,N_631,N_594);
or U1206 (N_1206,N_906,N_112);
xnor U1207 (N_1207,N_899,N_556);
nor U1208 (N_1208,N_816,N_957);
or U1209 (N_1209,N_860,N_866);
nand U1210 (N_1210,N_518,N_373);
nand U1211 (N_1211,N_478,N_823);
or U1212 (N_1212,N_135,N_465);
xnor U1213 (N_1213,N_645,N_382);
nand U1214 (N_1214,N_639,N_213);
xor U1215 (N_1215,N_36,N_692);
or U1216 (N_1216,N_759,N_456);
nand U1217 (N_1217,N_11,N_619);
and U1218 (N_1218,N_534,N_20);
xor U1219 (N_1219,N_319,N_724);
nand U1220 (N_1220,N_496,N_506);
or U1221 (N_1221,N_228,N_144);
xnor U1222 (N_1222,N_628,N_763);
and U1223 (N_1223,N_66,N_346);
and U1224 (N_1224,N_13,N_572);
and U1225 (N_1225,N_748,N_77);
nor U1226 (N_1226,N_91,N_687);
xnor U1227 (N_1227,N_625,N_158);
nand U1228 (N_1228,N_621,N_885);
and U1229 (N_1229,N_780,N_315);
xnor U1230 (N_1230,N_807,N_935);
nand U1231 (N_1231,N_185,N_155);
nor U1232 (N_1232,N_922,N_81);
and U1233 (N_1233,N_84,N_190);
nor U1234 (N_1234,N_222,N_274);
or U1235 (N_1235,N_421,N_936);
xor U1236 (N_1236,N_111,N_4);
or U1237 (N_1237,N_131,N_183);
nand U1238 (N_1238,N_9,N_299);
nor U1239 (N_1239,N_966,N_643);
xor U1240 (N_1240,N_288,N_98);
nor U1241 (N_1241,N_447,N_205);
xor U1242 (N_1242,N_926,N_500);
xnor U1243 (N_1243,N_683,N_115);
xnor U1244 (N_1244,N_279,N_708);
and U1245 (N_1245,N_983,N_472);
or U1246 (N_1246,N_814,N_148);
nor U1247 (N_1247,N_231,N_420);
or U1248 (N_1248,N_312,N_855);
nor U1249 (N_1249,N_208,N_716);
nand U1250 (N_1250,N_682,N_834);
xor U1251 (N_1251,N_387,N_101);
xnor U1252 (N_1252,N_731,N_163);
or U1253 (N_1253,N_876,N_490);
and U1254 (N_1254,N_969,N_428);
nand U1255 (N_1255,N_388,N_771);
or U1256 (N_1256,N_307,N_438);
or U1257 (N_1257,N_574,N_379);
and U1258 (N_1258,N_385,N_306);
nand U1259 (N_1259,N_974,N_339);
nor U1260 (N_1260,N_34,N_145);
or U1261 (N_1261,N_972,N_396);
or U1262 (N_1262,N_990,N_843);
nor U1263 (N_1263,N_861,N_245);
or U1264 (N_1264,N_844,N_201);
or U1265 (N_1265,N_530,N_12);
or U1266 (N_1266,N_961,N_837);
nand U1267 (N_1267,N_273,N_822);
nor U1268 (N_1268,N_555,N_730);
xor U1269 (N_1269,N_712,N_90);
or U1270 (N_1270,N_698,N_671);
and U1271 (N_1271,N_471,N_0);
nor U1272 (N_1272,N_87,N_227);
and U1273 (N_1273,N_747,N_776);
nor U1274 (N_1274,N_14,N_637);
and U1275 (N_1275,N_774,N_995);
nor U1276 (N_1276,N_267,N_293);
nor U1277 (N_1277,N_719,N_751);
nor U1278 (N_1278,N_681,N_23);
xnor U1279 (N_1279,N_821,N_988);
and U1280 (N_1280,N_336,N_845);
or U1281 (N_1281,N_237,N_128);
and U1282 (N_1282,N_524,N_103);
or U1283 (N_1283,N_950,N_203);
nor U1284 (N_1284,N_116,N_117);
xnor U1285 (N_1285,N_389,N_38);
nor U1286 (N_1286,N_300,N_335);
nand U1287 (N_1287,N_513,N_400);
or U1288 (N_1288,N_16,N_197);
xnor U1289 (N_1289,N_260,N_787);
xnor U1290 (N_1290,N_996,N_33);
xor U1291 (N_1291,N_85,N_207);
and U1292 (N_1292,N_820,N_311);
or U1293 (N_1293,N_129,N_786);
nand U1294 (N_1294,N_322,N_411);
or U1295 (N_1295,N_461,N_766);
nand U1296 (N_1296,N_241,N_783);
nand U1297 (N_1297,N_910,N_150);
and U1298 (N_1298,N_83,N_170);
and U1299 (N_1299,N_908,N_903);
or U1300 (N_1300,N_608,N_371);
nand U1301 (N_1301,N_790,N_220);
and U1302 (N_1302,N_588,N_762);
xor U1303 (N_1303,N_206,N_97);
and U1304 (N_1304,N_473,N_57);
and U1305 (N_1305,N_540,N_788);
nand U1306 (N_1306,N_357,N_494);
and U1307 (N_1307,N_579,N_276);
xnor U1308 (N_1308,N_324,N_407);
or U1309 (N_1309,N_605,N_833);
or U1310 (N_1310,N_593,N_99);
nor U1311 (N_1311,N_79,N_654);
nor U1312 (N_1312,N_100,N_520);
xor U1313 (N_1313,N_282,N_813);
nand U1314 (N_1314,N_932,N_136);
nor U1315 (N_1315,N_986,N_269);
nor U1316 (N_1316,N_286,N_964);
and U1317 (N_1317,N_498,N_226);
nor U1318 (N_1318,N_114,N_706);
xor U1319 (N_1319,N_657,N_734);
and U1320 (N_1320,N_949,N_24);
nor U1321 (N_1321,N_831,N_668);
and U1322 (N_1322,N_55,N_583);
xnor U1323 (N_1323,N_43,N_348);
or U1324 (N_1324,N_868,N_599);
and U1325 (N_1325,N_283,N_884);
or U1326 (N_1326,N_281,N_586);
nor U1327 (N_1327,N_688,N_924);
nor U1328 (N_1328,N_642,N_211);
and U1329 (N_1329,N_800,N_284);
nand U1330 (N_1330,N_366,N_181);
nor U1331 (N_1331,N_8,N_138);
and U1332 (N_1332,N_323,N_824);
and U1333 (N_1333,N_881,N_661);
or U1334 (N_1334,N_434,N_907);
and U1335 (N_1335,N_880,N_268);
nand U1336 (N_1336,N_653,N_329);
or U1337 (N_1337,N_606,N_76);
nor U1338 (N_1338,N_105,N_547);
nand U1339 (N_1339,N_247,N_756);
and U1340 (N_1340,N_123,N_793);
or U1341 (N_1341,N_512,N_452);
nand U1342 (N_1342,N_705,N_321);
nor U1343 (N_1343,N_917,N_872);
or U1344 (N_1344,N_806,N_404);
nor U1345 (N_1345,N_673,N_141);
xor U1346 (N_1346,N_180,N_640);
and U1347 (N_1347,N_603,N_869);
nor U1348 (N_1348,N_414,N_192);
xor U1349 (N_1349,N_744,N_951);
and U1350 (N_1350,N_463,N_596);
or U1351 (N_1351,N_64,N_914);
nor U1352 (N_1352,N_294,N_401);
nand U1353 (N_1353,N_612,N_156);
and U1354 (N_1354,N_427,N_727);
nor U1355 (N_1355,N_944,N_121);
nand U1356 (N_1356,N_740,N_537);
or U1357 (N_1357,N_272,N_539);
or U1358 (N_1358,N_528,N_200);
nand U1359 (N_1359,N_497,N_442);
nor U1360 (N_1360,N_229,N_449);
xnor U1361 (N_1361,N_650,N_854);
xor U1362 (N_1362,N_22,N_376);
and U1363 (N_1363,N_729,N_328);
and U1364 (N_1364,N_517,N_728);
or U1365 (N_1365,N_826,N_223);
or U1366 (N_1366,N_893,N_655);
nor U1367 (N_1367,N_474,N_50);
or U1368 (N_1368,N_610,N_558);
or U1369 (N_1369,N_667,N_977);
and U1370 (N_1370,N_753,N_784);
xnor U1371 (N_1371,N_5,N_723);
and U1372 (N_1372,N_811,N_457);
and U1373 (N_1373,N_810,N_342);
or U1374 (N_1374,N_1,N_3);
and U1375 (N_1375,N_130,N_796);
nor U1376 (N_1376,N_616,N_857);
and U1377 (N_1377,N_819,N_675);
nand U1378 (N_1378,N_828,N_72);
xnor U1379 (N_1379,N_614,N_501);
nand U1380 (N_1380,N_347,N_508);
and U1381 (N_1381,N_615,N_902);
nor U1382 (N_1382,N_109,N_403);
and U1383 (N_1383,N_510,N_848);
nand U1384 (N_1384,N_377,N_332);
or U1385 (N_1385,N_767,N_611);
and U1386 (N_1386,N_305,N_928);
nor U1387 (N_1387,N_142,N_533);
nor U1388 (N_1388,N_94,N_609);
xnor U1389 (N_1389,N_191,N_641);
and U1390 (N_1390,N_175,N_285);
xor U1391 (N_1391,N_52,N_867);
xor U1392 (N_1392,N_911,N_772);
nand U1393 (N_1393,N_168,N_840);
nor U1394 (N_1394,N_551,N_745);
nor U1395 (N_1395,N_40,N_925);
xnor U1396 (N_1396,N_359,N_839);
and U1397 (N_1397,N_721,N_689);
or U1398 (N_1398,N_122,N_51);
nand U1399 (N_1399,N_176,N_963);
and U1400 (N_1400,N_69,N_550);
or U1401 (N_1401,N_383,N_225);
and U1402 (N_1402,N_613,N_994);
nand U1403 (N_1403,N_309,N_486);
or U1404 (N_1404,N_781,N_62);
or U1405 (N_1405,N_587,N_458);
nor U1406 (N_1406,N_310,N_455);
xor U1407 (N_1407,N_720,N_580);
or U1408 (N_1408,N_308,N_709);
and U1409 (N_1409,N_363,N_451);
and U1410 (N_1410,N_29,N_552);
nand U1411 (N_1411,N_514,N_888);
xnor U1412 (N_1412,N_858,N_798);
nand U1413 (N_1413,N_42,N_397);
or U1414 (N_1414,N_469,N_157);
xor U1415 (N_1415,N_809,N_352);
xor U1416 (N_1416,N_257,N_519);
nand U1417 (N_1417,N_526,N_320);
nor U1418 (N_1418,N_154,N_345);
nor U1419 (N_1419,N_557,N_63);
xnor U1420 (N_1420,N_298,N_620);
or U1421 (N_1421,N_722,N_482);
xor U1422 (N_1422,N_446,N_849);
and U1423 (N_1423,N_981,N_804);
and U1424 (N_1424,N_941,N_601);
nand U1425 (N_1425,N_743,N_648);
or U1426 (N_1426,N_882,N_495);
or U1427 (N_1427,N_460,N_215);
or U1428 (N_1428,N_160,N_991);
xnor U1429 (N_1429,N_847,N_738);
nand U1430 (N_1430,N_302,N_736);
or U1431 (N_1431,N_718,N_794);
nand U1432 (N_1432,N_118,N_850);
nand U1433 (N_1433,N_317,N_484);
xor U1434 (N_1434,N_732,N_485);
nor U1435 (N_1435,N_423,N_742);
nor U1436 (N_1436,N_263,N_318);
nand U1437 (N_1437,N_812,N_409);
nand U1438 (N_1438,N_436,N_795);
or U1439 (N_1439,N_905,N_65);
nor U1440 (N_1440,N_663,N_93);
nor U1441 (N_1441,N_251,N_264);
nor U1442 (N_1442,N_965,N_585);
and U1443 (N_1443,N_775,N_127);
nand U1444 (N_1444,N_49,N_350);
nand U1445 (N_1445,N_146,N_913);
xnor U1446 (N_1446,N_862,N_443);
and U1447 (N_1447,N_542,N_567);
nor U1448 (N_1448,N_975,N_598);
nand U1449 (N_1449,N_554,N_939);
nand U1450 (N_1450,N_633,N_246);
nand U1451 (N_1451,N_92,N_916);
or U1452 (N_1452,N_304,N_416);
nand U1453 (N_1453,N_765,N_629);
nor U1454 (N_1454,N_475,N_777);
nand U1455 (N_1455,N_651,N_685);
or U1456 (N_1456,N_710,N_433);
nand U1457 (N_1457,N_44,N_412);
nor U1458 (N_1458,N_430,N_483);
nor U1459 (N_1459,N_536,N_46);
or U1460 (N_1460,N_295,N_779);
nand U1461 (N_1461,N_107,N_139);
nor U1462 (N_1462,N_15,N_746);
and U1463 (N_1463,N_271,N_992);
nand U1464 (N_1464,N_853,N_627);
and U1465 (N_1465,N_531,N_921);
and U1466 (N_1466,N_82,N_573);
and U1467 (N_1467,N_516,N_886);
xnor U1468 (N_1468,N_239,N_694);
and U1469 (N_1469,N_219,N_361);
nand U1470 (N_1470,N_750,N_21);
nor U1471 (N_1471,N_221,N_953);
nand U1472 (N_1472,N_337,N_956);
nand U1473 (N_1473,N_445,N_340);
or U1474 (N_1474,N_890,N_999);
and U1475 (N_1475,N_892,N_59);
nor U1476 (N_1476,N_560,N_334);
xor U1477 (N_1477,N_697,N_676);
nor U1478 (N_1478,N_262,N_940);
nand U1479 (N_1479,N_193,N_702);
nor U1480 (N_1480,N_527,N_883);
and U1481 (N_1481,N_755,N_415);
nand U1482 (N_1482,N_217,N_275);
nor U1483 (N_1483,N_665,N_707);
and U1484 (N_1484,N_693,N_68);
nand U1485 (N_1485,N_836,N_959);
and U1486 (N_1486,N_900,N_938);
or U1487 (N_1487,N_863,N_491);
nor U1488 (N_1488,N_189,N_30);
nor U1489 (N_1489,N_354,N_462);
or U1490 (N_1490,N_173,N_327);
and U1491 (N_1491,N_448,N_454);
or U1492 (N_1492,N_575,N_417);
or U1493 (N_1493,N_976,N_35);
nand U1494 (N_1494,N_277,N_73);
and U1495 (N_1495,N_859,N_945);
or U1496 (N_1496,N_946,N_31);
xnor U1497 (N_1497,N_877,N_19);
and U1498 (N_1498,N_236,N_934);
xor U1499 (N_1499,N_960,N_290);
and U1500 (N_1500,N_531,N_421);
nand U1501 (N_1501,N_421,N_647);
and U1502 (N_1502,N_46,N_841);
nor U1503 (N_1503,N_274,N_664);
nor U1504 (N_1504,N_51,N_803);
nand U1505 (N_1505,N_215,N_84);
or U1506 (N_1506,N_433,N_381);
xnor U1507 (N_1507,N_788,N_764);
nand U1508 (N_1508,N_705,N_309);
xor U1509 (N_1509,N_29,N_684);
or U1510 (N_1510,N_848,N_343);
and U1511 (N_1511,N_180,N_72);
and U1512 (N_1512,N_604,N_482);
or U1513 (N_1513,N_674,N_819);
and U1514 (N_1514,N_985,N_417);
nand U1515 (N_1515,N_945,N_184);
and U1516 (N_1516,N_29,N_427);
nand U1517 (N_1517,N_86,N_908);
nor U1518 (N_1518,N_98,N_669);
or U1519 (N_1519,N_800,N_468);
nand U1520 (N_1520,N_745,N_848);
xnor U1521 (N_1521,N_48,N_794);
or U1522 (N_1522,N_277,N_783);
and U1523 (N_1523,N_613,N_611);
nand U1524 (N_1524,N_495,N_30);
xor U1525 (N_1525,N_396,N_393);
and U1526 (N_1526,N_303,N_353);
or U1527 (N_1527,N_645,N_727);
nand U1528 (N_1528,N_989,N_303);
nor U1529 (N_1529,N_556,N_888);
xor U1530 (N_1530,N_675,N_996);
nor U1531 (N_1531,N_796,N_139);
and U1532 (N_1532,N_369,N_755);
xnor U1533 (N_1533,N_693,N_774);
nor U1534 (N_1534,N_572,N_57);
nand U1535 (N_1535,N_368,N_799);
nand U1536 (N_1536,N_98,N_803);
nor U1537 (N_1537,N_425,N_69);
xor U1538 (N_1538,N_86,N_635);
xor U1539 (N_1539,N_84,N_179);
and U1540 (N_1540,N_209,N_539);
and U1541 (N_1541,N_779,N_770);
nand U1542 (N_1542,N_520,N_454);
or U1543 (N_1543,N_239,N_618);
xnor U1544 (N_1544,N_846,N_258);
or U1545 (N_1545,N_686,N_942);
and U1546 (N_1546,N_287,N_794);
nand U1547 (N_1547,N_400,N_432);
or U1548 (N_1548,N_614,N_506);
nand U1549 (N_1549,N_205,N_962);
and U1550 (N_1550,N_441,N_288);
and U1551 (N_1551,N_42,N_218);
xor U1552 (N_1552,N_735,N_98);
and U1553 (N_1553,N_410,N_382);
or U1554 (N_1554,N_923,N_198);
and U1555 (N_1555,N_342,N_907);
nand U1556 (N_1556,N_928,N_267);
and U1557 (N_1557,N_186,N_6);
nand U1558 (N_1558,N_895,N_609);
xor U1559 (N_1559,N_551,N_607);
or U1560 (N_1560,N_718,N_159);
xor U1561 (N_1561,N_366,N_517);
and U1562 (N_1562,N_153,N_114);
xnor U1563 (N_1563,N_190,N_419);
xnor U1564 (N_1564,N_116,N_658);
xor U1565 (N_1565,N_715,N_975);
or U1566 (N_1566,N_334,N_834);
xnor U1567 (N_1567,N_100,N_219);
nor U1568 (N_1568,N_385,N_86);
and U1569 (N_1569,N_850,N_493);
nor U1570 (N_1570,N_172,N_682);
nand U1571 (N_1571,N_278,N_640);
nand U1572 (N_1572,N_112,N_788);
or U1573 (N_1573,N_53,N_387);
nand U1574 (N_1574,N_839,N_395);
or U1575 (N_1575,N_392,N_48);
xor U1576 (N_1576,N_663,N_179);
or U1577 (N_1577,N_646,N_977);
or U1578 (N_1578,N_633,N_932);
nor U1579 (N_1579,N_538,N_210);
and U1580 (N_1580,N_641,N_140);
or U1581 (N_1581,N_913,N_748);
xnor U1582 (N_1582,N_293,N_575);
nand U1583 (N_1583,N_406,N_216);
or U1584 (N_1584,N_408,N_962);
nand U1585 (N_1585,N_131,N_578);
nor U1586 (N_1586,N_343,N_938);
nor U1587 (N_1587,N_568,N_619);
nand U1588 (N_1588,N_162,N_424);
nand U1589 (N_1589,N_72,N_830);
xnor U1590 (N_1590,N_702,N_123);
nor U1591 (N_1591,N_73,N_383);
or U1592 (N_1592,N_132,N_771);
and U1593 (N_1593,N_837,N_679);
nand U1594 (N_1594,N_734,N_466);
nand U1595 (N_1595,N_819,N_407);
and U1596 (N_1596,N_451,N_464);
and U1597 (N_1597,N_752,N_980);
nand U1598 (N_1598,N_411,N_94);
nand U1599 (N_1599,N_419,N_23);
or U1600 (N_1600,N_252,N_83);
or U1601 (N_1601,N_946,N_584);
nor U1602 (N_1602,N_378,N_886);
nand U1603 (N_1603,N_286,N_944);
nor U1604 (N_1604,N_488,N_313);
and U1605 (N_1605,N_876,N_256);
nand U1606 (N_1606,N_31,N_649);
nand U1607 (N_1607,N_888,N_942);
and U1608 (N_1608,N_957,N_619);
nand U1609 (N_1609,N_972,N_130);
nor U1610 (N_1610,N_427,N_936);
nor U1611 (N_1611,N_869,N_340);
nor U1612 (N_1612,N_210,N_331);
and U1613 (N_1613,N_971,N_786);
nor U1614 (N_1614,N_90,N_840);
xor U1615 (N_1615,N_893,N_192);
nand U1616 (N_1616,N_928,N_223);
or U1617 (N_1617,N_827,N_160);
nor U1618 (N_1618,N_848,N_913);
and U1619 (N_1619,N_396,N_606);
nand U1620 (N_1620,N_170,N_506);
or U1621 (N_1621,N_819,N_497);
or U1622 (N_1622,N_969,N_282);
and U1623 (N_1623,N_633,N_44);
xnor U1624 (N_1624,N_285,N_334);
and U1625 (N_1625,N_704,N_349);
and U1626 (N_1626,N_963,N_370);
or U1627 (N_1627,N_272,N_19);
and U1628 (N_1628,N_338,N_935);
nor U1629 (N_1629,N_530,N_883);
and U1630 (N_1630,N_45,N_905);
nor U1631 (N_1631,N_971,N_153);
nor U1632 (N_1632,N_876,N_198);
xor U1633 (N_1633,N_458,N_202);
or U1634 (N_1634,N_274,N_584);
and U1635 (N_1635,N_335,N_917);
and U1636 (N_1636,N_277,N_198);
and U1637 (N_1637,N_973,N_945);
nor U1638 (N_1638,N_467,N_833);
and U1639 (N_1639,N_152,N_158);
nand U1640 (N_1640,N_213,N_98);
nand U1641 (N_1641,N_737,N_556);
nand U1642 (N_1642,N_68,N_759);
nor U1643 (N_1643,N_438,N_295);
xnor U1644 (N_1644,N_671,N_47);
or U1645 (N_1645,N_942,N_166);
and U1646 (N_1646,N_470,N_619);
and U1647 (N_1647,N_70,N_974);
nor U1648 (N_1648,N_991,N_424);
xnor U1649 (N_1649,N_407,N_640);
nand U1650 (N_1650,N_987,N_813);
and U1651 (N_1651,N_53,N_940);
nand U1652 (N_1652,N_28,N_154);
xnor U1653 (N_1653,N_773,N_270);
xor U1654 (N_1654,N_631,N_806);
and U1655 (N_1655,N_169,N_77);
or U1656 (N_1656,N_363,N_870);
xnor U1657 (N_1657,N_161,N_464);
and U1658 (N_1658,N_371,N_546);
xor U1659 (N_1659,N_319,N_263);
xor U1660 (N_1660,N_705,N_209);
or U1661 (N_1661,N_917,N_236);
nor U1662 (N_1662,N_327,N_609);
nor U1663 (N_1663,N_852,N_523);
xor U1664 (N_1664,N_51,N_120);
nand U1665 (N_1665,N_719,N_306);
xor U1666 (N_1666,N_485,N_677);
and U1667 (N_1667,N_482,N_620);
nand U1668 (N_1668,N_49,N_787);
nand U1669 (N_1669,N_571,N_570);
and U1670 (N_1670,N_4,N_739);
nor U1671 (N_1671,N_801,N_103);
xor U1672 (N_1672,N_9,N_309);
and U1673 (N_1673,N_257,N_914);
and U1674 (N_1674,N_432,N_784);
xnor U1675 (N_1675,N_34,N_815);
or U1676 (N_1676,N_958,N_367);
or U1677 (N_1677,N_943,N_870);
nor U1678 (N_1678,N_420,N_803);
xnor U1679 (N_1679,N_219,N_653);
and U1680 (N_1680,N_298,N_207);
nand U1681 (N_1681,N_43,N_946);
nor U1682 (N_1682,N_513,N_527);
nor U1683 (N_1683,N_31,N_239);
or U1684 (N_1684,N_419,N_14);
nor U1685 (N_1685,N_942,N_804);
and U1686 (N_1686,N_54,N_519);
nor U1687 (N_1687,N_917,N_345);
and U1688 (N_1688,N_245,N_808);
xor U1689 (N_1689,N_354,N_266);
nor U1690 (N_1690,N_112,N_464);
or U1691 (N_1691,N_104,N_221);
and U1692 (N_1692,N_822,N_248);
nand U1693 (N_1693,N_184,N_279);
or U1694 (N_1694,N_331,N_414);
xnor U1695 (N_1695,N_386,N_52);
nand U1696 (N_1696,N_742,N_198);
nor U1697 (N_1697,N_416,N_734);
nor U1698 (N_1698,N_117,N_171);
or U1699 (N_1699,N_429,N_166);
nand U1700 (N_1700,N_237,N_341);
nand U1701 (N_1701,N_864,N_106);
and U1702 (N_1702,N_193,N_180);
xor U1703 (N_1703,N_400,N_595);
xor U1704 (N_1704,N_883,N_805);
nor U1705 (N_1705,N_244,N_433);
nor U1706 (N_1706,N_766,N_843);
xnor U1707 (N_1707,N_108,N_839);
xor U1708 (N_1708,N_79,N_981);
xnor U1709 (N_1709,N_752,N_538);
xnor U1710 (N_1710,N_223,N_858);
xor U1711 (N_1711,N_506,N_644);
or U1712 (N_1712,N_713,N_807);
nor U1713 (N_1713,N_775,N_712);
and U1714 (N_1714,N_161,N_655);
nor U1715 (N_1715,N_30,N_666);
or U1716 (N_1716,N_393,N_115);
nor U1717 (N_1717,N_555,N_387);
nor U1718 (N_1718,N_600,N_982);
or U1719 (N_1719,N_273,N_809);
nand U1720 (N_1720,N_53,N_876);
and U1721 (N_1721,N_36,N_654);
nand U1722 (N_1722,N_481,N_943);
and U1723 (N_1723,N_578,N_174);
and U1724 (N_1724,N_83,N_452);
or U1725 (N_1725,N_665,N_832);
and U1726 (N_1726,N_128,N_443);
and U1727 (N_1727,N_51,N_249);
nand U1728 (N_1728,N_903,N_373);
nor U1729 (N_1729,N_197,N_967);
or U1730 (N_1730,N_394,N_367);
xor U1731 (N_1731,N_208,N_486);
nor U1732 (N_1732,N_252,N_333);
nor U1733 (N_1733,N_681,N_247);
nor U1734 (N_1734,N_176,N_502);
nor U1735 (N_1735,N_969,N_167);
and U1736 (N_1736,N_721,N_294);
nand U1737 (N_1737,N_311,N_145);
or U1738 (N_1738,N_953,N_932);
or U1739 (N_1739,N_842,N_12);
nor U1740 (N_1740,N_575,N_361);
and U1741 (N_1741,N_42,N_623);
or U1742 (N_1742,N_849,N_932);
and U1743 (N_1743,N_49,N_113);
nor U1744 (N_1744,N_180,N_775);
xnor U1745 (N_1745,N_93,N_544);
or U1746 (N_1746,N_0,N_755);
nand U1747 (N_1747,N_100,N_930);
nand U1748 (N_1748,N_932,N_96);
or U1749 (N_1749,N_986,N_7);
xor U1750 (N_1750,N_935,N_135);
nor U1751 (N_1751,N_489,N_577);
xor U1752 (N_1752,N_408,N_698);
and U1753 (N_1753,N_773,N_652);
or U1754 (N_1754,N_395,N_153);
and U1755 (N_1755,N_679,N_648);
nor U1756 (N_1756,N_135,N_605);
xor U1757 (N_1757,N_375,N_206);
and U1758 (N_1758,N_294,N_627);
and U1759 (N_1759,N_718,N_914);
nor U1760 (N_1760,N_861,N_130);
and U1761 (N_1761,N_829,N_449);
or U1762 (N_1762,N_706,N_363);
nand U1763 (N_1763,N_452,N_878);
nand U1764 (N_1764,N_408,N_158);
nand U1765 (N_1765,N_395,N_213);
xnor U1766 (N_1766,N_219,N_194);
and U1767 (N_1767,N_586,N_449);
or U1768 (N_1768,N_308,N_932);
and U1769 (N_1769,N_1,N_654);
xnor U1770 (N_1770,N_706,N_537);
and U1771 (N_1771,N_232,N_95);
or U1772 (N_1772,N_153,N_929);
and U1773 (N_1773,N_846,N_392);
or U1774 (N_1774,N_3,N_950);
xor U1775 (N_1775,N_802,N_411);
and U1776 (N_1776,N_351,N_962);
nand U1777 (N_1777,N_709,N_750);
nand U1778 (N_1778,N_743,N_546);
and U1779 (N_1779,N_892,N_108);
or U1780 (N_1780,N_386,N_441);
xor U1781 (N_1781,N_930,N_403);
and U1782 (N_1782,N_692,N_319);
xnor U1783 (N_1783,N_716,N_921);
and U1784 (N_1784,N_661,N_251);
nor U1785 (N_1785,N_696,N_473);
or U1786 (N_1786,N_462,N_485);
and U1787 (N_1787,N_426,N_541);
xnor U1788 (N_1788,N_941,N_278);
nor U1789 (N_1789,N_962,N_150);
and U1790 (N_1790,N_955,N_904);
xnor U1791 (N_1791,N_397,N_609);
or U1792 (N_1792,N_541,N_680);
xor U1793 (N_1793,N_663,N_495);
nand U1794 (N_1794,N_633,N_953);
nand U1795 (N_1795,N_616,N_800);
or U1796 (N_1796,N_573,N_804);
and U1797 (N_1797,N_913,N_33);
or U1798 (N_1798,N_141,N_201);
and U1799 (N_1799,N_151,N_908);
nand U1800 (N_1800,N_173,N_802);
and U1801 (N_1801,N_199,N_876);
xor U1802 (N_1802,N_997,N_913);
xor U1803 (N_1803,N_451,N_870);
and U1804 (N_1804,N_412,N_860);
nand U1805 (N_1805,N_325,N_262);
or U1806 (N_1806,N_958,N_407);
or U1807 (N_1807,N_600,N_35);
nor U1808 (N_1808,N_912,N_438);
or U1809 (N_1809,N_666,N_564);
or U1810 (N_1810,N_243,N_534);
or U1811 (N_1811,N_660,N_765);
and U1812 (N_1812,N_141,N_771);
nand U1813 (N_1813,N_823,N_778);
or U1814 (N_1814,N_976,N_820);
xor U1815 (N_1815,N_13,N_963);
nand U1816 (N_1816,N_615,N_828);
or U1817 (N_1817,N_686,N_290);
and U1818 (N_1818,N_602,N_285);
nor U1819 (N_1819,N_866,N_336);
and U1820 (N_1820,N_672,N_389);
nor U1821 (N_1821,N_950,N_397);
xnor U1822 (N_1822,N_397,N_767);
xor U1823 (N_1823,N_234,N_301);
nand U1824 (N_1824,N_162,N_507);
or U1825 (N_1825,N_865,N_658);
or U1826 (N_1826,N_576,N_505);
and U1827 (N_1827,N_334,N_506);
and U1828 (N_1828,N_627,N_888);
nor U1829 (N_1829,N_424,N_123);
or U1830 (N_1830,N_423,N_148);
nor U1831 (N_1831,N_737,N_685);
nor U1832 (N_1832,N_994,N_930);
and U1833 (N_1833,N_978,N_411);
and U1834 (N_1834,N_26,N_104);
nor U1835 (N_1835,N_161,N_826);
or U1836 (N_1836,N_385,N_778);
or U1837 (N_1837,N_44,N_624);
and U1838 (N_1838,N_856,N_667);
and U1839 (N_1839,N_560,N_956);
xnor U1840 (N_1840,N_376,N_470);
and U1841 (N_1841,N_330,N_125);
or U1842 (N_1842,N_698,N_365);
nand U1843 (N_1843,N_877,N_95);
nand U1844 (N_1844,N_744,N_753);
and U1845 (N_1845,N_334,N_220);
xnor U1846 (N_1846,N_792,N_600);
xor U1847 (N_1847,N_880,N_847);
nand U1848 (N_1848,N_214,N_154);
xnor U1849 (N_1849,N_322,N_748);
xor U1850 (N_1850,N_95,N_718);
xor U1851 (N_1851,N_744,N_849);
nand U1852 (N_1852,N_495,N_676);
nand U1853 (N_1853,N_594,N_893);
and U1854 (N_1854,N_633,N_856);
nor U1855 (N_1855,N_442,N_969);
and U1856 (N_1856,N_499,N_554);
or U1857 (N_1857,N_977,N_655);
or U1858 (N_1858,N_396,N_613);
xor U1859 (N_1859,N_558,N_907);
nand U1860 (N_1860,N_196,N_784);
or U1861 (N_1861,N_580,N_389);
nand U1862 (N_1862,N_829,N_599);
nand U1863 (N_1863,N_24,N_302);
and U1864 (N_1864,N_694,N_828);
xor U1865 (N_1865,N_222,N_7);
and U1866 (N_1866,N_207,N_694);
or U1867 (N_1867,N_650,N_797);
nor U1868 (N_1868,N_666,N_209);
xor U1869 (N_1869,N_593,N_670);
xnor U1870 (N_1870,N_158,N_518);
nor U1871 (N_1871,N_826,N_378);
xnor U1872 (N_1872,N_595,N_167);
or U1873 (N_1873,N_724,N_340);
or U1874 (N_1874,N_659,N_748);
nand U1875 (N_1875,N_577,N_387);
nor U1876 (N_1876,N_917,N_874);
nor U1877 (N_1877,N_60,N_15);
xnor U1878 (N_1878,N_851,N_692);
and U1879 (N_1879,N_546,N_187);
nor U1880 (N_1880,N_547,N_557);
nor U1881 (N_1881,N_388,N_514);
or U1882 (N_1882,N_783,N_37);
or U1883 (N_1883,N_322,N_999);
xnor U1884 (N_1884,N_730,N_91);
nor U1885 (N_1885,N_494,N_159);
xor U1886 (N_1886,N_83,N_873);
nor U1887 (N_1887,N_38,N_550);
xnor U1888 (N_1888,N_52,N_718);
and U1889 (N_1889,N_24,N_191);
and U1890 (N_1890,N_645,N_567);
nand U1891 (N_1891,N_408,N_948);
xnor U1892 (N_1892,N_365,N_697);
nand U1893 (N_1893,N_764,N_259);
nand U1894 (N_1894,N_262,N_46);
xor U1895 (N_1895,N_640,N_548);
xnor U1896 (N_1896,N_205,N_523);
and U1897 (N_1897,N_398,N_477);
xor U1898 (N_1898,N_914,N_771);
nand U1899 (N_1899,N_57,N_260);
or U1900 (N_1900,N_509,N_53);
and U1901 (N_1901,N_632,N_564);
nor U1902 (N_1902,N_77,N_865);
nor U1903 (N_1903,N_900,N_928);
nand U1904 (N_1904,N_192,N_861);
nand U1905 (N_1905,N_899,N_530);
or U1906 (N_1906,N_0,N_947);
nand U1907 (N_1907,N_106,N_880);
nor U1908 (N_1908,N_330,N_114);
nor U1909 (N_1909,N_201,N_809);
nand U1910 (N_1910,N_979,N_939);
xnor U1911 (N_1911,N_783,N_892);
xnor U1912 (N_1912,N_525,N_296);
xor U1913 (N_1913,N_679,N_139);
and U1914 (N_1914,N_839,N_414);
or U1915 (N_1915,N_688,N_163);
nand U1916 (N_1916,N_699,N_323);
xnor U1917 (N_1917,N_541,N_711);
nor U1918 (N_1918,N_935,N_119);
and U1919 (N_1919,N_486,N_910);
or U1920 (N_1920,N_906,N_881);
or U1921 (N_1921,N_915,N_625);
nor U1922 (N_1922,N_646,N_125);
nand U1923 (N_1923,N_738,N_530);
and U1924 (N_1924,N_821,N_775);
nand U1925 (N_1925,N_858,N_25);
nor U1926 (N_1926,N_561,N_129);
and U1927 (N_1927,N_670,N_703);
xor U1928 (N_1928,N_381,N_46);
xnor U1929 (N_1929,N_616,N_36);
xnor U1930 (N_1930,N_834,N_120);
or U1931 (N_1931,N_877,N_792);
or U1932 (N_1932,N_604,N_980);
nand U1933 (N_1933,N_749,N_140);
xor U1934 (N_1934,N_947,N_607);
nand U1935 (N_1935,N_950,N_802);
or U1936 (N_1936,N_754,N_508);
xor U1937 (N_1937,N_749,N_897);
and U1938 (N_1938,N_302,N_685);
xor U1939 (N_1939,N_816,N_679);
or U1940 (N_1940,N_667,N_870);
and U1941 (N_1941,N_757,N_239);
xor U1942 (N_1942,N_570,N_871);
and U1943 (N_1943,N_546,N_556);
and U1944 (N_1944,N_949,N_497);
nand U1945 (N_1945,N_761,N_171);
nor U1946 (N_1946,N_473,N_416);
nand U1947 (N_1947,N_549,N_154);
xor U1948 (N_1948,N_576,N_622);
or U1949 (N_1949,N_744,N_209);
nand U1950 (N_1950,N_243,N_216);
xnor U1951 (N_1951,N_468,N_989);
or U1952 (N_1952,N_450,N_170);
nand U1953 (N_1953,N_251,N_177);
xnor U1954 (N_1954,N_742,N_823);
and U1955 (N_1955,N_112,N_422);
nor U1956 (N_1956,N_531,N_703);
nand U1957 (N_1957,N_814,N_622);
nor U1958 (N_1958,N_978,N_706);
or U1959 (N_1959,N_977,N_74);
or U1960 (N_1960,N_670,N_52);
or U1961 (N_1961,N_192,N_860);
nor U1962 (N_1962,N_293,N_143);
nor U1963 (N_1963,N_361,N_527);
nand U1964 (N_1964,N_262,N_720);
and U1965 (N_1965,N_830,N_99);
or U1966 (N_1966,N_128,N_751);
nor U1967 (N_1967,N_734,N_412);
xor U1968 (N_1968,N_51,N_878);
or U1969 (N_1969,N_815,N_221);
or U1970 (N_1970,N_525,N_472);
nor U1971 (N_1971,N_925,N_299);
nor U1972 (N_1972,N_754,N_490);
nand U1973 (N_1973,N_580,N_170);
xor U1974 (N_1974,N_768,N_620);
xor U1975 (N_1975,N_572,N_541);
or U1976 (N_1976,N_227,N_291);
nor U1977 (N_1977,N_743,N_834);
nor U1978 (N_1978,N_946,N_27);
nor U1979 (N_1979,N_988,N_308);
xnor U1980 (N_1980,N_130,N_654);
nand U1981 (N_1981,N_109,N_161);
xor U1982 (N_1982,N_516,N_859);
nor U1983 (N_1983,N_671,N_836);
or U1984 (N_1984,N_580,N_777);
xor U1985 (N_1985,N_113,N_535);
nor U1986 (N_1986,N_100,N_920);
nand U1987 (N_1987,N_523,N_203);
or U1988 (N_1988,N_167,N_959);
nand U1989 (N_1989,N_623,N_587);
xnor U1990 (N_1990,N_448,N_634);
and U1991 (N_1991,N_355,N_560);
nand U1992 (N_1992,N_609,N_628);
nand U1993 (N_1993,N_232,N_667);
and U1994 (N_1994,N_901,N_409);
nor U1995 (N_1995,N_654,N_304);
and U1996 (N_1996,N_223,N_59);
nor U1997 (N_1997,N_294,N_701);
or U1998 (N_1998,N_189,N_909);
and U1999 (N_1999,N_999,N_293);
and U2000 (N_2000,N_1004,N_1792);
or U2001 (N_2001,N_1513,N_1774);
and U2002 (N_2002,N_1408,N_1080);
or U2003 (N_2003,N_1218,N_1463);
xnor U2004 (N_2004,N_1252,N_1144);
xor U2005 (N_2005,N_1723,N_1962);
and U2006 (N_2006,N_1928,N_1672);
xor U2007 (N_2007,N_1286,N_1251);
or U2008 (N_2008,N_1927,N_1013);
and U2009 (N_2009,N_1068,N_1323);
xor U2010 (N_2010,N_1247,N_1293);
nand U2011 (N_2011,N_1716,N_1757);
xnor U2012 (N_2012,N_1350,N_1507);
nand U2013 (N_2013,N_1549,N_1753);
xor U2014 (N_2014,N_1398,N_1747);
nor U2015 (N_2015,N_1869,N_1070);
nor U2016 (N_2016,N_1721,N_1977);
nand U2017 (N_2017,N_1645,N_1229);
xnor U2018 (N_2018,N_1582,N_1215);
nor U2019 (N_2019,N_1627,N_1801);
or U2020 (N_2020,N_1492,N_1494);
nor U2021 (N_2021,N_1578,N_1955);
xnor U2022 (N_2022,N_1301,N_1608);
xor U2023 (N_2023,N_1857,N_1698);
xor U2024 (N_2024,N_1356,N_1968);
nand U2025 (N_2025,N_1151,N_1586);
or U2026 (N_2026,N_1728,N_1490);
nand U2027 (N_2027,N_1925,N_1339);
and U2028 (N_2028,N_1148,N_1738);
or U2029 (N_2029,N_1106,N_1422);
and U2030 (N_2030,N_1466,N_1566);
nor U2031 (N_2031,N_1420,N_1793);
or U2032 (N_2032,N_1274,N_1732);
nor U2033 (N_2033,N_1481,N_1434);
nand U2034 (N_2034,N_1328,N_1146);
and U2035 (N_2035,N_1181,N_1918);
or U2036 (N_2036,N_1518,N_1132);
and U2037 (N_2037,N_1412,N_1527);
nor U2038 (N_2038,N_1805,N_1235);
nor U2039 (N_2039,N_1444,N_1005);
nand U2040 (N_2040,N_1242,N_1344);
nand U2041 (N_2041,N_1523,N_1543);
nor U2042 (N_2042,N_1307,N_1902);
and U2043 (N_2043,N_1631,N_1326);
and U2044 (N_2044,N_1419,N_1172);
or U2045 (N_2045,N_1401,N_1547);
nand U2046 (N_2046,N_1216,N_1312);
xor U2047 (N_2047,N_1266,N_1887);
nand U2048 (N_2048,N_1634,N_1358);
nand U2049 (N_2049,N_1874,N_1623);
nor U2050 (N_2050,N_1843,N_1833);
and U2051 (N_2051,N_1719,N_1019);
xor U2052 (N_2052,N_1439,N_1773);
nand U2053 (N_2053,N_1671,N_1253);
nor U2054 (N_2054,N_1361,N_1033);
or U2055 (N_2055,N_1249,N_1804);
xnor U2056 (N_2056,N_1550,N_1239);
xor U2057 (N_2057,N_1828,N_1539);
nand U2058 (N_2058,N_1935,N_1120);
and U2059 (N_2059,N_1739,N_1933);
nand U2060 (N_2060,N_1306,N_1016);
and U2061 (N_2061,N_1049,N_1505);
or U2062 (N_2062,N_1662,N_1090);
nor U2063 (N_2063,N_1687,N_1849);
nor U2064 (N_2064,N_1779,N_1017);
xnor U2065 (N_2065,N_1468,N_1820);
nand U2066 (N_2066,N_1467,N_1366);
nand U2067 (N_2067,N_1244,N_1960);
xnor U2068 (N_2068,N_1915,N_1708);
nor U2069 (N_2069,N_1911,N_1609);
xnor U2070 (N_2070,N_1325,N_1161);
and U2071 (N_2071,N_1152,N_1680);
and U2072 (N_2072,N_1938,N_1243);
and U2073 (N_2073,N_1959,N_1245);
nand U2074 (N_2074,N_1029,N_1159);
and U2075 (N_2075,N_1648,N_1473);
nor U2076 (N_2076,N_1612,N_1310);
nand U2077 (N_2077,N_1922,N_1409);
nand U2078 (N_2078,N_1688,N_1866);
and U2079 (N_2079,N_1103,N_1524);
and U2080 (N_2080,N_1559,N_1961);
xnor U2081 (N_2081,N_1093,N_1102);
nand U2082 (N_2082,N_1183,N_1411);
or U2083 (N_2083,N_1240,N_1569);
xor U2084 (N_2084,N_1149,N_1591);
or U2085 (N_2085,N_1607,N_1808);
and U2086 (N_2086,N_1273,N_1896);
and U2087 (N_2087,N_1290,N_1072);
xnor U2088 (N_2088,N_1329,N_1629);
xnor U2089 (N_2089,N_1397,N_1213);
xor U2090 (N_2090,N_1859,N_1652);
or U2091 (N_2091,N_1573,N_1173);
nor U2092 (N_2092,N_1864,N_1502);
and U2093 (N_2093,N_1063,N_1160);
or U2094 (N_2094,N_1075,N_1025);
xnor U2095 (N_2095,N_1296,N_1519);
or U2096 (N_2096,N_1875,N_1830);
xnor U2097 (N_2097,N_1291,N_1632);
nor U2098 (N_2098,N_1980,N_1435);
nor U2099 (N_2099,N_1856,N_1978);
xor U2100 (N_2100,N_1947,N_1641);
nor U2101 (N_2101,N_1186,N_1806);
nand U2102 (N_2102,N_1346,N_1135);
and U2103 (N_2103,N_1690,N_1362);
nand U2104 (N_2104,N_1895,N_1425);
xnor U2105 (N_2105,N_1086,N_1624);
and U2106 (N_2106,N_1258,N_1353);
or U2107 (N_2107,N_1416,N_1749);
or U2108 (N_2108,N_1133,N_1876);
xor U2109 (N_2109,N_1860,N_1796);
and U2110 (N_2110,N_1208,N_1143);
or U2111 (N_2111,N_1472,N_1261);
xor U2112 (N_2112,N_1081,N_1322);
nor U2113 (N_2113,N_1321,N_1180);
nand U2114 (N_2114,N_1458,N_1147);
nor U2115 (N_2115,N_1882,N_1803);
nor U2116 (N_2116,N_1610,N_1983);
nor U2117 (N_2117,N_1357,N_1555);
xnor U2118 (N_2118,N_1105,N_1126);
nor U2119 (N_2119,N_1574,N_1447);
nand U2120 (N_2120,N_1212,N_1130);
or U2121 (N_2121,N_1486,N_1592);
or U2122 (N_2122,N_1096,N_1389);
nor U2123 (N_2123,N_1127,N_1113);
nand U2124 (N_2124,N_1957,N_1210);
nor U2125 (N_2125,N_1171,N_1228);
or U2126 (N_2126,N_1585,N_1702);
and U2127 (N_2127,N_1538,N_1044);
and U2128 (N_2128,N_1751,N_1429);
or U2129 (N_2129,N_1192,N_1139);
nor U2130 (N_2130,N_1661,N_1972);
xnor U2131 (N_2131,N_1441,N_1021);
nand U2132 (N_2132,N_1289,N_1026);
xor U2133 (N_2133,N_1237,N_1780);
and U2134 (N_2134,N_1691,N_1885);
xor U2135 (N_2135,N_1720,N_1643);
and U2136 (N_2136,N_1998,N_1288);
xor U2137 (N_2137,N_1590,N_1975);
nor U2138 (N_2138,N_1039,N_1282);
xnor U2139 (N_2139,N_1639,N_1625);
xnor U2140 (N_2140,N_1224,N_1138);
and U2141 (N_2141,N_1658,N_1506);
nand U2142 (N_2142,N_1879,N_1987);
and U2143 (N_2143,N_1226,N_1755);
and U2144 (N_2144,N_1276,N_1685);
nand U2145 (N_2145,N_1563,N_1309);
and U2146 (N_2146,N_1571,N_1009);
and U2147 (N_2147,N_1000,N_1498);
nor U2148 (N_2148,N_1870,N_1400);
and U2149 (N_2149,N_1204,N_1758);
and U2150 (N_2150,N_1095,N_1199);
and U2151 (N_2151,N_1722,N_1230);
xnor U2152 (N_2152,N_1352,N_1724);
and U2153 (N_2153,N_1388,N_1031);
nand U2154 (N_2154,N_1012,N_1097);
xnor U2155 (N_2155,N_1710,N_1402);
and U2156 (N_2156,N_1917,N_1446);
nand U2157 (N_2157,N_1512,N_1117);
and U2158 (N_2158,N_1674,N_1287);
xor U2159 (N_2159,N_1684,N_1198);
or U2160 (N_2160,N_1540,N_1845);
and U2161 (N_2161,N_1331,N_1295);
nor U2162 (N_2162,N_1347,N_1734);
nor U2163 (N_2163,N_1487,N_1345);
xor U2164 (N_2164,N_1010,N_1602);
nor U2165 (N_2165,N_1509,N_1683);
and U2166 (N_2166,N_1971,N_1313);
nand U2167 (N_2167,N_1534,N_1053);
nand U2168 (N_2168,N_1881,N_1209);
xor U2169 (N_2169,N_1537,N_1851);
nand U2170 (N_2170,N_1891,N_1886);
and U2171 (N_2171,N_1707,N_1580);
nand U2172 (N_2172,N_1123,N_1587);
nor U2173 (N_2173,N_1514,N_1910);
or U2174 (N_2174,N_1638,N_1717);
nor U2175 (N_2175,N_1430,N_1363);
nand U2176 (N_2176,N_1759,N_1725);
and U2177 (N_2177,N_1837,N_1516);
nor U2178 (N_2178,N_1552,N_1170);
or U2179 (N_2179,N_1594,N_1640);
and U2180 (N_2180,N_1907,N_1630);
nor U2181 (N_2181,N_1766,N_1203);
or U2182 (N_2182,N_1320,N_1883);
or U2183 (N_2183,N_1715,N_1871);
xnor U2184 (N_2184,N_1562,N_1556);
or U2185 (N_2185,N_1692,N_1281);
and U2186 (N_2186,N_1219,N_1124);
or U2187 (N_2187,N_1669,N_1664);
or U2188 (N_2188,N_1054,N_1190);
nor U2189 (N_2189,N_1898,N_1262);
or U2190 (N_2190,N_1335,N_1179);
nor U2191 (N_2191,N_1848,N_1711);
xnor U2192 (N_2192,N_1992,N_1014);
nand U2193 (N_2193,N_1712,N_1056);
or U2194 (N_2194,N_1572,N_1989);
and U2195 (N_2195,N_1635,N_1386);
xnor U2196 (N_2196,N_1673,N_1155);
and U2197 (N_2197,N_1764,N_1726);
or U2198 (N_2198,N_1263,N_1600);
or U2199 (N_2199,N_1604,N_1951);
xnor U2200 (N_2200,N_1812,N_1696);
or U2201 (N_2201,N_1908,N_1618);
nand U2202 (N_2202,N_1488,N_1248);
xnor U2203 (N_2203,N_1340,N_1231);
or U2204 (N_2204,N_1432,N_1390);
nand U2205 (N_2205,N_1536,N_1076);
xnor U2206 (N_2206,N_1036,N_1062);
and U2207 (N_2207,N_1521,N_1375);
or U2208 (N_2208,N_1087,N_1164);
nand U2209 (N_2209,N_1840,N_1121);
nand U2210 (N_2210,N_1924,N_1651);
or U2211 (N_2211,N_1752,N_1069);
xnor U2212 (N_2212,N_1413,N_1847);
and U2213 (N_2213,N_1510,N_1465);
xor U2214 (N_2214,N_1763,N_1730);
xor U2215 (N_2215,N_1900,N_1916);
and U2216 (N_2216,N_1743,N_1381);
and U2217 (N_2217,N_1452,N_1831);
xnor U2218 (N_2218,N_1469,N_1660);
xor U2219 (N_2219,N_1890,N_1115);
nor U2220 (N_2220,N_1682,N_1937);
and U2221 (N_2221,N_1619,N_1169);
nand U2222 (N_2222,N_1541,N_1611);
nand U2223 (N_2223,N_1997,N_1305);
nor U2224 (N_2224,N_1066,N_1943);
xnor U2225 (N_2225,N_1740,N_1699);
nor U2226 (N_2226,N_1187,N_1995);
or U2227 (N_2227,N_1818,N_1395);
nand U2228 (N_2228,N_1868,N_1233);
or U2229 (N_2229,N_1786,N_1011);
nor U2230 (N_2230,N_1246,N_1116);
or U2231 (N_2231,N_1020,N_1166);
xnor U2232 (N_2232,N_1858,N_1626);
and U2233 (N_2233,N_1264,N_1084);
xor U2234 (N_2234,N_1359,N_1852);
or U2235 (N_2235,N_1649,N_1560);
and U2236 (N_2236,N_1349,N_1930);
nor U2237 (N_2237,N_1965,N_1050);
or U2238 (N_2238,N_1302,N_1109);
and U2239 (N_2239,N_1424,N_1431);
nor U2240 (N_2240,N_1259,N_1667);
or U2241 (N_2241,N_1677,N_1426);
xnor U2242 (N_2242,N_1200,N_1194);
and U2243 (N_2243,N_1168,N_1745);
and U2244 (N_2244,N_1823,N_1756);
nand U2245 (N_2245,N_1222,N_1558);
xnor U2246 (N_2246,N_1709,N_1636);
nor U2247 (N_2247,N_1034,N_1047);
nor U2248 (N_2248,N_1633,N_1396);
or U2249 (N_2249,N_1588,N_1731);
nand U2250 (N_2250,N_1675,N_1581);
or U2251 (N_2251,N_1889,N_1861);
or U2252 (N_2252,N_1944,N_1269);
or U2253 (N_2253,N_1182,N_1028);
and U2254 (N_2254,N_1531,N_1423);
nand U2255 (N_2255,N_1577,N_1846);
and U2256 (N_2256,N_1872,N_1002);
and U2257 (N_2257,N_1593,N_1491);
or U2258 (N_2258,N_1654,N_1921);
xnor U2259 (N_2259,N_1415,N_1942);
and U2260 (N_2260,N_1267,N_1901);
or U2261 (N_2261,N_1824,N_1460);
xor U2262 (N_2262,N_1813,N_1202);
nor U2263 (N_2263,N_1788,N_1969);
or U2264 (N_2264,N_1976,N_1526);
and U2265 (N_2265,N_1817,N_1374);
nor U2266 (N_2266,N_1158,N_1701);
nand U2267 (N_2267,N_1440,N_1175);
and U2268 (N_2268,N_1136,N_1771);
nand U2269 (N_2269,N_1255,N_1839);
or U2270 (N_2270,N_1232,N_1754);
and U2271 (N_2271,N_1548,N_1567);
nor U2272 (N_2272,N_1913,N_1250);
nand U2273 (N_2273,N_1829,N_1380);
nor U2274 (N_2274,N_1994,N_1744);
nand U2275 (N_2275,N_1819,N_1727);
xor U2276 (N_2276,N_1775,N_1271);
xor U2277 (N_2277,N_1003,N_1528);
nor U2278 (N_2278,N_1104,N_1535);
or U2279 (N_2279,N_1694,N_1832);
or U2280 (N_2280,N_1438,N_1079);
and U2281 (N_2281,N_1850,N_1118);
xnor U2282 (N_2282,N_1403,N_1365);
and U2283 (N_2283,N_1785,N_1088);
xnor U2284 (N_2284,N_1905,N_1532);
nand U2285 (N_2285,N_1570,N_1317);
or U2286 (N_2286,N_1733,N_1807);
nor U2287 (N_2287,N_1455,N_1973);
or U2288 (N_2288,N_1037,N_1892);
xor U2289 (N_2289,N_1663,N_1826);
and U2290 (N_2290,N_1433,N_1236);
and U2291 (N_2291,N_1211,N_1855);
nor U2292 (N_2292,N_1351,N_1545);
and U2293 (N_2293,N_1533,N_1367);
or U2294 (N_2294,N_1191,N_1984);
and U2295 (N_2295,N_1544,N_1330);
nand U2296 (N_2296,N_1450,N_1525);
and U2297 (N_2297,N_1098,N_1642);
and U2298 (N_2298,N_1101,N_1929);
or U2299 (N_2299,N_1777,N_1376);
nand U2300 (N_2300,N_1484,N_1299);
and U2301 (N_2301,N_1476,N_1620);
xor U2302 (N_2302,N_1713,N_1238);
and U2303 (N_2303,N_1379,N_1294);
nor U2304 (N_2304,N_1794,N_1043);
xnor U2305 (N_2305,N_1355,N_1300);
nor U2306 (N_2306,N_1427,N_1946);
nand U2307 (N_2307,N_1781,N_1797);
or U2308 (N_2308,N_1052,N_1999);
nand U2309 (N_2309,N_1704,N_1495);
xnor U2310 (N_2310,N_1954,N_1480);
xor U2311 (N_2311,N_1128,N_1140);
and U2312 (N_2312,N_1679,N_1145);
or U2313 (N_2313,N_1705,N_1884);
nand U2314 (N_2314,N_1214,N_1914);
nand U2315 (N_2315,N_1283,N_1670);
or U2316 (N_2316,N_1583,N_1893);
and U2317 (N_2317,N_1185,N_1737);
and U2318 (N_2318,N_1436,N_1967);
and U2319 (N_2319,N_1083,N_1167);
nand U2320 (N_2320,N_1844,N_1529);
and U2321 (N_2321,N_1931,N_1836);
nor U2322 (N_2322,N_1718,N_1500);
nor U2323 (N_2323,N_1815,N_1073);
or U2324 (N_2324,N_1067,N_1405);
nand U2325 (N_2325,N_1622,N_1314);
xnor U2326 (N_2326,N_1760,N_1697);
xnor U2327 (N_2327,N_1055,N_1018);
nand U2328 (N_2328,N_1920,N_1791);
nor U2329 (N_2329,N_1059,N_1765);
or U2330 (N_2330,N_1769,N_1477);
or U2331 (N_2331,N_1225,N_1048);
xnor U2332 (N_2332,N_1270,N_1926);
xnor U2333 (N_2333,N_1628,N_1561);
nand U2334 (N_2334,N_1517,N_1234);
nor U2335 (N_2335,N_1614,N_1129);
and U2336 (N_2336,N_1421,N_1008);
or U2337 (N_2337,N_1493,N_1094);
nand U2338 (N_2338,N_1564,N_1597);
or U2339 (N_2339,N_1919,N_1184);
nand U2340 (N_2340,N_1963,N_1051);
nor U2341 (N_2341,N_1221,N_1414);
nand U2342 (N_2342,N_1546,N_1382);
nand U2343 (N_2343,N_1162,N_1782);
or U2344 (N_2344,N_1207,N_1035);
or U2345 (N_2345,N_1280,N_1557);
or U2346 (N_2346,N_1195,N_1646);
or U2347 (N_2347,N_1030,N_1877);
and U2348 (N_2348,N_1193,N_1644);
nor U2349 (N_2349,N_1605,N_1277);
nand U2350 (N_2350,N_1948,N_1974);
nand U2351 (N_2351,N_1822,N_1551);
or U2352 (N_2352,N_1862,N_1841);
or U2353 (N_2353,N_1393,N_1964);
xor U2354 (N_2354,N_1197,N_1220);
and U2355 (N_2355,N_1107,N_1196);
xnor U2356 (N_2356,N_1163,N_1767);
xnor U2357 (N_2357,N_1077,N_1111);
or U2358 (N_2358,N_1873,N_1596);
nand U2359 (N_2359,N_1108,N_1297);
xnor U2360 (N_2360,N_1659,N_1568);
and U2361 (N_2361,N_1384,N_1598);
nor U2362 (N_2362,N_1789,N_1165);
and U2363 (N_2363,N_1327,N_1497);
nor U2364 (N_2364,N_1451,N_1986);
and U2365 (N_2365,N_1530,N_1736);
nor U2366 (N_2366,N_1324,N_1772);
nor U2367 (N_2367,N_1615,N_1150);
or U2368 (N_2368,N_1227,N_1385);
nor U2369 (N_2369,N_1853,N_1372);
xnor U2370 (N_2370,N_1176,N_1714);
nor U2371 (N_2371,N_1099,N_1040);
nand U2372 (N_2372,N_1337,N_1045);
or U2373 (N_2373,N_1368,N_1311);
and U2374 (N_2374,N_1936,N_1023);
nand U2375 (N_2375,N_1689,N_1336);
nor U2376 (N_2376,N_1142,N_1470);
and U2377 (N_2377,N_1064,N_1814);
nor U2378 (N_2378,N_1996,N_1678);
nor U2379 (N_2379,N_1483,N_1783);
xnor U2380 (N_2380,N_1778,N_1956);
nor U2381 (N_2381,N_1981,N_1428);
nor U2382 (N_2382,N_1453,N_1332);
nand U2383 (N_2383,N_1776,N_1201);
nand U2384 (N_2384,N_1579,N_1575);
nand U2385 (N_2385,N_1653,N_1906);
or U2386 (N_2386,N_1341,N_1599);
xor U2387 (N_2387,N_1122,N_1985);
xnor U2388 (N_2388,N_1982,N_1417);
or U2389 (N_2389,N_1693,N_1205);
nand U2390 (N_2390,N_1316,N_1650);
nor U2391 (N_2391,N_1810,N_1656);
nand U2392 (N_2392,N_1279,N_1260);
and U2393 (N_2393,N_1206,N_1442);
and U2394 (N_2394,N_1223,N_1795);
nor U2395 (N_2395,N_1178,N_1798);
or U2396 (N_2396,N_1156,N_1923);
or U2397 (N_2397,N_1038,N_1904);
or U2398 (N_2398,N_1348,N_1770);
and U2399 (N_2399,N_1681,N_1085);
nor U2400 (N_2400,N_1304,N_1407);
nor U2401 (N_2401,N_1647,N_1100);
or U2402 (N_2402,N_1448,N_1909);
or U2403 (N_2403,N_1177,N_1241);
or U2404 (N_2404,N_1945,N_1006);
nand U2405 (N_2405,N_1784,N_1899);
xor U2406 (N_2406,N_1338,N_1496);
and U2407 (N_2407,N_1508,N_1058);
or U2408 (N_2408,N_1787,N_1189);
xnor U2409 (N_2409,N_1703,N_1668);
xor U2410 (N_2410,N_1676,N_1371);
nor U2411 (N_2411,N_1990,N_1576);
or U2412 (N_2412,N_1119,N_1750);
xor U2413 (N_2413,N_1595,N_1952);
nor U2414 (N_2414,N_1254,N_1941);
nand U2415 (N_2415,N_1790,N_1520);
and U2416 (N_2416,N_1657,N_1057);
or U2417 (N_2417,N_1666,N_1392);
xnor U2418 (N_2418,N_1024,N_1292);
nand U2419 (N_2419,N_1655,N_1988);
nand U2420 (N_2420,N_1589,N_1272);
xor U2421 (N_2421,N_1318,N_1027);
nor U2422 (N_2422,N_1141,N_1342);
nor U2423 (N_2423,N_1617,N_1445);
and U2424 (N_2424,N_1482,N_1522);
xnor U2425 (N_2425,N_1334,N_1542);
nor U2426 (N_2426,N_1979,N_1489);
nand U2427 (N_2427,N_1621,N_1834);
and U2428 (N_2428,N_1912,N_1333);
xnor U2429 (N_2429,N_1700,N_1838);
and U2430 (N_2430,N_1474,N_1966);
nand U2431 (N_2431,N_1157,N_1842);
or U2432 (N_2432,N_1940,N_1802);
or U2433 (N_2433,N_1112,N_1827);
nand U2434 (N_2434,N_1553,N_1042);
or U2435 (N_2435,N_1761,N_1046);
xnor U2436 (N_2436,N_1449,N_1809);
xor U2437 (N_2437,N_1373,N_1364);
nor U2438 (N_2438,N_1811,N_1799);
or U2439 (N_2439,N_1565,N_1284);
or U2440 (N_2440,N_1137,N_1706);
nor U2441 (N_2441,N_1134,N_1735);
and U2442 (N_2442,N_1499,N_1485);
nor U2443 (N_2443,N_1880,N_1071);
nor U2444 (N_2444,N_1503,N_1863);
nand U2445 (N_2445,N_1603,N_1695);
and U2446 (N_2446,N_1748,N_1742);
nor U2447 (N_2447,N_1471,N_1953);
and U2448 (N_2448,N_1082,N_1800);
nand U2449 (N_2449,N_1686,N_1378);
nor U2450 (N_2450,N_1970,N_1613);
and U2451 (N_2451,N_1894,N_1041);
nand U2452 (N_2452,N_1383,N_1394);
nand U2453 (N_2453,N_1174,N_1939);
nor U2454 (N_2454,N_1456,N_1457);
and U2455 (N_2455,N_1406,N_1464);
nand U2456 (N_2456,N_1554,N_1131);
or U2457 (N_2457,N_1515,N_1410);
and U2458 (N_2458,N_1854,N_1601);
nor U2459 (N_2459,N_1888,N_1268);
nand U2460 (N_2460,N_1479,N_1092);
or U2461 (N_2461,N_1768,N_1354);
and U2462 (N_2462,N_1903,N_1443);
xor U2463 (N_2463,N_1459,N_1377);
nor U2464 (N_2464,N_1015,N_1303);
or U2465 (N_2465,N_1278,N_1501);
and U2466 (N_2466,N_1878,N_1370);
xnor U2467 (N_2467,N_1418,N_1991);
and U2468 (N_2468,N_1217,N_1404);
or U2469 (N_2469,N_1154,N_1399);
nor U2470 (N_2470,N_1369,N_1285);
nor U2471 (N_2471,N_1091,N_1001);
or U2472 (N_2472,N_1257,N_1637);
xnor U2473 (N_2473,N_1950,N_1007);
xnor U2474 (N_2474,N_1816,N_1032);
xnor U2475 (N_2475,N_1078,N_1308);
nand U2476 (N_2476,N_1616,N_1478);
and U2477 (N_2477,N_1746,N_1060);
nand U2478 (N_2478,N_1387,N_1391);
xor U2479 (N_2479,N_1865,N_1821);
nand U2480 (N_2480,N_1949,N_1825);
xnor U2481 (N_2481,N_1343,N_1153);
nand U2482 (N_2482,N_1993,N_1074);
nand U2483 (N_2483,N_1089,N_1315);
and U2484 (N_2484,N_1958,N_1762);
nand U2485 (N_2485,N_1360,N_1897);
nand U2486 (N_2486,N_1437,N_1125);
and U2487 (N_2487,N_1256,N_1932);
nand U2488 (N_2488,N_1835,N_1511);
nand U2489 (N_2489,N_1114,N_1061);
and U2490 (N_2490,N_1461,N_1934);
nand U2491 (N_2491,N_1584,N_1110);
nand U2492 (N_2492,N_1665,N_1022);
nand U2493 (N_2493,N_1298,N_1319);
or U2494 (N_2494,N_1275,N_1504);
nor U2495 (N_2495,N_1606,N_1867);
or U2496 (N_2496,N_1729,N_1741);
and U2497 (N_2497,N_1065,N_1265);
or U2498 (N_2498,N_1475,N_1454);
xor U2499 (N_2499,N_1462,N_1188);
nand U2500 (N_2500,N_1006,N_1100);
or U2501 (N_2501,N_1921,N_1626);
and U2502 (N_2502,N_1581,N_1034);
or U2503 (N_2503,N_1748,N_1200);
or U2504 (N_2504,N_1303,N_1049);
xor U2505 (N_2505,N_1245,N_1920);
xor U2506 (N_2506,N_1249,N_1669);
xnor U2507 (N_2507,N_1789,N_1364);
xnor U2508 (N_2508,N_1030,N_1221);
xor U2509 (N_2509,N_1289,N_1897);
nand U2510 (N_2510,N_1153,N_1130);
nand U2511 (N_2511,N_1374,N_1119);
xor U2512 (N_2512,N_1179,N_1694);
nor U2513 (N_2513,N_1103,N_1926);
xnor U2514 (N_2514,N_1185,N_1640);
and U2515 (N_2515,N_1261,N_1157);
xor U2516 (N_2516,N_1585,N_1537);
and U2517 (N_2517,N_1377,N_1317);
nand U2518 (N_2518,N_1388,N_1806);
xor U2519 (N_2519,N_1068,N_1547);
and U2520 (N_2520,N_1226,N_1962);
or U2521 (N_2521,N_1152,N_1605);
xor U2522 (N_2522,N_1343,N_1364);
and U2523 (N_2523,N_1489,N_1940);
nand U2524 (N_2524,N_1601,N_1792);
or U2525 (N_2525,N_1600,N_1679);
xnor U2526 (N_2526,N_1506,N_1595);
nor U2527 (N_2527,N_1050,N_1490);
or U2528 (N_2528,N_1776,N_1802);
and U2529 (N_2529,N_1481,N_1950);
xnor U2530 (N_2530,N_1598,N_1918);
or U2531 (N_2531,N_1713,N_1221);
nor U2532 (N_2532,N_1335,N_1596);
nand U2533 (N_2533,N_1182,N_1598);
or U2534 (N_2534,N_1657,N_1725);
xnor U2535 (N_2535,N_1055,N_1247);
nand U2536 (N_2536,N_1898,N_1308);
xor U2537 (N_2537,N_1302,N_1787);
and U2538 (N_2538,N_1292,N_1294);
nor U2539 (N_2539,N_1389,N_1590);
or U2540 (N_2540,N_1055,N_1265);
or U2541 (N_2541,N_1411,N_1887);
nor U2542 (N_2542,N_1059,N_1028);
and U2543 (N_2543,N_1026,N_1262);
and U2544 (N_2544,N_1436,N_1499);
nor U2545 (N_2545,N_1908,N_1139);
nor U2546 (N_2546,N_1128,N_1924);
and U2547 (N_2547,N_1404,N_1904);
and U2548 (N_2548,N_1306,N_1800);
nand U2549 (N_2549,N_1987,N_1795);
or U2550 (N_2550,N_1129,N_1187);
xnor U2551 (N_2551,N_1896,N_1820);
or U2552 (N_2552,N_1892,N_1113);
xnor U2553 (N_2553,N_1082,N_1496);
or U2554 (N_2554,N_1628,N_1347);
and U2555 (N_2555,N_1249,N_1198);
xor U2556 (N_2556,N_1213,N_1710);
or U2557 (N_2557,N_1962,N_1220);
and U2558 (N_2558,N_1247,N_1488);
and U2559 (N_2559,N_1525,N_1474);
or U2560 (N_2560,N_1823,N_1714);
xor U2561 (N_2561,N_1405,N_1647);
nor U2562 (N_2562,N_1133,N_1548);
nor U2563 (N_2563,N_1914,N_1808);
nor U2564 (N_2564,N_1646,N_1323);
nand U2565 (N_2565,N_1634,N_1720);
nor U2566 (N_2566,N_1659,N_1142);
and U2567 (N_2567,N_1387,N_1170);
nor U2568 (N_2568,N_1263,N_1445);
nand U2569 (N_2569,N_1906,N_1268);
and U2570 (N_2570,N_1532,N_1573);
and U2571 (N_2571,N_1533,N_1386);
xnor U2572 (N_2572,N_1796,N_1808);
and U2573 (N_2573,N_1659,N_1930);
and U2574 (N_2574,N_1595,N_1448);
xor U2575 (N_2575,N_1727,N_1635);
nor U2576 (N_2576,N_1294,N_1685);
nand U2577 (N_2577,N_1132,N_1877);
nor U2578 (N_2578,N_1628,N_1721);
and U2579 (N_2579,N_1593,N_1300);
nand U2580 (N_2580,N_1939,N_1896);
and U2581 (N_2581,N_1886,N_1458);
nand U2582 (N_2582,N_1040,N_1133);
nand U2583 (N_2583,N_1538,N_1215);
xnor U2584 (N_2584,N_1177,N_1565);
or U2585 (N_2585,N_1268,N_1869);
nand U2586 (N_2586,N_1114,N_1432);
and U2587 (N_2587,N_1867,N_1982);
or U2588 (N_2588,N_1631,N_1257);
and U2589 (N_2589,N_1192,N_1526);
nor U2590 (N_2590,N_1722,N_1347);
nor U2591 (N_2591,N_1652,N_1115);
nor U2592 (N_2592,N_1702,N_1959);
nand U2593 (N_2593,N_1724,N_1890);
nand U2594 (N_2594,N_1340,N_1121);
xnor U2595 (N_2595,N_1954,N_1148);
nand U2596 (N_2596,N_1380,N_1464);
and U2597 (N_2597,N_1143,N_1651);
or U2598 (N_2598,N_1062,N_1817);
or U2599 (N_2599,N_1724,N_1637);
nor U2600 (N_2600,N_1551,N_1922);
and U2601 (N_2601,N_1426,N_1189);
and U2602 (N_2602,N_1422,N_1053);
xor U2603 (N_2603,N_1938,N_1593);
nand U2604 (N_2604,N_1424,N_1062);
nand U2605 (N_2605,N_1162,N_1170);
xnor U2606 (N_2606,N_1937,N_1916);
xor U2607 (N_2607,N_1901,N_1647);
nor U2608 (N_2608,N_1138,N_1793);
xor U2609 (N_2609,N_1336,N_1942);
nand U2610 (N_2610,N_1284,N_1946);
or U2611 (N_2611,N_1698,N_1942);
and U2612 (N_2612,N_1924,N_1270);
or U2613 (N_2613,N_1024,N_1290);
or U2614 (N_2614,N_1300,N_1113);
nor U2615 (N_2615,N_1468,N_1953);
xnor U2616 (N_2616,N_1006,N_1459);
xor U2617 (N_2617,N_1638,N_1944);
nand U2618 (N_2618,N_1911,N_1236);
nor U2619 (N_2619,N_1247,N_1328);
nand U2620 (N_2620,N_1183,N_1803);
nand U2621 (N_2621,N_1702,N_1018);
and U2622 (N_2622,N_1752,N_1393);
and U2623 (N_2623,N_1155,N_1220);
xor U2624 (N_2624,N_1453,N_1648);
and U2625 (N_2625,N_1516,N_1441);
xor U2626 (N_2626,N_1830,N_1793);
or U2627 (N_2627,N_1345,N_1392);
nand U2628 (N_2628,N_1261,N_1317);
nor U2629 (N_2629,N_1569,N_1099);
nor U2630 (N_2630,N_1945,N_1185);
and U2631 (N_2631,N_1621,N_1133);
nor U2632 (N_2632,N_1739,N_1596);
nor U2633 (N_2633,N_1841,N_1523);
and U2634 (N_2634,N_1956,N_1768);
or U2635 (N_2635,N_1516,N_1566);
nand U2636 (N_2636,N_1903,N_1943);
nand U2637 (N_2637,N_1751,N_1778);
nand U2638 (N_2638,N_1414,N_1861);
or U2639 (N_2639,N_1984,N_1858);
nand U2640 (N_2640,N_1409,N_1200);
or U2641 (N_2641,N_1049,N_1698);
or U2642 (N_2642,N_1661,N_1695);
or U2643 (N_2643,N_1868,N_1436);
and U2644 (N_2644,N_1899,N_1766);
nand U2645 (N_2645,N_1898,N_1766);
and U2646 (N_2646,N_1411,N_1760);
or U2647 (N_2647,N_1535,N_1500);
and U2648 (N_2648,N_1750,N_1055);
or U2649 (N_2649,N_1882,N_1155);
and U2650 (N_2650,N_1195,N_1027);
nand U2651 (N_2651,N_1989,N_1410);
nand U2652 (N_2652,N_1879,N_1846);
xor U2653 (N_2653,N_1561,N_1304);
nand U2654 (N_2654,N_1087,N_1955);
nor U2655 (N_2655,N_1894,N_1950);
nor U2656 (N_2656,N_1815,N_1044);
xor U2657 (N_2657,N_1229,N_1427);
or U2658 (N_2658,N_1240,N_1536);
xnor U2659 (N_2659,N_1180,N_1565);
and U2660 (N_2660,N_1553,N_1196);
nand U2661 (N_2661,N_1087,N_1222);
nand U2662 (N_2662,N_1730,N_1642);
or U2663 (N_2663,N_1386,N_1107);
or U2664 (N_2664,N_1780,N_1527);
or U2665 (N_2665,N_1018,N_1991);
nor U2666 (N_2666,N_1288,N_1166);
or U2667 (N_2667,N_1854,N_1728);
xnor U2668 (N_2668,N_1313,N_1838);
nand U2669 (N_2669,N_1502,N_1348);
nor U2670 (N_2670,N_1396,N_1474);
or U2671 (N_2671,N_1148,N_1906);
nand U2672 (N_2672,N_1583,N_1728);
nor U2673 (N_2673,N_1270,N_1993);
nand U2674 (N_2674,N_1898,N_1214);
nor U2675 (N_2675,N_1569,N_1237);
xor U2676 (N_2676,N_1484,N_1963);
nor U2677 (N_2677,N_1925,N_1524);
xnor U2678 (N_2678,N_1208,N_1980);
nor U2679 (N_2679,N_1551,N_1197);
nand U2680 (N_2680,N_1827,N_1229);
nor U2681 (N_2681,N_1021,N_1420);
and U2682 (N_2682,N_1830,N_1757);
nor U2683 (N_2683,N_1981,N_1592);
nor U2684 (N_2684,N_1503,N_1763);
or U2685 (N_2685,N_1154,N_1139);
nand U2686 (N_2686,N_1774,N_1611);
or U2687 (N_2687,N_1350,N_1184);
and U2688 (N_2688,N_1562,N_1664);
xor U2689 (N_2689,N_1637,N_1099);
nor U2690 (N_2690,N_1288,N_1117);
and U2691 (N_2691,N_1309,N_1928);
xnor U2692 (N_2692,N_1664,N_1581);
nor U2693 (N_2693,N_1280,N_1965);
and U2694 (N_2694,N_1534,N_1381);
nand U2695 (N_2695,N_1221,N_1680);
and U2696 (N_2696,N_1831,N_1303);
nor U2697 (N_2697,N_1667,N_1727);
and U2698 (N_2698,N_1211,N_1156);
xnor U2699 (N_2699,N_1537,N_1616);
nand U2700 (N_2700,N_1721,N_1509);
nor U2701 (N_2701,N_1259,N_1476);
nand U2702 (N_2702,N_1545,N_1014);
and U2703 (N_2703,N_1669,N_1521);
xnor U2704 (N_2704,N_1009,N_1935);
xor U2705 (N_2705,N_1202,N_1426);
nand U2706 (N_2706,N_1187,N_1083);
and U2707 (N_2707,N_1376,N_1451);
nor U2708 (N_2708,N_1385,N_1092);
nor U2709 (N_2709,N_1010,N_1341);
nand U2710 (N_2710,N_1171,N_1498);
nor U2711 (N_2711,N_1965,N_1433);
or U2712 (N_2712,N_1188,N_1898);
nand U2713 (N_2713,N_1799,N_1543);
and U2714 (N_2714,N_1447,N_1686);
nand U2715 (N_2715,N_1561,N_1322);
nand U2716 (N_2716,N_1870,N_1927);
nor U2717 (N_2717,N_1452,N_1538);
xnor U2718 (N_2718,N_1614,N_1916);
or U2719 (N_2719,N_1974,N_1281);
nand U2720 (N_2720,N_1646,N_1748);
and U2721 (N_2721,N_1237,N_1241);
or U2722 (N_2722,N_1835,N_1889);
nor U2723 (N_2723,N_1840,N_1709);
and U2724 (N_2724,N_1701,N_1270);
or U2725 (N_2725,N_1384,N_1250);
or U2726 (N_2726,N_1651,N_1929);
or U2727 (N_2727,N_1219,N_1526);
nand U2728 (N_2728,N_1260,N_1197);
nand U2729 (N_2729,N_1492,N_1605);
xnor U2730 (N_2730,N_1073,N_1695);
or U2731 (N_2731,N_1600,N_1067);
nor U2732 (N_2732,N_1006,N_1067);
and U2733 (N_2733,N_1102,N_1123);
nand U2734 (N_2734,N_1202,N_1634);
or U2735 (N_2735,N_1770,N_1441);
and U2736 (N_2736,N_1742,N_1262);
xor U2737 (N_2737,N_1024,N_1534);
or U2738 (N_2738,N_1741,N_1557);
and U2739 (N_2739,N_1199,N_1823);
xnor U2740 (N_2740,N_1221,N_1555);
nor U2741 (N_2741,N_1538,N_1890);
xnor U2742 (N_2742,N_1762,N_1527);
or U2743 (N_2743,N_1722,N_1556);
or U2744 (N_2744,N_1999,N_1278);
nor U2745 (N_2745,N_1827,N_1712);
or U2746 (N_2746,N_1428,N_1364);
nand U2747 (N_2747,N_1261,N_1798);
nor U2748 (N_2748,N_1861,N_1589);
nor U2749 (N_2749,N_1474,N_1324);
and U2750 (N_2750,N_1127,N_1913);
xor U2751 (N_2751,N_1660,N_1493);
nor U2752 (N_2752,N_1793,N_1131);
or U2753 (N_2753,N_1196,N_1632);
or U2754 (N_2754,N_1833,N_1971);
nand U2755 (N_2755,N_1400,N_1862);
or U2756 (N_2756,N_1572,N_1071);
or U2757 (N_2757,N_1272,N_1563);
and U2758 (N_2758,N_1856,N_1119);
xor U2759 (N_2759,N_1554,N_1051);
or U2760 (N_2760,N_1387,N_1231);
and U2761 (N_2761,N_1298,N_1376);
and U2762 (N_2762,N_1336,N_1776);
nor U2763 (N_2763,N_1576,N_1627);
or U2764 (N_2764,N_1839,N_1822);
nor U2765 (N_2765,N_1510,N_1867);
and U2766 (N_2766,N_1357,N_1085);
and U2767 (N_2767,N_1781,N_1504);
nor U2768 (N_2768,N_1662,N_1005);
xor U2769 (N_2769,N_1218,N_1137);
nand U2770 (N_2770,N_1203,N_1825);
or U2771 (N_2771,N_1661,N_1074);
nand U2772 (N_2772,N_1093,N_1727);
nand U2773 (N_2773,N_1336,N_1518);
nand U2774 (N_2774,N_1557,N_1617);
xnor U2775 (N_2775,N_1583,N_1956);
or U2776 (N_2776,N_1304,N_1946);
xor U2777 (N_2777,N_1369,N_1878);
nand U2778 (N_2778,N_1284,N_1160);
xnor U2779 (N_2779,N_1965,N_1295);
and U2780 (N_2780,N_1518,N_1750);
nand U2781 (N_2781,N_1676,N_1658);
or U2782 (N_2782,N_1284,N_1697);
nor U2783 (N_2783,N_1572,N_1031);
nor U2784 (N_2784,N_1146,N_1597);
and U2785 (N_2785,N_1716,N_1001);
xor U2786 (N_2786,N_1962,N_1173);
or U2787 (N_2787,N_1083,N_1441);
nand U2788 (N_2788,N_1626,N_1279);
xnor U2789 (N_2789,N_1455,N_1157);
or U2790 (N_2790,N_1443,N_1858);
or U2791 (N_2791,N_1537,N_1539);
or U2792 (N_2792,N_1875,N_1448);
xor U2793 (N_2793,N_1699,N_1601);
or U2794 (N_2794,N_1640,N_1191);
xor U2795 (N_2795,N_1692,N_1682);
nor U2796 (N_2796,N_1878,N_1338);
nand U2797 (N_2797,N_1118,N_1982);
nor U2798 (N_2798,N_1951,N_1978);
or U2799 (N_2799,N_1469,N_1623);
nor U2800 (N_2800,N_1689,N_1988);
nor U2801 (N_2801,N_1208,N_1693);
nand U2802 (N_2802,N_1903,N_1113);
nand U2803 (N_2803,N_1945,N_1451);
xnor U2804 (N_2804,N_1692,N_1018);
nor U2805 (N_2805,N_1244,N_1768);
xor U2806 (N_2806,N_1949,N_1499);
nor U2807 (N_2807,N_1390,N_1902);
and U2808 (N_2808,N_1048,N_1355);
xor U2809 (N_2809,N_1376,N_1827);
xnor U2810 (N_2810,N_1732,N_1541);
and U2811 (N_2811,N_1403,N_1487);
and U2812 (N_2812,N_1195,N_1351);
xor U2813 (N_2813,N_1756,N_1905);
or U2814 (N_2814,N_1538,N_1175);
or U2815 (N_2815,N_1942,N_1485);
xor U2816 (N_2816,N_1773,N_1713);
and U2817 (N_2817,N_1696,N_1603);
nor U2818 (N_2818,N_1527,N_1064);
and U2819 (N_2819,N_1736,N_1021);
and U2820 (N_2820,N_1024,N_1949);
or U2821 (N_2821,N_1833,N_1609);
nand U2822 (N_2822,N_1768,N_1006);
nand U2823 (N_2823,N_1763,N_1585);
nor U2824 (N_2824,N_1050,N_1722);
and U2825 (N_2825,N_1460,N_1924);
nor U2826 (N_2826,N_1930,N_1026);
or U2827 (N_2827,N_1384,N_1549);
nor U2828 (N_2828,N_1799,N_1042);
nand U2829 (N_2829,N_1898,N_1057);
nand U2830 (N_2830,N_1782,N_1099);
nand U2831 (N_2831,N_1166,N_1173);
or U2832 (N_2832,N_1788,N_1122);
or U2833 (N_2833,N_1313,N_1113);
nor U2834 (N_2834,N_1773,N_1769);
and U2835 (N_2835,N_1266,N_1476);
nor U2836 (N_2836,N_1356,N_1433);
nor U2837 (N_2837,N_1051,N_1781);
nor U2838 (N_2838,N_1975,N_1182);
nor U2839 (N_2839,N_1682,N_1534);
xor U2840 (N_2840,N_1206,N_1083);
or U2841 (N_2841,N_1634,N_1892);
and U2842 (N_2842,N_1251,N_1788);
nor U2843 (N_2843,N_1500,N_1797);
nor U2844 (N_2844,N_1904,N_1612);
nand U2845 (N_2845,N_1546,N_1277);
and U2846 (N_2846,N_1012,N_1203);
xnor U2847 (N_2847,N_1435,N_1412);
nor U2848 (N_2848,N_1446,N_1990);
or U2849 (N_2849,N_1252,N_1467);
xor U2850 (N_2850,N_1029,N_1215);
nand U2851 (N_2851,N_1840,N_1320);
nand U2852 (N_2852,N_1559,N_1330);
nand U2853 (N_2853,N_1396,N_1783);
nor U2854 (N_2854,N_1992,N_1520);
nor U2855 (N_2855,N_1343,N_1895);
nor U2856 (N_2856,N_1735,N_1066);
nor U2857 (N_2857,N_1597,N_1733);
nor U2858 (N_2858,N_1997,N_1125);
or U2859 (N_2859,N_1043,N_1609);
nor U2860 (N_2860,N_1907,N_1049);
or U2861 (N_2861,N_1470,N_1791);
xnor U2862 (N_2862,N_1625,N_1751);
and U2863 (N_2863,N_1203,N_1264);
or U2864 (N_2864,N_1680,N_1777);
nand U2865 (N_2865,N_1258,N_1080);
nand U2866 (N_2866,N_1249,N_1781);
nor U2867 (N_2867,N_1416,N_1921);
nand U2868 (N_2868,N_1996,N_1942);
nor U2869 (N_2869,N_1976,N_1249);
and U2870 (N_2870,N_1509,N_1016);
and U2871 (N_2871,N_1552,N_1887);
and U2872 (N_2872,N_1736,N_1433);
nand U2873 (N_2873,N_1878,N_1528);
or U2874 (N_2874,N_1264,N_1886);
and U2875 (N_2875,N_1279,N_1199);
nand U2876 (N_2876,N_1035,N_1792);
or U2877 (N_2877,N_1952,N_1947);
nor U2878 (N_2878,N_1640,N_1171);
nand U2879 (N_2879,N_1491,N_1311);
and U2880 (N_2880,N_1426,N_1850);
and U2881 (N_2881,N_1419,N_1121);
or U2882 (N_2882,N_1757,N_1548);
nor U2883 (N_2883,N_1763,N_1483);
nand U2884 (N_2884,N_1563,N_1388);
nor U2885 (N_2885,N_1296,N_1327);
nand U2886 (N_2886,N_1912,N_1346);
and U2887 (N_2887,N_1603,N_1168);
nor U2888 (N_2888,N_1656,N_1632);
nand U2889 (N_2889,N_1166,N_1201);
and U2890 (N_2890,N_1786,N_1430);
and U2891 (N_2891,N_1936,N_1967);
and U2892 (N_2892,N_1402,N_1314);
nand U2893 (N_2893,N_1054,N_1322);
nand U2894 (N_2894,N_1983,N_1809);
nor U2895 (N_2895,N_1412,N_1713);
nor U2896 (N_2896,N_1647,N_1447);
nor U2897 (N_2897,N_1334,N_1431);
and U2898 (N_2898,N_1959,N_1151);
nor U2899 (N_2899,N_1215,N_1919);
nor U2900 (N_2900,N_1866,N_1311);
and U2901 (N_2901,N_1744,N_1688);
nor U2902 (N_2902,N_1411,N_1281);
nand U2903 (N_2903,N_1275,N_1589);
and U2904 (N_2904,N_1741,N_1329);
nor U2905 (N_2905,N_1549,N_1431);
xor U2906 (N_2906,N_1276,N_1871);
xor U2907 (N_2907,N_1818,N_1656);
and U2908 (N_2908,N_1215,N_1192);
and U2909 (N_2909,N_1837,N_1037);
and U2910 (N_2910,N_1593,N_1093);
xor U2911 (N_2911,N_1828,N_1069);
and U2912 (N_2912,N_1748,N_1321);
nand U2913 (N_2913,N_1031,N_1479);
nor U2914 (N_2914,N_1942,N_1507);
or U2915 (N_2915,N_1449,N_1348);
or U2916 (N_2916,N_1286,N_1862);
nor U2917 (N_2917,N_1363,N_1569);
and U2918 (N_2918,N_1956,N_1358);
nand U2919 (N_2919,N_1923,N_1549);
nand U2920 (N_2920,N_1379,N_1433);
and U2921 (N_2921,N_1251,N_1241);
xnor U2922 (N_2922,N_1510,N_1593);
xnor U2923 (N_2923,N_1566,N_1967);
nand U2924 (N_2924,N_1532,N_1446);
xnor U2925 (N_2925,N_1322,N_1916);
nand U2926 (N_2926,N_1965,N_1071);
xnor U2927 (N_2927,N_1654,N_1058);
xnor U2928 (N_2928,N_1140,N_1900);
nand U2929 (N_2929,N_1486,N_1287);
and U2930 (N_2930,N_1968,N_1676);
nand U2931 (N_2931,N_1400,N_1307);
and U2932 (N_2932,N_1598,N_1624);
nand U2933 (N_2933,N_1963,N_1983);
xor U2934 (N_2934,N_1371,N_1751);
xor U2935 (N_2935,N_1378,N_1964);
or U2936 (N_2936,N_1125,N_1341);
or U2937 (N_2937,N_1195,N_1925);
nor U2938 (N_2938,N_1349,N_1013);
and U2939 (N_2939,N_1198,N_1489);
nor U2940 (N_2940,N_1123,N_1367);
or U2941 (N_2941,N_1981,N_1208);
nand U2942 (N_2942,N_1071,N_1450);
nor U2943 (N_2943,N_1474,N_1643);
or U2944 (N_2944,N_1941,N_1574);
xnor U2945 (N_2945,N_1669,N_1511);
nor U2946 (N_2946,N_1312,N_1410);
nand U2947 (N_2947,N_1397,N_1969);
and U2948 (N_2948,N_1146,N_1327);
or U2949 (N_2949,N_1745,N_1934);
and U2950 (N_2950,N_1728,N_1935);
or U2951 (N_2951,N_1807,N_1933);
nand U2952 (N_2952,N_1410,N_1959);
xnor U2953 (N_2953,N_1712,N_1438);
and U2954 (N_2954,N_1404,N_1512);
nor U2955 (N_2955,N_1405,N_1733);
xor U2956 (N_2956,N_1432,N_1089);
nor U2957 (N_2957,N_1658,N_1938);
nand U2958 (N_2958,N_1063,N_1059);
and U2959 (N_2959,N_1550,N_1478);
xor U2960 (N_2960,N_1860,N_1514);
nor U2961 (N_2961,N_1967,N_1872);
or U2962 (N_2962,N_1022,N_1037);
or U2963 (N_2963,N_1474,N_1786);
or U2964 (N_2964,N_1022,N_1687);
nand U2965 (N_2965,N_1769,N_1214);
nor U2966 (N_2966,N_1613,N_1193);
and U2967 (N_2967,N_1735,N_1304);
and U2968 (N_2968,N_1486,N_1448);
or U2969 (N_2969,N_1878,N_1512);
nand U2970 (N_2970,N_1109,N_1832);
xnor U2971 (N_2971,N_1487,N_1189);
nor U2972 (N_2972,N_1978,N_1852);
and U2973 (N_2973,N_1543,N_1284);
or U2974 (N_2974,N_1752,N_1473);
and U2975 (N_2975,N_1481,N_1311);
xnor U2976 (N_2976,N_1477,N_1929);
nand U2977 (N_2977,N_1154,N_1133);
or U2978 (N_2978,N_1276,N_1656);
nand U2979 (N_2979,N_1653,N_1626);
or U2980 (N_2980,N_1599,N_1536);
nor U2981 (N_2981,N_1962,N_1955);
nand U2982 (N_2982,N_1096,N_1030);
nor U2983 (N_2983,N_1008,N_1125);
nand U2984 (N_2984,N_1959,N_1980);
and U2985 (N_2985,N_1793,N_1068);
xnor U2986 (N_2986,N_1594,N_1542);
nor U2987 (N_2987,N_1843,N_1551);
nand U2988 (N_2988,N_1129,N_1549);
nand U2989 (N_2989,N_1669,N_1379);
nand U2990 (N_2990,N_1987,N_1924);
and U2991 (N_2991,N_1855,N_1837);
nor U2992 (N_2992,N_1946,N_1372);
nand U2993 (N_2993,N_1626,N_1508);
and U2994 (N_2994,N_1660,N_1778);
nor U2995 (N_2995,N_1685,N_1840);
nor U2996 (N_2996,N_1476,N_1363);
and U2997 (N_2997,N_1348,N_1610);
nor U2998 (N_2998,N_1972,N_1986);
nand U2999 (N_2999,N_1311,N_1204);
nor U3000 (N_3000,N_2086,N_2984);
xor U3001 (N_3001,N_2521,N_2531);
and U3002 (N_3002,N_2378,N_2854);
nand U3003 (N_3003,N_2816,N_2811);
or U3004 (N_3004,N_2848,N_2921);
or U3005 (N_3005,N_2817,N_2852);
and U3006 (N_3006,N_2255,N_2863);
and U3007 (N_3007,N_2159,N_2657);
and U3008 (N_3008,N_2526,N_2296);
nor U3009 (N_3009,N_2719,N_2520);
or U3010 (N_3010,N_2654,N_2669);
xor U3011 (N_3011,N_2192,N_2310);
nand U3012 (N_3012,N_2146,N_2877);
nor U3013 (N_3013,N_2263,N_2011);
and U3014 (N_3014,N_2043,N_2812);
and U3015 (N_3015,N_2470,N_2939);
nor U3016 (N_3016,N_2494,N_2433);
xnor U3017 (N_3017,N_2686,N_2254);
nor U3018 (N_3018,N_2892,N_2336);
nand U3019 (N_3019,N_2682,N_2701);
xor U3020 (N_3020,N_2393,N_2519);
or U3021 (N_3021,N_2437,N_2618);
nand U3022 (N_3022,N_2483,N_2400);
and U3023 (N_3023,N_2027,N_2387);
xnor U3024 (N_3024,N_2063,N_2133);
nand U3025 (N_3025,N_2777,N_2860);
or U3026 (N_3026,N_2136,N_2834);
xnor U3027 (N_3027,N_2611,N_2893);
nor U3028 (N_3028,N_2622,N_2584);
nor U3029 (N_3029,N_2194,N_2826);
nand U3030 (N_3030,N_2839,N_2179);
or U3031 (N_3031,N_2850,N_2218);
or U3032 (N_3032,N_2452,N_2468);
or U3033 (N_3033,N_2900,N_2183);
nor U3034 (N_3034,N_2022,N_2971);
and U3035 (N_3035,N_2069,N_2078);
nor U3036 (N_3036,N_2660,N_2357);
or U3037 (N_3037,N_2407,N_2328);
or U3038 (N_3038,N_2420,N_2666);
nand U3039 (N_3039,N_2766,N_2829);
nor U3040 (N_3040,N_2227,N_2912);
or U3041 (N_3041,N_2004,N_2072);
nor U3042 (N_3042,N_2607,N_2486);
nor U3043 (N_3043,N_2754,N_2538);
and U3044 (N_3044,N_2942,N_2205);
nor U3045 (N_3045,N_2124,N_2201);
and U3046 (N_3046,N_2469,N_2785);
and U3047 (N_3047,N_2074,N_2096);
or U3048 (N_3048,N_2640,N_2768);
xnor U3049 (N_3049,N_2722,N_2335);
and U3050 (N_3050,N_2650,N_2623);
or U3051 (N_3051,N_2954,N_2792);
and U3052 (N_3052,N_2738,N_2464);
and U3053 (N_3053,N_2139,N_2130);
nand U3054 (N_3054,N_2188,N_2976);
xnor U3055 (N_3055,N_2454,N_2555);
or U3056 (N_3056,N_2889,N_2182);
nand U3057 (N_3057,N_2964,N_2858);
nor U3058 (N_3058,N_2597,N_2292);
xor U3059 (N_3059,N_2102,N_2569);
and U3060 (N_3060,N_2117,N_2511);
xnor U3061 (N_3061,N_2311,N_2392);
xor U3062 (N_3062,N_2616,N_2228);
or U3063 (N_3063,N_2568,N_2356);
xor U3064 (N_3064,N_2421,N_2406);
and U3065 (N_3065,N_2677,N_2794);
nand U3066 (N_3066,N_2489,N_2633);
nand U3067 (N_3067,N_2054,N_2248);
nand U3068 (N_3068,N_2718,N_2985);
and U3069 (N_3069,N_2068,N_2523);
nor U3070 (N_3070,N_2095,N_2636);
nor U3071 (N_3071,N_2176,N_2859);
and U3072 (N_3072,N_2385,N_2541);
nand U3073 (N_3073,N_2294,N_2259);
xor U3074 (N_3074,N_2527,N_2331);
nand U3075 (N_3075,N_2771,N_2325);
and U3076 (N_3076,N_2951,N_2522);
nand U3077 (N_3077,N_2560,N_2989);
or U3078 (N_3078,N_2021,N_2838);
nand U3079 (N_3079,N_2953,N_2429);
and U3080 (N_3080,N_2288,N_2362);
nand U3081 (N_3081,N_2591,N_2846);
nor U3082 (N_3082,N_2815,N_2390);
nand U3083 (N_3083,N_2023,N_2656);
nand U3084 (N_3084,N_2342,N_2033);
and U3085 (N_3085,N_2167,N_2424);
nand U3086 (N_3086,N_2317,N_2564);
nand U3087 (N_3087,N_2714,N_2732);
or U3088 (N_3088,N_2014,N_2036);
and U3089 (N_3089,N_2477,N_2217);
nor U3090 (N_3090,N_2155,N_2386);
nand U3091 (N_3091,N_2134,N_2059);
nor U3092 (N_3092,N_2352,N_2673);
nand U3093 (N_3093,N_2642,N_2837);
or U3094 (N_3094,N_2810,N_2933);
nor U3095 (N_3095,N_2937,N_2580);
nand U3096 (N_3096,N_2824,N_2741);
nor U3097 (N_3097,N_2710,N_2243);
and U3098 (N_3098,N_2371,N_2046);
nand U3099 (N_3099,N_2676,N_2170);
and U3100 (N_3100,N_2482,N_2554);
nand U3101 (N_3101,N_2299,N_2641);
nand U3102 (N_3102,N_2195,N_2475);
or U3103 (N_3103,N_2467,N_2045);
or U3104 (N_3104,N_2037,N_2465);
nand U3105 (N_3105,N_2298,N_2143);
nand U3106 (N_3106,N_2952,N_2729);
nor U3107 (N_3107,N_2605,N_2213);
nor U3108 (N_3108,N_2587,N_2319);
nand U3109 (N_3109,N_2051,N_2236);
and U3110 (N_3110,N_2105,N_2232);
nand U3111 (N_3111,N_2290,N_2833);
nand U3112 (N_3112,N_2664,N_2637);
nor U3113 (N_3113,N_2830,N_2935);
xnor U3114 (N_3114,N_2670,N_2349);
xor U3115 (N_3115,N_2518,N_2355);
xnor U3116 (N_3116,N_2125,N_2745);
xor U3117 (N_3117,N_2481,N_2153);
xor U3118 (N_3118,N_2450,N_2551);
xor U3119 (N_3119,N_2044,N_2338);
nor U3120 (N_3120,N_2016,N_2244);
and U3121 (N_3121,N_2679,N_2277);
or U3122 (N_3122,N_2535,N_2770);
and U3123 (N_3123,N_2737,N_2160);
nand U3124 (N_3124,N_2408,N_2561);
xor U3125 (N_3125,N_2533,N_2559);
nor U3126 (N_3126,N_2997,N_2229);
xnor U3127 (N_3127,N_2844,N_2870);
xor U3128 (N_3128,N_2060,N_2867);
xnor U3129 (N_3129,N_2749,N_2760);
and U3130 (N_3130,N_2261,N_2425);
nor U3131 (N_3131,N_2113,N_2142);
nor U3132 (N_3132,N_2586,N_2085);
or U3133 (N_3133,N_2916,N_2361);
or U3134 (N_3134,N_2906,N_2499);
nand U3135 (N_3135,N_2093,N_2208);
xor U3136 (N_3136,N_2164,N_2963);
xnor U3137 (N_3137,N_2266,N_2376);
nor U3138 (N_3138,N_2757,N_2969);
and U3139 (N_3139,N_2825,N_2725);
nor U3140 (N_3140,N_2126,N_2999);
xnor U3141 (N_3141,N_2540,N_2665);
and U3142 (N_3142,N_2012,N_2430);
xnor U3143 (N_3143,N_2603,N_2238);
and U3144 (N_3144,N_2222,N_2226);
xor U3145 (N_3145,N_2695,N_2571);
or U3146 (N_3146,N_2927,N_2365);
and U3147 (N_3147,N_2956,N_2765);
and U3148 (N_3148,N_2747,N_2274);
or U3149 (N_3149,N_2783,N_2127);
or U3150 (N_3150,N_2857,N_2663);
xor U3151 (N_3151,N_2536,N_2493);
xor U3152 (N_3152,N_2211,N_2849);
nor U3153 (N_3153,N_2391,N_2284);
nor U3154 (N_3154,N_2318,N_2048);
xnor U3155 (N_3155,N_2472,N_2874);
xnor U3156 (N_3156,N_2862,N_2478);
nor U3157 (N_3157,N_2786,N_2065);
nor U3158 (N_3158,N_2831,N_2716);
nor U3159 (N_3159,N_2109,N_2853);
and U3160 (N_3160,N_2256,N_2260);
and U3161 (N_3161,N_2692,N_2721);
nor U3162 (N_3162,N_2556,N_2509);
or U3163 (N_3163,N_2806,N_2052);
or U3164 (N_3164,N_2449,N_2247);
and U3165 (N_3165,N_2131,N_2885);
or U3166 (N_3166,N_2621,N_2647);
xor U3167 (N_3167,N_2345,N_2156);
nor U3168 (N_3168,N_2643,N_2461);
nand U3169 (N_3169,N_2517,N_2735);
xor U3170 (N_3170,N_2351,N_2726);
xnor U3171 (N_3171,N_2138,N_2098);
and U3172 (N_3172,N_2545,N_2928);
xnor U3173 (N_3173,N_2306,N_2106);
nand U3174 (N_3174,N_2053,N_2110);
nor U3175 (N_3175,N_2638,N_2791);
or U3176 (N_3176,N_2058,N_2491);
and U3177 (N_3177,N_2653,N_2974);
and U3178 (N_3178,N_2377,N_2122);
nor U3179 (N_3179,N_2304,N_2764);
nor U3180 (N_3180,N_2769,N_2381);
or U3181 (N_3181,N_2932,N_2734);
xor U3182 (N_3182,N_2414,N_2685);
or U3183 (N_3183,N_2428,N_2364);
xnor U3184 (N_3184,N_2197,N_2804);
nor U3185 (N_3185,N_2905,N_2574);
and U3186 (N_3186,N_2013,N_2209);
xor U3187 (N_3187,N_2823,N_2782);
nor U3188 (N_3188,N_2150,N_2432);
nor U3189 (N_3189,N_2819,N_2998);
or U3190 (N_3190,N_2083,N_2447);
or U3191 (N_3191,N_2443,N_2329);
and U3192 (N_3192,N_2359,N_2525);
or U3193 (N_3193,N_2832,N_2925);
or U3194 (N_3194,N_2909,N_2042);
nand U3195 (N_3195,N_2978,N_2700);
xor U3196 (N_3196,N_2258,N_2994);
nor U3197 (N_3197,N_2774,N_2417);
nand U3198 (N_3198,N_2005,N_2191);
xnor U3199 (N_3199,N_2582,N_2444);
xor U3200 (N_3200,N_2972,N_2748);
nor U3201 (N_3201,N_2610,N_2820);
nand U3202 (N_3202,N_2115,N_2594);
xnor U3203 (N_3203,N_2202,N_2471);
xnor U3204 (N_3204,N_2092,N_2703);
or U3205 (N_3205,N_2308,N_2613);
nand U3206 (N_3206,N_2856,N_2091);
and U3207 (N_3207,N_2029,N_2672);
xnor U3208 (N_3208,N_2436,N_2715);
xnor U3209 (N_3209,N_2300,N_2918);
and U3210 (N_3210,N_2632,N_2712);
nand U3211 (N_3211,N_2347,N_2171);
or U3212 (N_3212,N_2917,N_2612);
xnor U3213 (N_3213,N_2809,N_2223);
and U3214 (N_3214,N_2773,N_2941);
nand U3215 (N_3215,N_2872,N_2101);
xor U3216 (N_3216,N_2512,N_2090);
nand U3217 (N_3217,N_2088,N_2990);
or U3218 (N_3218,N_2314,N_2901);
nor U3219 (N_3219,N_2462,N_2007);
nand U3220 (N_3220,N_2082,N_2445);
or U3221 (N_3221,N_2221,N_2619);
nor U3222 (N_3222,N_2711,N_2674);
and U3223 (N_3223,N_2675,N_2966);
nand U3224 (N_3224,N_2010,N_2544);
and U3225 (N_3225,N_2434,N_2693);
nand U3226 (N_3226,N_2358,N_2890);
or U3227 (N_3227,N_2111,N_2546);
or U3228 (N_3228,N_2458,N_2476);
nand U3229 (N_3229,N_2084,N_2780);
and U3230 (N_3230,N_2842,N_2626);
and U3231 (N_3231,N_2845,N_2168);
nand U3232 (N_3232,N_2077,N_2380);
and U3233 (N_3233,N_2724,N_2129);
nor U3234 (N_3234,N_2455,N_2373);
and U3235 (N_3235,N_2898,N_2363);
or U3236 (N_3236,N_2869,N_2140);
nor U3237 (N_3237,N_2062,N_2354);
nor U3238 (N_3238,N_2879,N_2422);
nand U3239 (N_3239,N_2828,N_2814);
nor U3240 (N_3240,N_2000,N_2270);
xnor U3241 (N_3241,N_2755,N_2061);
xor U3242 (N_3242,N_2799,N_2220);
and U3243 (N_3243,N_2320,N_2793);
nor U3244 (N_3244,N_2507,N_2655);
nand U3245 (N_3245,N_2257,N_2868);
or U3246 (N_3246,N_2936,N_2697);
or U3247 (N_3247,N_2698,N_2880);
xnor U3248 (N_3248,N_2303,N_2914);
or U3249 (N_3249,N_2350,N_2104);
nand U3250 (N_3250,N_2949,N_2330);
and U3251 (N_3251,N_2911,N_2463);
or U3252 (N_3252,N_2137,N_2239);
nand U3253 (N_3253,N_2702,N_2961);
xnor U3254 (N_3254,N_2441,N_2075);
nand U3255 (N_3255,N_2505,N_2267);
nand U3256 (N_3256,N_2798,N_2460);
nor U3257 (N_3257,N_2415,N_2973);
or U3258 (N_3258,N_2279,N_2614);
nand U3259 (N_3259,N_2479,N_2323);
xor U3260 (N_3260,N_2409,N_2808);
and U3261 (N_3261,N_2038,N_2861);
and U3262 (N_3262,N_2305,N_2631);
nor U3263 (N_3263,N_2278,N_2658);
or U3264 (N_3264,N_2864,N_2931);
xnor U3265 (N_3265,N_2602,N_2787);
nand U3266 (N_3266,N_2181,N_2235);
and U3267 (N_3267,N_2435,N_2592);
or U3268 (N_3268,N_2600,N_2070);
xor U3269 (N_3269,N_2596,N_2206);
xor U3270 (N_3270,N_2652,N_2339);
xor U3271 (N_3271,N_2426,N_2573);
nand U3272 (N_3272,N_2583,N_2903);
xnor U3273 (N_3273,N_2529,N_2418);
xnor U3274 (N_3274,N_2416,N_2813);
and U3275 (N_3275,N_2283,N_2207);
or U3276 (N_3276,N_2297,N_2291);
nand U3277 (N_3277,N_2788,N_2410);
nor U3278 (N_3278,N_2524,N_2601);
and U3279 (N_3279,N_2411,N_2929);
and U3280 (N_3280,N_2480,N_2558);
xor U3281 (N_3281,N_2246,N_2694);
or U3282 (N_3282,N_2488,N_2172);
or U3283 (N_3283,N_2097,N_2431);
nand U3284 (N_3284,N_2412,N_2187);
nor U3285 (N_3285,N_2135,N_2174);
nand U3286 (N_3286,N_2562,N_2485);
xnor U3287 (N_3287,N_2980,N_2696);
xor U3288 (N_3288,N_2539,N_2372);
and U3289 (N_3289,N_2624,N_2326);
or U3290 (N_3290,N_2039,N_2606);
or U3291 (N_3291,N_2103,N_2275);
nand U3292 (N_3292,N_2720,N_2731);
nand U3293 (N_3293,N_2822,N_2967);
xor U3294 (N_3294,N_2908,N_2934);
or U3295 (N_3295,N_2293,N_2996);
or U3296 (N_3296,N_2646,N_2727);
or U3297 (N_3297,N_2215,N_2026);
and U3298 (N_3298,N_2289,N_2369);
or U3299 (N_3299,N_2958,N_2549);
nor U3300 (N_3300,N_2145,N_2413);
xnor U3301 (N_3301,N_2552,N_2923);
and U3302 (N_3302,N_2821,N_2500);
or U3303 (N_3303,N_2730,N_2767);
xnor U3304 (N_3304,N_2661,N_2891);
or U3305 (N_3305,N_2119,N_2706);
or U3306 (N_3306,N_2570,N_2805);
nor U3307 (N_3307,N_2132,N_2047);
and U3308 (N_3308,N_2177,N_2881);
or U3309 (N_3309,N_2678,N_2855);
nand U3310 (N_3310,N_2800,N_2883);
nor U3311 (N_3311,N_2576,N_2286);
xnor U3312 (N_3312,N_2018,N_2273);
nand U3313 (N_3313,N_2991,N_2717);
xnor U3314 (N_3314,N_2884,N_2548);
xnor U3315 (N_3315,N_2144,N_2920);
xor U3316 (N_3316,N_2055,N_2272);
nor U3317 (N_3317,N_2598,N_2282);
nand U3318 (N_3318,N_2644,N_2002);
nor U3319 (N_3319,N_2687,N_2309);
nand U3320 (N_3320,N_2240,N_2108);
xnor U3321 (N_3321,N_2690,N_2397);
or U3322 (N_3322,N_2689,N_2375);
nor U3323 (N_3323,N_2629,N_2200);
and U3324 (N_3324,N_2180,N_2490);
nand U3325 (N_3325,N_2402,N_2079);
xor U3326 (N_3326,N_2684,N_2620);
or U3327 (N_3327,N_2389,N_2346);
nand U3328 (N_3328,N_2818,N_2913);
nand U3329 (N_3329,N_2370,N_2563);
nor U3330 (N_3330,N_2019,N_2383);
xor U3331 (N_3331,N_2216,N_2340);
or U3332 (N_3332,N_2959,N_2659);
nand U3333 (N_3333,N_2020,N_2333);
or U3334 (N_3334,N_2532,N_2957);
nand U3335 (N_3335,N_2344,N_2926);
or U3336 (N_3336,N_2705,N_2199);
and U3337 (N_3337,N_2271,N_2713);
nand U3338 (N_3338,N_2341,N_2944);
xnor U3339 (N_3339,N_2185,N_2161);
xor U3340 (N_3340,N_2699,N_2154);
nor U3341 (N_3341,N_2789,N_2743);
xnor U3342 (N_3342,N_2634,N_2025);
nor U3343 (N_3343,N_2752,N_2628);
and U3344 (N_3344,N_2190,N_2955);
nor U3345 (N_3345,N_2827,N_2847);
or U3346 (N_3346,N_2151,N_2457);
and U3347 (N_3347,N_2865,N_2803);
xnor U3348 (N_3348,N_2099,N_2948);
or U3349 (N_3349,N_2453,N_2353);
nor U3350 (N_3350,N_2986,N_2017);
xnor U3351 (N_3351,N_2534,N_2506);
or U3352 (N_3352,N_2401,N_2938);
nand U3353 (N_3353,N_2593,N_2028);
nor U3354 (N_3354,N_2924,N_2495);
or U3355 (N_3355,N_2427,N_2440);
nand U3356 (N_3356,N_2112,N_2742);
or U3357 (N_3357,N_2797,N_2671);
nor U3358 (N_3358,N_2439,N_2899);
and U3359 (N_3359,N_2873,N_2423);
and U3360 (N_3360,N_2578,N_2588);
nor U3361 (N_3361,N_2975,N_2565);
xnor U3362 (N_3362,N_2313,N_2076);
xor U3363 (N_3363,N_2683,N_2250);
nand U3364 (N_3364,N_2759,N_2904);
xor U3365 (N_3365,N_2639,N_2231);
nand U3366 (N_3366,N_2395,N_2530);
xor U3367 (N_3367,N_2128,N_2031);
nand U3368 (N_3368,N_2466,N_2049);
nor U3369 (N_3369,N_2006,N_2508);
nor U3370 (N_3370,N_2977,N_2550);
nor U3371 (N_3371,N_2368,N_2513);
xnor U3372 (N_3372,N_2995,N_2241);
or U3373 (N_3373,N_2709,N_2089);
nand U3374 (N_3374,N_2148,N_2035);
nand U3375 (N_3375,N_2744,N_2772);
xnor U3376 (N_3376,N_2739,N_2504);
nand U3377 (N_3377,N_2635,N_2212);
xnor U3378 (N_3378,N_2123,N_2790);
nand U3379 (N_3379,N_2776,N_2152);
nand U3380 (N_3380,N_2875,N_2147);
xnor U3381 (N_3381,N_2166,N_2141);
xor U3382 (N_3382,N_2316,N_2866);
xor U3383 (N_3383,N_2723,N_2178);
nor U3384 (N_3384,N_2287,N_2301);
or U3385 (N_3385,N_2446,N_2557);
or U3386 (N_3386,N_2982,N_2740);
nand U3387 (N_3387,N_2149,N_2579);
or U3388 (N_3388,N_2992,N_2252);
nand U3389 (N_3389,N_2514,N_2915);
nor U3390 (N_3390,N_2708,N_2327);
and U3391 (N_3391,N_2394,N_2919);
nor U3392 (N_3392,N_2572,N_2662);
nand U3393 (N_3393,N_2897,N_2253);
and U3394 (N_3394,N_2750,N_2886);
or U3395 (N_3395,N_2030,N_2081);
or U3396 (N_3396,N_2210,N_2057);
nand U3397 (N_3397,N_2173,N_2071);
or U3398 (N_3398,N_2382,N_2567);
nor U3399 (N_3399,N_2746,N_2040);
or U3400 (N_3400,N_2302,N_2736);
nor U3401 (N_3401,N_2566,N_2324);
nand U3402 (N_3402,N_2264,N_2484);
and U3403 (N_3403,N_2487,N_2474);
xor U3404 (N_3404,N_2196,N_2778);
xor U3405 (N_3405,N_2775,N_2801);
xor U3406 (N_3406,N_2322,N_2163);
or U3407 (N_3407,N_2668,N_2896);
xnor U3408 (N_3408,N_2003,N_2249);
nor U3409 (N_3409,N_2728,N_2366);
nand U3410 (N_3410,N_2276,N_2073);
and U3411 (N_3411,N_2094,N_2280);
xnor U3412 (N_3412,N_2459,N_2064);
nand U3413 (N_3413,N_2761,N_2503);
and U3414 (N_3414,N_2186,N_2492);
nor U3415 (N_3415,N_2399,N_2510);
or U3416 (N_3416,N_2707,N_2608);
xnor U3417 (N_3417,N_2100,N_2515);
or U3418 (N_3418,N_2802,N_2553);
or U3419 (N_3419,N_2496,N_2876);
or U3420 (N_3420,N_2080,N_2945);
nor U3421 (N_3421,N_2056,N_2981);
xor U3422 (N_3422,N_2871,N_2807);
nor U3423 (N_3423,N_2041,N_2251);
xor U3424 (N_3424,N_2922,N_2645);
and U3425 (N_3425,N_2691,N_2547);
xnor U3426 (N_3426,N_2763,N_2988);
nand U3427 (N_3427,N_2681,N_2947);
xnor U3428 (N_3428,N_2169,N_2950);
nand U3429 (N_3429,N_2343,N_2979);
and U3430 (N_3430,N_2204,N_2498);
nor U3431 (N_3431,N_2184,N_2379);
nand U3432 (N_3432,N_2295,N_2087);
or U3433 (N_3433,N_2067,N_2840);
xor U3434 (N_3434,N_2285,N_2970);
nand U3435 (N_3435,N_2116,N_2599);
nor U3436 (N_3436,N_2015,N_2265);
and U3437 (N_3437,N_2965,N_2404);
or U3438 (N_3438,N_2269,N_2009);
nor U3439 (N_3439,N_2193,N_2882);
or U3440 (N_3440,N_2940,N_2625);
nand U3441 (N_3441,N_2337,N_2451);
and U3442 (N_3442,N_2367,N_2751);
nand U3443 (N_3443,N_2024,N_2907);
or U3444 (N_3444,N_2784,N_2242);
or U3445 (N_3445,N_2581,N_2118);
or U3446 (N_3446,N_2595,N_2237);
nor U3447 (N_3447,N_2157,N_2501);
nor U3448 (N_3448,N_2543,N_2312);
and U3449 (N_3449,N_2442,N_2983);
xnor U3450 (N_3450,N_2050,N_2419);
or U3451 (N_3451,N_2262,N_2680);
nor U3452 (N_3452,N_2497,N_2609);
nand U3453 (N_3453,N_2396,N_2120);
nor U3454 (N_3454,N_2398,N_2943);
nand U3455 (N_3455,N_2667,N_2034);
and U3456 (N_3456,N_2307,N_2245);
xnor U3457 (N_3457,N_2651,N_2374);
xnor U3458 (N_3458,N_2756,N_2894);
xnor U3459 (N_3459,N_2203,N_2528);
and U3460 (N_3460,N_2281,N_2836);
nand U3461 (N_3461,N_2032,N_2649);
nor U3462 (N_3462,N_2960,N_2175);
nor U3463 (N_3463,N_2888,N_2604);
xor U3464 (N_3464,N_2930,N_2438);
nand U3465 (N_3465,N_2615,N_2733);
and U3466 (N_3466,N_2781,N_2502);
nor U3467 (N_3467,N_2225,N_2585);
and U3468 (N_3468,N_2158,N_2162);
and U3469 (N_3469,N_2946,N_2851);
nand U3470 (N_3470,N_2334,N_2910);
or U3471 (N_3471,N_2688,N_2779);
and U3472 (N_3472,N_2796,N_2704);
nand U3473 (N_3473,N_2001,N_2987);
or U3474 (N_3474,N_2230,N_2887);
xor U3475 (N_3475,N_2473,N_2405);
or U3476 (N_3476,N_2233,N_2758);
nor U3477 (N_3477,N_2843,N_2360);
xnor U3478 (N_3478,N_2968,N_2268);
or U3479 (N_3479,N_2648,N_2577);
nand U3480 (N_3480,N_2448,N_2575);
and U3481 (N_3481,N_2388,N_2214);
xor U3482 (N_3482,N_2962,N_2008);
nor U3483 (N_3483,N_2993,N_2542);
xor U3484 (N_3484,N_2321,N_2198);
nor U3485 (N_3485,N_2234,N_2121);
xor U3486 (N_3486,N_2630,N_2753);
or U3487 (N_3487,N_2795,N_2617);
nor U3488 (N_3488,N_2114,N_2066);
and U3489 (N_3489,N_2403,N_2627);
nor U3490 (N_3490,N_2841,N_2878);
nor U3491 (N_3491,N_2384,N_2590);
or U3492 (N_3492,N_2219,N_2107);
or U3493 (N_3493,N_2835,N_2589);
nand U3494 (N_3494,N_2224,N_2189);
nand U3495 (N_3495,N_2762,N_2456);
or U3496 (N_3496,N_2537,N_2315);
nor U3497 (N_3497,N_2902,N_2332);
nor U3498 (N_3498,N_2165,N_2895);
or U3499 (N_3499,N_2348,N_2516);
or U3500 (N_3500,N_2570,N_2333);
or U3501 (N_3501,N_2688,N_2129);
or U3502 (N_3502,N_2292,N_2383);
xor U3503 (N_3503,N_2774,N_2371);
nand U3504 (N_3504,N_2285,N_2535);
xnor U3505 (N_3505,N_2560,N_2718);
or U3506 (N_3506,N_2704,N_2586);
xor U3507 (N_3507,N_2519,N_2011);
nor U3508 (N_3508,N_2018,N_2410);
nand U3509 (N_3509,N_2932,N_2137);
or U3510 (N_3510,N_2087,N_2954);
xnor U3511 (N_3511,N_2066,N_2459);
nor U3512 (N_3512,N_2913,N_2836);
and U3513 (N_3513,N_2105,N_2194);
nor U3514 (N_3514,N_2278,N_2598);
xnor U3515 (N_3515,N_2272,N_2498);
nor U3516 (N_3516,N_2088,N_2499);
nor U3517 (N_3517,N_2387,N_2301);
and U3518 (N_3518,N_2706,N_2717);
nand U3519 (N_3519,N_2724,N_2214);
or U3520 (N_3520,N_2313,N_2406);
xor U3521 (N_3521,N_2570,N_2411);
nand U3522 (N_3522,N_2718,N_2808);
or U3523 (N_3523,N_2686,N_2063);
nand U3524 (N_3524,N_2818,N_2417);
and U3525 (N_3525,N_2878,N_2116);
nand U3526 (N_3526,N_2767,N_2696);
or U3527 (N_3527,N_2528,N_2259);
or U3528 (N_3528,N_2669,N_2034);
or U3529 (N_3529,N_2471,N_2195);
xor U3530 (N_3530,N_2309,N_2122);
nor U3531 (N_3531,N_2613,N_2207);
nor U3532 (N_3532,N_2599,N_2843);
nand U3533 (N_3533,N_2353,N_2051);
nand U3534 (N_3534,N_2720,N_2179);
nand U3535 (N_3535,N_2656,N_2569);
nand U3536 (N_3536,N_2316,N_2928);
xor U3537 (N_3537,N_2614,N_2841);
or U3538 (N_3538,N_2250,N_2435);
nor U3539 (N_3539,N_2903,N_2144);
and U3540 (N_3540,N_2794,N_2139);
nor U3541 (N_3541,N_2241,N_2326);
and U3542 (N_3542,N_2083,N_2783);
and U3543 (N_3543,N_2938,N_2792);
or U3544 (N_3544,N_2493,N_2679);
or U3545 (N_3545,N_2673,N_2692);
xnor U3546 (N_3546,N_2144,N_2332);
or U3547 (N_3547,N_2998,N_2402);
xnor U3548 (N_3548,N_2188,N_2917);
xnor U3549 (N_3549,N_2442,N_2823);
nand U3550 (N_3550,N_2320,N_2242);
xnor U3551 (N_3551,N_2980,N_2160);
or U3552 (N_3552,N_2765,N_2002);
and U3553 (N_3553,N_2426,N_2247);
or U3554 (N_3554,N_2587,N_2952);
and U3555 (N_3555,N_2904,N_2069);
xor U3556 (N_3556,N_2326,N_2749);
or U3557 (N_3557,N_2676,N_2273);
or U3558 (N_3558,N_2297,N_2550);
nor U3559 (N_3559,N_2959,N_2166);
xor U3560 (N_3560,N_2264,N_2110);
nor U3561 (N_3561,N_2566,N_2115);
nor U3562 (N_3562,N_2774,N_2343);
nor U3563 (N_3563,N_2794,N_2787);
nand U3564 (N_3564,N_2247,N_2138);
and U3565 (N_3565,N_2562,N_2862);
xnor U3566 (N_3566,N_2985,N_2335);
nor U3567 (N_3567,N_2133,N_2278);
and U3568 (N_3568,N_2013,N_2127);
or U3569 (N_3569,N_2368,N_2227);
or U3570 (N_3570,N_2724,N_2678);
and U3571 (N_3571,N_2866,N_2449);
and U3572 (N_3572,N_2190,N_2906);
nor U3573 (N_3573,N_2962,N_2885);
or U3574 (N_3574,N_2880,N_2198);
nand U3575 (N_3575,N_2446,N_2509);
or U3576 (N_3576,N_2564,N_2444);
and U3577 (N_3577,N_2061,N_2813);
nor U3578 (N_3578,N_2893,N_2445);
nor U3579 (N_3579,N_2857,N_2920);
xor U3580 (N_3580,N_2950,N_2888);
xnor U3581 (N_3581,N_2633,N_2325);
and U3582 (N_3582,N_2927,N_2969);
nor U3583 (N_3583,N_2577,N_2216);
and U3584 (N_3584,N_2318,N_2395);
or U3585 (N_3585,N_2227,N_2101);
xor U3586 (N_3586,N_2394,N_2319);
and U3587 (N_3587,N_2663,N_2172);
xor U3588 (N_3588,N_2187,N_2906);
nor U3589 (N_3589,N_2706,N_2689);
or U3590 (N_3590,N_2672,N_2863);
nor U3591 (N_3591,N_2857,N_2319);
and U3592 (N_3592,N_2954,N_2448);
or U3593 (N_3593,N_2204,N_2408);
and U3594 (N_3594,N_2599,N_2287);
or U3595 (N_3595,N_2156,N_2898);
nor U3596 (N_3596,N_2502,N_2325);
or U3597 (N_3597,N_2934,N_2546);
xnor U3598 (N_3598,N_2273,N_2555);
nor U3599 (N_3599,N_2836,N_2544);
nand U3600 (N_3600,N_2013,N_2036);
nor U3601 (N_3601,N_2271,N_2718);
and U3602 (N_3602,N_2364,N_2488);
nand U3603 (N_3603,N_2195,N_2890);
and U3604 (N_3604,N_2264,N_2889);
and U3605 (N_3605,N_2022,N_2415);
and U3606 (N_3606,N_2761,N_2087);
and U3607 (N_3607,N_2204,N_2291);
or U3608 (N_3608,N_2504,N_2899);
nand U3609 (N_3609,N_2541,N_2980);
xnor U3610 (N_3610,N_2810,N_2414);
or U3611 (N_3611,N_2740,N_2112);
nor U3612 (N_3612,N_2913,N_2642);
or U3613 (N_3613,N_2080,N_2790);
nor U3614 (N_3614,N_2902,N_2306);
or U3615 (N_3615,N_2572,N_2466);
and U3616 (N_3616,N_2032,N_2254);
or U3617 (N_3617,N_2817,N_2606);
or U3618 (N_3618,N_2293,N_2980);
nor U3619 (N_3619,N_2031,N_2979);
nor U3620 (N_3620,N_2895,N_2931);
nand U3621 (N_3621,N_2701,N_2099);
xor U3622 (N_3622,N_2743,N_2541);
nand U3623 (N_3623,N_2068,N_2100);
nor U3624 (N_3624,N_2975,N_2522);
or U3625 (N_3625,N_2722,N_2279);
nor U3626 (N_3626,N_2895,N_2498);
and U3627 (N_3627,N_2781,N_2350);
and U3628 (N_3628,N_2121,N_2511);
xnor U3629 (N_3629,N_2985,N_2245);
nand U3630 (N_3630,N_2831,N_2241);
nor U3631 (N_3631,N_2246,N_2253);
xnor U3632 (N_3632,N_2436,N_2052);
xor U3633 (N_3633,N_2455,N_2316);
or U3634 (N_3634,N_2322,N_2109);
nor U3635 (N_3635,N_2048,N_2651);
or U3636 (N_3636,N_2550,N_2998);
nand U3637 (N_3637,N_2325,N_2130);
nand U3638 (N_3638,N_2105,N_2786);
xor U3639 (N_3639,N_2500,N_2871);
nand U3640 (N_3640,N_2605,N_2040);
and U3641 (N_3641,N_2423,N_2554);
or U3642 (N_3642,N_2881,N_2748);
nand U3643 (N_3643,N_2176,N_2886);
nor U3644 (N_3644,N_2832,N_2937);
nand U3645 (N_3645,N_2002,N_2172);
and U3646 (N_3646,N_2070,N_2697);
and U3647 (N_3647,N_2377,N_2907);
nor U3648 (N_3648,N_2501,N_2723);
and U3649 (N_3649,N_2591,N_2481);
nand U3650 (N_3650,N_2345,N_2614);
xor U3651 (N_3651,N_2987,N_2337);
and U3652 (N_3652,N_2993,N_2637);
nor U3653 (N_3653,N_2724,N_2006);
xnor U3654 (N_3654,N_2243,N_2811);
and U3655 (N_3655,N_2590,N_2145);
nor U3656 (N_3656,N_2857,N_2435);
xor U3657 (N_3657,N_2975,N_2970);
and U3658 (N_3658,N_2438,N_2553);
nand U3659 (N_3659,N_2463,N_2551);
or U3660 (N_3660,N_2348,N_2615);
xnor U3661 (N_3661,N_2534,N_2626);
and U3662 (N_3662,N_2396,N_2343);
nand U3663 (N_3663,N_2346,N_2587);
xor U3664 (N_3664,N_2502,N_2339);
and U3665 (N_3665,N_2125,N_2084);
xor U3666 (N_3666,N_2461,N_2251);
and U3667 (N_3667,N_2541,N_2793);
nor U3668 (N_3668,N_2356,N_2480);
nand U3669 (N_3669,N_2888,N_2314);
and U3670 (N_3670,N_2579,N_2582);
nor U3671 (N_3671,N_2834,N_2296);
nor U3672 (N_3672,N_2043,N_2186);
or U3673 (N_3673,N_2146,N_2645);
xor U3674 (N_3674,N_2847,N_2695);
nor U3675 (N_3675,N_2188,N_2434);
xor U3676 (N_3676,N_2990,N_2648);
and U3677 (N_3677,N_2771,N_2001);
and U3678 (N_3678,N_2397,N_2003);
nor U3679 (N_3679,N_2587,N_2193);
nor U3680 (N_3680,N_2292,N_2481);
xor U3681 (N_3681,N_2363,N_2465);
xor U3682 (N_3682,N_2050,N_2454);
nor U3683 (N_3683,N_2671,N_2972);
or U3684 (N_3684,N_2074,N_2464);
nor U3685 (N_3685,N_2375,N_2355);
or U3686 (N_3686,N_2656,N_2310);
nor U3687 (N_3687,N_2871,N_2348);
nand U3688 (N_3688,N_2318,N_2561);
nor U3689 (N_3689,N_2880,N_2977);
and U3690 (N_3690,N_2893,N_2303);
and U3691 (N_3691,N_2269,N_2257);
or U3692 (N_3692,N_2605,N_2352);
and U3693 (N_3693,N_2173,N_2031);
or U3694 (N_3694,N_2532,N_2166);
nand U3695 (N_3695,N_2889,N_2230);
nor U3696 (N_3696,N_2724,N_2436);
or U3697 (N_3697,N_2919,N_2003);
xor U3698 (N_3698,N_2627,N_2905);
or U3699 (N_3699,N_2220,N_2065);
xnor U3700 (N_3700,N_2538,N_2218);
nand U3701 (N_3701,N_2424,N_2895);
or U3702 (N_3702,N_2892,N_2095);
nor U3703 (N_3703,N_2579,N_2305);
xor U3704 (N_3704,N_2547,N_2068);
or U3705 (N_3705,N_2614,N_2182);
nor U3706 (N_3706,N_2913,N_2821);
xor U3707 (N_3707,N_2902,N_2900);
xnor U3708 (N_3708,N_2657,N_2987);
nor U3709 (N_3709,N_2207,N_2801);
xor U3710 (N_3710,N_2577,N_2933);
nand U3711 (N_3711,N_2042,N_2540);
or U3712 (N_3712,N_2075,N_2069);
and U3713 (N_3713,N_2049,N_2492);
nor U3714 (N_3714,N_2483,N_2953);
and U3715 (N_3715,N_2422,N_2606);
xor U3716 (N_3716,N_2891,N_2599);
xnor U3717 (N_3717,N_2204,N_2424);
or U3718 (N_3718,N_2235,N_2332);
nor U3719 (N_3719,N_2553,N_2840);
and U3720 (N_3720,N_2263,N_2487);
nand U3721 (N_3721,N_2692,N_2454);
or U3722 (N_3722,N_2437,N_2691);
xor U3723 (N_3723,N_2255,N_2432);
and U3724 (N_3724,N_2177,N_2056);
and U3725 (N_3725,N_2321,N_2692);
nand U3726 (N_3726,N_2704,N_2589);
nand U3727 (N_3727,N_2755,N_2005);
and U3728 (N_3728,N_2005,N_2429);
xnor U3729 (N_3729,N_2943,N_2030);
nor U3730 (N_3730,N_2838,N_2654);
xnor U3731 (N_3731,N_2269,N_2831);
or U3732 (N_3732,N_2924,N_2151);
nor U3733 (N_3733,N_2367,N_2889);
xor U3734 (N_3734,N_2618,N_2684);
or U3735 (N_3735,N_2359,N_2878);
xnor U3736 (N_3736,N_2353,N_2890);
nor U3737 (N_3737,N_2291,N_2517);
or U3738 (N_3738,N_2039,N_2761);
and U3739 (N_3739,N_2509,N_2063);
and U3740 (N_3740,N_2616,N_2231);
nor U3741 (N_3741,N_2696,N_2324);
nand U3742 (N_3742,N_2800,N_2163);
and U3743 (N_3743,N_2635,N_2362);
nand U3744 (N_3744,N_2863,N_2468);
xnor U3745 (N_3745,N_2548,N_2843);
or U3746 (N_3746,N_2956,N_2674);
xnor U3747 (N_3747,N_2060,N_2008);
xor U3748 (N_3748,N_2352,N_2057);
nor U3749 (N_3749,N_2377,N_2666);
nand U3750 (N_3750,N_2405,N_2427);
nor U3751 (N_3751,N_2229,N_2540);
nand U3752 (N_3752,N_2103,N_2825);
nand U3753 (N_3753,N_2522,N_2857);
or U3754 (N_3754,N_2673,N_2948);
or U3755 (N_3755,N_2306,N_2394);
and U3756 (N_3756,N_2557,N_2975);
or U3757 (N_3757,N_2295,N_2718);
or U3758 (N_3758,N_2361,N_2428);
and U3759 (N_3759,N_2572,N_2115);
or U3760 (N_3760,N_2751,N_2048);
and U3761 (N_3761,N_2548,N_2547);
or U3762 (N_3762,N_2423,N_2514);
or U3763 (N_3763,N_2625,N_2279);
or U3764 (N_3764,N_2127,N_2462);
nor U3765 (N_3765,N_2106,N_2844);
nor U3766 (N_3766,N_2885,N_2843);
nand U3767 (N_3767,N_2244,N_2603);
nand U3768 (N_3768,N_2300,N_2057);
and U3769 (N_3769,N_2471,N_2870);
or U3770 (N_3770,N_2550,N_2148);
xor U3771 (N_3771,N_2738,N_2192);
nor U3772 (N_3772,N_2606,N_2758);
nor U3773 (N_3773,N_2373,N_2377);
nand U3774 (N_3774,N_2256,N_2658);
and U3775 (N_3775,N_2238,N_2954);
xor U3776 (N_3776,N_2606,N_2920);
or U3777 (N_3777,N_2859,N_2985);
xnor U3778 (N_3778,N_2046,N_2824);
xor U3779 (N_3779,N_2066,N_2279);
nor U3780 (N_3780,N_2022,N_2521);
or U3781 (N_3781,N_2988,N_2155);
nand U3782 (N_3782,N_2542,N_2691);
nor U3783 (N_3783,N_2023,N_2869);
or U3784 (N_3784,N_2971,N_2562);
nor U3785 (N_3785,N_2122,N_2635);
nand U3786 (N_3786,N_2066,N_2711);
nand U3787 (N_3787,N_2751,N_2131);
and U3788 (N_3788,N_2947,N_2566);
or U3789 (N_3789,N_2868,N_2748);
nor U3790 (N_3790,N_2721,N_2265);
and U3791 (N_3791,N_2278,N_2172);
xor U3792 (N_3792,N_2712,N_2000);
and U3793 (N_3793,N_2875,N_2801);
xnor U3794 (N_3794,N_2310,N_2542);
nand U3795 (N_3795,N_2559,N_2268);
nor U3796 (N_3796,N_2852,N_2188);
nor U3797 (N_3797,N_2988,N_2630);
xnor U3798 (N_3798,N_2151,N_2068);
and U3799 (N_3799,N_2625,N_2160);
nand U3800 (N_3800,N_2274,N_2431);
and U3801 (N_3801,N_2053,N_2411);
xor U3802 (N_3802,N_2474,N_2160);
nor U3803 (N_3803,N_2552,N_2926);
nor U3804 (N_3804,N_2854,N_2381);
or U3805 (N_3805,N_2858,N_2597);
or U3806 (N_3806,N_2007,N_2641);
and U3807 (N_3807,N_2704,N_2610);
or U3808 (N_3808,N_2681,N_2979);
xor U3809 (N_3809,N_2865,N_2730);
nand U3810 (N_3810,N_2373,N_2092);
and U3811 (N_3811,N_2858,N_2631);
nand U3812 (N_3812,N_2829,N_2068);
nor U3813 (N_3813,N_2452,N_2409);
xnor U3814 (N_3814,N_2922,N_2327);
nor U3815 (N_3815,N_2194,N_2230);
nor U3816 (N_3816,N_2605,N_2787);
nand U3817 (N_3817,N_2501,N_2641);
nor U3818 (N_3818,N_2639,N_2403);
or U3819 (N_3819,N_2175,N_2892);
nor U3820 (N_3820,N_2025,N_2074);
xor U3821 (N_3821,N_2220,N_2597);
nand U3822 (N_3822,N_2758,N_2145);
and U3823 (N_3823,N_2215,N_2473);
nor U3824 (N_3824,N_2687,N_2573);
or U3825 (N_3825,N_2174,N_2786);
xor U3826 (N_3826,N_2606,N_2822);
xor U3827 (N_3827,N_2448,N_2362);
or U3828 (N_3828,N_2167,N_2102);
or U3829 (N_3829,N_2803,N_2324);
xnor U3830 (N_3830,N_2401,N_2576);
xor U3831 (N_3831,N_2714,N_2839);
and U3832 (N_3832,N_2260,N_2521);
or U3833 (N_3833,N_2521,N_2172);
xnor U3834 (N_3834,N_2482,N_2462);
xnor U3835 (N_3835,N_2319,N_2173);
and U3836 (N_3836,N_2568,N_2229);
nand U3837 (N_3837,N_2811,N_2192);
and U3838 (N_3838,N_2979,N_2585);
nand U3839 (N_3839,N_2147,N_2749);
nand U3840 (N_3840,N_2952,N_2479);
and U3841 (N_3841,N_2574,N_2482);
nand U3842 (N_3842,N_2774,N_2837);
nor U3843 (N_3843,N_2931,N_2206);
nor U3844 (N_3844,N_2502,N_2683);
nor U3845 (N_3845,N_2346,N_2496);
or U3846 (N_3846,N_2240,N_2280);
or U3847 (N_3847,N_2133,N_2549);
or U3848 (N_3848,N_2005,N_2745);
or U3849 (N_3849,N_2820,N_2827);
xnor U3850 (N_3850,N_2731,N_2738);
nand U3851 (N_3851,N_2980,N_2953);
nand U3852 (N_3852,N_2739,N_2553);
xnor U3853 (N_3853,N_2218,N_2580);
nand U3854 (N_3854,N_2542,N_2701);
xor U3855 (N_3855,N_2274,N_2687);
nand U3856 (N_3856,N_2053,N_2073);
xor U3857 (N_3857,N_2926,N_2741);
xnor U3858 (N_3858,N_2210,N_2586);
nand U3859 (N_3859,N_2516,N_2757);
nand U3860 (N_3860,N_2112,N_2123);
nand U3861 (N_3861,N_2807,N_2077);
nor U3862 (N_3862,N_2309,N_2111);
nor U3863 (N_3863,N_2928,N_2371);
and U3864 (N_3864,N_2749,N_2815);
and U3865 (N_3865,N_2867,N_2027);
xor U3866 (N_3866,N_2040,N_2345);
or U3867 (N_3867,N_2283,N_2584);
or U3868 (N_3868,N_2078,N_2879);
xnor U3869 (N_3869,N_2304,N_2526);
or U3870 (N_3870,N_2240,N_2818);
nand U3871 (N_3871,N_2949,N_2259);
or U3872 (N_3872,N_2015,N_2592);
nand U3873 (N_3873,N_2930,N_2673);
or U3874 (N_3874,N_2212,N_2587);
or U3875 (N_3875,N_2916,N_2510);
nand U3876 (N_3876,N_2373,N_2368);
and U3877 (N_3877,N_2433,N_2306);
and U3878 (N_3878,N_2854,N_2244);
and U3879 (N_3879,N_2762,N_2875);
and U3880 (N_3880,N_2099,N_2282);
nor U3881 (N_3881,N_2777,N_2154);
and U3882 (N_3882,N_2164,N_2681);
nor U3883 (N_3883,N_2578,N_2048);
nand U3884 (N_3884,N_2239,N_2045);
nor U3885 (N_3885,N_2214,N_2323);
xor U3886 (N_3886,N_2388,N_2632);
nand U3887 (N_3887,N_2373,N_2856);
or U3888 (N_3888,N_2406,N_2213);
and U3889 (N_3889,N_2132,N_2075);
and U3890 (N_3890,N_2128,N_2866);
nor U3891 (N_3891,N_2979,N_2678);
and U3892 (N_3892,N_2049,N_2005);
nand U3893 (N_3893,N_2396,N_2528);
nand U3894 (N_3894,N_2636,N_2103);
or U3895 (N_3895,N_2399,N_2358);
nor U3896 (N_3896,N_2842,N_2390);
and U3897 (N_3897,N_2459,N_2892);
nand U3898 (N_3898,N_2786,N_2570);
and U3899 (N_3899,N_2168,N_2468);
and U3900 (N_3900,N_2445,N_2667);
or U3901 (N_3901,N_2488,N_2289);
or U3902 (N_3902,N_2590,N_2088);
nor U3903 (N_3903,N_2859,N_2962);
nand U3904 (N_3904,N_2105,N_2561);
nor U3905 (N_3905,N_2556,N_2596);
nor U3906 (N_3906,N_2323,N_2777);
nand U3907 (N_3907,N_2177,N_2055);
nand U3908 (N_3908,N_2100,N_2775);
xor U3909 (N_3909,N_2864,N_2724);
or U3910 (N_3910,N_2396,N_2696);
and U3911 (N_3911,N_2098,N_2308);
or U3912 (N_3912,N_2277,N_2203);
nor U3913 (N_3913,N_2870,N_2759);
and U3914 (N_3914,N_2863,N_2557);
nor U3915 (N_3915,N_2882,N_2498);
and U3916 (N_3916,N_2194,N_2709);
and U3917 (N_3917,N_2034,N_2795);
or U3918 (N_3918,N_2319,N_2588);
and U3919 (N_3919,N_2996,N_2314);
nor U3920 (N_3920,N_2494,N_2403);
and U3921 (N_3921,N_2210,N_2137);
xnor U3922 (N_3922,N_2471,N_2679);
nor U3923 (N_3923,N_2865,N_2441);
nor U3924 (N_3924,N_2266,N_2830);
and U3925 (N_3925,N_2507,N_2028);
nand U3926 (N_3926,N_2063,N_2953);
xor U3927 (N_3927,N_2593,N_2022);
nand U3928 (N_3928,N_2678,N_2957);
or U3929 (N_3929,N_2639,N_2994);
nand U3930 (N_3930,N_2117,N_2423);
nor U3931 (N_3931,N_2669,N_2990);
nor U3932 (N_3932,N_2387,N_2351);
and U3933 (N_3933,N_2684,N_2694);
and U3934 (N_3934,N_2215,N_2993);
or U3935 (N_3935,N_2596,N_2020);
nor U3936 (N_3936,N_2165,N_2913);
or U3937 (N_3937,N_2778,N_2018);
or U3938 (N_3938,N_2618,N_2354);
nor U3939 (N_3939,N_2493,N_2283);
nor U3940 (N_3940,N_2182,N_2465);
nand U3941 (N_3941,N_2185,N_2075);
xor U3942 (N_3942,N_2811,N_2557);
nand U3943 (N_3943,N_2952,N_2228);
or U3944 (N_3944,N_2895,N_2203);
nor U3945 (N_3945,N_2543,N_2217);
or U3946 (N_3946,N_2075,N_2979);
and U3947 (N_3947,N_2762,N_2041);
and U3948 (N_3948,N_2505,N_2891);
and U3949 (N_3949,N_2666,N_2290);
and U3950 (N_3950,N_2880,N_2611);
nor U3951 (N_3951,N_2152,N_2294);
nor U3952 (N_3952,N_2860,N_2565);
xnor U3953 (N_3953,N_2942,N_2752);
xnor U3954 (N_3954,N_2079,N_2375);
nand U3955 (N_3955,N_2819,N_2750);
nor U3956 (N_3956,N_2863,N_2575);
nand U3957 (N_3957,N_2618,N_2536);
or U3958 (N_3958,N_2106,N_2489);
nor U3959 (N_3959,N_2829,N_2777);
or U3960 (N_3960,N_2961,N_2901);
nand U3961 (N_3961,N_2095,N_2666);
xnor U3962 (N_3962,N_2968,N_2811);
and U3963 (N_3963,N_2762,N_2218);
nand U3964 (N_3964,N_2402,N_2690);
and U3965 (N_3965,N_2614,N_2851);
xnor U3966 (N_3966,N_2891,N_2148);
nand U3967 (N_3967,N_2682,N_2228);
nor U3968 (N_3968,N_2366,N_2013);
xnor U3969 (N_3969,N_2312,N_2912);
and U3970 (N_3970,N_2957,N_2766);
nor U3971 (N_3971,N_2204,N_2713);
and U3972 (N_3972,N_2669,N_2631);
nor U3973 (N_3973,N_2234,N_2404);
or U3974 (N_3974,N_2370,N_2598);
and U3975 (N_3975,N_2364,N_2325);
nand U3976 (N_3976,N_2038,N_2734);
nand U3977 (N_3977,N_2044,N_2991);
nand U3978 (N_3978,N_2591,N_2862);
and U3979 (N_3979,N_2355,N_2099);
and U3980 (N_3980,N_2956,N_2297);
or U3981 (N_3981,N_2856,N_2039);
nand U3982 (N_3982,N_2758,N_2735);
nand U3983 (N_3983,N_2140,N_2703);
xnor U3984 (N_3984,N_2934,N_2489);
nor U3985 (N_3985,N_2801,N_2415);
xnor U3986 (N_3986,N_2700,N_2716);
nor U3987 (N_3987,N_2967,N_2206);
nor U3988 (N_3988,N_2823,N_2259);
nor U3989 (N_3989,N_2531,N_2177);
nand U3990 (N_3990,N_2345,N_2204);
xor U3991 (N_3991,N_2760,N_2071);
or U3992 (N_3992,N_2513,N_2710);
xor U3993 (N_3993,N_2237,N_2272);
nor U3994 (N_3994,N_2162,N_2175);
xor U3995 (N_3995,N_2551,N_2194);
nand U3996 (N_3996,N_2311,N_2879);
or U3997 (N_3997,N_2141,N_2847);
xor U3998 (N_3998,N_2842,N_2254);
xor U3999 (N_3999,N_2918,N_2343);
and U4000 (N_4000,N_3380,N_3865);
xor U4001 (N_4001,N_3496,N_3144);
nor U4002 (N_4002,N_3797,N_3356);
nand U4003 (N_4003,N_3152,N_3094);
nand U4004 (N_4004,N_3187,N_3163);
xor U4005 (N_4005,N_3641,N_3150);
or U4006 (N_4006,N_3710,N_3278);
and U4007 (N_4007,N_3201,N_3204);
nor U4008 (N_4008,N_3822,N_3998);
xor U4009 (N_4009,N_3104,N_3951);
xnor U4010 (N_4010,N_3596,N_3444);
or U4011 (N_4011,N_3165,N_3989);
xor U4012 (N_4012,N_3394,N_3243);
or U4013 (N_4013,N_3302,N_3699);
xnor U4014 (N_4014,N_3910,N_3116);
xnor U4015 (N_4015,N_3944,N_3727);
nor U4016 (N_4016,N_3584,N_3238);
xor U4017 (N_4017,N_3816,N_3233);
and U4018 (N_4018,N_3098,N_3218);
xor U4019 (N_4019,N_3782,N_3658);
xor U4020 (N_4020,N_3520,N_3425);
nand U4021 (N_4021,N_3527,N_3567);
or U4022 (N_4022,N_3849,N_3839);
nand U4023 (N_4023,N_3478,N_3331);
nor U4024 (N_4024,N_3723,N_3420);
nor U4025 (N_4025,N_3220,N_3739);
nand U4026 (N_4026,N_3623,N_3733);
xnor U4027 (N_4027,N_3117,N_3524);
or U4028 (N_4028,N_3054,N_3052);
nand U4029 (N_4029,N_3621,N_3476);
xnor U4030 (N_4030,N_3216,N_3731);
and U4031 (N_4031,N_3192,N_3337);
and U4032 (N_4032,N_3265,N_3109);
nand U4033 (N_4033,N_3426,N_3683);
nand U4034 (N_4034,N_3872,N_3259);
or U4035 (N_4035,N_3032,N_3452);
xnor U4036 (N_4036,N_3945,N_3361);
xor U4037 (N_4037,N_3007,N_3513);
and U4038 (N_4038,N_3210,N_3574);
nor U4039 (N_4039,N_3502,N_3501);
nand U4040 (N_4040,N_3770,N_3895);
or U4041 (N_4041,N_3294,N_3033);
and U4042 (N_4042,N_3393,N_3266);
nand U4043 (N_4043,N_3055,N_3140);
nor U4044 (N_4044,N_3362,N_3642);
xnor U4045 (N_4045,N_3647,N_3395);
nand U4046 (N_4046,N_3978,N_3948);
or U4047 (N_4047,N_3279,N_3020);
nand U4048 (N_4048,N_3328,N_3981);
and U4049 (N_4049,N_3592,N_3211);
and U4050 (N_4050,N_3219,N_3962);
nor U4051 (N_4051,N_3015,N_3301);
and U4052 (N_4052,N_3234,N_3409);
xor U4053 (N_4053,N_3445,N_3692);
nand U4054 (N_4054,N_3644,N_3453);
or U4055 (N_4055,N_3695,N_3235);
nor U4056 (N_4056,N_3806,N_3793);
nand U4057 (N_4057,N_3075,N_3977);
xnor U4058 (N_4058,N_3631,N_3406);
nand U4059 (N_4059,N_3374,N_3249);
or U4060 (N_4060,N_3350,N_3329);
or U4061 (N_4061,N_3252,N_3807);
and U4062 (N_4062,N_3611,N_3047);
and U4063 (N_4063,N_3506,N_3222);
xor U4064 (N_4064,N_3833,N_3427);
nand U4065 (N_4065,N_3118,N_3011);
nor U4066 (N_4066,N_3464,N_3071);
xnor U4067 (N_4067,N_3154,N_3775);
nor U4068 (N_4068,N_3515,N_3121);
and U4069 (N_4069,N_3964,N_3758);
and U4070 (N_4070,N_3143,N_3465);
or U4071 (N_4071,N_3435,N_3493);
xor U4072 (N_4072,N_3297,N_3049);
xnor U4073 (N_4073,N_3028,N_3325);
or U4074 (N_4074,N_3935,N_3480);
and U4075 (N_4075,N_3588,N_3084);
or U4076 (N_4076,N_3076,N_3538);
xnor U4077 (N_4077,N_3965,N_3198);
or U4078 (N_4078,N_3669,N_3382);
nand U4079 (N_4079,N_3751,N_3561);
or U4080 (N_4080,N_3682,N_3304);
or U4081 (N_4081,N_3954,N_3191);
xnor U4082 (N_4082,N_3283,N_3193);
xor U4083 (N_4083,N_3221,N_3859);
and U4084 (N_4084,N_3858,N_3158);
xor U4085 (N_4085,N_3196,N_3292);
nand U4086 (N_4086,N_3537,N_3558);
and U4087 (N_4087,N_3431,N_3311);
xor U4088 (N_4088,N_3971,N_3583);
or U4089 (N_4089,N_3825,N_3424);
nor U4090 (N_4090,N_3940,N_3194);
nor U4091 (N_4091,N_3632,N_3707);
nor U4092 (N_4092,N_3990,N_3375);
or U4093 (N_4093,N_3885,N_3309);
and U4094 (N_4094,N_3421,N_3817);
or U4095 (N_4095,N_3289,N_3556);
or U4096 (N_4096,N_3156,N_3418);
and U4097 (N_4097,N_3050,N_3587);
xor U4098 (N_4098,N_3860,N_3185);
or U4099 (N_4099,N_3326,N_3615);
or U4100 (N_4100,N_3730,N_3113);
or U4101 (N_4101,N_3153,N_3850);
or U4102 (N_4102,N_3923,N_3368);
nor U4103 (N_4103,N_3653,N_3072);
xnor U4104 (N_4104,N_3892,N_3392);
nand U4105 (N_4105,N_3914,N_3549);
nor U4106 (N_4106,N_3305,N_3687);
xnor U4107 (N_4107,N_3284,N_3794);
nand U4108 (N_4108,N_3928,N_3874);
nand U4109 (N_4109,N_3995,N_3876);
nand U4110 (N_4110,N_3798,N_3224);
xnor U4111 (N_4111,N_3771,N_3503);
xnor U4112 (N_4112,N_3791,N_3160);
or U4113 (N_4113,N_3159,N_3170);
xor U4114 (N_4114,N_3411,N_3510);
or U4115 (N_4115,N_3371,N_3044);
or U4116 (N_4116,N_3280,N_3061);
nor U4117 (N_4117,N_3299,N_3164);
or U4118 (N_4118,N_3236,N_3462);
nor U4119 (N_4119,N_3842,N_3030);
nor U4120 (N_4120,N_3397,N_3461);
nand U4121 (N_4121,N_3447,N_3122);
nor U4122 (N_4122,N_3343,N_3713);
or U4123 (N_4123,N_3572,N_3369);
and U4124 (N_4124,N_3268,N_3786);
and U4125 (N_4125,N_3638,N_3700);
or U4126 (N_4126,N_3626,N_3327);
or U4127 (N_4127,N_3991,N_3207);
xnor U4128 (N_4128,N_3927,N_3353);
nand U4129 (N_4129,N_3423,N_3985);
or U4130 (N_4130,N_3486,N_3704);
nor U4131 (N_4131,N_3800,N_3547);
nand U4132 (N_4132,N_3067,N_3245);
nand U4133 (N_4133,N_3296,N_3171);
nor U4134 (N_4134,N_3082,N_3021);
nor U4135 (N_4135,N_3999,N_3290);
or U4136 (N_4136,N_3488,N_3933);
or U4137 (N_4137,N_3231,N_3582);
or U4138 (N_4138,N_3808,N_3796);
and U4139 (N_4139,N_3780,N_3081);
nand U4140 (N_4140,N_3129,N_3186);
and U4141 (N_4141,N_3149,N_3594);
or U4142 (N_4142,N_3916,N_3525);
nand U4143 (N_4143,N_3332,N_3947);
or U4144 (N_4144,N_3479,N_3912);
xor U4145 (N_4145,N_3318,N_3407);
xor U4146 (N_4146,N_3260,N_3414);
xor U4147 (N_4147,N_3773,N_3509);
nand U4148 (N_4148,N_3039,N_3286);
nand U4149 (N_4149,N_3439,N_3251);
and U4150 (N_4150,N_3986,N_3018);
or U4151 (N_4151,N_3815,N_3718);
and U4152 (N_4152,N_3352,N_3811);
and U4153 (N_4153,N_3430,N_3667);
nand U4154 (N_4154,N_3016,N_3087);
xor U4155 (N_4155,N_3785,N_3778);
and U4156 (N_4156,N_3958,N_3390);
xnor U4157 (N_4157,N_3176,N_3686);
and U4158 (N_4158,N_3890,N_3013);
or U4159 (N_4159,N_3258,N_3612);
nor U4160 (N_4160,N_3378,N_3209);
or U4161 (N_4161,N_3672,N_3804);
xnor U4162 (N_4162,N_3455,N_3484);
xnor U4163 (N_4163,N_3038,N_3089);
nor U4164 (N_4164,N_3281,N_3115);
and U4165 (N_4165,N_3593,N_3119);
xnor U4166 (N_4166,N_3697,N_3080);
nor U4167 (N_4167,N_3491,N_3898);
or U4168 (N_4168,N_3357,N_3988);
xor U4169 (N_4169,N_3777,N_3400);
or U4170 (N_4170,N_3969,N_3341);
or U4171 (N_4171,N_3058,N_3078);
and U4172 (N_4172,N_3391,N_3000);
and U4173 (N_4173,N_3066,N_3381);
nand U4174 (N_4174,N_3415,N_3575);
nor U4175 (N_4175,N_3436,N_3789);
nand U4176 (N_4176,N_3629,N_3042);
nand U4177 (N_4177,N_3295,N_3319);
and U4178 (N_4178,N_3472,N_3528);
nor U4179 (N_4179,N_3511,N_3714);
nor U4180 (N_4180,N_3840,N_3984);
nand U4181 (N_4181,N_3536,N_3563);
nor U4182 (N_4182,N_3566,N_3889);
xnor U4183 (N_4183,N_3433,N_3440);
xnor U4184 (N_4184,N_3835,N_3086);
and U4185 (N_4185,N_3589,N_3834);
and U4186 (N_4186,N_3202,N_3130);
nor U4187 (N_4187,N_3215,N_3316);
or U4188 (N_4188,N_3045,N_3333);
xor U4189 (N_4189,N_3812,N_3399);
nand U4190 (N_4190,N_3725,N_3841);
xnor U4191 (N_4191,N_3899,N_3469);
and U4192 (N_4192,N_3110,N_3540);
nor U4193 (N_4193,N_3532,N_3652);
nand U4194 (N_4194,N_3728,N_3530);
nor U4195 (N_4195,N_3734,N_3470);
xor U4196 (N_4196,N_3174,N_3814);
nor U4197 (N_4197,N_3387,N_3801);
and U4198 (N_4198,N_3845,N_3358);
nor U4199 (N_4199,N_3206,N_3830);
xor U4200 (N_4200,N_3405,N_3344);
nor U4201 (N_4201,N_3046,N_3041);
nor U4202 (N_4202,N_3451,N_3712);
nor U4203 (N_4203,N_3499,N_3673);
xnor U4204 (N_4204,N_3006,N_3114);
xnor U4205 (N_4205,N_3595,N_3264);
nor U4206 (N_4206,N_3416,N_3868);
or U4207 (N_4207,N_3448,N_3471);
nand U4208 (N_4208,N_3880,N_3053);
or U4209 (N_4209,N_3485,N_3124);
or U4210 (N_4210,N_3157,N_3627);
xor U4211 (N_4211,N_3715,N_3239);
nand U4212 (N_4212,N_3008,N_3025);
nor U4213 (N_4213,N_3489,N_3674);
and U4214 (N_4214,N_3903,N_3136);
or U4215 (N_4215,N_3059,N_3494);
and U4216 (N_4216,N_3247,N_3126);
nor U4217 (N_4217,N_3636,N_3709);
nor U4218 (N_4218,N_3475,N_3383);
nor U4219 (N_4219,N_3272,N_3591);
nand U4220 (N_4220,N_3579,N_3742);
and U4221 (N_4221,N_3904,N_3883);
nor U4222 (N_4222,N_3586,N_3546);
or U4223 (N_4223,N_3966,N_3514);
nor U4224 (N_4224,N_3681,N_3274);
and U4225 (N_4225,N_3398,N_3303);
or U4226 (N_4226,N_3873,N_3208);
or U4227 (N_4227,N_3458,N_3377);
nand U4228 (N_4228,N_3861,N_3668);
xnor U4229 (N_4229,N_3237,N_3805);
or U4230 (N_4230,N_3459,N_3516);
nand U4231 (N_4231,N_3246,N_3911);
and U4232 (N_4232,N_3824,N_3766);
and U4233 (N_4233,N_3610,N_3323);
xor U4234 (N_4234,N_3602,N_3401);
xnor U4235 (N_4235,N_3922,N_3664);
nand U4236 (N_4236,N_3498,N_3155);
nand U4237 (N_4237,N_3034,N_3759);
and U4238 (N_4238,N_3146,N_3077);
xnor U4239 (N_4239,N_3744,N_3973);
or U4240 (N_4240,N_3635,N_3037);
nand U4241 (N_4241,N_3419,N_3917);
and U4242 (N_4242,N_3663,N_3483);
and U4243 (N_4243,N_3836,N_3607);
nand U4244 (N_4244,N_3359,N_3022);
nor U4245 (N_4245,N_3996,N_3500);
nor U4246 (N_4246,N_3570,N_3665);
and U4247 (N_4247,N_3705,N_3148);
and U4248 (N_4248,N_3616,N_3870);
and U4249 (N_4249,N_3783,N_3014);
xor U4250 (N_4250,N_3887,N_3769);
nor U4251 (N_4251,N_3460,N_3189);
or U4252 (N_4252,N_3363,N_3724);
or U4253 (N_4253,N_3671,N_3346);
and U4254 (N_4254,N_3852,N_3963);
nor U4255 (N_4255,N_3659,N_3949);
xor U4256 (N_4256,N_3388,N_3467);
nor U4257 (N_4257,N_3275,N_3925);
nor U4258 (N_4258,N_3776,N_3023);
xnor U4259 (N_4259,N_3543,N_3446);
or U4260 (N_4260,N_3504,N_3490);
or U4261 (N_4261,N_3934,N_3505);
nor U4262 (N_4262,N_3366,N_3262);
xor U4263 (N_4263,N_3466,N_3818);
or U4264 (N_4264,N_3897,N_3879);
nor U4265 (N_4265,N_3657,N_3799);
nand U4266 (N_4266,N_3468,N_3810);
or U4267 (N_4267,N_3248,N_3866);
or U4268 (N_4268,N_3142,N_3666);
nor U4269 (N_4269,N_3097,N_3195);
nand U4270 (N_4270,N_3961,N_3254);
or U4271 (N_4271,N_3312,N_3355);
or U4272 (N_4272,N_3307,N_3994);
nand U4273 (N_4273,N_3902,N_3980);
or U4274 (N_4274,N_3070,N_3372);
and U4275 (N_4275,N_3179,N_3967);
and U4276 (N_4276,N_3685,N_3477);
nand U4277 (N_4277,N_3267,N_3828);
or U4278 (N_4278,N_3088,N_3955);
or U4279 (N_4279,N_3747,N_3227);
nor U4280 (N_4280,N_3906,N_3120);
nor U4281 (N_4281,N_3442,N_3974);
nor U4282 (N_4282,N_3753,N_3823);
nand U4283 (N_4283,N_3924,N_3600);
nand U4284 (N_4284,N_3716,N_3057);
xnor U4285 (N_4285,N_3677,N_3622);
nor U4286 (N_4286,N_3907,N_3633);
and U4287 (N_4287,N_3107,N_3761);
nor U4288 (N_4288,N_3676,N_3133);
nor U4289 (N_4289,N_3410,N_3645);
nor U4290 (N_4290,N_3535,N_3027);
or U4291 (N_4291,N_3743,N_3637);
and U4292 (N_4292,N_3310,N_3099);
nand U4293 (N_4293,N_3779,N_3959);
xnor U4294 (N_4294,N_3765,N_3920);
nand U4295 (N_4295,N_3412,N_3190);
or U4296 (N_4296,N_3482,N_3930);
and U4297 (N_4297,N_3205,N_3590);
xor U4298 (N_4298,N_3606,N_3886);
or U4299 (N_4299,N_3757,N_3749);
and U4300 (N_4300,N_3560,N_3919);
and U4301 (N_4301,N_3905,N_3909);
nor U4302 (N_4302,N_3772,N_3123);
nand U4303 (N_4303,N_3649,N_3619);
nor U4304 (N_4304,N_3257,N_3893);
xnor U4305 (N_4305,N_3223,N_3228);
nor U4306 (N_4306,N_3417,N_3557);
xnor U4307 (N_4307,N_3151,N_3703);
or U4308 (N_4308,N_3443,N_3571);
nor U4309 (N_4309,N_3878,N_3609);
nor U4310 (N_4310,N_3533,N_3968);
nor U4311 (N_4311,N_3214,N_3270);
nand U4312 (N_4312,N_3012,N_3002);
nand U4313 (N_4313,N_3108,N_3729);
nor U4314 (N_4314,N_3300,N_3217);
nor U4315 (N_4315,N_3017,N_3679);
and U4316 (N_4316,N_3813,N_3131);
nor U4317 (N_4317,N_3379,N_3970);
or U4318 (N_4318,N_3351,N_3877);
nor U4319 (N_4319,N_3085,N_3565);
or U4320 (N_4320,N_3691,N_3182);
and U4321 (N_4321,N_3869,N_3932);
or U4322 (N_4322,N_3882,N_3349);
or U4323 (N_4323,N_3550,N_3752);
nand U4324 (N_4324,N_3846,N_3213);
and U4325 (N_4325,N_3226,N_3347);
nor U4326 (N_4326,N_3438,N_3678);
nor U4327 (N_4327,N_3137,N_3976);
nor U4328 (N_4328,N_3764,N_3173);
xnor U4329 (N_4329,N_3203,N_3437);
nand U4330 (N_4330,N_3062,N_3867);
and U4331 (N_4331,N_3063,N_3428);
nor U4332 (N_4332,N_3127,N_3413);
and U4333 (N_4333,N_3957,N_3523);
nor U4334 (N_4334,N_3396,N_3269);
xnor U4335 (N_4335,N_3979,N_3857);
nand U4336 (N_4336,N_3983,N_3624);
and U4337 (N_4337,N_3162,N_3250);
nand U4338 (N_4338,N_3982,N_3112);
or U4339 (N_4339,N_3891,N_3096);
or U4340 (N_4340,N_3581,N_3009);
or U4341 (N_4341,N_3992,N_3314);
and U4342 (N_4342,N_3386,N_3161);
or U4343 (N_4343,N_3939,N_3620);
nand U4344 (N_4344,N_3936,N_3255);
xnor U4345 (N_4345,N_3763,N_3754);
and U4346 (N_4346,N_3855,N_3942);
nand U4347 (N_4347,N_3340,N_3617);
nor U4348 (N_4348,N_3741,N_3913);
xor U4349 (N_4349,N_3888,N_3908);
nand U4350 (N_4350,N_3074,N_3694);
and U4351 (N_4351,N_3402,N_3884);
nand U4352 (N_4352,N_3900,N_3004);
nand U4353 (N_4353,N_3313,N_3745);
nand U4354 (N_4354,N_3838,N_3225);
nand U4355 (N_4355,N_3894,N_3864);
xor U4356 (N_4356,N_3670,N_3564);
nor U4357 (N_4357,N_3348,N_3282);
xnor U4358 (N_4358,N_3060,N_3956);
nand U4359 (N_4359,N_3141,N_3507);
and U4360 (N_4360,N_3809,N_3851);
and U4361 (N_4361,N_3106,N_3628);
or U4362 (N_4362,N_3792,N_3597);
and U4363 (N_4363,N_3688,N_3315);
and U4364 (N_4364,N_3360,N_3298);
xor U4365 (N_4365,N_3722,N_3843);
nor U4366 (N_4366,N_3921,N_3901);
and U4367 (N_4367,N_3784,N_3831);
or U4368 (N_4368,N_3518,N_3181);
or U4369 (N_4369,N_3696,N_3263);
and U4370 (N_4370,N_3139,N_3625);
or U4371 (N_4371,N_3338,N_3972);
nor U4372 (N_4372,N_3125,N_3091);
and U4373 (N_4373,N_3345,N_3684);
or U4374 (N_4374,N_3738,N_3577);
nand U4375 (N_4375,N_3103,N_3403);
or U4376 (N_4376,N_3495,N_3335);
nand U4377 (N_4377,N_3844,N_3544);
or U4378 (N_4378,N_3997,N_3706);
nor U4379 (N_4379,N_3083,N_3285);
and U4380 (N_4380,N_3829,N_3229);
and U4381 (N_4381,N_3241,N_3760);
nand U4382 (N_4382,N_3232,N_3324);
and U4383 (N_4383,N_3702,N_3661);
xnor U4384 (N_4384,N_3853,N_3317);
nand U4385 (N_4385,N_3102,N_3559);
xnor U4386 (N_4386,N_3145,N_3711);
xor U4387 (N_4387,N_3463,N_3277);
or U4388 (N_4388,N_3662,N_3365);
or U4389 (N_4389,N_3618,N_3946);
xnor U4390 (N_4390,N_3240,N_3184);
and U4391 (N_4391,N_3854,N_3166);
nor U4392 (N_4392,N_3079,N_3199);
and U4393 (N_4393,N_3253,N_3929);
nand U4394 (N_4394,N_3698,N_3943);
or U4395 (N_4395,N_3508,N_3975);
xor U4396 (N_4396,N_3640,N_3212);
and U4397 (N_4397,N_3643,N_3481);
nand U4398 (N_4398,N_3519,N_3605);
xor U4399 (N_4399,N_3404,N_3178);
xor U4400 (N_4400,N_3660,N_3512);
nor U4401 (N_4401,N_3555,N_3862);
nand U4402 (N_4402,N_3069,N_3261);
and U4403 (N_4403,N_3603,N_3111);
nor U4404 (N_4404,N_3848,N_3651);
nand U4405 (N_4405,N_3787,N_3613);
nand U4406 (N_4406,N_3756,N_3750);
nor U4407 (N_4407,N_3580,N_3048);
and U4408 (N_4408,N_3521,N_3432);
nand U4409 (N_4409,N_3554,N_3169);
nand U4410 (N_4410,N_3429,N_3701);
and U4411 (N_4411,N_3821,N_3654);
or U4412 (N_4412,N_3029,N_3373);
xor U4413 (N_4413,N_3719,N_3768);
and U4414 (N_4414,N_3024,N_3293);
and U4415 (N_4415,N_3376,N_3950);
nor U4416 (N_4416,N_3762,N_3384);
nor U4417 (N_4417,N_3599,N_3531);
xor U4418 (N_4418,N_3271,N_3056);
xnor U4419 (N_4419,N_3826,N_3693);
or U4420 (N_4420,N_3551,N_3562);
nand U4421 (N_4421,N_3308,N_3200);
xor U4422 (N_4422,N_3450,N_3915);
and U4423 (N_4423,N_3336,N_3526);
and U4424 (N_4424,N_3802,N_3576);
and U4425 (N_4425,N_3389,N_3721);
or U4426 (N_4426,N_3708,N_3492);
or U4427 (N_4427,N_3737,N_3736);
or U4428 (N_4428,N_3863,N_3542);
nor U4429 (N_4429,N_3101,N_3306);
xnor U4430 (N_4430,N_3517,N_3100);
nor U4431 (N_4431,N_3578,N_3330);
nand U4432 (N_4432,N_3422,N_3740);
xor U4433 (N_4433,N_3896,N_3321);
nor U4434 (N_4434,N_3457,N_3180);
or U4435 (N_4435,N_3604,N_3680);
and U4436 (N_4436,N_3342,N_3675);
nand U4437 (N_4437,N_3952,N_3320);
or U4438 (N_4438,N_3138,N_3953);
nand U4439 (N_4439,N_3441,N_3364);
or U4440 (N_4440,N_3043,N_3552);
xnor U4441 (N_4441,N_3827,N_3937);
and U4442 (N_4442,N_3134,N_3188);
and U4443 (N_4443,N_3090,N_3689);
nor U4444 (N_4444,N_3026,N_3573);
or U4445 (N_4445,N_3276,N_3803);
xnor U4446 (N_4446,N_3717,N_3230);
and U4447 (N_4447,N_3790,N_3569);
nand U4448 (N_4448,N_3781,N_3522);
nand U4449 (N_4449,N_3454,N_3367);
xnor U4450 (N_4450,N_3732,N_3132);
and U4451 (N_4451,N_3881,N_3646);
nand U4452 (N_4452,N_3608,N_3339);
nor U4453 (N_4453,N_3175,N_3598);
xor U4454 (N_4454,N_3820,N_3197);
nor U4455 (N_4455,N_3035,N_3748);
and U4456 (N_4456,N_3601,N_3795);
or U4457 (N_4457,N_3183,N_3005);
nor U4458 (N_4458,N_3847,N_3064);
or U4459 (N_4459,N_3068,N_3639);
nand U4460 (N_4460,N_3545,N_3147);
nand U4461 (N_4461,N_3726,N_3105);
xnor U4462 (N_4462,N_3449,N_3774);
and U4463 (N_4463,N_3487,N_3287);
and U4464 (N_4464,N_3720,N_3001);
and U4465 (N_4465,N_3987,N_3918);
nand U4466 (N_4466,N_3242,N_3456);
and U4467 (N_4467,N_3003,N_3539);
and U4468 (N_4468,N_3529,N_3354);
and U4469 (N_4469,N_3093,N_3065);
and U4470 (N_4470,N_3095,N_3568);
nand U4471 (N_4471,N_3073,N_3735);
xnor U4472 (N_4472,N_3092,N_3256);
nand U4473 (N_4473,N_3288,N_3434);
nor U4474 (N_4474,N_3385,N_3656);
or U4475 (N_4475,N_3655,N_3370);
xnor U4476 (N_4476,N_3837,N_3755);
nor U4477 (N_4477,N_3788,N_3291);
and U4478 (N_4478,N_3474,N_3534);
and U4479 (N_4479,N_3541,N_3585);
and U4480 (N_4480,N_3650,N_3938);
nand U4481 (N_4481,N_3548,N_3051);
and U4482 (N_4482,N_3553,N_3019);
nand U4483 (N_4483,N_3690,N_3172);
nand U4484 (N_4484,N_3819,N_3832);
or U4485 (N_4485,N_3941,N_3871);
xor U4486 (N_4486,N_3634,N_3473);
nand U4487 (N_4487,N_3960,N_3614);
nor U4488 (N_4488,N_3167,N_3408);
nor U4489 (N_4489,N_3875,N_3993);
or U4490 (N_4490,N_3031,N_3177);
xor U4491 (N_4491,N_3244,N_3630);
xor U4492 (N_4492,N_3036,N_3856);
nand U4493 (N_4493,N_3040,N_3010);
nand U4494 (N_4494,N_3334,N_3168);
xor U4495 (N_4495,N_3648,N_3128);
nor U4496 (N_4496,N_3767,N_3746);
nor U4497 (N_4497,N_3926,N_3273);
nor U4498 (N_4498,N_3497,N_3322);
or U4499 (N_4499,N_3135,N_3931);
and U4500 (N_4500,N_3848,N_3530);
or U4501 (N_4501,N_3244,N_3582);
and U4502 (N_4502,N_3183,N_3031);
nor U4503 (N_4503,N_3942,N_3304);
and U4504 (N_4504,N_3225,N_3373);
nand U4505 (N_4505,N_3433,N_3379);
xor U4506 (N_4506,N_3155,N_3945);
and U4507 (N_4507,N_3727,N_3133);
and U4508 (N_4508,N_3272,N_3670);
or U4509 (N_4509,N_3460,N_3389);
or U4510 (N_4510,N_3010,N_3579);
xnor U4511 (N_4511,N_3699,N_3044);
and U4512 (N_4512,N_3729,N_3554);
and U4513 (N_4513,N_3534,N_3628);
xor U4514 (N_4514,N_3603,N_3568);
nand U4515 (N_4515,N_3760,N_3995);
nor U4516 (N_4516,N_3199,N_3318);
nand U4517 (N_4517,N_3387,N_3533);
or U4518 (N_4518,N_3637,N_3052);
nor U4519 (N_4519,N_3107,N_3066);
nand U4520 (N_4520,N_3000,N_3702);
nor U4521 (N_4521,N_3862,N_3942);
xnor U4522 (N_4522,N_3942,N_3619);
xor U4523 (N_4523,N_3796,N_3892);
nor U4524 (N_4524,N_3946,N_3323);
and U4525 (N_4525,N_3884,N_3685);
or U4526 (N_4526,N_3166,N_3467);
nor U4527 (N_4527,N_3415,N_3493);
and U4528 (N_4528,N_3817,N_3174);
nor U4529 (N_4529,N_3220,N_3502);
xnor U4530 (N_4530,N_3643,N_3812);
xnor U4531 (N_4531,N_3620,N_3466);
or U4532 (N_4532,N_3291,N_3687);
xnor U4533 (N_4533,N_3078,N_3846);
or U4534 (N_4534,N_3703,N_3465);
nand U4535 (N_4535,N_3627,N_3794);
or U4536 (N_4536,N_3867,N_3855);
nand U4537 (N_4537,N_3150,N_3760);
nor U4538 (N_4538,N_3054,N_3873);
nor U4539 (N_4539,N_3637,N_3406);
and U4540 (N_4540,N_3731,N_3933);
and U4541 (N_4541,N_3645,N_3274);
nor U4542 (N_4542,N_3654,N_3922);
nor U4543 (N_4543,N_3858,N_3320);
nor U4544 (N_4544,N_3772,N_3299);
or U4545 (N_4545,N_3783,N_3701);
or U4546 (N_4546,N_3432,N_3378);
and U4547 (N_4547,N_3488,N_3625);
or U4548 (N_4548,N_3988,N_3789);
xnor U4549 (N_4549,N_3061,N_3204);
and U4550 (N_4550,N_3067,N_3862);
xor U4551 (N_4551,N_3528,N_3661);
nand U4552 (N_4552,N_3801,N_3292);
nand U4553 (N_4553,N_3141,N_3838);
nor U4554 (N_4554,N_3460,N_3837);
nor U4555 (N_4555,N_3650,N_3973);
nor U4556 (N_4556,N_3809,N_3846);
nand U4557 (N_4557,N_3120,N_3159);
xor U4558 (N_4558,N_3198,N_3264);
and U4559 (N_4559,N_3734,N_3152);
or U4560 (N_4560,N_3619,N_3304);
and U4561 (N_4561,N_3108,N_3054);
and U4562 (N_4562,N_3661,N_3590);
nor U4563 (N_4563,N_3944,N_3088);
nor U4564 (N_4564,N_3178,N_3556);
nor U4565 (N_4565,N_3849,N_3562);
xnor U4566 (N_4566,N_3776,N_3772);
nand U4567 (N_4567,N_3535,N_3008);
nand U4568 (N_4568,N_3355,N_3066);
xor U4569 (N_4569,N_3892,N_3484);
or U4570 (N_4570,N_3297,N_3173);
xnor U4571 (N_4571,N_3130,N_3230);
or U4572 (N_4572,N_3289,N_3566);
nand U4573 (N_4573,N_3981,N_3062);
or U4574 (N_4574,N_3234,N_3695);
nand U4575 (N_4575,N_3349,N_3378);
and U4576 (N_4576,N_3430,N_3536);
nor U4577 (N_4577,N_3298,N_3256);
and U4578 (N_4578,N_3953,N_3164);
xor U4579 (N_4579,N_3187,N_3350);
nor U4580 (N_4580,N_3208,N_3568);
xor U4581 (N_4581,N_3716,N_3971);
nand U4582 (N_4582,N_3713,N_3310);
nor U4583 (N_4583,N_3319,N_3537);
nor U4584 (N_4584,N_3500,N_3709);
or U4585 (N_4585,N_3876,N_3056);
nand U4586 (N_4586,N_3908,N_3198);
nand U4587 (N_4587,N_3490,N_3791);
xor U4588 (N_4588,N_3046,N_3012);
and U4589 (N_4589,N_3596,N_3975);
nand U4590 (N_4590,N_3976,N_3407);
or U4591 (N_4591,N_3746,N_3039);
nor U4592 (N_4592,N_3220,N_3913);
or U4593 (N_4593,N_3061,N_3733);
nand U4594 (N_4594,N_3006,N_3725);
nand U4595 (N_4595,N_3735,N_3890);
nor U4596 (N_4596,N_3093,N_3123);
nor U4597 (N_4597,N_3418,N_3045);
nand U4598 (N_4598,N_3196,N_3050);
and U4599 (N_4599,N_3142,N_3385);
nor U4600 (N_4600,N_3071,N_3050);
nand U4601 (N_4601,N_3840,N_3083);
nor U4602 (N_4602,N_3874,N_3808);
xnor U4603 (N_4603,N_3889,N_3278);
nor U4604 (N_4604,N_3006,N_3339);
nor U4605 (N_4605,N_3104,N_3200);
or U4606 (N_4606,N_3535,N_3200);
or U4607 (N_4607,N_3924,N_3770);
or U4608 (N_4608,N_3495,N_3460);
nor U4609 (N_4609,N_3809,N_3797);
and U4610 (N_4610,N_3669,N_3174);
nand U4611 (N_4611,N_3579,N_3712);
nor U4612 (N_4612,N_3104,N_3491);
nor U4613 (N_4613,N_3071,N_3643);
and U4614 (N_4614,N_3460,N_3788);
and U4615 (N_4615,N_3651,N_3073);
nor U4616 (N_4616,N_3764,N_3203);
or U4617 (N_4617,N_3482,N_3632);
and U4618 (N_4618,N_3211,N_3866);
nor U4619 (N_4619,N_3625,N_3324);
or U4620 (N_4620,N_3782,N_3994);
xor U4621 (N_4621,N_3574,N_3792);
and U4622 (N_4622,N_3204,N_3957);
or U4623 (N_4623,N_3373,N_3573);
nor U4624 (N_4624,N_3080,N_3146);
xor U4625 (N_4625,N_3988,N_3730);
and U4626 (N_4626,N_3963,N_3823);
xnor U4627 (N_4627,N_3900,N_3864);
nand U4628 (N_4628,N_3170,N_3665);
or U4629 (N_4629,N_3926,N_3039);
nand U4630 (N_4630,N_3208,N_3187);
nor U4631 (N_4631,N_3054,N_3095);
and U4632 (N_4632,N_3046,N_3929);
nand U4633 (N_4633,N_3840,N_3453);
nor U4634 (N_4634,N_3210,N_3233);
or U4635 (N_4635,N_3896,N_3174);
nand U4636 (N_4636,N_3993,N_3415);
or U4637 (N_4637,N_3053,N_3603);
and U4638 (N_4638,N_3047,N_3707);
nand U4639 (N_4639,N_3429,N_3899);
or U4640 (N_4640,N_3545,N_3411);
xor U4641 (N_4641,N_3882,N_3037);
nand U4642 (N_4642,N_3037,N_3907);
nor U4643 (N_4643,N_3352,N_3566);
xor U4644 (N_4644,N_3512,N_3087);
and U4645 (N_4645,N_3571,N_3023);
xnor U4646 (N_4646,N_3898,N_3440);
and U4647 (N_4647,N_3839,N_3825);
nor U4648 (N_4648,N_3784,N_3636);
and U4649 (N_4649,N_3326,N_3571);
nand U4650 (N_4650,N_3327,N_3088);
or U4651 (N_4651,N_3319,N_3420);
xnor U4652 (N_4652,N_3141,N_3417);
nand U4653 (N_4653,N_3611,N_3717);
nor U4654 (N_4654,N_3237,N_3290);
xor U4655 (N_4655,N_3602,N_3385);
nand U4656 (N_4656,N_3193,N_3211);
xor U4657 (N_4657,N_3649,N_3873);
nor U4658 (N_4658,N_3518,N_3359);
and U4659 (N_4659,N_3335,N_3121);
nor U4660 (N_4660,N_3295,N_3803);
nand U4661 (N_4661,N_3948,N_3099);
nand U4662 (N_4662,N_3143,N_3246);
nor U4663 (N_4663,N_3595,N_3968);
and U4664 (N_4664,N_3981,N_3922);
nand U4665 (N_4665,N_3389,N_3298);
and U4666 (N_4666,N_3131,N_3876);
or U4667 (N_4667,N_3327,N_3522);
or U4668 (N_4668,N_3932,N_3263);
or U4669 (N_4669,N_3384,N_3226);
xnor U4670 (N_4670,N_3808,N_3926);
xnor U4671 (N_4671,N_3954,N_3238);
nor U4672 (N_4672,N_3744,N_3383);
or U4673 (N_4673,N_3270,N_3296);
nor U4674 (N_4674,N_3967,N_3092);
xnor U4675 (N_4675,N_3985,N_3240);
xnor U4676 (N_4676,N_3014,N_3674);
xor U4677 (N_4677,N_3487,N_3324);
or U4678 (N_4678,N_3009,N_3666);
or U4679 (N_4679,N_3496,N_3726);
or U4680 (N_4680,N_3818,N_3609);
xor U4681 (N_4681,N_3416,N_3345);
or U4682 (N_4682,N_3437,N_3615);
or U4683 (N_4683,N_3584,N_3832);
nor U4684 (N_4684,N_3470,N_3827);
nand U4685 (N_4685,N_3120,N_3235);
xnor U4686 (N_4686,N_3455,N_3773);
and U4687 (N_4687,N_3914,N_3303);
xor U4688 (N_4688,N_3680,N_3802);
nor U4689 (N_4689,N_3026,N_3240);
nor U4690 (N_4690,N_3628,N_3370);
nand U4691 (N_4691,N_3710,N_3376);
nand U4692 (N_4692,N_3555,N_3705);
or U4693 (N_4693,N_3996,N_3415);
xor U4694 (N_4694,N_3659,N_3865);
and U4695 (N_4695,N_3547,N_3099);
xnor U4696 (N_4696,N_3485,N_3747);
nor U4697 (N_4697,N_3372,N_3923);
or U4698 (N_4698,N_3334,N_3576);
or U4699 (N_4699,N_3536,N_3499);
nor U4700 (N_4700,N_3173,N_3135);
or U4701 (N_4701,N_3066,N_3883);
xnor U4702 (N_4702,N_3163,N_3714);
nand U4703 (N_4703,N_3775,N_3590);
and U4704 (N_4704,N_3683,N_3712);
nand U4705 (N_4705,N_3003,N_3491);
nor U4706 (N_4706,N_3140,N_3993);
xnor U4707 (N_4707,N_3579,N_3573);
or U4708 (N_4708,N_3704,N_3628);
or U4709 (N_4709,N_3650,N_3158);
or U4710 (N_4710,N_3440,N_3674);
nor U4711 (N_4711,N_3957,N_3685);
and U4712 (N_4712,N_3455,N_3120);
and U4713 (N_4713,N_3720,N_3278);
xor U4714 (N_4714,N_3783,N_3328);
or U4715 (N_4715,N_3404,N_3893);
xnor U4716 (N_4716,N_3170,N_3468);
and U4717 (N_4717,N_3694,N_3282);
nor U4718 (N_4718,N_3988,N_3553);
xor U4719 (N_4719,N_3172,N_3004);
nand U4720 (N_4720,N_3555,N_3878);
and U4721 (N_4721,N_3525,N_3330);
and U4722 (N_4722,N_3579,N_3859);
and U4723 (N_4723,N_3326,N_3171);
xor U4724 (N_4724,N_3286,N_3972);
nor U4725 (N_4725,N_3614,N_3237);
or U4726 (N_4726,N_3542,N_3879);
or U4727 (N_4727,N_3590,N_3675);
xor U4728 (N_4728,N_3174,N_3419);
xor U4729 (N_4729,N_3854,N_3511);
or U4730 (N_4730,N_3494,N_3121);
nor U4731 (N_4731,N_3891,N_3138);
and U4732 (N_4732,N_3900,N_3242);
xor U4733 (N_4733,N_3286,N_3104);
and U4734 (N_4734,N_3045,N_3923);
xnor U4735 (N_4735,N_3092,N_3406);
xor U4736 (N_4736,N_3008,N_3608);
and U4737 (N_4737,N_3291,N_3448);
and U4738 (N_4738,N_3928,N_3307);
xnor U4739 (N_4739,N_3699,N_3354);
or U4740 (N_4740,N_3145,N_3691);
nand U4741 (N_4741,N_3645,N_3615);
xnor U4742 (N_4742,N_3885,N_3371);
xnor U4743 (N_4743,N_3861,N_3317);
and U4744 (N_4744,N_3776,N_3960);
and U4745 (N_4745,N_3322,N_3488);
xor U4746 (N_4746,N_3428,N_3928);
and U4747 (N_4747,N_3601,N_3686);
xnor U4748 (N_4748,N_3416,N_3710);
nand U4749 (N_4749,N_3432,N_3306);
xor U4750 (N_4750,N_3481,N_3610);
xor U4751 (N_4751,N_3942,N_3545);
and U4752 (N_4752,N_3600,N_3543);
or U4753 (N_4753,N_3192,N_3539);
or U4754 (N_4754,N_3122,N_3499);
or U4755 (N_4755,N_3164,N_3988);
nand U4756 (N_4756,N_3200,N_3418);
and U4757 (N_4757,N_3450,N_3947);
xnor U4758 (N_4758,N_3174,N_3468);
xnor U4759 (N_4759,N_3344,N_3335);
and U4760 (N_4760,N_3262,N_3219);
or U4761 (N_4761,N_3389,N_3548);
nor U4762 (N_4762,N_3441,N_3780);
nor U4763 (N_4763,N_3335,N_3637);
nor U4764 (N_4764,N_3660,N_3832);
xor U4765 (N_4765,N_3623,N_3759);
and U4766 (N_4766,N_3365,N_3378);
nor U4767 (N_4767,N_3312,N_3285);
nand U4768 (N_4768,N_3423,N_3565);
nand U4769 (N_4769,N_3937,N_3579);
xnor U4770 (N_4770,N_3884,N_3624);
and U4771 (N_4771,N_3165,N_3695);
nor U4772 (N_4772,N_3056,N_3537);
nand U4773 (N_4773,N_3026,N_3048);
nand U4774 (N_4774,N_3302,N_3147);
or U4775 (N_4775,N_3895,N_3167);
or U4776 (N_4776,N_3544,N_3787);
and U4777 (N_4777,N_3893,N_3038);
nand U4778 (N_4778,N_3371,N_3191);
and U4779 (N_4779,N_3993,N_3176);
and U4780 (N_4780,N_3611,N_3380);
nor U4781 (N_4781,N_3463,N_3342);
or U4782 (N_4782,N_3412,N_3456);
or U4783 (N_4783,N_3661,N_3801);
nand U4784 (N_4784,N_3427,N_3770);
or U4785 (N_4785,N_3082,N_3049);
nand U4786 (N_4786,N_3845,N_3066);
nand U4787 (N_4787,N_3483,N_3478);
xnor U4788 (N_4788,N_3098,N_3335);
nand U4789 (N_4789,N_3292,N_3734);
xnor U4790 (N_4790,N_3865,N_3238);
or U4791 (N_4791,N_3462,N_3499);
nand U4792 (N_4792,N_3057,N_3244);
and U4793 (N_4793,N_3135,N_3938);
xor U4794 (N_4794,N_3418,N_3578);
or U4795 (N_4795,N_3266,N_3530);
nor U4796 (N_4796,N_3506,N_3101);
and U4797 (N_4797,N_3127,N_3847);
xnor U4798 (N_4798,N_3810,N_3255);
nor U4799 (N_4799,N_3997,N_3268);
nor U4800 (N_4800,N_3799,N_3126);
and U4801 (N_4801,N_3269,N_3683);
xnor U4802 (N_4802,N_3889,N_3582);
nor U4803 (N_4803,N_3548,N_3586);
or U4804 (N_4804,N_3174,N_3209);
nand U4805 (N_4805,N_3748,N_3800);
nand U4806 (N_4806,N_3977,N_3184);
or U4807 (N_4807,N_3036,N_3816);
or U4808 (N_4808,N_3650,N_3746);
nand U4809 (N_4809,N_3564,N_3507);
nand U4810 (N_4810,N_3580,N_3224);
nor U4811 (N_4811,N_3717,N_3312);
nand U4812 (N_4812,N_3400,N_3608);
nand U4813 (N_4813,N_3030,N_3539);
or U4814 (N_4814,N_3910,N_3852);
or U4815 (N_4815,N_3628,N_3328);
nand U4816 (N_4816,N_3401,N_3032);
xor U4817 (N_4817,N_3066,N_3995);
nand U4818 (N_4818,N_3366,N_3194);
nand U4819 (N_4819,N_3357,N_3385);
nand U4820 (N_4820,N_3839,N_3263);
or U4821 (N_4821,N_3804,N_3154);
xnor U4822 (N_4822,N_3013,N_3521);
or U4823 (N_4823,N_3233,N_3109);
nand U4824 (N_4824,N_3154,N_3586);
nor U4825 (N_4825,N_3489,N_3430);
and U4826 (N_4826,N_3631,N_3315);
nand U4827 (N_4827,N_3312,N_3396);
and U4828 (N_4828,N_3696,N_3835);
nand U4829 (N_4829,N_3614,N_3051);
nand U4830 (N_4830,N_3406,N_3472);
xnor U4831 (N_4831,N_3019,N_3485);
nor U4832 (N_4832,N_3072,N_3429);
nor U4833 (N_4833,N_3929,N_3118);
or U4834 (N_4834,N_3711,N_3236);
xnor U4835 (N_4835,N_3543,N_3576);
nand U4836 (N_4836,N_3715,N_3428);
nor U4837 (N_4837,N_3479,N_3824);
xnor U4838 (N_4838,N_3207,N_3513);
or U4839 (N_4839,N_3893,N_3674);
nor U4840 (N_4840,N_3510,N_3403);
and U4841 (N_4841,N_3826,N_3129);
and U4842 (N_4842,N_3921,N_3261);
nand U4843 (N_4843,N_3753,N_3157);
and U4844 (N_4844,N_3935,N_3503);
nor U4845 (N_4845,N_3803,N_3619);
xor U4846 (N_4846,N_3505,N_3633);
xor U4847 (N_4847,N_3467,N_3801);
nand U4848 (N_4848,N_3044,N_3920);
or U4849 (N_4849,N_3667,N_3068);
or U4850 (N_4850,N_3907,N_3616);
or U4851 (N_4851,N_3540,N_3965);
nand U4852 (N_4852,N_3182,N_3256);
xnor U4853 (N_4853,N_3636,N_3649);
and U4854 (N_4854,N_3299,N_3252);
or U4855 (N_4855,N_3858,N_3523);
nand U4856 (N_4856,N_3321,N_3840);
and U4857 (N_4857,N_3852,N_3698);
and U4858 (N_4858,N_3859,N_3188);
and U4859 (N_4859,N_3928,N_3310);
nor U4860 (N_4860,N_3572,N_3647);
and U4861 (N_4861,N_3616,N_3327);
and U4862 (N_4862,N_3706,N_3621);
nand U4863 (N_4863,N_3349,N_3461);
or U4864 (N_4864,N_3909,N_3904);
nor U4865 (N_4865,N_3597,N_3759);
and U4866 (N_4866,N_3212,N_3369);
nand U4867 (N_4867,N_3464,N_3583);
xor U4868 (N_4868,N_3430,N_3217);
nand U4869 (N_4869,N_3731,N_3086);
nand U4870 (N_4870,N_3550,N_3986);
nand U4871 (N_4871,N_3764,N_3189);
and U4872 (N_4872,N_3895,N_3490);
or U4873 (N_4873,N_3141,N_3654);
and U4874 (N_4874,N_3336,N_3683);
and U4875 (N_4875,N_3987,N_3538);
and U4876 (N_4876,N_3559,N_3405);
and U4877 (N_4877,N_3712,N_3260);
or U4878 (N_4878,N_3914,N_3943);
xor U4879 (N_4879,N_3075,N_3379);
nand U4880 (N_4880,N_3627,N_3744);
or U4881 (N_4881,N_3252,N_3348);
or U4882 (N_4882,N_3752,N_3741);
xnor U4883 (N_4883,N_3502,N_3213);
and U4884 (N_4884,N_3099,N_3718);
or U4885 (N_4885,N_3311,N_3144);
nor U4886 (N_4886,N_3171,N_3231);
xnor U4887 (N_4887,N_3551,N_3996);
nand U4888 (N_4888,N_3065,N_3809);
or U4889 (N_4889,N_3442,N_3995);
nand U4890 (N_4890,N_3215,N_3536);
xnor U4891 (N_4891,N_3579,N_3338);
nand U4892 (N_4892,N_3058,N_3502);
xor U4893 (N_4893,N_3507,N_3860);
nand U4894 (N_4894,N_3228,N_3054);
xnor U4895 (N_4895,N_3118,N_3290);
or U4896 (N_4896,N_3664,N_3474);
or U4897 (N_4897,N_3394,N_3293);
xnor U4898 (N_4898,N_3960,N_3687);
and U4899 (N_4899,N_3308,N_3500);
or U4900 (N_4900,N_3972,N_3814);
and U4901 (N_4901,N_3827,N_3534);
nor U4902 (N_4902,N_3706,N_3964);
or U4903 (N_4903,N_3823,N_3672);
nand U4904 (N_4904,N_3318,N_3645);
and U4905 (N_4905,N_3301,N_3469);
and U4906 (N_4906,N_3388,N_3276);
or U4907 (N_4907,N_3378,N_3288);
nand U4908 (N_4908,N_3683,N_3544);
or U4909 (N_4909,N_3269,N_3406);
or U4910 (N_4910,N_3835,N_3941);
nor U4911 (N_4911,N_3976,N_3677);
nand U4912 (N_4912,N_3525,N_3409);
and U4913 (N_4913,N_3569,N_3829);
xnor U4914 (N_4914,N_3221,N_3415);
or U4915 (N_4915,N_3705,N_3749);
and U4916 (N_4916,N_3454,N_3987);
xnor U4917 (N_4917,N_3769,N_3423);
or U4918 (N_4918,N_3758,N_3412);
nor U4919 (N_4919,N_3962,N_3143);
nor U4920 (N_4920,N_3811,N_3935);
xor U4921 (N_4921,N_3398,N_3334);
xnor U4922 (N_4922,N_3744,N_3355);
xnor U4923 (N_4923,N_3718,N_3547);
nor U4924 (N_4924,N_3795,N_3432);
and U4925 (N_4925,N_3947,N_3615);
nand U4926 (N_4926,N_3549,N_3171);
nor U4927 (N_4927,N_3550,N_3676);
xnor U4928 (N_4928,N_3633,N_3870);
and U4929 (N_4929,N_3846,N_3252);
or U4930 (N_4930,N_3667,N_3992);
nor U4931 (N_4931,N_3293,N_3855);
and U4932 (N_4932,N_3066,N_3538);
nand U4933 (N_4933,N_3617,N_3372);
nand U4934 (N_4934,N_3639,N_3131);
or U4935 (N_4935,N_3596,N_3959);
xor U4936 (N_4936,N_3660,N_3398);
and U4937 (N_4937,N_3630,N_3178);
nor U4938 (N_4938,N_3051,N_3846);
or U4939 (N_4939,N_3984,N_3450);
and U4940 (N_4940,N_3579,N_3544);
or U4941 (N_4941,N_3371,N_3771);
xnor U4942 (N_4942,N_3835,N_3771);
nand U4943 (N_4943,N_3583,N_3229);
nor U4944 (N_4944,N_3191,N_3628);
xor U4945 (N_4945,N_3106,N_3663);
xnor U4946 (N_4946,N_3136,N_3174);
or U4947 (N_4947,N_3672,N_3978);
or U4948 (N_4948,N_3082,N_3831);
xor U4949 (N_4949,N_3715,N_3635);
nor U4950 (N_4950,N_3940,N_3134);
or U4951 (N_4951,N_3804,N_3171);
nor U4952 (N_4952,N_3909,N_3143);
xnor U4953 (N_4953,N_3575,N_3806);
xnor U4954 (N_4954,N_3111,N_3572);
nor U4955 (N_4955,N_3097,N_3216);
and U4956 (N_4956,N_3104,N_3773);
xor U4957 (N_4957,N_3623,N_3048);
or U4958 (N_4958,N_3658,N_3615);
or U4959 (N_4959,N_3314,N_3406);
nor U4960 (N_4960,N_3914,N_3928);
nand U4961 (N_4961,N_3454,N_3865);
xnor U4962 (N_4962,N_3215,N_3402);
nand U4963 (N_4963,N_3146,N_3448);
xor U4964 (N_4964,N_3038,N_3149);
xor U4965 (N_4965,N_3887,N_3023);
or U4966 (N_4966,N_3454,N_3412);
nor U4967 (N_4967,N_3701,N_3969);
xor U4968 (N_4968,N_3067,N_3696);
or U4969 (N_4969,N_3370,N_3125);
and U4970 (N_4970,N_3386,N_3930);
and U4971 (N_4971,N_3182,N_3004);
nand U4972 (N_4972,N_3257,N_3386);
nand U4973 (N_4973,N_3227,N_3862);
and U4974 (N_4974,N_3425,N_3310);
nor U4975 (N_4975,N_3211,N_3852);
nor U4976 (N_4976,N_3726,N_3367);
nand U4977 (N_4977,N_3345,N_3101);
or U4978 (N_4978,N_3096,N_3123);
and U4979 (N_4979,N_3361,N_3827);
xor U4980 (N_4980,N_3701,N_3253);
xnor U4981 (N_4981,N_3362,N_3693);
xor U4982 (N_4982,N_3259,N_3126);
nand U4983 (N_4983,N_3571,N_3973);
or U4984 (N_4984,N_3978,N_3648);
or U4985 (N_4985,N_3229,N_3089);
nor U4986 (N_4986,N_3885,N_3343);
or U4987 (N_4987,N_3066,N_3407);
or U4988 (N_4988,N_3158,N_3761);
or U4989 (N_4989,N_3360,N_3784);
xnor U4990 (N_4990,N_3720,N_3983);
xor U4991 (N_4991,N_3951,N_3580);
nand U4992 (N_4992,N_3236,N_3533);
nand U4993 (N_4993,N_3429,N_3559);
nor U4994 (N_4994,N_3718,N_3409);
xor U4995 (N_4995,N_3351,N_3233);
nor U4996 (N_4996,N_3120,N_3568);
nor U4997 (N_4997,N_3771,N_3972);
and U4998 (N_4998,N_3523,N_3222);
or U4999 (N_4999,N_3544,N_3576);
nor U5000 (N_5000,N_4700,N_4370);
nand U5001 (N_5001,N_4800,N_4677);
or U5002 (N_5002,N_4132,N_4092);
xor U5003 (N_5003,N_4515,N_4076);
or U5004 (N_5004,N_4712,N_4701);
or U5005 (N_5005,N_4178,N_4436);
nand U5006 (N_5006,N_4763,N_4792);
or U5007 (N_5007,N_4441,N_4155);
or U5008 (N_5008,N_4880,N_4285);
nor U5009 (N_5009,N_4585,N_4380);
nand U5010 (N_5010,N_4140,N_4552);
nor U5011 (N_5011,N_4806,N_4799);
and U5012 (N_5012,N_4575,N_4022);
or U5013 (N_5013,N_4428,N_4730);
nand U5014 (N_5014,N_4098,N_4029);
xnor U5015 (N_5015,N_4936,N_4376);
nor U5016 (N_5016,N_4233,N_4562);
nand U5017 (N_5017,N_4391,N_4169);
and U5018 (N_5018,N_4829,N_4406);
nor U5019 (N_5019,N_4708,N_4044);
nor U5020 (N_5020,N_4726,N_4909);
nand U5021 (N_5021,N_4296,N_4264);
or U5022 (N_5022,N_4818,N_4058);
and U5023 (N_5023,N_4008,N_4652);
nor U5024 (N_5024,N_4422,N_4332);
xnor U5025 (N_5025,N_4702,N_4041);
nor U5026 (N_5026,N_4350,N_4364);
nand U5027 (N_5027,N_4717,N_4019);
nor U5028 (N_5028,N_4703,N_4995);
xor U5029 (N_5029,N_4868,N_4555);
nand U5030 (N_5030,N_4247,N_4479);
xnor U5031 (N_5031,N_4639,N_4776);
nand U5032 (N_5032,N_4601,N_4823);
nor U5033 (N_5033,N_4931,N_4745);
nor U5034 (N_5034,N_4579,N_4576);
or U5035 (N_5035,N_4068,N_4084);
xor U5036 (N_5036,N_4257,N_4609);
and U5037 (N_5037,N_4622,N_4172);
nor U5038 (N_5038,N_4779,N_4404);
nor U5039 (N_5039,N_4822,N_4293);
nor U5040 (N_5040,N_4542,N_4787);
nand U5041 (N_5041,N_4521,N_4720);
nand U5042 (N_5042,N_4281,N_4001);
or U5043 (N_5043,N_4419,N_4292);
nand U5044 (N_5044,N_4706,N_4036);
or U5045 (N_5045,N_4690,N_4594);
and U5046 (N_5046,N_4379,N_4308);
nor U5047 (N_5047,N_4989,N_4572);
nor U5048 (N_5048,N_4802,N_4060);
and U5049 (N_5049,N_4235,N_4105);
nor U5050 (N_5050,N_4213,N_4026);
and U5051 (N_5051,N_4516,N_4333);
and U5052 (N_5052,N_4083,N_4725);
or U5053 (N_5053,N_4948,N_4988);
and U5054 (N_5054,N_4094,N_4009);
xor U5055 (N_5055,N_4052,N_4306);
or U5056 (N_5056,N_4385,N_4063);
xor U5057 (N_5057,N_4569,N_4446);
nor U5058 (N_5058,N_4692,N_4961);
xnor U5059 (N_5059,N_4359,N_4927);
nor U5060 (N_5060,N_4892,N_4173);
and U5061 (N_5061,N_4015,N_4604);
nand U5062 (N_5062,N_4963,N_4170);
or U5063 (N_5063,N_4560,N_4512);
and U5064 (N_5064,N_4635,N_4828);
or U5065 (N_5065,N_4513,N_4163);
and U5066 (N_5066,N_4318,N_4917);
or U5067 (N_5067,N_4537,N_4672);
or U5068 (N_5068,N_4805,N_4118);
or U5069 (N_5069,N_4732,N_4856);
and U5070 (N_5070,N_4298,N_4532);
and U5071 (N_5071,N_4746,N_4326);
nor U5072 (N_5072,N_4231,N_4261);
xor U5073 (N_5073,N_4388,N_4045);
nand U5074 (N_5074,N_4352,N_4403);
nand U5075 (N_5075,N_4345,N_4288);
or U5076 (N_5076,N_4766,N_4518);
nor U5077 (N_5077,N_4028,N_4954);
nand U5078 (N_5078,N_4517,N_4279);
and U5079 (N_5079,N_4833,N_4251);
xor U5080 (N_5080,N_4638,N_4875);
nor U5081 (N_5081,N_4758,N_4151);
nand U5082 (N_5082,N_4459,N_4048);
nand U5083 (N_5083,N_4295,N_4487);
xor U5084 (N_5084,N_4874,N_4410);
and U5085 (N_5085,N_4003,N_4775);
or U5086 (N_5086,N_4119,N_4592);
or U5087 (N_5087,N_4112,N_4901);
or U5088 (N_5088,N_4080,N_4885);
xnor U5089 (N_5089,N_4738,N_4887);
and U5090 (N_5090,N_4584,N_4777);
nor U5091 (N_5091,N_4567,N_4733);
xor U5092 (N_5092,N_4207,N_4329);
xnor U5093 (N_5093,N_4696,N_4788);
xor U5094 (N_5094,N_4017,N_4774);
xor U5095 (N_5095,N_4244,N_4042);
xor U5096 (N_5096,N_4289,N_4801);
and U5097 (N_5097,N_4740,N_4239);
and U5098 (N_5098,N_4707,N_4387);
nand U5099 (N_5099,N_4016,N_4483);
nand U5100 (N_5100,N_4586,N_4934);
nor U5101 (N_5101,N_4946,N_4122);
nor U5102 (N_5102,N_4697,N_4375);
and U5103 (N_5103,N_4138,N_4915);
and U5104 (N_5104,N_4854,N_4368);
nor U5105 (N_5105,N_4103,N_4722);
xnor U5106 (N_5106,N_4808,N_4627);
or U5107 (N_5107,N_4574,N_4541);
nand U5108 (N_5108,N_4500,N_4291);
nand U5109 (N_5109,N_4599,N_4321);
or U5110 (N_5110,N_4014,N_4924);
and U5111 (N_5111,N_4844,N_4759);
or U5112 (N_5112,N_4495,N_4680);
xnor U5113 (N_5113,N_4011,N_4024);
or U5114 (N_5114,N_4167,N_4382);
nor U5115 (N_5115,N_4554,N_4784);
xor U5116 (N_5116,N_4331,N_4741);
xor U5117 (N_5117,N_4681,N_4614);
nand U5118 (N_5118,N_4234,N_4619);
nor U5119 (N_5119,N_4715,N_4424);
xnor U5120 (N_5120,N_4904,N_4222);
nor U5121 (N_5121,N_4872,N_4451);
nor U5122 (N_5122,N_4563,N_4663);
nand U5123 (N_5123,N_4837,N_4282);
or U5124 (N_5124,N_4952,N_4496);
xor U5125 (N_5125,N_4531,N_4748);
nor U5126 (N_5126,N_4623,N_4429);
or U5127 (N_5127,N_4863,N_4477);
or U5128 (N_5128,N_4378,N_4543);
or U5129 (N_5129,N_4883,N_4461);
nand U5130 (N_5130,N_4632,N_4353);
or U5131 (N_5131,N_4535,N_4152);
nor U5132 (N_5132,N_4618,N_4159);
and U5133 (N_5133,N_4457,N_4998);
nand U5134 (N_5134,N_4179,N_4107);
nor U5135 (N_5135,N_4010,N_4383);
xor U5136 (N_5136,N_4791,N_4462);
and U5137 (N_5137,N_4843,N_4216);
and U5138 (N_5138,N_4476,N_4488);
and U5139 (N_5139,N_4611,N_4896);
nor U5140 (N_5140,N_4301,N_4121);
and U5141 (N_5141,N_4556,N_4120);
nand U5142 (N_5142,N_4405,N_4492);
or U5143 (N_5143,N_4072,N_4069);
nor U5144 (N_5144,N_4208,N_4734);
xnor U5145 (N_5145,N_4037,N_4302);
or U5146 (N_5146,N_4276,N_4662);
nor U5147 (N_5147,N_4530,N_4499);
xnor U5148 (N_5148,N_4631,N_4714);
or U5149 (N_5149,N_4377,N_4034);
xnor U5150 (N_5150,N_4689,N_4830);
nand U5151 (N_5151,N_4249,N_4187);
xnor U5152 (N_5152,N_4253,N_4996);
nand U5153 (N_5153,N_4657,N_4294);
or U5154 (N_5154,N_4711,N_4900);
nor U5155 (N_5155,N_4994,N_4974);
or U5156 (N_5156,N_4633,N_4005);
xnor U5157 (N_5157,N_4894,N_4990);
or U5158 (N_5158,N_4547,N_4964);
and U5159 (N_5159,N_4897,N_4782);
xnor U5160 (N_5160,N_4686,N_4438);
or U5161 (N_5161,N_4643,N_4693);
or U5162 (N_5162,N_4440,N_4523);
nor U5163 (N_5163,N_4270,N_4608);
and U5164 (N_5164,N_4903,N_4030);
nand U5165 (N_5165,N_4205,N_4088);
nand U5166 (N_5166,N_4256,N_4570);
nor U5167 (N_5167,N_4344,N_4199);
or U5168 (N_5168,N_4636,N_4942);
nand U5169 (N_5169,N_4324,N_4360);
nor U5170 (N_5170,N_4735,N_4212);
and U5171 (N_5171,N_4668,N_4506);
and U5172 (N_5172,N_4816,N_4445);
xnor U5173 (N_5173,N_4685,N_4906);
nor U5174 (N_5174,N_4347,N_4300);
or U5175 (N_5175,N_4188,N_4947);
nand U5176 (N_5176,N_4136,N_4933);
xnor U5177 (N_5177,N_4842,N_4031);
xor U5178 (N_5178,N_4561,N_4878);
nor U5179 (N_5179,N_4907,N_4337);
nor U5180 (N_5180,N_4923,N_4620);
and U5181 (N_5181,N_4047,N_4831);
nand U5182 (N_5182,N_4412,N_4480);
nor U5183 (N_5183,N_4435,N_4507);
xnor U5184 (N_5184,N_4115,N_4126);
nor U5185 (N_5185,N_4443,N_4057);
and U5186 (N_5186,N_4351,N_4154);
and U5187 (N_5187,N_4168,N_4000);
xnor U5188 (N_5188,N_4241,N_4991);
and U5189 (N_5189,N_4284,N_4973);
xnor U5190 (N_5190,N_4665,N_4046);
xnor U5191 (N_5191,N_4390,N_4340);
nand U5192 (N_5192,N_4413,N_4919);
or U5193 (N_5193,N_4603,N_4316);
xor U5194 (N_5194,N_4583,N_4674);
xor U5195 (N_5195,N_4660,N_4983);
and U5196 (N_5196,N_4240,N_4882);
nor U5197 (N_5197,N_4846,N_4203);
nand U5198 (N_5198,N_4771,N_4097);
xor U5199 (N_5199,N_4021,N_4020);
xnor U5200 (N_5200,N_4976,N_4054);
nor U5201 (N_5201,N_4966,N_4040);
and U5202 (N_5202,N_4557,N_4006);
xnor U5203 (N_5203,N_4381,N_4165);
and U5204 (N_5204,N_4879,N_4104);
xnor U5205 (N_5205,N_4366,N_4566);
nand U5206 (N_5206,N_4079,N_4867);
and U5207 (N_5207,N_4613,N_4237);
or U5208 (N_5208,N_4486,N_4605);
nand U5209 (N_5209,N_4786,N_4204);
nand U5210 (N_5210,N_4941,N_4224);
nand U5211 (N_5211,N_4666,N_4400);
xnor U5212 (N_5212,N_4023,N_4073);
nor U5213 (N_5213,N_4025,N_4386);
or U5214 (N_5214,N_4481,N_4817);
nor U5215 (N_5215,N_4432,N_4433);
xor U5216 (N_5216,N_4891,N_4250);
nand U5217 (N_5217,N_4968,N_4218);
and U5218 (N_5218,N_4580,N_4625);
nand U5219 (N_5219,N_4893,N_4252);
and U5220 (N_5220,N_4414,N_4447);
nand U5221 (N_5221,N_4095,N_4290);
or U5222 (N_5222,N_4164,N_4191);
nand U5223 (N_5223,N_4049,N_4582);
nor U5224 (N_5224,N_4129,N_4194);
nor U5225 (N_5225,N_4669,N_4962);
nand U5226 (N_5226,N_4392,N_4033);
xor U5227 (N_5227,N_4472,N_4245);
and U5228 (N_5228,N_4754,N_4372);
and U5229 (N_5229,N_4491,N_4320);
or U5230 (N_5230,N_4463,N_4971);
and U5231 (N_5231,N_4789,N_4215);
xnor U5232 (N_5232,N_4145,N_4803);
xor U5233 (N_5233,N_4371,N_4160);
xor U5234 (N_5234,N_4478,N_4664);
or U5235 (N_5235,N_4313,N_4794);
nand U5236 (N_5236,N_4336,N_4408);
nand U5237 (N_5237,N_4474,N_4248);
and U5238 (N_5238,N_4813,N_4980);
or U5239 (N_5239,N_4865,N_4807);
nor U5240 (N_5240,N_4354,N_4394);
and U5241 (N_5241,N_4930,N_4004);
nor U5242 (N_5242,N_4260,N_4940);
nor U5243 (N_5243,N_4196,N_4373);
nor U5244 (N_5244,N_4007,N_4577);
and U5245 (N_5245,N_4658,N_4319);
or U5246 (N_5246,N_4910,N_4795);
and U5247 (N_5247,N_4545,N_4230);
nand U5248 (N_5248,N_4881,N_4065);
nand U5249 (N_5249,N_4415,N_4838);
nand U5250 (N_5250,N_4473,N_4314);
xor U5251 (N_5251,N_4287,N_4678);
xor U5252 (N_5252,N_4661,N_4420);
or U5253 (N_5253,N_4108,N_4258);
and U5254 (N_5254,N_4077,N_4699);
or U5255 (N_5255,N_4629,N_4993);
or U5256 (N_5256,N_4659,N_4465);
or U5257 (N_5257,N_4694,N_4695);
nor U5258 (N_5258,N_4475,N_4090);
or U5259 (N_5259,N_4796,N_4275);
and U5260 (N_5260,N_4853,N_4158);
or U5261 (N_5261,N_4862,N_4839);
nor U5262 (N_5262,N_4781,N_4427);
or U5263 (N_5263,N_4525,N_4851);
and U5264 (N_5264,N_4265,N_4467);
and U5265 (N_5265,N_4826,N_4626);
or U5266 (N_5266,N_4317,N_4790);
or U5267 (N_5267,N_4002,N_4425);
xor U5268 (N_5268,N_4602,N_4100);
nor U5269 (N_5269,N_4598,N_4731);
or U5270 (N_5270,N_4510,N_4769);
nand U5271 (N_5271,N_4895,N_4322);
and U5272 (N_5272,N_4624,N_4220);
nor U5273 (N_5273,N_4857,N_4819);
nand U5274 (N_5274,N_4217,N_4274);
nand U5275 (N_5275,N_4484,N_4667);
xnor U5276 (N_5276,N_4012,N_4013);
or U5277 (N_5277,N_4349,N_4655);
xor U5278 (N_5278,N_4367,N_4229);
and U5279 (N_5279,N_4809,N_4426);
xor U5280 (N_5280,N_4951,N_4106);
xnor U5281 (N_5281,N_4018,N_4630);
xnor U5282 (N_5282,N_4650,N_4460);
nor U5283 (N_5283,N_4744,N_4705);
nor U5284 (N_5284,N_4812,N_4442);
and U5285 (N_5285,N_4202,N_4185);
xnor U5286 (N_5286,N_4497,N_4634);
and U5287 (N_5287,N_4798,N_4847);
or U5288 (N_5288,N_4670,N_4710);
and U5289 (N_5289,N_4671,N_4965);
and U5290 (N_5290,N_4468,N_4223);
and U5291 (N_5291,N_4102,N_4133);
and U5292 (N_5292,N_4197,N_4698);
nor U5293 (N_5293,N_4395,N_4890);
and U5294 (N_5294,N_4482,N_4565);
and U5295 (N_5295,N_4780,N_4494);
or U5296 (N_5296,N_4228,N_4546);
nor U5297 (N_5297,N_4498,N_4960);
or U5298 (N_5298,N_4870,N_4551);
or U5299 (N_5299,N_4723,N_4315);
and U5300 (N_5300,N_4511,N_4299);
xnor U5301 (N_5301,N_4534,N_4417);
or U5302 (N_5302,N_4922,N_4981);
and U5303 (N_5303,N_4310,N_4593);
and U5304 (N_5304,N_4564,N_4211);
and U5305 (N_5305,N_4409,N_4356);
xnor U5306 (N_5306,N_4082,N_4682);
or U5307 (N_5307,N_4458,N_4135);
and U5308 (N_5308,N_4729,N_4673);
xnor U5309 (N_5309,N_4066,N_4820);
xnor U5310 (N_5310,N_4411,N_4157);
and U5311 (N_5311,N_4840,N_4762);
xnor U5312 (N_5312,N_4526,N_4921);
nor U5313 (N_5313,N_4263,N_4266);
or U5314 (N_5314,N_4821,N_4760);
and U5315 (N_5315,N_4254,N_4918);
xnor U5316 (N_5316,N_4027,N_4713);
xnor U5317 (N_5317,N_4724,N_4956);
or U5318 (N_5318,N_4550,N_4911);
and U5319 (N_5319,N_4825,N_4186);
and U5320 (N_5320,N_4286,N_4852);
nor U5321 (N_5321,N_4916,N_4062);
or U5322 (N_5322,N_4398,N_4876);
nor U5323 (N_5323,N_4501,N_4452);
nor U5324 (N_5324,N_4719,N_4268);
nor U5325 (N_5325,N_4110,N_4038);
nor U5326 (N_5326,N_4143,N_4978);
nor U5327 (N_5327,N_4437,N_4600);
xnor U5328 (N_5328,N_4397,N_4929);
nor U5329 (N_5329,N_4125,N_4166);
nand U5330 (N_5330,N_4520,N_4985);
nand U5331 (N_5331,N_4358,N_4573);
nor U5332 (N_5332,N_4146,N_4716);
nand U5333 (N_5333,N_4055,N_4174);
nand U5334 (N_5334,N_4553,N_4148);
nor U5335 (N_5335,N_4075,N_4841);
and U5336 (N_5336,N_4529,N_4908);
and U5337 (N_5337,N_4051,N_4768);
nand U5338 (N_5338,N_4325,N_4912);
xnor U5339 (N_5339,N_4621,N_4374);
xnor U5340 (N_5340,N_4928,N_4651);
or U5341 (N_5341,N_4312,N_4597);
or U5342 (N_5342,N_4053,N_4858);
nand U5343 (N_5343,N_4471,N_4195);
nor U5344 (N_5344,N_4640,N_4679);
and U5345 (N_5345,N_4539,N_4469);
nor U5346 (N_5346,N_4309,N_4259);
or U5347 (N_5347,N_4342,N_4935);
nor U5348 (N_5348,N_4992,N_4864);
or U5349 (N_5349,N_4176,N_4866);
xnor U5350 (N_5350,N_4454,N_4262);
or U5351 (N_5351,N_4430,N_4902);
xor U5352 (N_5352,N_4238,N_4363);
and U5353 (N_5353,N_4399,N_4607);
xor U5354 (N_5354,N_4718,N_4558);
nor U5355 (N_5355,N_4785,N_4641);
nor U5356 (N_5356,N_4721,N_4214);
and U5357 (N_5357,N_4849,N_4323);
nor U5358 (N_5358,N_4778,N_4226);
xnor U5359 (N_5359,N_4939,N_4704);
nor U5360 (N_5360,N_4749,N_4335);
and U5361 (N_5361,N_4615,N_4117);
xor U5362 (N_5362,N_4127,N_4078);
and U5363 (N_5363,N_4180,N_4855);
xnor U5364 (N_5364,N_4210,N_4134);
xor U5365 (N_5365,N_4764,N_4182);
and U5366 (N_5366,N_4987,N_4181);
or U5367 (N_5367,N_4977,N_4175);
nor U5368 (N_5368,N_4085,N_4861);
and U5369 (N_5369,N_4591,N_4765);
nand U5370 (N_5370,N_4848,N_4969);
or U5371 (N_5371,N_4743,N_4559);
nand U5372 (N_5372,N_4141,N_4389);
nand U5373 (N_5373,N_4815,N_4087);
nand U5374 (N_5374,N_4549,N_4177);
xnor U5375 (N_5375,N_4470,N_4957);
xnor U5376 (N_5376,N_4810,N_4431);
or U5377 (N_5377,N_4311,N_4691);
nor U5378 (N_5378,N_4937,N_4423);
nor U5379 (N_5379,N_4343,N_4114);
or U5380 (N_5380,N_4514,N_4944);
or U5381 (N_5381,N_4147,N_4225);
nand U5382 (N_5382,N_4889,N_4654);
xnor U5383 (N_5383,N_4967,N_4384);
or U5384 (N_5384,N_4035,N_4091);
xnor U5385 (N_5385,N_4756,N_4093);
or U5386 (N_5386,N_4219,N_4884);
or U5387 (N_5387,N_4124,N_4307);
nand U5388 (N_5388,N_4271,N_4544);
and U5389 (N_5389,N_4355,N_4571);
xor U5390 (N_5390,N_4074,N_4149);
and U5391 (N_5391,N_4131,N_4757);
or U5392 (N_5392,N_4606,N_4056);
or U5393 (N_5393,N_4059,N_4824);
nor U5394 (N_5394,N_4950,N_4836);
or U5395 (N_5395,N_4648,N_4039);
xnor U5396 (N_5396,N_4588,N_4772);
or U5397 (N_5397,N_4522,N_4505);
or U5398 (N_5398,N_4153,N_4297);
xor U5399 (N_5399,N_4502,N_4448);
nand U5400 (N_5400,N_4183,N_4061);
and U5401 (N_5401,N_4341,N_4267);
nand U5402 (N_5402,N_4396,N_4859);
nand U5403 (N_5403,N_4455,N_4596);
or U5404 (N_5404,N_4401,N_4783);
nor U5405 (N_5405,N_4914,N_4845);
or U5406 (N_5406,N_4687,N_4466);
nand U5407 (N_5407,N_4755,N_4305);
and U5408 (N_5408,N_4644,N_4653);
nor U5409 (N_5409,N_4972,N_4508);
nand U5410 (N_5410,N_4338,N_4444);
and U5411 (N_5411,N_4676,N_4303);
nand U5412 (N_5412,N_4421,N_4277);
xor U5413 (N_5413,N_4984,N_4886);
and U5414 (N_5414,N_4986,N_4450);
or U5415 (N_5415,N_4959,N_4926);
and U5416 (N_5416,N_4688,N_4835);
nor U5417 (N_5417,N_4278,N_4888);
and U5418 (N_5418,N_4871,N_4128);
or U5419 (N_5419,N_4970,N_4184);
nor U5420 (N_5420,N_4675,N_4099);
and U5421 (N_5421,N_4190,N_4590);
or U5422 (N_5422,N_4932,N_4348);
nor U5423 (N_5423,N_4761,N_4130);
nor U5424 (N_5424,N_4150,N_4346);
xnor U5425 (N_5425,N_4067,N_4171);
nand U5426 (N_5426,N_4628,N_4490);
nor U5427 (N_5427,N_4123,N_4209);
nor U5428 (N_5428,N_4357,N_4101);
nor U5429 (N_5429,N_4109,N_4709);
nand U5430 (N_5430,N_4905,N_4489);
nand U5431 (N_5431,N_4361,N_4945);
xnor U5432 (N_5432,N_4578,N_4834);
and U5433 (N_5433,N_4649,N_4485);
nand U5434 (N_5434,N_4739,N_4246);
xor U5435 (N_5435,N_4144,N_4873);
or U5436 (N_5436,N_4747,N_4943);
and U5437 (N_5437,N_4232,N_4524);
xor U5438 (N_5438,N_4587,N_4742);
and U5439 (N_5439,N_4434,N_4949);
nand U5440 (N_5440,N_4111,N_4767);
and U5441 (N_5441,N_4504,N_4439);
nand U5442 (N_5442,N_4979,N_4925);
and U5443 (N_5443,N_4750,N_4201);
nor U5444 (N_5444,N_4913,N_4527);
and U5445 (N_5445,N_4538,N_4200);
nand U5446 (N_5446,N_4533,N_4860);
xor U5447 (N_5447,N_4955,N_4221);
and U5448 (N_5448,N_4206,N_4850);
xnor U5449 (N_5449,N_4832,N_4242);
nor U5450 (N_5450,N_4683,N_4456);
or U5451 (N_5451,N_4064,N_4797);
and U5452 (N_5452,N_4161,N_4402);
or U5453 (N_5453,N_4548,N_4043);
or U5454 (N_5454,N_4814,N_4449);
xnor U5455 (N_5455,N_4568,N_4751);
xor U5456 (N_5456,N_4493,N_4595);
xor U5457 (N_5457,N_4137,N_4536);
nand U5458 (N_5458,N_4339,N_4938);
or U5459 (N_5459,N_4328,N_4139);
nand U5460 (N_5460,N_4958,N_4081);
xnor U5461 (N_5461,N_4645,N_4519);
nor U5462 (N_5462,N_4503,N_4273);
xor U5463 (N_5463,N_4727,N_4113);
nand U5464 (N_5464,N_4362,N_4617);
nand U5465 (N_5465,N_4243,N_4071);
and U5466 (N_5466,N_4581,N_4156);
nand U5467 (N_5467,N_4192,N_4616);
xnor U5468 (N_5468,N_4280,N_4330);
nand U5469 (N_5469,N_4684,N_4236);
nor U5470 (N_5470,N_4656,N_4975);
and U5471 (N_5471,N_4827,N_4464);
xnor U5472 (N_5472,N_4416,N_4198);
nor U5473 (N_5473,N_4283,N_4877);
nand U5474 (N_5474,N_4920,N_4982);
and U5475 (N_5475,N_4753,N_4142);
xnor U5476 (N_5476,N_4193,N_4811);
nor U5477 (N_5477,N_4773,N_4086);
nand U5478 (N_5478,N_4793,N_4869);
nor U5479 (N_5479,N_4646,N_4334);
xnor U5480 (N_5480,N_4637,N_4269);
nand U5481 (N_5481,N_4642,N_4162);
or U5482 (N_5482,N_4050,N_4032);
nor U5483 (N_5483,N_4189,N_4393);
or U5484 (N_5484,N_4736,N_4418);
xor U5485 (N_5485,N_4899,N_4770);
or U5486 (N_5486,N_4997,N_4610);
or U5487 (N_5487,N_4089,N_4953);
or U5488 (N_5488,N_4070,N_4804);
and U5489 (N_5489,N_4116,N_4509);
and U5490 (N_5490,N_4589,N_4304);
xnor U5491 (N_5491,N_4752,N_4272);
or U5492 (N_5492,N_4528,N_4369);
nand U5493 (N_5493,N_4737,N_4365);
or U5494 (N_5494,N_4898,N_4612);
nor U5495 (N_5495,N_4327,N_4999);
and U5496 (N_5496,N_4728,N_4255);
xor U5497 (N_5497,N_4647,N_4407);
and U5498 (N_5498,N_4453,N_4227);
xor U5499 (N_5499,N_4096,N_4540);
and U5500 (N_5500,N_4795,N_4351);
or U5501 (N_5501,N_4507,N_4895);
nand U5502 (N_5502,N_4052,N_4120);
xnor U5503 (N_5503,N_4111,N_4565);
xor U5504 (N_5504,N_4903,N_4122);
and U5505 (N_5505,N_4733,N_4905);
nand U5506 (N_5506,N_4248,N_4904);
and U5507 (N_5507,N_4502,N_4505);
or U5508 (N_5508,N_4846,N_4560);
nor U5509 (N_5509,N_4580,N_4570);
or U5510 (N_5510,N_4427,N_4553);
xnor U5511 (N_5511,N_4193,N_4945);
or U5512 (N_5512,N_4057,N_4787);
nand U5513 (N_5513,N_4000,N_4487);
and U5514 (N_5514,N_4331,N_4821);
and U5515 (N_5515,N_4216,N_4621);
xor U5516 (N_5516,N_4748,N_4670);
or U5517 (N_5517,N_4917,N_4576);
nand U5518 (N_5518,N_4146,N_4445);
and U5519 (N_5519,N_4511,N_4046);
and U5520 (N_5520,N_4001,N_4754);
or U5521 (N_5521,N_4176,N_4006);
nor U5522 (N_5522,N_4520,N_4507);
nand U5523 (N_5523,N_4021,N_4296);
nand U5524 (N_5524,N_4617,N_4740);
nand U5525 (N_5525,N_4120,N_4951);
xnor U5526 (N_5526,N_4832,N_4888);
xnor U5527 (N_5527,N_4864,N_4346);
xnor U5528 (N_5528,N_4886,N_4980);
and U5529 (N_5529,N_4339,N_4931);
nor U5530 (N_5530,N_4431,N_4067);
or U5531 (N_5531,N_4426,N_4854);
or U5532 (N_5532,N_4200,N_4542);
nand U5533 (N_5533,N_4418,N_4432);
nor U5534 (N_5534,N_4163,N_4141);
or U5535 (N_5535,N_4435,N_4856);
or U5536 (N_5536,N_4658,N_4220);
nand U5537 (N_5537,N_4560,N_4837);
or U5538 (N_5538,N_4012,N_4532);
nor U5539 (N_5539,N_4018,N_4241);
xnor U5540 (N_5540,N_4009,N_4594);
and U5541 (N_5541,N_4259,N_4748);
nand U5542 (N_5542,N_4864,N_4040);
nand U5543 (N_5543,N_4325,N_4611);
xor U5544 (N_5544,N_4453,N_4992);
nand U5545 (N_5545,N_4966,N_4882);
xor U5546 (N_5546,N_4787,N_4314);
nand U5547 (N_5547,N_4850,N_4201);
nor U5548 (N_5548,N_4551,N_4954);
or U5549 (N_5549,N_4576,N_4668);
nand U5550 (N_5550,N_4855,N_4978);
and U5551 (N_5551,N_4222,N_4829);
xnor U5552 (N_5552,N_4740,N_4085);
and U5553 (N_5553,N_4251,N_4446);
nor U5554 (N_5554,N_4022,N_4573);
xor U5555 (N_5555,N_4936,N_4687);
or U5556 (N_5556,N_4470,N_4273);
and U5557 (N_5557,N_4427,N_4770);
and U5558 (N_5558,N_4331,N_4574);
nor U5559 (N_5559,N_4725,N_4838);
nor U5560 (N_5560,N_4541,N_4650);
nor U5561 (N_5561,N_4759,N_4017);
nor U5562 (N_5562,N_4395,N_4853);
nor U5563 (N_5563,N_4459,N_4242);
nor U5564 (N_5564,N_4722,N_4473);
xnor U5565 (N_5565,N_4501,N_4907);
or U5566 (N_5566,N_4548,N_4444);
or U5567 (N_5567,N_4830,N_4013);
nand U5568 (N_5568,N_4820,N_4587);
xor U5569 (N_5569,N_4831,N_4813);
nor U5570 (N_5570,N_4739,N_4899);
xor U5571 (N_5571,N_4795,N_4763);
nand U5572 (N_5572,N_4576,N_4915);
and U5573 (N_5573,N_4156,N_4072);
and U5574 (N_5574,N_4516,N_4298);
nor U5575 (N_5575,N_4259,N_4564);
or U5576 (N_5576,N_4426,N_4950);
nand U5577 (N_5577,N_4185,N_4578);
nor U5578 (N_5578,N_4804,N_4702);
nand U5579 (N_5579,N_4251,N_4147);
and U5580 (N_5580,N_4066,N_4600);
nor U5581 (N_5581,N_4019,N_4295);
xor U5582 (N_5582,N_4630,N_4594);
nand U5583 (N_5583,N_4652,N_4971);
and U5584 (N_5584,N_4506,N_4571);
and U5585 (N_5585,N_4756,N_4642);
nand U5586 (N_5586,N_4689,N_4057);
or U5587 (N_5587,N_4840,N_4517);
or U5588 (N_5588,N_4701,N_4423);
or U5589 (N_5589,N_4015,N_4166);
or U5590 (N_5590,N_4489,N_4719);
nor U5591 (N_5591,N_4551,N_4298);
or U5592 (N_5592,N_4142,N_4319);
nor U5593 (N_5593,N_4466,N_4720);
and U5594 (N_5594,N_4701,N_4152);
and U5595 (N_5595,N_4873,N_4257);
nor U5596 (N_5596,N_4628,N_4976);
or U5597 (N_5597,N_4115,N_4455);
xor U5598 (N_5598,N_4359,N_4053);
xor U5599 (N_5599,N_4305,N_4519);
xor U5600 (N_5600,N_4246,N_4313);
nor U5601 (N_5601,N_4455,N_4419);
xnor U5602 (N_5602,N_4322,N_4386);
or U5603 (N_5603,N_4331,N_4190);
nor U5604 (N_5604,N_4398,N_4204);
and U5605 (N_5605,N_4876,N_4297);
nor U5606 (N_5606,N_4716,N_4598);
nand U5607 (N_5607,N_4638,N_4209);
and U5608 (N_5608,N_4525,N_4571);
nor U5609 (N_5609,N_4235,N_4489);
and U5610 (N_5610,N_4920,N_4383);
nand U5611 (N_5611,N_4232,N_4467);
xor U5612 (N_5612,N_4597,N_4683);
nor U5613 (N_5613,N_4497,N_4353);
nand U5614 (N_5614,N_4546,N_4429);
xnor U5615 (N_5615,N_4892,N_4969);
or U5616 (N_5616,N_4768,N_4647);
and U5617 (N_5617,N_4733,N_4939);
nand U5618 (N_5618,N_4467,N_4377);
xor U5619 (N_5619,N_4765,N_4920);
nor U5620 (N_5620,N_4194,N_4318);
and U5621 (N_5621,N_4646,N_4423);
nand U5622 (N_5622,N_4948,N_4021);
or U5623 (N_5623,N_4828,N_4705);
nand U5624 (N_5624,N_4225,N_4091);
and U5625 (N_5625,N_4152,N_4690);
nand U5626 (N_5626,N_4871,N_4947);
or U5627 (N_5627,N_4902,N_4713);
nand U5628 (N_5628,N_4061,N_4505);
xnor U5629 (N_5629,N_4852,N_4070);
xor U5630 (N_5630,N_4794,N_4739);
and U5631 (N_5631,N_4056,N_4164);
nor U5632 (N_5632,N_4066,N_4130);
xor U5633 (N_5633,N_4916,N_4034);
and U5634 (N_5634,N_4373,N_4297);
and U5635 (N_5635,N_4048,N_4069);
and U5636 (N_5636,N_4106,N_4608);
xnor U5637 (N_5637,N_4764,N_4101);
xor U5638 (N_5638,N_4999,N_4453);
or U5639 (N_5639,N_4837,N_4240);
xnor U5640 (N_5640,N_4990,N_4695);
nor U5641 (N_5641,N_4638,N_4823);
or U5642 (N_5642,N_4019,N_4598);
nand U5643 (N_5643,N_4139,N_4574);
nand U5644 (N_5644,N_4345,N_4472);
nand U5645 (N_5645,N_4647,N_4815);
or U5646 (N_5646,N_4060,N_4955);
or U5647 (N_5647,N_4040,N_4462);
nand U5648 (N_5648,N_4132,N_4469);
and U5649 (N_5649,N_4375,N_4682);
nand U5650 (N_5650,N_4752,N_4709);
xnor U5651 (N_5651,N_4102,N_4851);
xor U5652 (N_5652,N_4140,N_4352);
or U5653 (N_5653,N_4945,N_4773);
nor U5654 (N_5654,N_4038,N_4227);
and U5655 (N_5655,N_4399,N_4932);
nor U5656 (N_5656,N_4184,N_4089);
or U5657 (N_5657,N_4506,N_4127);
nand U5658 (N_5658,N_4505,N_4661);
nor U5659 (N_5659,N_4150,N_4120);
or U5660 (N_5660,N_4433,N_4008);
and U5661 (N_5661,N_4250,N_4162);
nand U5662 (N_5662,N_4883,N_4167);
or U5663 (N_5663,N_4184,N_4536);
and U5664 (N_5664,N_4612,N_4213);
xor U5665 (N_5665,N_4398,N_4899);
xnor U5666 (N_5666,N_4692,N_4083);
and U5667 (N_5667,N_4974,N_4025);
nand U5668 (N_5668,N_4941,N_4325);
nand U5669 (N_5669,N_4786,N_4658);
xor U5670 (N_5670,N_4098,N_4214);
xor U5671 (N_5671,N_4768,N_4676);
nor U5672 (N_5672,N_4693,N_4752);
and U5673 (N_5673,N_4898,N_4157);
or U5674 (N_5674,N_4702,N_4077);
xnor U5675 (N_5675,N_4187,N_4695);
and U5676 (N_5676,N_4491,N_4102);
or U5677 (N_5677,N_4594,N_4998);
xor U5678 (N_5678,N_4162,N_4154);
nand U5679 (N_5679,N_4943,N_4282);
nor U5680 (N_5680,N_4254,N_4237);
nor U5681 (N_5681,N_4585,N_4040);
xor U5682 (N_5682,N_4168,N_4110);
and U5683 (N_5683,N_4265,N_4910);
nor U5684 (N_5684,N_4198,N_4867);
xor U5685 (N_5685,N_4962,N_4363);
nor U5686 (N_5686,N_4328,N_4010);
xor U5687 (N_5687,N_4713,N_4740);
nand U5688 (N_5688,N_4056,N_4669);
and U5689 (N_5689,N_4236,N_4471);
or U5690 (N_5690,N_4947,N_4963);
and U5691 (N_5691,N_4960,N_4274);
or U5692 (N_5692,N_4171,N_4995);
xor U5693 (N_5693,N_4962,N_4242);
nor U5694 (N_5694,N_4728,N_4858);
and U5695 (N_5695,N_4655,N_4670);
xor U5696 (N_5696,N_4962,N_4818);
nor U5697 (N_5697,N_4975,N_4894);
xor U5698 (N_5698,N_4130,N_4991);
and U5699 (N_5699,N_4028,N_4497);
or U5700 (N_5700,N_4066,N_4552);
nand U5701 (N_5701,N_4572,N_4876);
and U5702 (N_5702,N_4792,N_4317);
nor U5703 (N_5703,N_4206,N_4656);
and U5704 (N_5704,N_4790,N_4922);
or U5705 (N_5705,N_4931,N_4123);
and U5706 (N_5706,N_4666,N_4405);
nand U5707 (N_5707,N_4012,N_4769);
nand U5708 (N_5708,N_4733,N_4350);
and U5709 (N_5709,N_4897,N_4148);
xnor U5710 (N_5710,N_4591,N_4358);
nand U5711 (N_5711,N_4851,N_4878);
nand U5712 (N_5712,N_4847,N_4088);
or U5713 (N_5713,N_4320,N_4397);
nand U5714 (N_5714,N_4118,N_4659);
nor U5715 (N_5715,N_4540,N_4672);
nor U5716 (N_5716,N_4168,N_4270);
nand U5717 (N_5717,N_4229,N_4613);
nand U5718 (N_5718,N_4418,N_4413);
and U5719 (N_5719,N_4469,N_4375);
xnor U5720 (N_5720,N_4591,N_4899);
nand U5721 (N_5721,N_4111,N_4882);
nand U5722 (N_5722,N_4949,N_4512);
xnor U5723 (N_5723,N_4957,N_4613);
nand U5724 (N_5724,N_4587,N_4505);
or U5725 (N_5725,N_4070,N_4215);
and U5726 (N_5726,N_4495,N_4900);
and U5727 (N_5727,N_4357,N_4122);
and U5728 (N_5728,N_4417,N_4810);
xor U5729 (N_5729,N_4743,N_4539);
or U5730 (N_5730,N_4778,N_4664);
and U5731 (N_5731,N_4415,N_4597);
and U5732 (N_5732,N_4119,N_4772);
and U5733 (N_5733,N_4195,N_4658);
nor U5734 (N_5734,N_4468,N_4212);
and U5735 (N_5735,N_4407,N_4929);
nand U5736 (N_5736,N_4669,N_4452);
nand U5737 (N_5737,N_4862,N_4664);
and U5738 (N_5738,N_4652,N_4770);
nor U5739 (N_5739,N_4449,N_4586);
and U5740 (N_5740,N_4280,N_4461);
nand U5741 (N_5741,N_4856,N_4640);
or U5742 (N_5742,N_4587,N_4932);
xnor U5743 (N_5743,N_4658,N_4838);
or U5744 (N_5744,N_4338,N_4021);
nor U5745 (N_5745,N_4838,N_4917);
or U5746 (N_5746,N_4798,N_4183);
and U5747 (N_5747,N_4803,N_4446);
nand U5748 (N_5748,N_4363,N_4711);
nor U5749 (N_5749,N_4016,N_4632);
or U5750 (N_5750,N_4345,N_4246);
and U5751 (N_5751,N_4534,N_4683);
and U5752 (N_5752,N_4478,N_4896);
nand U5753 (N_5753,N_4163,N_4517);
and U5754 (N_5754,N_4218,N_4008);
or U5755 (N_5755,N_4057,N_4624);
or U5756 (N_5756,N_4399,N_4289);
or U5757 (N_5757,N_4394,N_4808);
nor U5758 (N_5758,N_4167,N_4569);
or U5759 (N_5759,N_4903,N_4039);
nand U5760 (N_5760,N_4504,N_4237);
nand U5761 (N_5761,N_4134,N_4946);
xnor U5762 (N_5762,N_4118,N_4619);
xnor U5763 (N_5763,N_4011,N_4283);
or U5764 (N_5764,N_4227,N_4268);
xor U5765 (N_5765,N_4138,N_4775);
nand U5766 (N_5766,N_4931,N_4119);
nor U5767 (N_5767,N_4176,N_4633);
xnor U5768 (N_5768,N_4024,N_4163);
nand U5769 (N_5769,N_4271,N_4136);
nor U5770 (N_5770,N_4510,N_4901);
and U5771 (N_5771,N_4185,N_4060);
nand U5772 (N_5772,N_4809,N_4107);
nor U5773 (N_5773,N_4888,N_4953);
and U5774 (N_5774,N_4679,N_4587);
and U5775 (N_5775,N_4408,N_4669);
xor U5776 (N_5776,N_4931,N_4978);
or U5777 (N_5777,N_4924,N_4337);
xnor U5778 (N_5778,N_4438,N_4393);
nand U5779 (N_5779,N_4995,N_4669);
or U5780 (N_5780,N_4371,N_4067);
nor U5781 (N_5781,N_4801,N_4023);
nor U5782 (N_5782,N_4394,N_4666);
and U5783 (N_5783,N_4217,N_4007);
nand U5784 (N_5784,N_4642,N_4532);
xor U5785 (N_5785,N_4106,N_4843);
xor U5786 (N_5786,N_4196,N_4864);
and U5787 (N_5787,N_4354,N_4837);
nand U5788 (N_5788,N_4955,N_4128);
nand U5789 (N_5789,N_4752,N_4178);
or U5790 (N_5790,N_4983,N_4810);
nand U5791 (N_5791,N_4324,N_4595);
nand U5792 (N_5792,N_4006,N_4036);
nand U5793 (N_5793,N_4405,N_4241);
xor U5794 (N_5794,N_4379,N_4984);
or U5795 (N_5795,N_4363,N_4712);
xnor U5796 (N_5796,N_4847,N_4369);
xor U5797 (N_5797,N_4419,N_4427);
nand U5798 (N_5798,N_4921,N_4205);
and U5799 (N_5799,N_4196,N_4872);
and U5800 (N_5800,N_4712,N_4690);
xnor U5801 (N_5801,N_4920,N_4880);
xor U5802 (N_5802,N_4269,N_4740);
nor U5803 (N_5803,N_4869,N_4824);
nor U5804 (N_5804,N_4463,N_4922);
or U5805 (N_5805,N_4545,N_4789);
nor U5806 (N_5806,N_4175,N_4950);
xnor U5807 (N_5807,N_4343,N_4651);
or U5808 (N_5808,N_4895,N_4961);
and U5809 (N_5809,N_4734,N_4219);
xor U5810 (N_5810,N_4739,N_4910);
nand U5811 (N_5811,N_4457,N_4045);
and U5812 (N_5812,N_4745,N_4310);
nor U5813 (N_5813,N_4904,N_4127);
and U5814 (N_5814,N_4578,N_4971);
nor U5815 (N_5815,N_4722,N_4513);
xnor U5816 (N_5816,N_4328,N_4929);
xor U5817 (N_5817,N_4575,N_4676);
xnor U5818 (N_5818,N_4955,N_4349);
nor U5819 (N_5819,N_4814,N_4097);
and U5820 (N_5820,N_4715,N_4292);
nor U5821 (N_5821,N_4836,N_4451);
nor U5822 (N_5822,N_4098,N_4501);
and U5823 (N_5823,N_4080,N_4075);
and U5824 (N_5824,N_4818,N_4751);
or U5825 (N_5825,N_4895,N_4584);
xor U5826 (N_5826,N_4703,N_4973);
xnor U5827 (N_5827,N_4565,N_4332);
nand U5828 (N_5828,N_4475,N_4304);
and U5829 (N_5829,N_4315,N_4729);
nand U5830 (N_5830,N_4660,N_4014);
nor U5831 (N_5831,N_4511,N_4548);
xor U5832 (N_5832,N_4939,N_4532);
or U5833 (N_5833,N_4782,N_4978);
nor U5834 (N_5834,N_4866,N_4551);
nor U5835 (N_5835,N_4215,N_4479);
and U5836 (N_5836,N_4921,N_4484);
and U5837 (N_5837,N_4741,N_4795);
and U5838 (N_5838,N_4651,N_4291);
xor U5839 (N_5839,N_4044,N_4815);
xor U5840 (N_5840,N_4983,N_4126);
and U5841 (N_5841,N_4248,N_4995);
nor U5842 (N_5842,N_4606,N_4547);
nor U5843 (N_5843,N_4258,N_4896);
and U5844 (N_5844,N_4785,N_4973);
nand U5845 (N_5845,N_4463,N_4039);
or U5846 (N_5846,N_4248,N_4959);
nand U5847 (N_5847,N_4355,N_4963);
nand U5848 (N_5848,N_4756,N_4790);
nand U5849 (N_5849,N_4568,N_4744);
nor U5850 (N_5850,N_4818,N_4347);
nor U5851 (N_5851,N_4196,N_4335);
nand U5852 (N_5852,N_4675,N_4531);
and U5853 (N_5853,N_4475,N_4656);
nand U5854 (N_5854,N_4888,N_4862);
nand U5855 (N_5855,N_4791,N_4902);
nand U5856 (N_5856,N_4429,N_4843);
and U5857 (N_5857,N_4791,N_4255);
or U5858 (N_5858,N_4820,N_4992);
and U5859 (N_5859,N_4164,N_4688);
nor U5860 (N_5860,N_4744,N_4931);
or U5861 (N_5861,N_4393,N_4358);
and U5862 (N_5862,N_4279,N_4793);
and U5863 (N_5863,N_4968,N_4792);
xnor U5864 (N_5864,N_4082,N_4904);
nor U5865 (N_5865,N_4778,N_4793);
and U5866 (N_5866,N_4794,N_4829);
nor U5867 (N_5867,N_4727,N_4724);
or U5868 (N_5868,N_4210,N_4977);
or U5869 (N_5869,N_4419,N_4019);
nand U5870 (N_5870,N_4173,N_4568);
nand U5871 (N_5871,N_4676,N_4491);
nand U5872 (N_5872,N_4190,N_4633);
or U5873 (N_5873,N_4119,N_4139);
or U5874 (N_5874,N_4212,N_4785);
nand U5875 (N_5875,N_4651,N_4218);
or U5876 (N_5876,N_4222,N_4217);
nor U5877 (N_5877,N_4978,N_4079);
nand U5878 (N_5878,N_4329,N_4800);
nand U5879 (N_5879,N_4889,N_4671);
and U5880 (N_5880,N_4523,N_4606);
nor U5881 (N_5881,N_4461,N_4488);
nor U5882 (N_5882,N_4657,N_4427);
nand U5883 (N_5883,N_4369,N_4350);
nand U5884 (N_5884,N_4468,N_4898);
xor U5885 (N_5885,N_4212,N_4766);
or U5886 (N_5886,N_4720,N_4307);
nand U5887 (N_5887,N_4834,N_4233);
or U5888 (N_5888,N_4701,N_4779);
xor U5889 (N_5889,N_4789,N_4538);
nor U5890 (N_5890,N_4415,N_4892);
and U5891 (N_5891,N_4791,N_4569);
nor U5892 (N_5892,N_4323,N_4174);
and U5893 (N_5893,N_4944,N_4491);
nand U5894 (N_5894,N_4609,N_4721);
nand U5895 (N_5895,N_4578,N_4473);
nand U5896 (N_5896,N_4420,N_4385);
nand U5897 (N_5897,N_4555,N_4995);
nor U5898 (N_5898,N_4367,N_4596);
nand U5899 (N_5899,N_4879,N_4118);
nor U5900 (N_5900,N_4012,N_4063);
or U5901 (N_5901,N_4094,N_4602);
nand U5902 (N_5902,N_4625,N_4901);
xor U5903 (N_5903,N_4898,N_4387);
nand U5904 (N_5904,N_4012,N_4267);
and U5905 (N_5905,N_4249,N_4715);
nand U5906 (N_5906,N_4726,N_4081);
nor U5907 (N_5907,N_4791,N_4774);
xnor U5908 (N_5908,N_4029,N_4785);
nor U5909 (N_5909,N_4068,N_4799);
and U5910 (N_5910,N_4639,N_4434);
nand U5911 (N_5911,N_4647,N_4323);
nor U5912 (N_5912,N_4777,N_4823);
nor U5913 (N_5913,N_4665,N_4655);
and U5914 (N_5914,N_4634,N_4432);
nor U5915 (N_5915,N_4298,N_4033);
and U5916 (N_5916,N_4076,N_4604);
and U5917 (N_5917,N_4178,N_4554);
nor U5918 (N_5918,N_4420,N_4049);
or U5919 (N_5919,N_4852,N_4935);
xnor U5920 (N_5920,N_4025,N_4791);
xor U5921 (N_5921,N_4788,N_4823);
or U5922 (N_5922,N_4640,N_4645);
and U5923 (N_5923,N_4811,N_4497);
and U5924 (N_5924,N_4264,N_4860);
nor U5925 (N_5925,N_4689,N_4390);
or U5926 (N_5926,N_4387,N_4623);
xnor U5927 (N_5927,N_4148,N_4549);
and U5928 (N_5928,N_4608,N_4576);
xnor U5929 (N_5929,N_4112,N_4796);
xor U5930 (N_5930,N_4590,N_4618);
or U5931 (N_5931,N_4618,N_4338);
or U5932 (N_5932,N_4904,N_4889);
nor U5933 (N_5933,N_4223,N_4165);
nor U5934 (N_5934,N_4689,N_4821);
and U5935 (N_5935,N_4607,N_4628);
and U5936 (N_5936,N_4135,N_4477);
xnor U5937 (N_5937,N_4293,N_4833);
nor U5938 (N_5938,N_4407,N_4565);
or U5939 (N_5939,N_4618,N_4764);
nand U5940 (N_5940,N_4111,N_4694);
nand U5941 (N_5941,N_4049,N_4029);
nand U5942 (N_5942,N_4660,N_4314);
xnor U5943 (N_5943,N_4096,N_4651);
or U5944 (N_5944,N_4955,N_4305);
nor U5945 (N_5945,N_4584,N_4734);
nand U5946 (N_5946,N_4386,N_4425);
and U5947 (N_5947,N_4155,N_4366);
or U5948 (N_5948,N_4003,N_4247);
nand U5949 (N_5949,N_4423,N_4974);
nor U5950 (N_5950,N_4681,N_4430);
nor U5951 (N_5951,N_4857,N_4304);
and U5952 (N_5952,N_4890,N_4807);
nor U5953 (N_5953,N_4976,N_4553);
and U5954 (N_5954,N_4812,N_4743);
or U5955 (N_5955,N_4612,N_4089);
xnor U5956 (N_5956,N_4637,N_4190);
xor U5957 (N_5957,N_4420,N_4433);
nor U5958 (N_5958,N_4987,N_4102);
xor U5959 (N_5959,N_4932,N_4699);
and U5960 (N_5960,N_4029,N_4204);
nand U5961 (N_5961,N_4156,N_4365);
and U5962 (N_5962,N_4542,N_4531);
or U5963 (N_5963,N_4372,N_4790);
xor U5964 (N_5964,N_4825,N_4244);
nand U5965 (N_5965,N_4158,N_4624);
and U5966 (N_5966,N_4452,N_4542);
nand U5967 (N_5967,N_4150,N_4237);
and U5968 (N_5968,N_4298,N_4023);
and U5969 (N_5969,N_4145,N_4055);
xnor U5970 (N_5970,N_4806,N_4355);
or U5971 (N_5971,N_4068,N_4865);
xor U5972 (N_5972,N_4530,N_4455);
nor U5973 (N_5973,N_4491,N_4306);
and U5974 (N_5974,N_4073,N_4491);
nor U5975 (N_5975,N_4388,N_4408);
nand U5976 (N_5976,N_4086,N_4507);
and U5977 (N_5977,N_4410,N_4003);
or U5978 (N_5978,N_4495,N_4295);
nor U5979 (N_5979,N_4734,N_4453);
and U5980 (N_5980,N_4512,N_4574);
nor U5981 (N_5981,N_4367,N_4853);
nor U5982 (N_5982,N_4177,N_4601);
nor U5983 (N_5983,N_4451,N_4876);
nand U5984 (N_5984,N_4264,N_4826);
nor U5985 (N_5985,N_4892,N_4435);
xor U5986 (N_5986,N_4893,N_4947);
xor U5987 (N_5987,N_4486,N_4987);
xnor U5988 (N_5988,N_4900,N_4153);
or U5989 (N_5989,N_4487,N_4371);
nand U5990 (N_5990,N_4610,N_4225);
or U5991 (N_5991,N_4028,N_4356);
or U5992 (N_5992,N_4294,N_4286);
nand U5993 (N_5993,N_4701,N_4467);
and U5994 (N_5994,N_4591,N_4723);
xnor U5995 (N_5995,N_4641,N_4412);
or U5996 (N_5996,N_4325,N_4375);
or U5997 (N_5997,N_4277,N_4405);
and U5998 (N_5998,N_4582,N_4785);
xor U5999 (N_5999,N_4671,N_4213);
or U6000 (N_6000,N_5468,N_5479);
xnor U6001 (N_6001,N_5129,N_5414);
or U6002 (N_6002,N_5385,N_5121);
nand U6003 (N_6003,N_5357,N_5484);
or U6004 (N_6004,N_5411,N_5311);
or U6005 (N_6005,N_5421,N_5260);
xnor U6006 (N_6006,N_5042,N_5596);
nand U6007 (N_6007,N_5926,N_5838);
xor U6008 (N_6008,N_5512,N_5244);
and U6009 (N_6009,N_5112,N_5934);
nand U6010 (N_6010,N_5697,N_5417);
nand U6011 (N_6011,N_5921,N_5541);
or U6012 (N_6012,N_5241,N_5028);
xnor U6013 (N_6013,N_5320,N_5097);
and U6014 (N_6014,N_5654,N_5950);
xnor U6015 (N_6015,N_5165,N_5398);
nand U6016 (N_6016,N_5291,N_5927);
xor U6017 (N_6017,N_5547,N_5844);
and U6018 (N_6018,N_5239,N_5614);
or U6019 (N_6019,N_5147,N_5712);
xor U6020 (N_6020,N_5806,N_5497);
or U6021 (N_6021,N_5024,N_5508);
xor U6022 (N_6022,N_5161,N_5397);
xor U6023 (N_6023,N_5723,N_5388);
and U6024 (N_6024,N_5317,N_5036);
or U6025 (N_6025,N_5841,N_5336);
and U6026 (N_6026,N_5308,N_5115);
nor U6027 (N_6027,N_5245,N_5300);
nand U6028 (N_6028,N_5586,N_5879);
or U6029 (N_6029,N_5450,N_5002);
and U6030 (N_6030,N_5142,N_5815);
and U6031 (N_6031,N_5400,N_5642);
nor U6032 (N_6032,N_5882,N_5946);
or U6033 (N_6033,N_5328,N_5187);
nand U6034 (N_6034,N_5622,N_5383);
and U6035 (N_6035,N_5919,N_5659);
and U6036 (N_6036,N_5086,N_5158);
nand U6037 (N_6037,N_5418,N_5343);
nor U6038 (N_6038,N_5782,N_5326);
and U6039 (N_6039,N_5648,N_5183);
xnor U6040 (N_6040,N_5575,N_5790);
xor U6041 (N_6041,N_5848,N_5119);
nor U6042 (N_6042,N_5854,N_5764);
xnor U6043 (N_6043,N_5874,N_5981);
and U6044 (N_6044,N_5406,N_5208);
nand U6045 (N_6045,N_5840,N_5638);
xnor U6046 (N_6046,N_5608,N_5469);
xnor U6047 (N_6047,N_5702,N_5964);
xnor U6048 (N_6048,N_5817,N_5914);
nor U6049 (N_6049,N_5903,N_5756);
nor U6050 (N_6050,N_5196,N_5281);
nor U6051 (N_6051,N_5490,N_5857);
or U6052 (N_6052,N_5886,N_5564);
or U6053 (N_6053,N_5200,N_5538);
and U6054 (N_6054,N_5639,N_5683);
nand U6055 (N_6055,N_5849,N_5319);
nand U6056 (N_6056,N_5017,N_5082);
nand U6057 (N_6057,N_5068,N_5894);
nand U6058 (N_6058,N_5685,N_5120);
xnor U6059 (N_6059,N_5229,N_5922);
and U6060 (N_6060,N_5724,N_5796);
or U6061 (N_6061,N_5627,N_5652);
xnor U6062 (N_6062,N_5014,N_5525);
or U6063 (N_6063,N_5907,N_5667);
and U6064 (N_6064,N_5714,N_5626);
or U6065 (N_6065,N_5333,N_5118);
xnor U6066 (N_6066,N_5709,N_5759);
nor U6067 (N_6067,N_5440,N_5318);
xnor U6068 (N_6068,N_5783,N_5352);
and U6069 (N_6069,N_5855,N_5455);
xor U6070 (N_6070,N_5337,N_5277);
or U6071 (N_6071,N_5456,N_5993);
xor U6072 (N_6072,N_5961,N_5008);
nand U6073 (N_6073,N_5185,N_5100);
xnor U6074 (N_6074,N_5307,N_5314);
or U6075 (N_6075,N_5134,N_5792);
and U6076 (N_6076,N_5269,N_5688);
xnor U6077 (N_6077,N_5928,N_5303);
or U6078 (N_6078,N_5209,N_5049);
and U6079 (N_6079,N_5252,N_5482);
xor U6080 (N_6080,N_5433,N_5199);
nand U6081 (N_6081,N_5203,N_5560);
or U6082 (N_6082,N_5077,N_5368);
nor U6083 (N_6083,N_5713,N_5064);
or U6084 (N_6084,N_5016,N_5684);
nand U6085 (N_6085,N_5289,N_5734);
xor U6086 (N_6086,N_5628,N_5675);
nand U6087 (N_6087,N_5248,N_5195);
xor U6088 (N_6088,N_5325,N_5087);
or U6089 (N_6089,N_5565,N_5828);
nor U6090 (N_6090,N_5572,N_5571);
xnor U6091 (N_6091,N_5872,N_5415);
nor U6092 (N_6092,N_5348,N_5364);
xnor U6093 (N_6093,N_5693,N_5194);
or U6094 (N_6094,N_5753,N_5130);
nand U6095 (N_6095,N_5917,N_5589);
nor U6096 (N_6096,N_5265,N_5021);
and U6097 (N_6097,N_5833,N_5672);
and U6098 (N_6098,N_5069,N_5096);
nor U6099 (N_6099,N_5682,N_5650);
xnor U6100 (N_6100,N_5278,N_5284);
xnor U6101 (N_6101,N_5338,N_5076);
and U6102 (N_6102,N_5228,N_5808);
nand U6103 (N_6103,N_5148,N_5020);
nor U6104 (N_6104,N_5137,N_5197);
and U6105 (N_6105,N_5056,N_5553);
xor U6106 (N_6106,N_5823,N_5827);
nand U6107 (N_6107,N_5593,N_5190);
or U6108 (N_6108,N_5274,N_5795);
and U6109 (N_6109,N_5633,N_5821);
nand U6110 (N_6110,N_5491,N_5146);
nand U6111 (N_6111,N_5132,N_5671);
nor U6112 (N_6112,N_5880,N_5568);
nor U6113 (N_6113,N_5610,N_5286);
nor U6114 (N_6114,N_5972,N_5396);
nand U6115 (N_6115,N_5094,N_5166);
nand U6116 (N_6116,N_5381,N_5316);
nand U6117 (N_6117,N_5550,N_5775);
or U6118 (N_6118,N_5210,N_5900);
nand U6119 (N_6119,N_5302,N_5151);
nor U6120 (N_6120,N_5859,N_5150);
xor U6121 (N_6121,N_5973,N_5298);
or U6122 (N_6122,N_5407,N_5009);
xor U6123 (N_6123,N_5125,N_5389);
or U6124 (N_6124,N_5902,N_5606);
or U6125 (N_6125,N_5947,N_5634);
or U6126 (N_6126,N_5910,N_5409);
and U6127 (N_6127,N_5053,N_5279);
nand U6128 (N_6128,N_5386,N_5613);
or U6129 (N_6129,N_5694,N_5242);
nand U6130 (N_6130,N_5135,N_5149);
and U6131 (N_6131,N_5812,N_5976);
and U6132 (N_6132,N_5974,N_5435);
nand U6133 (N_6133,N_5991,N_5478);
nand U6134 (N_6134,N_5915,N_5530);
or U6135 (N_6135,N_5104,N_5537);
and U6136 (N_6136,N_5567,N_5350);
and U6137 (N_6137,N_5520,N_5816);
or U6138 (N_6138,N_5349,N_5853);
nor U6139 (N_6139,N_5445,N_5085);
nor U6140 (N_6140,N_5052,N_5519);
xor U6141 (N_6141,N_5123,N_5984);
xnor U6142 (N_6142,N_5515,N_5788);
nand U6143 (N_6143,N_5144,N_5138);
xor U6144 (N_6144,N_5594,N_5888);
and U6145 (N_6145,N_5360,N_5198);
and U6146 (N_6146,N_5040,N_5152);
nor U6147 (N_6147,N_5646,N_5356);
xor U6148 (N_6148,N_5920,N_5892);
or U6149 (N_6149,N_5354,N_5977);
nor U6150 (N_6150,N_5653,N_5958);
nor U6151 (N_6151,N_5620,N_5377);
nor U6152 (N_6152,N_5374,N_5404);
nor U6153 (N_6153,N_5342,N_5699);
xor U6154 (N_6154,N_5544,N_5952);
nor U6155 (N_6155,N_5539,N_5665);
xor U6156 (N_6156,N_5770,N_5091);
nor U6157 (N_6157,N_5391,N_5117);
or U6158 (N_6158,N_5563,N_5233);
xor U6159 (N_6159,N_5465,N_5163);
xor U6160 (N_6160,N_5630,N_5366);
and U6161 (N_6161,N_5640,N_5532);
and U6162 (N_6162,N_5836,N_5031);
nand U6163 (N_6163,N_5708,N_5645);
and U6164 (N_6164,N_5700,N_5358);
nand U6165 (N_6165,N_5800,N_5707);
nor U6166 (N_6166,N_5932,N_5073);
nor U6167 (N_6167,N_5136,N_5705);
nor U6168 (N_6168,N_5944,N_5765);
nor U6169 (N_6169,N_5215,N_5583);
and U6170 (N_6170,N_5636,N_5032);
and U6171 (N_6171,N_5526,N_5425);
or U6172 (N_6172,N_5592,N_5171);
nand U6173 (N_6173,N_5851,N_5698);
and U6174 (N_6174,N_5581,N_5732);
and U6175 (N_6175,N_5579,N_5048);
or U6176 (N_6176,N_5089,N_5726);
and U6177 (N_6177,N_5884,N_5290);
or U6178 (N_6178,N_5037,N_5677);
nand U6179 (N_6179,N_5191,N_5295);
nand U6180 (N_6180,N_5483,N_5457);
nor U6181 (N_6181,N_5585,N_5427);
and U6182 (N_6182,N_5113,N_5804);
nor U6183 (N_6183,N_5426,N_5704);
and U6184 (N_6184,N_5387,N_5246);
xnor U6185 (N_6185,N_5935,N_5780);
or U6186 (N_6186,N_5625,N_5438);
nor U6187 (N_6187,N_5255,N_5359);
nand U6188 (N_6188,N_5680,N_5858);
or U6189 (N_6189,N_5876,N_5503);
nand U6190 (N_6190,N_5691,N_5270);
and U6191 (N_6191,N_5754,N_5598);
xor U6192 (N_6192,N_5744,N_5924);
and U6193 (N_6193,N_5329,N_5401);
and U6194 (N_6194,N_5271,N_5088);
and U6195 (N_6195,N_5825,N_5826);
nand U6196 (N_6196,N_5220,N_5225);
or U6197 (N_6197,N_5803,N_5116);
or U6198 (N_6198,N_5181,N_5495);
nor U6199 (N_6199,N_5382,N_5078);
or U6200 (N_6200,N_5390,N_5339);
and U6201 (N_6201,N_5370,N_5987);
and U6202 (N_6202,N_5331,N_5590);
or U6203 (N_6203,N_5647,N_5745);
nor U6204 (N_6204,N_5706,N_5766);
and U6205 (N_6205,N_5601,N_5023);
nor U6206 (N_6206,N_5802,N_5408);
and U6207 (N_6207,N_5644,N_5101);
xnor U6208 (N_6208,N_5066,N_5217);
nand U6209 (N_6209,N_5504,N_5030);
nand U6210 (N_6210,N_5664,N_5752);
nand U6211 (N_6211,N_5847,N_5039);
or U6212 (N_6212,N_5868,N_5529);
nor U6213 (N_6213,N_5536,N_5441);
nor U6214 (N_6214,N_5605,N_5341);
nor U6215 (N_6215,N_5953,N_5092);
or U6216 (N_6216,N_5480,N_5025);
nor U6217 (N_6217,N_5862,N_5897);
or U6218 (N_6218,N_5813,N_5127);
nor U6219 (N_6219,N_5616,N_5211);
nand U6220 (N_6220,N_5378,N_5019);
nor U6221 (N_6221,N_5501,N_5548);
nand U6222 (N_6222,N_5943,N_5965);
or U6223 (N_6223,N_5580,N_5000);
or U6224 (N_6224,N_5980,N_5988);
or U6225 (N_6225,N_5686,N_5243);
xnor U6226 (N_6226,N_5600,N_5607);
nand U6227 (N_6227,N_5617,N_5182);
nand U6228 (N_6228,N_5176,N_5798);
xnor U6229 (N_6229,N_5710,N_5930);
and U6230 (N_6230,N_5735,N_5065);
xnor U6231 (N_6231,N_5084,N_5747);
or U6232 (N_6232,N_5736,N_5670);
or U6233 (N_6233,N_5948,N_5098);
and U6234 (N_6234,N_5256,N_5340);
nor U6235 (N_6235,N_5105,N_5971);
nand U6236 (N_6236,N_5452,N_5951);
xnor U6237 (N_6237,N_5463,N_5192);
nor U6238 (N_6238,N_5431,N_5929);
or U6239 (N_6239,N_5003,N_5489);
nor U6240 (N_6240,N_5678,N_5375);
and U6241 (N_6241,N_5263,N_5824);
or U6242 (N_6242,N_5749,N_5889);
and U6243 (N_6243,N_5599,N_5878);
nor U6244 (N_6244,N_5058,N_5496);
xor U6245 (N_6245,N_5554,N_5454);
nand U6246 (N_6246,N_5822,N_5777);
or U6247 (N_6247,N_5227,N_5621);
and U6248 (N_6248,N_5561,N_5543);
nand U6249 (N_6249,N_5361,N_5448);
nand U6250 (N_6250,N_5758,N_5811);
nand U6251 (N_6251,N_5247,N_5380);
xnor U6252 (N_6252,N_5327,N_5459);
nand U6253 (N_6253,N_5254,N_5424);
or U6254 (N_6254,N_5293,N_5801);
or U6255 (N_6255,N_5034,N_5835);
or U6256 (N_6256,N_5602,N_5786);
and U6257 (N_6257,N_5905,N_5873);
and U6258 (N_6258,N_5657,N_5470);
nor U6259 (N_6259,N_5818,N_5035);
nor U6260 (N_6260,N_5999,N_5522);
xnor U6261 (N_6261,N_5038,N_5346);
nor U6262 (N_6262,N_5591,N_5997);
nor U6263 (N_6263,N_5842,N_5867);
or U6264 (N_6264,N_5901,N_5666);
nor U6265 (N_6265,N_5060,N_5212);
xnor U6266 (N_6266,N_5224,N_5584);
nor U6267 (N_6267,N_5179,N_5369);
xor U6268 (N_6268,N_5124,N_5738);
or U6269 (N_6269,N_5405,N_5969);
and U6270 (N_6270,N_5985,N_5830);
or U6271 (N_6271,N_5933,N_5942);
nor U6272 (N_6272,N_5072,N_5502);
nor U6273 (N_6273,N_5345,N_5159);
or U6274 (N_6274,N_5177,N_5067);
nor U6275 (N_6275,N_5332,N_5283);
nor U6276 (N_6276,N_5362,N_5301);
nor U6277 (N_6277,N_5423,N_5222);
xor U6278 (N_6278,N_5416,N_5057);
xnor U6279 (N_6279,N_5762,N_5157);
nand U6280 (N_6280,N_5133,N_5347);
and U6281 (N_6281,N_5748,N_5784);
and U6282 (N_6282,N_5516,N_5443);
and U6283 (N_6283,N_5379,N_5287);
nand U6284 (N_6284,N_5351,N_5511);
nor U6285 (N_6285,N_5186,N_5310);
and U6286 (N_6286,N_5540,N_5912);
nand U6287 (N_6287,N_5629,N_5029);
nand U6288 (N_6288,N_5430,N_5799);
xor U6289 (N_6289,N_5778,N_5852);
and U6290 (N_6290,N_5051,N_5750);
or U6291 (N_6291,N_5558,N_5781);
and U6292 (N_6292,N_5050,N_5022);
nor U6293 (N_6293,N_5015,N_5918);
and U6294 (N_6294,N_5110,N_5820);
xnor U6295 (N_6295,N_5725,N_5845);
nor U6296 (N_6296,N_5174,N_5292);
or U6297 (N_6297,N_5962,N_5047);
and U6298 (N_6298,N_5485,N_5280);
nand U6299 (N_6299,N_5494,N_5395);
nor U6300 (N_6300,N_5837,N_5939);
nor U6301 (N_6301,N_5432,N_5975);
xor U6302 (N_6302,N_5990,N_5413);
nor U6303 (N_6303,N_5624,N_5372);
xnor U6304 (N_6304,N_5010,N_5559);
xnor U6305 (N_6305,N_5739,N_5566);
and U6306 (N_6306,N_5582,N_5170);
nor U6307 (N_6307,N_5080,N_5760);
or U6308 (N_6308,N_5216,N_5891);
nand U6309 (N_6309,N_5956,N_5403);
nand U6310 (N_6310,N_5552,N_5861);
and U6311 (N_6311,N_5692,N_5304);
nor U6312 (N_6312,N_5899,N_5488);
nand U6313 (N_6313,N_5221,N_5164);
and U6314 (N_6314,N_5658,N_5940);
xnor U6315 (N_6315,N_5871,N_5729);
xor U6316 (N_6316,N_5986,N_5925);
nand U6317 (N_6317,N_5906,N_5661);
or U6318 (N_6318,N_5772,N_5041);
nor U6319 (N_6319,N_5510,N_5419);
xor U6320 (N_6320,N_5505,N_5557);
or U6321 (N_6321,N_5498,N_5172);
or U6322 (N_6322,N_5730,N_5787);
and U6323 (N_6323,N_5676,N_5937);
and U6324 (N_6324,N_5306,N_5365);
and U6325 (N_6325,N_5534,N_5296);
xor U6326 (N_6326,N_5487,N_5979);
nor U6327 (N_6327,N_5453,N_5954);
and U6328 (N_6328,N_5513,N_5588);
or U6329 (N_6329,N_5773,N_5393);
nor U6330 (N_6330,N_5574,N_5865);
and U6331 (N_6331,N_5743,N_5353);
or U6332 (N_6332,N_5911,N_5959);
nor U6333 (N_6333,N_5083,N_5475);
nor U6334 (N_6334,N_5230,N_5079);
and U6335 (N_6335,N_5226,N_5061);
xnor U6336 (N_6336,N_5866,N_5687);
nand U6337 (N_6337,N_5322,N_5690);
nor U6338 (N_6338,N_5517,N_5721);
nor U6339 (N_6339,N_5492,N_5982);
and U6340 (N_6340,N_5931,N_5272);
or U6341 (N_6341,N_5446,N_5305);
xnor U6342 (N_6342,N_5481,N_5612);
and U6343 (N_6343,N_5623,N_5461);
xnor U6344 (N_6344,N_5055,N_5074);
nand U6345 (N_6345,N_5632,N_5012);
or U6346 (N_6346,N_5500,N_5774);
xor U6347 (N_6347,N_5001,N_5716);
nor U6348 (N_6348,N_5436,N_5462);
xor U6349 (N_6349,N_5081,N_5656);
nand U6350 (N_6350,N_5881,N_5167);
xor U6351 (N_6351,N_5733,N_5885);
nor U6352 (N_6352,N_5207,N_5949);
xor U6353 (N_6353,N_5896,N_5063);
and U6354 (N_6354,N_5850,N_5649);
and U6355 (N_6355,N_5893,N_5238);
nor U6356 (N_6356,N_5741,N_5324);
nor U6357 (N_6357,N_5033,N_5335);
nand U6358 (N_6358,N_5219,N_5887);
and U6359 (N_6359,N_5330,N_5545);
nand U6360 (N_6360,N_5235,N_5577);
xnor U6361 (N_6361,N_5437,N_5111);
nand U6362 (N_6362,N_5751,N_5477);
or U6363 (N_6363,N_5141,N_5202);
or U6364 (N_6364,N_5237,N_5631);
nor U6365 (N_6365,N_5908,N_5275);
xor U6366 (N_6366,N_5471,N_5718);
nor U6367 (N_6367,N_5662,N_5913);
and U6368 (N_6368,N_5261,N_5312);
xnor U6369 (N_6369,N_5533,N_5737);
nand U6370 (N_6370,N_5890,N_5250);
nand U6371 (N_6371,N_5978,N_5236);
or U6372 (N_6372,N_5819,N_5916);
xor U6373 (N_6373,N_5093,N_5655);
and U6374 (N_6374,N_5587,N_5995);
xnor U6375 (N_6375,N_5904,N_5755);
or U6376 (N_6376,N_5864,N_5994);
and U6377 (N_6377,N_5509,N_5006);
xnor U6378 (N_6378,N_5785,N_5562);
nand U6379 (N_6379,N_5472,N_5779);
and U6380 (N_6380,N_5178,N_5143);
or U6381 (N_6381,N_5273,N_5367);
nor U6382 (N_6382,N_5771,N_5102);
xnor U6383 (N_6383,N_5371,N_5344);
nand U6384 (N_6384,N_5717,N_5829);
nand U6385 (N_6385,N_5728,N_5323);
and U6386 (N_6386,N_5442,N_5262);
nor U6387 (N_6387,N_5573,N_5394);
and U6388 (N_6388,N_5188,N_5422);
or U6389 (N_6389,N_5259,N_5095);
and U6390 (N_6390,N_5107,N_5938);
nand U6391 (N_6391,N_5309,N_5731);
nor U6392 (N_6392,N_5619,N_5258);
or U6393 (N_6393,N_5412,N_5114);
or U6394 (N_6394,N_5679,N_5145);
nand U6395 (N_6395,N_5355,N_5420);
nand U6396 (N_6396,N_5609,N_5576);
xnor U6397 (N_6397,N_5527,N_5551);
or U6398 (N_6398,N_5473,N_5810);
nor U6399 (N_6399,N_5027,N_5282);
and U6400 (N_6400,N_5266,N_5789);
nand U6401 (N_6401,N_5807,N_5288);
or U6402 (N_6402,N_5402,N_5809);
or U6403 (N_6403,N_5054,N_5004);
or U6404 (N_6404,N_5460,N_5856);
xnor U6405 (N_6405,N_5140,N_5797);
nand U6406 (N_6406,N_5681,N_5410);
or U6407 (N_6407,N_5696,N_5615);
nor U6408 (N_6408,N_5875,N_5523);
or U6409 (N_6409,N_5218,N_5669);
and U6410 (N_6410,N_5466,N_5249);
xnor U6411 (N_6411,N_5719,N_5205);
xnor U6412 (N_6412,N_5805,N_5767);
nor U6413 (N_6413,N_5321,N_5791);
xor U6414 (N_6414,N_5429,N_5846);
xor U6415 (N_6415,N_5231,N_5071);
nand U6416 (N_6416,N_5740,N_5555);
or U6417 (N_6417,N_5674,N_5531);
or U6418 (N_6418,N_5831,N_5264);
or U6419 (N_6419,N_5376,N_5045);
nor U6420 (N_6420,N_5970,N_5153);
xor U6421 (N_6421,N_5597,N_5162);
and U6422 (N_6422,N_5711,N_5315);
nand U6423 (N_6423,N_5556,N_5668);
or U6424 (N_6424,N_5695,N_5514);
nand U6425 (N_6425,N_5139,N_5201);
or U6426 (N_6426,N_5635,N_5595);
nor U6427 (N_6427,N_5439,N_5793);
nand U6428 (N_6428,N_5059,N_5996);
nand U6429 (N_6429,N_5834,N_5106);
nand U6430 (N_6430,N_5869,N_5128);
xor U6431 (N_6431,N_5660,N_5447);
xor U6432 (N_6432,N_5449,N_5458);
or U6433 (N_6433,N_5070,N_5746);
and U6434 (N_6434,N_5257,N_5968);
and U6435 (N_6435,N_5499,N_5232);
nor U6436 (N_6436,N_5474,N_5005);
or U6437 (N_6437,N_5184,N_5535);
and U6438 (N_6438,N_5839,N_5966);
and U6439 (N_6439,N_5941,N_5007);
xnor U6440 (N_6440,N_5651,N_5168);
and U6441 (N_6441,N_5832,N_5549);
nor U6442 (N_6442,N_5294,N_5223);
or U6443 (N_6443,N_5570,N_5641);
xor U6444 (N_6444,N_5963,N_5936);
nor U6445 (N_6445,N_5524,N_5026);
xor U6446 (N_6446,N_5276,N_5603);
nor U6447 (N_6447,N_5701,N_5428);
xnor U6448 (N_6448,N_5154,N_5486);
xnor U6449 (N_6449,N_5507,N_5108);
or U6450 (N_6450,N_5173,N_5373);
nand U6451 (N_6451,N_5763,N_5578);
xnor U6452 (N_6452,N_5967,N_5109);
nor U6453 (N_6453,N_5992,N_5313);
nand U6454 (N_6454,N_5618,N_5895);
nor U6455 (N_6455,N_5769,N_5204);
and U6456 (N_6456,N_5722,N_5189);
or U6457 (N_6457,N_5213,N_5860);
nand U6458 (N_6458,N_5528,N_5175);
nand U6459 (N_6459,N_5090,N_5234);
xnor U6460 (N_6460,N_5018,N_5267);
nand U6461 (N_6461,N_5960,N_5689);
or U6462 (N_6462,N_5444,N_5663);
nor U6463 (N_6463,N_5251,N_5521);
nor U6464 (N_6464,N_5131,N_5493);
nand U6465 (N_6465,N_5776,N_5957);
and U6466 (N_6466,N_5285,N_5011);
nand U6467 (N_6467,N_5062,N_5464);
and U6468 (N_6468,N_5768,N_5955);
xnor U6469 (N_6469,N_5268,N_5122);
and U6470 (N_6470,N_5757,N_5451);
and U6471 (N_6471,N_5898,N_5193);
xor U6472 (N_6472,N_5945,N_5794);
and U6473 (N_6473,N_5870,N_5546);
xnor U6474 (N_6474,N_5604,N_5253);
or U6475 (N_6475,N_5814,N_5044);
nor U6476 (N_6476,N_5761,N_5542);
nand U6477 (N_6477,N_5673,N_5742);
nand U6478 (N_6478,N_5384,N_5013);
or U6479 (N_6479,N_5156,N_5434);
or U6480 (N_6480,N_5983,N_5883);
nor U6481 (N_6481,N_5299,N_5877);
nand U6482 (N_6482,N_5506,N_5518);
xor U6483 (N_6483,N_5297,N_5099);
or U6484 (N_6484,N_5126,N_5180);
or U6485 (N_6485,N_5843,N_5863);
nor U6486 (N_6486,N_5569,N_5643);
nand U6487 (N_6487,N_5909,N_5989);
xor U6488 (N_6488,N_5923,N_5160);
or U6489 (N_6489,N_5727,N_5998);
xor U6490 (N_6490,N_5169,N_5467);
nor U6491 (N_6491,N_5103,N_5334);
and U6492 (N_6492,N_5075,N_5715);
nor U6493 (N_6493,N_5214,N_5392);
and U6494 (N_6494,N_5476,N_5240);
or U6495 (N_6495,N_5637,N_5155);
or U6496 (N_6496,N_5046,N_5703);
or U6497 (N_6497,N_5043,N_5399);
nand U6498 (N_6498,N_5611,N_5206);
nand U6499 (N_6499,N_5363,N_5720);
and U6500 (N_6500,N_5142,N_5706);
or U6501 (N_6501,N_5729,N_5838);
or U6502 (N_6502,N_5288,N_5438);
nor U6503 (N_6503,N_5811,N_5073);
xor U6504 (N_6504,N_5995,N_5303);
or U6505 (N_6505,N_5334,N_5008);
nand U6506 (N_6506,N_5379,N_5819);
nand U6507 (N_6507,N_5332,N_5176);
or U6508 (N_6508,N_5881,N_5285);
xor U6509 (N_6509,N_5999,N_5559);
or U6510 (N_6510,N_5847,N_5379);
or U6511 (N_6511,N_5431,N_5732);
xnor U6512 (N_6512,N_5235,N_5182);
or U6513 (N_6513,N_5956,N_5608);
nor U6514 (N_6514,N_5473,N_5030);
and U6515 (N_6515,N_5920,N_5940);
and U6516 (N_6516,N_5645,N_5017);
and U6517 (N_6517,N_5921,N_5395);
nor U6518 (N_6518,N_5350,N_5777);
xor U6519 (N_6519,N_5773,N_5315);
nand U6520 (N_6520,N_5611,N_5585);
nand U6521 (N_6521,N_5325,N_5127);
and U6522 (N_6522,N_5641,N_5119);
or U6523 (N_6523,N_5754,N_5223);
nand U6524 (N_6524,N_5667,N_5167);
nor U6525 (N_6525,N_5812,N_5164);
nand U6526 (N_6526,N_5616,N_5073);
and U6527 (N_6527,N_5925,N_5940);
and U6528 (N_6528,N_5840,N_5551);
nand U6529 (N_6529,N_5042,N_5427);
nand U6530 (N_6530,N_5742,N_5555);
and U6531 (N_6531,N_5239,N_5573);
nand U6532 (N_6532,N_5520,N_5042);
and U6533 (N_6533,N_5644,N_5860);
or U6534 (N_6534,N_5541,N_5398);
xnor U6535 (N_6535,N_5140,N_5855);
nor U6536 (N_6536,N_5711,N_5183);
nand U6537 (N_6537,N_5027,N_5894);
xor U6538 (N_6538,N_5572,N_5436);
xor U6539 (N_6539,N_5570,N_5202);
xnor U6540 (N_6540,N_5074,N_5984);
nor U6541 (N_6541,N_5448,N_5867);
nand U6542 (N_6542,N_5473,N_5707);
nand U6543 (N_6543,N_5388,N_5287);
nor U6544 (N_6544,N_5743,N_5484);
nor U6545 (N_6545,N_5982,N_5522);
nor U6546 (N_6546,N_5996,N_5921);
xnor U6547 (N_6547,N_5756,N_5059);
or U6548 (N_6548,N_5281,N_5491);
xor U6549 (N_6549,N_5284,N_5740);
nand U6550 (N_6550,N_5801,N_5045);
nor U6551 (N_6551,N_5780,N_5182);
and U6552 (N_6552,N_5965,N_5179);
nand U6553 (N_6553,N_5815,N_5243);
and U6554 (N_6554,N_5143,N_5343);
xnor U6555 (N_6555,N_5688,N_5720);
xor U6556 (N_6556,N_5119,N_5670);
nor U6557 (N_6557,N_5724,N_5280);
nand U6558 (N_6558,N_5823,N_5054);
nand U6559 (N_6559,N_5327,N_5777);
or U6560 (N_6560,N_5121,N_5905);
nand U6561 (N_6561,N_5629,N_5041);
or U6562 (N_6562,N_5620,N_5479);
nor U6563 (N_6563,N_5123,N_5200);
xor U6564 (N_6564,N_5529,N_5785);
nand U6565 (N_6565,N_5350,N_5231);
xnor U6566 (N_6566,N_5965,N_5563);
and U6567 (N_6567,N_5936,N_5264);
nand U6568 (N_6568,N_5595,N_5044);
and U6569 (N_6569,N_5940,N_5892);
xor U6570 (N_6570,N_5431,N_5886);
and U6571 (N_6571,N_5741,N_5409);
and U6572 (N_6572,N_5005,N_5481);
nor U6573 (N_6573,N_5995,N_5020);
xnor U6574 (N_6574,N_5932,N_5386);
and U6575 (N_6575,N_5677,N_5114);
xor U6576 (N_6576,N_5162,N_5842);
or U6577 (N_6577,N_5251,N_5469);
and U6578 (N_6578,N_5611,N_5468);
nor U6579 (N_6579,N_5058,N_5404);
or U6580 (N_6580,N_5411,N_5481);
xor U6581 (N_6581,N_5557,N_5691);
and U6582 (N_6582,N_5350,N_5237);
nor U6583 (N_6583,N_5685,N_5080);
and U6584 (N_6584,N_5516,N_5691);
and U6585 (N_6585,N_5826,N_5934);
or U6586 (N_6586,N_5262,N_5354);
xor U6587 (N_6587,N_5147,N_5728);
or U6588 (N_6588,N_5839,N_5974);
nand U6589 (N_6589,N_5616,N_5807);
nand U6590 (N_6590,N_5404,N_5375);
xnor U6591 (N_6591,N_5691,N_5245);
and U6592 (N_6592,N_5371,N_5551);
and U6593 (N_6593,N_5981,N_5148);
xnor U6594 (N_6594,N_5555,N_5439);
nor U6595 (N_6595,N_5795,N_5782);
or U6596 (N_6596,N_5295,N_5331);
or U6597 (N_6597,N_5047,N_5766);
nand U6598 (N_6598,N_5960,N_5734);
and U6599 (N_6599,N_5924,N_5886);
nand U6600 (N_6600,N_5914,N_5484);
or U6601 (N_6601,N_5360,N_5384);
or U6602 (N_6602,N_5497,N_5220);
xnor U6603 (N_6603,N_5654,N_5368);
and U6604 (N_6604,N_5998,N_5996);
xor U6605 (N_6605,N_5394,N_5756);
or U6606 (N_6606,N_5612,N_5726);
or U6607 (N_6607,N_5559,N_5294);
nand U6608 (N_6608,N_5979,N_5191);
and U6609 (N_6609,N_5425,N_5199);
or U6610 (N_6610,N_5082,N_5252);
and U6611 (N_6611,N_5458,N_5169);
nor U6612 (N_6612,N_5305,N_5486);
or U6613 (N_6613,N_5895,N_5637);
or U6614 (N_6614,N_5738,N_5575);
nor U6615 (N_6615,N_5846,N_5885);
or U6616 (N_6616,N_5833,N_5580);
nand U6617 (N_6617,N_5893,N_5353);
and U6618 (N_6618,N_5433,N_5196);
xor U6619 (N_6619,N_5126,N_5307);
nor U6620 (N_6620,N_5182,N_5363);
or U6621 (N_6621,N_5408,N_5057);
nand U6622 (N_6622,N_5111,N_5549);
nand U6623 (N_6623,N_5996,N_5291);
nand U6624 (N_6624,N_5456,N_5523);
nor U6625 (N_6625,N_5480,N_5742);
xor U6626 (N_6626,N_5636,N_5283);
nor U6627 (N_6627,N_5130,N_5702);
or U6628 (N_6628,N_5362,N_5302);
xor U6629 (N_6629,N_5253,N_5122);
nand U6630 (N_6630,N_5668,N_5410);
xor U6631 (N_6631,N_5877,N_5682);
nand U6632 (N_6632,N_5841,N_5113);
xor U6633 (N_6633,N_5755,N_5923);
nand U6634 (N_6634,N_5436,N_5174);
and U6635 (N_6635,N_5731,N_5591);
nor U6636 (N_6636,N_5164,N_5680);
and U6637 (N_6637,N_5514,N_5079);
or U6638 (N_6638,N_5645,N_5951);
nor U6639 (N_6639,N_5104,N_5989);
xnor U6640 (N_6640,N_5138,N_5758);
nand U6641 (N_6641,N_5610,N_5337);
nand U6642 (N_6642,N_5477,N_5981);
or U6643 (N_6643,N_5217,N_5480);
nand U6644 (N_6644,N_5107,N_5298);
and U6645 (N_6645,N_5045,N_5864);
nand U6646 (N_6646,N_5039,N_5667);
and U6647 (N_6647,N_5498,N_5000);
nand U6648 (N_6648,N_5867,N_5536);
and U6649 (N_6649,N_5876,N_5046);
nand U6650 (N_6650,N_5419,N_5288);
xnor U6651 (N_6651,N_5409,N_5495);
nand U6652 (N_6652,N_5746,N_5358);
and U6653 (N_6653,N_5963,N_5762);
and U6654 (N_6654,N_5531,N_5691);
xnor U6655 (N_6655,N_5815,N_5108);
nor U6656 (N_6656,N_5988,N_5059);
and U6657 (N_6657,N_5868,N_5928);
nor U6658 (N_6658,N_5947,N_5642);
xnor U6659 (N_6659,N_5571,N_5456);
or U6660 (N_6660,N_5555,N_5652);
xnor U6661 (N_6661,N_5983,N_5350);
nand U6662 (N_6662,N_5329,N_5984);
nand U6663 (N_6663,N_5928,N_5235);
xnor U6664 (N_6664,N_5390,N_5823);
nor U6665 (N_6665,N_5862,N_5219);
nand U6666 (N_6666,N_5509,N_5588);
nor U6667 (N_6667,N_5548,N_5247);
xnor U6668 (N_6668,N_5602,N_5882);
xor U6669 (N_6669,N_5970,N_5528);
and U6670 (N_6670,N_5202,N_5088);
xor U6671 (N_6671,N_5844,N_5134);
xnor U6672 (N_6672,N_5880,N_5134);
or U6673 (N_6673,N_5869,N_5853);
or U6674 (N_6674,N_5791,N_5079);
nand U6675 (N_6675,N_5464,N_5476);
nand U6676 (N_6676,N_5389,N_5131);
xnor U6677 (N_6677,N_5175,N_5181);
or U6678 (N_6678,N_5116,N_5300);
or U6679 (N_6679,N_5605,N_5754);
nand U6680 (N_6680,N_5895,N_5936);
and U6681 (N_6681,N_5972,N_5013);
xor U6682 (N_6682,N_5494,N_5797);
nand U6683 (N_6683,N_5101,N_5153);
or U6684 (N_6684,N_5539,N_5309);
nor U6685 (N_6685,N_5630,N_5144);
xor U6686 (N_6686,N_5478,N_5085);
and U6687 (N_6687,N_5268,N_5140);
or U6688 (N_6688,N_5577,N_5762);
or U6689 (N_6689,N_5295,N_5137);
and U6690 (N_6690,N_5286,N_5929);
or U6691 (N_6691,N_5199,N_5750);
and U6692 (N_6692,N_5659,N_5271);
nor U6693 (N_6693,N_5138,N_5290);
or U6694 (N_6694,N_5654,N_5413);
or U6695 (N_6695,N_5564,N_5508);
nand U6696 (N_6696,N_5670,N_5183);
and U6697 (N_6697,N_5443,N_5203);
xnor U6698 (N_6698,N_5251,N_5633);
or U6699 (N_6699,N_5915,N_5120);
and U6700 (N_6700,N_5698,N_5560);
nor U6701 (N_6701,N_5679,N_5250);
nor U6702 (N_6702,N_5280,N_5308);
xor U6703 (N_6703,N_5279,N_5555);
nand U6704 (N_6704,N_5403,N_5140);
nand U6705 (N_6705,N_5224,N_5373);
nor U6706 (N_6706,N_5401,N_5909);
nor U6707 (N_6707,N_5165,N_5905);
or U6708 (N_6708,N_5846,N_5216);
and U6709 (N_6709,N_5039,N_5289);
or U6710 (N_6710,N_5559,N_5408);
and U6711 (N_6711,N_5465,N_5432);
and U6712 (N_6712,N_5414,N_5723);
and U6713 (N_6713,N_5064,N_5750);
nor U6714 (N_6714,N_5861,N_5110);
nor U6715 (N_6715,N_5503,N_5022);
and U6716 (N_6716,N_5237,N_5294);
nor U6717 (N_6717,N_5518,N_5743);
nor U6718 (N_6718,N_5159,N_5804);
and U6719 (N_6719,N_5314,N_5613);
and U6720 (N_6720,N_5125,N_5331);
xnor U6721 (N_6721,N_5059,N_5228);
or U6722 (N_6722,N_5348,N_5382);
or U6723 (N_6723,N_5659,N_5049);
nor U6724 (N_6724,N_5903,N_5643);
nand U6725 (N_6725,N_5372,N_5679);
and U6726 (N_6726,N_5068,N_5587);
xnor U6727 (N_6727,N_5518,N_5245);
nor U6728 (N_6728,N_5332,N_5600);
or U6729 (N_6729,N_5465,N_5962);
nand U6730 (N_6730,N_5625,N_5998);
and U6731 (N_6731,N_5874,N_5221);
xor U6732 (N_6732,N_5121,N_5991);
nand U6733 (N_6733,N_5439,N_5784);
xnor U6734 (N_6734,N_5472,N_5378);
or U6735 (N_6735,N_5269,N_5408);
or U6736 (N_6736,N_5332,N_5836);
or U6737 (N_6737,N_5100,N_5651);
nand U6738 (N_6738,N_5889,N_5689);
xnor U6739 (N_6739,N_5161,N_5761);
xnor U6740 (N_6740,N_5270,N_5940);
or U6741 (N_6741,N_5192,N_5135);
nor U6742 (N_6742,N_5767,N_5446);
or U6743 (N_6743,N_5260,N_5037);
or U6744 (N_6744,N_5953,N_5430);
xor U6745 (N_6745,N_5288,N_5962);
xor U6746 (N_6746,N_5106,N_5005);
nor U6747 (N_6747,N_5045,N_5639);
and U6748 (N_6748,N_5771,N_5790);
nor U6749 (N_6749,N_5229,N_5446);
and U6750 (N_6750,N_5756,N_5709);
nor U6751 (N_6751,N_5724,N_5648);
nor U6752 (N_6752,N_5042,N_5798);
nand U6753 (N_6753,N_5209,N_5698);
nand U6754 (N_6754,N_5307,N_5372);
and U6755 (N_6755,N_5265,N_5437);
or U6756 (N_6756,N_5363,N_5629);
or U6757 (N_6757,N_5554,N_5994);
xor U6758 (N_6758,N_5506,N_5956);
nor U6759 (N_6759,N_5367,N_5597);
or U6760 (N_6760,N_5554,N_5809);
xor U6761 (N_6761,N_5170,N_5878);
nor U6762 (N_6762,N_5255,N_5635);
nand U6763 (N_6763,N_5655,N_5211);
nor U6764 (N_6764,N_5376,N_5086);
xnor U6765 (N_6765,N_5735,N_5097);
and U6766 (N_6766,N_5951,N_5807);
nor U6767 (N_6767,N_5264,N_5110);
or U6768 (N_6768,N_5628,N_5074);
and U6769 (N_6769,N_5817,N_5384);
nor U6770 (N_6770,N_5139,N_5956);
nand U6771 (N_6771,N_5179,N_5169);
nor U6772 (N_6772,N_5148,N_5278);
nand U6773 (N_6773,N_5896,N_5474);
nand U6774 (N_6774,N_5205,N_5219);
xnor U6775 (N_6775,N_5036,N_5156);
nand U6776 (N_6776,N_5028,N_5830);
nand U6777 (N_6777,N_5873,N_5668);
and U6778 (N_6778,N_5076,N_5494);
nand U6779 (N_6779,N_5208,N_5019);
nand U6780 (N_6780,N_5891,N_5679);
or U6781 (N_6781,N_5565,N_5745);
nor U6782 (N_6782,N_5725,N_5154);
or U6783 (N_6783,N_5538,N_5341);
xnor U6784 (N_6784,N_5229,N_5038);
nand U6785 (N_6785,N_5081,N_5777);
xnor U6786 (N_6786,N_5447,N_5616);
xnor U6787 (N_6787,N_5447,N_5827);
nor U6788 (N_6788,N_5259,N_5522);
xor U6789 (N_6789,N_5342,N_5380);
nor U6790 (N_6790,N_5795,N_5133);
or U6791 (N_6791,N_5487,N_5691);
nor U6792 (N_6792,N_5151,N_5163);
or U6793 (N_6793,N_5008,N_5945);
xnor U6794 (N_6794,N_5092,N_5988);
xnor U6795 (N_6795,N_5167,N_5209);
nand U6796 (N_6796,N_5013,N_5584);
or U6797 (N_6797,N_5054,N_5973);
and U6798 (N_6798,N_5971,N_5222);
nor U6799 (N_6799,N_5310,N_5738);
and U6800 (N_6800,N_5003,N_5578);
nand U6801 (N_6801,N_5706,N_5613);
nor U6802 (N_6802,N_5333,N_5075);
nand U6803 (N_6803,N_5301,N_5509);
xor U6804 (N_6804,N_5656,N_5730);
nand U6805 (N_6805,N_5482,N_5039);
nand U6806 (N_6806,N_5733,N_5841);
xor U6807 (N_6807,N_5388,N_5951);
nand U6808 (N_6808,N_5943,N_5296);
or U6809 (N_6809,N_5771,N_5434);
nor U6810 (N_6810,N_5754,N_5056);
nor U6811 (N_6811,N_5318,N_5177);
xor U6812 (N_6812,N_5422,N_5998);
and U6813 (N_6813,N_5128,N_5791);
nand U6814 (N_6814,N_5505,N_5078);
nand U6815 (N_6815,N_5593,N_5891);
nand U6816 (N_6816,N_5955,N_5069);
or U6817 (N_6817,N_5767,N_5178);
xor U6818 (N_6818,N_5140,N_5737);
and U6819 (N_6819,N_5569,N_5449);
xnor U6820 (N_6820,N_5286,N_5647);
nor U6821 (N_6821,N_5500,N_5696);
xor U6822 (N_6822,N_5981,N_5795);
xor U6823 (N_6823,N_5374,N_5985);
and U6824 (N_6824,N_5098,N_5155);
nand U6825 (N_6825,N_5640,N_5562);
and U6826 (N_6826,N_5191,N_5583);
nand U6827 (N_6827,N_5042,N_5019);
xor U6828 (N_6828,N_5402,N_5544);
and U6829 (N_6829,N_5793,N_5067);
xor U6830 (N_6830,N_5802,N_5777);
xnor U6831 (N_6831,N_5278,N_5744);
xnor U6832 (N_6832,N_5752,N_5159);
and U6833 (N_6833,N_5488,N_5767);
or U6834 (N_6834,N_5139,N_5815);
or U6835 (N_6835,N_5796,N_5756);
xnor U6836 (N_6836,N_5171,N_5321);
or U6837 (N_6837,N_5282,N_5061);
xnor U6838 (N_6838,N_5174,N_5798);
and U6839 (N_6839,N_5366,N_5744);
nor U6840 (N_6840,N_5849,N_5823);
nor U6841 (N_6841,N_5555,N_5586);
and U6842 (N_6842,N_5977,N_5565);
nand U6843 (N_6843,N_5594,N_5938);
nand U6844 (N_6844,N_5861,N_5663);
nand U6845 (N_6845,N_5476,N_5910);
and U6846 (N_6846,N_5431,N_5113);
xnor U6847 (N_6847,N_5961,N_5023);
and U6848 (N_6848,N_5147,N_5135);
nor U6849 (N_6849,N_5553,N_5373);
nor U6850 (N_6850,N_5740,N_5304);
or U6851 (N_6851,N_5230,N_5490);
xnor U6852 (N_6852,N_5604,N_5424);
xor U6853 (N_6853,N_5822,N_5303);
xor U6854 (N_6854,N_5733,N_5795);
nor U6855 (N_6855,N_5430,N_5796);
nand U6856 (N_6856,N_5305,N_5091);
or U6857 (N_6857,N_5153,N_5421);
and U6858 (N_6858,N_5855,N_5232);
and U6859 (N_6859,N_5990,N_5877);
nand U6860 (N_6860,N_5661,N_5060);
xnor U6861 (N_6861,N_5605,N_5575);
nand U6862 (N_6862,N_5553,N_5948);
and U6863 (N_6863,N_5985,N_5186);
and U6864 (N_6864,N_5070,N_5838);
nor U6865 (N_6865,N_5878,N_5547);
nand U6866 (N_6866,N_5607,N_5282);
and U6867 (N_6867,N_5664,N_5243);
nor U6868 (N_6868,N_5662,N_5052);
and U6869 (N_6869,N_5469,N_5730);
and U6870 (N_6870,N_5252,N_5430);
xor U6871 (N_6871,N_5600,N_5418);
nor U6872 (N_6872,N_5759,N_5851);
and U6873 (N_6873,N_5174,N_5122);
nand U6874 (N_6874,N_5469,N_5238);
nor U6875 (N_6875,N_5701,N_5826);
or U6876 (N_6876,N_5675,N_5841);
nor U6877 (N_6877,N_5160,N_5482);
or U6878 (N_6878,N_5399,N_5491);
xor U6879 (N_6879,N_5967,N_5501);
and U6880 (N_6880,N_5617,N_5181);
or U6881 (N_6881,N_5765,N_5160);
nand U6882 (N_6882,N_5805,N_5923);
and U6883 (N_6883,N_5073,N_5326);
xnor U6884 (N_6884,N_5566,N_5315);
and U6885 (N_6885,N_5145,N_5039);
nor U6886 (N_6886,N_5170,N_5725);
nand U6887 (N_6887,N_5116,N_5208);
or U6888 (N_6888,N_5248,N_5637);
or U6889 (N_6889,N_5764,N_5763);
nand U6890 (N_6890,N_5233,N_5119);
and U6891 (N_6891,N_5166,N_5270);
xor U6892 (N_6892,N_5128,N_5565);
or U6893 (N_6893,N_5585,N_5241);
nand U6894 (N_6894,N_5685,N_5438);
or U6895 (N_6895,N_5943,N_5140);
nor U6896 (N_6896,N_5221,N_5593);
or U6897 (N_6897,N_5265,N_5783);
nand U6898 (N_6898,N_5557,N_5660);
nand U6899 (N_6899,N_5697,N_5862);
xnor U6900 (N_6900,N_5192,N_5486);
or U6901 (N_6901,N_5979,N_5862);
nand U6902 (N_6902,N_5621,N_5451);
nand U6903 (N_6903,N_5481,N_5027);
and U6904 (N_6904,N_5117,N_5700);
and U6905 (N_6905,N_5839,N_5871);
xor U6906 (N_6906,N_5485,N_5439);
nand U6907 (N_6907,N_5218,N_5733);
nand U6908 (N_6908,N_5674,N_5603);
nor U6909 (N_6909,N_5696,N_5766);
nor U6910 (N_6910,N_5975,N_5115);
nand U6911 (N_6911,N_5007,N_5644);
xor U6912 (N_6912,N_5630,N_5530);
xnor U6913 (N_6913,N_5643,N_5197);
nand U6914 (N_6914,N_5668,N_5940);
and U6915 (N_6915,N_5083,N_5379);
or U6916 (N_6916,N_5989,N_5218);
xor U6917 (N_6917,N_5560,N_5529);
xor U6918 (N_6918,N_5974,N_5036);
xnor U6919 (N_6919,N_5045,N_5635);
nor U6920 (N_6920,N_5411,N_5843);
or U6921 (N_6921,N_5309,N_5952);
xnor U6922 (N_6922,N_5695,N_5690);
nand U6923 (N_6923,N_5957,N_5267);
nand U6924 (N_6924,N_5546,N_5829);
nand U6925 (N_6925,N_5289,N_5982);
and U6926 (N_6926,N_5289,N_5426);
or U6927 (N_6927,N_5202,N_5966);
and U6928 (N_6928,N_5905,N_5099);
xnor U6929 (N_6929,N_5722,N_5885);
nand U6930 (N_6930,N_5940,N_5611);
xor U6931 (N_6931,N_5552,N_5657);
xnor U6932 (N_6932,N_5248,N_5435);
and U6933 (N_6933,N_5223,N_5952);
or U6934 (N_6934,N_5032,N_5338);
xnor U6935 (N_6935,N_5868,N_5996);
and U6936 (N_6936,N_5919,N_5260);
nand U6937 (N_6937,N_5442,N_5035);
or U6938 (N_6938,N_5071,N_5296);
and U6939 (N_6939,N_5570,N_5657);
or U6940 (N_6940,N_5862,N_5263);
and U6941 (N_6941,N_5565,N_5904);
nand U6942 (N_6942,N_5318,N_5888);
nor U6943 (N_6943,N_5866,N_5716);
and U6944 (N_6944,N_5622,N_5560);
nor U6945 (N_6945,N_5868,N_5570);
or U6946 (N_6946,N_5915,N_5797);
xnor U6947 (N_6947,N_5306,N_5262);
and U6948 (N_6948,N_5349,N_5159);
xnor U6949 (N_6949,N_5514,N_5551);
nand U6950 (N_6950,N_5183,N_5626);
or U6951 (N_6951,N_5834,N_5919);
nor U6952 (N_6952,N_5699,N_5921);
nor U6953 (N_6953,N_5721,N_5317);
and U6954 (N_6954,N_5955,N_5322);
xnor U6955 (N_6955,N_5818,N_5536);
or U6956 (N_6956,N_5533,N_5672);
xor U6957 (N_6957,N_5031,N_5243);
nor U6958 (N_6958,N_5437,N_5442);
nor U6959 (N_6959,N_5942,N_5017);
or U6960 (N_6960,N_5727,N_5522);
nand U6961 (N_6961,N_5887,N_5682);
or U6962 (N_6962,N_5350,N_5126);
xnor U6963 (N_6963,N_5690,N_5370);
nor U6964 (N_6964,N_5530,N_5773);
and U6965 (N_6965,N_5548,N_5782);
xnor U6966 (N_6966,N_5750,N_5211);
or U6967 (N_6967,N_5470,N_5778);
and U6968 (N_6968,N_5315,N_5041);
nor U6969 (N_6969,N_5477,N_5300);
nand U6970 (N_6970,N_5981,N_5449);
xor U6971 (N_6971,N_5578,N_5274);
nor U6972 (N_6972,N_5590,N_5519);
nor U6973 (N_6973,N_5616,N_5715);
nand U6974 (N_6974,N_5874,N_5199);
or U6975 (N_6975,N_5608,N_5916);
nand U6976 (N_6976,N_5012,N_5554);
nor U6977 (N_6977,N_5900,N_5757);
or U6978 (N_6978,N_5434,N_5272);
or U6979 (N_6979,N_5529,N_5693);
and U6980 (N_6980,N_5698,N_5957);
or U6981 (N_6981,N_5057,N_5038);
and U6982 (N_6982,N_5441,N_5993);
or U6983 (N_6983,N_5819,N_5283);
and U6984 (N_6984,N_5130,N_5165);
or U6985 (N_6985,N_5741,N_5093);
xor U6986 (N_6986,N_5962,N_5838);
xnor U6987 (N_6987,N_5700,N_5197);
nand U6988 (N_6988,N_5028,N_5701);
nand U6989 (N_6989,N_5635,N_5259);
nor U6990 (N_6990,N_5273,N_5948);
nand U6991 (N_6991,N_5683,N_5162);
nor U6992 (N_6992,N_5845,N_5294);
or U6993 (N_6993,N_5052,N_5148);
nand U6994 (N_6994,N_5626,N_5986);
nor U6995 (N_6995,N_5599,N_5894);
or U6996 (N_6996,N_5460,N_5581);
xor U6997 (N_6997,N_5559,N_5909);
nand U6998 (N_6998,N_5202,N_5356);
nor U6999 (N_6999,N_5266,N_5449);
and U7000 (N_7000,N_6937,N_6133);
and U7001 (N_7001,N_6155,N_6980);
and U7002 (N_7002,N_6029,N_6751);
nor U7003 (N_7003,N_6950,N_6544);
nand U7004 (N_7004,N_6457,N_6865);
xnor U7005 (N_7005,N_6374,N_6215);
and U7006 (N_7006,N_6774,N_6375);
and U7007 (N_7007,N_6110,N_6999);
nor U7008 (N_7008,N_6346,N_6019);
nand U7009 (N_7009,N_6419,N_6669);
xor U7010 (N_7010,N_6461,N_6316);
nor U7011 (N_7011,N_6629,N_6644);
nor U7012 (N_7012,N_6891,N_6422);
nor U7013 (N_7013,N_6895,N_6507);
nor U7014 (N_7014,N_6272,N_6717);
or U7015 (N_7015,N_6556,N_6979);
xor U7016 (N_7016,N_6403,N_6676);
or U7017 (N_7017,N_6801,N_6993);
or U7018 (N_7018,N_6291,N_6223);
nand U7019 (N_7019,N_6872,N_6516);
or U7020 (N_7020,N_6378,N_6615);
nand U7021 (N_7021,N_6884,N_6326);
nand U7022 (N_7022,N_6860,N_6677);
and U7023 (N_7023,N_6286,N_6084);
xor U7024 (N_7024,N_6162,N_6815);
nand U7025 (N_7025,N_6625,N_6092);
or U7026 (N_7026,N_6562,N_6941);
and U7027 (N_7027,N_6227,N_6639);
or U7028 (N_7028,N_6192,N_6067);
xor U7029 (N_7029,N_6696,N_6252);
and U7030 (N_7030,N_6515,N_6060);
nand U7031 (N_7031,N_6525,N_6087);
xor U7032 (N_7032,N_6078,N_6911);
or U7033 (N_7033,N_6915,N_6695);
and U7034 (N_7034,N_6976,N_6796);
and U7035 (N_7035,N_6064,N_6728);
nand U7036 (N_7036,N_6808,N_6267);
xor U7037 (N_7037,N_6641,N_6968);
xor U7038 (N_7038,N_6446,N_6988);
xnor U7039 (N_7039,N_6610,N_6497);
or U7040 (N_7040,N_6372,N_6298);
or U7041 (N_7041,N_6889,N_6052);
nor U7042 (N_7042,N_6727,N_6729);
xor U7043 (N_7043,N_6847,N_6704);
or U7044 (N_7044,N_6118,N_6673);
xnor U7045 (N_7045,N_6505,N_6528);
xor U7046 (N_7046,N_6720,N_6632);
and U7047 (N_7047,N_6420,N_6834);
nand U7048 (N_7048,N_6671,N_6113);
nor U7049 (N_7049,N_6906,N_6569);
nand U7050 (N_7050,N_6638,N_6954);
and U7051 (N_7051,N_6309,N_6255);
nand U7052 (N_7052,N_6091,N_6306);
and U7053 (N_7053,N_6536,N_6646);
xnor U7054 (N_7054,N_6836,N_6703);
nor U7055 (N_7055,N_6220,N_6264);
nor U7056 (N_7056,N_6804,N_6732);
nor U7057 (N_7057,N_6427,N_6382);
or U7058 (N_7058,N_6508,N_6230);
xor U7059 (N_7059,N_6718,N_6780);
nand U7060 (N_7060,N_6406,N_6755);
and U7061 (N_7061,N_6454,N_6885);
nand U7062 (N_7062,N_6626,N_6825);
nand U7063 (N_7063,N_6903,N_6604);
nor U7064 (N_7064,N_6771,N_6736);
nand U7065 (N_7065,N_6417,N_6095);
and U7066 (N_7066,N_6283,N_6691);
nor U7067 (N_7067,N_6074,N_6204);
nor U7068 (N_7068,N_6219,N_6452);
nand U7069 (N_7069,N_6408,N_6441);
nor U7070 (N_7070,N_6111,N_6928);
or U7071 (N_7071,N_6531,N_6085);
xnor U7072 (N_7072,N_6936,N_6036);
or U7073 (N_7073,N_6694,N_6278);
and U7074 (N_7074,N_6352,N_6555);
nor U7075 (N_7075,N_6684,N_6470);
xnor U7076 (N_7076,N_6429,N_6870);
xnor U7077 (N_7077,N_6701,N_6905);
and U7078 (N_7078,N_6044,N_6170);
nand U7079 (N_7079,N_6413,N_6894);
nor U7080 (N_7080,N_6243,N_6586);
xnor U7081 (N_7081,N_6975,N_6135);
or U7082 (N_7082,N_6476,N_6377);
or U7083 (N_7083,N_6921,N_6892);
nand U7084 (N_7084,N_6491,N_6105);
and U7085 (N_7085,N_6364,N_6404);
xnor U7086 (N_7086,N_6966,N_6425);
xnor U7087 (N_7087,N_6855,N_6200);
xor U7088 (N_7088,N_6482,N_6244);
and U7089 (N_7089,N_6518,N_6800);
nor U7090 (N_7090,N_6883,N_6866);
xnor U7091 (N_7091,N_6628,N_6089);
nand U7092 (N_7092,N_6764,N_6724);
xor U7093 (N_7093,N_6940,N_6480);
nand U7094 (N_7094,N_6198,N_6935);
nor U7095 (N_7095,N_6543,N_6462);
or U7096 (N_7096,N_6636,N_6414);
and U7097 (N_7097,N_6265,N_6650);
nand U7098 (N_7098,N_6459,N_6068);
or U7099 (N_7099,N_6767,N_6334);
nand U7100 (N_7100,N_6213,N_6897);
or U7101 (N_7101,N_6124,N_6581);
or U7102 (N_7102,N_6115,N_6246);
and U7103 (N_7103,N_6857,N_6489);
xnor U7104 (N_7104,N_6635,N_6401);
or U7105 (N_7105,N_6288,N_6472);
xor U7106 (N_7106,N_6498,N_6440);
or U7107 (N_7107,N_6754,N_6486);
or U7108 (N_7108,N_6260,N_6186);
or U7109 (N_7109,N_6805,N_6799);
nand U7110 (N_7110,N_6631,N_6465);
nor U7111 (N_7111,N_6978,N_6350);
or U7112 (N_7112,N_6914,N_6475);
or U7113 (N_7113,N_6154,N_6238);
or U7114 (N_7114,N_6959,N_6933);
nor U7115 (N_7115,N_6558,N_6623);
xnor U7116 (N_7116,N_6046,N_6202);
or U7117 (N_7117,N_6524,N_6387);
nor U7118 (N_7118,N_6930,N_6709);
xnor U7119 (N_7119,N_6742,N_6753);
and U7120 (N_7120,N_6484,N_6412);
nor U7121 (N_7121,N_6315,N_6953);
nand U7122 (N_7122,N_6297,N_6195);
nand U7123 (N_7123,N_6426,N_6974);
and U7124 (N_7124,N_6896,N_6149);
xor U7125 (N_7125,N_6539,N_6721);
xor U7126 (N_7126,N_6282,N_6450);
and U7127 (N_7127,N_6770,N_6605);
or U7128 (N_7128,N_6130,N_6136);
or U7129 (N_7129,N_6958,N_6102);
and U7130 (N_7130,N_6431,N_6699);
nand U7131 (N_7131,N_6168,N_6931);
nand U7132 (N_7132,N_6273,N_6062);
xor U7133 (N_7133,N_6416,N_6285);
nor U7134 (N_7134,N_6151,N_6253);
and U7135 (N_7135,N_6358,N_6410);
nand U7136 (N_7136,N_6448,N_6051);
and U7137 (N_7137,N_6494,N_6812);
and U7138 (N_7138,N_6707,N_6400);
nand U7139 (N_7139,N_6792,N_6613);
or U7140 (N_7140,N_6762,N_6349);
nand U7141 (N_7141,N_6787,N_6502);
nor U7142 (N_7142,N_6877,N_6070);
xor U7143 (N_7143,N_6094,N_6066);
and U7144 (N_7144,N_6409,N_6761);
or U7145 (N_7145,N_6561,N_6983);
and U7146 (N_7146,N_6888,N_6816);
nor U7147 (N_7147,N_6225,N_6268);
or U7148 (N_7148,N_6107,N_6361);
and U7149 (N_7149,N_6678,N_6823);
and U7150 (N_7150,N_6863,N_6559);
nor U7151 (N_7151,N_6428,N_6398);
or U7152 (N_7152,N_6777,N_6453);
nand U7153 (N_7153,N_6533,N_6363);
xnor U7154 (N_7154,N_6611,N_6271);
nor U7155 (N_7155,N_6101,N_6464);
and U7156 (N_7156,N_6961,N_6109);
nor U7157 (N_7157,N_6172,N_6584);
and U7158 (N_7158,N_6589,N_6396);
and U7159 (N_7159,N_6250,N_6281);
nor U7160 (N_7160,N_6006,N_6939);
nor U7161 (N_7161,N_6240,N_6784);
xnor U7162 (N_7162,N_6126,N_6967);
xnor U7163 (N_7163,N_6175,N_6634);
nand U7164 (N_7164,N_6045,N_6160);
nand U7165 (N_7165,N_6772,N_6828);
nand U7166 (N_7166,N_6354,N_6934);
or U7167 (N_7167,N_6726,N_6603);
nor U7168 (N_7168,N_6593,N_6367);
nor U7169 (N_7169,N_6547,N_6570);
nor U7170 (N_7170,N_6471,N_6529);
and U7171 (N_7171,N_6731,N_6766);
nor U7172 (N_7172,N_6868,N_6969);
xnor U7173 (N_7173,N_6247,N_6526);
and U7174 (N_7174,N_6768,N_6854);
nor U7175 (N_7175,N_6832,N_6700);
xnor U7176 (N_7176,N_6588,N_6838);
nand U7177 (N_7177,N_6495,N_6830);
or U7178 (N_7178,N_6263,N_6908);
nand U7179 (N_7179,N_6379,N_6577);
or U7180 (N_7180,N_6249,N_6088);
or U7181 (N_7181,N_6312,N_6279);
nand U7182 (N_7182,N_6532,N_6485);
nand U7183 (N_7183,N_6758,N_6234);
nor U7184 (N_7184,N_6948,N_6657);
or U7185 (N_7185,N_6241,N_6106);
nand U7186 (N_7186,N_6926,N_6002);
nor U7187 (N_7187,N_6340,N_6099);
nor U7188 (N_7188,N_6444,N_6519);
xnor U7189 (N_7189,N_6232,N_6293);
or U7190 (N_7190,N_6618,N_6318);
or U7191 (N_7191,N_6027,N_6852);
nand U7192 (N_7192,N_6734,N_6012);
nand U7193 (N_7193,N_6965,N_6917);
and U7194 (N_7194,N_6017,N_6776);
or U7195 (N_7195,N_6411,N_6567);
xnor U7196 (N_7196,N_6007,N_6275);
nor U7197 (N_7197,N_6566,N_6612);
or U7198 (N_7198,N_6276,N_6478);
xor U7199 (N_7199,N_6300,N_6167);
and U7200 (N_7200,N_6713,N_6096);
nor U7201 (N_7201,N_6021,N_6185);
nor U7202 (N_7202,N_6499,N_6919);
or U7203 (N_7203,N_6114,N_6506);
xnor U7204 (N_7204,N_6038,N_6075);
nor U7205 (N_7205,N_6112,N_6127);
nand U7206 (N_7206,N_6817,N_6342);
nor U7207 (N_7207,N_6009,N_6530);
nand U7208 (N_7208,N_6487,N_6756);
nand U7209 (N_7209,N_6209,N_6765);
nand U7210 (N_7210,N_6616,N_6343);
or U7211 (N_7211,N_6913,N_6322);
or U7212 (N_7212,N_6656,N_6233);
or U7213 (N_7213,N_6654,N_6537);
nor U7214 (N_7214,N_6496,N_6998);
nand U7215 (N_7215,N_6806,N_6011);
xor U7216 (N_7216,N_6706,N_6858);
or U7217 (N_7217,N_6191,N_6073);
xnor U7218 (N_7218,N_6097,N_6432);
xor U7219 (N_7219,N_6345,N_6147);
or U7220 (N_7220,N_6504,N_6355);
and U7221 (N_7221,N_6277,N_6134);
and U7222 (N_7222,N_6688,N_6887);
nor U7223 (N_7223,N_6159,N_6781);
xor U7224 (N_7224,N_6550,N_6438);
nor U7225 (N_7225,N_6653,N_6920);
nand U7226 (N_7226,N_6437,N_6090);
xnor U7227 (N_7227,N_6793,N_6189);
nor U7228 (N_7228,N_6982,N_6176);
or U7229 (N_7229,N_6393,N_6986);
and U7230 (N_7230,N_6660,N_6500);
xnor U7231 (N_7231,N_6574,N_6356);
or U7232 (N_7232,N_6128,N_6177);
nor U7233 (N_7233,N_6594,N_6261);
and U7234 (N_7234,N_6972,N_6456);
and U7235 (N_7235,N_6698,N_6788);
nor U7236 (N_7236,N_6809,N_6466);
nor U7237 (N_7237,N_6338,N_6418);
nor U7238 (N_7238,N_6842,N_6328);
nand U7239 (N_7239,N_6879,N_6571);
xor U7240 (N_7240,N_6630,N_6256);
and U7241 (N_7241,N_6757,N_6849);
and U7242 (N_7242,N_6206,N_6295);
or U7243 (N_7243,N_6900,N_6984);
xor U7244 (N_7244,N_6239,N_6122);
nor U7245 (N_7245,N_6037,N_6517);
xnor U7246 (N_7246,N_6479,N_6178);
and U7247 (N_7247,N_6783,N_6861);
nor U7248 (N_7248,N_6455,N_6575);
or U7249 (N_7249,N_6514,N_6080);
nor U7250 (N_7250,N_6150,N_6620);
and U7251 (N_7251,N_6018,N_6977);
xor U7252 (N_7252,N_6347,N_6786);
nand U7253 (N_7253,N_6157,N_6715);
xnor U7254 (N_7254,N_6851,N_6837);
nor U7255 (N_7255,N_6290,N_6014);
nor U7256 (N_7256,N_6296,N_6165);
or U7257 (N_7257,N_6778,N_6308);
nand U7258 (N_7258,N_6910,N_6221);
or U7259 (N_7259,N_6228,N_6633);
and U7260 (N_7260,N_6880,N_6392);
nand U7261 (N_7261,N_6474,N_6143);
xor U7262 (N_7262,N_6994,N_6659);
or U7263 (N_7263,N_6740,N_6946);
or U7264 (N_7264,N_6001,N_6224);
xnor U7265 (N_7265,N_6738,N_6590);
or U7266 (N_7266,N_6775,N_6874);
xor U7267 (N_7267,N_6733,N_6957);
or U7268 (N_7268,N_6871,N_6963);
or U7269 (N_7269,N_6744,N_6047);
or U7270 (N_7270,N_6760,N_6004);
or U7271 (N_7271,N_6752,N_6601);
nand U7272 (N_7272,N_6270,N_6655);
nand U7273 (N_7273,N_6152,N_6469);
nor U7274 (N_7274,N_6875,N_6648);
or U7275 (N_7275,N_6236,N_6840);
xor U7276 (N_7276,N_6680,N_6791);
nor U7277 (N_7277,N_6546,N_6158);
or U7278 (N_7278,N_6645,N_6987);
or U7279 (N_7279,N_6138,N_6811);
nor U7280 (N_7280,N_6366,N_6207);
nor U7281 (N_7281,N_6909,N_6672);
nand U7282 (N_7282,N_6424,N_6376);
xor U7283 (N_7283,N_6449,N_6120);
xnor U7284 (N_7284,N_6031,N_6697);
xnor U7285 (N_7285,N_6055,N_6503);
xnor U7286 (N_7286,N_6662,N_6619);
nand U7287 (N_7287,N_6030,N_6245);
xor U7288 (N_7288,N_6621,N_6063);
and U7289 (N_7289,N_6922,N_6579);
nand U7290 (N_7290,N_6714,N_6121);
and U7291 (N_7291,N_6564,N_6218);
or U7292 (N_7292,N_6082,N_6481);
nand U7293 (N_7293,N_6869,N_6582);
or U7294 (N_7294,N_6723,N_6208);
nand U7295 (N_7295,N_6310,N_6022);
xor U7296 (N_7296,N_6749,N_6553);
nand U7297 (N_7297,N_6527,N_6161);
nand U7298 (N_7298,N_6194,N_6596);
nand U7299 (N_7299,N_6841,N_6054);
and U7300 (N_7300,N_6059,N_6573);
xnor U7301 (N_7301,N_6501,N_6600);
or U7302 (N_7302,N_6899,N_6592);
xor U7303 (N_7303,N_6399,N_6826);
nand U7304 (N_7304,N_6477,N_6269);
and U7305 (N_7305,N_6890,N_6025);
xnor U7306 (N_7306,N_6705,N_6348);
or U7307 (N_7307,N_6551,N_6597);
xor U7308 (N_7308,N_6739,N_6169);
nand U7309 (N_7309,N_6242,N_6985);
nand U7310 (N_7310,N_6214,N_6927);
or U7311 (N_7311,N_6819,N_6443);
nand U7312 (N_7312,N_6490,N_6188);
nor U7313 (N_7313,N_6722,N_6587);
xor U7314 (N_7314,N_6370,N_6179);
nor U7315 (N_7315,N_6992,N_6995);
or U7316 (N_7316,N_6511,N_6435);
nand U7317 (N_7317,N_6302,N_6810);
or U7318 (N_7318,N_6173,N_6952);
xor U7319 (N_7319,N_6081,N_6020);
nor U7320 (N_7320,N_6132,N_6862);
and U7321 (N_7321,N_6026,N_6827);
nand U7322 (N_7322,N_6667,N_6005);
and U7323 (N_7323,N_6924,N_6795);
nand U7324 (N_7324,N_6226,N_6745);
or U7325 (N_7325,N_6434,N_6876);
nor U7326 (N_7326,N_6943,N_6652);
and U7327 (N_7327,N_6509,N_6835);
nor U7328 (N_7328,N_6098,N_6839);
or U7329 (N_7329,N_6436,N_6864);
nor U7330 (N_7330,N_6932,N_6844);
and U7331 (N_7331,N_6108,N_6294);
nor U7332 (N_7332,N_6759,N_6365);
xnor U7333 (N_7333,N_6304,N_6077);
xor U7334 (N_7334,N_6216,N_6665);
or U7335 (N_7335,N_6670,N_6690);
xnor U7336 (N_7336,N_6664,N_6923);
nand U7337 (N_7337,N_6171,N_6492);
xor U7338 (N_7338,N_6702,N_6820);
and U7339 (N_7339,N_6331,N_6708);
nand U7340 (N_7340,N_6327,N_6750);
nand U7341 (N_7341,N_6071,N_6843);
xor U7342 (N_7342,N_6576,N_6821);
or U7343 (N_7343,N_6803,N_6512);
and U7344 (N_7344,N_6148,N_6468);
or U7345 (N_7345,N_6560,N_6989);
nand U7346 (N_7346,N_6997,N_6397);
nor U7347 (N_7347,N_6303,N_6339);
or U7348 (N_7348,N_6488,N_6104);
nand U7349 (N_7349,N_6451,N_6990);
nand U7350 (N_7350,N_6960,N_6320);
or U7351 (N_7351,N_6578,N_6867);
and U7352 (N_7352,N_6853,N_6257);
or U7353 (N_7353,N_6039,N_6423);
or U7354 (N_7354,N_6797,N_6572);
and U7355 (N_7355,N_6146,N_6368);
nor U7356 (N_7356,N_6325,N_6049);
or U7357 (N_7357,N_6785,N_6292);
nor U7358 (N_7358,N_6617,N_6813);
or U7359 (N_7359,N_6510,N_6904);
nor U7360 (N_7360,N_6319,N_6057);
or U7361 (N_7361,N_6898,N_6741);
xor U7362 (N_7362,N_6737,N_6981);
or U7363 (N_7363,N_6607,N_6442);
nand U7364 (N_7364,N_6719,N_6313);
and U7365 (N_7365,N_6140,N_6086);
or U7366 (N_7366,N_6274,N_6061);
nand U7367 (N_7367,N_6802,N_6262);
nor U7368 (N_7368,N_6362,N_6180);
xor U7369 (N_7369,N_6048,N_6034);
xor U7370 (N_7370,N_6693,N_6568);
xnor U7371 (N_7371,N_6235,N_6534);
xnor U7372 (N_7372,N_6415,N_6523);
nor U7373 (N_7373,N_6153,N_6711);
xnor U7374 (N_7374,N_6123,N_6614);
nand U7375 (N_7375,N_6163,N_6380);
and U7376 (N_7376,N_6661,N_6685);
or U7377 (N_7377,N_6015,N_6833);
xor U7378 (N_7378,N_6119,N_6390);
or U7379 (N_7379,N_6773,N_6563);
nand U7380 (N_7380,N_6798,N_6137);
and U7381 (N_7381,N_6846,N_6344);
nand U7382 (N_7382,N_6371,N_6337);
xnor U7383 (N_7383,N_6237,N_6251);
or U7384 (N_7384,N_6254,N_6565);
xnor U7385 (N_7385,N_6217,N_6210);
xnor U7386 (N_7386,N_6712,N_6299);
and U7387 (N_7387,N_6129,N_6058);
and U7388 (N_7388,N_6942,N_6609);
or U7389 (N_7389,N_6807,N_6822);
nor U7390 (N_7390,N_6329,N_6918);
or U7391 (N_7391,N_6181,N_6324);
or U7392 (N_7392,N_6033,N_6013);
xnor U7393 (N_7393,N_6028,N_6043);
or U7394 (N_7394,N_6789,N_6335);
nand U7395 (N_7395,N_6141,N_6580);
nand U7396 (N_7396,N_6991,N_6385);
xor U7397 (N_7397,N_6323,N_6682);
and U7398 (N_7398,N_6203,N_6554);
and U7399 (N_7399,N_6381,N_6955);
xor U7400 (N_7400,N_6336,N_6608);
nand U7401 (N_7401,N_6542,N_6421);
or U7402 (N_7402,N_6683,N_6956);
nor U7403 (N_7403,N_6357,N_6447);
xor U7404 (N_7404,N_6540,N_6845);
xor U7405 (N_7405,N_6032,N_6769);
nor U7406 (N_7406,N_6735,N_6212);
or U7407 (N_7407,N_6710,N_6483);
nor U7408 (N_7408,N_6873,N_6902);
nand U7409 (N_7409,N_6599,N_6595);
and U7410 (N_7410,N_6321,N_6103);
nor U7411 (N_7411,N_6637,N_6301);
and U7412 (N_7412,N_6184,N_6222);
nor U7413 (N_7413,N_6284,N_6716);
and U7414 (N_7414,N_6794,N_6405);
nor U7415 (N_7415,N_6131,N_6395);
and U7416 (N_7416,N_6627,N_6386);
and U7417 (N_7417,N_6541,N_6460);
nor U7418 (N_7418,N_6643,N_6083);
xnor U7419 (N_7419,N_6971,N_6473);
and U7420 (N_7420,N_6287,N_6289);
or U7421 (N_7421,N_6394,N_6023);
or U7422 (N_7422,N_6522,N_6681);
nand U7423 (N_7423,N_6658,N_6231);
nand U7424 (N_7424,N_6763,N_6211);
nor U7425 (N_7425,N_6183,N_6647);
or U7426 (N_7426,N_6258,N_6687);
nor U7427 (N_7427,N_6259,N_6951);
nor U7428 (N_7428,N_6139,N_6583);
and U7429 (N_7429,N_6591,N_6351);
or U7430 (N_7430,N_6818,N_6008);
xor U7431 (N_7431,N_6391,N_6205);
and U7432 (N_7432,N_6886,N_6280);
and U7433 (N_7433,N_6266,N_6493);
nor U7434 (N_7434,N_6521,N_6675);
and U7435 (N_7435,N_6538,N_6445);
nor U7436 (N_7436,N_6925,N_6003);
and U7437 (N_7437,N_6916,N_6663);
xnor U7438 (N_7438,N_6144,N_6035);
or U7439 (N_7439,N_6882,N_6384);
nand U7440 (N_7440,N_6353,N_6166);
xor U7441 (N_7441,N_6467,N_6229);
xnor U7442 (N_7442,N_6407,N_6856);
xnor U7443 (N_7443,N_6458,N_6949);
nor U7444 (N_7444,N_6016,N_6402);
nor U7445 (N_7445,N_6748,N_6651);
nand U7446 (N_7446,N_6305,N_6944);
nor U7447 (N_7447,N_6196,N_6649);
nor U7448 (N_7448,N_6790,N_6042);
or U7449 (N_7449,N_6463,N_6053);
and U7450 (N_7450,N_6929,N_6848);
or U7451 (N_7451,N_6973,N_6624);
nor U7452 (N_7452,N_6557,N_6117);
xnor U7453 (N_7453,N_6193,N_6314);
xnor U7454 (N_7454,N_6552,N_6549);
nor U7455 (N_7455,N_6388,N_6041);
nand U7456 (N_7456,N_6622,N_6142);
nand U7457 (N_7457,N_6674,N_6606);
or U7458 (N_7458,N_6050,N_6640);
or U7459 (N_7459,N_6730,N_6430);
and U7460 (N_7460,N_6174,N_6859);
xnor U7461 (N_7461,N_6545,N_6996);
nor U7462 (N_7462,N_6125,N_6907);
nor U7463 (N_7463,N_6585,N_6182);
xor U7464 (N_7464,N_6201,N_6433);
or U7465 (N_7465,N_6076,N_6389);
and U7466 (N_7466,N_6513,N_6938);
xnor U7467 (N_7467,N_6945,N_6947);
and U7468 (N_7468,N_6330,N_6079);
and U7469 (N_7469,N_6116,N_6056);
or U7470 (N_7470,N_6439,N_6072);
nor U7471 (N_7471,N_6962,N_6850);
nand U7472 (N_7472,N_6598,N_6024);
nand U7473 (N_7473,N_6248,N_6535);
xor U7474 (N_7474,N_6341,N_6878);
or U7475 (N_7475,N_6666,N_6746);
or U7476 (N_7476,N_6197,N_6901);
nor U7477 (N_7477,N_6970,N_6686);
or U7478 (N_7478,N_6743,N_6692);
nor U7479 (N_7479,N_6100,N_6383);
and U7480 (N_7480,N_6782,N_6069);
and U7481 (N_7481,N_6156,N_6725);
nand U7482 (N_7482,N_6779,N_6187);
nand U7483 (N_7483,N_6332,N_6093);
nand U7484 (N_7484,N_6307,N_6145);
and U7485 (N_7485,N_6893,N_6360);
or U7486 (N_7486,N_6311,N_6359);
nand U7487 (N_7487,N_6602,N_6190);
xnor U7488 (N_7488,N_6199,N_6333);
or U7489 (N_7489,N_6668,N_6369);
nor U7490 (N_7490,N_6912,N_6831);
or U7491 (N_7491,N_6373,N_6747);
or U7492 (N_7492,N_6317,N_6824);
nor U7493 (N_7493,N_6548,N_6814);
and U7494 (N_7494,N_6000,N_6829);
nand U7495 (N_7495,N_6679,N_6040);
xor U7496 (N_7496,N_6642,N_6964);
nand U7497 (N_7497,N_6689,N_6065);
xnor U7498 (N_7498,N_6164,N_6881);
nor U7499 (N_7499,N_6010,N_6520);
or U7500 (N_7500,N_6636,N_6702);
nand U7501 (N_7501,N_6434,N_6288);
xnor U7502 (N_7502,N_6134,N_6086);
nand U7503 (N_7503,N_6875,N_6134);
xnor U7504 (N_7504,N_6473,N_6574);
or U7505 (N_7505,N_6273,N_6537);
or U7506 (N_7506,N_6533,N_6112);
or U7507 (N_7507,N_6152,N_6014);
nor U7508 (N_7508,N_6689,N_6713);
or U7509 (N_7509,N_6012,N_6692);
and U7510 (N_7510,N_6343,N_6900);
and U7511 (N_7511,N_6323,N_6042);
nand U7512 (N_7512,N_6978,N_6052);
or U7513 (N_7513,N_6783,N_6286);
and U7514 (N_7514,N_6480,N_6421);
and U7515 (N_7515,N_6236,N_6865);
xnor U7516 (N_7516,N_6537,N_6093);
xnor U7517 (N_7517,N_6677,N_6418);
nor U7518 (N_7518,N_6893,N_6127);
and U7519 (N_7519,N_6201,N_6462);
nor U7520 (N_7520,N_6438,N_6447);
xnor U7521 (N_7521,N_6417,N_6580);
xor U7522 (N_7522,N_6870,N_6449);
nand U7523 (N_7523,N_6149,N_6794);
nand U7524 (N_7524,N_6077,N_6352);
xnor U7525 (N_7525,N_6661,N_6533);
nand U7526 (N_7526,N_6470,N_6815);
nand U7527 (N_7527,N_6899,N_6111);
nor U7528 (N_7528,N_6983,N_6324);
or U7529 (N_7529,N_6860,N_6912);
or U7530 (N_7530,N_6462,N_6794);
xnor U7531 (N_7531,N_6607,N_6955);
and U7532 (N_7532,N_6135,N_6493);
nand U7533 (N_7533,N_6320,N_6560);
or U7534 (N_7534,N_6436,N_6003);
and U7535 (N_7535,N_6607,N_6636);
xnor U7536 (N_7536,N_6754,N_6063);
nor U7537 (N_7537,N_6018,N_6902);
nor U7538 (N_7538,N_6796,N_6977);
or U7539 (N_7539,N_6382,N_6584);
and U7540 (N_7540,N_6962,N_6319);
nor U7541 (N_7541,N_6348,N_6648);
nand U7542 (N_7542,N_6562,N_6646);
xor U7543 (N_7543,N_6773,N_6911);
nand U7544 (N_7544,N_6139,N_6734);
and U7545 (N_7545,N_6050,N_6197);
nand U7546 (N_7546,N_6033,N_6293);
and U7547 (N_7547,N_6723,N_6295);
xnor U7548 (N_7548,N_6626,N_6167);
nor U7549 (N_7549,N_6502,N_6454);
or U7550 (N_7550,N_6205,N_6410);
nand U7551 (N_7551,N_6509,N_6142);
nor U7552 (N_7552,N_6026,N_6997);
and U7553 (N_7553,N_6930,N_6304);
xnor U7554 (N_7554,N_6521,N_6302);
xor U7555 (N_7555,N_6928,N_6179);
xnor U7556 (N_7556,N_6913,N_6556);
nor U7557 (N_7557,N_6368,N_6733);
nor U7558 (N_7558,N_6093,N_6346);
xnor U7559 (N_7559,N_6753,N_6274);
nor U7560 (N_7560,N_6282,N_6352);
and U7561 (N_7561,N_6427,N_6480);
xnor U7562 (N_7562,N_6355,N_6619);
or U7563 (N_7563,N_6934,N_6544);
or U7564 (N_7564,N_6039,N_6061);
and U7565 (N_7565,N_6961,N_6178);
xor U7566 (N_7566,N_6240,N_6091);
nand U7567 (N_7567,N_6242,N_6804);
xor U7568 (N_7568,N_6460,N_6350);
and U7569 (N_7569,N_6194,N_6917);
or U7570 (N_7570,N_6262,N_6474);
and U7571 (N_7571,N_6912,N_6810);
xor U7572 (N_7572,N_6363,N_6344);
or U7573 (N_7573,N_6548,N_6565);
or U7574 (N_7574,N_6647,N_6655);
nor U7575 (N_7575,N_6810,N_6862);
nand U7576 (N_7576,N_6935,N_6584);
nand U7577 (N_7577,N_6877,N_6086);
xnor U7578 (N_7578,N_6464,N_6084);
nand U7579 (N_7579,N_6894,N_6177);
nand U7580 (N_7580,N_6232,N_6475);
nand U7581 (N_7581,N_6192,N_6791);
or U7582 (N_7582,N_6471,N_6789);
nor U7583 (N_7583,N_6232,N_6173);
xnor U7584 (N_7584,N_6624,N_6570);
nand U7585 (N_7585,N_6841,N_6342);
nand U7586 (N_7586,N_6389,N_6518);
xor U7587 (N_7587,N_6105,N_6176);
xnor U7588 (N_7588,N_6288,N_6650);
and U7589 (N_7589,N_6239,N_6864);
nor U7590 (N_7590,N_6843,N_6464);
or U7591 (N_7591,N_6343,N_6830);
and U7592 (N_7592,N_6343,N_6018);
xnor U7593 (N_7593,N_6168,N_6219);
or U7594 (N_7594,N_6544,N_6499);
nor U7595 (N_7595,N_6754,N_6936);
nand U7596 (N_7596,N_6168,N_6704);
nor U7597 (N_7597,N_6633,N_6732);
or U7598 (N_7598,N_6357,N_6121);
nand U7599 (N_7599,N_6492,N_6179);
nand U7600 (N_7600,N_6247,N_6234);
nand U7601 (N_7601,N_6613,N_6303);
or U7602 (N_7602,N_6134,N_6917);
or U7603 (N_7603,N_6379,N_6110);
or U7604 (N_7604,N_6845,N_6856);
and U7605 (N_7605,N_6140,N_6435);
xor U7606 (N_7606,N_6934,N_6115);
and U7607 (N_7607,N_6888,N_6589);
nor U7608 (N_7608,N_6724,N_6609);
nand U7609 (N_7609,N_6601,N_6491);
or U7610 (N_7610,N_6291,N_6511);
xor U7611 (N_7611,N_6145,N_6970);
xor U7612 (N_7612,N_6089,N_6035);
xnor U7613 (N_7613,N_6480,N_6612);
nor U7614 (N_7614,N_6053,N_6848);
nor U7615 (N_7615,N_6281,N_6116);
and U7616 (N_7616,N_6197,N_6812);
xnor U7617 (N_7617,N_6984,N_6477);
xnor U7618 (N_7618,N_6225,N_6303);
xor U7619 (N_7619,N_6903,N_6229);
nor U7620 (N_7620,N_6558,N_6691);
or U7621 (N_7621,N_6558,N_6503);
xor U7622 (N_7622,N_6371,N_6466);
nor U7623 (N_7623,N_6611,N_6126);
xnor U7624 (N_7624,N_6299,N_6174);
xor U7625 (N_7625,N_6629,N_6204);
nor U7626 (N_7626,N_6934,N_6901);
nor U7627 (N_7627,N_6939,N_6627);
and U7628 (N_7628,N_6312,N_6984);
and U7629 (N_7629,N_6164,N_6211);
or U7630 (N_7630,N_6066,N_6674);
nor U7631 (N_7631,N_6492,N_6500);
nor U7632 (N_7632,N_6147,N_6967);
nand U7633 (N_7633,N_6565,N_6818);
nand U7634 (N_7634,N_6057,N_6784);
nor U7635 (N_7635,N_6510,N_6578);
xnor U7636 (N_7636,N_6541,N_6918);
or U7637 (N_7637,N_6043,N_6236);
xnor U7638 (N_7638,N_6404,N_6566);
nand U7639 (N_7639,N_6115,N_6012);
nand U7640 (N_7640,N_6467,N_6439);
or U7641 (N_7641,N_6156,N_6918);
and U7642 (N_7642,N_6032,N_6207);
nand U7643 (N_7643,N_6160,N_6508);
xor U7644 (N_7644,N_6244,N_6446);
xnor U7645 (N_7645,N_6922,N_6327);
xnor U7646 (N_7646,N_6497,N_6072);
xor U7647 (N_7647,N_6984,N_6269);
xnor U7648 (N_7648,N_6369,N_6462);
and U7649 (N_7649,N_6927,N_6889);
xor U7650 (N_7650,N_6707,N_6742);
nor U7651 (N_7651,N_6571,N_6730);
xor U7652 (N_7652,N_6221,N_6506);
nor U7653 (N_7653,N_6261,N_6742);
or U7654 (N_7654,N_6459,N_6757);
nor U7655 (N_7655,N_6960,N_6951);
nand U7656 (N_7656,N_6749,N_6141);
xnor U7657 (N_7657,N_6975,N_6340);
or U7658 (N_7658,N_6563,N_6110);
or U7659 (N_7659,N_6367,N_6268);
nor U7660 (N_7660,N_6908,N_6079);
and U7661 (N_7661,N_6185,N_6377);
and U7662 (N_7662,N_6604,N_6442);
nor U7663 (N_7663,N_6791,N_6113);
nand U7664 (N_7664,N_6872,N_6971);
xnor U7665 (N_7665,N_6326,N_6481);
and U7666 (N_7666,N_6937,N_6748);
nor U7667 (N_7667,N_6349,N_6478);
and U7668 (N_7668,N_6086,N_6325);
xor U7669 (N_7669,N_6167,N_6059);
nor U7670 (N_7670,N_6845,N_6476);
xor U7671 (N_7671,N_6270,N_6654);
and U7672 (N_7672,N_6179,N_6125);
or U7673 (N_7673,N_6555,N_6956);
and U7674 (N_7674,N_6942,N_6798);
nand U7675 (N_7675,N_6119,N_6922);
nand U7676 (N_7676,N_6508,N_6074);
nand U7677 (N_7677,N_6190,N_6708);
and U7678 (N_7678,N_6277,N_6552);
xor U7679 (N_7679,N_6639,N_6184);
nor U7680 (N_7680,N_6488,N_6603);
nand U7681 (N_7681,N_6946,N_6608);
and U7682 (N_7682,N_6293,N_6977);
xor U7683 (N_7683,N_6339,N_6813);
and U7684 (N_7684,N_6343,N_6177);
or U7685 (N_7685,N_6846,N_6421);
nor U7686 (N_7686,N_6850,N_6288);
xor U7687 (N_7687,N_6304,N_6188);
nor U7688 (N_7688,N_6693,N_6998);
nand U7689 (N_7689,N_6759,N_6691);
and U7690 (N_7690,N_6063,N_6223);
or U7691 (N_7691,N_6374,N_6679);
nand U7692 (N_7692,N_6467,N_6767);
or U7693 (N_7693,N_6305,N_6457);
nand U7694 (N_7694,N_6155,N_6660);
and U7695 (N_7695,N_6237,N_6806);
nand U7696 (N_7696,N_6411,N_6445);
or U7697 (N_7697,N_6604,N_6618);
and U7698 (N_7698,N_6138,N_6105);
nand U7699 (N_7699,N_6392,N_6550);
nor U7700 (N_7700,N_6967,N_6036);
and U7701 (N_7701,N_6682,N_6554);
nor U7702 (N_7702,N_6253,N_6166);
nand U7703 (N_7703,N_6002,N_6944);
or U7704 (N_7704,N_6982,N_6378);
nand U7705 (N_7705,N_6130,N_6419);
and U7706 (N_7706,N_6181,N_6604);
and U7707 (N_7707,N_6418,N_6615);
nand U7708 (N_7708,N_6103,N_6608);
xor U7709 (N_7709,N_6381,N_6226);
nor U7710 (N_7710,N_6356,N_6977);
and U7711 (N_7711,N_6340,N_6355);
nor U7712 (N_7712,N_6384,N_6829);
nor U7713 (N_7713,N_6107,N_6321);
xnor U7714 (N_7714,N_6001,N_6047);
nand U7715 (N_7715,N_6313,N_6600);
and U7716 (N_7716,N_6135,N_6756);
and U7717 (N_7717,N_6951,N_6961);
nor U7718 (N_7718,N_6523,N_6721);
and U7719 (N_7719,N_6814,N_6820);
xnor U7720 (N_7720,N_6935,N_6655);
nand U7721 (N_7721,N_6702,N_6134);
and U7722 (N_7722,N_6802,N_6503);
nor U7723 (N_7723,N_6740,N_6004);
xor U7724 (N_7724,N_6114,N_6350);
xnor U7725 (N_7725,N_6081,N_6558);
and U7726 (N_7726,N_6559,N_6318);
and U7727 (N_7727,N_6661,N_6317);
nand U7728 (N_7728,N_6926,N_6338);
and U7729 (N_7729,N_6992,N_6049);
xnor U7730 (N_7730,N_6360,N_6563);
and U7731 (N_7731,N_6970,N_6988);
nand U7732 (N_7732,N_6831,N_6345);
xnor U7733 (N_7733,N_6771,N_6747);
nor U7734 (N_7734,N_6764,N_6195);
and U7735 (N_7735,N_6837,N_6303);
xor U7736 (N_7736,N_6138,N_6507);
nand U7737 (N_7737,N_6771,N_6624);
or U7738 (N_7738,N_6614,N_6598);
and U7739 (N_7739,N_6625,N_6627);
nand U7740 (N_7740,N_6600,N_6668);
nor U7741 (N_7741,N_6980,N_6028);
or U7742 (N_7742,N_6800,N_6153);
nand U7743 (N_7743,N_6974,N_6054);
or U7744 (N_7744,N_6777,N_6021);
nand U7745 (N_7745,N_6896,N_6482);
xor U7746 (N_7746,N_6605,N_6747);
nor U7747 (N_7747,N_6761,N_6143);
or U7748 (N_7748,N_6628,N_6255);
and U7749 (N_7749,N_6074,N_6454);
and U7750 (N_7750,N_6370,N_6877);
and U7751 (N_7751,N_6879,N_6081);
nor U7752 (N_7752,N_6636,N_6915);
xor U7753 (N_7753,N_6095,N_6394);
xor U7754 (N_7754,N_6777,N_6013);
or U7755 (N_7755,N_6006,N_6680);
nor U7756 (N_7756,N_6678,N_6256);
or U7757 (N_7757,N_6670,N_6086);
and U7758 (N_7758,N_6514,N_6569);
or U7759 (N_7759,N_6752,N_6375);
or U7760 (N_7760,N_6405,N_6336);
xor U7761 (N_7761,N_6694,N_6325);
and U7762 (N_7762,N_6793,N_6956);
nand U7763 (N_7763,N_6903,N_6732);
xnor U7764 (N_7764,N_6719,N_6992);
or U7765 (N_7765,N_6702,N_6672);
and U7766 (N_7766,N_6864,N_6096);
and U7767 (N_7767,N_6590,N_6650);
or U7768 (N_7768,N_6003,N_6362);
nor U7769 (N_7769,N_6537,N_6877);
nor U7770 (N_7770,N_6955,N_6851);
and U7771 (N_7771,N_6810,N_6529);
xnor U7772 (N_7772,N_6304,N_6797);
nand U7773 (N_7773,N_6953,N_6444);
nand U7774 (N_7774,N_6441,N_6524);
or U7775 (N_7775,N_6019,N_6276);
nor U7776 (N_7776,N_6813,N_6187);
nand U7777 (N_7777,N_6603,N_6765);
nand U7778 (N_7778,N_6798,N_6946);
nand U7779 (N_7779,N_6257,N_6210);
xnor U7780 (N_7780,N_6669,N_6814);
xor U7781 (N_7781,N_6046,N_6349);
and U7782 (N_7782,N_6596,N_6525);
nor U7783 (N_7783,N_6838,N_6491);
or U7784 (N_7784,N_6633,N_6752);
nor U7785 (N_7785,N_6350,N_6491);
xnor U7786 (N_7786,N_6389,N_6700);
nand U7787 (N_7787,N_6353,N_6697);
or U7788 (N_7788,N_6610,N_6312);
or U7789 (N_7789,N_6007,N_6815);
xor U7790 (N_7790,N_6530,N_6085);
nand U7791 (N_7791,N_6827,N_6204);
or U7792 (N_7792,N_6746,N_6336);
or U7793 (N_7793,N_6479,N_6522);
nand U7794 (N_7794,N_6221,N_6484);
or U7795 (N_7795,N_6590,N_6519);
and U7796 (N_7796,N_6804,N_6709);
nor U7797 (N_7797,N_6742,N_6353);
xnor U7798 (N_7798,N_6634,N_6798);
and U7799 (N_7799,N_6230,N_6879);
or U7800 (N_7800,N_6248,N_6478);
nand U7801 (N_7801,N_6013,N_6548);
and U7802 (N_7802,N_6159,N_6552);
nor U7803 (N_7803,N_6541,N_6317);
nand U7804 (N_7804,N_6760,N_6952);
nor U7805 (N_7805,N_6742,N_6224);
and U7806 (N_7806,N_6457,N_6633);
nor U7807 (N_7807,N_6349,N_6094);
xnor U7808 (N_7808,N_6456,N_6524);
xor U7809 (N_7809,N_6049,N_6489);
xor U7810 (N_7810,N_6267,N_6997);
and U7811 (N_7811,N_6469,N_6670);
nor U7812 (N_7812,N_6824,N_6198);
nor U7813 (N_7813,N_6840,N_6968);
nand U7814 (N_7814,N_6022,N_6507);
or U7815 (N_7815,N_6040,N_6921);
nand U7816 (N_7816,N_6904,N_6939);
xnor U7817 (N_7817,N_6516,N_6290);
xor U7818 (N_7818,N_6340,N_6858);
nor U7819 (N_7819,N_6626,N_6731);
nor U7820 (N_7820,N_6021,N_6757);
or U7821 (N_7821,N_6724,N_6944);
and U7822 (N_7822,N_6767,N_6128);
nor U7823 (N_7823,N_6611,N_6389);
nand U7824 (N_7824,N_6926,N_6344);
and U7825 (N_7825,N_6390,N_6798);
and U7826 (N_7826,N_6217,N_6953);
nand U7827 (N_7827,N_6873,N_6538);
and U7828 (N_7828,N_6931,N_6313);
xnor U7829 (N_7829,N_6465,N_6992);
xor U7830 (N_7830,N_6035,N_6188);
and U7831 (N_7831,N_6082,N_6204);
and U7832 (N_7832,N_6889,N_6952);
xnor U7833 (N_7833,N_6816,N_6814);
nand U7834 (N_7834,N_6758,N_6702);
or U7835 (N_7835,N_6591,N_6173);
nand U7836 (N_7836,N_6734,N_6305);
nand U7837 (N_7837,N_6600,N_6639);
nor U7838 (N_7838,N_6896,N_6302);
xnor U7839 (N_7839,N_6242,N_6301);
xor U7840 (N_7840,N_6224,N_6437);
and U7841 (N_7841,N_6520,N_6851);
or U7842 (N_7842,N_6897,N_6976);
nand U7843 (N_7843,N_6786,N_6072);
nor U7844 (N_7844,N_6261,N_6533);
nor U7845 (N_7845,N_6771,N_6203);
or U7846 (N_7846,N_6781,N_6413);
nand U7847 (N_7847,N_6779,N_6852);
or U7848 (N_7848,N_6634,N_6567);
nor U7849 (N_7849,N_6856,N_6788);
nand U7850 (N_7850,N_6962,N_6548);
and U7851 (N_7851,N_6671,N_6051);
or U7852 (N_7852,N_6323,N_6405);
nor U7853 (N_7853,N_6748,N_6882);
xor U7854 (N_7854,N_6622,N_6150);
and U7855 (N_7855,N_6740,N_6651);
nand U7856 (N_7856,N_6170,N_6637);
or U7857 (N_7857,N_6445,N_6841);
nor U7858 (N_7858,N_6035,N_6647);
xnor U7859 (N_7859,N_6257,N_6510);
nand U7860 (N_7860,N_6977,N_6128);
xnor U7861 (N_7861,N_6722,N_6669);
or U7862 (N_7862,N_6831,N_6358);
and U7863 (N_7863,N_6482,N_6301);
xor U7864 (N_7864,N_6862,N_6305);
nor U7865 (N_7865,N_6337,N_6812);
xor U7866 (N_7866,N_6008,N_6126);
and U7867 (N_7867,N_6233,N_6224);
and U7868 (N_7868,N_6910,N_6432);
nand U7869 (N_7869,N_6665,N_6737);
or U7870 (N_7870,N_6109,N_6340);
or U7871 (N_7871,N_6363,N_6295);
xor U7872 (N_7872,N_6796,N_6833);
nand U7873 (N_7873,N_6733,N_6878);
or U7874 (N_7874,N_6562,N_6900);
xor U7875 (N_7875,N_6076,N_6216);
nor U7876 (N_7876,N_6579,N_6052);
xor U7877 (N_7877,N_6936,N_6488);
and U7878 (N_7878,N_6368,N_6996);
or U7879 (N_7879,N_6707,N_6323);
nand U7880 (N_7880,N_6788,N_6013);
and U7881 (N_7881,N_6702,N_6126);
nand U7882 (N_7882,N_6401,N_6217);
and U7883 (N_7883,N_6644,N_6313);
xor U7884 (N_7884,N_6047,N_6592);
and U7885 (N_7885,N_6471,N_6888);
nand U7886 (N_7886,N_6080,N_6845);
xnor U7887 (N_7887,N_6863,N_6305);
nand U7888 (N_7888,N_6504,N_6736);
or U7889 (N_7889,N_6371,N_6512);
nor U7890 (N_7890,N_6057,N_6174);
or U7891 (N_7891,N_6988,N_6321);
or U7892 (N_7892,N_6797,N_6638);
or U7893 (N_7893,N_6620,N_6302);
nand U7894 (N_7894,N_6277,N_6495);
or U7895 (N_7895,N_6344,N_6282);
nor U7896 (N_7896,N_6097,N_6419);
xnor U7897 (N_7897,N_6372,N_6155);
xnor U7898 (N_7898,N_6834,N_6879);
or U7899 (N_7899,N_6168,N_6108);
nor U7900 (N_7900,N_6890,N_6558);
and U7901 (N_7901,N_6838,N_6427);
and U7902 (N_7902,N_6437,N_6022);
nand U7903 (N_7903,N_6715,N_6844);
or U7904 (N_7904,N_6730,N_6210);
and U7905 (N_7905,N_6779,N_6433);
and U7906 (N_7906,N_6148,N_6421);
nor U7907 (N_7907,N_6040,N_6347);
or U7908 (N_7908,N_6519,N_6346);
xor U7909 (N_7909,N_6227,N_6161);
xnor U7910 (N_7910,N_6366,N_6906);
xor U7911 (N_7911,N_6601,N_6822);
xnor U7912 (N_7912,N_6858,N_6195);
or U7913 (N_7913,N_6063,N_6396);
nand U7914 (N_7914,N_6249,N_6235);
xnor U7915 (N_7915,N_6024,N_6107);
nor U7916 (N_7916,N_6287,N_6636);
nand U7917 (N_7917,N_6189,N_6853);
xnor U7918 (N_7918,N_6182,N_6344);
nand U7919 (N_7919,N_6752,N_6030);
xor U7920 (N_7920,N_6723,N_6658);
and U7921 (N_7921,N_6869,N_6245);
xor U7922 (N_7922,N_6405,N_6498);
xor U7923 (N_7923,N_6602,N_6365);
nor U7924 (N_7924,N_6555,N_6125);
xnor U7925 (N_7925,N_6767,N_6600);
nor U7926 (N_7926,N_6562,N_6779);
nand U7927 (N_7927,N_6081,N_6625);
or U7928 (N_7928,N_6672,N_6253);
xor U7929 (N_7929,N_6439,N_6103);
and U7930 (N_7930,N_6542,N_6238);
and U7931 (N_7931,N_6409,N_6330);
nand U7932 (N_7932,N_6605,N_6827);
nand U7933 (N_7933,N_6494,N_6139);
nand U7934 (N_7934,N_6221,N_6272);
nor U7935 (N_7935,N_6914,N_6786);
and U7936 (N_7936,N_6911,N_6884);
nand U7937 (N_7937,N_6792,N_6079);
nor U7938 (N_7938,N_6223,N_6400);
xor U7939 (N_7939,N_6936,N_6496);
nand U7940 (N_7940,N_6522,N_6884);
xor U7941 (N_7941,N_6505,N_6379);
or U7942 (N_7942,N_6825,N_6210);
or U7943 (N_7943,N_6847,N_6528);
or U7944 (N_7944,N_6984,N_6754);
nor U7945 (N_7945,N_6026,N_6027);
or U7946 (N_7946,N_6694,N_6533);
xor U7947 (N_7947,N_6454,N_6923);
and U7948 (N_7948,N_6056,N_6416);
or U7949 (N_7949,N_6673,N_6384);
and U7950 (N_7950,N_6018,N_6643);
and U7951 (N_7951,N_6182,N_6615);
and U7952 (N_7952,N_6641,N_6738);
and U7953 (N_7953,N_6535,N_6739);
and U7954 (N_7954,N_6190,N_6272);
and U7955 (N_7955,N_6246,N_6845);
nor U7956 (N_7956,N_6195,N_6788);
nor U7957 (N_7957,N_6689,N_6458);
and U7958 (N_7958,N_6652,N_6418);
xnor U7959 (N_7959,N_6894,N_6756);
and U7960 (N_7960,N_6073,N_6323);
and U7961 (N_7961,N_6810,N_6682);
and U7962 (N_7962,N_6350,N_6207);
nand U7963 (N_7963,N_6829,N_6172);
and U7964 (N_7964,N_6891,N_6928);
nand U7965 (N_7965,N_6961,N_6877);
xor U7966 (N_7966,N_6136,N_6898);
or U7967 (N_7967,N_6381,N_6286);
or U7968 (N_7968,N_6765,N_6372);
or U7969 (N_7969,N_6776,N_6757);
and U7970 (N_7970,N_6764,N_6801);
nor U7971 (N_7971,N_6987,N_6970);
and U7972 (N_7972,N_6329,N_6180);
and U7973 (N_7973,N_6642,N_6919);
and U7974 (N_7974,N_6209,N_6428);
xnor U7975 (N_7975,N_6086,N_6618);
xor U7976 (N_7976,N_6066,N_6807);
nor U7977 (N_7977,N_6027,N_6227);
nand U7978 (N_7978,N_6571,N_6134);
nand U7979 (N_7979,N_6662,N_6076);
nand U7980 (N_7980,N_6818,N_6866);
or U7981 (N_7981,N_6574,N_6522);
nand U7982 (N_7982,N_6525,N_6878);
or U7983 (N_7983,N_6779,N_6219);
or U7984 (N_7984,N_6240,N_6516);
xnor U7985 (N_7985,N_6438,N_6981);
xnor U7986 (N_7986,N_6802,N_6011);
xnor U7987 (N_7987,N_6317,N_6482);
nor U7988 (N_7988,N_6737,N_6204);
and U7989 (N_7989,N_6133,N_6015);
xnor U7990 (N_7990,N_6717,N_6660);
xor U7991 (N_7991,N_6995,N_6930);
or U7992 (N_7992,N_6612,N_6710);
or U7993 (N_7993,N_6599,N_6933);
nand U7994 (N_7994,N_6801,N_6372);
nand U7995 (N_7995,N_6646,N_6948);
nand U7996 (N_7996,N_6704,N_6313);
nand U7997 (N_7997,N_6686,N_6856);
xnor U7998 (N_7998,N_6709,N_6531);
and U7999 (N_7999,N_6277,N_6301);
and U8000 (N_8000,N_7445,N_7079);
and U8001 (N_8001,N_7062,N_7148);
and U8002 (N_8002,N_7423,N_7766);
nor U8003 (N_8003,N_7071,N_7518);
and U8004 (N_8004,N_7789,N_7762);
xor U8005 (N_8005,N_7356,N_7939);
or U8006 (N_8006,N_7287,N_7696);
or U8007 (N_8007,N_7143,N_7885);
xnor U8008 (N_8008,N_7723,N_7452);
nand U8009 (N_8009,N_7398,N_7472);
or U8010 (N_8010,N_7305,N_7352);
nand U8011 (N_8011,N_7076,N_7146);
and U8012 (N_8012,N_7659,N_7857);
xor U8013 (N_8013,N_7643,N_7262);
nand U8014 (N_8014,N_7769,N_7375);
and U8015 (N_8015,N_7083,N_7029);
nor U8016 (N_8016,N_7973,N_7531);
nand U8017 (N_8017,N_7403,N_7566);
or U8018 (N_8018,N_7756,N_7955);
nand U8019 (N_8019,N_7249,N_7163);
and U8020 (N_8020,N_7603,N_7720);
or U8021 (N_8021,N_7416,N_7132);
xnor U8022 (N_8022,N_7883,N_7668);
and U8023 (N_8023,N_7000,N_7381);
or U8024 (N_8024,N_7161,N_7248);
nand U8025 (N_8025,N_7015,N_7677);
nor U8026 (N_8026,N_7158,N_7712);
xnor U8027 (N_8027,N_7821,N_7797);
xnor U8028 (N_8028,N_7642,N_7465);
xnor U8029 (N_8029,N_7688,N_7990);
nand U8030 (N_8030,N_7521,N_7820);
nor U8031 (N_8031,N_7063,N_7678);
xnor U8032 (N_8032,N_7611,N_7951);
or U8033 (N_8033,N_7920,N_7354);
or U8034 (N_8034,N_7830,N_7245);
or U8035 (N_8035,N_7285,N_7782);
nor U8036 (N_8036,N_7215,N_7372);
nand U8037 (N_8037,N_7446,N_7036);
and U8038 (N_8038,N_7815,N_7722);
or U8039 (N_8039,N_7099,N_7179);
and U8040 (N_8040,N_7469,N_7786);
and U8041 (N_8041,N_7599,N_7236);
nand U8042 (N_8042,N_7407,N_7186);
xnor U8043 (N_8043,N_7135,N_7093);
or U8044 (N_8044,N_7321,N_7116);
nor U8045 (N_8045,N_7238,N_7964);
nor U8046 (N_8046,N_7967,N_7713);
nand U8047 (N_8047,N_7208,N_7360);
xnor U8048 (N_8048,N_7441,N_7164);
xor U8049 (N_8049,N_7912,N_7960);
nor U8050 (N_8050,N_7202,N_7225);
nor U8051 (N_8051,N_7644,N_7073);
and U8052 (N_8052,N_7190,N_7685);
nand U8053 (N_8053,N_7418,N_7954);
nand U8054 (N_8054,N_7652,N_7796);
nand U8055 (N_8055,N_7223,N_7965);
xor U8056 (N_8056,N_7290,N_7589);
and U8057 (N_8057,N_7046,N_7098);
and U8058 (N_8058,N_7517,N_7201);
or U8059 (N_8059,N_7616,N_7408);
or U8060 (N_8060,N_7315,N_7218);
and U8061 (N_8061,N_7162,N_7676);
xnor U8062 (N_8062,N_7396,N_7667);
xnor U8063 (N_8063,N_7383,N_7868);
xor U8064 (N_8064,N_7590,N_7926);
xor U8065 (N_8065,N_7400,N_7673);
nor U8066 (N_8066,N_7972,N_7010);
and U8067 (N_8067,N_7822,N_7039);
and U8068 (N_8068,N_7368,N_7865);
xnor U8069 (N_8069,N_7543,N_7529);
and U8070 (N_8070,N_7255,N_7414);
xnor U8071 (N_8071,N_7622,N_7332);
xor U8072 (N_8072,N_7749,N_7580);
nand U8073 (N_8073,N_7500,N_7992);
nor U8074 (N_8074,N_7896,N_7573);
xnor U8075 (N_8075,N_7706,N_7933);
and U8076 (N_8076,N_7031,N_7623);
nand U8077 (N_8077,N_7376,N_7358);
nand U8078 (N_8078,N_7625,N_7806);
nand U8079 (N_8079,N_7867,N_7882);
nand U8080 (N_8080,N_7247,N_7264);
nand U8081 (N_8081,N_7359,N_7293);
nor U8082 (N_8082,N_7592,N_7107);
or U8083 (N_8083,N_7212,N_7773);
nand U8084 (N_8084,N_7870,N_7984);
nor U8085 (N_8085,N_7853,N_7856);
or U8086 (N_8086,N_7998,N_7800);
and U8087 (N_8087,N_7204,N_7909);
nor U8088 (N_8088,N_7895,N_7273);
nand U8089 (N_8089,N_7629,N_7008);
or U8090 (N_8090,N_7087,N_7417);
nand U8091 (N_8091,N_7829,N_7980);
and U8092 (N_8092,N_7075,N_7772);
xor U8093 (N_8093,N_7942,N_7138);
nor U8094 (N_8094,N_7096,N_7197);
nor U8095 (N_8095,N_7981,N_7144);
nand U8096 (N_8096,N_7373,N_7346);
and U8097 (N_8097,N_7350,N_7619);
and U8098 (N_8098,N_7489,N_7637);
xor U8099 (N_8099,N_7552,N_7567);
xnor U8100 (N_8100,N_7339,N_7838);
xnor U8101 (N_8101,N_7171,N_7721);
xor U8102 (N_8102,N_7732,N_7985);
xor U8103 (N_8103,N_7938,N_7977);
xnor U8104 (N_8104,N_7627,N_7081);
and U8105 (N_8105,N_7496,N_7279);
nor U8106 (N_8106,N_7934,N_7413);
and U8107 (N_8107,N_7412,N_7329);
or U8108 (N_8108,N_7320,N_7823);
or U8109 (N_8109,N_7549,N_7013);
nor U8110 (N_8110,N_7898,N_7178);
and U8111 (N_8111,N_7269,N_7511);
nor U8112 (N_8112,N_7054,N_7394);
nor U8113 (N_8113,N_7288,N_7494);
xnor U8114 (N_8114,N_7274,N_7594);
xor U8115 (N_8115,N_7251,N_7795);
and U8116 (N_8116,N_7017,N_7224);
nand U8117 (N_8117,N_7211,N_7842);
nor U8118 (N_8118,N_7863,N_7322);
or U8119 (N_8119,N_7940,N_7907);
xnor U8120 (N_8120,N_7957,N_7565);
nand U8121 (N_8121,N_7301,N_7462);
nor U8122 (N_8122,N_7425,N_7740);
nand U8123 (N_8123,N_7026,N_7809);
nand U8124 (N_8124,N_7843,N_7505);
nor U8125 (N_8125,N_7345,N_7207);
and U8126 (N_8126,N_7227,N_7804);
and U8127 (N_8127,N_7139,N_7744);
xnor U8128 (N_8128,N_7560,N_7640);
or U8129 (N_8129,N_7477,N_7457);
nor U8130 (N_8130,N_7378,N_7170);
nand U8131 (N_8131,N_7357,N_7935);
nor U8132 (N_8132,N_7056,N_7554);
xnor U8133 (N_8133,N_7150,N_7509);
nand U8134 (N_8134,N_7950,N_7326);
xnor U8135 (N_8135,N_7522,N_7878);
and U8136 (N_8136,N_7608,N_7600);
or U8137 (N_8137,N_7709,N_7717);
nor U8138 (N_8138,N_7873,N_7818);
xnor U8139 (N_8139,N_7385,N_7118);
nand U8140 (N_8140,N_7193,N_7528);
nor U8141 (N_8141,N_7088,N_7794);
xnor U8142 (N_8142,N_7596,N_7395);
or U8143 (N_8143,N_7695,N_7136);
or U8144 (N_8144,N_7999,N_7877);
nand U8145 (N_8145,N_7324,N_7651);
nor U8146 (N_8146,N_7958,N_7745);
nand U8147 (N_8147,N_7328,N_7239);
nor U8148 (N_8148,N_7149,N_7731);
nor U8149 (N_8149,N_7283,N_7988);
or U8150 (N_8150,N_7504,N_7669);
and U8151 (N_8151,N_7409,N_7854);
xnor U8152 (N_8152,N_7297,N_7100);
nand U8153 (N_8153,N_7012,N_7780);
xnor U8154 (N_8154,N_7027,N_7607);
nor U8155 (N_8155,N_7151,N_7656);
and U8156 (N_8156,N_7562,N_7121);
or U8157 (N_8157,N_7124,N_7181);
and U8158 (N_8158,N_7628,N_7436);
or U8159 (N_8159,N_7890,N_7751);
or U8160 (N_8160,N_7278,N_7473);
or U8161 (N_8161,N_7674,N_7006);
xnor U8162 (N_8162,N_7296,N_7834);
and U8163 (N_8163,N_7793,N_7258);
or U8164 (N_8164,N_7392,N_7771);
and U8165 (N_8165,N_7974,N_7111);
or U8166 (N_8166,N_7022,N_7948);
nor U8167 (N_8167,N_7810,N_7024);
xnor U8168 (N_8168,N_7959,N_7182);
nand U8169 (N_8169,N_7639,N_7591);
xnor U8170 (N_8170,N_7172,N_7754);
and U8171 (N_8171,N_7647,N_7927);
or U8172 (N_8172,N_7219,N_7109);
nand U8173 (N_8173,N_7449,N_7563);
nand U8174 (N_8174,N_7479,N_7739);
nand U8175 (N_8175,N_7270,N_7765);
nand U8176 (N_8176,N_7157,N_7879);
and U8177 (N_8177,N_7604,N_7295);
nand U8178 (N_8178,N_7515,N_7787);
and U8179 (N_8179,N_7750,N_7790);
nor U8180 (N_8180,N_7976,N_7825);
and U8181 (N_8181,N_7314,N_7903);
or U8182 (N_8182,N_7510,N_7388);
xnor U8183 (N_8183,N_7574,N_7451);
nor U8184 (N_8184,N_7911,N_7228);
and U8185 (N_8185,N_7915,N_7078);
and U8186 (N_8186,N_7490,N_7430);
nand U8187 (N_8187,N_7069,N_7516);
and U8188 (N_8188,N_7123,N_7450);
or U8189 (N_8189,N_7371,N_7177);
or U8190 (N_8190,N_7770,N_7011);
nor U8191 (N_8191,N_7281,N_7930);
nand U8192 (N_8192,N_7839,N_7363);
or U8193 (N_8193,N_7003,N_7294);
and U8194 (N_8194,N_7028,N_7606);
nor U8195 (N_8195,N_7620,N_7120);
and U8196 (N_8196,N_7134,N_7658);
nor U8197 (N_8197,N_7716,N_7663);
xnor U8198 (N_8198,N_7259,N_7213);
and U8199 (N_8199,N_7482,N_7798);
and U8200 (N_8200,N_7335,N_7747);
nand U8201 (N_8201,N_7564,N_7913);
nor U8202 (N_8202,N_7699,N_7499);
xor U8203 (N_8203,N_7065,N_7978);
xnor U8204 (N_8204,N_7131,N_7337);
nand U8205 (N_8205,N_7495,N_7308);
or U8206 (N_8206,N_7665,N_7548);
nor U8207 (N_8207,N_7467,N_7864);
xnor U8208 (N_8208,N_7814,N_7090);
nand U8209 (N_8209,N_7317,N_7832);
xnor U8210 (N_8210,N_7953,N_7086);
and U8211 (N_8211,N_7080,N_7544);
and U8212 (N_8212,N_7049,N_7764);
nor U8213 (N_8213,N_7561,N_7602);
xor U8214 (N_8214,N_7894,N_7660);
nand U8215 (N_8215,N_7613,N_7869);
and U8216 (N_8216,N_7682,N_7971);
nand U8217 (N_8217,N_7949,N_7859);
nor U8218 (N_8218,N_7550,N_7995);
or U8219 (N_8219,N_7460,N_7348);
or U8220 (N_8220,N_7817,N_7370);
nand U8221 (N_8221,N_7498,N_7007);
and U8222 (N_8222,N_7729,N_7276);
or U8223 (N_8223,N_7860,N_7167);
nor U8224 (N_8224,N_7897,N_7527);
nand U8225 (N_8225,N_7155,N_7737);
nand U8226 (N_8226,N_7195,N_7648);
and U8227 (N_8227,N_7748,N_7129);
nand U8228 (N_8228,N_7943,N_7066);
nand U8229 (N_8229,N_7827,N_7067);
or U8230 (N_8230,N_7040,N_7057);
and U8231 (N_8231,N_7875,N_7393);
nand U8232 (N_8232,N_7092,N_7196);
xnor U8233 (N_8233,N_7719,N_7921);
nand U8234 (N_8234,N_7997,N_7338);
or U8235 (N_8235,N_7630,N_7014);
or U8236 (N_8236,N_7456,N_7480);
or U8237 (N_8237,N_7657,N_7188);
nand U8238 (N_8238,N_7654,N_7064);
xnor U8239 (N_8239,N_7595,N_7847);
nand U8240 (N_8240,N_7159,N_7443);
and U8241 (N_8241,N_7578,N_7585);
nand U8242 (N_8242,N_7635,N_7519);
nor U8243 (N_8243,N_7174,N_7893);
nand U8244 (N_8244,N_7198,N_7470);
nor U8245 (N_8245,N_7351,N_7537);
or U8246 (N_8246,N_7390,N_7886);
xnor U8247 (N_8247,N_7513,N_7185);
nand U8248 (N_8248,N_7243,N_7979);
and U8249 (N_8249,N_7691,N_7784);
or U8250 (N_8250,N_7961,N_7377);
and U8251 (N_8251,N_7872,N_7240);
or U8252 (N_8252,N_7700,N_7618);
or U8253 (N_8253,N_7349,N_7380);
nor U8254 (N_8254,N_7047,N_7633);
nor U8255 (N_8255,N_7447,N_7914);
or U8256 (N_8256,N_7761,N_7030);
and U8257 (N_8257,N_7871,N_7816);
nand U8258 (N_8258,N_7881,N_7718);
or U8259 (N_8259,N_7636,N_7439);
and U8260 (N_8260,N_7127,N_7369);
xnor U8261 (N_8261,N_7032,N_7837);
and U8262 (N_8262,N_7779,N_7846);
xor U8263 (N_8263,N_7256,N_7753);
nor U8264 (N_8264,N_7097,N_7641);
xor U8265 (N_8265,N_7041,N_7675);
xor U8266 (N_8266,N_7391,N_7508);
and U8267 (N_8267,N_7632,N_7835);
xor U8268 (N_8268,N_7048,N_7267);
nand U8269 (N_8269,N_7891,N_7968);
nand U8270 (N_8270,N_7402,N_7250);
nand U8271 (N_8271,N_7226,N_7541);
xnor U8272 (N_8272,N_7542,N_7776);
and U8273 (N_8273,N_7154,N_7389);
and U8274 (N_8274,N_7956,N_7189);
xor U8275 (N_8275,N_7275,N_7680);
xor U8276 (N_8276,N_7848,N_7145);
nor U8277 (N_8277,N_7698,N_7461);
and U8278 (N_8278,N_7576,N_7952);
nor U8279 (N_8279,N_7438,N_7140);
xnor U8280 (N_8280,N_7852,N_7252);
nand U8281 (N_8281,N_7374,N_7662);
and U8282 (N_8282,N_7650,N_7671);
nand U8283 (N_8283,N_7768,N_7429);
xor U8284 (N_8284,N_7906,N_7001);
nor U8285 (N_8285,N_7191,N_7690);
xor U8286 (N_8286,N_7755,N_7353);
xor U8287 (N_8287,N_7683,N_7535);
and U8288 (N_8288,N_7887,N_7568);
or U8289 (N_8289,N_7432,N_7005);
or U8290 (N_8290,N_7582,N_7058);
xnor U8291 (N_8291,N_7899,N_7944);
nand U8292 (N_8292,N_7532,N_7323);
or U8293 (N_8293,N_7180,N_7733);
or U8294 (N_8294,N_7217,N_7307);
nor U8295 (N_8295,N_7533,N_7042);
nand U8296 (N_8296,N_7741,N_7133);
xnor U8297 (N_8297,N_7476,N_7234);
and U8298 (N_8298,N_7692,N_7593);
and U8299 (N_8299,N_7725,N_7114);
nor U8300 (N_8300,N_7464,N_7597);
and U8301 (N_8301,N_7917,N_7989);
or U8302 (N_8302,N_7319,N_7343);
nand U8303 (N_8303,N_7483,N_7889);
nand U8304 (N_8304,N_7016,N_7728);
xor U8305 (N_8305,N_7703,N_7707);
nand U8306 (N_8306,N_7074,N_7095);
or U8307 (N_8307,N_7840,N_7405);
nand U8308 (N_8308,N_7502,N_7803);
xor U8309 (N_8309,N_7055,N_7963);
xor U8310 (N_8310,N_7468,N_7923);
or U8311 (N_8311,N_7214,N_7849);
nor U8312 (N_8312,N_7697,N_7501);
and U8313 (N_8313,N_7572,N_7649);
nor U8314 (N_8314,N_7406,N_7540);
xor U8315 (N_8315,N_7488,N_7724);
nor U8316 (N_8316,N_7142,N_7993);
xnor U8317 (N_8317,N_7422,N_7702);
nand U8318 (N_8318,N_7059,N_7759);
nor U8319 (N_8319,N_7970,N_7105);
or U8320 (N_8320,N_7424,N_7801);
or U8321 (N_8321,N_7615,N_7002);
nor U8322 (N_8322,N_7404,N_7735);
xor U8323 (N_8323,N_7310,N_7117);
xor U8324 (N_8324,N_7617,N_7888);
nand U8325 (N_8325,N_7113,N_7559);
xnor U8326 (N_8326,N_7653,N_7033);
and U8327 (N_8327,N_7638,N_7525);
or U8328 (N_8328,N_7110,N_7130);
and U8329 (N_8329,N_7431,N_7503);
nor U8330 (N_8330,N_7996,N_7876);
xor U8331 (N_8331,N_7704,N_7126);
xor U8332 (N_8332,N_7119,N_7401);
xnor U8333 (N_8333,N_7426,N_7778);
xnor U8334 (N_8334,N_7428,N_7237);
nand U8335 (N_8335,N_7734,N_7481);
and U8336 (N_8336,N_7021,N_7836);
nand U8337 (N_8337,N_7598,N_7265);
and U8338 (N_8338,N_7601,N_7880);
nor U8339 (N_8339,N_7586,N_7726);
or U8340 (N_8340,N_7280,N_7156);
nor U8341 (N_8341,N_7037,N_7605);
or U8342 (N_8342,N_7901,N_7689);
and U8343 (N_8343,N_7714,N_7947);
nand U8344 (N_8344,N_7845,N_7785);
xor U8345 (N_8345,N_7101,N_7077);
or U8346 (N_8346,N_7813,N_7318);
xor U8347 (N_8347,N_7791,N_7435);
and U8348 (N_8348,N_7681,N_7569);
nand U8349 (N_8349,N_7386,N_7555);
or U8350 (N_8350,N_7742,N_7610);
nor U8351 (N_8351,N_7115,N_7084);
or U8352 (N_8352,N_7705,N_7313);
nor U8353 (N_8353,N_7679,N_7289);
nand U8354 (N_8354,N_7571,N_7106);
or U8355 (N_8355,N_7220,N_7819);
xor U8356 (N_8356,N_7539,N_7851);
and U8357 (N_8357,N_7298,N_7969);
nand U8358 (N_8358,N_7757,N_7327);
nor U8359 (N_8359,N_7112,N_7035);
and U8360 (N_8360,N_7841,N_7304);
nor U8361 (N_8361,N_7104,N_7486);
nor U8362 (N_8362,N_7070,N_7344);
xnor U8363 (N_8363,N_7577,N_7738);
or U8364 (N_8364,N_7900,N_7631);
nand U8365 (N_8365,N_7666,N_7715);
and U8366 (N_8366,N_7799,N_7484);
nand U8367 (N_8367,N_7018,N_7634);
nand U8368 (N_8368,N_7788,N_7254);
nand U8369 (N_8369,N_7986,N_7583);
nand U8370 (N_8370,N_7570,N_7760);
nand U8371 (N_8371,N_7588,N_7670);
nor U8372 (N_8372,N_7458,N_7743);
nand U8373 (N_8373,N_7176,N_7231);
nand U8374 (N_8374,N_7045,N_7205);
xor U8375 (N_8375,N_7340,N_7038);
and U8376 (N_8376,N_7455,N_7474);
or U8377 (N_8377,N_7918,N_7546);
nor U8378 (N_8378,N_7946,N_7165);
and U8379 (N_8379,N_7168,N_7727);
nor U8380 (N_8380,N_7858,N_7802);
or U8381 (N_8381,N_7536,N_7442);
and U8382 (N_8382,N_7526,N_7694);
xnor U8383 (N_8383,N_7701,N_7410);
nand U8384 (N_8384,N_7203,N_7102);
xor U8385 (N_8385,N_7844,N_7466);
and U8386 (N_8386,N_7932,N_7260);
nor U8387 (N_8387,N_7824,N_7050);
nor U8388 (N_8388,N_7922,N_7547);
xor U8389 (N_8389,N_7019,N_7929);
and U8390 (N_8390,N_7434,N_7487);
or U8391 (N_8391,N_7199,N_7708);
nor U8392 (N_8392,N_7299,N_7966);
nand U8393 (N_8393,N_7624,N_7268);
or U8394 (N_8394,N_7257,N_7147);
or U8395 (N_8395,N_7421,N_7261);
nor U8396 (N_8396,N_7085,N_7924);
and U8397 (N_8397,N_7361,N_7246);
nor U8398 (N_8398,N_7061,N_7330);
and U8399 (N_8399,N_7587,N_7686);
xnor U8400 (N_8400,N_7902,N_7684);
or U8401 (N_8401,N_7336,N_7284);
nand U8402 (N_8402,N_7387,N_7277);
xor U8403 (N_8403,N_7448,N_7173);
or U8404 (N_8404,N_7244,N_7614);
nand U8405 (N_8405,N_7263,N_7316);
or U8406 (N_8406,N_7850,N_7553);
xnor U8407 (N_8407,N_7200,N_7271);
nor U8408 (N_8408,N_7463,N_7043);
nor U8409 (N_8409,N_7655,N_7282);
xnor U8410 (N_8410,N_7928,N_7991);
or U8411 (N_8411,N_7538,N_7874);
or U8412 (N_8412,N_7556,N_7910);
xnor U8413 (N_8413,N_7664,N_7491);
nor U8414 (N_8414,N_7206,N_7783);
or U8415 (N_8415,N_7153,N_7411);
and U8416 (N_8416,N_7020,N_7807);
and U8417 (N_8417,N_7730,N_7919);
xor U8418 (N_8418,N_7306,N_7661);
xnor U8419 (N_8419,N_7302,N_7342);
nand U8420 (N_8420,N_7253,N_7053);
or U8421 (N_8421,N_7831,N_7209);
and U8422 (N_8422,N_7364,N_7774);
xor U8423 (N_8423,N_7781,N_7325);
nand U8424 (N_8424,N_7160,N_7497);
or U8425 (N_8425,N_7221,N_7169);
xor U8426 (N_8426,N_7866,N_7397);
nor U8427 (N_8427,N_7646,N_7767);
nor U8428 (N_8428,N_7471,N_7557);
or U8429 (N_8429,N_7621,N_7300);
nand U8430 (N_8430,N_7091,N_7945);
nor U8431 (N_8431,N_7855,N_7808);
xnor U8432 (N_8432,N_7025,N_7693);
nand U8433 (N_8433,N_7524,N_7530);
nand U8434 (N_8434,N_7520,N_7905);
or U8435 (N_8435,N_7506,N_7478);
and U8436 (N_8436,N_7485,N_7908);
and U8437 (N_8437,N_7331,N_7558);
xor U8438 (N_8438,N_7128,N_7068);
xnor U8439 (N_8439,N_7534,N_7379);
or U8440 (N_8440,N_7419,N_7004);
or U8441 (N_8441,N_7475,N_7828);
nand U8442 (N_8442,N_7612,N_7982);
and U8443 (N_8443,N_7312,N_7687);
and U8444 (N_8444,N_7672,N_7975);
xnor U8445 (N_8445,N_7812,N_7175);
nor U8446 (N_8446,N_7861,N_7235);
or U8447 (N_8447,N_7763,N_7232);
and U8448 (N_8448,N_7309,N_7266);
xnor U8449 (N_8449,N_7303,N_7384);
or U8450 (N_8450,N_7194,N_7711);
or U8451 (N_8451,N_7420,N_7453);
nor U8452 (N_8452,N_7184,N_7454);
nand U8453 (N_8453,N_7884,N_7437);
nand U8454 (N_8454,N_7507,N_7962);
xor U8455 (N_8455,N_7365,N_7805);
nor U8456 (N_8456,N_7183,N_7862);
xnor U8457 (N_8457,N_7272,N_7925);
nand U8458 (N_8458,N_7645,N_7433);
nand U8459 (N_8459,N_7366,N_7931);
or U8460 (N_8460,N_7286,N_7009);
xnor U8461 (N_8461,N_7125,N_7415);
xnor U8462 (N_8462,N_7034,N_7994);
nor U8463 (N_8463,N_7523,N_7492);
nor U8464 (N_8464,N_7052,N_7626);
xor U8465 (N_8465,N_7609,N_7459);
nor U8466 (N_8466,N_7108,N_7103);
xor U8467 (N_8467,N_7941,N_7192);
and U8468 (N_8468,N_7241,N_7752);
and U8469 (N_8469,N_7382,N_7233);
nand U8470 (N_8470,N_7579,N_7230);
or U8471 (N_8471,N_7216,N_7936);
nand U8472 (N_8472,N_7341,N_7089);
and U8473 (N_8473,N_7166,N_7427);
nand U8474 (N_8474,N_7347,N_7444);
nand U8475 (N_8475,N_7229,N_7334);
nand U8476 (N_8476,N_7833,N_7575);
and U8477 (N_8477,N_7362,N_7210);
nor U8478 (N_8478,N_7983,N_7367);
or U8479 (N_8479,N_7551,N_7937);
nor U8480 (N_8480,N_7122,N_7023);
nand U8481 (N_8481,N_7222,N_7892);
or U8482 (N_8482,N_7060,N_7584);
or U8483 (N_8483,N_7141,N_7545);
or U8484 (N_8484,N_7137,N_7072);
or U8485 (N_8485,N_7311,N_7811);
xor U8486 (N_8486,N_7493,N_7333);
or U8487 (N_8487,N_7746,N_7904);
and U8488 (N_8488,N_7082,N_7355);
and U8489 (N_8489,N_7792,N_7440);
or U8490 (N_8490,N_7291,N_7187);
or U8491 (N_8491,N_7051,N_7736);
nand U8492 (N_8492,N_7512,N_7152);
or U8493 (N_8493,N_7916,N_7242);
nor U8494 (N_8494,N_7758,N_7581);
xnor U8495 (N_8495,N_7987,N_7777);
xnor U8496 (N_8496,N_7292,N_7826);
nand U8497 (N_8497,N_7094,N_7044);
xnor U8498 (N_8498,N_7710,N_7514);
nor U8499 (N_8499,N_7775,N_7399);
xnor U8500 (N_8500,N_7684,N_7024);
nor U8501 (N_8501,N_7623,N_7186);
and U8502 (N_8502,N_7233,N_7982);
or U8503 (N_8503,N_7904,N_7958);
xor U8504 (N_8504,N_7087,N_7358);
nor U8505 (N_8505,N_7453,N_7675);
nand U8506 (N_8506,N_7741,N_7078);
nor U8507 (N_8507,N_7207,N_7179);
nor U8508 (N_8508,N_7173,N_7376);
nor U8509 (N_8509,N_7354,N_7993);
nand U8510 (N_8510,N_7316,N_7794);
or U8511 (N_8511,N_7662,N_7218);
or U8512 (N_8512,N_7825,N_7907);
or U8513 (N_8513,N_7694,N_7584);
and U8514 (N_8514,N_7101,N_7073);
xor U8515 (N_8515,N_7134,N_7696);
nand U8516 (N_8516,N_7832,N_7973);
or U8517 (N_8517,N_7967,N_7576);
nand U8518 (N_8518,N_7344,N_7341);
nor U8519 (N_8519,N_7864,N_7120);
xor U8520 (N_8520,N_7879,N_7242);
nor U8521 (N_8521,N_7493,N_7386);
and U8522 (N_8522,N_7769,N_7435);
nor U8523 (N_8523,N_7246,N_7868);
xor U8524 (N_8524,N_7276,N_7898);
and U8525 (N_8525,N_7882,N_7183);
and U8526 (N_8526,N_7996,N_7575);
nand U8527 (N_8527,N_7659,N_7771);
nand U8528 (N_8528,N_7820,N_7180);
nand U8529 (N_8529,N_7729,N_7851);
nor U8530 (N_8530,N_7301,N_7036);
or U8531 (N_8531,N_7587,N_7002);
xnor U8532 (N_8532,N_7539,N_7482);
nand U8533 (N_8533,N_7066,N_7913);
and U8534 (N_8534,N_7567,N_7914);
and U8535 (N_8535,N_7423,N_7601);
xnor U8536 (N_8536,N_7906,N_7961);
nand U8537 (N_8537,N_7542,N_7340);
and U8538 (N_8538,N_7641,N_7259);
nand U8539 (N_8539,N_7979,N_7263);
or U8540 (N_8540,N_7688,N_7424);
nand U8541 (N_8541,N_7425,N_7356);
nand U8542 (N_8542,N_7012,N_7777);
and U8543 (N_8543,N_7406,N_7240);
or U8544 (N_8544,N_7601,N_7827);
and U8545 (N_8545,N_7787,N_7553);
and U8546 (N_8546,N_7258,N_7969);
and U8547 (N_8547,N_7043,N_7772);
nor U8548 (N_8548,N_7391,N_7188);
xor U8549 (N_8549,N_7701,N_7453);
or U8550 (N_8550,N_7078,N_7869);
nor U8551 (N_8551,N_7059,N_7918);
nor U8552 (N_8552,N_7009,N_7497);
or U8553 (N_8553,N_7162,N_7830);
xnor U8554 (N_8554,N_7879,N_7213);
nor U8555 (N_8555,N_7291,N_7317);
nor U8556 (N_8556,N_7381,N_7616);
nor U8557 (N_8557,N_7968,N_7834);
xnor U8558 (N_8558,N_7530,N_7128);
xnor U8559 (N_8559,N_7657,N_7873);
and U8560 (N_8560,N_7045,N_7338);
and U8561 (N_8561,N_7821,N_7560);
nand U8562 (N_8562,N_7359,N_7369);
nor U8563 (N_8563,N_7358,N_7026);
nor U8564 (N_8564,N_7642,N_7360);
xor U8565 (N_8565,N_7888,N_7105);
xnor U8566 (N_8566,N_7868,N_7871);
and U8567 (N_8567,N_7077,N_7909);
and U8568 (N_8568,N_7828,N_7523);
nor U8569 (N_8569,N_7402,N_7769);
nand U8570 (N_8570,N_7760,N_7076);
or U8571 (N_8571,N_7391,N_7646);
and U8572 (N_8572,N_7558,N_7282);
or U8573 (N_8573,N_7545,N_7335);
xnor U8574 (N_8574,N_7408,N_7603);
and U8575 (N_8575,N_7597,N_7077);
and U8576 (N_8576,N_7859,N_7295);
nor U8577 (N_8577,N_7385,N_7964);
and U8578 (N_8578,N_7865,N_7900);
xnor U8579 (N_8579,N_7029,N_7458);
nand U8580 (N_8580,N_7700,N_7271);
nand U8581 (N_8581,N_7046,N_7101);
and U8582 (N_8582,N_7786,N_7481);
nor U8583 (N_8583,N_7198,N_7166);
or U8584 (N_8584,N_7155,N_7540);
xnor U8585 (N_8585,N_7633,N_7540);
and U8586 (N_8586,N_7463,N_7384);
and U8587 (N_8587,N_7576,N_7487);
nor U8588 (N_8588,N_7259,N_7488);
xor U8589 (N_8589,N_7261,N_7707);
or U8590 (N_8590,N_7983,N_7640);
and U8591 (N_8591,N_7732,N_7619);
nand U8592 (N_8592,N_7428,N_7518);
or U8593 (N_8593,N_7496,N_7249);
nand U8594 (N_8594,N_7474,N_7829);
nor U8595 (N_8595,N_7276,N_7783);
xor U8596 (N_8596,N_7044,N_7028);
nand U8597 (N_8597,N_7671,N_7806);
or U8598 (N_8598,N_7719,N_7173);
nand U8599 (N_8599,N_7424,N_7114);
and U8600 (N_8600,N_7305,N_7160);
and U8601 (N_8601,N_7451,N_7113);
nand U8602 (N_8602,N_7394,N_7786);
xnor U8603 (N_8603,N_7266,N_7990);
or U8604 (N_8604,N_7994,N_7534);
xor U8605 (N_8605,N_7245,N_7464);
xnor U8606 (N_8606,N_7046,N_7128);
nor U8607 (N_8607,N_7749,N_7408);
xnor U8608 (N_8608,N_7139,N_7964);
or U8609 (N_8609,N_7165,N_7436);
and U8610 (N_8610,N_7411,N_7073);
xor U8611 (N_8611,N_7293,N_7232);
nand U8612 (N_8612,N_7799,N_7598);
or U8613 (N_8613,N_7201,N_7116);
or U8614 (N_8614,N_7074,N_7794);
or U8615 (N_8615,N_7367,N_7098);
or U8616 (N_8616,N_7943,N_7330);
nor U8617 (N_8617,N_7409,N_7843);
and U8618 (N_8618,N_7777,N_7538);
or U8619 (N_8619,N_7930,N_7029);
and U8620 (N_8620,N_7631,N_7419);
nand U8621 (N_8621,N_7712,N_7113);
and U8622 (N_8622,N_7915,N_7477);
nand U8623 (N_8623,N_7256,N_7733);
nand U8624 (N_8624,N_7801,N_7176);
or U8625 (N_8625,N_7029,N_7312);
or U8626 (N_8626,N_7108,N_7027);
nand U8627 (N_8627,N_7971,N_7101);
and U8628 (N_8628,N_7550,N_7531);
and U8629 (N_8629,N_7947,N_7233);
and U8630 (N_8630,N_7380,N_7465);
nor U8631 (N_8631,N_7693,N_7164);
nand U8632 (N_8632,N_7077,N_7641);
or U8633 (N_8633,N_7608,N_7110);
or U8634 (N_8634,N_7963,N_7890);
nor U8635 (N_8635,N_7598,N_7947);
nand U8636 (N_8636,N_7882,N_7481);
and U8637 (N_8637,N_7412,N_7555);
nor U8638 (N_8638,N_7662,N_7373);
and U8639 (N_8639,N_7672,N_7923);
xnor U8640 (N_8640,N_7438,N_7281);
nor U8641 (N_8641,N_7346,N_7176);
xnor U8642 (N_8642,N_7476,N_7080);
and U8643 (N_8643,N_7082,N_7822);
and U8644 (N_8644,N_7855,N_7783);
nand U8645 (N_8645,N_7022,N_7496);
nor U8646 (N_8646,N_7296,N_7521);
or U8647 (N_8647,N_7251,N_7738);
nor U8648 (N_8648,N_7630,N_7944);
or U8649 (N_8649,N_7285,N_7499);
and U8650 (N_8650,N_7367,N_7638);
nor U8651 (N_8651,N_7334,N_7287);
or U8652 (N_8652,N_7981,N_7990);
xnor U8653 (N_8653,N_7002,N_7859);
xor U8654 (N_8654,N_7891,N_7203);
and U8655 (N_8655,N_7899,N_7406);
xnor U8656 (N_8656,N_7040,N_7379);
xnor U8657 (N_8657,N_7347,N_7114);
xor U8658 (N_8658,N_7311,N_7731);
or U8659 (N_8659,N_7737,N_7361);
and U8660 (N_8660,N_7743,N_7681);
nor U8661 (N_8661,N_7756,N_7800);
or U8662 (N_8662,N_7300,N_7213);
or U8663 (N_8663,N_7314,N_7259);
nor U8664 (N_8664,N_7792,N_7333);
nor U8665 (N_8665,N_7107,N_7494);
and U8666 (N_8666,N_7088,N_7756);
and U8667 (N_8667,N_7091,N_7171);
xor U8668 (N_8668,N_7352,N_7593);
and U8669 (N_8669,N_7646,N_7780);
nand U8670 (N_8670,N_7102,N_7985);
or U8671 (N_8671,N_7135,N_7574);
xnor U8672 (N_8672,N_7553,N_7608);
and U8673 (N_8673,N_7556,N_7525);
nand U8674 (N_8674,N_7035,N_7628);
and U8675 (N_8675,N_7906,N_7045);
xnor U8676 (N_8676,N_7041,N_7279);
xnor U8677 (N_8677,N_7955,N_7626);
nand U8678 (N_8678,N_7266,N_7248);
or U8679 (N_8679,N_7319,N_7511);
nor U8680 (N_8680,N_7774,N_7570);
xnor U8681 (N_8681,N_7524,N_7595);
or U8682 (N_8682,N_7660,N_7968);
nand U8683 (N_8683,N_7608,N_7542);
nand U8684 (N_8684,N_7985,N_7207);
xnor U8685 (N_8685,N_7931,N_7992);
xor U8686 (N_8686,N_7793,N_7587);
or U8687 (N_8687,N_7753,N_7743);
nand U8688 (N_8688,N_7211,N_7004);
nor U8689 (N_8689,N_7314,N_7726);
and U8690 (N_8690,N_7259,N_7921);
nand U8691 (N_8691,N_7630,N_7113);
nor U8692 (N_8692,N_7117,N_7971);
nand U8693 (N_8693,N_7088,N_7702);
nor U8694 (N_8694,N_7199,N_7289);
nor U8695 (N_8695,N_7300,N_7161);
nand U8696 (N_8696,N_7157,N_7888);
or U8697 (N_8697,N_7681,N_7040);
and U8698 (N_8698,N_7218,N_7071);
nand U8699 (N_8699,N_7928,N_7725);
xor U8700 (N_8700,N_7212,N_7226);
and U8701 (N_8701,N_7230,N_7679);
and U8702 (N_8702,N_7073,N_7945);
or U8703 (N_8703,N_7485,N_7892);
nand U8704 (N_8704,N_7201,N_7619);
or U8705 (N_8705,N_7580,N_7791);
nand U8706 (N_8706,N_7644,N_7165);
or U8707 (N_8707,N_7690,N_7412);
nor U8708 (N_8708,N_7783,N_7738);
nor U8709 (N_8709,N_7411,N_7167);
or U8710 (N_8710,N_7862,N_7852);
or U8711 (N_8711,N_7219,N_7431);
xnor U8712 (N_8712,N_7503,N_7809);
nand U8713 (N_8713,N_7056,N_7714);
and U8714 (N_8714,N_7549,N_7911);
nand U8715 (N_8715,N_7310,N_7285);
xor U8716 (N_8716,N_7196,N_7733);
and U8717 (N_8717,N_7162,N_7053);
xnor U8718 (N_8718,N_7585,N_7154);
xnor U8719 (N_8719,N_7653,N_7464);
and U8720 (N_8720,N_7177,N_7232);
nand U8721 (N_8721,N_7342,N_7946);
or U8722 (N_8722,N_7943,N_7184);
nor U8723 (N_8723,N_7898,N_7730);
xor U8724 (N_8724,N_7965,N_7240);
xnor U8725 (N_8725,N_7214,N_7361);
and U8726 (N_8726,N_7893,N_7153);
nor U8727 (N_8727,N_7839,N_7931);
nand U8728 (N_8728,N_7969,N_7599);
or U8729 (N_8729,N_7372,N_7580);
xnor U8730 (N_8730,N_7513,N_7610);
nor U8731 (N_8731,N_7553,N_7700);
nor U8732 (N_8732,N_7292,N_7527);
nand U8733 (N_8733,N_7298,N_7122);
and U8734 (N_8734,N_7320,N_7231);
xor U8735 (N_8735,N_7243,N_7663);
nand U8736 (N_8736,N_7444,N_7165);
or U8737 (N_8737,N_7529,N_7302);
nor U8738 (N_8738,N_7953,N_7287);
nand U8739 (N_8739,N_7395,N_7628);
xor U8740 (N_8740,N_7716,N_7309);
or U8741 (N_8741,N_7388,N_7357);
nand U8742 (N_8742,N_7969,N_7195);
and U8743 (N_8743,N_7166,N_7743);
or U8744 (N_8744,N_7350,N_7533);
and U8745 (N_8745,N_7847,N_7205);
or U8746 (N_8746,N_7147,N_7507);
nand U8747 (N_8747,N_7783,N_7235);
nand U8748 (N_8748,N_7495,N_7122);
and U8749 (N_8749,N_7283,N_7669);
nor U8750 (N_8750,N_7589,N_7697);
and U8751 (N_8751,N_7244,N_7808);
nand U8752 (N_8752,N_7660,N_7773);
nand U8753 (N_8753,N_7782,N_7737);
nand U8754 (N_8754,N_7516,N_7150);
nor U8755 (N_8755,N_7236,N_7797);
xnor U8756 (N_8756,N_7280,N_7601);
nor U8757 (N_8757,N_7382,N_7163);
and U8758 (N_8758,N_7791,N_7182);
or U8759 (N_8759,N_7462,N_7979);
and U8760 (N_8760,N_7309,N_7084);
nand U8761 (N_8761,N_7017,N_7788);
or U8762 (N_8762,N_7658,N_7095);
xnor U8763 (N_8763,N_7317,N_7170);
or U8764 (N_8764,N_7322,N_7005);
nand U8765 (N_8765,N_7892,N_7625);
or U8766 (N_8766,N_7681,N_7757);
nand U8767 (N_8767,N_7058,N_7635);
or U8768 (N_8768,N_7585,N_7317);
xor U8769 (N_8769,N_7154,N_7547);
and U8770 (N_8770,N_7245,N_7553);
nor U8771 (N_8771,N_7267,N_7912);
xnor U8772 (N_8772,N_7554,N_7371);
nand U8773 (N_8773,N_7844,N_7106);
nand U8774 (N_8774,N_7338,N_7873);
xor U8775 (N_8775,N_7861,N_7934);
nor U8776 (N_8776,N_7848,N_7565);
and U8777 (N_8777,N_7560,N_7431);
nor U8778 (N_8778,N_7756,N_7806);
nand U8779 (N_8779,N_7578,N_7659);
nand U8780 (N_8780,N_7503,N_7328);
nor U8781 (N_8781,N_7912,N_7199);
xor U8782 (N_8782,N_7425,N_7342);
nand U8783 (N_8783,N_7463,N_7412);
and U8784 (N_8784,N_7296,N_7955);
and U8785 (N_8785,N_7724,N_7951);
and U8786 (N_8786,N_7921,N_7087);
or U8787 (N_8787,N_7153,N_7776);
nor U8788 (N_8788,N_7633,N_7457);
nand U8789 (N_8789,N_7882,N_7634);
and U8790 (N_8790,N_7626,N_7260);
nand U8791 (N_8791,N_7764,N_7258);
xor U8792 (N_8792,N_7615,N_7975);
nand U8793 (N_8793,N_7315,N_7012);
or U8794 (N_8794,N_7844,N_7599);
and U8795 (N_8795,N_7748,N_7314);
or U8796 (N_8796,N_7879,N_7117);
and U8797 (N_8797,N_7304,N_7199);
or U8798 (N_8798,N_7967,N_7715);
nor U8799 (N_8799,N_7407,N_7272);
or U8800 (N_8800,N_7511,N_7023);
xor U8801 (N_8801,N_7968,N_7486);
or U8802 (N_8802,N_7653,N_7770);
nor U8803 (N_8803,N_7825,N_7856);
or U8804 (N_8804,N_7912,N_7239);
nor U8805 (N_8805,N_7357,N_7257);
nand U8806 (N_8806,N_7412,N_7032);
or U8807 (N_8807,N_7340,N_7513);
or U8808 (N_8808,N_7507,N_7817);
nor U8809 (N_8809,N_7671,N_7346);
xor U8810 (N_8810,N_7760,N_7597);
or U8811 (N_8811,N_7087,N_7222);
and U8812 (N_8812,N_7683,N_7577);
nand U8813 (N_8813,N_7266,N_7484);
xnor U8814 (N_8814,N_7583,N_7528);
nor U8815 (N_8815,N_7592,N_7318);
or U8816 (N_8816,N_7568,N_7792);
nor U8817 (N_8817,N_7518,N_7249);
nor U8818 (N_8818,N_7439,N_7527);
xnor U8819 (N_8819,N_7013,N_7350);
nand U8820 (N_8820,N_7752,N_7598);
xor U8821 (N_8821,N_7074,N_7900);
nor U8822 (N_8822,N_7697,N_7154);
nor U8823 (N_8823,N_7825,N_7828);
nor U8824 (N_8824,N_7452,N_7820);
xnor U8825 (N_8825,N_7375,N_7006);
nor U8826 (N_8826,N_7958,N_7254);
nand U8827 (N_8827,N_7128,N_7488);
nor U8828 (N_8828,N_7595,N_7328);
and U8829 (N_8829,N_7207,N_7678);
nor U8830 (N_8830,N_7003,N_7968);
and U8831 (N_8831,N_7474,N_7037);
and U8832 (N_8832,N_7639,N_7618);
and U8833 (N_8833,N_7907,N_7930);
and U8834 (N_8834,N_7394,N_7804);
nor U8835 (N_8835,N_7075,N_7831);
or U8836 (N_8836,N_7191,N_7046);
or U8837 (N_8837,N_7855,N_7623);
xor U8838 (N_8838,N_7969,N_7812);
xor U8839 (N_8839,N_7979,N_7745);
or U8840 (N_8840,N_7851,N_7960);
nor U8841 (N_8841,N_7582,N_7700);
nand U8842 (N_8842,N_7355,N_7185);
nand U8843 (N_8843,N_7996,N_7897);
xnor U8844 (N_8844,N_7710,N_7647);
and U8845 (N_8845,N_7291,N_7012);
xor U8846 (N_8846,N_7805,N_7654);
nor U8847 (N_8847,N_7268,N_7103);
xnor U8848 (N_8848,N_7458,N_7850);
nand U8849 (N_8849,N_7081,N_7393);
nand U8850 (N_8850,N_7630,N_7736);
nand U8851 (N_8851,N_7121,N_7316);
xor U8852 (N_8852,N_7455,N_7926);
or U8853 (N_8853,N_7050,N_7883);
nand U8854 (N_8854,N_7209,N_7215);
nor U8855 (N_8855,N_7946,N_7346);
and U8856 (N_8856,N_7384,N_7701);
or U8857 (N_8857,N_7208,N_7988);
xor U8858 (N_8858,N_7672,N_7232);
or U8859 (N_8859,N_7929,N_7175);
and U8860 (N_8860,N_7127,N_7687);
nor U8861 (N_8861,N_7232,N_7686);
nor U8862 (N_8862,N_7041,N_7203);
or U8863 (N_8863,N_7140,N_7187);
and U8864 (N_8864,N_7284,N_7943);
xor U8865 (N_8865,N_7105,N_7869);
nor U8866 (N_8866,N_7103,N_7904);
or U8867 (N_8867,N_7420,N_7896);
xnor U8868 (N_8868,N_7778,N_7070);
xor U8869 (N_8869,N_7366,N_7632);
nor U8870 (N_8870,N_7606,N_7815);
and U8871 (N_8871,N_7378,N_7501);
or U8872 (N_8872,N_7063,N_7056);
nor U8873 (N_8873,N_7015,N_7186);
xor U8874 (N_8874,N_7155,N_7902);
and U8875 (N_8875,N_7330,N_7378);
xnor U8876 (N_8876,N_7336,N_7976);
or U8877 (N_8877,N_7023,N_7299);
or U8878 (N_8878,N_7389,N_7764);
and U8879 (N_8879,N_7593,N_7040);
or U8880 (N_8880,N_7137,N_7115);
or U8881 (N_8881,N_7478,N_7489);
or U8882 (N_8882,N_7159,N_7600);
nand U8883 (N_8883,N_7492,N_7864);
nor U8884 (N_8884,N_7769,N_7452);
nor U8885 (N_8885,N_7251,N_7503);
nor U8886 (N_8886,N_7551,N_7995);
xnor U8887 (N_8887,N_7641,N_7844);
and U8888 (N_8888,N_7796,N_7532);
or U8889 (N_8889,N_7428,N_7252);
nor U8890 (N_8890,N_7316,N_7839);
nand U8891 (N_8891,N_7865,N_7942);
xnor U8892 (N_8892,N_7884,N_7170);
or U8893 (N_8893,N_7801,N_7324);
and U8894 (N_8894,N_7887,N_7547);
xnor U8895 (N_8895,N_7522,N_7280);
or U8896 (N_8896,N_7424,N_7920);
nand U8897 (N_8897,N_7017,N_7242);
and U8898 (N_8898,N_7284,N_7566);
xor U8899 (N_8899,N_7938,N_7837);
nor U8900 (N_8900,N_7791,N_7887);
or U8901 (N_8901,N_7445,N_7350);
nor U8902 (N_8902,N_7264,N_7516);
or U8903 (N_8903,N_7887,N_7679);
nor U8904 (N_8904,N_7224,N_7873);
nor U8905 (N_8905,N_7412,N_7757);
xnor U8906 (N_8906,N_7650,N_7708);
and U8907 (N_8907,N_7146,N_7299);
and U8908 (N_8908,N_7301,N_7564);
xor U8909 (N_8909,N_7833,N_7646);
and U8910 (N_8910,N_7036,N_7213);
nand U8911 (N_8911,N_7551,N_7928);
and U8912 (N_8912,N_7025,N_7982);
xnor U8913 (N_8913,N_7076,N_7293);
and U8914 (N_8914,N_7055,N_7951);
nand U8915 (N_8915,N_7318,N_7826);
nor U8916 (N_8916,N_7526,N_7747);
nand U8917 (N_8917,N_7798,N_7648);
and U8918 (N_8918,N_7948,N_7111);
and U8919 (N_8919,N_7821,N_7901);
nand U8920 (N_8920,N_7915,N_7077);
or U8921 (N_8921,N_7790,N_7157);
xor U8922 (N_8922,N_7768,N_7383);
and U8923 (N_8923,N_7791,N_7988);
nand U8924 (N_8924,N_7508,N_7766);
nand U8925 (N_8925,N_7036,N_7461);
or U8926 (N_8926,N_7057,N_7568);
nand U8927 (N_8927,N_7998,N_7334);
nand U8928 (N_8928,N_7784,N_7008);
and U8929 (N_8929,N_7262,N_7520);
nand U8930 (N_8930,N_7718,N_7135);
and U8931 (N_8931,N_7410,N_7324);
nand U8932 (N_8932,N_7420,N_7219);
nand U8933 (N_8933,N_7051,N_7855);
or U8934 (N_8934,N_7698,N_7363);
xor U8935 (N_8935,N_7586,N_7090);
xor U8936 (N_8936,N_7907,N_7170);
nand U8937 (N_8937,N_7881,N_7873);
nand U8938 (N_8938,N_7778,N_7348);
nand U8939 (N_8939,N_7890,N_7018);
or U8940 (N_8940,N_7918,N_7056);
xnor U8941 (N_8941,N_7253,N_7162);
nor U8942 (N_8942,N_7985,N_7155);
nor U8943 (N_8943,N_7668,N_7199);
and U8944 (N_8944,N_7039,N_7574);
nand U8945 (N_8945,N_7579,N_7537);
and U8946 (N_8946,N_7179,N_7200);
xnor U8947 (N_8947,N_7521,N_7517);
and U8948 (N_8948,N_7751,N_7289);
and U8949 (N_8949,N_7968,N_7341);
and U8950 (N_8950,N_7728,N_7292);
and U8951 (N_8951,N_7801,N_7531);
nand U8952 (N_8952,N_7634,N_7129);
xor U8953 (N_8953,N_7550,N_7842);
nand U8954 (N_8954,N_7961,N_7883);
xor U8955 (N_8955,N_7211,N_7724);
nand U8956 (N_8956,N_7510,N_7589);
nor U8957 (N_8957,N_7705,N_7455);
nor U8958 (N_8958,N_7148,N_7610);
or U8959 (N_8959,N_7303,N_7724);
and U8960 (N_8960,N_7243,N_7083);
or U8961 (N_8961,N_7307,N_7780);
nand U8962 (N_8962,N_7014,N_7597);
nand U8963 (N_8963,N_7567,N_7238);
xnor U8964 (N_8964,N_7763,N_7111);
nor U8965 (N_8965,N_7362,N_7976);
or U8966 (N_8966,N_7521,N_7316);
nand U8967 (N_8967,N_7925,N_7788);
nor U8968 (N_8968,N_7250,N_7562);
xnor U8969 (N_8969,N_7684,N_7801);
and U8970 (N_8970,N_7887,N_7413);
xnor U8971 (N_8971,N_7142,N_7738);
or U8972 (N_8972,N_7694,N_7177);
and U8973 (N_8973,N_7379,N_7062);
nand U8974 (N_8974,N_7321,N_7214);
xor U8975 (N_8975,N_7245,N_7688);
nand U8976 (N_8976,N_7891,N_7092);
or U8977 (N_8977,N_7837,N_7034);
or U8978 (N_8978,N_7352,N_7223);
nor U8979 (N_8979,N_7030,N_7858);
nand U8980 (N_8980,N_7526,N_7852);
and U8981 (N_8981,N_7196,N_7124);
nor U8982 (N_8982,N_7136,N_7246);
or U8983 (N_8983,N_7990,N_7558);
or U8984 (N_8984,N_7979,N_7202);
xnor U8985 (N_8985,N_7092,N_7342);
xor U8986 (N_8986,N_7829,N_7434);
xnor U8987 (N_8987,N_7331,N_7738);
nor U8988 (N_8988,N_7516,N_7616);
xnor U8989 (N_8989,N_7168,N_7040);
or U8990 (N_8990,N_7693,N_7417);
xor U8991 (N_8991,N_7198,N_7459);
xor U8992 (N_8992,N_7839,N_7943);
nand U8993 (N_8993,N_7063,N_7717);
and U8994 (N_8994,N_7983,N_7473);
and U8995 (N_8995,N_7417,N_7798);
nand U8996 (N_8996,N_7365,N_7963);
nand U8997 (N_8997,N_7947,N_7896);
xnor U8998 (N_8998,N_7357,N_7862);
xnor U8999 (N_8999,N_7771,N_7614);
or U9000 (N_9000,N_8210,N_8469);
and U9001 (N_9001,N_8723,N_8604);
or U9002 (N_9002,N_8146,N_8700);
or U9003 (N_9003,N_8853,N_8292);
nor U9004 (N_9004,N_8257,N_8219);
xor U9005 (N_9005,N_8211,N_8589);
xnor U9006 (N_9006,N_8784,N_8035);
and U9007 (N_9007,N_8578,N_8092);
or U9008 (N_9008,N_8980,N_8125);
xor U9009 (N_9009,N_8037,N_8098);
and U9010 (N_9010,N_8790,N_8242);
and U9011 (N_9011,N_8188,N_8820);
nand U9012 (N_9012,N_8278,N_8975);
nand U9013 (N_9013,N_8521,N_8648);
and U9014 (N_9014,N_8132,N_8281);
or U9015 (N_9015,N_8566,N_8195);
xnor U9016 (N_9016,N_8361,N_8798);
xor U9017 (N_9017,N_8499,N_8434);
and U9018 (N_9018,N_8363,N_8465);
nor U9019 (N_9019,N_8246,N_8355);
or U9020 (N_9020,N_8071,N_8576);
and U9021 (N_9021,N_8942,N_8580);
nand U9022 (N_9022,N_8957,N_8719);
or U9023 (N_9023,N_8844,N_8796);
nand U9024 (N_9024,N_8238,N_8344);
and U9025 (N_9025,N_8059,N_8922);
and U9026 (N_9026,N_8476,N_8187);
and U9027 (N_9027,N_8228,N_8792);
or U9028 (N_9028,N_8209,N_8058);
and U9029 (N_9029,N_8207,N_8738);
nor U9030 (N_9030,N_8430,N_8946);
and U9031 (N_9031,N_8764,N_8452);
nor U9032 (N_9032,N_8901,N_8658);
or U9033 (N_9033,N_8845,N_8777);
and U9034 (N_9034,N_8220,N_8688);
and U9035 (N_9035,N_8105,N_8787);
and U9036 (N_9036,N_8695,N_8339);
xor U9037 (N_9037,N_8051,N_8742);
nor U9038 (N_9038,N_8221,N_8159);
xnor U9039 (N_9039,N_8919,N_8786);
or U9040 (N_9040,N_8822,N_8256);
and U9041 (N_9041,N_8028,N_8879);
nor U9042 (N_9042,N_8735,N_8460);
nand U9043 (N_9043,N_8495,N_8655);
nor U9044 (N_9044,N_8108,N_8538);
nor U9045 (N_9045,N_8873,N_8736);
nand U9046 (N_9046,N_8231,N_8439);
xor U9047 (N_9047,N_8009,N_8643);
xnor U9048 (N_9048,N_8124,N_8849);
nor U9049 (N_9049,N_8630,N_8485);
or U9050 (N_9050,N_8198,N_8064);
nor U9051 (N_9051,N_8008,N_8878);
xor U9052 (N_9052,N_8110,N_8842);
and U9053 (N_9053,N_8733,N_8940);
nor U9054 (N_9054,N_8459,N_8584);
nand U9055 (N_9055,N_8837,N_8240);
nand U9056 (N_9056,N_8480,N_8772);
nand U9057 (N_9057,N_8974,N_8606);
and U9058 (N_9058,N_8097,N_8793);
xnor U9059 (N_9059,N_8675,N_8809);
and U9060 (N_9060,N_8299,N_8954);
xnor U9061 (N_9061,N_8520,N_8970);
nand U9062 (N_9062,N_8565,N_8237);
nor U9063 (N_9063,N_8399,N_8794);
xor U9064 (N_9064,N_8501,N_8621);
or U9065 (N_9065,N_8366,N_8341);
or U9066 (N_9066,N_8571,N_8867);
nand U9067 (N_9067,N_8596,N_8270);
xor U9068 (N_9068,N_8425,N_8511);
xor U9069 (N_9069,N_8271,N_8681);
nand U9070 (N_9070,N_8711,N_8085);
nor U9071 (N_9071,N_8585,N_8561);
nor U9072 (N_9072,N_8697,N_8552);
nand U9073 (N_9073,N_8212,N_8562);
xor U9074 (N_9074,N_8770,N_8079);
or U9075 (N_9075,N_8614,N_8456);
nand U9076 (N_9076,N_8704,N_8007);
and U9077 (N_9077,N_8996,N_8951);
or U9078 (N_9078,N_8194,N_8300);
or U9079 (N_9079,N_8682,N_8966);
nor U9080 (N_9080,N_8789,N_8056);
nand U9081 (N_9081,N_8583,N_8810);
xor U9082 (N_9082,N_8141,N_8807);
xor U9083 (N_9083,N_8156,N_8239);
or U9084 (N_9084,N_8023,N_8507);
and U9085 (N_9085,N_8780,N_8717);
nor U9086 (N_9086,N_8702,N_8165);
or U9087 (N_9087,N_8289,N_8619);
nand U9088 (N_9088,N_8597,N_8889);
or U9089 (N_9089,N_8450,N_8973);
nor U9090 (N_9090,N_8687,N_8959);
nand U9091 (N_9091,N_8884,N_8369);
or U9092 (N_9092,N_8080,N_8123);
nand U9093 (N_9093,N_8864,N_8752);
nand U9094 (N_9094,N_8855,N_8699);
nand U9095 (N_9095,N_8865,N_8145);
xnor U9096 (N_9096,N_8761,N_8749);
or U9097 (N_9097,N_8164,N_8517);
nor U9098 (N_9098,N_8380,N_8320);
nand U9099 (N_9099,N_8273,N_8985);
nand U9100 (N_9100,N_8312,N_8082);
and U9101 (N_9101,N_8535,N_8850);
xor U9102 (N_9102,N_8118,N_8177);
nand U9103 (N_9103,N_8947,N_8559);
xnor U9104 (N_9104,N_8757,N_8374);
nor U9105 (N_9105,N_8902,N_8229);
or U9106 (N_9106,N_8261,N_8781);
and U9107 (N_9107,N_8275,N_8731);
and U9108 (N_9108,N_8714,N_8721);
or U9109 (N_9109,N_8414,N_8342);
and U9110 (N_9110,N_8963,N_8838);
nand U9111 (N_9111,N_8431,N_8055);
xor U9112 (N_9112,N_8030,N_8831);
xor U9113 (N_9113,N_8815,N_8642);
or U9114 (N_9114,N_8052,N_8436);
xnor U9115 (N_9115,N_8692,N_8326);
nand U9116 (N_9116,N_8601,N_8100);
nand U9117 (N_9117,N_8564,N_8607);
nand U9118 (N_9118,N_8244,N_8277);
and U9119 (N_9119,N_8771,N_8746);
nand U9120 (N_9120,N_8078,N_8316);
nor U9121 (N_9121,N_8814,N_8147);
xnor U9122 (N_9122,N_8819,N_8824);
xor U9123 (N_9123,N_8540,N_8068);
or U9124 (N_9124,N_8451,N_8612);
xor U9125 (N_9125,N_8259,N_8722);
xnor U9126 (N_9126,N_8650,N_8926);
nand U9127 (N_9127,N_8785,N_8429);
xor U9128 (N_9128,N_8408,N_8512);
or U9129 (N_9129,N_8783,N_8302);
nand U9130 (N_9130,N_8915,N_8218);
or U9131 (N_9131,N_8148,N_8545);
nor U9132 (N_9132,N_8489,N_8575);
or U9133 (N_9133,N_8018,N_8245);
or U9134 (N_9134,N_8544,N_8943);
nand U9135 (N_9135,N_8063,N_8860);
nor U9136 (N_9136,N_8006,N_8911);
or U9137 (N_9137,N_8154,N_8801);
nand U9138 (N_9138,N_8338,N_8936);
or U9139 (N_9139,N_8336,N_8728);
nand U9140 (N_9140,N_8554,N_8641);
nand U9141 (N_9141,N_8720,N_8982);
and U9142 (N_9142,N_8362,N_8400);
or U9143 (N_9143,N_8625,N_8269);
xor U9144 (N_9144,N_8811,N_8712);
nor U9145 (N_9145,N_8492,N_8223);
and U9146 (N_9146,N_8284,N_8365);
and U9147 (N_9147,N_8350,N_8703);
or U9148 (N_9148,N_8532,N_8441);
or U9149 (N_9149,N_8230,N_8135);
nor U9150 (N_9150,N_8823,N_8698);
nor U9151 (N_9151,N_8043,N_8547);
and U9152 (N_9152,N_8529,N_8689);
or U9153 (N_9153,N_8002,N_8137);
nor U9154 (N_9154,N_8000,N_8183);
nand U9155 (N_9155,N_8560,N_8376);
xor U9156 (N_9156,N_8993,N_8073);
xor U9157 (N_9157,N_8635,N_8295);
or U9158 (N_9158,N_8402,N_8170);
and U9159 (N_9159,N_8310,N_8314);
nor U9160 (N_9160,N_8727,N_8760);
and U9161 (N_9161,N_8778,N_8461);
and U9162 (N_9162,N_8907,N_8404);
nand U9163 (N_9163,N_8906,N_8570);
and U9164 (N_9164,N_8286,N_8482);
nor U9165 (N_9165,N_8611,N_8249);
and U9166 (N_9166,N_8426,N_8550);
nand U9167 (N_9167,N_8972,N_8042);
xor U9168 (N_9168,N_8303,N_8328);
and U9169 (N_9169,N_8679,N_8033);
nor U9170 (N_9170,N_8917,N_8836);
nor U9171 (N_9171,N_8318,N_8638);
nor U9172 (N_9172,N_8739,N_8861);
and U9173 (N_9173,N_8029,N_8537);
or U9174 (N_9174,N_8962,N_8881);
xor U9175 (N_9175,N_8397,N_8225);
xnor U9176 (N_9176,N_8890,N_8317);
or U9177 (N_9177,N_8967,N_8074);
or U9178 (N_9178,N_8885,N_8826);
nor U9179 (N_9179,N_8984,N_8081);
nand U9180 (N_9180,N_8817,N_8367);
and U9181 (N_9181,N_8031,N_8255);
nor U9182 (N_9182,N_8252,N_8877);
xnor U9183 (N_9183,N_8563,N_8644);
xor U9184 (N_9184,N_8140,N_8931);
and U9185 (N_9185,N_8613,N_8045);
nor U9186 (N_9186,N_8453,N_8224);
nor U9187 (N_9187,N_8396,N_8676);
or U9188 (N_9188,N_8047,N_8519);
nand U9189 (N_9189,N_8473,N_8927);
nand U9190 (N_9190,N_8041,N_8715);
nor U9191 (N_9191,N_8184,N_8484);
nor U9192 (N_9192,N_8395,N_8191);
nor U9193 (N_9193,N_8851,N_8568);
xor U9194 (N_9194,N_8965,N_8083);
nor U9195 (N_9195,N_8010,N_8910);
nand U9196 (N_9196,N_8513,N_8623);
nand U9197 (N_9197,N_8754,N_8114);
nand U9198 (N_9198,N_8263,N_8274);
nor U9199 (N_9199,N_8038,N_8151);
xnor U9200 (N_9200,N_8744,N_8173);
and U9201 (N_9201,N_8933,N_8542);
and U9202 (N_9202,N_8490,N_8593);
and U9203 (N_9203,N_8581,N_8574);
and U9204 (N_9204,N_8454,N_8639);
xnor U9205 (N_9205,N_8048,N_8032);
or U9206 (N_9206,N_8181,N_8179);
nand U9207 (N_9207,N_8264,N_8072);
xor U9208 (N_9208,N_8516,N_8149);
xor U9209 (N_9209,N_8693,N_8634);
and U9210 (N_9210,N_8444,N_8375);
and U9211 (N_9211,N_8357,N_8446);
or U9212 (N_9212,N_8653,N_8335);
and U9213 (N_9213,N_8440,N_8088);
nor U9214 (N_9214,N_8398,N_8918);
and U9215 (N_9215,N_8267,N_8325);
xnor U9216 (N_9216,N_8351,N_8153);
nand U9217 (N_9217,N_8816,N_8981);
xor U9218 (N_9218,N_8020,N_8729);
and U9219 (N_9219,N_8157,N_8629);
nand U9220 (N_9220,N_8497,N_8882);
nand U9221 (N_9221,N_8769,N_8724);
nand U9222 (N_9222,N_8379,N_8600);
nand U9223 (N_9223,N_8961,N_8858);
xnor U9224 (N_9224,N_8678,N_8812);
xor U9225 (N_9225,N_8458,N_8285);
xnor U9226 (N_9226,N_8017,N_8825);
nand U9227 (N_9227,N_8869,N_8791);
nor U9228 (N_9228,N_8603,N_8701);
nor U9229 (N_9229,N_8233,N_8661);
nand U9230 (N_9230,N_8691,N_8830);
or U9231 (N_9231,N_8232,N_8654);
xnor U9232 (N_9232,N_8610,N_8775);
xnor U9233 (N_9233,N_8382,N_8841);
nand U9234 (N_9234,N_8373,N_8839);
nand U9235 (N_9235,N_8352,N_8553);
nor U9236 (N_9236,N_8543,N_8416);
and U9237 (N_9237,N_8340,N_8011);
or U9238 (N_9238,N_8437,N_8279);
xor U9239 (N_9239,N_8671,N_8204);
and U9240 (N_9240,N_8403,N_8205);
or U9241 (N_9241,N_8174,N_8734);
xor U9242 (N_9242,N_8636,N_8445);
xnor U9243 (N_9243,N_8549,N_8854);
or U9244 (N_9244,N_8832,N_8863);
nand U9245 (N_9245,N_8948,N_8628);
nand U9246 (N_9246,N_8572,N_8903);
xnor U9247 (N_9247,N_8526,N_8912);
nor U9248 (N_9248,N_8364,N_8093);
or U9249 (N_9249,N_8664,N_8514);
nor U9250 (N_9250,N_8925,N_8143);
nand U9251 (N_9251,N_8806,N_8457);
and U9252 (N_9252,N_8523,N_8062);
or U9253 (N_9253,N_8905,N_8419);
nor U9254 (N_9254,N_8828,N_8637);
or U9255 (N_9255,N_8478,N_8496);
and U9256 (N_9256,N_8986,N_8904);
nand U9257 (N_9257,N_8803,N_8958);
and U9258 (N_9258,N_8356,N_8272);
nand U9259 (N_9259,N_8932,N_8094);
nand U9260 (N_9260,N_8133,N_8260);
xor U9261 (N_9261,N_8737,N_8420);
or U9262 (N_9262,N_8747,N_8095);
xnor U9263 (N_9263,N_8150,N_8608);
and U9264 (N_9264,N_8856,N_8012);
or U9265 (N_9265,N_8805,N_8646);
and U9266 (N_9266,N_8886,N_8117);
nor U9267 (N_9267,N_8106,N_8944);
nand U9268 (N_9268,N_8663,N_8305);
or U9269 (N_9269,N_8716,N_8280);
nand U9270 (N_9270,N_8337,N_8569);
nand U9271 (N_9271,N_8536,N_8616);
nor U9272 (N_9272,N_8534,N_8577);
xnor U9273 (N_9273,N_8502,N_8586);
and U9274 (N_9274,N_8776,N_8428);
xor U9275 (N_9275,N_8852,N_8500);
and U9276 (N_9276,N_8309,N_8527);
xor U9277 (N_9277,N_8180,N_8371);
nand U9278 (N_9278,N_8347,N_8955);
nand U9279 (N_9279,N_8950,N_8102);
and U9280 (N_9280,N_8290,N_8683);
nand U9281 (N_9281,N_8992,N_8053);
nand U9282 (N_9282,N_8065,N_8657);
nand U9283 (N_9283,N_8163,N_8107);
or U9284 (N_9284,N_8160,N_8243);
xor U9285 (N_9285,N_8740,N_8732);
and U9286 (N_9286,N_8196,N_8504);
nand U9287 (N_9287,N_8176,N_8713);
nor U9288 (N_9288,N_8136,N_8378);
or U9289 (N_9289,N_8413,N_8401);
xor U9290 (N_9290,N_8090,N_8880);
xor U9291 (N_9291,N_8509,N_8468);
nor U9292 (N_9292,N_8186,N_8266);
nor U9293 (N_9293,N_8169,N_8096);
and U9294 (N_9294,N_8421,N_8498);
nor U9295 (N_9295,N_8202,N_8923);
and U9296 (N_9296,N_8888,N_8518);
and U9297 (N_9297,N_8493,N_8372);
and U9298 (N_9298,N_8329,N_8144);
or U9299 (N_9299,N_8390,N_8598);
nor U9300 (N_9300,N_8892,N_8175);
nor U9301 (N_9301,N_8026,N_8087);
nand U9302 (N_9302,N_8743,N_8192);
nor U9303 (N_9303,N_8674,N_8387);
or U9304 (N_9304,N_8346,N_8591);
and U9305 (N_9305,N_8185,N_8934);
xnor U9306 (N_9306,N_8914,N_8127);
nand U9307 (N_9307,N_8077,N_8443);
or U9308 (N_9308,N_8427,N_8381);
and U9309 (N_9309,N_8620,N_8158);
and U9310 (N_9310,N_8573,N_8034);
or U9311 (N_9311,N_8193,N_8875);
xor U9312 (N_9312,N_8442,N_8594);
nand U9313 (N_9313,N_8515,N_8883);
or U9314 (N_9314,N_8475,N_8234);
or U9315 (N_9315,N_8938,N_8990);
or U9316 (N_9316,N_8359,N_8510);
nor U9317 (N_9317,N_8960,N_8908);
xnor U9318 (N_9318,N_8206,N_8168);
or U9319 (N_9319,N_8306,N_8227);
nor U9320 (N_9320,N_8659,N_8748);
xor U9321 (N_9321,N_8615,N_8236);
nand U9322 (N_9322,N_8119,N_8684);
nand U9323 (N_9323,N_8935,N_8991);
xor U9324 (N_9324,N_8321,N_8921);
nor U9325 (N_9325,N_8779,N_8296);
nand U9326 (N_9326,N_8131,N_8040);
or U9327 (N_9327,N_8353,N_8293);
nand U9328 (N_9328,N_8166,N_8322);
nor U9329 (N_9329,N_8319,N_8672);
xor U9330 (N_9330,N_8546,N_8874);
xnor U9331 (N_9331,N_8800,N_8308);
nor U9332 (N_9332,N_8235,N_8756);
and U9333 (N_9333,N_8969,N_8152);
or U9334 (N_9334,N_8287,N_8622);
xnor U9335 (N_9335,N_8751,N_8848);
nor U9336 (N_9336,N_8019,N_8755);
nand U9337 (N_9337,N_8021,N_8411);
nor U9338 (N_9338,N_8887,N_8708);
xnor U9339 (N_9339,N_8182,N_8197);
nand U9340 (N_9340,N_8360,N_8802);
nor U9341 (N_9341,N_8226,N_8897);
and U9342 (N_9342,N_8968,N_8670);
nor U9343 (N_9343,N_8348,N_8945);
xor U9344 (N_9344,N_8005,N_8409);
nor U9345 (N_9345,N_8994,N_8334);
nand U9346 (N_9346,N_8455,N_8758);
nor U9347 (N_9347,N_8104,N_8291);
nand U9348 (N_9348,N_8645,N_8753);
xor U9349 (N_9349,N_8307,N_8330);
or U9350 (N_9350,N_8189,N_8588);
or U9351 (N_9351,N_8774,N_8999);
nor U9352 (N_9352,N_8036,N_8412);
or U9353 (N_9353,N_8016,N_8354);
or U9354 (N_9354,N_8432,N_8894);
and U9355 (N_9355,N_8632,N_8686);
nor U9356 (N_9356,N_8463,N_8989);
or U9357 (N_9357,N_8385,N_8909);
and U9358 (N_9358,N_8384,N_8506);
or U9359 (N_9359,N_8422,N_8386);
nand U9360 (N_9360,N_8987,N_8530);
nor U9361 (N_9361,N_8988,N_8015);
and U9362 (N_9362,N_8258,N_8759);
nor U9363 (N_9363,N_8685,N_8111);
and U9364 (N_9364,N_8673,N_8470);
or U9365 (N_9365,N_8750,N_8139);
and U9366 (N_9366,N_8827,N_8767);
or U9367 (N_9367,N_8998,N_8649);
and U9368 (N_9368,N_8406,N_8392);
xnor U9369 (N_9369,N_8762,N_8924);
nand U9370 (N_9370,N_8254,N_8370);
nand U9371 (N_9371,N_8115,N_8358);
or U9372 (N_9372,N_8126,N_8069);
nand U9373 (N_9373,N_8423,N_8155);
or U9374 (N_9374,N_8528,N_8389);
and U9375 (N_9375,N_8626,N_8706);
and U9376 (N_9376,N_8294,N_8555);
nor U9377 (N_9377,N_8208,N_8680);
nor U9378 (N_9378,N_8592,N_8248);
xnor U9379 (N_9379,N_8788,N_8640);
and U9380 (N_9380,N_8595,N_8101);
and U9381 (N_9381,N_8808,N_8718);
xor U9382 (N_9382,N_8134,N_8061);
nand U9383 (N_9383,N_8847,N_8324);
nand U9384 (N_9384,N_8870,N_8677);
xor U9385 (N_9385,N_8447,N_8567);
and U9386 (N_9386,N_8505,N_8773);
and U9387 (N_9387,N_8696,N_8618);
or U9388 (N_9388,N_8862,N_8690);
nand U9389 (N_9389,N_8871,N_8178);
nand U9390 (N_9390,N_8025,N_8941);
nor U9391 (N_9391,N_8913,N_8474);
xnor U9392 (N_9392,N_8027,N_8405);
xor U9393 (N_9393,N_8730,N_8129);
xnor U9394 (N_9394,N_8726,N_8813);
xnor U9395 (N_9395,N_8524,N_8297);
or U9396 (N_9396,N_8647,N_8548);
nor U9397 (N_9397,N_8768,N_8253);
or U9398 (N_9398,N_8896,N_8304);
nand U9399 (N_9399,N_8332,N_8930);
xor U9400 (N_9400,N_8741,N_8044);
and U9401 (N_9401,N_8582,N_8167);
nand U9402 (N_9402,N_8843,N_8368);
nand U9403 (N_9403,N_8669,N_8213);
and U9404 (N_9404,N_8956,N_8250);
and U9405 (N_9405,N_8418,N_8001);
or U9406 (N_9406,N_8605,N_8834);
nand U9407 (N_9407,N_8609,N_8121);
and U9408 (N_9408,N_8745,N_8109);
nand U9409 (N_9409,N_8433,N_8709);
xor U9410 (N_9410,N_8556,N_8013);
xor U9411 (N_9411,N_8086,N_8138);
nor U9412 (N_9412,N_8503,N_8471);
and U9413 (N_9413,N_8804,N_8763);
or U9414 (N_9414,N_8066,N_8891);
xnor U9415 (N_9415,N_8142,N_8200);
and U9416 (N_9416,N_8694,N_8089);
xnor U9417 (N_9417,N_8953,N_8551);
and U9418 (N_9418,N_8070,N_8276);
nor U9419 (N_9419,N_8103,N_8262);
or U9420 (N_9420,N_8391,N_8665);
xor U9421 (N_9421,N_8162,N_8539);
and U9422 (N_9422,N_8898,N_8216);
nand U9423 (N_9423,N_8039,N_8487);
xor U9424 (N_9424,N_8383,N_8464);
xor U9425 (N_9425,N_8315,N_8631);
nor U9426 (N_9426,N_8203,N_8172);
nand U9427 (N_9427,N_8531,N_8199);
or U9428 (N_9428,N_8014,N_8099);
and U9429 (N_9429,N_8003,N_8483);
nor U9430 (N_9430,N_8004,N_8161);
and U9431 (N_9431,N_8113,N_8668);
and U9432 (N_9432,N_8821,N_8928);
and U9433 (N_9433,N_8876,N_8964);
and U9434 (N_9434,N_8394,N_8313);
nor U9435 (N_9435,N_8920,N_8449);
xor U9436 (N_9436,N_8846,N_8084);
nor U9437 (N_9437,N_8868,N_8301);
nor U9438 (N_9438,N_8481,N_8590);
nor U9439 (N_9439,N_8054,N_8417);
nor U9440 (N_9440,N_8331,N_8949);
nand U9441 (N_9441,N_8283,N_8190);
nand U9442 (N_9442,N_8599,N_8494);
and U9443 (N_9443,N_8265,N_8333);
xnor U9444 (N_9444,N_8617,N_8525);
nand U9445 (N_9445,N_8491,N_8782);
nor U9446 (N_9446,N_8895,N_8508);
nand U9447 (N_9447,N_8122,N_8766);
and U9448 (N_9448,N_8268,N_8076);
xor U9449 (N_9449,N_8438,N_8977);
xnor U9450 (N_9450,N_8247,N_8835);
or U9451 (N_9451,N_8049,N_8979);
nand U9452 (N_9452,N_8091,N_8660);
nand U9453 (N_9453,N_8112,N_8833);
and U9454 (N_9454,N_8799,N_8651);
and U9455 (N_9455,N_8050,N_8024);
and U9456 (N_9456,N_8857,N_8349);
nand U9457 (N_9457,N_8067,N_8214);
xor U9458 (N_9458,N_8710,N_8311);
nor U9459 (N_9459,N_8075,N_8840);
or U9460 (N_9460,N_8667,N_8899);
and U9461 (N_9461,N_8707,N_8558);
nand U9462 (N_9462,N_8633,N_8345);
or U9463 (N_9463,N_8997,N_8116);
xor U9464 (N_9464,N_8288,N_8533);
nor U9465 (N_9465,N_8624,N_8388);
xnor U9466 (N_9466,N_8477,N_8217);
nor U9467 (N_9467,N_8557,N_8215);
nand U9468 (N_9468,N_8893,N_8488);
xnor U9469 (N_9469,N_8795,N_8602);
or U9470 (N_9470,N_8022,N_8393);
or U9471 (N_9471,N_8128,N_8929);
and U9472 (N_9472,N_8201,N_8424);
or U9473 (N_9473,N_8462,N_8120);
nor U9474 (N_9474,N_8479,N_8343);
xnor U9475 (N_9475,N_8797,N_8976);
xnor U9476 (N_9476,N_8866,N_8448);
xnor U9477 (N_9477,N_8327,N_8377);
nand U9478 (N_9478,N_8046,N_8579);
nand U9479 (N_9479,N_8725,N_8995);
nand U9480 (N_9480,N_8765,N_8939);
xor U9481 (N_9481,N_8916,N_8818);
xor U9482 (N_9482,N_8829,N_8057);
or U9483 (N_9483,N_8171,N_8060);
nor U9484 (N_9484,N_8407,N_8222);
nor U9485 (N_9485,N_8435,N_8472);
and U9486 (N_9486,N_8282,N_8662);
nand U9487 (N_9487,N_8971,N_8652);
and U9488 (N_9488,N_8522,N_8541);
xnor U9489 (N_9489,N_8467,N_8466);
xnor U9490 (N_9490,N_8587,N_8900);
or U9491 (N_9491,N_8298,N_8323);
nand U9492 (N_9492,N_8241,N_8656);
or U9493 (N_9493,N_8415,N_8627);
nand U9494 (N_9494,N_8952,N_8983);
xor U9495 (N_9495,N_8872,N_8705);
nand U9496 (N_9496,N_8410,N_8978);
or U9497 (N_9497,N_8130,N_8937);
nand U9498 (N_9498,N_8666,N_8859);
nor U9499 (N_9499,N_8251,N_8486);
nand U9500 (N_9500,N_8747,N_8833);
nor U9501 (N_9501,N_8167,N_8726);
and U9502 (N_9502,N_8085,N_8729);
nor U9503 (N_9503,N_8796,N_8163);
or U9504 (N_9504,N_8098,N_8594);
or U9505 (N_9505,N_8143,N_8801);
nand U9506 (N_9506,N_8706,N_8083);
nand U9507 (N_9507,N_8813,N_8255);
and U9508 (N_9508,N_8361,N_8204);
xnor U9509 (N_9509,N_8949,N_8399);
nor U9510 (N_9510,N_8611,N_8051);
and U9511 (N_9511,N_8088,N_8480);
nor U9512 (N_9512,N_8427,N_8347);
or U9513 (N_9513,N_8723,N_8111);
or U9514 (N_9514,N_8352,N_8318);
xor U9515 (N_9515,N_8097,N_8618);
xor U9516 (N_9516,N_8119,N_8973);
nor U9517 (N_9517,N_8680,N_8594);
or U9518 (N_9518,N_8598,N_8790);
and U9519 (N_9519,N_8943,N_8885);
nand U9520 (N_9520,N_8178,N_8293);
or U9521 (N_9521,N_8696,N_8008);
or U9522 (N_9522,N_8682,N_8466);
or U9523 (N_9523,N_8543,N_8691);
xnor U9524 (N_9524,N_8670,N_8790);
or U9525 (N_9525,N_8606,N_8510);
and U9526 (N_9526,N_8009,N_8337);
or U9527 (N_9527,N_8334,N_8391);
or U9528 (N_9528,N_8532,N_8948);
or U9529 (N_9529,N_8529,N_8034);
or U9530 (N_9530,N_8276,N_8647);
xor U9531 (N_9531,N_8275,N_8956);
or U9532 (N_9532,N_8833,N_8735);
nand U9533 (N_9533,N_8520,N_8530);
or U9534 (N_9534,N_8941,N_8288);
xor U9535 (N_9535,N_8854,N_8036);
nor U9536 (N_9536,N_8103,N_8397);
or U9537 (N_9537,N_8319,N_8381);
nand U9538 (N_9538,N_8402,N_8871);
nor U9539 (N_9539,N_8964,N_8793);
xor U9540 (N_9540,N_8344,N_8660);
and U9541 (N_9541,N_8761,N_8101);
xnor U9542 (N_9542,N_8376,N_8172);
xnor U9543 (N_9543,N_8186,N_8820);
nand U9544 (N_9544,N_8382,N_8032);
or U9545 (N_9545,N_8317,N_8808);
or U9546 (N_9546,N_8322,N_8043);
nand U9547 (N_9547,N_8052,N_8502);
and U9548 (N_9548,N_8686,N_8456);
or U9549 (N_9549,N_8459,N_8206);
and U9550 (N_9550,N_8846,N_8220);
nand U9551 (N_9551,N_8617,N_8846);
and U9552 (N_9552,N_8718,N_8360);
nand U9553 (N_9553,N_8593,N_8550);
xor U9554 (N_9554,N_8996,N_8301);
nand U9555 (N_9555,N_8181,N_8050);
xnor U9556 (N_9556,N_8607,N_8137);
nand U9557 (N_9557,N_8581,N_8812);
xnor U9558 (N_9558,N_8463,N_8636);
nor U9559 (N_9559,N_8403,N_8814);
nor U9560 (N_9560,N_8551,N_8582);
and U9561 (N_9561,N_8237,N_8178);
or U9562 (N_9562,N_8783,N_8697);
nor U9563 (N_9563,N_8493,N_8996);
nor U9564 (N_9564,N_8873,N_8151);
nor U9565 (N_9565,N_8864,N_8485);
nor U9566 (N_9566,N_8484,N_8209);
nor U9567 (N_9567,N_8792,N_8105);
nor U9568 (N_9568,N_8250,N_8825);
or U9569 (N_9569,N_8104,N_8804);
nand U9570 (N_9570,N_8257,N_8914);
nand U9571 (N_9571,N_8467,N_8474);
nor U9572 (N_9572,N_8935,N_8040);
nor U9573 (N_9573,N_8906,N_8730);
and U9574 (N_9574,N_8781,N_8466);
nand U9575 (N_9575,N_8458,N_8844);
xnor U9576 (N_9576,N_8599,N_8797);
xor U9577 (N_9577,N_8856,N_8730);
nor U9578 (N_9578,N_8045,N_8921);
and U9579 (N_9579,N_8157,N_8687);
or U9580 (N_9580,N_8520,N_8472);
xnor U9581 (N_9581,N_8424,N_8315);
or U9582 (N_9582,N_8814,N_8536);
and U9583 (N_9583,N_8624,N_8197);
and U9584 (N_9584,N_8064,N_8874);
xnor U9585 (N_9585,N_8647,N_8466);
nand U9586 (N_9586,N_8700,N_8637);
and U9587 (N_9587,N_8211,N_8968);
nand U9588 (N_9588,N_8888,N_8222);
and U9589 (N_9589,N_8621,N_8785);
and U9590 (N_9590,N_8158,N_8097);
nand U9591 (N_9591,N_8775,N_8743);
and U9592 (N_9592,N_8976,N_8372);
xnor U9593 (N_9593,N_8751,N_8386);
or U9594 (N_9594,N_8783,N_8207);
nor U9595 (N_9595,N_8938,N_8520);
xor U9596 (N_9596,N_8056,N_8768);
or U9597 (N_9597,N_8842,N_8278);
nand U9598 (N_9598,N_8995,N_8788);
nand U9599 (N_9599,N_8786,N_8692);
nand U9600 (N_9600,N_8437,N_8586);
or U9601 (N_9601,N_8149,N_8396);
nand U9602 (N_9602,N_8916,N_8283);
and U9603 (N_9603,N_8548,N_8429);
xnor U9604 (N_9604,N_8125,N_8166);
nor U9605 (N_9605,N_8593,N_8861);
and U9606 (N_9606,N_8503,N_8456);
or U9607 (N_9607,N_8089,N_8709);
nand U9608 (N_9608,N_8906,N_8001);
and U9609 (N_9609,N_8381,N_8436);
nand U9610 (N_9610,N_8832,N_8028);
or U9611 (N_9611,N_8206,N_8101);
nor U9612 (N_9612,N_8311,N_8500);
xor U9613 (N_9613,N_8684,N_8614);
xnor U9614 (N_9614,N_8142,N_8094);
xnor U9615 (N_9615,N_8941,N_8144);
and U9616 (N_9616,N_8583,N_8648);
xnor U9617 (N_9617,N_8044,N_8854);
xor U9618 (N_9618,N_8512,N_8182);
or U9619 (N_9619,N_8765,N_8847);
nor U9620 (N_9620,N_8534,N_8569);
nand U9621 (N_9621,N_8063,N_8624);
xor U9622 (N_9622,N_8166,N_8788);
or U9623 (N_9623,N_8822,N_8148);
nor U9624 (N_9624,N_8623,N_8956);
and U9625 (N_9625,N_8851,N_8512);
and U9626 (N_9626,N_8563,N_8544);
or U9627 (N_9627,N_8249,N_8616);
xor U9628 (N_9628,N_8868,N_8309);
or U9629 (N_9629,N_8113,N_8924);
xor U9630 (N_9630,N_8645,N_8979);
xnor U9631 (N_9631,N_8976,N_8291);
or U9632 (N_9632,N_8550,N_8200);
xor U9633 (N_9633,N_8715,N_8741);
nand U9634 (N_9634,N_8453,N_8896);
and U9635 (N_9635,N_8288,N_8472);
xnor U9636 (N_9636,N_8678,N_8190);
nand U9637 (N_9637,N_8778,N_8210);
nor U9638 (N_9638,N_8961,N_8719);
nand U9639 (N_9639,N_8138,N_8661);
nor U9640 (N_9640,N_8567,N_8357);
or U9641 (N_9641,N_8978,N_8599);
nor U9642 (N_9642,N_8326,N_8787);
or U9643 (N_9643,N_8389,N_8848);
or U9644 (N_9644,N_8035,N_8595);
xor U9645 (N_9645,N_8623,N_8212);
xor U9646 (N_9646,N_8966,N_8247);
nor U9647 (N_9647,N_8967,N_8795);
and U9648 (N_9648,N_8176,N_8234);
or U9649 (N_9649,N_8606,N_8180);
nand U9650 (N_9650,N_8809,N_8630);
and U9651 (N_9651,N_8629,N_8585);
or U9652 (N_9652,N_8872,N_8863);
and U9653 (N_9653,N_8304,N_8782);
and U9654 (N_9654,N_8045,N_8006);
or U9655 (N_9655,N_8933,N_8365);
xor U9656 (N_9656,N_8766,N_8986);
nor U9657 (N_9657,N_8320,N_8139);
or U9658 (N_9658,N_8412,N_8397);
xnor U9659 (N_9659,N_8166,N_8454);
xnor U9660 (N_9660,N_8874,N_8083);
xnor U9661 (N_9661,N_8926,N_8457);
or U9662 (N_9662,N_8652,N_8023);
nor U9663 (N_9663,N_8247,N_8260);
xor U9664 (N_9664,N_8915,N_8190);
nand U9665 (N_9665,N_8364,N_8107);
or U9666 (N_9666,N_8142,N_8998);
nand U9667 (N_9667,N_8912,N_8377);
or U9668 (N_9668,N_8731,N_8910);
nand U9669 (N_9669,N_8404,N_8050);
and U9670 (N_9670,N_8214,N_8046);
nor U9671 (N_9671,N_8854,N_8478);
nand U9672 (N_9672,N_8136,N_8015);
or U9673 (N_9673,N_8473,N_8685);
and U9674 (N_9674,N_8087,N_8540);
xor U9675 (N_9675,N_8524,N_8070);
or U9676 (N_9676,N_8635,N_8668);
nor U9677 (N_9677,N_8590,N_8675);
nand U9678 (N_9678,N_8730,N_8934);
nor U9679 (N_9679,N_8399,N_8418);
and U9680 (N_9680,N_8271,N_8086);
and U9681 (N_9681,N_8146,N_8207);
or U9682 (N_9682,N_8940,N_8260);
xor U9683 (N_9683,N_8893,N_8167);
and U9684 (N_9684,N_8624,N_8308);
nor U9685 (N_9685,N_8893,N_8274);
nand U9686 (N_9686,N_8003,N_8000);
or U9687 (N_9687,N_8826,N_8768);
xor U9688 (N_9688,N_8915,N_8374);
and U9689 (N_9689,N_8824,N_8542);
nand U9690 (N_9690,N_8574,N_8985);
nand U9691 (N_9691,N_8758,N_8042);
nand U9692 (N_9692,N_8608,N_8207);
or U9693 (N_9693,N_8847,N_8546);
nand U9694 (N_9694,N_8646,N_8967);
nand U9695 (N_9695,N_8929,N_8176);
or U9696 (N_9696,N_8275,N_8806);
and U9697 (N_9697,N_8363,N_8692);
nor U9698 (N_9698,N_8403,N_8555);
nand U9699 (N_9699,N_8809,N_8653);
and U9700 (N_9700,N_8883,N_8872);
nor U9701 (N_9701,N_8774,N_8595);
and U9702 (N_9702,N_8367,N_8090);
or U9703 (N_9703,N_8735,N_8983);
and U9704 (N_9704,N_8131,N_8968);
nor U9705 (N_9705,N_8987,N_8854);
and U9706 (N_9706,N_8910,N_8716);
nor U9707 (N_9707,N_8878,N_8662);
and U9708 (N_9708,N_8564,N_8346);
nand U9709 (N_9709,N_8378,N_8456);
nor U9710 (N_9710,N_8532,N_8177);
and U9711 (N_9711,N_8103,N_8842);
and U9712 (N_9712,N_8051,N_8157);
nand U9713 (N_9713,N_8401,N_8728);
and U9714 (N_9714,N_8463,N_8618);
and U9715 (N_9715,N_8117,N_8687);
nand U9716 (N_9716,N_8860,N_8145);
or U9717 (N_9717,N_8255,N_8872);
nand U9718 (N_9718,N_8722,N_8916);
or U9719 (N_9719,N_8514,N_8948);
nand U9720 (N_9720,N_8558,N_8074);
and U9721 (N_9721,N_8359,N_8276);
or U9722 (N_9722,N_8222,N_8121);
or U9723 (N_9723,N_8094,N_8529);
and U9724 (N_9724,N_8056,N_8665);
xor U9725 (N_9725,N_8934,N_8498);
nor U9726 (N_9726,N_8678,N_8067);
and U9727 (N_9727,N_8988,N_8187);
nor U9728 (N_9728,N_8696,N_8816);
nor U9729 (N_9729,N_8996,N_8900);
or U9730 (N_9730,N_8446,N_8825);
and U9731 (N_9731,N_8591,N_8173);
and U9732 (N_9732,N_8817,N_8751);
xor U9733 (N_9733,N_8416,N_8439);
nor U9734 (N_9734,N_8977,N_8942);
or U9735 (N_9735,N_8345,N_8201);
xor U9736 (N_9736,N_8642,N_8089);
and U9737 (N_9737,N_8181,N_8631);
xor U9738 (N_9738,N_8143,N_8808);
or U9739 (N_9739,N_8109,N_8142);
nor U9740 (N_9740,N_8223,N_8920);
nand U9741 (N_9741,N_8951,N_8676);
and U9742 (N_9742,N_8841,N_8343);
and U9743 (N_9743,N_8416,N_8945);
and U9744 (N_9744,N_8026,N_8530);
xor U9745 (N_9745,N_8938,N_8030);
nor U9746 (N_9746,N_8516,N_8183);
and U9747 (N_9747,N_8972,N_8663);
nor U9748 (N_9748,N_8887,N_8392);
or U9749 (N_9749,N_8392,N_8221);
xnor U9750 (N_9750,N_8625,N_8626);
and U9751 (N_9751,N_8376,N_8397);
nor U9752 (N_9752,N_8362,N_8474);
nor U9753 (N_9753,N_8003,N_8768);
or U9754 (N_9754,N_8432,N_8361);
xor U9755 (N_9755,N_8730,N_8252);
and U9756 (N_9756,N_8869,N_8334);
nand U9757 (N_9757,N_8710,N_8578);
or U9758 (N_9758,N_8393,N_8130);
or U9759 (N_9759,N_8165,N_8934);
xnor U9760 (N_9760,N_8606,N_8614);
nor U9761 (N_9761,N_8060,N_8803);
xor U9762 (N_9762,N_8188,N_8486);
xor U9763 (N_9763,N_8476,N_8921);
or U9764 (N_9764,N_8177,N_8450);
or U9765 (N_9765,N_8617,N_8072);
and U9766 (N_9766,N_8777,N_8717);
xor U9767 (N_9767,N_8498,N_8973);
nor U9768 (N_9768,N_8104,N_8800);
or U9769 (N_9769,N_8723,N_8993);
nor U9770 (N_9770,N_8229,N_8088);
and U9771 (N_9771,N_8218,N_8089);
nor U9772 (N_9772,N_8135,N_8142);
or U9773 (N_9773,N_8516,N_8971);
xor U9774 (N_9774,N_8278,N_8417);
nand U9775 (N_9775,N_8250,N_8261);
nand U9776 (N_9776,N_8830,N_8203);
nand U9777 (N_9777,N_8051,N_8636);
nor U9778 (N_9778,N_8502,N_8334);
nor U9779 (N_9779,N_8870,N_8609);
nor U9780 (N_9780,N_8336,N_8307);
nand U9781 (N_9781,N_8380,N_8792);
and U9782 (N_9782,N_8010,N_8020);
xor U9783 (N_9783,N_8044,N_8649);
xnor U9784 (N_9784,N_8324,N_8629);
xnor U9785 (N_9785,N_8102,N_8343);
and U9786 (N_9786,N_8613,N_8614);
and U9787 (N_9787,N_8162,N_8587);
xnor U9788 (N_9788,N_8005,N_8568);
and U9789 (N_9789,N_8830,N_8329);
or U9790 (N_9790,N_8193,N_8490);
and U9791 (N_9791,N_8180,N_8270);
and U9792 (N_9792,N_8875,N_8856);
nor U9793 (N_9793,N_8323,N_8158);
xnor U9794 (N_9794,N_8871,N_8955);
or U9795 (N_9795,N_8086,N_8238);
nor U9796 (N_9796,N_8970,N_8480);
nor U9797 (N_9797,N_8448,N_8974);
nand U9798 (N_9798,N_8685,N_8703);
and U9799 (N_9799,N_8981,N_8660);
xor U9800 (N_9800,N_8722,N_8933);
nor U9801 (N_9801,N_8675,N_8819);
and U9802 (N_9802,N_8411,N_8492);
nor U9803 (N_9803,N_8622,N_8184);
nand U9804 (N_9804,N_8429,N_8101);
and U9805 (N_9805,N_8172,N_8403);
and U9806 (N_9806,N_8728,N_8084);
and U9807 (N_9807,N_8439,N_8696);
and U9808 (N_9808,N_8252,N_8758);
nand U9809 (N_9809,N_8674,N_8971);
nand U9810 (N_9810,N_8554,N_8774);
nor U9811 (N_9811,N_8987,N_8087);
nand U9812 (N_9812,N_8090,N_8000);
nand U9813 (N_9813,N_8683,N_8986);
and U9814 (N_9814,N_8017,N_8926);
xnor U9815 (N_9815,N_8978,N_8989);
nor U9816 (N_9816,N_8689,N_8545);
xor U9817 (N_9817,N_8493,N_8415);
or U9818 (N_9818,N_8596,N_8859);
and U9819 (N_9819,N_8724,N_8335);
or U9820 (N_9820,N_8748,N_8370);
and U9821 (N_9821,N_8078,N_8525);
and U9822 (N_9822,N_8236,N_8261);
or U9823 (N_9823,N_8934,N_8405);
nand U9824 (N_9824,N_8383,N_8474);
xnor U9825 (N_9825,N_8371,N_8284);
nand U9826 (N_9826,N_8806,N_8092);
and U9827 (N_9827,N_8734,N_8553);
and U9828 (N_9828,N_8837,N_8255);
nor U9829 (N_9829,N_8214,N_8196);
nand U9830 (N_9830,N_8950,N_8713);
nor U9831 (N_9831,N_8551,N_8196);
and U9832 (N_9832,N_8522,N_8351);
nand U9833 (N_9833,N_8041,N_8947);
xnor U9834 (N_9834,N_8142,N_8053);
nor U9835 (N_9835,N_8142,N_8227);
nor U9836 (N_9836,N_8006,N_8540);
or U9837 (N_9837,N_8433,N_8753);
nand U9838 (N_9838,N_8669,N_8012);
xor U9839 (N_9839,N_8457,N_8610);
xnor U9840 (N_9840,N_8860,N_8199);
and U9841 (N_9841,N_8192,N_8366);
or U9842 (N_9842,N_8303,N_8325);
xnor U9843 (N_9843,N_8759,N_8842);
and U9844 (N_9844,N_8983,N_8057);
and U9845 (N_9845,N_8839,N_8935);
nand U9846 (N_9846,N_8419,N_8700);
xnor U9847 (N_9847,N_8812,N_8256);
or U9848 (N_9848,N_8120,N_8654);
xnor U9849 (N_9849,N_8029,N_8385);
xnor U9850 (N_9850,N_8256,N_8169);
and U9851 (N_9851,N_8224,N_8048);
and U9852 (N_9852,N_8660,N_8749);
and U9853 (N_9853,N_8326,N_8993);
nor U9854 (N_9854,N_8078,N_8498);
and U9855 (N_9855,N_8204,N_8632);
and U9856 (N_9856,N_8840,N_8495);
nand U9857 (N_9857,N_8404,N_8877);
or U9858 (N_9858,N_8103,N_8298);
and U9859 (N_9859,N_8504,N_8541);
or U9860 (N_9860,N_8841,N_8010);
or U9861 (N_9861,N_8158,N_8230);
nand U9862 (N_9862,N_8550,N_8985);
nor U9863 (N_9863,N_8735,N_8199);
nand U9864 (N_9864,N_8463,N_8906);
nor U9865 (N_9865,N_8568,N_8921);
nand U9866 (N_9866,N_8823,N_8674);
nor U9867 (N_9867,N_8277,N_8460);
nand U9868 (N_9868,N_8076,N_8611);
or U9869 (N_9869,N_8548,N_8327);
and U9870 (N_9870,N_8564,N_8029);
nand U9871 (N_9871,N_8435,N_8785);
nor U9872 (N_9872,N_8561,N_8381);
and U9873 (N_9873,N_8705,N_8317);
and U9874 (N_9874,N_8688,N_8840);
or U9875 (N_9875,N_8195,N_8553);
or U9876 (N_9876,N_8764,N_8063);
xnor U9877 (N_9877,N_8616,N_8118);
nand U9878 (N_9878,N_8790,N_8899);
and U9879 (N_9879,N_8028,N_8467);
nor U9880 (N_9880,N_8638,N_8934);
or U9881 (N_9881,N_8627,N_8766);
or U9882 (N_9882,N_8515,N_8758);
nand U9883 (N_9883,N_8983,N_8180);
and U9884 (N_9884,N_8356,N_8623);
nor U9885 (N_9885,N_8810,N_8887);
nor U9886 (N_9886,N_8343,N_8953);
nand U9887 (N_9887,N_8119,N_8267);
xor U9888 (N_9888,N_8281,N_8761);
or U9889 (N_9889,N_8529,N_8726);
xor U9890 (N_9890,N_8043,N_8237);
nand U9891 (N_9891,N_8031,N_8639);
nand U9892 (N_9892,N_8168,N_8790);
nand U9893 (N_9893,N_8426,N_8125);
xor U9894 (N_9894,N_8225,N_8728);
and U9895 (N_9895,N_8756,N_8607);
nor U9896 (N_9896,N_8774,N_8060);
and U9897 (N_9897,N_8075,N_8378);
nor U9898 (N_9898,N_8125,N_8966);
nand U9899 (N_9899,N_8390,N_8772);
or U9900 (N_9900,N_8414,N_8567);
or U9901 (N_9901,N_8379,N_8599);
xnor U9902 (N_9902,N_8364,N_8636);
or U9903 (N_9903,N_8589,N_8243);
nand U9904 (N_9904,N_8327,N_8460);
nor U9905 (N_9905,N_8568,N_8699);
nand U9906 (N_9906,N_8479,N_8877);
nand U9907 (N_9907,N_8617,N_8185);
nor U9908 (N_9908,N_8190,N_8075);
or U9909 (N_9909,N_8173,N_8877);
or U9910 (N_9910,N_8873,N_8104);
or U9911 (N_9911,N_8623,N_8911);
or U9912 (N_9912,N_8654,N_8540);
nand U9913 (N_9913,N_8931,N_8784);
xnor U9914 (N_9914,N_8459,N_8854);
or U9915 (N_9915,N_8898,N_8398);
and U9916 (N_9916,N_8532,N_8463);
and U9917 (N_9917,N_8297,N_8736);
nor U9918 (N_9918,N_8893,N_8544);
nand U9919 (N_9919,N_8192,N_8931);
or U9920 (N_9920,N_8837,N_8913);
nand U9921 (N_9921,N_8911,N_8796);
nand U9922 (N_9922,N_8203,N_8400);
or U9923 (N_9923,N_8699,N_8408);
xor U9924 (N_9924,N_8674,N_8879);
or U9925 (N_9925,N_8283,N_8945);
or U9926 (N_9926,N_8655,N_8910);
or U9927 (N_9927,N_8729,N_8546);
nor U9928 (N_9928,N_8551,N_8693);
and U9929 (N_9929,N_8600,N_8156);
nand U9930 (N_9930,N_8795,N_8787);
nor U9931 (N_9931,N_8585,N_8722);
nand U9932 (N_9932,N_8211,N_8891);
and U9933 (N_9933,N_8235,N_8054);
xnor U9934 (N_9934,N_8499,N_8368);
and U9935 (N_9935,N_8699,N_8322);
nand U9936 (N_9936,N_8735,N_8093);
and U9937 (N_9937,N_8630,N_8197);
nand U9938 (N_9938,N_8553,N_8837);
or U9939 (N_9939,N_8014,N_8344);
and U9940 (N_9940,N_8565,N_8607);
xnor U9941 (N_9941,N_8954,N_8093);
nand U9942 (N_9942,N_8244,N_8650);
and U9943 (N_9943,N_8507,N_8585);
nor U9944 (N_9944,N_8962,N_8219);
and U9945 (N_9945,N_8080,N_8421);
nand U9946 (N_9946,N_8976,N_8699);
nor U9947 (N_9947,N_8913,N_8115);
nor U9948 (N_9948,N_8052,N_8417);
nor U9949 (N_9949,N_8545,N_8463);
or U9950 (N_9950,N_8995,N_8617);
or U9951 (N_9951,N_8494,N_8285);
and U9952 (N_9952,N_8796,N_8308);
nand U9953 (N_9953,N_8504,N_8162);
or U9954 (N_9954,N_8705,N_8321);
and U9955 (N_9955,N_8753,N_8124);
xor U9956 (N_9956,N_8755,N_8734);
or U9957 (N_9957,N_8974,N_8840);
nand U9958 (N_9958,N_8912,N_8179);
nand U9959 (N_9959,N_8284,N_8662);
and U9960 (N_9960,N_8396,N_8135);
xnor U9961 (N_9961,N_8580,N_8459);
nand U9962 (N_9962,N_8236,N_8302);
nor U9963 (N_9963,N_8774,N_8454);
xor U9964 (N_9964,N_8400,N_8035);
xnor U9965 (N_9965,N_8377,N_8678);
and U9966 (N_9966,N_8524,N_8444);
or U9967 (N_9967,N_8480,N_8474);
nor U9968 (N_9968,N_8634,N_8297);
and U9969 (N_9969,N_8893,N_8843);
xnor U9970 (N_9970,N_8143,N_8725);
nor U9971 (N_9971,N_8797,N_8865);
and U9972 (N_9972,N_8647,N_8654);
and U9973 (N_9973,N_8904,N_8792);
xor U9974 (N_9974,N_8948,N_8108);
nand U9975 (N_9975,N_8096,N_8792);
nor U9976 (N_9976,N_8440,N_8796);
and U9977 (N_9977,N_8164,N_8824);
and U9978 (N_9978,N_8957,N_8414);
and U9979 (N_9979,N_8393,N_8195);
and U9980 (N_9980,N_8039,N_8432);
xor U9981 (N_9981,N_8799,N_8732);
xnor U9982 (N_9982,N_8638,N_8898);
and U9983 (N_9983,N_8459,N_8114);
xnor U9984 (N_9984,N_8271,N_8633);
nor U9985 (N_9985,N_8814,N_8741);
and U9986 (N_9986,N_8539,N_8583);
and U9987 (N_9987,N_8789,N_8627);
nand U9988 (N_9988,N_8900,N_8181);
or U9989 (N_9989,N_8276,N_8327);
nand U9990 (N_9990,N_8278,N_8106);
or U9991 (N_9991,N_8605,N_8969);
nor U9992 (N_9992,N_8302,N_8919);
nand U9993 (N_9993,N_8368,N_8717);
or U9994 (N_9994,N_8090,N_8165);
nand U9995 (N_9995,N_8700,N_8443);
nand U9996 (N_9996,N_8567,N_8844);
nor U9997 (N_9997,N_8661,N_8077);
nand U9998 (N_9998,N_8927,N_8911);
xor U9999 (N_9999,N_8663,N_8948);
and UO_0 (O_0,N_9657,N_9969);
xor UO_1 (O_1,N_9352,N_9158);
nor UO_2 (O_2,N_9424,N_9722);
nand UO_3 (O_3,N_9420,N_9936);
nand UO_4 (O_4,N_9023,N_9426);
nand UO_5 (O_5,N_9759,N_9307);
or UO_6 (O_6,N_9091,N_9959);
nor UO_7 (O_7,N_9731,N_9473);
nor UO_8 (O_8,N_9752,N_9392);
or UO_9 (O_9,N_9806,N_9428);
and UO_10 (O_10,N_9646,N_9043);
and UO_11 (O_11,N_9773,N_9166);
nor UO_12 (O_12,N_9130,N_9522);
or UO_13 (O_13,N_9248,N_9461);
or UO_14 (O_14,N_9183,N_9826);
nand UO_15 (O_15,N_9179,N_9174);
nand UO_16 (O_16,N_9111,N_9156);
xnor UO_17 (O_17,N_9405,N_9421);
nand UO_18 (O_18,N_9438,N_9830);
nor UO_19 (O_19,N_9744,N_9126);
or UO_20 (O_20,N_9104,N_9062);
nand UO_21 (O_21,N_9547,N_9412);
nand UO_22 (O_22,N_9884,N_9184);
nand UO_23 (O_23,N_9114,N_9264);
xor UO_24 (O_24,N_9889,N_9801);
xor UO_25 (O_25,N_9790,N_9131);
nand UO_26 (O_26,N_9384,N_9343);
nor UO_27 (O_27,N_9751,N_9758);
nand UO_28 (O_28,N_9573,N_9194);
xnor UO_29 (O_29,N_9280,N_9219);
nor UO_30 (O_30,N_9479,N_9150);
xor UO_31 (O_31,N_9193,N_9148);
or UO_32 (O_32,N_9778,N_9504);
nor UO_33 (O_33,N_9821,N_9814);
xor UO_34 (O_34,N_9227,N_9332);
xnor UO_35 (O_35,N_9222,N_9747);
nor UO_36 (O_36,N_9923,N_9318);
or UO_37 (O_37,N_9932,N_9305);
nor UO_38 (O_38,N_9609,N_9035);
xor UO_39 (O_39,N_9455,N_9441);
or UO_40 (O_40,N_9781,N_9764);
and UO_41 (O_41,N_9797,N_9724);
and UO_42 (O_42,N_9624,N_9729);
nor UO_43 (O_43,N_9047,N_9966);
nand UO_44 (O_44,N_9268,N_9386);
or UO_45 (O_45,N_9559,N_9477);
nand UO_46 (O_46,N_9917,N_9979);
nand UO_47 (O_47,N_9914,N_9703);
or UO_48 (O_48,N_9768,N_9659);
or UO_49 (O_49,N_9353,N_9937);
xor UO_50 (O_50,N_9031,N_9333);
and UO_51 (O_51,N_9776,N_9257);
nor UO_52 (O_52,N_9246,N_9635);
nor UO_53 (O_53,N_9511,N_9075);
or UO_54 (O_54,N_9896,N_9338);
nand UO_55 (O_55,N_9162,N_9548);
nand UO_56 (O_56,N_9086,N_9367);
and UO_57 (O_57,N_9563,N_9024);
nand UO_58 (O_58,N_9355,N_9039);
and UO_59 (O_59,N_9991,N_9871);
or UO_60 (O_60,N_9147,N_9170);
and UO_61 (O_61,N_9300,N_9551);
or UO_62 (O_62,N_9572,N_9775);
or UO_63 (O_63,N_9198,N_9944);
xnor UO_64 (O_64,N_9651,N_9348);
and UO_65 (O_65,N_9665,N_9427);
nor UO_66 (O_66,N_9452,N_9688);
xnor UO_67 (O_67,N_9383,N_9272);
xor UO_68 (O_68,N_9533,N_9525);
or UO_69 (O_69,N_9457,N_9127);
nand UO_70 (O_70,N_9517,N_9822);
xor UO_71 (O_71,N_9082,N_9143);
xnor UO_72 (O_72,N_9231,N_9520);
or UO_73 (O_73,N_9701,N_9949);
and UO_74 (O_74,N_9341,N_9481);
xnor UO_75 (O_75,N_9065,N_9656);
xor UO_76 (O_76,N_9016,N_9197);
or UO_77 (O_77,N_9259,N_9337);
nand UO_78 (O_78,N_9313,N_9626);
nand UO_79 (O_79,N_9578,N_9209);
nand UO_80 (O_80,N_9850,N_9851);
or UO_81 (O_81,N_9360,N_9908);
or UO_82 (O_82,N_9738,N_9807);
or UO_83 (O_83,N_9238,N_9686);
nor UO_84 (O_84,N_9900,N_9017);
xnor UO_85 (O_85,N_9597,N_9435);
xor UO_86 (O_86,N_9395,N_9458);
and UO_87 (O_87,N_9811,N_9109);
xor UO_88 (O_88,N_9645,N_9403);
nand UO_89 (O_89,N_9630,N_9160);
and UO_90 (O_90,N_9216,N_9014);
and UO_91 (O_91,N_9566,N_9087);
nand UO_92 (O_92,N_9293,N_9494);
xnor UO_93 (O_93,N_9610,N_9555);
xnor UO_94 (O_94,N_9265,N_9389);
and UO_95 (O_95,N_9311,N_9507);
xnor UO_96 (O_96,N_9116,N_9957);
nor UO_97 (O_97,N_9855,N_9402);
nor UO_98 (O_98,N_9967,N_9927);
and UO_99 (O_99,N_9837,N_9954);
and UO_100 (O_100,N_9106,N_9004);
or UO_101 (O_101,N_9053,N_9748);
xnor UO_102 (O_102,N_9363,N_9545);
nand UO_103 (O_103,N_9943,N_9560);
nand UO_104 (O_104,N_9585,N_9780);
xnor UO_105 (O_105,N_9078,N_9097);
nor UO_106 (O_106,N_9877,N_9139);
nor UO_107 (O_107,N_9152,N_9978);
nor UO_108 (O_108,N_9653,N_9115);
xor UO_109 (O_109,N_9103,N_9336);
nor UO_110 (O_110,N_9298,N_9169);
xor UO_111 (O_111,N_9044,N_9051);
nor UO_112 (O_112,N_9490,N_9750);
nand UO_113 (O_113,N_9398,N_9240);
or UO_114 (O_114,N_9819,N_9244);
xnor UO_115 (O_115,N_9813,N_9502);
xnor UO_116 (O_116,N_9330,N_9678);
or UO_117 (O_117,N_9213,N_9679);
or UO_118 (O_118,N_9326,N_9981);
or UO_119 (O_119,N_9207,N_9418);
xnor UO_120 (O_120,N_9045,N_9680);
or UO_121 (O_121,N_9377,N_9171);
or UO_122 (O_122,N_9590,N_9269);
and UO_123 (O_123,N_9327,N_9296);
and UO_124 (O_124,N_9281,N_9677);
xor UO_125 (O_125,N_9536,N_9867);
nand UO_126 (O_126,N_9445,N_9998);
nor UO_127 (O_127,N_9587,N_9380);
or UO_128 (O_128,N_9832,N_9134);
xnor UO_129 (O_129,N_9369,N_9612);
xnor UO_130 (O_130,N_9342,N_9366);
nand UO_131 (O_131,N_9647,N_9549);
nand UO_132 (O_132,N_9436,N_9793);
and UO_133 (O_133,N_9681,N_9586);
nand UO_134 (O_134,N_9770,N_9180);
and UO_135 (O_135,N_9989,N_9382);
nand UO_136 (O_136,N_9655,N_9685);
nand UO_137 (O_137,N_9066,N_9589);
or UO_138 (O_138,N_9081,N_9709);
and UO_139 (O_139,N_9186,N_9829);
nor UO_140 (O_140,N_9123,N_9375);
xor UO_141 (O_141,N_9029,N_9234);
nand UO_142 (O_142,N_9718,N_9915);
or UO_143 (O_143,N_9054,N_9239);
xor UO_144 (O_144,N_9317,N_9093);
nand UO_145 (O_145,N_9245,N_9250);
xnor UO_146 (O_146,N_9279,N_9601);
or UO_147 (O_147,N_9467,N_9926);
and UO_148 (O_148,N_9095,N_9810);
nand UO_149 (O_149,N_9637,N_9475);
or UO_150 (O_150,N_9726,N_9308);
xnor UO_151 (O_151,N_9287,N_9886);
and UO_152 (O_152,N_9059,N_9892);
nand UO_153 (O_153,N_9746,N_9159);
nand UO_154 (O_154,N_9594,N_9975);
or UO_155 (O_155,N_9510,N_9088);
or UO_156 (O_156,N_9816,N_9498);
nand UO_157 (O_157,N_9912,N_9669);
and UO_158 (O_158,N_9530,N_9735);
or UO_159 (O_159,N_9662,N_9113);
nor UO_160 (O_160,N_9101,N_9495);
xnor UO_161 (O_161,N_9956,N_9515);
xor UO_162 (O_162,N_9921,N_9958);
or UO_163 (O_163,N_9357,N_9593);
or UO_164 (O_164,N_9771,N_9523);
nand UO_165 (O_165,N_9347,N_9456);
nand UO_166 (O_166,N_9876,N_9411);
and UO_167 (O_167,N_9579,N_9472);
nor UO_168 (O_168,N_9497,N_9861);
nor UO_169 (O_169,N_9060,N_9191);
or UO_170 (O_170,N_9107,N_9503);
xnor UO_171 (O_171,N_9569,N_9334);
or UO_172 (O_172,N_9464,N_9018);
and UO_173 (O_173,N_9061,N_9026);
xor UO_174 (O_174,N_9805,N_9212);
nand UO_175 (O_175,N_9774,N_9020);
nand UO_176 (O_176,N_9794,N_9391);
nor UO_177 (O_177,N_9521,N_9299);
nand UO_178 (O_178,N_9745,N_9302);
nand UO_179 (O_179,N_9328,N_9310);
and UO_180 (O_180,N_9036,N_9749);
xor UO_181 (O_181,N_9702,N_9903);
nor UO_182 (O_182,N_9815,N_9570);
or UO_183 (O_183,N_9151,N_9725);
xnor UO_184 (O_184,N_9451,N_9071);
nand UO_185 (O_185,N_9176,N_9717);
and UO_186 (O_186,N_9951,N_9195);
and UO_187 (O_187,N_9079,N_9080);
nor UO_188 (O_188,N_9450,N_9527);
and UO_189 (O_189,N_9002,N_9631);
nand UO_190 (O_190,N_9820,N_9836);
and UO_191 (O_191,N_9190,N_9404);
xor UO_192 (O_192,N_9552,N_9543);
xnor UO_193 (O_193,N_9396,N_9072);
or UO_194 (O_194,N_9633,N_9947);
and UO_195 (O_195,N_9682,N_9410);
and UO_196 (O_196,N_9433,N_9406);
or UO_197 (O_197,N_9754,N_9439);
xnor UO_198 (O_198,N_9674,N_9273);
or UO_199 (O_199,N_9690,N_9730);
nor UO_200 (O_200,N_9478,N_9964);
nor UO_201 (O_201,N_9693,N_9262);
nand UO_202 (O_202,N_9182,N_9037);
xnor UO_203 (O_203,N_9137,N_9437);
or UO_204 (O_204,N_9067,N_9295);
xor UO_205 (O_205,N_9303,N_9188);
nor UO_206 (O_206,N_9627,N_9422);
nor UO_207 (O_207,N_9898,N_9972);
nand UO_208 (O_208,N_9835,N_9499);
nand UO_209 (O_209,N_9827,N_9562);
or UO_210 (O_210,N_9909,N_9344);
nand UO_211 (O_211,N_9762,N_9030);
nand UO_212 (O_212,N_9275,N_9432);
nor UO_213 (O_213,N_9987,N_9973);
xor UO_214 (O_214,N_9110,N_9938);
and UO_215 (O_215,N_9666,N_9225);
nand UO_216 (O_216,N_9895,N_9695);
xor UO_217 (O_217,N_9133,N_9741);
xnor UO_218 (O_218,N_9100,N_9581);
and UO_219 (O_219,N_9469,N_9138);
nand UO_220 (O_220,N_9846,N_9795);
xor UO_221 (O_221,N_9173,N_9482);
or UO_222 (O_222,N_9140,N_9644);
nand UO_223 (O_223,N_9052,N_9859);
nand UO_224 (O_224,N_9529,N_9901);
nand UO_225 (O_225,N_9168,N_9471);
xor UO_226 (O_226,N_9615,N_9288);
xor UO_227 (O_227,N_9187,N_9935);
or UO_228 (O_228,N_9924,N_9550);
xor UO_229 (O_229,N_9860,N_9611);
nor UO_230 (O_230,N_9124,N_9955);
or UO_231 (O_231,N_9934,N_9145);
nand UO_232 (O_232,N_9697,N_9509);
and UO_233 (O_233,N_9628,N_9335);
nand UO_234 (O_234,N_9331,N_9387);
nand UO_235 (O_235,N_9112,N_9779);
xnor UO_236 (O_236,N_9144,N_9668);
xor UO_237 (O_237,N_9474,N_9890);
nor UO_238 (O_238,N_9416,N_9099);
nand UO_239 (O_239,N_9089,N_9997);
or UO_240 (O_240,N_9349,N_9493);
and UO_241 (O_241,N_9906,N_9430);
xnor UO_242 (O_242,N_9157,N_9622);
xor UO_243 (O_243,N_9825,N_9289);
and UO_244 (O_244,N_9041,N_9799);
and UO_245 (O_245,N_9266,N_9713);
and UO_246 (O_246,N_9463,N_9316);
nor UO_247 (O_247,N_9962,N_9442);
nor UO_248 (O_248,N_9230,N_9518);
or UO_249 (O_249,N_9519,N_9514);
nor UO_250 (O_250,N_9415,N_9496);
nor UO_251 (O_251,N_9155,N_9417);
and UO_252 (O_252,N_9785,N_9119);
xnor UO_253 (O_253,N_9304,N_9220);
xor UO_254 (O_254,N_9378,N_9325);
and UO_255 (O_255,N_9390,N_9715);
nor UO_256 (O_256,N_9358,N_9643);
and UO_257 (O_257,N_9704,N_9802);
and UO_258 (O_258,N_9929,N_9032);
xnor UO_259 (O_259,N_9397,N_9165);
nor UO_260 (O_260,N_9542,N_9893);
or UO_261 (O_261,N_9034,N_9649);
and UO_262 (O_262,N_9919,N_9648);
or UO_263 (O_263,N_9714,N_9322);
xnor UO_264 (O_264,N_9175,N_9638);
and UO_265 (O_265,N_9995,N_9008);
nand UO_266 (O_266,N_9629,N_9982);
xnor UO_267 (O_267,N_9664,N_9361);
xnor UO_268 (O_268,N_9460,N_9636);
and UO_269 (O_269,N_9146,N_9883);
nand UO_270 (O_270,N_9948,N_9654);
xor UO_271 (O_271,N_9640,N_9761);
nand UO_272 (O_272,N_9185,N_9226);
or UO_273 (O_273,N_9596,N_9940);
or UO_274 (O_274,N_9694,N_9930);
nor UO_275 (O_275,N_9670,N_9491);
and UO_276 (O_276,N_9619,N_9512);
nand UO_277 (O_277,N_9235,N_9800);
nand UO_278 (O_278,N_9723,N_9946);
xor UO_279 (O_279,N_9576,N_9784);
or UO_280 (O_280,N_9808,N_9639);
nor UO_281 (O_281,N_9364,N_9189);
or UO_282 (O_282,N_9920,N_9121);
xor UO_283 (O_283,N_9600,N_9000);
nand UO_284 (O_284,N_9178,N_9447);
xnor UO_285 (O_285,N_9842,N_9215);
xor UO_286 (O_286,N_9323,N_9853);
nor UO_287 (O_287,N_9049,N_9315);
nand UO_288 (O_288,N_9783,N_9076);
xnor UO_289 (O_289,N_9329,N_9069);
xor UO_290 (O_290,N_9362,N_9862);
or UO_291 (O_291,N_9258,N_9271);
and UO_292 (O_292,N_9255,N_9960);
nor UO_293 (O_293,N_9015,N_9534);
nand UO_294 (O_294,N_9869,N_9849);
and UO_295 (O_295,N_9575,N_9561);
and UO_296 (O_296,N_9993,N_9057);
xor UO_297 (O_297,N_9122,N_9873);
xor UO_298 (O_298,N_9286,N_9284);
or UO_299 (O_299,N_9096,N_9251);
and UO_300 (O_300,N_9734,N_9602);
nor UO_301 (O_301,N_9580,N_9848);
or UO_302 (O_302,N_9249,N_9620);
nand UO_303 (O_303,N_9009,N_9218);
or UO_304 (O_304,N_9125,N_9592);
xnor UO_305 (O_305,N_9485,N_9064);
and UO_306 (O_306,N_9388,N_9824);
xnor UO_307 (O_307,N_9028,N_9006);
and UO_308 (O_308,N_9013,N_9261);
or UO_309 (O_309,N_9865,N_9074);
nor UO_310 (O_310,N_9370,N_9046);
or UO_311 (O_311,N_9149,N_9221);
xnor UO_312 (O_312,N_9346,N_9818);
xor UO_313 (O_313,N_9707,N_9831);
nand UO_314 (O_314,N_9988,N_9712);
xor UO_315 (O_315,N_9446,N_9634);
or UO_316 (O_316,N_9894,N_9291);
or UO_317 (O_317,N_9385,N_9449);
and UO_318 (O_318,N_9683,N_9419);
and UO_319 (O_319,N_9990,N_9870);
nor UO_320 (O_320,N_9660,N_9376);
nor UO_321 (O_321,N_9401,N_9443);
or UO_322 (O_322,N_9931,N_9760);
xor UO_323 (O_323,N_9928,N_9732);
and UO_324 (O_324,N_9614,N_9804);
and UO_325 (O_325,N_9070,N_9698);
or UO_326 (O_326,N_9772,N_9274);
or UO_327 (O_327,N_9513,N_9661);
xnor UO_328 (O_328,N_9202,N_9984);
nor UO_329 (O_329,N_9038,N_9902);
or UO_330 (O_330,N_9285,N_9823);
and UO_331 (O_331,N_9073,N_9736);
or UO_332 (O_332,N_9721,N_9650);
xor UO_333 (O_333,N_9618,N_9719);
and UO_334 (O_334,N_9236,N_9623);
or UO_335 (O_335,N_9365,N_9983);
nand UO_336 (O_336,N_9866,N_9206);
nor UO_337 (O_337,N_9834,N_9868);
or UO_338 (O_338,N_9465,N_9658);
or UO_339 (O_339,N_9068,N_9706);
and UO_340 (O_340,N_9933,N_9787);
or UO_341 (O_341,N_9588,N_9217);
and UO_342 (O_342,N_9691,N_9118);
or UO_343 (O_343,N_9526,N_9699);
nor UO_344 (O_344,N_9667,N_9911);
and UO_345 (O_345,N_9440,N_9263);
and UO_346 (O_346,N_9789,N_9223);
or UO_347 (O_347,N_9812,N_9606);
and UO_348 (O_348,N_9994,N_9524);
nand UO_349 (O_349,N_9393,N_9027);
nand UO_350 (O_350,N_9021,N_9407);
nor UO_351 (O_351,N_9083,N_9117);
and UO_352 (O_352,N_9557,N_9408);
nand UO_353 (O_353,N_9373,N_9976);
or UO_354 (O_354,N_9005,N_9753);
and UO_355 (O_355,N_9381,N_9056);
or UO_356 (O_356,N_9192,N_9505);
nor UO_357 (O_357,N_9756,N_9345);
and UO_358 (O_358,N_9539,N_9399);
or UO_359 (O_359,N_9229,N_9181);
nand UO_360 (O_360,N_9444,N_9796);
and UO_361 (O_361,N_9925,N_9888);
xnor UO_362 (O_362,N_9201,N_9564);
or UO_363 (O_363,N_9577,N_9372);
and UO_364 (O_364,N_9306,N_9309);
and UO_365 (O_365,N_9211,N_9875);
xnor UO_366 (O_366,N_9882,N_9922);
xor UO_367 (O_367,N_9292,N_9142);
and UO_368 (O_368,N_9501,N_9558);
nand UO_369 (O_369,N_9048,N_9872);
or UO_370 (O_370,N_9453,N_9058);
nand UO_371 (O_371,N_9094,N_9319);
nor UO_372 (O_372,N_9368,N_9913);
nand UO_373 (O_373,N_9720,N_9077);
nand UO_374 (O_374,N_9809,N_9556);
and UO_375 (O_375,N_9765,N_9843);
or UO_376 (O_376,N_9672,N_9210);
or UO_377 (O_377,N_9102,N_9085);
nor UO_378 (O_378,N_9544,N_9632);
nor UO_379 (O_379,N_9961,N_9232);
nor UO_380 (O_380,N_9763,N_9120);
or UO_381 (O_381,N_9839,N_9742);
or UO_382 (O_382,N_9092,N_9132);
xnor UO_383 (O_383,N_9591,N_9484);
nor UO_384 (O_384,N_9012,N_9791);
nand UO_385 (O_385,N_9583,N_9459);
and UO_386 (O_386,N_9356,N_9727);
nand UO_387 (O_387,N_9425,N_9769);
nor UO_388 (O_388,N_9243,N_9608);
or UO_389 (O_389,N_9625,N_9642);
xnor UO_390 (O_390,N_9007,N_9128);
nor UO_391 (O_391,N_9400,N_9033);
nand UO_392 (O_392,N_9604,N_9878);
and UO_393 (O_393,N_9090,N_9833);
and UO_394 (O_394,N_9616,N_9025);
nor UO_395 (O_395,N_9603,N_9766);
and UO_396 (O_396,N_9199,N_9880);
and UO_397 (O_397,N_9276,N_9413);
xor UO_398 (O_398,N_9571,N_9084);
nor UO_399 (O_399,N_9980,N_9598);
and UO_400 (O_400,N_9354,N_9506);
nand UO_401 (O_401,N_9857,N_9671);
nand UO_402 (O_402,N_9663,N_9595);
and UO_403 (O_403,N_9716,N_9965);
nor UO_404 (O_404,N_9737,N_9001);
xnor UO_405 (O_405,N_9945,N_9242);
nor UO_406 (O_406,N_9105,N_9468);
and UO_407 (O_407,N_9710,N_9177);
xnor UO_408 (O_408,N_9541,N_9108);
xor UO_409 (O_409,N_9500,N_9214);
xnor UO_410 (O_410,N_9740,N_9379);
nor UO_411 (O_411,N_9196,N_9584);
xnor UO_412 (O_412,N_9394,N_9817);
nand UO_413 (O_413,N_9567,N_9905);
xor UO_414 (O_414,N_9696,N_9885);
xnor UO_415 (O_415,N_9055,N_9782);
and UO_416 (O_416,N_9568,N_9767);
or UO_417 (O_417,N_9856,N_9641);
nand UO_418 (O_418,N_9516,N_9454);
xor UO_419 (O_419,N_9466,N_9374);
or UO_420 (O_420,N_9897,N_9700);
and UO_421 (O_421,N_9996,N_9999);
nor UO_422 (O_422,N_9952,N_9711);
xor UO_423 (O_423,N_9540,N_9963);
or UO_424 (O_424,N_9844,N_9350);
or UO_425 (O_425,N_9129,N_9448);
nand UO_426 (O_426,N_9605,N_9260);
nor UO_427 (O_427,N_9554,N_9278);
and UO_428 (O_428,N_9487,N_9879);
or UO_429 (O_429,N_9939,N_9918);
xnor UO_430 (O_430,N_9841,N_9163);
nor UO_431 (O_431,N_9042,N_9204);
xnor UO_432 (O_432,N_9743,N_9968);
and UO_433 (O_433,N_9532,N_9153);
or UO_434 (O_434,N_9786,N_9488);
nor UO_435 (O_435,N_9161,N_9537);
xnor UO_436 (O_436,N_9480,N_9063);
or UO_437 (O_437,N_9253,N_9247);
and UO_438 (O_438,N_9237,N_9010);
nand UO_439 (O_439,N_9953,N_9845);
and UO_440 (O_440,N_9154,N_9907);
nand UO_441 (O_441,N_9970,N_9705);
nor UO_442 (O_442,N_9256,N_9941);
and UO_443 (O_443,N_9891,N_9546);
xnor UO_444 (O_444,N_9676,N_9301);
nand UO_445 (O_445,N_9689,N_9371);
or UO_446 (O_446,N_9254,N_9167);
nand UO_447 (O_447,N_9798,N_9011);
nand UO_448 (O_448,N_9565,N_9476);
nand UO_449 (O_449,N_9205,N_9040);
xnor UO_450 (O_450,N_9904,N_9838);
or UO_451 (O_451,N_9312,N_9486);
xor UO_452 (O_452,N_9692,N_9172);
nor UO_453 (O_453,N_9788,N_9434);
nor UO_454 (O_454,N_9019,N_9423);
nand UO_455 (O_455,N_9224,N_9228);
nor UO_456 (O_456,N_9431,N_9321);
xnor UO_457 (O_457,N_9351,N_9916);
xor UO_458 (O_458,N_9864,N_9673);
nand UO_459 (O_459,N_9582,N_9950);
xnor UO_460 (O_460,N_9733,N_9652);
or UO_461 (O_461,N_9208,N_9599);
nor UO_462 (O_462,N_9409,N_9992);
nor UO_463 (O_463,N_9282,N_9359);
nor UO_464 (O_464,N_9977,N_9852);
nand UO_465 (O_465,N_9863,N_9429);
and UO_466 (O_466,N_9971,N_9270);
and UO_467 (O_467,N_9050,N_9854);
nand UO_468 (O_468,N_9141,N_9290);
and UO_469 (O_469,N_9022,N_9617);
nand UO_470 (O_470,N_9553,N_9607);
xnor UO_471 (O_471,N_9233,N_9320);
nor UO_472 (O_472,N_9755,N_9986);
xnor UO_473 (O_473,N_9470,N_9528);
nor UO_474 (O_474,N_9483,N_9538);
nor UO_475 (O_475,N_9881,N_9899);
nor UO_476 (O_476,N_9098,N_9847);
or UO_477 (O_477,N_9203,N_9492);
nand UO_478 (O_478,N_9340,N_9283);
or UO_479 (O_479,N_9462,N_9414);
or UO_480 (O_480,N_9277,N_9252);
or UO_481 (O_481,N_9136,N_9687);
xor UO_482 (O_482,N_9241,N_9684);
xnor UO_483 (O_483,N_9858,N_9200);
and UO_484 (O_484,N_9792,N_9675);
or UO_485 (O_485,N_9297,N_9613);
nor UO_486 (O_486,N_9708,N_9339);
nor UO_487 (O_487,N_9985,N_9294);
and UO_488 (O_488,N_9757,N_9003);
nand UO_489 (O_489,N_9531,N_9728);
nor UO_490 (O_490,N_9828,N_9267);
and UO_491 (O_491,N_9910,N_9974);
nor UO_492 (O_492,N_9508,N_9535);
nand UO_493 (O_493,N_9164,N_9739);
nor UO_494 (O_494,N_9314,N_9574);
xnor UO_495 (O_495,N_9489,N_9840);
nor UO_496 (O_496,N_9942,N_9621);
nand UO_497 (O_497,N_9777,N_9803);
or UO_498 (O_498,N_9135,N_9874);
or UO_499 (O_499,N_9324,N_9887);
xor UO_500 (O_500,N_9558,N_9560);
and UO_501 (O_501,N_9351,N_9321);
xnor UO_502 (O_502,N_9196,N_9057);
nand UO_503 (O_503,N_9814,N_9981);
xor UO_504 (O_504,N_9725,N_9226);
and UO_505 (O_505,N_9933,N_9418);
xor UO_506 (O_506,N_9316,N_9505);
or UO_507 (O_507,N_9431,N_9114);
or UO_508 (O_508,N_9465,N_9593);
xnor UO_509 (O_509,N_9332,N_9572);
nand UO_510 (O_510,N_9327,N_9791);
or UO_511 (O_511,N_9646,N_9016);
xor UO_512 (O_512,N_9830,N_9907);
nor UO_513 (O_513,N_9687,N_9440);
nor UO_514 (O_514,N_9971,N_9747);
and UO_515 (O_515,N_9285,N_9690);
nand UO_516 (O_516,N_9141,N_9460);
nor UO_517 (O_517,N_9567,N_9469);
or UO_518 (O_518,N_9642,N_9835);
nand UO_519 (O_519,N_9377,N_9162);
nand UO_520 (O_520,N_9370,N_9619);
or UO_521 (O_521,N_9638,N_9602);
nand UO_522 (O_522,N_9545,N_9800);
xor UO_523 (O_523,N_9452,N_9477);
nor UO_524 (O_524,N_9358,N_9029);
nor UO_525 (O_525,N_9828,N_9356);
xnor UO_526 (O_526,N_9498,N_9194);
nand UO_527 (O_527,N_9041,N_9065);
xor UO_528 (O_528,N_9220,N_9369);
xnor UO_529 (O_529,N_9843,N_9749);
nor UO_530 (O_530,N_9582,N_9641);
nor UO_531 (O_531,N_9263,N_9452);
xor UO_532 (O_532,N_9556,N_9091);
nor UO_533 (O_533,N_9430,N_9806);
nand UO_534 (O_534,N_9678,N_9595);
nand UO_535 (O_535,N_9627,N_9034);
and UO_536 (O_536,N_9726,N_9696);
nor UO_537 (O_537,N_9800,N_9239);
nor UO_538 (O_538,N_9488,N_9909);
nor UO_539 (O_539,N_9114,N_9543);
and UO_540 (O_540,N_9748,N_9598);
nor UO_541 (O_541,N_9293,N_9654);
or UO_542 (O_542,N_9243,N_9864);
and UO_543 (O_543,N_9556,N_9854);
and UO_544 (O_544,N_9648,N_9162);
nand UO_545 (O_545,N_9112,N_9777);
nand UO_546 (O_546,N_9852,N_9010);
and UO_547 (O_547,N_9649,N_9550);
xor UO_548 (O_548,N_9252,N_9237);
xnor UO_549 (O_549,N_9646,N_9609);
nand UO_550 (O_550,N_9425,N_9876);
or UO_551 (O_551,N_9766,N_9618);
and UO_552 (O_552,N_9572,N_9014);
nand UO_553 (O_553,N_9417,N_9849);
nand UO_554 (O_554,N_9683,N_9830);
and UO_555 (O_555,N_9966,N_9690);
and UO_556 (O_556,N_9809,N_9223);
nand UO_557 (O_557,N_9579,N_9876);
xnor UO_558 (O_558,N_9410,N_9690);
and UO_559 (O_559,N_9317,N_9873);
nand UO_560 (O_560,N_9325,N_9508);
nor UO_561 (O_561,N_9853,N_9063);
and UO_562 (O_562,N_9409,N_9087);
xnor UO_563 (O_563,N_9804,N_9083);
xor UO_564 (O_564,N_9385,N_9798);
and UO_565 (O_565,N_9426,N_9102);
nand UO_566 (O_566,N_9152,N_9172);
nand UO_567 (O_567,N_9821,N_9015);
nor UO_568 (O_568,N_9116,N_9478);
and UO_569 (O_569,N_9204,N_9962);
and UO_570 (O_570,N_9605,N_9547);
nor UO_571 (O_571,N_9636,N_9716);
and UO_572 (O_572,N_9085,N_9459);
xor UO_573 (O_573,N_9986,N_9811);
nor UO_574 (O_574,N_9620,N_9824);
xnor UO_575 (O_575,N_9377,N_9749);
xnor UO_576 (O_576,N_9373,N_9551);
xnor UO_577 (O_577,N_9734,N_9308);
nor UO_578 (O_578,N_9806,N_9481);
nor UO_579 (O_579,N_9280,N_9484);
and UO_580 (O_580,N_9658,N_9848);
xnor UO_581 (O_581,N_9353,N_9488);
nand UO_582 (O_582,N_9142,N_9837);
and UO_583 (O_583,N_9635,N_9425);
and UO_584 (O_584,N_9064,N_9757);
nand UO_585 (O_585,N_9608,N_9299);
nand UO_586 (O_586,N_9324,N_9411);
or UO_587 (O_587,N_9302,N_9562);
or UO_588 (O_588,N_9546,N_9069);
or UO_589 (O_589,N_9561,N_9099);
nand UO_590 (O_590,N_9783,N_9584);
xor UO_591 (O_591,N_9770,N_9049);
nor UO_592 (O_592,N_9125,N_9583);
nand UO_593 (O_593,N_9611,N_9407);
or UO_594 (O_594,N_9519,N_9484);
and UO_595 (O_595,N_9343,N_9762);
nor UO_596 (O_596,N_9037,N_9649);
nand UO_597 (O_597,N_9205,N_9241);
or UO_598 (O_598,N_9487,N_9408);
nor UO_599 (O_599,N_9911,N_9769);
and UO_600 (O_600,N_9021,N_9387);
or UO_601 (O_601,N_9652,N_9961);
and UO_602 (O_602,N_9776,N_9983);
and UO_603 (O_603,N_9021,N_9749);
nand UO_604 (O_604,N_9077,N_9269);
xnor UO_605 (O_605,N_9234,N_9290);
or UO_606 (O_606,N_9367,N_9525);
nand UO_607 (O_607,N_9689,N_9854);
xor UO_608 (O_608,N_9153,N_9493);
or UO_609 (O_609,N_9474,N_9850);
and UO_610 (O_610,N_9703,N_9157);
and UO_611 (O_611,N_9689,N_9282);
xor UO_612 (O_612,N_9058,N_9966);
nand UO_613 (O_613,N_9645,N_9780);
or UO_614 (O_614,N_9664,N_9914);
nor UO_615 (O_615,N_9510,N_9648);
xor UO_616 (O_616,N_9552,N_9643);
or UO_617 (O_617,N_9976,N_9043);
nor UO_618 (O_618,N_9046,N_9719);
and UO_619 (O_619,N_9534,N_9487);
or UO_620 (O_620,N_9765,N_9346);
nor UO_621 (O_621,N_9017,N_9655);
and UO_622 (O_622,N_9791,N_9928);
or UO_623 (O_623,N_9368,N_9819);
or UO_624 (O_624,N_9242,N_9590);
nand UO_625 (O_625,N_9553,N_9576);
or UO_626 (O_626,N_9331,N_9125);
and UO_627 (O_627,N_9856,N_9373);
and UO_628 (O_628,N_9186,N_9881);
or UO_629 (O_629,N_9298,N_9483);
and UO_630 (O_630,N_9952,N_9723);
and UO_631 (O_631,N_9995,N_9336);
xor UO_632 (O_632,N_9012,N_9728);
nor UO_633 (O_633,N_9122,N_9990);
xnor UO_634 (O_634,N_9172,N_9552);
xnor UO_635 (O_635,N_9366,N_9005);
and UO_636 (O_636,N_9748,N_9575);
or UO_637 (O_637,N_9687,N_9912);
or UO_638 (O_638,N_9560,N_9991);
and UO_639 (O_639,N_9848,N_9184);
xnor UO_640 (O_640,N_9445,N_9319);
or UO_641 (O_641,N_9275,N_9101);
and UO_642 (O_642,N_9422,N_9771);
xnor UO_643 (O_643,N_9276,N_9416);
nor UO_644 (O_644,N_9553,N_9798);
and UO_645 (O_645,N_9792,N_9966);
xnor UO_646 (O_646,N_9859,N_9761);
xnor UO_647 (O_647,N_9297,N_9024);
nor UO_648 (O_648,N_9617,N_9661);
xor UO_649 (O_649,N_9252,N_9622);
nor UO_650 (O_650,N_9662,N_9580);
nor UO_651 (O_651,N_9318,N_9271);
nor UO_652 (O_652,N_9974,N_9283);
and UO_653 (O_653,N_9583,N_9808);
or UO_654 (O_654,N_9655,N_9241);
and UO_655 (O_655,N_9296,N_9233);
nand UO_656 (O_656,N_9505,N_9941);
or UO_657 (O_657,N_9172,N_9946);
nand UO_658 (O_658,N_9623,N_9171);
xnor UO_659 (O_659,N_9307,N_9647);
xor UO_660 (O_660,N_9329,N_9622);
nand UO_661 (O_661,N_9014,N_9032);
nand UO_662 (O_662,N_9631,N_9204);
or UO_663 (O_663,N_9016,N_9078);
or UO_664 (O_664,N_9880,N_9949);
and UO_665 (O_665,N_9036,N_9631);
or UO_666 (O_666,N_9729,N_9609);
xnor UO_667 (O_667,N_9393,N_9433);
and UO_668 (O_668,N_9027,N_9108);
and UO_669 (O_669,N_9312,N_9452);
xnor UO_670 (O_670,N_9377,N_9776);
nand UO_671 (O_671,N_9729,N_9058);
or UO_672 (O_672,N_9185,N_9252);
xnor UO_673 (O_673,N_9525,N_9883);
and UO_674 (O_674,N_9374,N_9349);
nand UO_675 (O_675,N_9873,N_9436);
nand UO_676 (O_676,N_9893,N_9348);
or UO_677 (O_677,N_9367,N_9022);
nor UO_678 (O_678,N_9900,N_9042);
and UO_679 (O_679,N_9443,N_9329);
nor UO_680 (O_680,N_9824,N_9108);
nor UO_681 (O_681,N_9595,N_9090);
xnor UO_682 (O_682,N_9308,N_9352);
nor UO_683 (O_683,N_9358,N_9010);
nand UO_684 (O_684,N_9221,N_9410);
xor UO_685 (O_685,N_9888,N_9211);
and UO_686 (O_686,N_9074,N_9741);
nor UO_687 (O_687,N_9676,N_9579);
nand UO_688 (O_688,N_9575,N_9939);
and UO_689 (O_689,N_9220,N_9483);
nor UO_690 (O_690,N_9014,N_9956);
or UO_691 (O_691,N_9291,N_9664);
xor UO_692 (O_692,N_9175,N_9210);
and UO_693 (O_693,N_9299,N_9326);
or UO_694 (O_694,N_9584,N_9193);
or UO_695 (O_695,N_9613,N_9615);
nor UO_696 (O_696,N_9233,N_9507);
or UO_697 (O_697,N_9071,N_9165);
nand UO_698 (O_698,N_9223,N_9284);
nand UO_699 (O_699,N_9001,N_9460);
xnor UO_700 (O_700,N_9010,N_9687);
xnor UO_701 (O_701,N_9055,N_9050);
nand UO_702 (O_702,N_9798,N_9550);
or UO_703 (O_703,N_9033,N_9514);
xor UO_704 (O_704,N_9861,N_9867);
nor UO_705 (O_705,N_9129,N_9070);
nor UO_706 (O_706,N_9411,N_9517);
nand UO_707 (O_707,N_9700,N_9761);
nand UO_708 (O_708,N_9012,N_9149);
nor UO_709 (O_709,N_9599,N_9682);
nand UO_710 (O_710,N_9588,N_9599);
and UO_711 (O_711,N_9020,N_9289);
and UO_712 (O_712,N_9924,N_9863);
and UO_713 (O_713,N_9654,N_9227);
nor UO_714 (O_714,N_9745,N_9727);
xor UO_715 (O_715,N_9964,N_9877);
xor UO_716 (O_716,N_9854,N_9410);
and UO_717 (O_717,N_9447,N_9397);
xor UO_718 (O_718,N_9504,N_9370);
xnor UO_719 (O_719,N_9191,N_9580);
xnor UO_720 (O_720,N_9779,N_9128);
xor UO_721 (O_721,N_9095,N_9797);
nand UO_722 (O_722,N_9943,N_9581);
or UO_723 (O_723,N_9036,N_9769);
nand UO_724 (O_724,N_9252,N_9422);
xor UO_725 (O_725,N_9247,N_9552);
nor UO_726 (O_726,N_9819,N_9278);
xnor UO_727 (O_727,N_9484,N_9832);
or UO_728 (O_728,N_9429,N_9714);
and UO_729 (O_729,N_9223,N_9808);
xnor UO_730 (O_730,N_9580,N_9992);
nand UO_731 (O_731,N_9620,N_9408);
and UO_732 (O_732,N_9400,N_9120);
xnor UO_733 (O_733,N_9291,N_9362);
or UO_734 (O_734,N_9702,N_9530);
nand UO_735 (O_735,N_9235,N_9686);
or UO_736 (O_736,N_9076,N_9082);
or UO_737 (O_737,N_9654,N_9344);
and UO_738 (O_738,N_9821,N_9014);
xnor UO_739 (O_739,N_9072,N_9461);
xor UO_740 (O_740,N_9375,N_9713);
nand UO_741 (O_741,N_9463,N_9528);
xor UO_742 (O_742,N_9652,N_9948);
xnor UO_743 (O_743,N_9158,N_9024);
and UO_744 (O_744,N_9396,N_9385);
nand UO_745 (O_745,N_9769,N_9768);
or UO_746 (O_746,N_9499,N_9121);
xor UO_747 (O_747,N_9978,N_9110);
nand UO_748 (O_748,N_9678,N_9991);
xnor UO_749 (O_749,N_9551,N_9003);
or UO_750 (O_750,N_9031,N_9023);
nor UO_751 (O_751,N_9593,N_9991);
xnor UO_752 (O_752,N_9651,N_9124);
nor UO_753 (O_753,N_9807,N_9288);
or UO_754 (O_754,N_9074,N_9467);
and UO_755 (O_755,N_9785,N_9406);
nand UO_756 (O_756,N_9151,N_9365);
and UO_757 (O_757,N_9298,N_9450);
and UO_758 (O_758,N_9156,N_9389);
nand UO_759 (O_759,N_9532,N_9792);
or UO_760 (O_760,N_9553,N_9870);
and UO_761 (O_761,N_9843,N_9482);
nor UO_762 (O_762,N_9366,N_9989);
nor UO_763 (O_763,N_9972,N_9848);
xnor UO_764 (O_764,N_9624,N_9804);
nand UO_765 (O_765,N_9738,N_9690);
nor UO_766 (O_766,N_9860,N_9145);
or UO_767 (O_767,N_9075,N_9716);
and UO_768 (O_768,N_9610,N_9033);
and UO_769 (O_769,N_9853,N_9725);
nand UO_770 (O_770,N_9901,N_9493);
nor UO_771 (O_771,N_9542,N_9603);
and UO_772 (O_772,N_9817,N_9863);
nand UO_773 (O_773,N_9887,N_9290);
nor UO_774 (O_774,N_9070,N_9767);
xor UO_775 (O_775,N_9219,N_9385);
xor UO_776 (O_776,N_9781,N_9990);
or UO_777 (O_777,N_9191,N_9954);
xor UO_778 (O_778,N_9126,N_9902);
or UO_779 (O_779,N_9222,N_9087);
xnor UO_780 (O_780,N_9875,N_9833);
nor UO_781 (O_781,N_9127,N_9669);
nand UO_782 (O_782,N_9804,N_9296);
nor UO_783 (O_783,N_9676,N_9103);
xor UO_784 (O_784,N_9471,N_9550);
nor UO_785 (O_785,N_9489,N_9868);
xor UO_786 (O_786,N_9238,N_9478);
or UO_787 (O_787,N_9204,N_9975);
and UO_788 (O_788,N_9798,N_9887);
and UO_789 (O_789,N_9570,N_9805);
nor UO_790 (O_790,N_9259,N_9326);
xor UO_791 (O_791,N_9408,N_9568);
nand UO_792 (O_792,N_9714,N_9318);
xnor UO_793 (O_793,N_9100,N_9902);
nor UO_794 (O_794,N_9527,N_9615);
xnor UO_795 (O_795,N_9437,N_9399);
and UO_796 (O_796,N_9781,N_9723);
nand UO_797 (O_797,N_9618,N_9751);
or UO_798 (O_798,N_9876,N_9803);
or UO_799 (O_799,N_9402,N_9810);
and UO_800 (O_800,N_9288,N_9779);
and UO_801 (O_801,N_9660,N_9357);
nand UO_802 (O_802,N_9212,N_9381);
nand UO_803 (O_803,N_9142,N_9471);
or UO_804 (O_804,N_9679,N_9487);
nand UO_805 (O_805,N_9556,N_9623);
or UO_806 (O_806,N_9809,N_9600);
nor UO_807 (O_807,N_9529,N_9091);
nand UO_808 (O_808,N_9689,N_9075);
and UO_809 (O_809,N_9452,N_9673);
nand UO_810 (O_810,N_9821,N_9917);
and UO_811 (O_811,N_9344,N_9429);
and UO_812 (O_812,N_9449,N_9887);
and UO_813 (O_813,N_9603,N_9636);
nor UO_814 (O_814,N_9680,N_9027);
and UO_815 (O_815,N_9468,N_9746);
and UO_816 (O_816,N_9962,N_9330);
or UO_817 (O_817,N_9864,N_9498);
or UO_818 (O_818,N_9623,N_9242);
or UO_819 (O_819,N_9271,N_9937);
or UO_820 (O_820,N_9996,N_9500);
xnor UO_821 (O_821,N_9303,N_9658);
xnor UO_822 (O_822,N_9655,N_9874);
or UO_823 (O_823,N_9610,N_9646);
and UO_824 (O_824,N_9940,N_9373);
or UO_825 (O_825,N_9345,N_9437);
or UO_826 (O_826,N_9626,N_9318);
or UO_827 (O_827,N_9793,N_9359);
xnor UO_828 (O_828,N_9907,N_9922);
xor UO_829 (O_829,N_9740,N_9557);
xor UO_830 (O_830,N_9167,N_9006);
or UO_831 (O_831,N_9860,N_9128);
or UO_832 (O_832,N_9842,N_9504);
xnor UO_833 (O_833,N_9722,N_9532);
nand UO_834 (O_834,N_9353,N_9397);
nor UO_835 (O_835,N_9169,N_9007);
nand UO_836 (O_836,N_9225,N_9601);
xnor UO_837 (O_837,N_9783,N_9379);
xor UO_838 (O_838,N_9052,N_9729);
xor UO_839 (O_839,N_9481,N_9657);
nor UO_840 (O_840,N_9045,N_9880);
nor UO_841 (O_841,N_9632,N_9954);
and UO_842 (O_842,N_9523,N_9551);
and UO_843 (O_843,N_9978,N_9964);
xor UO_844 (O_844,N_9946,N_9481);
nand UO_845 (O_845,N_9167,N_9680);
and UO_846 (O_846,N_9109,N_9072);
nor UO_847 (O_847,N_9124,N_9573);
nand UO_848 (O_848,N_9866,N_9845);
or UO_849 (O_849,N_9339,N_9855);
nor UO_850 (O_850,N_9493,N_9564);
nor UO_851 (O_851,N_9087,N_9351);
nor UO_852 (O_852,N_9668,N_9143);
nand UO_853 (O_853,N_9346,N_9452);
xnor UO_854 (O_854,N_9132,N_9311);
nand UO_855 (O_855,N_9482,N_9779);
nand UO_856 (O_856,N_9070,N_9082);
xnor UO_857 (O_857,N_9418,N_9821);
nand UO_858 (O_858,N_9678,N_9797);
and UO_859 (O_859,N_9614,N_9621);
xor UO_860 (O_860,N_9921,N_9177);
nand UO_861 (O_861,N_9089,N_9143);
xnor UO_862 (O_862,N_9439,N_9630);
nor UO_863 (O_863,N_9219,N_9310);
or UO_864 (O_864,N_9440,N_9866);
or UO_865 (O_865,N_9115,N_9735);
nor UO_866 (O_866,N_9513,N_9419);
or UO_867 (O_867,N_9723,N_9108);
xor UO_868 (O_868,N_9172,N_9655);
or UO_869 (O_869,N_9637,N_9126);
and UO_870 (O_870,N_9872,N_9571);
nand UO_871 (O_871,N_9591,N_9178);
xor UO_872 (O_872,N_9085,N_9568);
and UO_873 (O_873,N_9538,N_9744);
nor UO_874 (O_874,N_9661,N_9313);
and UO_875 (O_875,N_9129,N_9301);
and UO_876 (O_876,N_9441,N_9348);
nor UO_877 (O_877,N_9837,N_9829);
or UO_878 (O_878,N_9532,N_9292);
and UO_879 (O_879,N_9095,N_9275);
nor UO_880 (O_880,N_9814,N_9508);
or UO_881 (O_881,N_9836,N_9278);
xor UO_882 (O_882,N_9341,N_9067);
xnor UO_883 (O_883,N_9592,N_9599);
nor UO_884 (O_884,N_9259,N_9126);
xnor UO_885 (O_885,N_9540,N_9460);
xor UO_886 (O_886,N_9648,N_9357);
and UO_887 (O_887,N_9364,N_9959);
xor UO_888 (O_888,N_9260,N_9852);
or UO_889 (O_889,N_9623,N_9235);
nand UO_890 (O_890,N_9818,N_9502);
xor UO_891 (O_891,N_9447,N_9935);
nand UO_892 (O_892,N_9945,N_9827);
xnor UO_893 (O_893,N_9090,N_9332);
nor UO_894 (O_894,N_9672,N_9226);
or UO_895 (O_895,N_9580,N_9428);
or UO_896 (O_896,N_9320,N_9553);
and UO_897 (O_897,N_9959,N_9171);
or UO_898 (O_898,N_9144,N_9091);
nor UO_899 (O_899,N_9033,N_9988);
and UO_900 (O_900,N_9401,N_9851);
nor UO_901 (O_901,N_9962,N_9525);
nor UO_902 (O_902,N_9972,N_9277);
nand UO_903 (O_903,N_9071,N_9257);
nor UO_904 (O_904,N_9298,N_9504);
xnor UO_905 (O_905,N_9168,N_9508);
and UO_906 (O_906,N_9874,N_9136);
nor UO_907 (O_907,N_9692,N_9971);
nor UO_908 (O_908,N_9816,N_9262);
nand UO_909 (O_909,N_9353,N_9600);
and UO_910 (O_910,N_9645,N_9893);
nand UO_911 (O_911,N_9570,N_9488);
nor UO_912 (O_912,N_9530,N_9168);
or UO_913 (O_913,N_9414,N_9883);
nand UO_914 (O_914,N_9384,N_9493);
and UO_915 (O_915,N_9405,N_9977);
or UO_916 (O_916,N_9676,N_9949);
or UO_917 (O_917,N_9024,N_9656);
and UO_918 (O_918,N_9524,N_9185);
or UO_919 (O_919,N_9038,N_9414);
xor UO_920 (O_920,N_9636,N_9303);
xor UO_921 (O_921,N_9667,N_9644);
and UO_922 (O_922,N_9776,N_9181);
or UO_923 (O_923,N_9185,N_9608);
nor UO_924 (O_924,N_9395,N_9387);
xor UO_925 (O_925,N_9621,N_9112);
or UO_926 (O_926,N_9375,N_9614);
and UO_927 (O_927,N_9783,N_9359);
or UO_928 (O_928,N_9438,N_9767);
or UO_929 (O_929,N_9122,N_9287);
and UO_930 (O_930,N_9079,N_9191);
xor UO_931 (O_931,N_9216,N_9784);
nand UO_932 (O_932,N_9496,N_9389);
nor UO_933 (O_933,N_9242,N_9841);
xor UO_934 (O_934,N_9012,N_9216);
xnor UO_935 (O_935,N_9057,N_9875);
nand UO_936 (O_936,N_9032,N_9218);
and UO_937 (O_937,N_9569,N_9226);
nor UO_938 (O_938,N_9348,N_9968);
nor UO_939 (O_939,N_9529,N_9241);
nor UO_940 (O_940,N_9617,N_9433);
or UO_941 (O_941,N_9668,N_9847);
xnor UO_942 (O_942,N_9995,N_9657);
nor UO_943 (O_943,N_9265,N_9936);
or UO_944 (O_944,N_9468,N_9704);
nand UO_945 (O_945,N_9341,N_9705);
or UO_946 (O_946,N_9641,N_9668);
or UO_947 (O_947,N_9596,N_9271);
nand UO_948 (O_948,N_9147,N_9894);
nor UO_949 (O_949,N_9367,N_9885);
and UO_950 (O_950,N_9063,N_9043);
xor UO_951 (O_951,N_9792,N_9276);
or UO_952 (O_952,N_9311,N_9930);
nand UO_953 (O_953,N_9630,N_9443);
xor UO_954 (O_954,N_9261,N_9498);
nand UO_955 (O_955,N_9792,N_9225);
nor UO_956 (O_956,N_9802,N_9846);
nand UO_957 (O_957,N_9600,N_9753);
xnor UO_958 (O_958,N_9146,N_9778);
and UO_959 (O_959,N_9756,N_9076);
xor UO_960 (O_960,N_9740,N_9920);
xnor UO_961 (O_961,N_9641,N_9182);
nand UO_962 (O_962,N_9777,N_9641);
xor UO_963 (O_963,N_9392,N_9072);
or UO_964 (O_964,N_9454,N_9729);
nand UO_965 (O_965,N_9124,N_9978);
xor UO_966 (O_966,N_9397,N_9269);
or UO_967 (O_967,N_9511,N_9462);
xor UO_968 (O_968,N_9298,N_9117);
nor UO_969 (O_969,N_9881,N_9180);
nor UO_970 (O_970,N_9252,N_9114);
and UO_971 (O_971,N_9840,N_9600);
and UO_972 (O_972,N_9135,N_9176);
and UO_973 (O_973,N_9129,N_9946);
and UO_974 (O_974,N_9952,N_9205);
and UO_975 (O_975,N_9328,N_9316);
nand UO_976 (O_976,N_9022,N_9028);
nor UO_977 (O_977,N_9110,N_9566);
and UO_978 (O_978,N_9680,N_9702);
nand UO_979 (O_979,N_9349,N_9269);
nor UO_980 (O_980,N_9849,N_9215);
nor UO_981 (O_981,N_9281,N_9988);
xnor UO_982 (O_982,N_9780,N_9222);
nand UO_983 (O_983,N_9745,N_9127);
xnor UO_984 (O_984,N_9761,N_9552);
nor UO_985 (O_985,N_9117,N_9518);
nand UO_986 (O_986,N_9781,N_9553);
and UO_987 (O_987,N_9480,N_9040);
xnor UO_988 (O_988,N_9358,N_9519);
nand UO_989 (O_989,N_9696,N_9819);
and UO_990 (O_990,N_9478,N_9071);
or UO_991 (O_991,N_9166,N_9347);
nand UO_992 (O_992,N_9075,N_9319);
and UO_993 (O_993,N_9891,N_9705);
xor UO_994 (O_994,N_9237,N_9602);
or UO_995 (O_995,N_9896,N_9620);
and UO_996 (O_996,N_9958,N_9342);
nand UO_997 (O_997,N_9477,N_9919);
xnor UO_998 (O_998,N_9936,N_9404);
or UO_999 (O_999,N_9691,N_9537);
and UO_1000 (O_1000,N_9106,N_9176);
xor UO_1001 (O_1001,N_9638,N_9347);
and UO_1002 (O_1002,N_9814,N_9862);
and UO_1003 (O_1003,N_9301,N_9141);
nor UO_1004 (O_1004,N_9628,N_9488);
xnor UO_1005 (O_1005,N_9024,N_9979);
and UO_1006 (O_1006,N_9738,N_9352);
nand UO_1007 (O_1007,N_9948,N_9119);
nand UO_1008 (O_1008,N_9855,N_9306);
nand UO_1009 (O_1009,N_9757,N_9344);
xor UO_1010 (O_1010,N_9002,N_9721);
and UO_1011 (O_1011,N_9834,N_9844);
nor UO_1012 (O_1012,N_9377,N_9783);
nor UO_1013 (O_1013,N_9118,N_9214);
and UO_1014 (O_1014,N_9708,N_9071);
nand UO_1015 (O_1015,N_9239,N_9514);
and UO_1016 (O_1016,N_9022,N_9114);
xor UO_1017 (O_1017,N_9382,N_9467);
nand UO_1018 (O_1018,N_9924,N_9575);
nor UO_1019 (O_1019,N_9443,N_9856);
nand UO_1020 (O_1020,N_9954,N_9278);
and UO_1021 (O_1021,N_9715,N_9427);
nand UO_1022 (O_1022,N_9159,N_9284);
xor UO_1023 (O_1023,N_9690,N_9231);
and UO_1024 (O_1024,N_9514,N_9003);
nor UO_1025 (O_1025,N_9225,N_9937);
nand UO_1026 (O_1026,N_9807,N_9139);
and UO_1027 (O_1027,N_9460,N_9419);
nor UO_1028 (O_1028,N_9181,N_9015);
xnor UO_1029 (O_1029,N_9119,N_9340);
and UO_1030 (O_1030,N_9511,N_9530);
xor UO_1031 (O_1031,N_9733,N_9427);
xnor UO_1032 (O_1032,N_9940,N_9320);
and UO_1033 (O_1033,N_9656,N_9542);
and UO_1034 (O_1034,N_9688,N_9653);
nand UO_1035 (O_1035,N_9344,N_9026);
or UO_1036 (O_1036,N_9146,N_9413);
or UO_1037 (O_1037,N_9551,N_9053);
nor UO_1038 (O_1038,N_9422,N_9728);
nor UO_1039 (O_1039,N_9128,N_9348);
nor UO_1040 (O_1040,N_9827,N_9225);
and UO_1041 (O_1041,N_9318,N_9237);
and UO_1042 (O_1042,N_9048,N_9072);
nand UO_1043 (O_1043,N_9761,N_9119);
xor UO_1044 (O_1044,N_9499,N_9896);
nor UO_1045 (O_1045,N_9364,N_9014);
nor UO_1046 (O_1046,N_9003,N_9737);
nor UO_1047 (O_1047,N_9635,N_9156);
or UO_1048 (O_1048,N_9629,N_9768);
nor UO_1049 (O_1049,N_9137,N_9353);
xor UO_1050 (O_1050,N_9140,N_9787);
nor UO_1051 (O_1051,N_9181,N_9940);
nor UO_1052 (O_1052,N_9390,N_9006);
or UO_1053 (O_1053,N_9363,N_9945);
and UO_1054 (O_1054,N_9753,N_9986);
nand UO_1055 (O_1055,N_9015,N_9166);
nand UO_1056 (O_1056,N_9795,N_9984);
xnor UO_1057 (O_1057,N_9665,N_9026);
nor UO_1058 (O_1058,N_9569,N_9770);
xor UO_1059 (O_1059,N_9011,N_9097);
nor UO_1060 (O_1060,N_9775,N_9148);
nor UO_1061 (O_1061,N_9271,N_9921);
nor UO_1062 (O_1062,N_9008,N_9296);
nand UO_1063 (O_1063,N_9093,N_9407);
nor UO_1064 (O_1064,N_9324,N_9658);
nor UO_1065 (O_1065,N_9117,N_9925);
nand UO_1066 (O_1066,N_9329,N_9335);
nor UO_1067 (O_1067,N_9982,N_9153);
and UO_1068 (O_1068,N_9651,N_9443);
or UO_1069 (O_1069,N_9879,N_9475);
and UO_1070 (O_1070,N_9540,N_9761);
nand UO_1071 (O_1071,N_9041,N_9552);
and UO_1072 (O_1072,N_9152,N_9289);
xnor UO_1073 (O_1073,N_9425,N_9094);
nand UO_1074 (O_1074,N_9051,N_9567);
or UO_1075 (O_1075,N_9881,N_9803);
or UO_1076 (O_1076,N_9066,N_9457);
nand UO_1077 (O_1077,N_9384,N_9359);
and UO_1078 (O_1078,N_9781,N_9061);
and UO_1079 (O_1079,N_9994,N_9876);
nand UO_1080 (O_1080,N_9426,N_9247);
or UO_1081 (O_1081,N_9043,N_9700);
or UO_1082 (O_1082,N_9660,N_9121);
nor UO_1083 (O_1083,N_9798,N_9513);
nand UO_1084 (O_1084,N_9258,N_9339);
nor UO_1085 (O_1085,N_9178,N_9614);
and UO_1086 (O_1086,N_9260,N_9776);
or UO_1087 (O_1087,N_9956,N_9655);
or UO_1088 (O_1088,N_9822,N_9689);
nand UO_1089 (O_1089,N_9527,N_9109);
and UO_1090 (O_1090,N_9847,N_9521);
xor UO_1091 (O_1091,N_9143,N_9572);
and UO_1092 (O_1092,N_9173,N_9702);
or UO_1093 (O_1093,N_9994,N_9495);
nand UO_1094 (O_1094,N_9583,N_9633);
or UO_1095 (O_1095,N_9321,N_9586);
nor UO_1096 (O_1096,N_9142,N_9028);
and UO_1097 (O_1097,N_9145,N_9827);
and UO_1098 (O_1098,N_9616,N_9432);
xnor UO_1099 (O_1099,N_9866,N_9920);
nor UO_1100 (O_1100,N_9536,N_9979);
nand UO_1101 (O_1101,N_9684,N_9459);
xor UO_1102 (O_1102,N_9072,N_9471);
or UO_1103 (O_1103,N_9785,N_9049);
nand UO_1104 (O_1104,N_9999,N_9401);
xor UO_1105 (O_1105,N_9676,N_9371);
and UO_1106 (O_1106,N_9469,N_9998);
and UO_1107 (O_1107,N_9776,N_9179);
or UO_1108 (O_1108,N_9204,N_9130);
nor UO_1109 (O_1109,N_9544,N_9306);
xor UO_1110 (O_1110,N_9952,N_9493);
xnor UO_1111 (O_1111,N_9765,N_9390);
and UO_1112 (O_1112,N_9411,N_9254);
xnor UO_1113 (O_1113,N_9387,N_9423);
and UO_1114 (O_1114,N_9719,N_9393);
xnor UO_1115 (O_1115,N_9831,N_9906);
or UO_1116 (O_1116,N_9897,N_9889);
xnor UO_1117 (O_1117,N_9922,N_9584);
nor UO_1118 (O_1118,N_9408,N_9613);
xor UO_1119 (O_1119,N_9822,N_9064);
nand UO_1120 (O_1120,N_9903,N_9040);
xnor UO_1121 (O_1121,N_9976,N_9656);
and UO_1122 (O_1122,N_9308,N_9408);
or UO_1123 (O_1123,N_9060,N_9487);
xnor UO_1124 (O_1124,N_9991,N_9046);
xor UO_1125 (O_1125,N_9992,N_9764);
xnor UO_1126 (O_1126,N_9409,N_9893);
and UO_1127 (O_1127,N_9486,N_9499);
nor UO_1128 (O_1128,N_9672,N_9384);
or UO_1129 (O_1129,N_9542,N_9766);
and UO_1130 (O_1130,N_9291,N_9613);
nand UO_1131 (O_1131,N_9957,N_9850);
nor UO_1132 (O_1132,N_9317,N_9852);
or UO_1133 (O_1133,N_9831,N_9229);
and UO_1134 (O_1134,N_9662,N_9484);
or UO_1135 (O_1135,N_9041,N_9307);
xnor UO_1136 (O_1136,N_9586,N_9244);
or UO_1137 (O_1137,N_9358,N_9306);
or UO_1138 (O_1138,N_9681,N_9971);
or UO_1139 (O_1139,N_9853,N_9976);
nor UO_1140 (O_1140,N_9720,N_9744);
xnor UO_1141 (O_1141,N_9308,N_9183);
nand UO_1142 (O_1142,N_9420,N_9644);
or UO_1143 (O_1143,N_9706,N_9957);
or UO_1144 (O_1144,N_9137,N_9722);
nand UO_1145 (O_1145,N_9736,N_9860);
nor UO_1146 (O_1146,N_9397,N_9964);
and UO_1147 (O_1147,N_9237,N_9342);
nor UO_1148 (O_1148,N_9608,N_9883);
xnor UO_1149 (O_1149,N_9398,N_9740);
nand UO_1150 (O_1150,N_9217,N_9465);
nor UO_1151 (O_1151,N_9740,N_9439);
nor UO_1152 (O_1152,N_9886,N_9420);
nand UO_1153 (O_1153,N_9039,N_9541);
and UO_1154 (O_1154,N_9355,N_9602);
nand UO_1155 (O_1155,N_9886,N_9015);
nand UO_1156 (O_1156,N_9601,N_9420);
and UO_1157 (O_1157,N_9797,N_9766);
xor UO_1158 (O_1158,N_9289,N_9940);
and UO_1159 (O_1159,N_9377,N_9468);
or UO_1160 (O_1160,N_9157,N_9012);
and UO_1161 (O_1161,N_9901,N_9161);
or UO_1162 (O_1162,N_9339,N_9107);
or UO_1163 (O_1163,N_9620,N_9175);
or UO_1164 (O_1164,N_9604,N_9420);
nand UO_1165 (O_1165,N_9693,N_9138);
and UO_1166 (O_1166,N_9699,N_9308);
nor UO_1167 (O_1167,N_9999,N_9454);
and UO_1168 (O_1168,N_9046,N_9625);
and UO_1169 (O_1169,N_9627,N_9235);
and UO_1170 (O_1170,N_9853,N_9007);
nand UO_1171 (O_1171,N_9380,N_9764);
xnor UO_1172 (O_1172,N_9336,N_9351);
and UO_1173 (O_1173,N_9948,N_9863);
nand UO_1174 (O_1174,N_9680,N_9609);
nor UO_1175 (O_1175,N_9497,N_9650);
xor UO_1176 (O_1176,N_9831,N_9466);
or UO_1177 (O_1177,N_9830,N_9399);
nor UO_1178 (O_1178,N_9646,N_9192);
nor UO_1179 (O_1179,N_9306,N_9709);
xor UO_1180 (O_1180,N_9141,N_9614);
xor UO_1181 (O_1181,N_9182,N_9621);
nor UO_1182 (O_1182,N_9368,N_9451);
and UO_1183 (O_1183,N_9290,N_9285);
nor UO_1184 (O_1184,N_9450,N_9481);
xor UO_1185 (O_1185,N_9098,N_9834);
or UO_1186 (O_1186,N_9626,N_9055);
or UO_1187 (O_1187,N_9412,N_9236);
and UO_1188 (O_1188,N_9212,N_9125);
or UO_1189 (O_1189,N_9383,N_9539);
xor UO_1190 (O_1190,N_9221,N_9819);
nand UO_1191 (O_1191,N_9277,N_9044);
xnor UO_1192 (O_1192,N_9123,N_9317);
nor UO_1193 (O_1193,N_9654,N_9970);
nor UO_1194 (O_1194,N_9249,N_9565);
or UO_1195 (O_1195,N_9718,N_9488);
xnor UO_1196 (O_1196,N_9962,N_9349);
and UO_1197 (O_1197,N_9826,N_9345);
or UO_1198 (O_1198,N_9382,N_9446);
nand UO_1199 (O_1199,N_9261,N_9857);
xnor UO_1200 (O_1200,N_9281,N_9194);
nor UO_1201 (O_1201,N_9085,N_9926);
and UO_1202 (O_1202,N_9827,N_9382);
or UO_1203 (O_1203,N_9107,N_9696);
nor UO_1204 (O_1204,N_9059,N_9566);
xnor UO_1205 (O_1205,N_9318,N_9965);
nor UO_1206 (O_1206,N_9788,N_9950);
nor UO_1207 (O_1207,N_9614,N_9459);
xor UO_1208 (O_1208,N_9175,N_9009);
nor UO_1209 (O_1209,N_9217,N_9708);
xor UO_1210 (O_1210,N_9406,N_9951);
nor UO_1211 (O_1211,N_9401,N_9073);
and UO_1212 (O_1212,N_9472,N_9651);
nor UO_1213 (O_1213,N_9238,N_9872);
nand UO_1214 (O_1214,N_9554,N_9018);
xor UO_1215 (O_1215,N_9901,N_9460);
or UO_1216 (O_1216,N_9075,N_9640);
nand UO_1217 (O_1217,N_9103,N_9361);
nand UO_1218 (O_1218,N_9278,N_9842);
xor UO_1219 (O_1219,N_9109,N_9919);
or UO_1220 (O_1220,N_9646,N_9067);
nor UO_1221 (O_1221,N_9431,N_9050);
or UO_1222 (O_1222,N_9882,N_9057);
xor UO_1223 (O_1223,N_9270,N_9979);
nand UO_1224 (O_1224,N_9046,N_9890);
nor UO_1225 (O_1225,N_9910,N_9107);
nand UO_1226 (O_1226,N_9420,N_9041);
or UO_1227 (O_1227,N_9622,N_9156);
and UO_1228 (O_1228,N_9680,N_9492);
nand UO_1229 (O_1229,N_9373,N_9384);
xor UO_1230 (O_1230,N_9422,N_9339);
nand UO_1231 (O_1231,N_9995,N_9867);
and UO_1232 (O_1232,N_9094,N_9412);
nor UO_1233 (O_1233,N_9080,N_9978);
xnor UO_1234 (O_1234,N_9054,N_9745);
nand UO_1235 (O_1235,N_9469,N_9163);
nand UO_1236 (O_1236,N_9125,N_9011);
nand UO_1237 (O_1237,N_9246,N_9384);
or UO_1238 (O_1238,N_9601,N_9253);
and UO_1239 (O_1239,N_9467,N_9626);
and UO_1240 (O_1240,N_9541,N_9599);
xor UO_1241 (O_1241,N_9248,N_9078);
or UO_1242 (O_1242,N_9195,N_9608);
nand UO_1243 (O_1243,N_9337,N_9169);
nand UO_1244 (O_1244,N_9040,N_9012);
nand UO_1245 (O_1245,N_9847,N_9246);
or UO_1246 (O_1246,N_9349,N_9628);
nor UO_1247 (O_1247,N_9557,N_9764);
xnor UO_1248 (O_1248,N_9602,N_9863);
and UO_1249 (O_1249,N_9088,N_9897);
xor UO_1250 (O_1250,N_9454,N_9535);
xnor UO_1251 (O_1251,N_9545,N_9142);
and UO_1252 (O_1252,N_9702,N_9978);
and UO_1253 (O_1253,N_9320,N_9115);
xor UO_1254 (O_1254,N_9126,N_9690);
nor UO_1255 (O_1255,N_9006,N_9283);
nor UO_1256 (O_1256,N_9729,N_9638);
nor UO_1257 (O_1257,N_9178,N_9445);
nor UO_1258 (O_1258,N_9928,N_9214);
nand UO_1259 (O_1259,N_9924,N_9727);
xor UO_1260 (O_1260,N_9119,N_9991);
nor UO_1261 (O_1261,N_9302,N_9555);
and UO_1262 (O_1262,N_9917,N_9128);
nor UO_1263 (O_1263,N_9985,N_9326);
xnor UO_1264 (O_1264,N_9433,N_9769);
nand UO_1265 (O_1265,N_9949,N_9427);
or UO_1266 (O_1266,N_9858,N_9687);
nand UO_1267 (O_1267,N_9142,N_9804);
and UO_1268 (O_1268,N_9938,N_9324);
nor UO_1269 (O_1269,N_9323,N_9014);
or UO_1270 (O_1270,N_9844,N_9707);
xor UO_1271 (O_1271,N_9373,N_9320);
nand UO_1272 (O_1272,N_9676,N_9165);
nand UO_1273 (O_1273,N_9973,N_9944);
nor UO_1274 (O_1274,N_9762,N_9120);
or UO_1275 (O_1275,N_9230,N_9213);
nor UO_1276 (O_1276,N_9333,N_9593);
xnor UO_1277 (O_1277,N_9598,N_9385);
nor UO_1278 (O_1278,N_9974,N_9867);
nor UO_1279 (O_1279,N_9567,N_9637);
nand UO_1280 (O_1280,N_9827,N_9868);
and UO_1281 (O_1281,N_9590,N_9423);
and UO_1282 (O_1282,N_9236,N_9445);
xor UO_1283 (O_1283,N_9027,N_9806);
nand UO_1284 (O_1284,N_9142,N_9789);
xor UO_1285 (O_1285,N_9741,N_9089);
nor UO_1286 (O_1286,N_9053,N_9854);
xor UO_1287 (O_1287,N_9982,N_9859);
nand UO_1288 (O_1288,N_9687,N_9178);
and UO_1289 (O_1289,N_9815,N_9556);
nand UO_1290 (O_1290,N_9004,N_9261);
nand UO_1291 (O_1291,N_9428,N_9322);
or UO_1292 (O_1292,N_9225,N_9529);
xnor UO_1293 (O_1293,N_9039,N_9139);
nand UO_1294 (O_1294,N_9459,N_9540);
nand UO_1295 (O_1295,N_9350,N_9509);
nand UO_1296 (O_1296,N_9732,N_9983);
and UO_1297 (O_1297,N_9530,N_9268);
xor UO_1298 (O_1298,N_9208,N_9320);
or UO_1299 (O_1299,N_9338,N_9193);
nand UO_1300 (O_1300,N_9505,N_9202);
xor UO_1301 (O_1301,N_9579,N_9077);
nor UO_1302 (O_1302,N_9315,N_9074);
nor UO_1303 (O_1303,N_9227,N_9314);
or UO_1304 (O_1304,N_9462,N_9411);
and UO_1305 (O_1305,N_9495,N_9748);
nand UO_1306 (O_1306,N_9685,N_9211);
nor UO_1307 (O_1307,N_9498,N_9671);
nor UO_1308 (O_1308,N_9897,N_9962);
nand UO_1309 (O_1309,N_9256,N_9307);
nand UO_1310 (O_1310,N_9942,N_9939);
and UO_1311 (O_1311,N_9157,N_9968);
nand UO_1312 (O_1312,N_9878,N_9861);
xnor UO_1313 (O_1313,N_9277,N_9501);
nand UO_1314 (O_1314,N_9085,N_9631);
and UO_1315 (O_1315,N_9023,N_9859);
or UO_1316 (O_1316,N_9175,N_9518);
nand UO_1317 (O_1317,N_9939,N_9996);
nand UO_1318 (O_1318,N_9439,N_9841);
xnor UO_1319 (O_1319,N_9255,N_9223);
or UO_1320 (O_1320,N_9899,N_9777);
nor UO_1321 (O_1321,N_9400,N_9390);
and UO_1322 (O_1322,N_9569,N_9832);
xnor UO_1323 (O_1323,N_9842,N_9444);
xor UO_1324 (O_1324,N_9967,N_9463);
xor UO_1325 (O_1325,N_9363,N_9921);
and UO_1326 (O_1326,N_9842,N_9600);
and UO_1327 (O_1327,N_9597,N_9449);
and UO_1328 (O_1328,N_9092,N_9422);
and UO_1329 (O_1329,N_9352,N_9362);
or UO_1330 (O_1330,N_9290,N_9491);
xor UO_1331 (O_1331,N_9365,N_9774);
nand UO_1332 (O_1332,N_9802,N_9486);
nor UO_1333 (O_1333,N_9557,N_9328);
or UO_1334 (O_1334,N_9313,N_9096);
or UO_1335 (O_1335,N_9960,N_9392);
or UO_1336 (O_1336,N_9643,N_9211);
or UO_1337 (O_1337,N_9654,N_9535);
xnor UO_1338 (O_1338,N_9938,N_9081);
xor UO_1339 (O_1339,N_9030,N_9793);
and UO_1340 (O_1340,N_9585,N_9332);
nor UO_1341 (O_1341,N_9493,N_9784);
xor UO_1342 (O_1342,N_9217,N_9387);
xnor UO_1343 (O_1343,N_9132,N_9919);
or UO_1344 (O_1344,N_9698,N_9055);
or UO_1345 (O_1345,N_9881,N_9954);
or UO_1346 (O_1346,N_9075,N_9071);
and UO_1347 (O_1347,N_9527,N_9061);
nor UO_1348 (O_1348,N_9521,N_9854);
nor UO_1349 (O_1349,N_9653,N_9555);
nand UO_1350 (O_1350,N_9617,N_9679);
and UO_1351 (O_1351,N_9347,N_9068);
nor UO_1352 (O_1352,N_9756,N_9906);
nand UO_1353 (O_1353,N_9823,N_9287);
xnor UO_1354 (O_1354,N_9752,N_9789);
or UO_1355 (O_1355,N_9828,N_9628);
xor UO_1356 (O_1356,N_9445,N_9141);
xor UO_1357 (O_1357,N_9157,N_9846);
nand UO_1358 (O_1358,N_9572,N_9846);
nor UO_1359 (O_1359,N_9770,N_9254);
nand UO_1360 (O_1360,N_9219,N_9124);
nand UO_1361 (O_1361,N_9781,N_9295);
nor UO_1362 (O_1362,N_9448,N_9034);
nand UO_1363 (O_1363,N_9560,N_9705);
or UO_1364 (O_1364,N_9420,N_9663);
nand UO_1365 (O_1365,N_9258,N_9156);
or UO_1366 (O_1366,N_9883,N_9645);
nor UO_1367 (O_1367,N_9239,N_9353);
nor UO_1368 (O_1368,N_9289,N_9196);
nand UO_1369 (O_1369,N_9148,N_9233);
xor UO_1370 (O_1370,N_9245,N_9819);
xnor UO_1371 (O_1371,N_9760,N_9732);
nand UO_1372 (O_1372,N_9476,N_9399);
or UO_1373 (O_1373,N_9508,N_9503);
nor UO_1374 (O_1374,N_9522,N_9122);
nor UO_1375 (O_1375,N_9762,N_9382);
nor UO_1376 (O_1376,N_9984,N_9459);
nor UO_1377 (O_1377,N_9403,N_9479);
and UO_1378 (O_1378,N_9834,N_9969);
and UO_1379 (O_1379,N_9150,N_9624);
xor UO_1380 (O_1380,N_9820,N_9765);
nor UO_1381 (O_1381,N_9811,N_9945);
xor UO_1382 (O_1382,N_9746,N_9504);
nor UO_1383 (O_1383,N_9075,N_9379);
xor UO_1384 (O_1384,N_9047,N_9763);
or UO_1385 (O_1385,N_9818,N_9109);
nand UO_1386 (O_1386,N_9043,N_9120);
and UO_1387 (O_1387,N_9037,N_9468);
nand UO_1388 (O_1388,N_9362,N_9962);
or UO_1389 (O_1389,N_9961,N_9077);
or UO_1390 (O_1390,N_9584,N_9944);
xnor UO_1391 (O_1391,N_9105,N_9352);
nor UO_1392 (O_1392,N_9957,N_9464);
and UO_1393 (O_1393,N_9663,N_9125);
and UO_1394 (O_1394,N_9452,N_9918);
nand UO_1395 (O_1395,N_9512,N_9610);
nor UO_1396 (O_1396,N_9358,N_9823);
nand UO_1397 (O_1397,N_9801,N_9587);
xor UO_1398 (O_1398,N_9560,N_9868);
nand UO_1399 (O_1399,N_9626,N_9545);
and UO_1400 (O_1400,N_9434,N_9192);
xnor UO_1401 (O_1401,N_9839,N_9378);
and UO_1402 (O_1402,N_9467,N_9264);
xor UO_1403 (O_1403,N_9242,N_9473);
nand UO_1404 (O_1404,N_9417,N_9099);
or UO_1405 (O_1405,N_9864,N_9957);
nand UO_1406 (O_1406,N_9162,N_9097);
nand UO_1407 (O_1407,N_9329,N_9305);
and UO_1408 (O_1408,N_9473,N_9803);
or UO_1409 (O_1409,N_9464,N_9836);
nor UO_1410 (O_1410,N_9986,N_9393);
xnor UO_1411 (O_1411,N_9355,N_9238);
and UO_1412 (O_1412,N_9299,N_9681);
or UO_1413 (O_1413,N_9763,N_9218);
and UO_1414 (O_1414,N_9258,N_9295);
xnor UO_1415 (O_1415,N_9021,N_9054);
and UO_1416 (O_1416,N_9262,N_9220);
or UO_1417 (O_1417,N_9725,N_9959);
nand UO_1418 (O_1418,N_9992,N_9305);
or UO_1419 (O_1419,N_9681,N_9753);
xnor UO_1420 (O_1420,N_9557,N_9864);
nor UO_1421 (O_1421,N_9977,N_9683);
and UO_1422 (O_1422,N_9001,N_9168);
nor UO_1423 (O_1423,N_9113,N_9298);
and UO_1424 (O_1424,N_9658,N_9283);
nor UO_1425 (O_1425,N_9451,N_9504);
nand UO_1426 (O_1426,N_9528,N_9078);
or UO_1427 (O_1427,N_9529,N_9983);
or UO_1428 (O_1428,N_9717,N_9584);
or UO_1429 (O_1429,N_9759,N_9593);
or UO_1430 (O_1430,N_9832,N_9349);
nor UO_1431 (O_1431,N_9992,N_9280);
and UO_1432 (O_1432,N_9560,N_9251);
or UO_1433 (O_1433,N_9052,N_9572);
or UO_1434 (O_1434,N_9162,N_9140);
nand UO_1435 (O_1435,N_9754,N_9249);
nor UO_1436 (O_1436,N_9647,N_9016);
and UO_1437 (O_1437,N_9855,N_9383);
nor UO_1438 (O_1438,N_9340,N_9837);
nand UO_1439 (O_1439,N_9707,N_9475);
and UO_1440 (O_1440,N_9245,N_9267);
nor UO_1441 (O_1441,N_9914,N_9893);
nand UO_1442 (O_1442,N_9714,N_9378);
nand UO_1443 (O_1443,N_9967,N_9906);
and UO_1444 (O_1444,N_9137,N_9968);
nor UO_1445 (O_1445,N_9496,N_9480);
xnor UO_1446 (O_1446,N_9535,N_9126);
xor UO_1447 (O_1447,N_9716,N_9206);
or UO_1448 (O_1448,N_9776,N_9626);
or UO_1449 (O_1449,N_9030,N_9471);
xnor UO_1450 (O_1450,N_9776,N_9258);
or UO_1451 (O_1451,N_9122,N_9095);
nor UO_1452 (O_1452,N_9761,N_9604);
nand UO_1453 (O_1453,N_9094,N_9940);
or UO_1454 (O_1454,N_9788,N_9387);
or UO_1455 (O_1455,N_9435,N_9083);
or UO_1456 (O_1456,N_9332,N_9708);
nand UO_1457 (O_1457,N_9580,N_9198);
and UO_1458 (O_1458,N_9181,N_9755);
nand UO_1459 (O_1459,N_9095,N_9910);
nor UO_1460 (O_1460,N_9020,N_9213);
or UO_1461 (O_1461,N_9183,N_9110);
or UO_1462 (O_1462,N_9784,N_9401);
nor UO_1463 (O_1463,N_9333,N_9288);
or UO_1464 (O_1464,N_9894,N_9537);
nor UO_1465 (O_1465,N_9828,N_9697);
and UO_1466 (O_1466,N_9737,N_9681);
nand UO_1467 (O_1467,N_9112,N_9016);
xor UO_1468 (O_1468,N_9749,N_9330);
and UO_1469 (O_1469,N_9856,N_9727);
and UO_1470 (O_1470,N_9609,N_9014);
nand UO_1471 (O_1471,N_9879,N_9311);
xnor UO_1472 (O_1472,N_9500,N_9318);
and UO_1473 (O_1473,N_9562,N_9339);
nor UO_1474 (O_1474,N_9011,N_9003);
xnor UO_1475 (O_1475,N_9137,N_9704);
nor UO_1476 (O_1476,N_9832,N_9116);
nor UO_1477 (O_1477,N_9612,N_9321);
or UO_1478 (O_1478,N_9965,N_9269);
nor UO_1479 (O_1479,N_9402,N_9374);
and UO_1480 (O_1480,N_9244,N_9663);
xnor UO_1481 (O_1481,N_9454,N_9689);
or UO_1482 (O_1482,N_9292,N_9967);
and UO_1483 (O_1483,N_9131,N_9150);
or UO_1484 (O_1484,N_9928,N_9564);
nor UO_1485 (O_1485,N_9599,N_9772);
nor UO_1486 (O_1486,N_9639,N_9879);
nand UO_1487 (O_1487,N_9157,N_9881);
nand UO_1488 (O_1488,N_9013,N_9481);
xor UO_1489 (O_1489,N_9389,N_9870);
nand UO_1490 (O_1490,N_9751,N_9364);
or UO_1491 (O_1491,N_9864,N_9399);
nor UO_1492 (O_1492,N_9913,N_9104);
or UO_1493 (O_1493,N_9176,N_9801);
xor UO_1494 (O_1494,N_9145,N_9426);
nor UO_1495 (O_1495,N_9840,N_9596);
or UO_1496 (O_1496,N_9806,N_9086);
xnor UO_1497 (O_1497,N_9593,N_9168);
xor UO_1498 (O_1498,N_9523,N_9177);
and UO_1499 (O_1499,N_9105,N_9858);
endmodule